
module biu32_axi(rstn, clk, write_req, write_ack, write_data, write_sz, write_msk
		, read_req, read_ack, read_data, read_sz, Daddr, code_req, code_ack
		, code_data, code_addr, code_wreq, code_wack, code_wdata, readio_req
		, writeio_req, readio_ack, writeio_ack, writeio_data, readio_data
		, io_add, axi_AW, axi_AWVALID, axi_AWREADY, axi_AWBURST, axi_AWLEN
		, axi_AWSIZE, axi_W, axi_WVALID, axi_WREADY, axi_WSTRB, axi_WLAST
		, axi_AR, axi_ARVALID, axi_ARREADY, axi_ARBURST, axi_ARLEN, axi_ARSIZE
		, axi_R, axi_RVALID, axi_RREADY, axi_RLAST, axi_io_AW, axi_io_AWVALID
		, axi_io_AWREADY, axi_io_AWBURST, axi_io_AWLEN, axi_io_AWSIZE, axi_io_W
		, axi_io_WVALID, axi_io_WREADY, axi_io_WSTRB, axi_io_WLAST, axi_io_AR
		, axi_io_ARVALID, axi_io_ARREADY, axi_io_ARBURST, axi_io_ARLEN, axi_io_ARSIZE
		, axi_io_R, axi_io_RVALID, axi_io_RREADY, axi_io_RLAST, busy, outstanding
		);

	input rstn;
	input clk;
	input write_req;
	output write_ack;
	input [31:0] write_data;
	input [1:0] write_sz;
	input [3:0] write_msk;
	input read_req;
	output read_ack;
	output [31:0] read_data;
	input [1:0] read_sz;
	input [31:0] Daddr;
	input code_req;
	output code_ack;
	output [127:0] code_data;
	input [31:0] code_addr;
	input code_wreq;
	output code_wack;
	input [31:0] code_wdata;
	input readio_req;
	input writeio_req;
	output readio_ack;
	output writeio_ack;
	input [31:0] writeio_data;
	output [31:0] readio_data;
	input [31:0] io_add;
	output [31:0] axi_AW;
	output axi_AWVALID;
	input axi_AWREADY;
	output [1:0] axi_AWBURST;
	output [7:0] axi_AWLEN;
	output [2:0] axi_AWSIZE;
	output [31:0] axi_W;
	output axi_WVALID;
	input axi_WREADY;
	output [3:0] axi_WSTRB;
	output axi_WLAST;
	output [31:0] axi_AR;
	output axi_ARVALID;
	input axi_ARREADY;
	output [1:0] axi_ARBURST;
	output [7:0] axi_ARLEN;
	output [2:0] axi_ARSIZE;
	input [31:0] axi_R;
	input axi_RVALID;
	output axi_RREADY;
	input axi_RLAST;
	output [31:0] axi_io_AW;
	output axi_io_AWVALID;
	input axi_io_AWREADY;
	output [1:0] axi_io_AWBURST;
	output [7:0] axi_io_AWLEN;
	output [2:0] axi_io_AWSIZE;
	output [31:0] axi_io_W;
	output axi_io_WVALID;
	input axi_io_WREADY;
	output [3:0] axi_io_WSTRB;
	output axi_io_WLAST;
	output [31:0] axi_io_AR;
	output axi_io_ARVALID;
	input axi_io_ARREADY;
	output [1:0] axi_io_ARBURST;
	output [7:0] axi_io_ARLEN;
	output [2:0] axi_io_ARSIZE;
	input [31:0] axi_io_R;
	input axi_io_RVALID;
	output axi_io_RREADY;
	input axi_io_RLAST;
	output busy;
	input outstanding;

	wire [1:0] A4;
	wire [4:0] fsm;
	wire [4:0] burst_idx;
	wire [9:0] cacheA;
	wire [149:0] cacheQ;
	wire [149:0] cacheD;
	wire [15:0] cacheM;



	notech_inv i_15669(.A(n_62423), .Z(n_62424));
	notech_inv i_15668(.A(n_62416), .Z(n_62423));
	notech_inv i_15667(.A(n_62421), .Z(n_62422));
	notech_inv i_15666(.A(n_62408), .Z(n_62421));
	notech_inv i_15665(.A(n_62419), .Z(n_62420));
	notech_inv i_15664(.A(n_62404), .Z(n_62419));
	notech_inv i_15663(.A(n_62417), .Z(n_62418));
	notech_inv i_15662(.A(n_62402), .Z(n_62417));
	notech_inv i_15661(.A(n_62415), .Z(n_62416));
	notech_inv i_15660(.A(n_62400), .Z(n_62415));
	notech_inv i_15659(.A(n_62413), .Z(n_62414));
	notech_inv i_15658(.A(n_62392), .Z(n_62413));
	notech_inv i_15657(.A(n_62411), .Z(n_62412));
	notech_inv i_15656(.A(n_62390), .Z(n_62411));
	notech_inv i_15655(.A(n_62409), .Z(n_62410));
	notech_inv i_15654(.A(n_62388), .Z(n_62409));
	notech_inv i_15653(.A(n_62407), .Z(n_62408));
	notech_inv i_15652(.A(n_62386), .Z(n_62407));
	notech_inv i_15651(.A(n_62405), .Z(n_62406));
	notech_inv i_15650(.A(n_62384), .Z(n_62405));
	notech_inv i_15649(.A(n_62403), .Z(n_62404));
	notech_inv i_15648(.A(n_62382), .Z(n_62403));
	notech_inv i_15647(.A(n_62401), .Z(n_62402));
	notech_inv i_15646(.A(n_62380), .Z(n_62401));
	notech_inv i_15645(.A(n_62399), .Z(n_62400));
	notech_inv i_15644(.A(n_62418), .Z(n_62399));
	notech_inv i_15643(.A(n_62397), .Z(n_62398));
	notech_inv i_15642(.A(n_62374), .Z(n_62397));
	notech_inv i_15641(.A(n_62395), .Z(n_62396));
	notech_inv i_15640(.A(n_62370), .Z(n_62395));
	notech_inv i_15639(.A(n_62393), .Z(n_62394));
	notech_inv i_15638(.A(n_62368), .Z(n_62393));
	notech_inv i_15637(.A(n_62391), .Z(n_62392));
	notech_inv i_15636(.A(n_62394), .Z(n_62391));
	notech_inv i_15635(.A(n_62389), .Z(n_62390));
	notech_inv i_15634(.A(n_62364), .Z(n_62389));
	notech_inv i_15633(.A(n_62387), .Z(n_62388));
	notech_inv i_15632(.A(n_62362), .Z(n_62387));
	notech_inv i_15631(.A(n_62385), .Z(n_62386));
	notech_inv i_15630(.A(n_62410), .Z(n_62385));
	notech_inv i_15629(.A(n_62383), .Z(n_62384));
	notech_inv i_15628(.A(n_62360), .Z(n_62383));
	notech_inv i_15627(.A(n_62381), .Z(n_62382));
	notech_inv i_15626(.A(n_62406), .Z(n_62381));
	notech_inv i_15625(.A(n_62379), .Z(n_62380));
	notech_inv i_15624(.A(n_62420), .Z(n_62379));
	notech_inv i_15623(.A(n_62377), .Z(n_62378));
	notech_inv i_15622(.A(n_62356), .Z(n_62377));
	notech_inv i_15621(.A(n_62375), .Z(n_62376));
	notech_inv i_15620(.A(n_62354), .Z(n_62375));
	notech_inv i_15619(.A(n_62373), .Z(n_62374));
	notech_inv i_15618(.A(n_62376), .Z(n_62373));
	notech_inv i_15617(.A(n_62371), .Z(n_62372));
	notech_inv i_15616(.A(n_62352), .Z(n_62371));
	notech_inv i_15615(.A(n_62369), .Z(n_62370));
	notech_inv i_15614(.A(n_62372), .Z(n_62369));
	notech_inv i_15613(.A(n_62367), .Z(n_62368));
	notech_inv i_15612(.A(n_62396), .Z(n_62367));
	notech_inv i_15611(.A(n_62365), .Z(n_62366));
	notech_inv i_15610(.A(n_62350), .Z(n_62365));
	notech_inv i_15609(.A(n_62363), .Z(n_62364));
	notech_inv i_15608(.A(n_62366), .Z(n_62363));
	notech_inv i_15607(.A(n_62361), .Z(n_62362));
	notech_inv i_15606(.A(n_62412), .Z(n_62361));
	notech_inv i_15605(.A(n_62359), .Z(n_62360));
	notech_inv i_15604(.A(n_62422), .Z(n_62359));
	notech_inv i_15603(.A(n_62357), .Z(n_62358));
	notech_inv i_15602(.A(clk), .Z(n_62357));
	notech_inv i_15601(.A(n_62355), .Z(n_62356));
	notech_inv i_15600(.A(n_62358), .Z(n_62355));
	notech_inv i_15599(.A(n_62353), .Z(n_62354));
	notech_inv i_15598(.A(n_62378), .Z(n_62353));
	notech_inv i_15597(.A(n_62351), .Z(n_62352));
	notech_inv i_15596(.A(n_62398), .Z(n_62351));
	notech_inv i_15595(.A(n_62349), .Z(n_62350));
	notech_inv i_15594(.A(n_62414), .Z(n_62349));
	notech_inv i_15213(.A(n_61967), .Z(n_61972));
	notech_inv i_15209(.A(n_61967), .Z(n_61968));
	notech_inv i_15208(.A(n_1996), .Z(n_61967));
	notech_inv i_15201(.A(n_61958), .Z(n_61959));
	notech_inv i_15200(.A(n_967), .Z(n_61958));
	notech_inv i_14834(.A(n_61881), .Z(n_61895));
	notech_inv i_14833(.A(n_61881), .Z(n_61894));
	notech_inv i_14827(.A(n_61881), .Z(n_61888));
	notech_inv i_14821(.A(n_61881), .Z(n_61882));
	notech_inv i_14820(.A(n_2008), .Z(n_61881));
	notech_inv i_14813(.A(n_61872), .Z(n_61873));
	notech_inv i_14812(.A(n_28023), .Z(n_61872));
	notech_inv i_14809(.A(n_61856), .Z(n_61868));
	notech_inv i_14808(.A(n_61856), .Z(n_61867));
	notech_inv i_14803(.A(n_61856), .Z(n_61862));
	notech_inv i_14798(.A(n_61856), .Z(n_61857));
	notech_inv i_14797(.A(n_970), .Z(n_61856));
	notech_inv i_14771(.A(n_61820), .Z(n_61826));
	notech_inv i_14770(.A(n_61820), .Z(n_61825));
	notech_inv i_14766(.A(n_61820), .Z(n_61821));
	notech_inv i_14765(.A(n_2003), .Z(n_61820));
	notech_inv i_14764(.A(n_61798), .Z(n_61818));
	notech_inv i_14763(.A(n_61798), .Z(n_61817));
	notech_inv i_14762(.A(n_61798), .Z(n_61816));
	notech_inv i_14761(.A(n_61798), .Z(n_61815));
	notech_inv i_14760(.A(n_61798), .Z(n_61814));
	notech_inv i_14759(.A(n_61798), .Z(n_61813));
	notech_inv i_14757(.A(n_61798), .Z(n_61811));
	notech_inv i_14756(.A(n_61798), .Z(n_61810));
	notech_inv i_14755(.A(n_61798), .Z(n_61809));
	notech_inv i_14754(.A(n_61798), .Z(n_61808));
	notech_inv i_14753(.A(n_61798), .Z(n_61807));
	notech_inv i_14752(.A(n_61798), .Z(n_61806));
	notech_inv i_14750(.A(n_61798), .Z(n_61804));
	notech_inv i_14749(.A(n_61798), .Z(n_61803));
	notech_inv i_14748(.A(n_61798), .Z(n_61802));
	notech_inv i_14747(.A(n_61798), .Z(n_61801));
	notech_inv i_14746(.A(n_61798), .Z(n_61800));
	notech_inv i_14745(.A(n_61798), .Z(n_61799));
	notech_inv i_14744(.A(rstn), .Z(n_61798));
	notech_inv i_14208(.A(n_61256), .Z(n_61257));
	notech_inv i_14207(.A(n_2010), .Z(n_61256));
	notech_inv i_14198(.A(n_61245), .Z(n_61246));
	notech_inv i_14197(.A(n_1065), .Z(n_61245));
	notech_inv i_14190(.A(n_61236), .Z(n_61237));
	notech_inv i_14189(.A(n_1059), .Z(n_61236));
	notech_inv i_14182(.A(n_61223), .Z(n_61228));
	notech_inv i_14178(.A(n_61223), .Z(n_61224));
	notech_inv i_14177(.A(n_2024), .Z(n_61223));
	notech_inv i_14170(.A(n_61214), .Z(n_61215));
	notech_inv i_14169(.A(n_6629), .Z(n_61214));
	notech_inv i_14162(.A(n_61201), .Z(n_61206));
	notech_inv i_14158(.A(n_61201), .Z(n_61202));
	notech_inv i_14157(.A(\nbus_11686[0] ), .Z(n_61201));
	notech_inv i_13760(.A(n_60805), .Z(n_60807));
	notech_inv i_13759(.A(n_60805), .Z(code_data[0]));
	notech_inv i_13758(.A(\nbus_14527[0] ), .Z(n_60805));
	notech_inv i_12970(.A(n_59929), .Z(n_59930));
	notech_inv i_12969(.A(n_1277), .Z(n_59929));
	notech_inv i_12962(.A(n_59920), .Z(n_59921));
	notech_inv i_12961(.A(n_2071), .Z(n_59920));
	notech_inv i_12952(.A(n_59909), .Z(n_59910));
	notech_inv i_12951(.A(n_1375), .Z(n_59909));
	notech_inv i_12949(.A(n_59884), .Z(n_59906));
	notech_inv i_12947(.A(n_59884), .Z(n_59904));
	notech_inv i_12946(.A(n_59884), .Z(n_59903));
	notech_inv i_12942(.A(n_59884), .Z(n_59899));
	notech_inv i_12940(.A(n_59884), .Z(n_59897));
	notech_inv i_12937(.A(n_59884), .Z(n_59894));
	notech_inv i_12935(.A(n_59884), .Z(n_59892));
	notech_inv i_12934(.A(n_59884), .Z(n_59891));
	notech_inv i_12930(.A(n_59884), .Z(n_59887));
	notech_inv i_12928(.A(n_59884), .Z(n_59885));
	notech_inv i_12927(.A(A4[0]), .Z(n_59884));
	notech_inv i_12923(.A(n_59865), .Z(n_59879));
	notech_inv i_12922(.A(n_59865), .Z(n_59878));
	notech_inv i_12916(.A(n_59865), .Z(n_59872));
	notech_inv i_12910(.A(n_59865), .Z(n_59866));
	notech_inv i_12909(.A(n_2074), .Z(n_59865));
	notech_inv i_12905(.A(n_59846), .Z(n_59860));
	notech_inv i_12904(.A(n_59846), .Z(n_59859));
	notech_inv i_12898(.A(n_59846), .Z(n_59853));
	notech_inv i_12892(.A(n_59846), .Z(n_59847));
	notech_inv i_12891(.A(n_2076), .Z(n_59846));
	notech_inv i_12882(.A(n_59835), .Z(n_59836));
	notech_inv i_12881(.A(n_1377), .Z(n_59835));
	notech_inv i_12872(.A(n_59824), .Z(n_59825));
	notech_inv i_12871(.A(n_1474), .Z(n_59824));
	notech_inv i_12862(.A(n_59813), .Z(n_59814));
	notech_inv i_12861(.A(n_1476), .Z(n_59813));
	notech_inv i_12852(.A(n_59802), .Z(n_59803));
	notech_inv i_12851(.A(n_1573), .Z(n_59802));
	notech_inv i_12842(.A(n_59791), .Z(n_59792));
	notech_inv i_12841(.A(n_1575), .Z(n_59791));
	notech_inv i_12832(.A(n_59780), .Z(n_59781));
	notech_inv i_12831(.A(n_1703), .Z(n_59780));
	notech_inv i_12822(.A(n_59769), .Z(n_59770));
	notech_inv i_12821(.A(n_1705), .Z(n_59769));
	notech_inv i_10457(.A(n_57109), .Z(n_57110));
	notech_inv i_10456(.A(n_6743), .Z(n_57109));
	notech_inv i_8337(.A(n_54993), .Z(n_54994));
	notech_inv i_8336(.A(\nbus_11696[0] ), .Z(n_54993));
	notech_inv i_7910(.A(n_54523), .Z(n_54524));
	notech_inv i_7909(.A(n_6746), .Z(n_54523));
	notech_inv i_7900(.A(n_54512), .Z(n_54513));
	notech_inv i_7899(.A(n_6745), .Z(n_54512));
	notech_inv i_7890(.A(n_54501), .Z(n_54502));
	notech_inv i_7889(.A(n_6744), .Z(n_54501));
	notech_inv i_7800(.A(n_54368), .Z(n_54369));
	notech_inv i_7799(.A(n_2245), .Z(n_54368));
	notech_inv i_7790(.A(n_54357), .Z(n_54358));
	notech_inv i_7789(.A(n_224057077), .Z(n_54357));
	notech_inv i_7782(.A(n_54348), .Z(n_54349));
	notech_inv i_7781(.A(n_223857075), .Z(n_54348));
	notech_inv i_7772(.A(n_54293), .Z(n_54294));
	notech_inv i_7771(.A(n_224357080), .Z(n_54293));
	notech_ao4 i_57723(.A(n_1059), .B(n_6807), .C(n_2010), .D(n_6845), .Z(n_990
		));
	notech_ao4 i_57729(.A(n_1059), .B(n_6808), .C(n_2010), .D(n_6846), .Z(n_987
		));
	notech_ao4 i_57735(.A(n_1059), .B(n_6809), .C(n_2010), .D(n_6847), .Z(n_984
		));
	notech_ao4 i_57741(.A(n_1059), .B(n_6810), .C(n_2010), .D(n_6848), .Z(n_981
		));
	notech_ao4 i_57747(.A(n_1059), .B(n_6811), .C(n_2010), .D(n_6849), .Z(n_978
		));
	notech_and4 i_58879(.A(n_61894), .B(n_61825), .C(n_971), .D(n_974), .Z(n_975
		));
	notech_nand3 i_151(.A(axi_RVALID), .B(axi_RLAST), .C(n_27143), .Z(n_974)
		);
	notech_and4 i_59961(.A(n_61894), .B(n_61825), .C(n_971), .D(n_972), .Z(n_973
		));
	notech_nand2 i_148(.A(axi_WREADY), .B(n_29767), .Z(n_972));
	notech_and2 i_43(.A(n_1218), .B(n_2010), .Z(n_971));
	notech_and3 i_48(.A(n_967), .B(n_61894), .C(n_28023), .Z(n_970));
	notech_nor2 i_138(.A(code_ack), .B(n_6979), .Z(n_969));
	notech_or4 i_62(.A(fsm[1]), .B(fsm[3]), .C(n_6630), .D(fsm[2]), .Z(busy)
		);
	notech_and2 i_5(.A(n_1996), .B(n_6636), .Z(n_967));
	notech_xor2 i_133(.A(burst_idx[4]), .B(n_2028), .Z(n_966));
	notech_xor2 i_132(.A(burst_idx[3]), .B(n_2027), .Z(n_965));
	notech_xor2 i_131(.A(burst_idx[2]), .B(n_2026), .Z(n_964));
	notech_xor2 i_130(.A(burst_idx[1]), .B(burst_idx[0]), .Z(n_963));
	notech_nand2 i_128(.A(n_1218), .B(n_28023), .Z(n_962));
	notech_xor2 i_1880101(.A(axi_AR[14]), .B(cacheQ[128]), .Z(n_959));
	notech_xor2 i_1980102(.A(axi_AR[15]), .B(cacheQ[129]), .Z(n_958));
	notech_xor2 i_20(.A(axi_AR[16]), .B(cacheQ[130]), .Z(n_957));
	notech_xor2 i_2180103(.A(axi_AR[17]), .B(cacheQ[131]), .Z(n_956));
	notech_xor2 i_2280104(.A(axi_AR[18]), .B(cacheQ[132]), .Z(n_955));
	notech_xor2 i_2380105(.A(axi_AR[19]), .B(cacheQ[133]), .Z(n_954));
	notech_xor2 i_2480106(.A(axi_AR[20]), .B(cacheQ[134]), .Z(n_953));
	notech_xor2 i_2580107(.A(axi_AR[21]), .B(cacheQ[135]), .Z(n_952));
	notech_xor2 i_2680108(.A(axi_AR[22]), .B(cacheQ[136]), .Z(n_951));
	notech_xor2 i_2780109(.A(axi_AR[23]), .B(cacheQ[137]), .Z(n_950));
	notech_xor2 i_28(.A(axi_AR[24]), .B(cacheQ[138]), .Z(n_949));
	notech_xor2 i_2980110(.A(axi_AR[25]), .B(cacheQ[139]), .Z(n_948));
	notech_xor2 i_3080111(.A(axi_AR[26]), .B(cacheQ[140]), .Z(n_947));
	notech_xor2 i_3180112(.A(axi_AR[27]), .B(cacheQ[141]), .Z(n_946));
	notech_xor2 i_3280113(.A(axi_AR[28]), .B(cacheQ[142]), .Z(n_945));
	notech_xor2 i_3380114(.A(axi_AR[29]), .B(cacheQ[143]), .Z(n_944));
	notech_xor2 i_3480115(.A(axi_AR[30]), .B(cacheQ[144]), .Z(n_943));
	notech_xor2 i_3580116(.A(axi_AR[31]), .B(cacheQ[145]), .Z(n_942));
	notech_or4 i_4780126(.A(n_959), .B(n_958), .C(n_957), .D(n_956), .Z(n_933
		));
	notech_or4 i_4880127(.A(n_955), .B(n_954), .C(n_953), .D(n_952), .Z(n_932
		));
	notech_or4 i_4980128(.A(n_951), .B(n_950), .C(n_949), .D(n_948), .Z(n_931
		));
	notech_or4 i_5080129(.A(n_947), .B(n_946), .C(n_945), .D(n_944), .Z(n_930
		));
	notech_or4 i_5580132(.A(n_933), .B(n_932), .C(n_931), .D(n_930), .Z(n_927
		));
	notech_xor2 i_1880152(.A(cacheQ[128]), .B(axi_AW[14]), .Z(n_925));
	notech_xor2 i_1980153(.A(cacheQ[129]), .B(axi_AW[15]), .Z(n_924));
	notech_xor2 i_2080154(.A(cacheQ[130]), .B(axi_AW[16]), .Z(n_923));
	notech_xor2 i_2180155(.A(cacheQ[131]), .B(axi_AW[17]), .Z(n_922));
	notech_xor2 i_2280156(.A(cacheQ[132]), .B(axi_AW[18]), .Z(n_921));
	notech_xor2 i_2380157(.A(cacheQ[133]), .B(axi_AW[19]), .Z(n_920));
	notech_xor2 i_2480158(.A(cacheQ[134]), .B(axi_AW[20]), .Z(n_919));
	notech_xor2 i_2580159(.A(cacheQ[135]), .B(axi_AW[21]), .Z(n_918));
	notech_xor2 i_2680160(.A(cacheQ[136]), .B(axi_AW[22]), .Z(n_917));
	notech_xor2 i_2780161(.A(cacheQ[137]), .B(axi_AW[23]), .Z(n_916));
	notech_xor2 i_2880162(.A(cacheQ[138]), .B(axi_AW[24]), .Z(n_915));
	notech_xor2 i_2980163(.A(cacheQ[139]), .B(axi_AW[25]), .Z(n_914));
	notech_xor2 i_3080164(.A(cacheQ[140]), .B(axi_AW[26]), .Z(n_913));
	notech_xor2 i_3180165(.A(cacheQ[141]), .B(axi_AW[27]), .Z(n_912));
	notech_xor2 i_3280166(.A(cacheQ[142]), .B(axi_AW[28]), .Z(n_911));
	notech_xor2 i_3380167(.A(cacheQ[143]), .B(axi_AW[29]), .Z(n_910));
	notech_xor2 i_3480168(.A(n_6970), .B(axi_AW[30]), .Z(n_909));
	notech_xor2 i_3580169(.A(n_6971), .B(axi_AW[31]), .Z(n_908));
	notech_or4 i_4780179(.A(n_925), .B(n_924), .C(n_923), .D(n_922), .Z(n_899
		));
	notech_or4 i_4880180(.A(n_921), .B(n_920), .C(n_919), .D(n_918), .Z(n_898
		));
	notech_or4 i_4980181(.A(n_917), .B(n_916), .C(n_915), .D(n_914), .Z(n_897
		));
	notech_or4 i_5080182(.A(n_913), .B(n_912), .C(n_911), .D(n_910), .Z(n_896
		));
	notech_or4 i_5580185(.A(n_899), .B(n_898), .C(n_897), .D(n_896), .Z(n_893
		));
	notech_ao4 i_57717(.A(n_1059), .B(n_6806), .C(n_2010), .D(n_6844), .Z(n_993
		));
	notech_ao4 i_57711(.A(n_1059), .B(n_6805), .C(n_2010), .D(n_6843), .Z(n_996
		));
	notech_ao4 i_57705(.A(n_1059), .B(n_6804), .C(n_2010), .D(n_6842), .Z(n_999
		));
	notech_ao4 i_57699(.A(n_1059), .B(n_6803), .C(n_2010), .D(n_6841), .Z(n_1002
		));
	notech_ao4 i_57693(.A(n_1059), .B(n_6802), .C(n_2010), .D(n_6840), .Z(n_1005
		));
	notech_ao4 i_57687(.A(n_1059), .B(n_6801), .C(n_2010), .D(n_6839), .Z(n_1008
		));
	notech_ao4 i_57681(.A(n_1059), .B(n_6800), .C(n_2010), .D(n_6838), .Z(n_1011
		));
	notech_ao4 i_57675(.A(n_1059), .B(n_6799), .C(n_2010), .D(n_6837), .Z(n_1014
		));
	notech_ao4 i_57669(.A(n_1059), .B(n_6798), .C(n_2010), .D(n_6836), .Z(n_1017
		));
	notech_ao4 i_57663(.A(n_61237), .B(n_6797), .C(n_2010), .D(n_6835), .Z(n_1020
		));
	notech_ao4 i_57657(.A(n_61237), .B(n_6796), .C(n_2010), .D(n_6834), .Z(n_1023
		));
	notech_ao4 i_57651(.A(n_61237), .B(n_6795), .C(n_2010), .D(n_6833), .Z(n_1026
		));
	notech_ao4 i_57645(.A(n_61237), .B(n_6794), .C(n_61257), .D(n_6832), .Z(n_1029
		));
	notech_ao4 i_57639(.A(n_61237), .B(n_6784), .C(n_61257), .D(n_6831), .Z(n_1032
		));
	notech_ao4 i_57633(.A(n_61237), .B(n_6785), .C(n_61257), .D(n_6830), .Z(n_1035
		));
	notech_ao4 i_57627(.A(n_61237), .B(n_6786), .C(n_61257), .D(n_6829), .Z(n_1038
		));
	notech_ao4 i_57621(.A(n_61237), .B(n_6787), .C(n_61257), .D(n_6828), .Z(n_1041
		));
	notech_ao4 i_57615(.A(n_61237), .B(n_6788), .C(n_61257), .D(n_6827), .Z(n_1044
		));
	notech_ao4 i_57609(.A(n_1059), .B(n_6789), .C(n_61257), .D(n_6826), .Z(n_1047
		));
	notech_ao4 i_57603(.A(n_61237), .B(n_6790), .C(n_61257), .D(n_6825), .Z(n_1050
		));
	notech_ao4 i_57597(.A(n_61237), .B(n_6791), .C(n_61257), .D(n_6824), .Z(n_1053
		));
	notech_ao4 i_57591(.A(n_61237), .B(n_6792), .C(n_61257), .D(n_6823), .Z(n_1056
		));
	notech_and3 i_30(.A(n_967), .B(n_2020), .C(n_1218), .Z(n_1059));
	notech_ao4 i_57585(.A(n_61237), .B(n_6793), .C(n_61257), .D(n_6822), .Z(n_1060
		));
	notech_ao4 i_57579(.A(n_2021), .B(n_6783), .C(n_61257), .D(n_6821), .Z(n_1063
		));
	notech_or4 i_242(.A(n_2019), .B(n_2016), .C(axi_AR[31]), .D(n_6974), .Z(n_1064
		));
	notech_and4 i_59898(.A(n_1218), .B(n_61257), .C(n_967), .D(n_1064), .Z(n_1065
		));
	notech_ao4 i_57574(.A(n_2021), .B(n_6782), .C(n_61257), .D(n_6820), .Z(n_1068
		));
	notech_ao4 i_57898(.A(n_61894), .B(n_6849), .C(n_61826), .D(n_6811), .Z(n_1071
		));
	notech_ao4 i_57893(.A(n_61894), .B(n_6848), .C(n_61826), .D(n_6810), .Z(n_1074
		));
	notech_ao4 i_57888(.A(n_61894), .B(n_6847), .C(n_61826), .D(n_6809), .Z(n_1077
		));
	notech_ao4 i_57883(.A(n_61895), .B(n_6846), .C(n_61825), .D(n_6808), .Z(n_1080
		));
	notech_ao4 i_57878(.A(n_61894), .B(n_6845), .C(n_61825), .D(n_6807), .Z(n_1083
		));
	notech_ao4 i_57873(.A(n_61894), .B(n_6844), .C(n_61825), .D(n_6806), .Z(n_1086
		));
	notech_ao4 i_57868(.A(n_61894), .B(n_6843), .C(n_61825), .D(n_6805), .Z(n_1089
		));
	notech_ao4 i_57863(.A(n_61894), .B(n_6842), .C(n_61825), .D(n_6804), .Z(n_1092
		));
	notech_ao4 i_57858(.A(n_61894), .B(n_6841), .C(n_61826), .D(n_6803), .Z(n_1095
		));
	notech_ao4 i_57853(.A(n_61894), .B(n_6840), .C(n_61826), .D(n_6802), .Z(n_1098
		));
	notech_ao4 i_57848(.A(n_61894), .B(n_6839), .C(n_61826), .D(n_6801), .Z(n_1101
		));
	notech_ao4 i_57843(.A(n_61894), .B(n_6838), .C(n_61826), .D(n_6800), .Z(n_1104
		));
	notech_ao4 i_57838(.A(n_61894), .B(n_6837), .C(n_61826), .D(n_6799), .Z(n_1107
		));
	notech_ao4 i_57833(.A(n_61894), .B(n_6836), .C(n_61826), .D(n_6798), .Z(n_1110
		));
	notech_ao4 i_57828(.A(n_61894), .B(n_6835), .C(n_61826), .D(n_6797), .Z(n_1113
		));
	notech_ao4 i_57823(.A(n_61895), .B(n_6834), .C(n_61826), .D(n_6796), .Z(n_1116
		));
	notech_ao4 i_57818(.A(n_61895), .B(n_6833), .C(n_61826), .D(n_6795), .Z(n_1119
		));
	notech_ao4 i_57813(.A(n_61895), .B(n_6832), .C(n_61826), .D(n_6794), .Z(n_1122
		));
	notech_ao4 i_57808(.A(n_61895), .B(n_6831), .C(n_61826), .D(n_6784), .Z(n_1125
		));
	notech_ao4 i_57803(.A(n_61895), .B(n_6830), .C(n_61821), .D(n_6785), .Z(n_1128
		));
	notech_ao4 i_57798(.A(n_61895), .B(n_6829), .C(n_61821), .D(n_6786), .Z(n_1131
		));
	notech_ao4 i_57793(.A(n_61895), .B(n_6828), .C(n_61821), .D(n_6787), .Z(n_1134
		));
	notech_ao4 i_57788(.A(n_61895), .B(n_6827), .C(n_61821), .D(n_6788), .Z(n_1137
		));
	notech_ao4 i_57783(.A(n_61895), .B(n_6826), .C(n_61821), .D(n_6789), .Z(n_1140
		));
	notech_ao4 i_57778(.A(n_61895), .B(n_6825), .C(n_61821), .D(n_6790), .Z(n_1143
		));
	notech_ao4 i_57773(.A(n_61895), .B(n_6824), .C(n_61821), .D(n_6791), .Z(n_1146
		));
	notech_ao4 i_57768(.A(n_61895), .B(n_6823), .C(n_61821), .D(n_6792), .Z(n_1149
		));
	notech_ao4 i_57763(.A(n_61895), .B(n_6822), .C(n_61821), .D(n_6793), .Z(n_1152
		));
	notech_ao4 i_57758(.A(n_61895), .B(n_6821), .C(n_61821), .D(n_6783), .Z(n_1155
		));
	notech_ao4 i_57753(.A(n_61895), .B(n_6820), .C(n_61821), .D(n_6782), .Z(n_1158
		));
	notech_or2 i_345(.A(n_2032), .B(n_2040), .Z(n_1166));
	notech_and3 i_127(.A(n_28023), .B(n_1166), .C(n_971), .Z(n_1169));
	notech_ao4 i_60225(.A(n_1169), .B(n_6976), .C(n_2025), .D(n_2030), .Z(n_1170
		));
	notech_ao4 i_57903(.A(n_2025), .B(burst_idx[0]), .C(n_2017), .D(n_1998),
		 .Z(n_1172));
	notech_ao4 i_57963(.A(n_61895), .B(n_6819), .C(n_61825), .D(n_6857), .Z(n_1175
		));
	notech_ao4 i_57958(.A(n_61895), .B(n_6818), .C(n_61825), .D(n_6856), .Z(n_1178
		));
	notech_ao4 i_57953(.A(n_61895), .B(n_6817), .C(n_61825), .D(n_6855), .Z(n_1181
		));
	notech_ao4 i_57948(.A(n_61895), .B(n_6816), .C(n_61825), .D(n_6854), .Z(n_1184
		));
	notech_ao4 i_57943(.A(n_61882), .B(n_6815), .C(n_61825), .D(n_6853), .Z(n_1187
		));
	notech_ao4 i_57938(.A(n_61882), .B(n_6814), .C(n_61821), .D(n_6852), .Z(n_1190
		));
	notech_ao4 i_57933(.A(n_61882), .B(n_6813), .C(n_61821), .D(n_6851), .Z(n_1193
		));
	notech_ao4 i_57928(.A(n_61882), .B(n_6812), .C(n_61821), .D(n_6850), .Z(n_1196
		));
	notech_nand2 i_381(.A(axi_ARREADY), .B(n_6647), .Z(n_1201));
	notech_and4 i_59890(.A(n_967), .B(n_971), .C(n_2045), .D(n_1201), .Z(n_1202
		));
	notech_nand2 i_58067(.A(n_61257), .B(n_2046), .Z(n_1203));
	notech_and4 i_60389(.A(n_967), .B(n_2049), .C(n_28023), .D(n_971), .Z(n_1206
		));
	notech_nand2 i_58070(.A(n_6677), .B(n_6625), .Z(n_1207));
	notech_or4 i_392(.A(fsm[0]), .B(fsm[4]), .C(fsm[2]), .D(n_6634), .Z(n_1208
		));
	notech_nand3 i_394(.A(read_req), .B(n_2044), .C(n_2043), .Z(n_1210));
	notech_and4 i_59206(.A(n_61867), .B(n_971), .C(n_2054), .D(n_1210), .Z(n_1211
		));
	notech_or2 i_399(.A(abort), .B(n_6625), .Z(n_1212));
	notech_nand3 i_58073(.A(n_2020), .B(n_1208), .C(n_1212), .Z(n_1213));
	notech_and4 i_59148(.A(n_61882), .B(n_61825), .C(n_2032), .D(n_971), .Z(n_1214
		));
	notech_nand3 i_58084(.A(n_61257), .B(n_61888), .C(n_2061), .Z(n_1215));
	notech_and4 i_58082(.A(n_2064), .B(n_61888), .C(n_2059), .D(n_2025), .Z(n_1216
		));
	notech_nand2 i_58081(.A(n_1064), .B(n_2061), .Z(n_1217));
	notech_nao3 i_61(.A(read_req), .B(n_6978), .C(n_2004), .Z(n_1218));
	notech_nand3 i_58079(.A(n_1218), .B(n_2061), .C(n_1750), .Z(n_1219));
	notech_nand2 i_413(.A(axi_WREADY), .B(n_2058), .Z(n_1220));
	notech_and4 i_58889(.A(n_967), .B(n_61888), .C(n_1220), .D(n_28023), .Z(n_1221
		));
	notech_and4 i_59369(.A(n_61867), .B(n_2068), .C(n_2045), .D(n_1220), .Z(n_1222
		));
	notech_and4 i_58077(.A(n_2025), .B(n_2060), .C(n_28023), .D(n_971), .Z(n_1223
		));
	notech_nand2 i_58553(.A(n_2024), .B(n_2071), .Z(n_1224));
	notech_ao4 i_58547(.A(n_2024), .B(n_6811), .C(n_2071), .D(n_6971), .Z(n_1227
		));
	notech_ao4 i_58544(.A(n_61228), .B(n_6810), .C(n_2071), .D(n_6970), .Z(n_1230
		));
	notech_ao4 i_58541(.A(n_2024), .B(n_6809), .C(n_2071), .D(n_6969), .Z(n_1233
		));
	notech_ao4 i_58538(.A(n_2024), .B(n_6808), .C(n_2071), .D(n_6968), .Z(n_1236
		));
	notech_ao4 i_58535(.A(n_2024), .B(n_6807), .C(n_2071), .D(n_6967), .Z(n_1239
		));
	notech_ao4 i_58532(.A(n_61228), .B(n_6806), .C(n_2071), .D(n_6966), .Z(n_1242
		));
	notech_ao4 i_58529(.A(n_61228), .B(n_6805), .C(n_2071), .D(n_6965), .Z(n_1245
		));
	notech_ao4 i_58526(.A(n_61228), .B(n_6804), .C(n_2071), .D(n_6964), .Z(n_1248
		));
	notech_ao4 i_58523(.A(n_61228), .B(n_6803), .C(n_2071), .D(n_6963), .Z(n_1251
		));
	notech_ao4 i_58520(.A(n_61228), .B(n_6802), .C(n_2071), .D(n_6962), .Z(n_1254
		));
	notech_ao4 i_58517(.A(n_61228), .B(n_6801), .C(n_59921), .D(n_6961), .Z(n_1257
		));
	notech_ao4 i_58514(.A(n_61228), .B(n_6800), .C(n_59921), .D(n_6960), .Z(n_1260
		));
	notech_ao4 i_58511(.A(n_2024), .B(n_6799), .C(n_59921), .D(n_6959), .Z(n_1263
		));
	notech_ao4 i_58508(.A(n_2024), .B(n_6798), .C(n_59921), .D(n_6958), .Z(n_1266
		));
	notech_ao4 i_58505(.A(n_2024), .B(n_6797), .C(n_59921), .D(n_6957), .Z(n_1269
		));
	notech_ao4 i_58502(.A(n_2024), .B(n_6796), .C(n_59921), .D(n_6956), .Z(n_1272
		));
	notech_ao4 i_58499(.A(n_2024), .B(n_6795), .C(n_59921), .D(n_6955), .Z(n_1275
		));
	notech_ao4 i_58979(.A(n_2073), .B(n_6983), .C(n_2072), .D(n_6976), .Z(n_1277
		));
	notech_ao4 i_58496(.A(n_2024), .B(n_6794), .C(n_2071), .D(n_6954), .Z(n_1280
		));
	notech_nand2 i_480(.A(cacheQ[127]), .B(n_1377), .Z(n_1281));
	notech_nand3 i_479(.A(n_59899), .B(n_59878), .C(axi_W[31]), .Z(n_1282)
		);
	notech_nao3 i_58493(.A(n_1282), .B(n_1281), .C(n_1579), .Z(n_1283));
	notech_nand2 i_484(.A(n_1377), .B(cacheQ[126]), .Z(n_1284));
	notech_nand3 i_483(.A(n_59899), .B(n_59878), .C(axi_W[30]), .Z(n_1285)
		);
	notech_nao3 i_58490(.A(n_1285), .B(n_1284), .C(n_1583), .Z(n_1286));
	notech_nand2 i_488(.A(n_1377), .B(cacheQ[125]), .Z(n_1287));
	notech_nand3 i_487(.A(n_59899), .B(n_59878), .C(axi_W[29]), .Z(n_1288)
		);
	notech_nao3 i_58487(.A(n_1288), .B(n_1287), .C(n_1587), .Z(n_1289));
	notech_nand2 i_492(.A(n_1377), .B(cacheQ[124]), .Z(n_1290));
	notech_nand3 i_491(.A(n_59899), .B(n_59878), .C(axi_W[28]), .Z(n_1291)
		);
	notech_nao3 i_58484(.A(n_1291), .B(n_1290), .C(n_1591), .Z(n_1292));
	notech_nand2 i_496(.A(n_1377), .B(cacheQ[123]), .Z(n_1293));
	notech_nand3 i_495(.A(n_59899), .B(n_59878), .C(axi_W[27]), .Z(n_1294)
		);
	notech_nao3 i_58481(.A(n_1294), .B(n_1293), .C(n_1595), .Z(n_1295));
	notech_nand2 i_500(.A(n_1377), .B(cacheQ[122]), .Z(n_1296));
	notech_nand3 i_499(.A(n_59899), .B(n_59879), .C(axi_W[26]), .Z(n_1297)
		);
	notech_nao3 i_58478(.A(n_1297), .B(n_1296), .C(n_1599), .Z(n_1298));
	notech_nand2 i_504(.A(n_1377), .B(cacheQ[121]), .Z(n_1299));
	notech_nand3 i_503(.A(n_59899), .B(n_59879), .C(axi_W[25]), .Z(n_1300)
		);
	notech_nao3 i_58475(.A(n_1300), .B(n_1299), .C(n_1603), .Z(n_1301));
	notech_nand2 i_508(.A(n_1377), .B(cacheQ[120]), .Z(n_1302));
	notech_nand3 i_507(.A(n_59899), .B(n_59878), .C(axi_W[24]), .Z(n_1303)
		);
	notech_nao3 i_58472(.A(n_1303), .B(n_1302), .C(n_1607), .Z(n_1304));
	notech_nand2 i_512(.A(n_1377), .B(cacheQ[119]), .Z(n_1305));
	notech_nand3 i_511(.A(n_59899), .B(n_59878), .C(axi_W[23]), .Z(n_1306)
		);
	notech_nao3 i_58469(.A(n_1306), .B(n_1305), .C(n_1611), .Z(n_1307));
	notech_nand2 i_516(.A(n_1377), .B(cacheQ[118]), .Z(n_1308));
	notech_nand3 i_515(.A(n_59903), .B(n_59878), .C(axi_W[22]), .Z(n_1309)
		);
	notech_nao3 i_58466(.A(n_1309), .B(n_1308), .C(n_1615), .Z(n_1310));
	notech_nand2 i_520(.A(n_1377), .B(cacheQ[117]), .Z(n_1311));
	notech_nand3 i_519(.A(n_59903), .B(n_59878), .C(axi_W[21]), .Z(n_1312)
		);
	notech_nao3 i_58463(.A(n_1312), .B(n_1311), .C(n_1619), .Z(n_1313));
	notech_nand2 i_524(.A(n_1377), .B(cacheQ[116]), .Z(n_1314));
	notech_nand3 i_523(.A(n_59903), .B(n_59878), .C(axi_W[20]), .Z(n_1315)
		);
	notech_nao3 i_58460(.A(n_1315), .B(n_1314), .C(n_1623), .Z(n_1316));
	notech_nand2 i_528(.A(n_1377), .B(cacheQ[115]), .Z(n_1317));
	notech_nand3 i_527(.A(n_59903), .B(n_59878), .C(axi_W[19]), .Z(n_1318)
		);
	notech_nao3 i_58457(.A(n_1318), .B(n_1317), .C(n_1627), .Z(n_1319));
	notech_nand2 i_532(.A(n_1377), .B(cacheQ[114]), .Z(n_1320));
	notech_nand3 i_531(.A(n_59903), .B(n_59878), .C(axi_W[18]), .Z(n_1321)
		);
	notech_nao3 i_58454(.A(n_1321), .B(n_1320), .C(n_1631), .Z(n_1322));
	notech_nand2 i_536(.A(n_1377), .B(cacheQ[113]), .Z(n_1323));
	notech_nand3 i_535(.A(n_59903), .B(n_59878), .C(axi_W[17]), .Z(n_1324)
		);
	notech_nao3 i_58451(.A(n_1324), .B(n_1323), .C(n_1635), .Z(n_1325));
	notech_nand2 i_540(.A(n_1377), .B(cacheQ[112]), .Z(n_1326));
	notech_nand3 i_539(.A(n_59903), .B(n_59878), .C(axi_W[16]), .Z(n_1327)
		);
	notech_nao3 i_58448(.A(n_1327), .B(n_1326), .C(n_1639), .Z(n_1328));
	notech_nand2 i_544(.A(n_59836), .B(cacheQ[111]), .Z(n_1329));
	notech_nand3 i_543(.A(n_59903), .B(n_59878), .C(axi_W[15]), .Z(n_1330)
		);
	notech_nao3 i_58445(.A(n_1330), .B(n_1329), .C(n_1643), .Z(n_1331));
	notech_nand2 i_548(.A(n_59836), .B(cacheQ[110]), .Z(n_1332));
	notech_nand3 i_547(.A(n_59903), .B(n_59878), .C(axi_W[14]), .Z(n_1333)
		);
	notech_nao3 i_58442(.A(n_1333), .B(n_1332), .C(n_1647), .Z(n_1334));
	notech_nand2 i_552(.A(n_59836), .B(cacheQ[109]), .Z(n_1335));
	notech_nand3 i_551(.A(n_59903), .B(n_59879), .C(axi_W[13]), .Z(n_1336)
		);
	notech_nao3 i_58439(.A(n_1336), .B(n_1335), .C(n_1651), .Z(n_1337));
	notech_nand2 i_556(.A(n_59836), .B(cacheQ[108]), .Z(n_1338));
	notech_nand3 i_555(.A(n_59897), .B(n_59879), .C(axi_W[12]), .Z(n_1339)
		);
	notech_nao3 i_58436(.A(n_1339), .B(n_1338), .C(n_1655), .Z(n_1340));
	notech_nand2 i_560(.A(n_59836), .B(cacheQ[107]), .Z(n_1341));
	notech_nand3 i_559(.A(n_59897), .B(n_59879), .C(axi_W[11]), .Z(n_1342)
		);
	notech_nao3 i_58433(.A(n_1342), .B(n_1341), .C(n_1659), .Z(n_1343));
	notech_nand2 i_564(.A(n_59836), .B(cacheQ[106]), .Z(n_1344));
	notech_nand3 i_563(.A(n_59897), .B(n_59879), .C(axi_W[10]), .Z(n_1345)
		);
	notech_nao3 i_58430(.A(n_1345), .B(n_1344), .C(n_1663), .Z(n_1346));
	notech_nand2 i_568(.A(n_59836), .B(cacheQ[105]), .Z(n_1347));
	notech_nand3 i_567(.A(n_59897), .B(n_59879), .C(axi_W[9]), .Z(n_1348));
	notech_nao3 i_58427(.A(n_1348), .B(n_1347), .C(n_1667), .Z(n_1349));
	notech_nand2 i_572(.A(n_59836), .B(cacheQ[104]), .Z(n_1350));
	notech_nand3 i_571(.A(n_59897), .B(n_59879), .C(axi_W[8]), .Z(n_1351));
	notech_nao3 i_58424(.A(n_1351), .B(n_1350), .C(n_1671), .Z(n_1352));
	notech_nand2 i_576(.A(n_59836), .B(cacheQ[103]), .Z(n_1353));
	notech_nand3 i_575(.A(n_59897), .B(n_59879), .C(axi_W[7]), .Z(n_1354));
	notech_nao3 i_58421(.A(n_1354), .B(n_1353), .C(n_1675), .Z(n_1355));
	notech_nand2 i_580(.A(n_59836), .B(cacheQ[102]), .Z(n_1356));
	notech_nand3 i_579(.A(n_59897), .B(n_59879), .C(axi_W[6]), .Z(n_1357));
	notech_nao3 i_58418(.A(n_1357), .B(n_1356), .C(n_1679), .Z(n_1358));
	notech_nand2 i_584(.A(n_59836), .B(cacheQ[101]), .Z(n_1359));
	notech_nand3 i_583(.A(n_59897), .B(n_59879), .C(axi_W[5]), .Z(n_1360));
	notech_nao3 i_58415(.A(n_1360), .B(n_1359), .C(n_1683), .Z(n_1361));
	notech_nand2 i_588(.A(n_59836), .B(cacheQ[100]), .Z(n_1362));
	notech_nand3 i_587(.A(n_59897), .B(n_59879), .C(axi_W[4]), .Z(n_1363));
	notech_nao3 i_58412(.A(n_1363), .B(n_1362), .C(n_1687), .Z(n_1364));
	notech_nand2 i_592(.A(n_59836), .B(cacheQ[99]), .Z(n_1365));
	notech_nand3 i_591(.A(n_59897), .B(n_59879), .C(axi_W[3]), .Z(n_1366));
	notech_nao3 i_58409(.A(n_1366), .B(n_1365), .C(n_1691), .Z(n_1367));
	notech_nand2 i_596(.A(n_59836), .B(cacheQ[98]), .Z(n_1368));
	notech_nand3 i_595(.A(n_59899), .B(n_59879), .C(axi_W[2]), .Z(n_1369));
	notech_nao3 i_58406(.A(n_1369), .B(n_1368), .C(n_1695), .Z(n_1370));
	notech_nand2 i_600(.A(n_59836), .B(cacheQ[97]), .Z(n_1371));
	notech_nand3 i_599(.A(n_59899), .B(n_59879), .C(axi_W[1]), .Z(n_1372));
	notech_nao3 i_58403(.A(n_1372), .B(n_1371), .C(n_1699), .Z(n_1373));
	notech_ao4 i_58978(.A(n_2073), .B(n_2109), .C(n_2072), .D(n_6976), .Z(n_1375
		));
	notech_nand2 i_607(.A(n_59836), .B(cacheQ[96]), .Z(n_1376));
	notech_or2 i_18(.A(n_59859), .B(n_2075), .Z(n_1377));
	notech_nand3 i_606(.A(n_59899), .B(n_59879), .C(axi_W[0]), .Z(n_1378));
	notech_nao3 i_58400(.A(n_1378), .B(n_1376), .C(n_1706), .Z(n_1379));
	notech_nand2 i_611(.A(cacheQ[95]), .B(n_1476), .Z(n_1380));
	notech_nao3 i_610(.A(n_59879), .B(axi_W[31]), .C(n_59899), .Z(n_1381));
	notech_nao3 i_58397(.A(n_1381), .B(n_1380), .C(n_1579), .Z(n_1382));
	notech_nand2 i_615(.A(n_1476), .B(cacheQ[94]), .Z(n_1383));
	notech_nao3 i_614(.A(n_59879), .B(axi_W[30]), .C(n_59899), .Z(n_1384));
	notech_nao3 i_58394(.A(n_1384), .B(n_1383), .C(n_1583), .Z(n_1385));
	notech_nand2 i_619(.A(n_1476), .B(cacheQ[93]), .Z(n_1386));
	notech_nao3 i_618(.A(n_59879), .B(axi_W[29]), .C(n_59897), .Z(n_1387));
	notech_nao3 i_58391(.A(n_1387), .B(n_1386), .C(n_1587), .Z(n_1388));
	notech_nand2 i_623(.A(n_1476), .B(cacheQ[92]), .Z(n_1389));
	notech_nao3 i_622(.A(n_59879), .B(axi_W[28]), .C(n_59897), .Z(n_1390));
	notech_nao3 i_58388(.A(n_1390), .B(n_1389), .C(n_1591), .Z(n_1391));
	notech_nand2 i_627(.A(n_1476), .B(cacheQ[91]), .Z(n_1392));
	notech_nao3 i_626(.A(n_59878), .B(axi_W[27]), .C(n_59899), .Z(n_1393));
	notech_nao3 i_58385(.A(n_1393), .B(n_1392), .C(n_1595), .Z(n_1394));
	notech_nand2 i_631(.A(n_1476), .B(cacheQ[90]), .Z(n_1395));
	notech_nao3 i_630(.A(n_59866), .B(axi_W[26]), .C(n_59899), .Z(n_1396));
	notech_nao3 i_58382(.A(n_1396), .B(n_1395), .C(n_1599), .Z(n_1397));
	notech_nand2 i_635(.A(n_1476), .B(cacheQ[89]), .Z(n_1398));
	notech_nao3 i_634(.A(n_59866), .B(axi_W[25]), .C(n_59906), .Z(n_1399));
	notech_nao3 i_58379(.A(n_1399), .B(n_1398), .C(n_1603), .Z(n_1400));
	notech_nand2 i_639(.A(n_1476), .B(cacheQ[88]), .Z(n_1401));
	notech_nao3 i_638(.A(n_59866), .B(axi_W[24]), .C(n_59906), .Z(n_1402));
	notech_nao3 i_58376(.A(n_1402), .B(n_1401), .C(n_1607), .Z(n_1403));
	notech_nand2 i_643(.A(n_1476), .B(cacheQ[87]), .Z(n_1404));
	notech_nao3 i_642(.A(n_59866), .B(axi_W[23]), .C(n_59906), .Z(n_1405));
	notech_nao3 i_58373(.A(n_1405), .B(n_1404), .C(n_1611), .Z(n_1406));
	notech_nand2 i_647(.A(n_1476), .B(cacheQ[86]), .Z(n_1407));
	notech_nao3 i_646(.A(n_59872), .B(axi_W[22]), .C(n_59906), .Z(n_1408));
	notech_nao3 i_58370(.A(n_1408), .B(n_1407), .C(n_1615), .Z(n_1409));
	notech_nand2 i_651(.A(n_1476), .B(cacheQ[85]), .Z(n_1410));
	notech_nao3 i_650(.A(n_59872), .B(axi_W[21]), .C(n_59906), .Z(n_1411));
	notech_nao3 i_58367(.A(n_1411), .B(n_1410), .C(n_1619), .Z(n_1412));
	notech_nand2 i_655(.A(n_1476), .B(cacheQ[84]), .Z(n_1413));
	notech_nao3 i_654(.A(n_59872), .B(axi_W[20]), .C(n_59904), .Z(n_1414));
	notech_nao3 i_58364(.A(n_1414), .B(n_1413), .C(n_1623), .Z(n_1415));
	notech_nand2 i_659(.A(n_1476), .B(cacheQ[83]), .Z(n_1416));
	notech_nao3 i_658(.A(n_59872), .B(axi_W[19]), .C(n_59904), .Z(n_1417));
	notech_nao3 i_58361(.A(n_1417), .B(n_1416), .C(n_1627), .Z(n_1418));
	notech_nand2 i_663(.A(n_1476), .B(cacheQ[82]), .Z(n_1419));
	notech_nao3 i_662(.A(n_59872), .B(axi_W[18]), .C(n_59906), .Z(n_1420));
	notech_nao3 i_58358(.A(n_1420), .B(n_1419), .C(n_1631), .Z(n_1421));
	notech_nand2 i_667(.A(n_1476), .B(cacheQ[81]), .Z(n_1422));
	notech_nao3 i_666(.A(n_59866), .B(axi_W[17]), .C(n_59904), .Z(n_1423));
	notech_nao3 i_58355(.A(n_1423), .B(n_1422), .C(n_1635), .Z(n_1424));
	notech_nand2 i_671(.A(n_1476), .B(cacheQ[80]), .Z(n_1425));
	notech_nao3 i_670(.A(n_59866), .B(axi_W[16]), .C(n_59906), .Z(n_1426));
	notech_nao3 i_58352(.A(n_1426), .B(n_1425), .C(n_1639), .Z(n_1427));
	notech_nand2 i_675(.A(n_59814), .B(cacheQ[79]), .Z(n_1428));
	notech_nao3 i_674(.A(n_59866), .B(axi_W[15]), .C(n_59906), .Z(n_1429));
	notech_nao3 i_58349(.A(n_1429), .B(n_1428), .C(n_1643), .Z(n_1430));
	notech_nand2 i_679(.A(n_59814), .B(cacheQ[78]), .Z(n_1431));
	notech_nao3 i_678(.A(n_59866), .B(axi_W[14]), .C(n_59906), .Z(n_1432));
	notech_nao3 i_58346(.A(n_1432), .B(n_1431), .C(n_1647), .Z(n_1433));
	notech_nand2 i_683(.A(n_59814), .B(cacheQ[77]), .Z(n_1434));
	notech_nao3 i_682(.A(n_59866), .B(axi_W[13]), .C(n_59906), .Z(n_1435));
	notech_nao3 i_58343(.A(n_1435), .B(n_1434), .C(n_1651), .Z(n_1436));
	notech_nand2 i_687(.A(n_59814), .B(cacheQ[76]), .Z(n_1437));
	notech_nao3 i_686(.A(n_59866), .B(axi_W[12]), .C(n_59906), .Z(n_1438));
	notech_nao3 i_58340(.A(n_1438), .B(n_1437), .C(n_1655), .Z(n_1439));
	notech_nand2 i_691(.A(n_59814), .B(cacheQ[75]), .Z(n_1440));
	notech_nao3 i_690(.A(n_59866), .B(axi_W[11]), .C(n_59906), .Z(n_1441));
	notech_nao3 i_58337(.A(n_1441), .B(n_1440), .C(n_1659), .Z(n_1442));
	notech_nand2 i_695(.A(n_59814), .B(cacheQ[74]), .Z(n_1443));
	notech_nao3 i_694(.A(n_59866), .B(axi_W[10]), .C(n_59906), .Z(n_1444));
	notech_nao3 i_58334(.A(n_1444), .B(n_1443), .C(n_1663), .Z(n_1445));
	notech_nand2 i_699(.A(n_59814), .B(cacheQ[73]), .Z(n_1446));
	notech_nao3 i_698(.A(n_59866), .B(axi_W[9]), .C(n_59906), .Z(n_1447));
	notech_nao3 i_58331(.A(n_1447), .B(n_1446), .C(n_1667), .Z(n_1448));
	notech_nand2 i_703(.A(n_59814), .B(cacheQ[72]), .Z(n_1449));
	notech_nao3 i_702(.A(n_59872), .B(axi_W[8]), .C(n_59906), .Z(n_1450));
	notech_nao3 i_58328(.A(n_1450), .B(n_1449), .C(n_1671), .Z(n_1451));
	notech_nand2 i_707(.A(n_59814), .B(cacheQ[71]), .Z(n_1452));
	notech_nao3 i_706(.A(n_59872), .B(axi_W[7]), .C(n_59906), .Z(n_1453));
	notech_nao3 i_58325(.A(n_1453), .B(n_1452), .C(n_1675), .Z(n_1454));
	notech_nand2 i_711(.A(n_59814), .B(cacheQ[70]), .Z(n_1455));
	notech_nao3 i_710(.A(n_59872), .B(axi_W[6]), .C(n_59904), .Z(n_1456));
	notech_nao3 i_58322(.A(n_1456), .B(n_1455), .C(n_1679), .Z(n_1457));
	notech_nand2 i_715(.A(n_59814), .B(cacheQ[69]), .Z(n_1458));
	notech_nao3 i_714(.A(n_59872), .B(axi_W[5]), .C(n_59903), .Z(n_1459));
	notech_nao3 i_58319(.A(n_1459), .B(n_1458), .C(n_1683), .Z(n_1460));
	notech_nand2 i_719(.A(n_59814), .B(cacheQ[68]), .Z(n_1461));
	notech_nao3 i_718(.A(n_59872), .B(axi_W[4]), .C(n_59904), .Z(n_1462));
	notech_nao3 i_58316(.A(n_1462), .B(n_1461), .C(n_1687), .Z(n_1463));
	notech_nand2 i_723(.A(n_59814), .B(cacheQ[67]), .Z(n_1464));
	notech_nao3 i_722(.A(n_59878), .B(axi_W[3]), .C(n_59904), .Z(n_1465));
	notech_nao3 i_58313(.A(n_1465), .B(n_1464), .C(n_1691), .Z(n_1466));
	notech_nand2 i_727(.A(n_59814), .B(cacheQ[66]), .Z(n_1467));
	notech_nao3 i_726(.A(n_59878), .B(axi_W[2]), .C(n_59903), .Z(n_1468));
	notech_nao3 i_58310(.A(n_1468), .B(n_1467), .C(n_1695), .Z(n_1469));
	notech_nand2 i_731(.A(n_59814), .B(cacheQ[65]), .Z(n_1470));
	notech_nao3 i_730(.A(n_59872), .B(axi_W[1]), .C(n_59903), .Z(n_1471));
	notech_nao3 i_58307(.A(n_1471), .B(n_1470), .C(n_1699), .Z(n_1472));
	notech_ao4 i_58977(.A(n_2073), .B(n_214256979), .C(n_2072), .D(n_6976), 
		.Z(n_1474));
	notech_nand2 i_738(.A(n_59814), .B(cacheQ[64]), .Z(n_1475));
	notech_or2 i_17(.A(n_59859), .B(n_2077), .Z(n_1476));
	notech_nao3 i_737(.A(n_59878), .B(axi_W[0]), .C(n_59903), .Z(n_1477));
	notech_nao3 i_58304(.A(n_1477), .B(n_1475), .C(n_1706), .Z(n_1478));
	notech_nand2 i_742(.A(cacheQ[63]), .B(n_1575), .Z(n_1479));
	notech_nand3 i_741(.A(n_59903), .B(n_59859), .C(axi_W[31]), .Z(n_1480)
		);
	notech_nao3 i_58301(.A(n_1480), .B(n_1479), .C(n_1579), .Z(n_1481));
	notech_nand2 i_746(.A(n_1575), .B(cacheQ[62]), .Z(n_1482));
	notech_nand3 i_745(.A(n_59903), .B(n_59859), .C(axi_W[30]), .Z(n_1483)
		);
	notech_nao3 i_58298(.A(n_1483), .B(n_1482), .C(n_1583), .Z(n_1484));
	notech_nand2 i_750(.A(n_1575), .B(cacheQ[61]), .Z(n_1485));
	notech_nand3 i_749(.A(n_59904), .B(n_59859), .C(axi_W[29]), .Z(n_1486)
		);
	notech_nao3 i_58295(.A(n_1486), .B(n_1485), .C(n_1587), .Z(n_1487));
	notech_nand2 i_754(.A(n_1575), .B(cacheQ[60]), .Z(n_1488));
	notech_nand3 i_753(.A(n_59904), .B(n_59859), .C(axi_W[28]), .Z(n_1489)
		);
	notech_nao3 i_58292(.A(n_1489), .B(n_1488), .C(n_1591), .Z(n_1490));
	notech_nand2 i_758(.A(n_1575), .B(cacheQ[59]), .Z(n_1491));
	notech_nand3 i_757(.A(n_59904), .B(n_59860), .C(axi_W[27]), .Z(n_1492)
		);
	notech_nao3 i_58289(.A(n_1492), .B(n_1491), .C(n_1595), .Z(n_1493));
	notech_nand2 i_762(.A(n_1575), .B(cacheQ[58]), .Z(n_1494));
	notech_nand3 i_761(.A(n_59904), .B(n_59859), .C(axi_W[26]), .Z(n_1495)
		);
	notech_nao3 i_58286(.A(n_1495), .B(n_1494), .C(n_1599), .Z(n_1496));
	notech_nand2 i_766(.A(n_1575), .B(cacheQ[57]), .Z(n_1497));
	notech_nand3 i_765(.A(n_59904), .B(n_59859), .C(axi_W[25]), .Z(n_1498)
		);
	notech_nao3 i_58283(.A(n_1498), .B(n_1497), .C(n_1603), .Z(n_1499));
	notech_nand2 i_770(.A(n_1575), .B(cacheQ[56]), .Z(n_1500));
	notech_nand3 i_769(.A(n_59904), .B(n_59859), .C(axi_W[24]), .Z(n_1501)
		);
	notech_nao3 i_58280(.A(n_1501), .B(n_1500), .C(n_1607), .Z(n_1502));
	notech_nand2 i_774(.A(n_1575), .B(cacheQ[55]), .Z(n_1503));
	notech_nand3 i_773(.A(n_59904), .B(n_59859), .C(axi_W[23]), .Z(n_1504)
		);
	notech_nao3 i_58277(.A(n_1504), .B(n_1503), .C(n_1611), .Z(n_1505));
	notech_nand2 i_778(.A(n_1575), .B(cacheQ[54]), .Z(n_1506));
	notech_nand3 i_777(.A(n_59904), .B(n_59859), .C(axi_W[22]), .Z(n_1507)
		);
	notech_nao3 i_58274(.A(n_1507), .B(n_1506), .C(n_1615), .Z(n_1508));
	notech_nand2 i_782(.A(n_1575), .B(cacheQ[53]), .Z(n_1509));
	notech_nand3 i_781(.A(n_59904), .B(n_59859), .C(axi_W[21]), .Z(n_1510)
		);
	notech_nao3 i_58271(.A(n_1510), .B(n_1509), .C(n_1619), .Z(n_1511));
	notech_nand2 i_786(.A(n_1575), .B(cacheQ[52]), .Z(n_1512));
	notech_nand3 i_785(.A(n_59904), .B(n_59859), .C(axi_W[20]), .Z(n_1513)
		);
	notech_nao3 i_58268(.A(n_1513), .B(n_1512), .C(n_1623), .Z(n_1514));
	notech_nand2 i_790(.A(n_1575), .B(cacheQ[51]), .Z(n_1515));
	notech_nand3 i_789(.A(n_59887), .B(n_59859), .C(axi_W[19]), .Z(n_1516)
		);
	notech_nao3 i_58265(.A(n_1516), .B(n_1515), .C(n_1627), .Z(n_1517));
	notech_nand2 i_794(.A(n_1575), .B(cacheQ[50]), .Z(n_1518));
	notech_nand3 i_793(.A(n_59887), .B(n_59859), .C(axi_W[18]), .Z(n_1519)
		);
	notech_nao3 i_58262(.A(n_1519), .B(n_1518), .C(n_1631), .Z(n_1520));
	notech_nand2 i_798(.A(n_1575), .B(cacheQ[49]), .Z(n_1521));
	notech_nand3 i_797(.A(n_59887), .B(n_59859), .C(axi_W[17]), .Z(n_1522)
		);
	notech_nao3 i_58259(.A(n_1522), .B(n_1521), .C(n_1635), .Z(n_1523));
	notech_nand2 i_802(.A(n_1575), .B(cacheQ[48]), .Z(n_1524));
	notech_nand3 i_801(.A(n_59887), .B(n_59859), .C(axi_W[16]), .Z(n_1525)
		);
	notech_nao3 i_58256(.A(n_1525), .B(n_1524), .C(n_1639), .Z(n_1526));
	notech_nand2 i_806(.A(n_59792), .B(cacheQ[47]), .Z(n_1527));
	notech_nand3 i_805(.A(n_59887), .B(n_59860), .C(axi_W[15]), .Z(n_1528)
		);
	notech_nao3 i_58253(.A(n_1528), .B(n_1527), .C(n_1643), .Z(n_1529));
	notech_nand2 i_810(.A(n_59792), .B(cacheQ[46]), .Z(n_1530));
	notech_nand3 i_809(.A(n_59887), .B(n_59860), .C(axi_W[14]), .Z(n_1531)
		);
	notech_nao3 i_58250(.A(n_1531), .B(n_1530), .C(n_1647), .Z(n_1532));
	notech_nand2 i_814(.A(n_59792), .B(cacheQ[45]), .Z(n_1533));
	notech_nand3 i_813(.A(n_59887), .B(n_59860), .C(axi_W[13]), .Z(n_1534)
		);
	notech_nao3 i_58247(.A(n_1534), .B(n_1533), .C(n_1651), .Z(n_1535));
	notech_nand2 i_818(.A(n_59792), .B(cacheQ[44]), .Z(n_1536));
	notech_nand3 i_817(.A(n_59887), .B(n_59860), .C(axi_W[12]), .Z(n_1537)
		);
	notech_nao3 i_58244(.A(n_1537), .B(n_1536), .C(n_1655), .Z(n_1538));
	notech_nand2 i_822(.A(n_59792), .B(cacheQ[43]), .Z(n_1539));
	notech_nand3 i_821(.A(n_59887), .B(n_59860), .C(axi_W[11]), .Z(n_1540)
		);
	notech_nao3 i_58241(.A(n_1540), .B(n_1539), .C(n_1659), .Z(n_1541));
	notech_nand2 i_826(.A(n_59792), .B(cacheQ[42]), .Z(n_1542));
	notech_nand3 i_825(.A(n_59887), .B(n_59860), .C(axi_W[10]), .Z(n_1543)
		);
	notech_nao3 i_58238(.A(n_1543), .B(n_1542), .C(n_1663), .Z(n_1544));
	notech_nand2 i_830(.A(n_59792), .B(cacheQ[41]), .Z(n_1545));
	notech_nand3 i_829(.A(n_59891), .B(n_59860), .C(axi_W[9]), .Z(n_1546));
	notech_nao3 i_58235(.A(n_1546), .B(n_1545), .C(n_1667), .Z(n_1547));
	notech_nand2 i_834(.A(n_59792), .B(cacheQ[40]), .Z(n_1548));
	notech_nand3 i_833(.A(n_59891), .B(n_59860), .C(axi_W[8]), .Z(n_1549));
	notech_nao3 i_58232(.A(n_1549), .B(n_1548), .C(n_1671), .Z(n_1550));
	notech_nand2 i_838(.A(n_59792), .B(cacheQ[39]), .Z(n_1551));
	notech_nand3 i_837(.A(n_59891), .B(n_59860), .C(axi_W[7]), .Z(n_1552));
	notech_nao3 i_58229(.A(n_1552), .B(n_1551), .C(n_1675), .Z(n_1553));
	notech_nand2 i_842(.A(n_59792), .B(cacheQ[38]), .Z(n_1554));
	notech_nand3 i_841(.A(n_59891), .B(n_59860), .C(axi_W[6]), .Z(n_1555));
	notech_nao3 i_58226(.A(n_1555), .B(n_1554), .C(n_1679), .Z(n_1556));
	notech_nand2 i_846(.A(n_59792), .B(cacheQ[37]), .Z(n_1557));
	notech_nand3 i_845(.A(n_59891), .B(n_59860), .C(axi_W[5]), .Z(n_1558));
	notech_nao3 i_58223(.A(n_1558), .B(n_1557), .C(n_1683), .Z(n_1559));
	notech_nand2 i_850(.A(n_59792), .B(cacheQ[36]), .Z(n_1560));
	notech_nand3 i_849(.A(n_59891), .B(n_59860), .C(axi_W[4]), .Z(n_1561));
	notech_nao3 i_58220(.A(n_1561), .B(n_1560), .C(n_1687), .Z(n_1562));
	notech_nand2 i_854(.A(n_59792), .B(cacheQ[35]), .Z(n_1563));
	notech_nand3 i_853(.A(n_59891), .B(n_59860), .C(axi_W[3]), .Z(n_1564));
	notech_nao3 i_58217(.A(n_1564), .B(n_1563), .C(n_1691), .Z(n_1565));
	notech_nand2 i_858(.A(n_59792), .B(cacheQ[34]), .Z(n_1566));
	notech_nand3 i_857(.A(n_59891), .B(n_59860), .C(axi_W[2]), .Z(n_1567));
	notech_nao3 i_58214(.A(n_1567), .B(n_1566), .C(n_1695), .Z(n_1568));
	notech_nand2 i_862(.A(n_59792), .B(cacheQ[33]), .Z(n_1569));
	notech_nand3 i_861(.A(n_59891), .B(n_59860), .C(axi_W[1]), .Z(n_1570));
	notech_nao3 i_58211(.A(n_1570), .B(n_1569), .C(n_1699), .Z(n_1571));
	notech_ao4 i_58976(.A(n_2073), .B(n_217757014), .C(n_2072), .D(n_6976), 
		.Z(n_1573));
	notech_nand2 i_869(.A(n_59792), .B(cacheQ[32]), .Z(n_1574));
	notech_nand2 i_16(.A(n_214456981), .B(n_6633), .Z(n_1575));
	notech_nand3 i_868(.A(n_59885), .B(n_59860), .C(axi_W[0]), .Z(n_1576));
	notech_nao3 i_58208(.A(n_1576), .B(n_1574), .C(n_1706), .Z(n_1577));
	notech_nand2 i_873(.A(cacheQ[31]), .B(n_1705), .Z(n_1578));
	notech_nor2 i_111(.A(n_2024), .B(n_6781), .Z(n_1579));
	notech_nao3 i_872(.A(n_59860), .B(axi_W[31]), .C(n_59885), .Z(n_1580));
	notech_nao3 i_58205(.A(n_1580), .B(n_1578), .C(n_1579), .Z(n_1581));
	notech_nand2 i_877(.A(n_1705), .B(cacheQ[30]), .Z(n_1582));
	notech_nor2 i_81(.A(n_2024), .B(n_6780), .Z(n_1583));
	notech_nao3 i_876(.A(n_59860), .B(axi_W[30]), .C(n_59885), .Z(n_1584));
	notech_nao3 i_58202(.A(n_1584), .B(n_1582), .C(n_1583), .Z(n_1585));
	notech_nand2 i_881(.A(n_1705), .B(cacheQ[29]), .Z(n_1586));
	notech_nor2 i_105(.A(n_2024), .B(n_6779), .Z(n_1587));
	notech_nao3 i_880(.A(n_59860), .B(axi_W[29]), .C(n_59885), .Z(n_1588));
	notech_nao3 i_58199(.A(n_1588), .B(n_1586), .C(n_1587), .Z(n_1589));
	notech_nand2 i_885(.A(n_1705), .B(cacheQ[28]), .Z(n_1590));
	notech_nor2 i_82(.A(n_2024), .B(n_6778), .Z(n_1591));
	notech_nao3 i_884(.A(n_59847), .B(axi_W[28]), .C(n_59885), .Z(n_1592));
	notech_nao3 i_58196(.A(n_1592), .B(n_1590), .C(n_1591), .Z(n_1593));
	notech_nand2 i_889(.A(n_1705), .B(cacheQ[27]), .Z(n_1594));
	notech_nor2 i_83(.A(n_2024), .B(n_6777), .Z(n_1595));
	notech_nao3 i_888(.A(n_59847), .B(axi_W[27]), .C(n_59885), .Z(n_1596));
	notech_nao3 i_58193(.A(n_1596), .B(n_1594), .C(n_1595), .Z(n_1597));
	notech_nand2 i_893(.A(n_1705), .B(cacheQ[26]), .Z(n_1598));
	notech_nor2 i_84(.A(n_2024), .B(n_6776), .Z(n_1599));
	notech_nao3 i_892(.A(n_59847), .B(axi_W[26]), .C(n_59885), .Z(n_1600));
	notech_nao3 i_58190(.A(n_1600), .B(n_1598), .C(n_1599), .Z(n_1601));
	notech_nand2 i_903(.A(n_1705), .B(cacheQ[25]), .Z(n_1602));
	notech_nor2 i_107(.A(n_2024), .B(n_6775), .Z(n_1603));
	notech_nao3 i_902(.A(n_59847), .B(axi_W[25]), .C(n_59885), .Z(n_1604));
	notech_nao3 i_58187(.A(n_1604), .B(n_1602), .C(n_1603), .Z(n_1605));
	notech_nand2 i_908(.A(n_1705), .B(cacheQ[24]), .Z(n_1606));
	notech_nor2 i_85(.A(n_61228), .B(n_6774), .Z(n_1607));
	notech_nao3 i_907(.A(n_59847), .B(axi_W[24]), .C(n_59885), .Z(n_1608));
	notech_nao3 i_58184(.A(n_1608), .B(n_1606), .C(n_1607), .Z(n_1609));
	notech_nand2 i_912(.A(n_1705), .B(cacheQ[23]), .Z(n_1610));
	notech_nor2 i_110(.A(n_61224), .B(n_6773), .Z(n_1611));
	notech_nao3 i_911(.A(n_59853), .B(axi_W[23]), .C(n_59885), .Z(n_1612));
	notech_nao3 i_58181(.A(n_1612), .B(n_1610), .C(n_1611), .Z(n_1613));
	notech_nand2 i_919(.A(n_1705), .B(cacheQ[22]), .Z(n_1614));
	notech_nor2 i_87(.A(n_61224), .B(n_6772), .Z(n_1615));
	notech_nao3 i_915(.A(n_59853), .B(axi_W[22]), .C(n_59887), .Z(n_1616));
	notech_nao3 i_58178(.A(n_1616), .B(n_1614), .C(n_1615), .Z(n_1617));
	notech_nand2 i_923(.A(n_1705), .B(cacheQ[21]), .Z(n_1618));
	notech_nor2 i_109(.A(n_61224), .B(n_6771), .Z(n_1619));
	notech_nao3 i_922(.A(n_59853), .B(axi_W[21]), .C(n_59887), .Z(n_1620));
	notech_nao3 i_58175(.A(n_1620), .B(n_1618), .C(n_1619), .Z(n_1621));
	notech_nand2 i_927(.A(n_1705), .B(cacheQ[20]), .Z(n_1622));
	notech_nor2 i_89(.A(n_61224), .B(n_6770), .Z(n_1623));
	notech_nao3 i_926(.A(n_59853), .B(axi_W[20]), .C(n_59887), .Z(n_1624));
	notech_nao3 i_58172(.A(n_1624), .B(n_1622), .C(n_1623), .Z(n_1625));
	notech_nand2 i_931(.A(n_1705), .B(cacheQ[19]), .Z(n_1626));
	notech_nor2 i_90(.A(n_61224), .B(n_6769), .Z(n_1627));
	notech_nao3 i_930(.A(n_59847), .B(axi_W[19]), .C(n_59887), .Z(n_1628));
	notech_nao3 i_58169(.A(n_1628), .B(n_1626), .C(n_1627), .Z(n_1629));
	notech_nand2 i_935(.A(n_1705), .B(cacheQ[18]), .Z(n_1630));
	notech_nor2 i_91(.A(n_61224), .B(n_6768), .Z(n_1631));
	notech_nao3 i_934(.A(n_59847), .B(axi_W[18]), .C(n_59885), .Z(n_1632));
	notech_nao3 i_58166(.A(n_1632), .B(n_1630), .C(n_1631), .Z(n_1633));
	notech_nand2 i_939(.A(n_1705), .B(cacheQ[17]), .Z(n_1634));
	notech_nor2 i_98(.A(n_61224), .B(n_6767), .Z(n_1635));
	notech_nao3 i_938(.A(n_59847), .B(axi_W[17]), .C(n_59885), .Z(n_1636));
	notech_nao3 i_58163(.A(n_1636), .B(n_1634), .C(n_1635), .Z(n_1637));
	notech_nand2 i_943(.A(n_1705), .B(cacheQ[16]), .Z(n_1638));
	notech_nor2 i_93(.A(n_61224), .B(n_6766), .Z(n_1639));
	notech_nao3 i_942(.A(n_59847), .B(axi_W[16]), .C(n_59885), .Z(n_1640));
	notech_nao3 i_58160(.A(n_1640), .B(n_1638), .C(n_1639), .Z(n_1641));
	notech_nand2 i_947(.A(n_59770), .B(cacheQ[15]), .Z(n_1642));
	notech_nor2 i_97(.A(n_61224), .B(n_6765), .Z(n_1643));
	notech_nao3 i_946(.A(n_59847), .B(axi_W[15]), .C(n_59885), .Z(n_1644));
	notech_nao3 i_58157(.A(n_1644), .B(n_1642), .C(n_1643), .Z(n_1645));
	notech_nand2 i_951(.A(n_59770), .B(cacheQ[14]), .Z(n_1646));
	notech_nor2 i_96(.A(n_61224), .B(n_6764), .Z(n_1647));
	notech_nao3 i_950(.A(n_59847), .B(axi_W[14]), .C(n_59885), .Z(n_1648));
	notech_nao3 i_58154(.A(n_1648), .B(n_1646), .C(n_1647), .Z(n_1649));
	notech_nand2 i_955(.A(n_59770), .B(cacheQ[13]), .Z(n_1650));
	notech_nor2 i_95(.A(n_61224), .B(n_6763), .Z(n_1651));
	notech_nao3 i_954(.A(n_59847), .B(axi_W[13]), .C(n_59894), .Z(n_1652));
	notech_nao3 i_58151(.A(n_1652), .B(n_1650), .C(n_1651), .Z(n_1653));
	notech_nand2 i_959(.A(n_59770), .B(cacheQ[12]), .Z(n_1654));
	notech_nor2 i_94(.A(n_61224), .B(n_6762), .Z(n_1655));
	notech_nao3 i_958(.A(n_59847), .B(axi_W[12]), .C(n_59894), .Z(n_1656));
	notech_nao3 i_58148(.A(n_1656), .B(n_1654), .C(n_1655), .Z(n_1657));
	notech_nand2 i_963(.A(n_59770), .B(cacheQ[11]), .Z(n_1658));
	notech_nor2 i_92(.A(n_61224), .B(n_6761), .Z(n_1659));
	notech_nao3 i_962(.A(n_59847), .B(axi_W[11]), .C(n_59894), .Z(n_1660));
	notech_nao3 i_58145(.A(n_1660), .B(n_1658), .C(n_1659), .Z(n_1661));
	notech_nand2 i_967(.A(n_59770), .B(cacheQ[10]), .Z(n_1662));
	notech_nor2 i_88(.A(n_61228), .B(n_6760), .Z(n_1663));
	notech_nao3 i_966(.A(n_59853), .B(axi_W[10]), .C(n_59894), .Z(n_1664));
	notech_nao3 i_58142(.A(n_1664), .B(n_1662), .C(n_1663), .Z(n_1665));
	notech_nand2 i_971(.A(n_59770), .B(cacheQ[9]), .Z(n_1666));
	notech_nor2 i_86(.A(n_61228), .B(n_6759), .Z(n_1667));
	notech_nao3 i_970(.A(n_59853), .B(axi_W[9]), .C(n_59894), .Z(n_1668));
	notech_nao3 i_58139(.A(n_1668), .B(n_1666), .C(n_1667), .Z(n_1669));
	notech_nand2 i_975(.A(n_59770), .B(cacheQ[8]), .Z(n_1670));
	notech_nor2 i_100(.A(n_61228), .B(n_6758), .Z(n_1671));
	notech_nao3 i_974(.A(n_59853), .B(axi_W[8]), .C(n_59894), .Z(n_1672));
	notech_nao3 i_58136(.A(n_1672), .B(n_1670), .C(n_1671), .Z(n_1673));
	notech_nand2 i_979(.A(n_59770), .B(cacheQ[7]), .Z(n_1674));
	notech_nor2 i_115(.A(n_61228), .B(n_6757), .Z(n_1675));
	notech_nao3 i_978(.A(n_59853), .B(axi_W[7]), .C(n_59894), .Z(n_1676));
	notech_nao3 i_58133(.A(n_1676), .B(n_1674), .C(n_1675), .Z(n_1677));
	notech_nand2 i_983(.A(n_59770), .B(cacheQ[6]), .Z(n_1678));
	notech_nor2 i_101(.A(n_61228), .B(n_6756), .Z(n_1679));
	notech_nao3 i_982(.A(n_59853), .B(axi_W[6]), .C(n_59894), .Z(n_1680));
	notech_nao3 i_58130(.A(n_1680), .B(n_1678), .C(n_1679), .Z(n_1681));
	notech_nand2 i_987(.A(n_59770), .B(cacheQ[5]), .Z(n_1682));
	notech_nor2 i_114(.A(n_61228), .B(n_6755), .Z(n_1683));
	notech_nao3 i_986(.A(n_59853), .B(axi_W[5]), .C(n_59894), .Z(n_1684));
	notech_nao3 i_58127(.A(n_1684), .B(n_1682), .C(n_1683), .Z(n_1685));
	notech_nand2 i_991(.A(n_59770), .B(cacheQ[4]), .Z(n_1686));
	notech_nor2 i_79(.A(n_61228), .B(n_6754), .Z(n_1687));
	notech_nao3 i_990(.A(n_59859), .B(axi_W[4]), .C(n_59894), .Z(n_1688));
	notech_nao3 i_58124(.A(n_1688), .B(n_1686), .C(n_1687), .Z(n_1689));
	notech_nand2 i_995(.A(n_59770), .B(cacheQ[3]), .Z(n_1690));
	notech_nor2 i_104(.A(n_61224), .B(n_6753), .Z(n_1691));
	notech_nao3 i_994(.A(n_59859), .B(axi_W[3]), .C(n_59897), .Z(n_1692));
	notech_nao3 i_58121(.A(n_1692), .B(n_1690), .C(n_1691), .Z(n_1693));
	notech_nand2 i_999(.A(n_59770), .B(cacheQ[2]), .Z(n_1694));
	notech_nor2 i_106(.A(n_61224), .B(n_6752), .Z(n_1695));
	notech_nao3 i_998(.A(n_59853), .B(axi_W[2]), .C(n_59897), .Z(n_1696));
	notech_nao3 i_58118(.A(n_1696), .B(n_1694), .C(n_1695), .Z(n_1697));
	notech_nand2 i_1003(.A(n_59770), .B(cacheQ[1]), .Z(n_1698));
	notech_nor2 i_112(.A(n_61224), .B(n_6751), .Z(n_1699));
	notech_nao3 i_1002(.A(n_59859), .B(axi_W[1]), .C(n_59897), .Z(n_1700));
	notech_nao3 i_58115(.A(n_1700), .B(n_1698), .C(n_1699), .Z(n_1701));
	notech_ao4 i_58975(.A(n_2038), .B(n_2073), .C(n_2072), .D(n_6976), .Z(n_1703
		));
	notech_nand2 i_1009(.A(n_59770), .B(cacheQ[0]), .Z(n_1704));
	notech_nand2 i_15(.A(n_6633), .B(n_214556982), .Z(n_1705));
	notech_nor2 i_103(.A(n_61228), .B(n_6750), .Z(n_1706));
	notech_nao3 i_1008(.A(n_59853), .B(axi_W[0]), .C(n_59897), .Z(n_1707));
	notech_nao3 i_58112(.A(n_1707), .B(n_1704), .C(n_1706), .Z(n_1708));
	notech_ao4 i_57522(.A(n_28023), .B(n_6973), .C(n_2004), .D(n_2007), .Z(n_1710
		));
	notech_or2 i_1014(.A(n_2032), .B(n_6977), .Z(n_1711));
	notech_nand3 i_1017(.A(n_59894), .B(n_59872), .C(axi_WSTRB[3]), .Z(n_1712
		));
	notech_nand3 i_58589(.A(n_61888), .B(n_221257049), .C(n_1712), .Z(n_1713
		));
	notech_nand3 i_1019(.A(n_59894), .B(n_59872), .C(axi_WSTRB[2]), .Z(n_1714
		));
	notech_nand3 i_58587(.A(n_61882), .B(n_221257049), .C(n_1714), .Z(n_1715
		));
	notech_nand3 i_1021(.A(n_59894), .B(n_59872), .C(axi_WSTRB[1]), .Z(n_1716
		));
	notech_nand3 i_58585(.A(n_61882), .B(n_221257049), .C(n_1716), .Z(n_1717
		));
	notech_nand3 i_1023(.A(n_59894), .B(axi_WSTRB[0]), .C(n_59872), .Z(n_1718
		));
	notech_nand3 i_58583(.A(n_61882), .B(n_221257049), .C(n_1718), .Z(n_1719
		));
	notech_nao3 i_1025(.A(n_59872), .B(axi_WSTRB[3]), .C(n_59894), .Z(n_1720
		));
	notech_nand3 i_58581(.A(n_61882), .B(n_221257049), .C(n_1720), .Z(n_1721
		));
	notech_nao3 i_1027(.A(n_59872), .B(axi_WSTRB[2]), .C(n_59892), .Z(n_1722
		));
	notech_nand3 i_58579(.A(n_61882), .B(n_221257049), .C(n_1722), .Z(n_1723
		));
	notech_nao3 i_1029(.A(n_59872), .B(axi_WSTRB[1]), .C(n_59892), .Z(n_1724
		));
	notech_nand3 i_58577(.A(n_61882), .B(n_221257049), .C(n_1724), .Z(n_1725
		));
	notech_nao3 i_1031(.A(n_59872), .B(axi_WSTRB[0]), .C(n_59892), .Z(n_1726
		));
	notech_nand3 i_58575(.A(n_61882), .B(n_221257049), .C(n_1726), .Z(n_1727
		));
	notech_nand3 i_1033(.A(n_59892), .B(n_59853), .C(axi_WSTRB[3]), .Z(n_1728
		));
	notech_nand3 i_58573(.A(n_61882), .B(n_221257049), .C(n_1728), .Z(n_1729
		));
	notech_nand3 i_1035(.A(n_59891), .B(n_59853), .C(axi_WSTRB[2]), .Z(n_1730
		));
	notech_nand3 i_58571(.A(n_61882), .B(n_221257049), .C(n_1730), .Z(n_1731
		));
	notech_nand3 i_1037(.A(n_59891), .B(n_59853), .C(axi_WSTRB[1]), .Z(n_1732
		));
	notech_nand3 i_58569(.A(n_61888), .B(n_221257049), .C(n_1732), .Z(n_1733
		));
	notech_nand3 i_1039(.A(n_59891), .B(n_59853), .C(axi_WSTRB[0]), .Z(n_1734
		));
	notech_nand3 i_58567(.A(n_61888), .B(n_221257049), .C(n_1734), .Z(n_1735
		));
	notech_nao3 i_1041(.A(n_59853), .B(axi_WSTRB[3]), .C(n_59891), .Z(n_1736
		));
	notech_nand3 i_58565(.A(n_61888), .B(n_221257049), .C(n_1736), .Z(n_1737
		));
	notech_nao3 i_1043(.A(n_59853), .B(axi_WSTRB[2]), .C(n_59891), .Z(n_1738
		));
	notech_nand3 i_58563(.A(n_61888), .B(n_221257049), .C(n_1738), .Z(n_1739
		));
	notech_nao3 i_1045(.A(n_59853), .B(axi_WSTRB[1]), .C(n_59892), .Z(n_1740
		));
	notech_nand3 i_58561(.A(n_61888), .B(n_221257049), .C(n_1740), .Z(n_1741
		));
	notech_and4 i_123(.A(fsm[2]), .B(fsm[4]), .C(fsm[0]), .D(n_1993), .Z(n_1742
		));
	notech_nand2 i_1047(.A(n_2052), .B(n_6624), .Z(n_1743));
	notech_ao3 i_60092(.A(n_2072), .B(n_1743), .C(n_1742), .Z(n_1744));
	notech_or4 i_1053(.A(A4[1]), .B(n_59921), .C(n_59892), .D(n_6749), .Z(n_1745
		));
	notech_nand3 i_58559(.A(n_61888), .B(n_221257049), .C(n_1745), .Z(n_1746
		));
	notech_or4 i_1057(.A(fsm[0]), .B(fsm[4]), .C(n_2012), .D(n_6632), .Z(n_1748
		));
	notech_and4 i_60404(.A(n_2032), .B(n_221657053), .C(n_1748), .D(n_221557052
		), .Z(n_1749));
	notech_nao3 i_63(.A(fsm[0]), .B(n_6738), .C(n_2012), .Z(n_1750));
	notech_nand2 i_58594(.A(n_221957056), .B(n_221557052), .Z(n_1752));
	notech_nand2 i_1066(.A(axi_ARREADY), .B(n_1754), .Z(n_1753));
	notech_nand3 i_129(.A(n_61228), .B(n_6677), .C(n_6625), .Z(n_1754));
	notech_and4 i_60377(.A(n_61257), .B(n_1743), .C(n_2023), .D(n_1753), .Z(n_1755
		));
	notech_nand2 i_58596(.A(n_61257), .B(n_2020), .Z(n_1756));
	notech_ao4 i_59139(.A(n_222957066), .B(n_222857065), .C(n_6747), .D(n_222257059
		), .Z(n_1758));
	notech_ao4 i_68(.A(n_222457061), .B(n_222357060), .C(n_222257059), .D(n_6747
		), .Z(n_1760));
	notech_ao4 i_58901(.A(n_222857065), .B(n_223157068), .C(n_6740), .D(n_222557062
		), .Z(n_1762));
	notech_ao4 i_59165(.A(n_6628), .B(n_6627), .C(n_222557062), .D(n_6740), 
		.Z(n_1763));
	notech_ao4 i_60234(.A(readio_ack), .B(n_6975), .C(n_222457061), .D(n_222357060
		), .Z(n_1766));
	notech_nand2 i_108(.A(n_61894), .B(n_28023), .Z(n_1767));
	notech_nand2 i_1121(.A(n_2058), .B(axi_AWREADY), .Z(n_1768));
	notech_and4 i_58635(.A(n_967), .B(n_61894), .C(n_28023), .D(n_1768), .Z(n_1769
		));
	notech_or4 i_1123(.A(fsm[3]), .B(n_6630), .C(fsm[2]), .D(n_6736), .Z(n_1770
		));
	notech_mux2 i_1(.S(n_223657073), .A(axi_AW[4]), .B(Daddr[4]), .Z(cacheA[
		0]));
	notech_mux2 i_211496(.S(n_223657073), .A(axi_AW[5]), .B(Daddr[5]), .Z(cacheA
		[1]));
	notech_mux2 i_3(.S(n_223657073), .A(axi_AW[6]), .B(Daddr[6]), .Z(cacheA[
		2]));
	notech_mux2 i_4(.S(n_223657073), .A(axi_AW[7]), .B(Daddr[7]), .Z(cacheA[
		3]));
	notech_mux2 i_511497(.S(n_223657073), .A(axi_AW[8]), .B(Daddr[8]), .Z(cacheA
		[4]));
	notech_mux2 i_6(.S(n_223657073), .A(axi_AW[9]), .B(Daddr[9]), .Z(cacheA[
		5]));
	notech_mux2 i_7(.S(n_223657073), .A(axi_AW[10]), .B(Daddr[10]), .Z(cacheA
		[6]));
	notech_mux2 i_8(.S(n_223657073), .A(axi_AW[11]), .B(Daddr[11]), .Z(cacheA
		[7]));
	notech_mux2 i_9(.S(n_223657073), .A(axi_AW[12]), .B(Daddr[12]), .Z(cacheA
		[8]));
	notech_mux2 i_10(.S(n_223657073), .A(axi_AW[13]), .B(Daddr[13]), .Z(cacheA
		[9]));
	notech_nand2 i_1163(.A(cacheQ[64]), .B(n_224357080), .Z(n_1805));
	notech_nand3 i_122038(.A(n_2246), .B(n_224157078), .C(n_1805), .Z(read_data
		[0]));
	notech_nand2 i_1172(.A(n_224357080), .B(cacheQ[65]), .Z(n_1811));
	notech_reg code_wack_reg(.CP(n_62350), .D(n_3152), .CD(n_61813), .Q(code_wack
		));
	notech_mux2 i_2328(.S(n_973), .A(n_29767), .B(code_wack), .Z(n_3152));
	notech_nand3 i_222039(.A(n_2249), .B(n_2248), .C(n_1811), .Z(read_data[1
		]));
	notech_reg code_ack_slow_reg(.CP(n_62350), .D(n_3158), .CD(n_61813), .Q(code_ack
		));
	notech_mux2 i_2336(.S(n_975), .A(n_27143), .B(code_ack), .Z(n_3158));
	notech_reg axi_AR_reg_0(.CP(n_62350), .D(n_3167), .CD(n_61813), .Q(axi_AR
		[0]));
	notech_and4 i_2346(.A(axi_AR[0]), .B(n_967), .C(n_1064), .D(n_971), .Z(n_3167
		));
	notech_reg axi_AR_reg_1(.CP(n_62350), .D(n_3173), .CD(n_61813), .Q(axi_AR
		[1]));
	notech_and4 i_2354(.A(n_967), .B(n_1064), .C(n_971), .D(axi_AR[1]), .Z(n_3173
		));
	notech_reg axi_AR_reg_2(.CP(n_62350), .D(n_3176), .CD(n_61813), .Q(axi_AR
		[2]));
	notech_mux2 i_2360(.S(n_1065), .A(n_6669), .B(axi_AR[2]), .Z(n_3176));
	notech_reg axi_AR_reg_3(.CP(n_62350), .D(n_3182), .CD(n_61813), .Q(axi_AR
		[3]));
	notech_mux2 i_2368(.S(n_1065), .A(n_6668), .B(axi_AR[3]), .Z(n_3182));
	notech_nand2 i_1181(.A(n_224357080), .B(cacheQ[66]), .Z(n_1817));
	notech_reg axi_AR_reg_4(.CP(n_62350), .D(n_3188), .CD(n_61813), .Q(axi_AR
		[4]));
	notech_mux2 i_2376(.S(n_1065), .A(n_6667), .B(axi_AR[4]), .Z(n_3188));
	notech_nand3 i_322040(.A(n_2252), .B(n_2251), .C(n_1817), .Z(read_data[2
		]));
	notech_reg axi_AR_reg_5(.CP(n_62350), .D(n_3194), .CD(n_61813), .Q(axi_AR
		[5]));
	notech_mux2 i_2384(.S(n_1065), .A(n_6666), .B(axi_AR[5]), .Z(n_3194));
	notech_reg axi_AR_reg_6(.CP(n_62350), .D(n_3200), .CD(n_61811), .Q(axi_AR
		[6]));
	notech_mux2 i_2392(.S(n_1065), .A(n_6665), .B(axi_AR[6]), .Z(n_3200));
	notech_reg axi_AR_reg_7(.CP(n_62350), .D(n_3206), .CD(n_61811), .Q(axi_AR
		[7]));
	notech_mux2 i_2400(.S(n_1065), .A(n_6664), .B(axi_AR[7]), .Z(n_3206));
	notech_reg axi_AR_reg_8(.CP(n_62350), .D(n_3212), .CD(n_61811), .Q(axi_AR
		[8]));
	notech_mux2 i_2408(.S(n_1065), .A(n_6663), .B(axi_AR[8]), .Z(n_3212));
	notech_reg axi_AR_reg_9(.CP(n_62350), .D(n_3218), .CD(n_61811), .Q(axi_AR
		[9]));
	notech_mux2 i_2416(.S(n_1065), .A(n_6662), .B(axi_AR[9]), .Z(n_3218));
	notech_nand2 i_1190(.A(n_224357080), .B(cacheQ[67]), .Z(n_1823));
	notech_reg axi_AR_reg_10(.CP(n_62350), .D(n_3224), .CD(n_61811), .Q(axi_AR
		[10]));
	notech_mux2 i_2424(.S(n_1065), .A(n_6661), .B(axi_AR[10]), .Z(n_3224));
	notech_nand3 i_422041(.A(n_2255), .B(n_2254), .C(n_1823), .Z(read_data[3
		]));
	notech_reg axi_AR_reg_11(.CP(n_62350), .D(n_3230), .CD(n_61813), .Q(axi_AR
		[11]));
	notech_mux2 i_2432(.S(n_1065), .A(n_6660), .B(axi_AR[11]), .Z(n_3230));
	notech_reg axi_AR_reg_12(.CP(n_62350), .D(n_3236), .CD(n_61811), .Q(axi_AR
		[12]));
	notech_mux2 i_2440(.S(n_1065), .A(n_6659), .B(axi_AR[12]), .Z(n_3236));
	notech_reg axi_AR_reg_13(.CP(n_62350), .D(n_3242), .CD(n_61811), .Q(axi_AR
		[13]));
	notech_mux2 i_2448(.S(n_1065), .A(n_6658), .B(axi_AR[13]), .Z(n_3242));
	notech_reg axi_AR_reg_14(.CP(n_62350), .D(n_3248), .CD(n_61813), .Q(axi_AR
		[14]));
	notech_mux2 i_2456(.S(n_1065), .A(n_6657), .B(axi_AR[14]), .Z(n_3248));
	notech_reg axi_AR_reg_15(.CP(n_62350), .D(n_3254), .CD(n_61814), .Q(axi_AR
		[15]));
	notech_mux2 i_2464(.S(n_1065), .A(n_6656), .B(axi_AR[15]), .Z(n_3254));
	notech_nand2 i_1199(.A(n_224357080), .B(cacheQ[68]), .Z(n_1829));
	notech_reg axi_AR_reg_16(.CP(n_62350), .D(n_3260), .CD(n_61814), .Q(axi_AR
		[16]));
	notech_mux2 i_2472(.S(n_1065), .A(n_6655), .B(axi_AR[16]), .Z(n_3260));
	notech_nand3 i_522042(.A(n_2258), .B(n_2257), .C(n_1829), .Z(read_data[4
		]));
	notech_reg axi_AR_reg_17(.CP(n_62366), .D(n_3266), .CD(n_61814), .Q(axi_AR
		[17]));
	notech_mux2 i_2480(.S(n_1065), .A(n_6654), .B(axi_AR[17]), .Z(n_3266));
	notech_reg axi_AR_reg_18(.CP(n_62366), .D(n_3272), .CD(n_61814), .Q(axi_AR
		[18]));
	notech_mux2 i_2488(.S(n_61246), .A(n_6653), .B(axi_AR[18]), .Z(n_3272)
		);
	notech_reg axi_AR_reg_19(.CP(n_62366), .D(n_3278), .CD(n_61814), .Q(axi_AR
		[19]));
	notech_mux2 i_2496(.S(n_61246), .A(n_6652), .B(axi_AR[19]), .Z(n_3278)
		);
	notech_reg axi_AR_reg_20(.CP(n_62366), .D(n_3284), .CD(n_61814), .Q(axi_AR
		[20]));
	notech_mux2 i_2504(.S(n_61246), .A(n_6651), .B(axi_AR[20]), .Z(n_3284)
		);
	notech_reg axi_AR_reg_21(.CP(n_62366), .D(n_3290), .CD(n_61814), .Q(axi_AR
		[21]));
	notech_mux2 i_2512(.S(n_61246), .A(n_6650), .B(axi_AR[21]), .Z(n_3290)
		);
	notech_nand2 i_1208(.A(n_224357080), .B(cacheQ[69]), .Z(n_1835));
	notech_reg axi_AR_reg_22(.CP(n_62366), .D(n_3296), .CD(n_61814), .Q(axi_AR
		[22]));
	notech_mux2 i_2520(.S(n_61246), .A(n_6649), .B(axi_AR[22]), .Z(n_3296)
		);
	notech_nand3 i_622043(.A(n_2261), .B(n_2260), .C(n_1835), .Z(read_data[5
		]));
	notech_reg axi_AR_reg_23(.CP(n_62366), .D(n_3302), .CD(n_61813), .Q(axi_AR
		[23]));
	notech_mux2 i_2528(.S(n_61246), .A(n_6648), .B(axi_AR[23]), .Z(n_3302)
		);
	notech_reg axi_AR_reg_24(.CP(n_62366), .D(n_3308), .CD(n_61813), .Q(axi_AR
		[24]));
	notech_mux2 i_2536(.S(n_61246), .A(n_6646), .B(axi_AR[24]), .Z(n_3308)
		);
	notech_reg axi_AR_reg_25(.CP(n_62366), .D(n_3314), .CD(n_61813), .Q(axi_AR
		[25]));
	notech_mux2 i_2544(.S(n_61246), .A(n_6645), .B(axi_AR[25]), .Z(n_3314)
		);
	notech_reg axi_AR_reg_26(.CP(n_62366), .D(n_3320), .CD(n_61813), .Q(axi_AR
		[26]));
	notech_mux2 i_2552(.S(n_61246), .A(n_6644), .B(axi_AR[26]), .Z(n_3320)
		);
	notech_reg axi_AR_reg_27(.CP(n_62366), .D(n_3326), .CD(n_61814), .Q(axi_AR
		[27]));
	notech_mux2 i_2560(.S(n_61246), .A(n_6643), .B(axi_AR[27]), .Z(n_3326)
		);
	notech_nand2 i_1217(.A(n_224357080), .B(cacheQ[70]), .Z(n_1841));
	notech_reg axi_AR_reg_28(.CP(n_62366), .D(n_3332), .CD(n_61814), .Q(axi_AR
		[28]));
	notech_mux2 i_2568(.S(n_61246), .A(n_6641), .B(axi_AR[28]), .Z(n_3332)
		);
	notech_nand3 i_722044(.A(n_2264), .B(n_2263), .C(n_1841), .Z(read_data[6
		]));
	notech_reg axi_AR_reg_29(.CP(n_62366), .D(n_3338), .CD(n_61813), .Q(axi_AR
		[29]));
	notech_mux2 i_2576(.S(n_61246), .A(n_6640), .B(axi_AR[29]), .Z(n_3338)
		);
	notech_reg axi_AR_reg_30(.CP(n_62366), .D(n_3344), .CD(n_61814), .Q(axi_AR
		[30]));
	notech_mux2 i_2584(.S(n_61246), .A(n_6639), .B(axi_AR[30]), .Z(n_3344)
		);
	notech_reg axi_AR_reg_31(.CP(n_62366), .D(n_3350), .CD(n_61810), .Q(axi_AR
		[31]));
	notech_mux2 i_2592(.S(n_61246), .A(n_6638), .B(axi_AR[31]), .Z(n_3350)
		);
	notech_reg axi_AW_reg_0(.CP(n_62366), .D(n_3359), .CD(n_61810), .Q(axi_AW
		[0]));
	notech_and4 i_2602(.A(n_967), .B(n_28023), .C(n_61888), .D(axi_AW[0]), .Z
		(n_3359));
	notech_reg axi_AW_reg_1(.CP(n_62366), .D(n_3365), .CD(n_61809), .Q(axi_AW
		[1]));
	notech_and4 i_2610(.A(n_967), .B(n_28023), .C(n_61894), .D(axi_AW[1]), .Z
		(n_3365));
	notech_nand2 i_1226(.A(n_224357080), .B(cacheQ[71]), .Z(n_1847));
	notech_reg axi_AW_reg_2(.CP(n_62366), .D(n_3368), .CD(n_61809), .Q(axi_AW
		[2]));
	notech_mux2 i_2616(.S(n_61867), .A(n_6701), .B(axi_AW[2]), .Z(n_3368));
	notech_nand3 i_822045(.A(n_2267), .B(n_2266), .C(n_1847), .Z(read_data[7
		]));
	notech_reg axi_AW_reg_3(.CP(n_62366), .D(n_3374), .CD(n_61810), .Q(axi_AW
		[3]));
	notech_mux2 i_2624(.S(n_61867), .A(n_6700), .B(axi_AW[3]), .Z(n_3374));
	notech_reg axi_AW_reg_4(.CP(n_62412), .D(n_3380), .CD(n_61810), .Q(axi_AW
		[4]));
	notech_mux2 i_2632(.S(n_61867), .A(n_6699), .B(axi_AW[4]), .Z(n_3380));
	notech_reg axi_AW_reg_5(.CP(n_62364), .D(n_3386), .CD(n_61810), .Q(axi_AW
		[5]));
	notech_mux2 i_2640(.S(n_61868), .A(n_6698), .B(axi_AW[5]), .Z(n_3386));
	notech_reg axi_AW_reg_6(.CP(n_62412), .D(n_3392), .CD(n_61810), .Q(axi_AW
		[6]));
	notech_mux2 i_2648(.S(n_61867), .A(n_6697), .B(axi_AW[6]), .Z(n_3392));
	notech_reg axi_AW_reg_7(.CP(n_62412), .D(n_3398), .CD(n_61809), .Q(axi_AW
		[7]));
	notech_mux2 i_2656(.S(n_61867), .A(n_6696), .B(axi_AW[7]), .Z(n_3398));
	notech_nand2 i_1235(.A(n_224357080), .B(cacheQ[72]), .Z(n_1853));
	notech_reg axi_AW_reg_8(.CP(n_62412), .D(n_3404), .CD(n_61809), .Q(axi_AW
		[8]));
	notech_mux2 i_2664(.S(n_61867), .A(n_6695), .B(axi_AW[8]), .Z(n_3404));
	notech_nand3 i_922046(.A(n_2270), .B(n_2269), .C(n_1853), .Z(read_data[8
		]));
	notech_reg axi_AW_reg_9(.CP(n_62412), .D(n_3410), .CD(n_61809), .Q(axi_AW
		[9]));
	notech_mux2 i_2672(.S(n_61867), .A(n_6694), .B(axi_AW[9]), .Z(n_3410));
	notech_reg axi_AW_reg_10(.CP(n_62412), .D(n_3416), .CD(n_61809), .Q(axi_AW
		[10]));
	notech_mux2 i_2680(.S(n_61867), .A(n_6693), .B(axi_AW[10]), .Z(n_3416)
		);
	notech_reg axi_AW_reg_11(.CP(n_62412), .D(n_3422), .CD(n_61809), .Q(axi_AW
		[11]));
	notech_mux2 i_2688(.S(n_61867), .A(n_6692), .B(axi_AW[11]), .Z(n_3422)
		);
	notech_reg axi_AW_reg_12(.CP(n_62412), .D(n_3428), .CD(n_61809), .Q(axi_AW
		[12]));
	notech_mux2 i_2696(.S(n_61867), .A(n_6691), .B(axi_AW[12]), .Z(n_3428)
		);
	notech_reg axi_AW_reg_13(.CP(n_62412), .D(n_3434), .CD(n_61809), .Q(axi_AW
		[13]));
	notech_mux2 i_2704(.S(n_61867), .A(n_6690), .B(axi_AW[13]), .Z(n_3434)
		);
	notech_nand2 i_1244(.A(n_224357080), .B(cacheQ[73]), .Z(n_1859));
	notech_reg axi_AW_reg_14(.CP(n_62412), .D(n_3440), .CD(n_61809), .Q(axi_AW
		[14]));
	notech_mux2 i_2712(.S(n_61867), .A(n_6689), .B(axi_AW[14]), .Z(n_3440)
		);
	notech_nand3 i_1022047(.A(n_2273), .B(n_2272), .C(n_1859), .Z(read_data[
		9]));
	notech_reg axi_AW_reg_15(.CP(n_62412), .D(n_3446), .CD(n_61810), .Q(axi_AW
		[15]));
	notech_mux2 i_2720(.S(n_61867), .A(n_6688), .B(axi_AW[15]), .Z(n_3446)
		);
	notech_reg axi_AW_reg_16(.CP(n_62412), .D(n_3452), .CD(n_61811), .Q(axi_AW
		[16]));
	notech_mux2 i_2728(.S(n_61867), .A(n_6687), .B(axi_AW[16]), .Z(n_3452)
		);
	notech_reg axi_AW_reg_17(.CP(n_62412), .D(n_3458), .CD(n_61811), .Q(axi_AW
		[17]));
	notech_mux2 i_2736(.S(n_61868), .A(n_6686), .B(axi_AW[17]), .Z(n_3458)
		);
	notech_reg axi_AW_reg_18(.CP(n_62412), .D(n_3464), .CD(n_61811), .Q(axi_AW
		[18]));
	notech_mux2 i_2744(.S(n_61868), .A(n_6685), .B(axi_AW[18]), .Z(n_3464)
		);
	notech_reg axi_AW_reg_19(.CP(n_62412), .D(n_3470), .CD(n_61811), .Q(axi_AW
		[19]));
	notech_mux2 i_2752(.S(n_61868), .A(n_6684), .B(axi_AW[19]), .Z(n_3470)
		);
	notech_nand2 i_1253(.A(n_224357080), .B(cacheQ[74]), .Z(n_1865));
	notech_reg axi_AW_reg_20(.CP(n_62412), .D(n_3476), .CD(n_61811), .Q(axi_AW
		[20]));
	notech_mux2 i_2760(.S(n_61868), .A(n_6683), .B(axi_AW[20]), .Z(n_3476)
		);
	notech_nand3 i_1122048(.A(n_2276), .B(n_2275), .C(n_1865), .Z(read_data[
		10]));
	notech_reg axi_AW_reg_21(.CP(n_62412), .D(n_3482), .CD(n_61811), .Q(axi_AW
		[21]));
	notech_mux2 i_2768(.S(n_61868), .A(n_6682), .B(axi_AW[21]), .Z(n_3482)
		);
	notech_reg axi_AW_reg_22(.CP(n_62412), .D(n_3488), .CD(n_61811), .Q(axi_AW
		[22]));
	notech_mux2 i_2776(.S(n_61868), .A(n_6681), .B(axi_AW[22]), .Z(n_3488)
		);
	notech_reg axi_AW_reg_23(.CP(n_62390), .D(n_3494), .CD(n_61811), .Q(axi_AW
		[23]));
	notech_mux2 i_2784(.S(n_61868), .A(n_6680), .B(axi_AW[23]), .Z(n_3494)
		);
	notech_reg axi_AW_reg_24(.CP(n_62364), .D(n_3500), .CD(n_61810), .Q(axi_AW
		[24]));
	notech_mux2 i_2792(.S(n_61868), .A(n_6679), .B(axi_AW[24]), .Z(n_3500)
		);
	notech_reg axi_AW_reg_25(.CP(n_62364), .D(n_3506), .CD(n_61810), .Q(axi_AW
		[25]));
	notech_mux2 i_2800(.S(n_61868), .A(n_6678), .B(axi_AW[25]), .Z(n_3506)
		);
	notech_nand2 i_1262(.A(n_224357080), .B(cacheQ[75]), .Z(n_1871));
	notech_reg axi_AW_reg_26(.CP(n_62364), .D(n_3512), .CD(n_61810), .Q(axi_AW
		[26]));
	notech_mux2 i_2808(.S(n_61868), .A(n_6676), .B(axi_AW[26]), .Z(n_3512)
		);
	notech_nand3 i_1222049(.A(n_2279), .B(n_2278), .C(n_1871), .Z(read_data[
		11]));
	notech_reg axi_AW_reg_27(.CP(n_62364), .D(n_3518), .CD(n_61810), .Q(axi_AW
		[27]));
	notech_mux2 i_2816(.S(n_61868), .A(n_6674), .B(axi_AW[27]), .Z(n_3518)
		);
	notech_reg axi_AW_reg_28(.CP(n_62364), .D(n_3524), .CD(n_61810), .Q(axi_AW
		[28]));
	notech_mux2 i_2824(.S(n_61868), .A(n_6673), .B(axi_AW[28]), .Z(n_3524)
		);
	notech_reg axi_AW_reg_29(.CP(n_62364), .D(n_3530), .CD(n_61810), .Q(axi_AW
		[29]));
	notech_mux2 i_2832(.S(n_61868), .A(n_6672), .B(axi_AW[29]), .Z(n_3530)
		);
	notech_reg axi_AW_reg_30(.CP(n_62364), .D(n_3536), .CD(n_61810), .Q(axi_AW
		[30]));
	notech_mux2 i_2840(.S(n_61868), .A(n_6671), .B(axi_AW[30]), .Z(n_3536)
		);
	notech_reg axi_AW_reg_31(.CP(n_62364), .D(n_3542), .CD(n_61810), .Q(axi_AW
		[31]));
	notech_mux2 i_2848(.S(n_61868), .A(n_6670), .B(axi_AW[31]), .Z(n_3542)
		);
	notech_nand2 i_1271(.A(n_224357080), .B(cacheQ[76]), .Z(n_1877));
	notech_reg_set burst_idx_reg_0(.CP(n_62364), .D(n_3548), .SD(1'b1), .Q(burst_idx
		[0]));
	notech_mux2 i_2856(.S(n_1170), .A(n_6702), .B(burst_idx[0]), .Z(n_3548)
		);
	notech_nand3 i_1322050(.A(n_2282), .B(n_2281), .C(n_1877), .Z(read_data[
		12]));
	notech_reg_set burst_idx_reg_1(.CP(n_62364), .D(n_3554), .SD(1'b1), .Q(burst_idx
		[1]));
	notech_mux2 i_2864(.S(n_1170), .A(n_30150), .B(burst_idx[1]), .Z(n_3554)
		);
	notech_reg_set burst_idx_reg_2(.CP(n_62364), .D(n_3560), .SD(1'b1), .Q(burst_idx
		[2]));
	notech_mux2 i_2872(.S(n_1170), .A(n_30155), .B(burst_idx[2]), .Z(n_3560)
		);
	notech_reg_set burst_idx_reg_3(.CP(n_62364), .D(n_3566), .SD(1'b1), .Q(burst_idx
		[3]));
	notech_mux2 i_2880(.S(n_1170), .A(n_30160), .B(burst_idx[3]), .Z(n_3566)
		);
	notech_reg_set burst_idx_reg_4(.CP(n_62364), .D(n_3572), .SD(1'b1), .Q(burst_idx
		[4]));
	notech_mux2 i_2888(.S(n_1170), .A(n_30165), .B(burst_idx[4]), .Z(n_3572)
		);
	notech_reg_set A4_reg_0(.CP(n_62364), .D(n_3578), .SD(1'b1), .Q(A4[0])
		);
	notech_mux2 i_2896(.S(\nbus_11697[0] ), .A(n_59892), .B(Daddr[2]), .Z(n_3578
		));
	notech_nand2 i_1280(.A(n_224357080), .B(cacheQ[77]), .Z(n_1883));
	notech_reg_set A4_reg_1(.CP(n_62364), .D(n_3584), .SD(1'b1), .Q(A4[1])
		);
	notech_mux2 i_2904(.S(\nbus_11697[0] ), .A(A4[1]), .B(Daddr[3]), .Z(n_3584
		));
	notech_nand3 i_1422051(.A(n_2285), .B(n_2284), .C(n_1883), .Z(read_data[
		13]));
	notech_reg axi_W_reg_0(.CP(n_62364), .D(n_3590), .CD(n_61814), .Q(axi_W[
		0]));
	notech_mux2 i_2912(.S(n_61868), .A(n_6710), .B(axi_W[0]), .Z(n_3590));
	notech_reg axi_W_reg_1(.CP(n_62364), .D(n_3596), .CD(n_61817), .Q(axi_W[
		1]));
	notech_mux2 i_2920(.S(n_61868), .A(n_6709), .B(axi_W[1]), .Z(n_3596));
	notech_reg axi_W_reg_2(.CP(n_62364), .D(n_3602), .CD(n_61817), .Q(axi_W[
		2]));
	notech_mux2 i_2928(.S(n_61867), .A(n_6708), .B(axi_W[2]), .Z(n_3602));
	notech_reg axi_W_reg_3(.CP(n_62412), .D(n_3608), .CD(n_61817), .Q(axi_W[
		3]));
	notech_mux2 i_2936(.S(n_61857), .A(n_6707), .B(axi_W[3]), .Z(n_3608));
	notech_reg axi_W_reg_4(.CP(n_62386), .D(n_3614), .CD(n_61817), .Q(axi_W[
		4]));
	notech_mux2 i_2944(.S(n_61857), .A(n_6706), .B(axi_W[4]), .Z(n_3614));
	notech_nand2 i_1289(.A(n_224357080), .B(cacheQ[78]), .Z(n_1889));
	notech_reg axi_W_reg_5(.CP(n_62362), .D(n_3620), .CD(n_61817), .Q(axi_W[
		5]));
	notech_mux2 i_2952(.S(n_61857), .A(n_6705), .B(axi_W[5]), .Z(n_3620));
	notech_nand3 i_1522052(.A(n_2288), .B(n_2287), .C(n_1889), .Z(read_data[
		14]));
	notech_reg axi_W_reg_6(.CP(n_62386), .D(n_3626), .CD(n_61817), .Q(axi_W[
		6]));
	notech_mux2 i_2960(.S(n_61857), .A(n_6704), .B(axi_W[6]), .Z(n_3626));
	notech_reg axi_W_reg_7(.CP(n_62386), .D(n_3632), .CD(n_61817), .Q(axi_W[
		7]));
	notech_mux2 i_2968(.S(n_61862), .A(n_6703), .B(axi_W[7]), .Z(n_3632));
	notech_reg axi_W_reg_8(.CP(n_62386), .D(n_3638), .CD(n_61817), .Q(axi_W[
		8]));
	notech_mux2 i_2976(.S(n_61862), .A(n_29532), .B(axi_W[8]), .Z(n_3638));
	notech_reg axi_W_reg_9(.CP(n_62386), .D(n_3644), .CD(n_61817), .Q(axi_W[
		9]));
	notech_mux2 i_2984(.S(n_61857), .A(n_29538), .B(axi_W[9]), .Z(n_3644));
	notech_reg axi_W_reg_10(.CP(n_62386), .D(n_3650), .CD(n_61817), .Q(axi_W
		[10]));
	notech_mux2 i_2992(.S(n_61857), .A(n_29544), .B(axi_W[10]), .Z(n_3650)
		);
	notech_nand2 i_1298(.A(n_224357080), .B(cacheQ[79]), .Z(n_1895));
	notech_reg axi_W_reg_11(.CP(n_62386), .D(n_3656), .CD(n_61817), .Q(axi_W
		[11]));
	notech_mux2 i_3000(.S(n_61857), .A(n_29550), .B(axi_W[11]), .Z(n_3656)
		);
	notech_nand3 i_1622053(.A(n_2291), .B(n_2290), .C(n_1895), .Z(read_data[
		15]));
	notech_reg axi_W_reg_12(.CP(n_62386), .D(n_3662), .CD(n_61817), .Q(axi_W
		[12]));
	notech_mux2 i_3008(.S(n_61857), .A(n_29556), .B(axi_W[12]), .Z(n_3662)
		);
	notech_reg axi_W_reg_13(.CP(n_62386), .D(n_3668), .CD(n_61817), .Q(axi_W
		[13]));
	notech_mux2 i_3016(.S(n_61857), .A(n_29562), .B(axi_W[13]), .Z(n_3668)
		);
	notech_reg axi_W_reg_14(.CP(n_62386), .D(n_3674), .CD(n_61817), .Q(axi_W
		[14]));
	notech_mux2 i_3024(.S(n_61857), .A(n_29568), .B(axi_W[14]), .Z(n_3674)
		);
	notech_reg axi_W_reg_15(.CP(n_62386), .D(n_3680), .CD(n_61817), .Q(axi_W
		[15]));
	notech_mux2 i_3032(.S(n_61857), .A(n_29574), .B(axi_W[15]), .Z(n_3680)
		);
	notech_reg axi_W_reg_16(.CP(n_62386), .D(n_3686), .CD(n_61817), .Q(axi_W
		[16]));
	notech_mux2 i_3040(.S(n_61857), .A(n_29580), .B(axi_W[16]), .Z(n_3686)
		);
	notech_nand2 i_1307(.A(n_54294), .B(cacheQ[80]), .Z(n_1901));
	notech_reg axi_W_reg_17(.CP(n_62386), .D(n_3692), .CD(n_61818), .Q(axi_W
		[17]));
	notech_mux2 i_3048(.S(n_61857), .A(n_29586), .B(axi_W[17]), .Z(n_3692)
		);
	notech_nand3 i_1722054(.A(n_2294), .B(n_2293), .C(n_1901), .Z(read_data[
		16]));
	notech_reg axi_W_reg_18(.CP(n_62386), .D(n_3698), .CD(n_61818), .Q(axi_W
		[18]));
	notech_mux2 i_3056(.S(n_61857), .A(n_29592), .B(axi_W[18]), .Z(n_3698)
		);
	notech_reg axi_W_reg_19(.CP(n_62386), .D(n_3704), .CD(n_61818), .Q(axi_W
		[19]));
	notech_mux2 i_3064(.S(n_61857), .A(n_29598), .B(axi_W[19]), .Z(n_3704)
		);
	notech_reg axi_W_reg_20(.CP(n_62386), .D(n_3710), .CD(n_61818), .Q(axi_W
		[20]));
	notech_mux2 i_3072(.S(n_61862), .A(n_29604), .B(axi_W[20]), .Z(n_3710)
		);
	notech_reg axi_W_reg_21(.CP(n_62386), .D(n_3716), .CD(n_61818), .Q(axi_W
		[21]));
	notech_mux2 i_3080(.S(n_61862), .A(n_29610), .B(axi_W[21]), .Z(n_3716)
		);
	notech_reg axi_W_reg_22(.CP(n_62386), .D(n_3722), .CD(n_61818), .Q(axi_W
		[22]));
	notech_mux2 i_3088(.S(n_61862), .A(n_29616), .B(axi_W[22]), .Z(n_3722)
		);
	notech_nand2 i_1316(.A(n_54294), .B(cacheQ[81]), .Z(n_1907));
	notech_reg axi_W_reg_23(.CP(n_62422), .D(n_3728), .CD(n_61818), .Q(axi_W
		[23]));
	notech_mux2 i_3096(.S(n_61862), .A(n_29622), .B(axi_W[23]), .Z(n_3728)
		);
	notech_nand3 i_1822055(.A(n_2297), .B(n_2296), .C(n_1907), .Z(read_data[
		17]));
	notech_reg axi_W_reg_24(.CP(n_62408), .D(n_3734), .CD(n_61818), .Q(axi_W
		[24]));
	notech_mux2 i_3104(.S(n_61862), .A(n_29628), .B(axi_W[24]), .Z(n_3734)
		);
	notech_reg axi_W_reg_25(.CP(n_62422), .D(n_3740), .CD(n_61818), .Q(axi_W
		[25]));
	notech_mux2 i_3112(.S(n_61867), .A(n_29634), .B(axi_W[25]), .Z(n_3740)
		);
	notech_reg axi_W_reg_26(.CP(n_62422), .D(n_3746), .CD(n_61818), .Q(axi_W
		[26]));
	notech_mux2 i_3120(.S(n_61862), .A(n_29640), .B(axi_W[26]), .Z(n_3746)
		);
	notech_reg axi_W_reg_27(.CP(n_62422), .D(n_3752), .CD(n_61818), .Q(axi_W
		[27]));
	notech_mux2 i_3128(.S(n_61862), .A(n_29646), .B(axi_W[27]), .Z(n_3752)
		);
	notech_reg axi_W_reg_28(.CP(n_62422), .D(n_3758), .CD(n_61818), .Q(axi_W
		[28]));
	notech_mux2 i_3136(.S(n_61862), .A(n_29652), .B(axi_W[28]), .Z(n_3758)
		);
	notech_nand2 i_1325(.A(n_54294), .B(cacheQ[82]), .Z(n_1913));
	notech_reg axi_W_reg_29(.CP(n_62422), .D(n_3764), .CD(n_61818), .Q(axi_W
		[29]));
	notech_mux2 i_3144(.S(n_61862), .A(n_29658), .B(axi_W[29]), .Z(n_3764)
		);
	notech_nand3 i_1922056(.A(n_2300), .B(n_2299), .C(n_1913), .Z(read_data[
		18]));
	notech_reg axi_W_reg_30(.CP(n_62422), .D(n_3770), .CD(n_61818), .Q(axi_W
		[30]));
	notech_mux2 i_3152(.S(n_61862), .A(n_29664), .B(axi_W[30]), .Z(n_3770)
		);
	notech_reg axi_W_reg_31(.CP(n_62422), .D(n_3776), .CD(n_61818), .Q(axi_W
		[31]));
	notech_mux2 i_3160(.S(n_61862), .A(n_29670), .B(axi_W[31]), .Z(n_3776)
		);
	notech_reg axi_RREADY_reg(.CP(n_62422), .D(n_3782), .CD(n_61818), .Q(axi_RREADY
		));
	notech_mux2 i_3168(.S(n_1202), .A(n_1203), .B(axi_RREADY), .Z(n_3782));
	notech_reg abort_reg(.CP(n_62422), .D(n_3788), .CD(n_61818), .Q(abort)
		);
	notech_mux2 i_3176(.S(n_1206), .A(n_1207), .B(abort), .Z(n_3788));
	notech_reg read_ack_slow_reg(.CP(n_62422), .D(n_3794), .CD(n_61815), .Q(read_ack
		));
	notech_mux2 i_3184(.S(n_1211), .A(n_1213), .B(read_ack), .Z(n_3794));
	notech_nand2 i_1334(.A(n_54294), .B(cacheQ[83]), .Z(n_1919));
	notech_reg wrint_ack_reg(.CP(n_62422), .D(n_3800), .CD(n_61815), .Q(write_ack
		));
	notech_mux2 i_3192(.S(n_1214), .A(n_6733), .B(write_ack), .Z(n_3800));
	notech_nand3 i_2022057(.A(n_2303), .B(n_2302), .C(n_1919), .Z(read_data[
		19]));
	notech_reg fsm_reg_0(.CP(n_62422), .D(n_3806), .CD(n_61815), .Q(fsm[0])
		);
	notech_mux2 i_3200(.S(n_1222), .A(n_6713), .B(fsm[0]), .Z(n_3806));
	notech_reg fsm_reg_1(.CP(n_62422), .D(n_3812), .CD(n_61815), .Q(fsm[1])
		);
	notech_mux2 i_3208(.S(n_1222), .A(n_1219), .B(fsm[1]), .Z(n_3812));
	notech_reg fsm_reg_2(.CP(n_62422), .D(n_3818), .CD(n_61815), .Q(fsm[2])
		);
	notech_mux2 i_3216(.S(n_1222), .A(n_1217), .B(fsm[2]), .Z(n_3818));
	notech_reg fsm_reg_3(.CP(n_62422), .D(n_3824), .CD(n_61815), .Q(fsm[3])
		);
	notech_mux2 i_3224(.S(n_1222), .A(n_6711), .B(fsm[3]), .Z(n_3824));
	notech_reg fsm_reg_4(.CP(n_62422), .D(n_3830), .CD(n_61815), .Q(fsm[4])
		);
	notech_mux2 i_3232(.S(n_1222), .A(n_1215), .B(fsm[4]), .Z(n_3830));
	notech_nand2 i_1343(.A(n_54294), .B(cacheQ[84]), .Z(n_1925));
	notech_reg_set cacheD_reg_0(.CP(n_62422), .D(n_3836), .SD(1'b1), .Q(cacheD
		[0]));
	notech_mux2 i_3240(.S(n_1703), .A(n_1708), .B(cacheD[0]), .Z(n_3836));
	notech_nand3 i_2122058(.A(n_2306), .B(n_2305), .C(n_1925), .Z(read_data[
		20]));
	notech_reg_set cacheD_reg_1(.CP(n_62386), .D(n_3842), .SD(1'b1), .Q(cacheD
		[1]));
	notech_mux2 i_3248(.S(n_1703), .A(n_1701), .B(cacheD[1]), .Z(n_3842));
	notech_reg_set cacheD_reg_2(.CP(n_62422), .D(n_3848), .SD(1'b1), .Q(cacheD
		[2]));
	notech_mux2 i_3256(.S(n_1703), .A(n_1697), .B(cacheD[2]), .Z(n_3848));
	notech_reg_set cacheD_reg_3(.CP(n_62410), .D(n_3854), .SD(1'b1), .Q(cacheD
		[3]));
	notech_mux2 i_3264(.S(n_1703), .A(n_1693), .B(cacheD[3]), .Z(n_3854));
	notech_reg_set cacheD_reg_4(.CP(n_62410), .D(n_3860), .SD(1'b1), .Q(cacheD
		[4]));
	notech_mux2 i_3272(.S(n_1703), .A(n_1689), .B(cacheD[4]), .Z(n_3860));
	notech_reg_set cacheD_reg_5(.CP(n_62410), .D(n_3866), .SD(1'b1), .Q(cacheD
		[5]));
	notech_mux2 i_3280(.S(n_1703), .A(n_1685), .B(cacheD[5]), .Z(n_3866));
	notech_nand2 i_1352(.A(n_54294), .B(cacheQ[85]), .Z(n_1931));
	notech_reg_set cacheD_reg_6(.CP(n_62410), .D(n_3872), .SD(1'b1), .Q(cacheD
		[6]));
	notech_mux2 i_3288(.S(n_1703), .A(n_1681), .B(cacheD[6]), .Z(n_3872));
	notech_nand3 i_2222059(.A(n_2309), .B(n_2308), .C(n_1931), .Z(read_data[
		21]));
	notech_reg_set cacheD_reg_7(.CP(n_62410), .D(n_3878), .SD(1'b1), .Q(cacheD
		[7]));
	notech_mux2 i_3296(.S(n_1703), .A(n_1677), .B(cacheD[7]), .Z(n_3878));
	notech_reg_set cacheD_reg_8(.CP(n_62410), .D(n_3884), .SD(1'b1), .Q(cacheD
		[8]));
	notech_mux2 i_3304(.S(n_1703), .A(n_1673), .B(cacheD[8]), .Z(n_3884));
	notech_reg_set cacheD_reg_9(.CP(n_62410), .D(n_3890), .SD(1'b1), .Q(cacheD
		[9]));
	notech_mux2 i_3312(.S(n_1703), .A(n_1669), .B(cacheD[9]), .Z(n_3890));
	notech_reg_set cacheD_reg_10(.CP(n_62410), .D(n_3896), .SD(1'b1), .Q(cacheD
		[10]));
	notech_mux2 i_3320(.S(n_1703), .A(n_1665), .B(cacheD[10]), .Z(n_3896));
	notech_reg_set cacheD_reg_11(.CP(n_62410), .D(n_3902), .SD(1'b1), .Q(cacheD
		[11]));
	notech_mux2 i_3328(.S(n_1703), .A(n_1661), .B(cacheD[11]), .Z(n_3902));
	notech_nand2 i_1361(.A(n_54294), .B(cacheQ[86]), .Z(n_1937));
	notech_reg_set cacheD_reg_12(.CP(n_62410), .D(n_3908), .SD(1'b1), .Q(cacheD
		[12]));
	notech_mux2 i_3336(.S(n_1703), .A(n_1657), .B(cacheD[12]), .Z(n_3908));
	notech_nand3 i_2322060(.A(n_2312), .B(n_2311), .C(n_1937), .Z(read_data[
		22]));
	notech_reg_set cacheD_reg_13(.CP(n_62410), .D(n_3914), .SD(1'b1), .Q(cacheD
		[13]));
	notech_mux2 i_3344(.S(n_1703), .A(n_1653), .B(cacheD[13]), .Z(n_3914));
	notech_reg_set cacheD_reg_14(.CP(n_62410), .D(n_3920), .SD(1'b1), .Q(cacheD
		[14]));
	notech_mux2 i_3352(.S(n_1703), .A(n_1649), .B(cacheD[14]), .Z(n_3920));
	notech_reg_set cacheD_reg_15(.CP(n_62410), .D(n_3926), .SD(1'b1), .Q(cacheD
		[15]));
	notech_mux2 i_3360(.S(n_1703), .A(n_1645), .B(cacheD[15]), .Z(n_3926));
	notech_reg_set cacheD_reg_16(.CP(n_62410), .D(n_3932), .SD(1'b1), .Q(cacheD
		[16]));
	notech_mux2 i_3368(.S(n_59781), .A(n_1641), .B(cacheD[16]), .Z(n_3932)
		);
	notech_reg_set cacheD_reg_17(.CP(n_62410), .D(n_3938), .SD(1'b1), .Q(cacheD
		[17]));
	notech_mux2 i_3376(.S(n_59781), .A(n_1637), .B(cacheD[17]), .Z(n_3938)
		);
	notech_nand2 i_1370(.A(n_54294), .B(cacheQ[87]), .Z(n_1943));
	notech_reg_set cacheD_reg_18(.CP(n_62410), .D(n_3944), .SD(1'b1), .Q(cacheD
		[18]));
	notech_mux2 i_3384(.S(n_59781), .A(n_1633), .B(cacheD[18]), .Z(n_3944)
		);
	notech_nand3 i_2422061(.A(n_2315), .B(n_2314), .C(n_1943), .Z(read_data[
		23]));
	notech_reg_set cacheD_reg_19(.CP(n_62410), .D(n_3950), .SD(1'b1), .Q(cacheD
		[19]));
	notech_mux2 i_3392(.S(n_59781), .A(n_1629), .B(cacheD[19]), .Z(n_3950)
		);
	notech_reg_set cacheD_reg_20(.CP(n_62410), .D(n_3956), .SD(1'b1), .Q(cacheD
		[20]));
	notech_mux2 i_3400(.S(n_59781), .A(n_1625), .B(cacheD[20]), .Z(n_3956)
		);
	notech_reg_set cacheD_reg_21(.CP(n_62388), .D(n_3962), .SD(1'b1), .Q(cacheD
		[21]));
	notech_mux2 i_3408(.S(n_59781), .A(n_1621), .B(cacheD[21]), .Z(n_3962)
		);
	notech_reg_set cacheD_reg_22(.CP(n_62362), .D(n_3968), .SD(1'b1), .Q(cacheD
		[22]));
	notech_mux2 i_3416(.S(n_59781), .A(n_1617), .B(cacheD[22]), .Z(n_3968)
		);
	notech_reg_set cacheD_reg_23(.CP(n_62362), .D(n_3974), .SD(1'b1), .Q(cacheD
		[23]));
	notech_mux2 i_3424(.S(n_59781), .A(n_1613), .B(cacheD[23]), .Z(n_3974)
		);
	notech_nand2 i_1379(.A(n_54294), .B(cacheQ[88]), .Z(n_1949));
	notech_reg_set cacheD_reg_24(.CP(n_62362), .D(n_3980), .SD(1'b1), .Q(cacheD
		[24]));
	notech_mux2 i_3432(.S(n_59781), .A(n_1609), .B(cacheD[24]), .Z(n_3980)
		);
	notech_nand3 i_2522062(.A(n_2318), .B(n_2317), .C(n_1949), .Z(read_data[
		24]));
	notech_reg_set cacheD_reg_25(.CP(n_62362), .D(n_3986), .SD(1'b1), .Q(cacheD
		[25]));
	notech_mux2 i_3440(.S(n_59781), .A(n_1605), .B(cacheD[25]), .Z(n_3986)
		);
	notech_reg_set cacheD_reg_26(.CP(n_62362), .D(n_3992), .SD(1'b1), .Q(cacheD
		[26]));
	notech_mux2 i_3448(.S(n_59781), .A(n_1601), .B(cacheD[26]), .Z(n_3992)
		);
	notech_reg_set cacheD_reg_27(.CP(n_62362), .D(n_3998), .SD(1'b1), .Q(cacheD
		[27]));
	notech_mux2 i_3456(.S(n_59781), .A(n_1597), .B(cacheD[27]), .Z(n_3998)
		);
	notech_reg_set cacheD_reg_28(.CP(n_62362), .D(n_4004), .SD(1'b1), .Q(cacheD
		[28]));
	notech_mux2 i_3464(.S(n_59781), .A(n_1593), .B(cacheD[28]), .Z(n_4004)
		);
	notech_reg_set cacheD_reg_29(.CP(n_62362), .D(n_4010), .SD(1'b1), .Q(cacheD
		[29]));
	notech_mux2 i_3472(.S(n_59781), .A(n_1589), .B(cacheD[29]), .Z(n_4010)
		);
	notech_nand2 i_1388(.A(n_54294), .B(cacheQ[89]), .Z(n_1955));
	notech_reg_set cacheD_reg_30(.CP(n_62362), .D(n_4016), .SD(1'b1), .Q(cacheD
		[30]));
	notech_mux2 i_3480(.S(n_59781), .A(n_1585), .B(cacheD[30]), .Z(n_4016)
		);
	notech_nand3 i_2622063(.A(n_2321), .B(n_2320), .C(n_1955), .Z(read_data[
		25]));
	notech_reg_set cacheD_reg_31(.CP(n_62362), .D(n_4022), .SD(1'b1), .Q(cacheD
		[31]));
	notech_mux2 i_3488(.S(n_59781), .A(n_1581), .B(cacheD[31]), .Z(n_4022)
		);
	notech_reg_set cacheD_reg_32(.CP(n_62362), .D(n_4028), .SD(1'b1), .Q(cacheD
		[32]));
	notech_mux2 i_3496(.S(n_1573), .A(n_1577), .B(cacheD[32]), .Z(n_4028));
	notech_reg_set cacheD_reg_33(.CP(n_62362), .D(n_4034), .SD(1'b1), .Q(cacheD
		[33]));
	notech_mux2 i_3504(.S(n_1573), .A(n_1571), .B(cacheD[33]), .Z(n_4034));
	notech_reg_set cacheD_reg_34(.CP(n_62362), .D(n_4040), .SD(1'b1), .Q(cacheD
		[34]));
	notech_mux2 i_3512(.S(n_1573), .A(n_1568), .B(cacheD[34]), .Z(n_4040));
	notech_reg_set cacheD_reg_35(.CP(n_62362), .D(n_4046), .SD(1'b1), .Q(cacheD
		[35]));
	notech_mux2 i_3520(.S(n_1573), .A(n_1565), .B(cacheD[35]), .Z(n_4046));
	notech_nand2 i_1397(.A(n_54294), .B(cacheQ[90]), .Z(n_1961));
	notech_reg_set cacheD_reg_36(.CP(n_62362), .D(n_4052), .SD(1'b1), .Q(cacheD
		[36]));
	notech_mux2 i_3528(.S(n_1573), .A(n_1562), .B(cacheD[36]), .Z(n_4052));
	notech_nand3 i_2722064(.A(n_2324), .B(n_2323), .C(n_1961), .Z(read_data[
		26]));
	notech_reg_set cacheD_reg_37(.CP(n_62362), .D(n_4058), .SD(1'b1), .Q(cacheD
		[37]));
	notech_mux2 i_3536(.S(n_1573), .A(n_1559), .B(cacheD[37]), .Z(n_4058));
	notech_reg_set cacheD_reg_38(.CP(n_62362), .D(n_4064), .SD(1'b1), .Q(cacheD
		[38]));
	notech_mux2 i_3544(.S(n_1573), .A(n_1556), .B(cacheD[38]), .Z(n_4064));
	notech_reg_set cacheD_reg_39(.CP(n_62362), .D(n_4070), .SD(1'b1), .Q(cacheD
		[39]));
	notech_mux2 i_3552(.S(n_1573), .A(n_1553), .B(cacheD[39]), .Z(n_4070));
	notech_reg_set cacheD_reg_40(.CP(n_62410), .D(n_4076), .SD(1'b1), .Q(cacheD
		[40]));
	notech_mux2 i_3560(.S(n_1573), .A(n_1550), .B(cacheD[40]), .Z(n_4076));
	notech_reg_set cacheD_reg_41(.CP(n_62380), .D(n_4082), .SD(1'b1), .Q(cacheD
		[41]));
	notech_mux2 i_3568(.S(n_1573), .A(n_1547), .B(cacheD[41]), .Z(n_4082));
	notech_nand2 i_1406(.A(n_54294), .B(cacheQ[91]), .Z(n_1967));
	notech_reg_set cacheD_reg_42(.CP(n_62380), .D(n_4088), .SD(1'b1), .Q(cacheD
		[42]));
	notech_mux2 i_3576(.S(n_1573), .A(n_1544), .B(cacheD[42]), .Z(n_4088));
	notech_nand3 i_2822065(.A(n_2327), .B(n_2326), .C(n_1967), .Z(read_data[
		27]));
	notech_reg_set cacheD_reg_43(.CP(n_62380), .D(n_4094), .SD(1'b1), .Q(cacheD
		[43]));
	notech_mux2 i_3584(.S(n_1573), .A(n_1541), .B(cacheD[43]), .Z(n_4094));
	notech_reg_set cacheD_reg_44(.CP(n_62380), .D(n_4100), .SD(1'b1), .Q(cacheD
		[44]));
	notech_mux2 i_3592(.S(n_1573), .A(n_1538), .B(cacheD[44]), .Z(n_4100));
	notech_reg_set cacheD_reg_45(.CP(n_62380), .D(n_4106), .SD(1'b1), .Q(cacheD
		[45]));
	notech_mux2 i_3600(.S(n_1573), .A(n_1535), .B(cacheD[45]), .Z(n_4106));
	notech_reg_set cacheD_reg_46(.CP(n_62380), .D(n_4112), .SD(1'b1), .Q(cacheD
		[46]));
	notech_mux2 i_3608(.S(n_1573), .A(n_1532), .B(cacheD[46]), .Z(n_4112));
	notech_reg_set cacheD_reg_47(.CP(n_62380), .D(n_4118), .SD(1'b1), .Q(cacheD
		[47]));
	notech_mux2 i_3616(.S(n_1573), .A(n_1529), .B(cacheD[47]), .Z(n_4118));
	notech_nand2 i_1415(.A(n_54294), .B(cacheQ[92]), .Z(n_1973));
	notech_reg_set cacheD_reg_48(.CP(n_62380), .D(n_4124), .SD(1'b1), .Q(cacheD
		[48]));
	notech_mux2 i_3624(.S(n_59803), .A(n_1526), .B(cacheD[48]), .Z(n_4124)
		);
	notech_nand3 i_2922066(.A(n_2330), .B(n_2329), .C(n_1973), .Z(read_data[
		28]));
	notech_reg_set cacheD_reg_49(.CP(n_62380), .D(n_4130), .SD(1'b1), .Q(cacheD
		[49]));
	notech_mux2 i_3632(.S(n_59803), .A(n_1523), .B(cacheD[49]), .Z(n_4130)
		);
	notech_reg_set cacheD_reg_50(.CP(n_62380), .D(n_4136), .SD(1'b1), .Q(cacheD
		[50]));
	notech_mux2 i_3640(.S(n_59803), .A(n_1520), .B(cacheD[50]), .Z(n_4136)
		);
	notech_reg_set cacheD_reg_51(.CP(n_62380), .D(n_4142), .SD(1'b1), .Q(cacheD
		[51]));
	notech_mux2 i_3648(.S(n_59803), .A(n_1517), .B(cacheD[51]), .Z(n_4142)
		);
	notech_reg_set cacheD_reg_52(.CP(n_62380), .D(n_4148), .SD(1'b1), .Q(cacheD
		[52]));
	notech_mux2 i_3656(.S(n_59803), .A(n_1514), .B(cacheD[52]), .Z(n_4148)
		);
	notech_reg_set cacheD_reg_53(.CP(n_62380), .D(n_4154), .SD(1'b1), .Q(cacheD
		[53]));
	notech_mux2 i_3664(.S(n_59803), .A(n_1511), .B(cacheD[53]), .Z(n_4154)
		);
	notech_nand2 i_1424(.A(n_54294), .B(cacheQ[93]), .Z(n_1979));
	notech_reg_set cacheD_reg_54(.CP(n_62380), .D(n_4160), .SD(1'b1), .Q(cacheD
		[54]));
	notech_mux2 i_3672(.S(n_59803), .A(n_1508), .B(cacheD[54]), .Z(n_4160)
		);
	notech_nand3 i_3022067(.A(n_2333), .B(n_2332), .C(n_1979), .Z(read_data[
		29]));
	notech_reg_set cacheD_reg_55(.CP(n_62380), .D(n_4166), .SD(1'b1), .Q(cacheD
		[55]));
	notech_mux2 i_3680(.S(n_59803), .A(n_1505), .B(cacheD[55]), .Z(n_4166)
		);
	notech_reg_set cacheD_reg_56(.CP(n_62380), .D(n_4172), .SD(1'b1), .Q(cacheD
		[56]));
	notech_mux2 i_3688(.S(n_59803), .A(n_1502), .B(cacheD[56]), .Z(n_4172)
		);
	notech_reg_set cacheD_reg_57(.CP(n_62380), .D(n_4178), .SD(1'b1), .Q(cacheD
		[57]));
	notech_mux2 i_3696(.S(n_59803), .A(n_1499), .B(cacheD[57]), .Z(n_4178)
		);
	notech_reg_set cacheD_reg_58(.CP(n_62380), .D(n_4184), .SD(1'b1), .Q(cacheD
		[58]));
	notech_mux2 i_3704(.S(n_59803), .A(n_1496), .B(cacheD[58]), .Z(n_4184)
		);
	notech_reg_set cacheD_reg_59(.CP(n_62380), .D(n_4190), .SD(1'b1), .Q(cacheD
		[59]));
	notech_mux2 i_3712(.S(n_59803), .A(n_1493), .B(cacheD[59]), .Z(n_4190)
		);
	notech_nand2 i_1433(.A(n_54294), .B(cacheQ[94]), .Z(n_1985));
	notech_reg_set cacheD_reg_60(.CP(n_62418), .D(n_4196), .SD(1'b1), .Q(cacheD
		[60]));
	notech_mux2 i_3720(.S(n_59803), .A(n_1490), .B(cacheD[60]), .Z(n_4196)
		);
	notech_nand3 i_3122068(.A(n_2336), .B(n_2335), .C(n_1985), .Z(read_data[
		30]));
	notech_reg_set cacheD_reg_61(.CP(n_62402), .D(n_4202), .SD(1'b1), .Q(cacheD
		[61]));
	notech_mux2 i_3728(.S(n_59803), .A(n_1487), .B(cacheD[61]), .Z(n_4202)
		);
	notech_reg_set cacheD_reg_62(.CP(n_62418), .D(n_4208), .SD(1'b1), .Q(cacheD
		[62]));
	notech_mux2 i_3736(.S(n_59803), .A(n_1484), .B(cacheD[62]), .Z(n_4208)
		);
	notech_reg_set cacheD_reg_63(.CP(n_62418), .D(n_4214), .SD(1'b1), .Q(cacheD
		[63]));
	notech_mux2 i_3744(.S(n_59803), .A(n_1481), .B(cacheD[63]), .Z(n_4214)
		);
	notech_reg_set cacheD_reg_64(.CP(n_62418), .D(n_4220), .SD(1'b1), .Q(cacheD
		[64]));
	notech_mux2 i_3752(.S(n_1474), .A(n_1478), .B(cacheD[64]), .Z(n_4220));
	notech_reg_set cacheD_reg_65(.CP(n_62418), .D(n_4226), .SD(1'b1), .Q(cacheD
		[65]));
	notech_mux2 i_3760(.S(n_1474), .A(n_1472), .B(cacheD[65]), .Z(n_4226));
	notech_nand2 i_1442(.A(cacheQ[95]), .B(n_54294), .Z(n_1991));
	notech_reg_set cacheD_reg_66(.CP(n_62418), .D(n_4232), .SD(1'b1), .Q(cacheD
		[66]));
	notech_mux2 i_3768(.S(n_1474), .A(n_1469), .B(cacheD[66]), .Z(n_4232));
	notech_nand3 i_3222069(.A(n_2339), .B(n_2338), .C(n_1991), .Z(read_data[
		31]));
	notech_reg_set cacheD_reg_67(.CP(n_62418), .D(n_4238), .SD(1'b1), .Q(cacheD
		[67]));
	notech_mux2 i_3776(.S(n_1474), .A(n_1466), .B(cacheD[67]), .Z(n_4238));
	notech_and2 i_64(.A(fsm[3]), .B(fsm[1]), .Z(n_1993));
	notech_reg_set cacheD_reg_68(.CP(n_62418), .D(n_4244), .SD(1'b1), .Q(cacheD
		[68]));
	notech_mux2 i_3784(.S(n_1474), .A(n_1463), .B(cacheD[68]), .Z(n_4244));
	notech_reg_set cacheD_reg_69(.CP(n_62418), .D(n_4250), .SD(1'b1), .Q(cacheD
		[69]));
	notech_mux2 i_3792(.S(n_1474), .A(n_1460), .B(cacheD[69]), .Z(n_4250));
	notech_reg_set cacheD_reg_70(.CP(n_62418), .D(n_4256), .SD(1'b1), .Q(cacheD
		[70]));
	notech_mux2 i_3800(.S(n_1474), .A(n_1457), .B(cacheD[70]), .Z(n_4256));
	notech_or4 i_1329639(.A(fsm[0]), .B(n_6634), .C(n_6737), .D(n_6738), .Z(n_1996
		));
	notech_reg_set cacheD_reg_71(.CP(n_62418), .D(n_4262), .SD(1'b1), .Q(cacheD
		[71]));
	notech_mux2 i_3808(.S(n_1474), .A(n_1454), .B(cacheD[71]), .Z(n_4262));
	notech_reg_set cacheD_reg_72(.CP(n_62418), .D(n_4268), .SD(1'b1), .Q(cacheD
		[72]));
	notech_mux2 i_3816(.S(n_1474), .A(n_1451), .B(cacheD[72]), .Z(n_4268));
	notech_nao3 i_56(.A(n_6737), .B(n_6736), .C(fsm[3]), .Z(n_1998));
	notech_reg_set cacheD_reg_73(.CP(n_62418), .D(n_4274), .SD(1'b1), .Q(cacheD
		[73]));
	notech_mux2 i_3824(.S(n_1474), .A(n_1448), .B(cacheD[73]), .Z(n_4274));
	notech_and2 i_45(.A(n_6735), .B(n_6738), .Z(n_1999));
	notech_reg_set cacheD_reg_74(.CP(n_62418), .D(n_4280), .SD(1'b1), .Q(cacheD
		[74]));
	notech_mux2 i_3832(.S(n_1474), .A(n_1445), .B(cacheD[74]), .Z(n_4280));
	notech_nor2 i_57399(.A(write_ack), .B(n_6982), .Z(n_2000));
	notech_reg_set cacheD_reg_75(.CP(n_62418), .D(n_4286), .SD(1'b1), .Q(cacheD
		[75]));
	notech_mux2 i_3840(.S(n_1474), .A(n_1442), .B(cacheD[75]), .Z(n_4286));
	notech_and2 i_23(.A(n_6978), .B(read_req), .Z(n_2001));
	notech_reg_set cacheD_reg_76(.CP(n_62418), .D(n_4292), .SD(1'b1), .Q(cacheD
		[76]));
	notech_mux2 i_3848(.S(n_1474), .A(n_1439), .B(cacheD[76]), .Z(n_4292));
	notech_reg_set cacheD_reg_77(.CP(n_62418), .D(n_4298), .SD(1'b1), .Q(cacheD
		[77]));
	notech_mux2 i_3856(.S(n_1474), .A(n_1436), .B(cacheD[77]), .Z(n_4298));
	notech_ao3 i_13(.A(n_61972), .B(n_61873), .C(n_1742), .Z(n_2003));
	notech_reg_set cacheD_reg_78(.CP(n_62418), .D(n_4304), .SD(1'b1), .Q(cacheD
		[78]));
	notech_mux2 i_3864(.S(n_1474), .A(n_1433), .B(cacheD[78]), .Z(n_4304));
	notech_or4 i_40(.A(fsm[0]), .B(fsm[4]), .C(n_1998), .D(n_2000), .Z(n_2004
		));
	notech_reg_set cacheD_reg_79(.CP(n_62418), .D(n_4310), .SD(1'b1), .Q(cacheD
		[79]));
	notech_mux2 i_3872(.S(n_1474), .A(n_1430), .B(cacheD[79]), .Z(n_4310));
	notech_reg_set cacheD_reg_80(.CP(n_62416), .D(n_4316), .SD(1'b1), .Q(cacheD
		[80]));
	notech_mux2 i_3880(.S(n_59825), .A(n_1427), .B(cacheD[80]), .Z(n_4316)
		);
	notech_reg_set cacheD_reg_81(.CP(n_62424), .D(n_4322), .SD(1'b1), .Q(cacheD
		[81]));
	notech_mux2 i_3888(.S(n_59825), .A(n_1424), .B(cacheD[81]), .Z(n_4322)
		);
	notech_or4 i_141(.A(code_wack), .B(n_969), .C(n_2001), .D(n_6981), .Z(n_2007
		));
	notech_reg_set cacheD_reg_82(.CP(n_62424), .D(n_4328), .SD(1'b1), .Q(cacheD
		[82]));
	notech_mux2 i_3896(.S(n_59825), .A(n_1421), .B(cacheD[82]), .Z(n_4328)
		);
	notech_or2 i_57510(.A(n_2007), .B(n_2004), .Z(n_2008));
	notech_reg_set cacheD_reg_83(.CP(n_62424), .D(n_4334), .SD(1'b1), .Q(cacheD
		[83]));
	notech_mux2 i_3904(.S(n_59825), .A(n_1418), .B(cacheD[83]), .Z(n_4334)
		);
	notech_reg_set cacheD_reg_84(.CP(n_62424), .D(n_4340), .SD(1'b1), .Q(cacheD
		[84]));
	notech_mux2 i_3912(.S(n_59825), .A(n_1415), .B(cacheD[84]), .Z(n_4340)
		);
	notech_or4 i_57497(.A(code_ack), .B(n_2001), .C(n_2004), .D(n_6979), .Z(n_2010
		));
	notech_reg_set cacheD_reg_85(.CP(n_62424), .D(n_4346), .SD(1'b1), .Q(cacheD
		[85]));
	notech_mux2 i_3920(.S(n_59825), .A(n_1412), .B(cacheD[85]), .Z(n_4346)
		);
	notech_reg_set cacheD_reg_86(.CP(n_62424), .D(n_4352), .SD(1'b1), .Q(cacheD
		[86]));
	notech_mux2 i_3928(.S(n_59825), .A(n_1409), .B(cacheD[86]), .Z(n_4352)
		);
	notech_nand3 i_102(.A(fsm[3]), .B(n_6737), .C(n_6736), .Z(n_2012));
	notech_reg_set cacheD_reg_87(.CP(n_62424), .D(n_4358), .SD(1'b1), .Q(cacheD
		[87]));
	notech_mux2 i_3936(.S(n_59825), .A(n_1406), .B(cacheD[87]), .Z(n_4358)
		);
	notech_reg_set cacheD_reg_88(.CP(n_62424), .D(n_4364), .SD(1'b1), .Q(cacheD
		[88]));
	notech_mux2 i_3944(.S(n_59825), .A(n_1403), .B(cacheD[88]), .Z(n_4364)
		);
	notech_nand2 i_150(.A(fsm[0]), .B(fsm[4]), .Z(n_2014));
	notech_reg_set cacheD_reg_89(.CP(n_62424), .D(n_4370), .SD(1'b1), .Q(cacheD
		[89]));
	notech_mux2 i_3952(.S(n_59825), .A(n_1400), .B(cacheD[89]), .Z(n_4370)
		);
	notech_and2 i_21(.A(axi_RVALID), .B(axi_RLAST), .Z(n_2015));
	notech_reg_set cacheD_reg_90(.CP(n_62424), .D(n_4376), .SD(1'b1), .Q(cacheD
		[90]));
	notech_mux2 i_3960(.S(n_59825), .A(n_1397), .B(cacheD[90]), .Z(n_4376)
		);
	notech_nand3 i_119(.A(fsm[3]), .B(fsm[1]), .C(n_6737), .Z(n_2016));
	notech_reg_set cacheD_reg_91(.CP(n_62424), .D(n_4382), .SD(1'b1), .Q(cacheD
		[91]));
	notech_mux2 i_3968(.S(n_59825), .A(n_1394), .B(cacheD[91]), .Z(n_4382)
		);
	notech_nand2 i_99(.A(n_6738), .B(fsm[0]), .Z(n_2017));
	notech_reg_set cacheD_reg_92(.CP(n_62424), .D(n_4388), .SD(1'b1), .Q(cacheD
		[92]));
	notech_mux2 i_3976(.S(n_59825), .A(n_1391), .B(cacheD[92]), .Z(n_4388)
		);
	notech_reg_set cacheD_reg_93(.CP(n_62424), .D(n_4394), .SD(1'b1), .Q(cacheD
		[93]));
	notech_mux2 i_3984(.S(n_59825), .A(n_1388), .B(cacheD[93]), .Z(n_4394)
		);
	notech_or4 i_154(.A(n_2000), .B(n_2017), .C(read_ack), .D(n_6980), .Z(n_2019
		));
	notech_reg_set cacheD_reg_94(.CP(n_62424), .D(n_4400), .SD(1'b1), .Q(cacheD
		[94]));
	notech_mux2 i_3992(.S(n_59825), .A(n_1385), .B(cacheD[94]), .Z(n_4400)
		);
	notech_nao3 i_57472(.A(n_6737), .B(n_1993), .C(n_2019), .Z(n_2020));
	notech_reg_set cacheD_reg_95(.CP(n_62424), .D(n_4406), .SD(1'b1), .Q(cacheD
		[95]));
	notech_mux2 i_4000(.S(n_59825), .A(n_1382), .B(cacheD[95]), .Z(n_4406)
		);
	notech_ao3 i_53(.A(n_1996), .B(n_2020), .C(n_1742), .Z(n_2021));
	notech_reg_set cacheD_reg_96(.CP(n_62424), .D(n_4412), .SD(1'b1), .Q(cacheD
		[96]));
	notech_mux2 i_4008(.S(n_1375), .A(n_1379), .B(cacheD[96]), .Z(n_4412));
	notech_nor2 i_11(.A(axi_AR[31]), .B(n_6974), .Z(n_2022));
	notech_reg_set cacheD_reg_97(.CP(n_62424), .D(n_4418), .SD(1'b1), .Q(cacheD
		[97]));
	notech_mux2 i_4016(.S(n_1375), .A(n_1373), .B(cacheD[97]), .Z(n_4418));
	notech_and2 i_116(.A(n_967), .B(n_1064), .Z(n_2023));
	notech_reg_set cacheD_reg_98(.CP(n_62424), .D(n_4424), .SD(1'b1), .Q(cacheD
		[98]));
	notech_mux2 i_4024(.S(n_1375), .A(n_1370), .B(cacheD[98]), .Z(n_4424));
	notech_nao3 i_57477(.A(n_6735), .B(n_6738), .C(n_2012), .Z(n_2024));
	notech_reg_set cacheD_reg_99(.CP(n_62424), .D(n_4430), .SD(1'b1), .Q(cacheD
		[99]));
	notech_mux2 i_4032(.S(n_1375), .A(n_1367), .B(cacheD[99]), .Z(n_4430));
	notech_ao4 i_31(.A(n_1998), .B(n_2014), .C(n_2012), .D(n_6630), .Z(n_2025
		));
	notech_reg_set cacheD_reg_100(.CP(n_62424), .D(n_4436), .SD(1'b1), .Q(cacheD
		[100]));
	notech_mux2 i_4040(.S(n_1375), .A(n_1364), .B(cacheD[100]), .Z(n_4436)
		);
	notech_and2 i_12(.A(burst_idx[0]), .B(burst_idx[1]), .Z(n_2026));
	notech_reg_set cacheD_reg_101(.CP(n_62400), .D(n_4442), .SD(1'b1), .Q(cacheD
		[101]));
	notech_mux2 i_4048(.S(n_1375), .A(n_1361), .B(cacheD[101]), .Z(n_4442)
		);
	notech_and3 i_27(.A(burst_idx[0]), .B(burst_idx[1]), .C(burst_idx[2]), .Z
		(n_2027));
	notech_reg_set cacheD_reg_102(.CP(n_62400), .D(n_4448), .SD(1'b1), .Q(cacheD
		[102]));
	notech_mux2 i_4056(.S(n_1375), .A(n_1358), .B(cacheD[102]), .Z(n_4448)
		);
	notech_and4 i_74(.A(burst_idx[0]), .B(burst_idx[1]), .C(burst_idx[2]), .D
		(burst_idx[3]), .Z(n_2028));
	notech_reg_set cacheD_reg_103(.CP(n_62400), .D(n_4454), .SD(1'b1), .Q(cacheD
		[103]));
	notech_mux2 i_4064(.S(n_1375), .A(n_1355), .B(cacheD[103]), .Z(n_4454)
		);
	notech_reg_set cacheD_reg_104(.CP(n_62400), .D(n_4460), .SD(1'b1), .Q(cacheD
		[104]));
	notech_mux2 i_4072(.S(n_1375), .A(n_1352), .B(cacheD[104]), .Z(n_4460)
		);
	notech_nand2 i_51(.A(axi_RVALID), .B(n_61815), .Z(n_2030));
	notech_reg_set cacheD_reg_105(.CP(n_62400), .D(n_4466), .SD(1'b1), .Q(cacheD
		[105]));
	notech_mux2 i_4080(.S(n_1375), .A(n_1349), .B(cacheD[105]), .Z(n_4466)
		);
	notech_reg_set cacheD_reg_106(.CP(n_62400), .D(n_4472), .SD(1'b1), .Q(cacheD
		[106]));
	notech_mux2 i_4088(.S(n_1375), .A(n_1346), .B(cacheD[106]), .Z(n_4472)
		);
	notech_nao3 i_14(.A(fsm[0]), .B(n_6738), .C(n_1998), .Z(n_2032));
	notech_reg_set cacheD_reg_107(.CP(n_62400), .D(n_4478), .SD(1'b1), .Q(cacheD
		[107]));
	notech_mux2 i_4096(.S(n_1375), .A(n_1343), .B(cacheD[107]), .Z(n_4478)
		);
	notech_nao3 i_5780186(.A(n_909), .B(n_908), .C(n_893), .Z(n_2033));
	notech_reg_set cacheD_reg_108(.CP(n_62400), .D(n_4484), .SD(1'b1), .Q(cacheD
		[108]));
	notech_mux2 i_4104(.S(n_1375), .A(n_1340), .B(cacheD[108]), .Z(n_4484)
		);
	notech_reg_set cacheD_reg_109(.CP(n_62400), .D(n_4490), .SD(1'b1), .Q(cacheD
		[109]));
	notech_mux2 i_4112(.S(n_1375), .A(n_1337), .B(cacheD[109]), .Z(n_4490)
		);
	notech_or2 i_344(.A(burst_idx[2]), .B(burst_idx[3]), .Z(n_2035));
	notech_reg_set cacheD_reg_110(.CP(n_62400), .D(n_4496), .SD(1'b1), .Q(cacheD
		[110]));
	notech_mux2 i_4120(.S(n_1375), .A(n_1334), .B(cacheD[110]), .Z(n_4496)
		);
	notech_reg_set cacheD_reg_111(.CP(n_62400), .D(n_4502), .SD(1'b1), .Q(cacheD
		[111]));
	notech_mux2 i_4128(.S(n_1375), .A(n_1331), .B(cacheD[111]), .Z(n_4502)
		);
	notech_reg_set cacheD_reg_112(.CP(n_62400), .D(n_4508), .SD(1'b1), .Q(cacheD
		[112]));
	notech_mux2 i_4136(.S(n_59910), .A(n_1328), .B(cacheD[112]), .Z(n_4508)
		);
	notech_or4 i_46(.A(burst_idx[4]), .B(burst_idx[1]), .C(burst_idx[0]), .D
		(n_2035), .Z(n_2038));
	notech_reg_set cacheD_reg_113(.CP(n_62400), .D(n_4514), .SD(1'b1), .Q(cacheD
		[113]));
	notech_mux2 i_4144(.S(n_59910), .A(n_1325), .B(cacheD[113]), .Z(n_4514)
		);
	notech_reg_set cacheD_reg_114(.CP(n_62400), .D(n_4520), .SD(1'b1), .Q(cacheD
		[114]));
	notech_mux2 i_4152(.S(n_59910), .A(n_1322), .B(cacheD[114]), .Z(n_4520)
		);
	notech_or4 i_78(.A(axi_WREADY), .B(n_2038), .C(n_2033), .D(n_6972), .Z(n_2040
		));
	notech_reg_set cacheD_reg_115(.CP(n_62400), .D(n_4526), .SD(1'b1), .Q(cacheD
		[115]));
	notech_mux2 i_4160(.S(n_59910), .A(n_1319), .B(cacheD[115]), .Z(n_4526)
		);
	notech_reg_set cacheD_reg_116(.CP(n_62400), .D(n_4532), .SD(1'b1), .Q(cacheD
		[116]));
	notech_mux2 i_4168(.S(n_59910), .A(n_1316), .B(cacheD[116]), .Z(n_4532)
		);
	notech_reg_set cacheD_reg_117(.CP(n_62400), .D(n_4538), .SD(1'b1), .Q(cacheD
		[117]));
	notech_mux2 i_4176(.S(n_59910), .A(n_1313), .B(cacheD[117]), .Z(n_4538)
		);
	notech_and4 i_57489(.A(fsm[3]), .B(n_6736), .C(fsm[2]), .D(n_1999), .Z(n_2043
		));
	notech_reg_set cacheD_reg_118(.CP(n_62400), .D(n_4544), .SD(1'b1), .Q(cacheD
		[118]));
	notech_mux2 i_4184(.S(n_59910), .A(n_1310), .B(cacheD[118]), .Z(n_4544)
		);
	notech_and2 i_24(.A(axi_RREADY), .B(axi_RVALID), .Z(n_2044));
	notech_reg_set cacheD_reg_119(.CP(n_62400), .D(n_4550), .SD(1'b1), .Q(cacheD
		[119]));
	notech_mux2 i_4192(.S(n_59910), .A(n_1307), .B(cacheD[119]), .Z(n_4550)
		);
	notech_ao4 i_73(.A(n_6642), .B(n_6625), .C(n_2025), .D(n_6632), .Z(n_2045
		));
	notech_reg_set cacheD_reg_120(.CP(n_62420), .D(n_4556), .SD(1'b1), .Q(cacheD
		[120]));
	notech_mux2 i_4200(.S(n_59910), .A(n_1304), .B(cacheD[120]), .Z(n_4556)
		);
	notech_ao4 i_58(.A(n_6625), .B(n_2044), .C(n_61224), .D(n_2015), .Z(n_2046
		));
	notech_reg_set cacheD_reg_121(.CP(n_62382), .D(n_4562), .SD(1'b1), .Q(cacheD
		[121]));
	notech_mux2 i_4208(.S(n_59910), .A(n_1301), .B(cacheD[121]), .Z(n_4562)
		);
	notech_reg_set cacheD_reg_122(.CP(n_62382), .D(n_4568), .SD(1'b1), .Q(cacheD
		[122]));
	notech_mux2 i_4216(.S(n_59910), .A(n_1298), .B(cacheD[122]), .Z(n_4568)
		);
	notech_reg_set cacheD_reg_123(.CP(n_62382), .D(n_4574), .SD(1'b1), .Q(cacheD
		[123]));
	notech_mux2 i_4224(.S(n_59910), .A(n_1295), .B(cacheD[123]), .Z(n_4574)
		);
	notech_ao4 i_388(.A(code_req), .B(n_6677), .C(read_req), .D(n_6625), .Z(n_2049
		));
	notech_reg_set cacheD_reg_124(.CP(n_62382), .D(n_4580), .SD(1'b1), .Q(cacheD
		[124]));
	notech_mux2 i_4232(.S(n_59910), .A(n_1292), .B(cacheD[124]), .Z(n_4580)
		);
	notech_reg_set cacheD_reg_125(.CP(n_62382), .D(n_4586), .SD(1'b1), .Q(cacheD
		[125]));
	notech_mux2 i_4240(.S(n_59910), .A(n_1289), .B(cacheD[125]), .Z(n_4586)
		);
	notech_reg_set cacheD_reg_126(.CP(n_62382), .D(n_4592), .SD(1'b1), .Q(cacheD
		[126]));
	notech_mux2 i_4248(.S(n_59910), .A(n_1286), .B(cacheD[126]), .Z(n_4592)
		);
	notech_or4 i_42(.A(n_927), .B(n_943), .C(n_942), .D(n_6972), .Z(n_2052)
		);
	notech_reg_set cacheD_reg_127(.CP(n_62382), .D(n_4598), .SD(1'b1), .Q(cacheD
		[127]));
	notech_mux2 i_4256(.S(n_59910), .A(n_1283), .B(cacheD[127]), .Z(n_4598)
		);
	notech_or4 i_126(.A(fsm[2]), .B(n_2019), .C(n_6634), .D(n_2022), .Z(n_2053
		));
	notech_reg_set cacheD_reg_128(.CP(n_62382), .D(n_4604), .SD(1'b1), .Q(cacheD
		[128]));
	notech_mux2 i_4264(.S(n_1277), .A(n_6734), .B(cacheD[128]), .Z(n_4604)
		);
	notech_ao4 i_44(.A(n_2053), .B(n_2052), .C(n_6630), .D(n_2016), .Z(n_2054
		));
	notech_reg_set cacheD_reg_129(.CP(n_62382), .D(n_4610), .SD(1'b1), .Q(cacheD
		[129]));
	notech_mux2 i_4272(.S(n_1277), .A(n_6732), .B(cacheD[129]), .Z(n_4610)
		);
	notech_reg_set cacheD_reg_130(.CP(n_62382), .D(n_4616), .SD(1'b1), .Q(cacheD
		[130]));
	notech_mux2 i_4280(.S(n_1277), .A(n_6731), .B(cacheD[130]), .Z(n_4616)
		);
	notech_reg_set cacheD_reg_131(.CP(n_62382), .D(n_4622), .SD(1'b1), .Q(cacheD
		[131]));
	notech_mux2 i_4288(.S(n_1277), .A(n_6730), .B(cacheD[131]), .Z(n_4622)
		);
	notech_reg_set cacheD_reg_132(.CP(n_62382), .D(n_4628), .SD(1'b1), .Q(cacheD
		[132]));
	notech_mux2 i_4296(.S(n_1277), .A(n_6729), .B(cacheD[132]), .Z(n_4628)
		);
	notech_nand2 i_47(.A(n_2032), .B(n_6675), .Z(n_2058));
	notech_reg_set cacheD_reg_133(.CP(n_62382), .D(n_4634), .SD(1'b1), .Q(cacheD
		[133]));
	notech_mux2 i_4304(.S(n_1277), .A(n_6728), .B(cacheD[133]), .Z(n_4634)
		);
	notech_and3 i_50(.A(n_2032), .B(n_6675), .C(n_6625), .Z(n_2059));
	notech_reg_set cacheD_reg_134(.CP(n_62382), .D(n_4640), .SD(1'b1), .Q(cacheD
		[134]));
	notech_mux2 i_4312(.S(n_1277), .A(n_6727), .B(cacheD[134]), .Z(n_4640)
		);
	notech_and4 i_76(.A(n_2032), .B(n_6675), .C(n_2054), .D(n_6625), .Z(n_2060
		));
	notech_reg_set cacheD_reg_135(.CP(n_62382), .D(n_4646), .SD(1'b1), .Q(cacheD
		[135]));
	notech_mux2 i_4320(.S(n_1277), .A(n_6726), .B(cacheD[135]), .Z(n_4646)
		);
	notech_and2 i_121(.A(n_2060), .B(n_6677), .Z(n_2061));
	notech_reg_set cacheD_reg_136(.CP(n_62382), .D(n_4652), .SD(1'b1), .Q(cacheD
		[136]));
	notech_mux2 i_4328(.S(n_1277), .A(n_6725), .B(cacheD[136]), .Z(n_4652)
		);
	notech_reg_set cacheD_reg_137(.CP(n_62382), .D(n_4658), .SD(1'b1), .Q(cacheD
		[137]));
	notech_mux2 i_4336(.S(n_1277), .A(n_6724), .B(cacheD[137]), .Z(n_4658)
		);
	notech_reg_set cacheD_reg_138(.CP(n_62420), .D(n_4664), .SD(1'b1), .Q(cacheD
		[138]));
	notech_mux2 i_4344(.S(n_1277), .A(n_6723), .B(cacheD[138]), .Z(n_4664)
		);
	notech_and4 i_405(.A(n_2020), .B(n_1208), .C(n_1750), .D(n_1218), .Z(n_2064
		));
	notech_reg_set cacheD_reg_139(.CP(n_62404), .D(n_4670), .SD(1'b1), .Q(cacheD
		[139]));
	notech_mux2 i_4352(.S(n_59930), .A(n_6722), .B(cacheD[139]), .Z(n_4670)
		);
	notech_reg_set cacheD_reg_140(.CP(n_62420), .D(n_4676), .SD(1'b1), .Q(cacheD
		[140]));
	notech_mux2 i_4360(.S(n_59930), .A(n_6721), .B(cacheD[140]), .Z(n_4676)
		);
	notech_reg_set cacheD_reg_141(.CP(n_62420), .D(n_4682), .SD(1'b1), .Q(cacheD
		[141]));
	notech_mux2 i_4368(.S(n_59930), .A(n_6720), .B(cacheD[141]), .Z(n_4682)
		);
	notech_reg_set cacheD_reg_142(.CP(n_62420), .D(n_4688), .SD(1'b1), .Q(cacheD
		[142]));
	notech_mux2 i_4376(.S(n_59930), .A(n_6719), .B(cacheD[142]), .Z(n_4688)
		);
	notech_and4 i_416(.A(n_1750), .B(n_2020), .C(n_1208), .D(n_971), .Z(n_2068
		));
	notech_reg_set cacheD_reg_143(.CP(n_62420), .D(n_4694), .SD(1'b1), .Q(cacheD
		[143]));
	notech_mux2 i_4384(.S(n_59930), .A(n_6718), .B(cacheD[143]), .Z(n_4694)
		);
	notech_reg_set cacheD_reg_144(.CP(n_62420), .D(n_4700), .SD(1'b1), .Q(cacheD
		[144]));
	notech_mux2 i_4392(.S(n_59930), .A(n_6717), .B(cacheD[144]), .Z(n_4700)
		);
	notech_reg_set cacheD_reg_145(.CP(n_62420), .D(n_4706), .SD(1'b1), .Q(cacheD
		[145]));
	notech_mux2 i_4400(.S(n_59930), .A(n_6715), .B(cacheD[145]), .Z(n_4706)
		);
	notech_or2 i_0(.A(n_2032), .B(n_26108), .Z(n_2071));
	notech_reg_set cacheD_reg_146(.CP(n_62420), .D(n_4712), .SD(1'b1), .Q(cacheD
		[146]));
	notech_mux2 i_4408(.S(n_1277), .A(n_27983), .B(cacheD[146]), .Z(n_4712)
		);
	notech_and2 i_49(.A(n_61888), .B(n_1166), .Z(n_2072));
	notech_reg_set cacheD_reg_147(.CP(n_62420), .D(n_4718), .SD(1'b1), .Q(cacheD
		[147]));
	notech_mux2 i_4416(.S(n_59930), .A(n_27988), .B(cacheD[147]), .Z(n_4718)
		);
	notech_or4 i_60(.A(fsm[0]), .B(fsm[4]), .C(n_2012), .D(n_2030), .Z(n_2073
		));
	notech_reg_set cacheD_reg_148(.CP(n_62420), .D(n_4724), .SD(1'b1), .Q(cacheD
		[148]));
	notech_mux2 i_4424(.S(n_59930), .A(n_1224), .B(cacheD[148]), .Z(n_4724)
		);
	notech_ao3 i_71(.A(A4[1]), .B(n_6977), .C(n_2032), .Z(n_2074));
	notech_reg_set cacheD_reg_149(.CP(n_62420), .D(n_4730), .SD(1'b1), .Q(cacheD
		[149]));
	notech_mux2 i_4432(.S(n_59930), .A(n_27998), .B(cacheD[149]), .Z(n_4730)
		);
	notech_nor2 i_35(.A(n_59892), .B(n_6633), .Z(n_2075));
	notech_reg axi_WSTRB_reg_0(.CP(n_62420), .D(n_4736), .CD(n_61814), .Q(axi_WSTRB
		[0]));
	notech_mux2 i_4440(.S(n_61862), .A(n_6741), .B(axi_WSTRB[0]), .Z(n_4736)
		);
	notech_nor2 i_70(.A(A4[1]), .B(n_59921), .Z(n_2076));
	notech_reg axi_WSTRB_reg_1(.CP(n_62420), .D(n_4742), .CD(n_61815), .Q(axi_WSTRB
		[1]));
	notech_mux2 i_4448(.S(n_61862), .A(n_28066), .B(axi_WSTRB[1]), .Z(n_4742
		));
	notech_ao3 i_33(.A(A4[1]), .B(n_59892), .C(n_59921), .Z(n_2077));
	notech_reg axi_WSTRB_reg_2(.CP(n_62420), .D(n_4748), .CD(n_61814), .Q(axi_WSTRB
		[2]));
	notech_mux2 i_4456(.S(n_61862), .A(n_28072), .B(axi_WSTRB[2]), .Z(n_4748
		));
	notech_reg axi_WSTRB_reg_3(.CP(n_62420), .D(n_4754), .CD(n_61814), .Q(axi_WSTRB
		[3]));
	notech_mux2 i_4464(.S(n_61862), .A(n_28078), .B(axi_WSTRB[3]), .Z(n_4754
		));
	notech_reg_set cacheM_reg_0(.CP(n_62420), .D(n_4760), .SD(n_61815), .Q(cacheM
		[0]));
	notech_mux2 i_4472(.S(n_1744), .A(n_1746), .B(cacheM[0]), .Z(n_4760));
	notech_reg_set cacheM_reg_1(.CP(n_62420), .D(n_4766), .SD(n_61815), .Q(cacheM
		[1]));
	notech_mux2 i_4480(.S(n_1744), .A(n_1741), .B(cacheM[1]), .Z(n_4766));
	notech_reg_set cacheM_reg_2(.CP(n_62420), .D(n_4772), .SD(n_61815), .Q(cacheM
		[2]));
	notech_mux2 i_4488(.S(n_1744), .A(n_1739), .B(cacheM[2]), .Z(n_4772));
	notech_reg_set cacheM_reg_3(.CP(n_62382), .D(n_4778), .SD(n_61815), .Q(cacheM
		[3]));
	notech_mux2 i_4496(.S(n_1744), .A(n_1737), .B(cacheM[3]), .Z(n_4778));
	notech_reg_set cacheM_reg_4(.CP(n_62382), .D(n_4784), .SD(n_61815), .Q(cacheM
		[4]));
	notech_mux2 i_4504(.S(n_1744), .A(n_1735), .B(cacheM[4]), .Z(n_4784));
	notech_reg_set cacheM_reg_5(.CP(n_62406), .D(n_4790), .SD(n_61816), .Q(cacheM
		[5]));
	notech_mux2 i_4512(.S(n_1744), .A(n_1733), .B(cacheM[5]), .Z(n_4790));
	notech_reg_set cacheM_reg_6(.CP(n_62406), .D(n_4796), .SD(n_61816), .Q(cacheM
		[6]));
	notech_mux2 i_4520(.S(n_1744), .A(n_1731), .B(cacheM[6]), .Z(n_4796));
	notech_reg_set cacheM_reg_7(.CP(n_62406), .D(n_4802), .SD(n_61816), .Q(cacheM
		[7]));
	notech_mux2 i_4528(.S(n_1744), .A(n_1729), .B(cacheM[7]), .Z(n_4802));
	notech_reg_set cacheM_reg_8(.CP(n_62406), .D(n_4808), .SD(n_61816), .Q(cacheM
		[8]));
	notech_mux2 i_4536(.S(n_1744), .A(n_1727), .B(cacheM[8]), .Z(n_4808));
	notech_reg_set cacheM_reg_9(.CP(n_62406), .D(n_4814), .SD(n_61816), .Q(cacheM
		[9]));
	notech_mux2 i_4544(.S(n_1744), .A(n_1725), .B(cacheM[9]), .Z(n_4814));
	notech_reg_set cacheM_reg_10(.CP(n_62406), .D(n_4820), .SD(n_61816), .Q(cacheM
		[10]));
	notech_mux2 i_4552(.S(n_1744), .A(n_1723), .B(cacheM[10]), .Z(n_4820));
	notech_reg_set cacheM_reg_11(.CP(n_62406), .D(n_4826), .SD(n_61816), .Q(cacheM
		[11]));
	notech_mux2 i_4560(.S(n_1744), .A(n_1721), .B(cacheM[11]), .Z(n_4826));
	notech_reg_set cacheM_reg_12(.CP(n_62406), .D(n_4832), .SD(n_61816), .Q(cacheM
		[12]));
	notech_mux2 i_4568(.S(n_1744), .A(n_1719), .B(cacheM[12]), .Z(n_4832));
	notech_reg_set cacheM_reg_13(.CP(n_62406), .D(n_4838), .SD(n_61816), .Q(cacheM
		[13]));
	notech_mux2 i_4576(.S(n_1744), .A(n_1717), .B(cacheM[13]), .Z(n_4838));
	notech_reg_set cacheM_reg_14(.CP(n_62406), .D(n_4844), .SD(n_61816), .Q(cacheM
		[14]));
	notech_mux2 i_4584(.S(n_1744), .A(n_1715), .B(cacheM[14]), .Z(n_4844));
	notech_reg_set cacheM_reg_15(.CP(n_62406), .D(n_4850), .SD(n_61816), .Q(cacheM
		[15]));
	notech_mux2 i_4592(.S(n_1744), .A(n_1713), .B(cacheM[15]), .Z(n_4850));
	notech_reg_set cacheWEN_reg(.CP(n_62406), .D(n_4856), .SD(n_61816), .Q(cacheWEN
		));
	notech_mux2 i_4600(.S(n_1749), .A(n_1752), .B(cacheWEN), .Z(n_4856));
	notech_reg axi_ARVALID_reg(.CP(n_62406), .D(n_4862), .CD(n_61816), .Q(axi_ARVALID
		));
	notech_mux2 i_4608(.S(n_1755), .A(n_1756), .B(axi_ARVALID), .Z(n_4862)
		);
	notech_reg wf_reg(.CP(n_62406), .D(writeio_req), .CD(n_61816), .Q(wf));
	notech_reg axi_io_AWVALID_reg(.CP(n_62406), .D(n_4870), .CD(n_61816), .Q
		(axi_io_AWVALID));
	notech_mux2 i_4620(.S(n_1758), .A(n_6747), .B(axi_io_AWVALID), .Z(n_4870
		));
	notech_reg axi_io_WVALID_reg(.CP(n_62406), .D(n_4876), .CD(n_61816), .Q(axi_io_WVALID
		));
	notech_mux2 i_4628(.S(n_1760), .A(n_27181), .B(axi_io_WVALID), .Z(n_4876
		));
	notech_reg rf_reg(.CP(n_62406), .D(readio_req), .CD(n_61809), .Q(rf));
	notech_reg axi_io_ARVALID_reg(.CP(n_62406), .D(n_4884), .CD(n_61802), .Q
		(axi_io_ARVALID));
	notech_mux2 i_4640(.S(n_1762), .A(n_6740), .B(axi_io_ARVALID), .Z(n_4884
		));
	notech_reg axi_io_RREADY_reg(.CP(n_62384), .D(n_4890), .CD(n_61802), .Q(axi_io_RREADY
		));
	notech_mux2 i_4648(.S(n_1763), .A(n_28035), .B(axi_io_RREADY), .Z(n_4890
		));
	notech_reg readio_ack_reg(.CP(n_62406), .D(n_4898), .CD(n_61801), .Q(readio_ack
		));
	notech_ao3 i_4657(.A(n_222757064), .B(n_222657063), .C(readio_ack), .Z(n_4898
		));
	notech_reg writeio_ack_reg(.CP(n_62360), .D(n_4902), .CD(n_61802), .Q(writeio_ack
		));
	notech_xor2 i_4664(.A(n_6975), .B(n_1766), .Z(n_4902));
	notech_reg axi_ARSIZE_reg_0(.CP(n_62360), .D(n_4911), .CD(n_61802), .Q(axi_ARSIZE
		[0]));
	notech_and2 i_4674(.A(n_967), .B(axi_ARSIZE[0]), .Z(n_4911));
	notech_reg_set axi_ARSIZE_reg_1(.CP(n_62360), .D(n_4919), .SD(n_61802), 
		.Q(axi_ARSIZE[1]));
	notech_nao3 i_4685(.A(n_967), .B(1'b1), .C(axi_ARSIZE[1]), .Z(n_4919));
	notech_reg axi_ARSIZE_reg_2(.CP(n_62360), .D(n_4923), .CD(n_61802), .Q(axi_ARSIZE
		[2]));
	notech_and2 i_4690(.A(n_967), .B(axi_ARSIZE[2]), .Z(n_4923));
	notech_reg axi_WLAST_reg(.CP(n_62360), .D(n_4926), .CD(n_61802), .Q(axi_WLAST
		));
	notech_mux2 i_4696(.S(n_61862), .A(n_1767), .B(axi_WLAST), .Z(n_4926));
	notech_reg axi_io_AW_reg_0(.CP(n_62360), .D(n_4935), .CD(n_61801), .Q(axi_io_AW
		[0]));
	notech_and2 i_4706(.A(axi_io_AW[0]), .B(n_6748), .Z(n_4935));
	notech_reg axi_io_AW_reg_1(.CP(n_62360), .D(n_4941), .CD(n_61801), .Q(axi_io_AW
		[1]));
	notech_and2 i_4714(.A(n_6748), .B(axi_io_AW[1]), .Z(n_4941));
	notech_or4 i_604(.A(burst_idx[2]), .B(burst_idx[3]), .C(burst_idx[4]), .D
		(n_6635), .Z(n_2109));
	notech_reg axi_io_AW_reg_2(.CP(n_62360), .D(n_4944), .CD(n_61801), .Q(axi_io_AW
		[2]));
	notech_mux2 i_4720(.S(\nbus_11686[0] ), .A(axi_io_AW[2]), .B(io_add[0]),
		 .Z(n_4944));
	notech_reg axi_io_AW_reg_3(.CP(n_62360), .D(n_4950), .CD(n_61801), .Q(axi_io_AW
		[3]));
	notech_mux2 i_4728(.S(\nbus_11686[0] ), .A(axi_io_AW[3]), .B(io_add[1]),
		 .Z(n_4950));
	notech_reg axi_io_AW_reg_4(.CP(n_62360), .D(n_4956), .CD(n_61801), .Q(axi_io_AW
		[4]));
	notech_mux2 i_4736(.S(\nbus_11686[0] ), .A(axi_io_AW[4]), .B(io_add[2]),
		 .Z(n_4956));
	notech_reg axi_io_AW_reg_5(.CP(n_62360), .D(n_4962), .CD(n_61801), .Q(axi_io_AW
		[5]));
	notech_mux2 i_4744(.S(\nbus_11686[0] ), .A(axi_io_AW[5]), .B(io_add[3]),
		 .Z(n_4962));
	notech_reg axi_io_AW_reg_6(.CP(n_62360), .D(n_4968), .CD(n_61801), .Q(axi_io_AW
		[6]));
	notech_mux2 i_4752(.S(\nbus_11686[0] ), .A(axi_io_AW[6]), .B(io_add[4]),
		 .Z(n_4968));
	notech_reg axi_io_AW_reg_7(.CP(n_62360), .D(n_4974), .CD(n_61801), .Q(axi_io_AW
		[7]));
	notech_mux2 i_4760(.S(\nbus_11686[0] ), .A(axi_io_AW[7]), .B(io_add[5]),
		 .Z(n_4974));
	notech_reg axi_io_AW_reg_8(.CP(n_62360), .D(n_4980), .CD(n_61802), .Q(axi_io_AW
		[8]));
	notech_mux2 i_4768(.S(n_61206), .A(axi_io_AW[8]), .B(io_add[6]), .Z(n_4980
		));
	notech_reg axi_io_AW_reg_9(.CP(n_62360), .D(n_4986), .CD(n_61803), .Q(axi_io_AW
		[9]));
	notech_mux2 i_4776(.S(n_61206), .A(axi_io_AW[9]), .B(io_add[7]), .Z(n_4986
		));
	notech_reg axi_io_AW_reg_10(.CP(n_62360), .D(n_4992), .CD(n_61803), .Q(axi_io_AW
		[10]));
	notech_mux2 i_4784(.S(n_61206), .A(axi_io_AW[10]), .B(io_add[8]), .Z(n_4992
		));
	notech_reg axi_io_AW_reg_11(.CP(n_62360), .D(n_4998), .CD(n_61803), .Q(axi_io_AW
		[11]));
	notech_mux2 i_4792(.S(n_61206), .A(axi_io_AW[11]), .B(io_add[9]), .Z(n_4998
		));
	notech_reg axi_io_AW_reg_12(.CP(n_62360), .D(n_5004), .CD(n_61803), .Q(axi_io_AW
		[12]));
	notech_mux2 i_4800(.S(n_61206), .A(axi_io_AW[12]), .B(io_add[10]), .Z(n_5004
		));
	notech_reg axi_io_AW_reg_13(.CP(n_62360), .D(n_5010), .CD(n_61803), .Q(axi_io_AW
		[13]));
	notech_mux2 i_4808(.S(n_61206), .A(axi_io_AW[13]), .B(io_add[11]), .Z(n_5010
		));
	notech_reg axi_io_AW_reg_14(.CP(n_62368), .D(n_5016), .CD(n_61803), .Q(axi_io_AW
		[14]));
	notech_mux2 i_4816(.S(\nbus_11686[0] ), .A(axi_io_AW[14]), .B(io_add[12]
		), .Z(n_5016));
	notech_reg axi_io_AW_reg_15(.CP(n_62352), .D(n_5022), .CD(n_61803), .Q(axi_io_AW
		[15]));
	notech_mux2 i_4824(.S(\nbus_11686[0] ), .A(axi_io_AW[15]), .B(io_add[13]
		), .Z(n_5022));
	notech_reg axi_io_AW_reg_16(.CP(n_62352), .D(n_5028), .CD(n_61803), .Q(axi_io_AW
		[16]));
	notech_mux2 i_4832(.S(\nbus_11686[0] ), .A(axi_io_AW[16]), .B(io_add[14]
		), .Z(n_5028));
	notech_reg axi_io_AW_reg_17(.CP(n_62352), .D(n_5034), .CD(n_61802), .Q(axi_io_AW
		[17]));
	notech_mux2 i_4840(.S(\nbus_11686[0] ), .A(axi_io_AW[17]), .B(io_add[15]
		), .Z(n_5034));
	notech_reg axi_io_AW_reg_18(.CP(n_62352), .D(n_5043), .CD(n_61802), .Q(axi_io_AW
		[18]));
	notech_and2 i_4850(.A(axi_io_AW[18]), .B(n_6748), .Z(n_5043));
	notech_reg axi_io_AW_reg_19(.CP(n_62352), .D(n_5049), .CD(n_61802), .Q(axi_io_AW
		[19]));
	notech_and2 i_4858(.A(axi_io_AW[19]), .B(n_6748), .Z(n_5049));
	notech_reg axi_io_AW_reg_20(.CP(n_62352), .D(n_5055), .CD(n_61802), .Q(axi_io_AW
		[20]));
	notech_and2 i_4866(.A(axi_io_AW[20]), .B(n_6748), .Z(n_5055));
	notech_reg axi_io_AW_reg_21(.CP(n_62352), .D(n_5061), .CD(n_61802), .Q(axi_io_AW
		[21]));
	notech_and2 i_4874(.A(axi_io_AW[21]), .B(n_6748), .Z(n_5061));
	notech_reg axi_io_AW_reg_22(.CP(n_62352), .D(n_5067), .CD(n_61803), .Q(axi_io_AW
		[22]));
	notech_and2 i_4882(.A(axi_io_AW[22]), .B(n_6748), .Z(n_5067));
	notech_reg axi_io_AW_reg_23(.CP(n_62352), .D(n_5073), .CD(n_61802), .Q(axi_io_AW
		[23]));
	notech_and2 i_4890(.A(axi_io_AW[23]), .B(n_6748), .Z(n_5073));
	notech_reg axi_io_AW_reg_24(.CP(n_62352), .D(n_5079), .CD(n_61802), .Q(axi_io_AW
		[24]));
	notech_and2 i_4898(.A(axi_io_AW[24]), .B(n_6748), .Z(n_5079));
	notech_reg axi_io_AW_reg_25(.CP(n_62352), .D(n_5085), .CD(n_61799), .Q(axi_io_AW
		[25]));
	notech_and2 i_4906(.A(axi_io_AW[25]), .B(n_6748), .Z(n_5085));
	notech_reg axi_io_AW_reg_26(.CP(n_62352), .D(n_5091), .CD(n_61799), .Q(axi_io_AW
		[26]));
	notech_and2 i_4914(.A(axi_io_AW[26]), .B(n_6748), .Z(n_5091));
	notech_reg axi_io_AW_reg_27(.CP(n_62352), .D(n_5097), .CD(n_61799), .Q(axi_io_AW
		[27]));
	notech_and2 i_4922(.A(axi_io_AW[27]), .B(n_6748), .Z(n_5097));
	notech_reg axi_io_AW_reg_28(.CP(n_62352), .D(n_5103), .CD(n_61799), .Q(axi_io_AW
		[28]));
	notech_and2 i_4930(.A(axi_io_AW[28]), .B(n_6748), .Z(n_5103));
	notech_reg axi_io_AW_reg_29(.CP(n_62352), .D(n_5109), .CD(n_61800), .Q(axi_io_AW
		[29]));
	notech_and2 i_4938(.A(axi_io_AW[29]), .B(n_6748), .Z(n_5109));
	notech_reg axi_io_AW_reg_30(.CP(n_62372), .D(n_5115), .CD(n_61800), .Q(axi_io_AW
		[30]));
	notech_and2 i_4946(.A(axi_io_AW[30]), .B(n_6748), .Z(n_5115));
	notech_reg axi_io_AW_reg_31(.CP(n_62372), .D(n_5121), .CD(n_61799), .Q(axi_io_AW
		[31]));
	notech_and2 i_4954(.A(axi_io_AW[31]), .B(n_6748), .Z(n_5121));
	notech_reg axi_ARLEN_reg_0(.CP(n_62372), .D(n_5124), .CD(n_61799), .Q(axi_ARLEN
		[0]));
	notech_mux2 i_4960(.S(n_61246), .A(n_6637), .B(axi_ARLEN[0]), .Z(n_5124)
		);
	notech_reg axi_ARLEN_reg_1(.CP(n_62372), .D(n_5130), .CD(n_61799), .Q(axi_ARLEN
		[1]));
	notech_mux2 i_4968(.S(n_61246), .A(n_6637), .B(axi_ARLEN[1]), .Z(n_5130)
		);
	notech_reg axi_ARLEN_reg_2(.CP(n_62372), .D(n_5139), .CD(n_61799), .Q(axi_ARLEN
		[2]));
	notech_and4 i_4978(.A(n_967), .B(n_1064), .C(axi_ARLEN[2]), .D(n_971), .Z
		(n_5139));
	notech_or4 i_735(.A(burst_idx[4]), .B(n_2035), .C(burst_idx[0]), .D(n_6714
		), .Z(n_214256979));
	notech_reg axi_ARLEN_reg_3(.CP(n_62372), .D(n_5145), .CD(n_61799), .Q(axi_ARLEN
		[3]));
	notech_and4 i_4986(.A(n_967), .B(n_1064), .C(axi_ARLEN[3]), .D(n_971), .Z
		(n_5145));
	notech_reg axi_ARLEN_reg_4(.CP(n_62372), .D(n_5151), .CD(n_61799), .Q(axi_ARLEN
		[4]));
	notech_and4 i_4994(.A(n_61959), .B(n_1064), .C(axi_ARLEN[4]), .D(n_971),
		 .Z(n_5151));
	notech_or4 i_34(.A(n_26108), .B(n_2032), .C(A4[1]), .D(n_59892), .Z(n_214456981
		));
	notech_reg axi_ARLEN_reg_5(.CP(n_62372), .D(n_5157), .CD(n_61799), .Q(axi_ARLEN
		[5]));
	notech_and4 i_5002(.A(n_61959), .B(n_1064), .C(axi_ARLEN[5]), .D(n_971),
		 .Z(n_5157));
	notech_nand2 i_32(.A(n_59892), .B(n_59853), .Z(n_214556982));
	notech_reg axi_ARLEN_reg_6(.CP(n_62372), .D(n_5163), .CD(n_61799), .Q(axi_ARLEN
		[6]));
	notech_and4 i_5010(.A(n_61959), .B(n_1064), .C(axi_ARLEN[6]), .D(n_971),
		 .Z(n_5163));
	notech_reg axi_ARLEN_reg_7(.CP(n_62372), .D(n_5169), .CD(n_61799), .Q(axi_ARLEN
		[7]));
	notech_and4 i_5018(.A(n_61959), .B(n_1064), .C(axi_ARLEN[7]), .D(n_971),
		 .Z(n_5169));
	notech_reg axi_io_AR_reg_0(.CP(n_62372), .D(n_5175), .CD(n_61799), .Q(axi_io_AR
		[0]));
	notech_and2 i_5026(.A(axi_io_AR[0]), .B(n_6742), .Z(n_5175));
	notech_reg axi_io_AR_reg_1(.CP(n_62372), .D(n_5181), .CD(n_61800), .Q(axi_io_AR
		[1]));
	notech_and2 i_5034(.A(n_6742), .B(axi_io_AR[1]), .Z(n_5181));
	notech_reg axi_io_AR_reg_2(.CP(n_62372), .D(n_5184), .CD(n_61800), .Q(axi_io_AR
		[2]));
	notech_mux2 i_5040(.S(\nbus_11699[0] ), .A(axi_io_AR[2]), .B(io_add[0]),
		 .Z(n_5184));
	notech_reg axi_io_AR_reg_3(.CP(n_62372), .D(n_5190), .CD(n_61801), .Q(axi_io_AR
		[3]));
	notech_mux2 i_5048(.S(\nbus_11699[0] ), .A(axi_io_AR[3]), .B(io_add[1]),
		 .Z(n_5190));
	notech_reg axi_io_AR_reg_4(.CP(n_62372), .D(n_5196), .CD(n_61800), .Q(axi_io_AR
		[4]));
	notech_mux2 i_5056(.S(\nbus_11699[0] ), .A(axi_io_AR[4]), .B(io_add[2]),
		 .Z(n_5196));
	notech_reg axi_io_AR_reg_5(.CP(n_62372), .D(n_5202), .CD(n_61800), .Q(axi_io_AR
		[5]));
	notech_mux2 i_5064(.S(\nbus_11699[0] ), .A(axi_io_AR[5]), .B(io_add[3]),
		 .Z(n_5202));
	notech_reg axi_io_AR_reg_6(.CP(n_62372), .D(n_5208), .CD(n_61801), .Q(axi_io_AR
		[6]));
	notech_mux2 i_5072(.S(\nbus_11699[0] ), .A(axi_io_AR[6]), .B(io_add[4]),
		 .Z(n_5208));
	notech_reg axi_io_AR_reg_7(.CP(n_62372), .D(n_5214), .CD(n_61801), .Q(axi_io_AR
		[7]));
	notech_mux2 i_5080(.S(\nbus_11699[0] ), .A(axi_io_AR[7]), .B(io_add[5]),
		 .Z(n_5214));
	notech_reg axi_io_AR_reg_8(.CP(n_62372), .D(n_5220), .CD(n_61801), .Q(axi_io_AR
		[8]));
	notech_mux2 i_5088(.S(\nbus_11699[0] ), .A(axi_io_AR[8]), .B(io_add[6]),
		 .Z(n_5220));
	notech_reg axi_io_AR_reg_9(.CP(n_62370), .D(n_5226), .CD(n_61801), .Q(axi_io_AR
		[9]));
	notech_mux2 i_5096(.S(\nbus_11699[0] ), .A(axi_io_AR[9]), .B(io_add[7]),
		 .Z(n_5226));
	notech_reg axi_io_AR_reg_10(.CP(n_62370), .D(n_5232), .CD(n_61800), .Q(axi_io_AR
		[10]));
	notech_mux2 i_5104(.S(\nbus_11699[0] ), .A(axi_io_AR[10]), .B(io_add[8])
		, .Z(n_5232));
	notech_reg axi_io_AR_reg_11(.CP(n_62396), .D(n_5238), .CD(n_61800), .Q(axi_io_AR
		[11]));
	notech_mux2 i_5112(.S(\nbus_11699[0] ), .A(axi_io_AR[11]), .B(io_add[9])
		, .Z(n_5238));
	notech_reg axi_io_AR_reg_12(.CP(n_62396), .D(n_5244), .CD(n_61800), .Q(axi_io_AR
		[12]));
	notech_mux2 i_5120(.S(\nbus_11699[0] ), .A(axi_io_AR[12]), .B(io_add[10]
		), .Z(n_5244));
	notech_reg axi_io_AR_reg_13(.CP(n_62396), .D(n_5250), .CD(n_61800), .Q(axi_io_AR
		[13]));
	notech_mux2 i_5128(.S(\nbus_11699[0] ), .A(axi_io_AR[13]), .B(io_add[11]
		), .Z(n_5250));
	notech_reg axi_io_AR_reg_14(.CP(n_62396), .D(n_5256), .CD(n_61800), .Q(axi_io_AR
		[14]));
	notech_mux2 i_5136(.S(\nbus_11699[0] ), .A(axi_io_AR[14]), .B(io_add[12]
		), .Z(n_5256));
	notech_reg axi_io_AR_reg_15(.CP(n_62396), .D(n_5262), .CD(n_61800), .Q(axi_io_AR
		[15]));
	notech_mux2 i_5144(.S(\nbus_11699[0] ), .A(axi_io_AR[15]), .B(io_add[13]
		), .Z(n_5262));
	notech_reg axi_io_AR_reg_16(.CP(n_62396), .D(n_5268), .CD(n_61800), .Q(axi_io_AR
		[16]));
	notech_mux2 i_5152(.S(\nbus_11699[0] ), .A(axi_io_AR[16]), .B(io_add[14]
		), .Z(n_5268));
	notech_reg axi_io_AR_reg_17(.CP(n_62396), .D(n_5274), .CD(n_61800), .Q(axi_io_AR
		[17]));
	notech_mux2 i_5160(.S(\nbus_11699[0] ), .A(axi_io_AR[17]), .B(io_add[15]
		), .Z(n_5274));
	notech_reg axi_io_AR_reg_18(.CP(n_62396), .D(n_5283), .CD(n_61803), .Q(axi_io_AR
		[18]));
	notech_and2 i_5170(.A(axi_io_AR[18]), .B(n_6742), .Z(n_5283));
	notech_reg axi_io_AR_reg_19(.CP(n_62396), .D(n_5289), .CD(n_61807), .Q(axi_io_AR
		[19]));
	notech_and2 i_5178(.A(axi_io_AR[19]), .B(n_6742), .Z(n_5289));
	notech_reg axi_io_AR_reg_20(.CP(n_62396), .D(n_5295), .CD(n_61807), .Q(axi_io_AR
		[20]));
	notech_and2 i_5186(.A(axi_io_AR[20]), .B(n_6742), .Z(n_5295));
	notech_reg axi_io_AR_reg_21(.CP(n_62396), .D(n_5301), .CD(n_61807), .Q(axi_io_AR
		[21]));
	notech_and2 i_5194(.A(axi_io_AR[21]), .B(n_6742), .Z(n_5301));
	notech_reg axi_io_AR_reg_22(.CP(n_62396), .D(n_5307), .CD(n_61807), .Q(axi_io_AR
		[22]));
	notech_and2 i_5202(.A(axi_io_AR[22]), .B(n_6742), .Z(n_5307));
	notech_reg axi_io_AR_reg_23(.CP(n_62396), .D(n_5313), .CD(n_61807), .Q(axi_io_AR
		[23]));
	notech_and2 i_5210(.A(axi_io_AR[23]), .B(n_6742), .Z(n_5313));
	notech_reg axi_io_AR_reg_24(.CP(n_62396), .D(n_5319), .CD(n_61807), .Q(axi_io_AR
		[24]));
	notech_and2 i_5218(.A(axi_io_AR[24]), .B(n_6742), .Z(n_5319));
	notech_reg axi_io_AR_reg_25(.CP(n_62396), .D(n_5325), .CD(n_61807), .Q(axi_io_AR
		[25]));
	notech_and2 i_5226(.A(axi_io_AR[25]), .B(n_6742), .Z(n_5325));
	notech_reg axi_io_AR_reg_26(.CP(n_62396), .D(n_5331), .CD(n_61807), .Q(axi_io_AR
		[26]));
	notech_and2 i_5234(.A(axi_io_AR[26]), .B(n_6742), .Z(n_5331));
	notech_reg axi_io_AR_reg_27(.CP(n_62396), .D(n_5337), .CD(n_61807), .Q(axi_io_AR
		[27]));
	notech_and2 i_5242(.A(axi_io_AR[27]), .B(n_6742), .Z(n_5337));
	notech_reg axi_io_AR_reg_28(.CP(n_62396), .D(n_5343), .CD(n_61807), .Q(axi_io_AR
		[28]));
	notech_and2 i_5250(.A(axi_io_AR[28]), .B(n_6742), .Z(n_5343));
	notech_reg axi_io_AR_reg_29(.CP(n_62370), .D(n_5349), .CD(n_61806), .Q(axi_io_AR
		[29]));
	notech_and2 i_5258(.A(axi_io_AR[29]), .B(n_6742), .Z(n_5349));
	notech_or4 i_866(.A(burst_idx[4]), .B(n_2035), .C(burst_idx[1]), .D(n_6712
		), .Z(n_217757014));
	notech_reg axi_io_AR_reg_30(.CP(n_62370), .D(n_5355), .CD(n_61807), .Q(axi_io_AR
		[30]));
	notech_and2 i_5266(.A(axi_io_AR[30]), .B(n_6742), .Z(n_5355));
	notech_reg axi_io_AR_reg_31(.CP(n_62370), .D(n_5361), .CD(n_61807), .Q(axi_io_AR
		[31]));
	notech_and2 i_5274(.A(axi_io_AR[31]), .B(n_6742), .Z(n_5361));
	notech_reg_set readio_data_reg_0(.CP(n_62370), .D(n_5364), .SD(1'b1), .Q
		(readio_data[0]));
	notech_mux2 i_5280(.S(\nbus_11696[0] ), .A(readio_data[0]), .B(axi_io_R[
		0]), .Z(n_5364));
	notech_reg_set readio_data_reg_1(.CP(n_62370), .D(n_5370), .SD(1'b1), .Q
		(readio_data[1]));
	notech_mux2 i_5288(.S(\nbus_11696[0] ), .A(readio_data[1]), .B(axi_io_R[
		1]), .Z(n_5370));
	notech_reg_set readio_data_reg_2(.CP(n_62370), .D(n_5376), .SD(1'b1), .Q
		(readio_data[2]));
	notech_mux2 i_5296(.S(\nbus_11696[0] ), .A(readio_data[2]), .B(axi_io_R[
		2]), .Z(n_5376));
	notech_reg_set readio_data_reg_3(.CP(n_62370), .D(n_5382), .SD(1'b1), .Q
		(readio_data[3]));
	notech_mux2 i_5304(.S(\nbus_11696[0] ), .A(readio_data[3]), .B(axi_io_R[
		3]), .Z(n_5382));
	notech_reg_set readio_data_reg_4(.CP(n_62370), .D(n_5388), .SD(1'b1), .Q
		(readio_data[4]));
	notech_mux2 i_5312(.S(\nbus_11696[0] ), .A(readio_data[4]), .B(axi_io_R[
		4]), .Z(n_5388));
	notech_reg_set readio_data_reg_5(.CP(n_62370), .D(n_5394), .SD(1'b1), .Q
		(readio_data[5]));
	notech_mux2 i_5320(.S(\nbus_11696[0] ), .A(readio_data[5]), .B(axi_io_R[
		5]), .Z(n_5394));
	notech_reg_set readio_data_reg_6(.CP(n_62370), .D(n_5400), .SD(1'b1), .Q
		(readio_data[6]));
	notech_mux2 i_5328(.S(\nbus_11696[0] ), .A(readio_data[6]), .B(axi_io_R[
		6]), .Z(n_5400));
	notech_reg_set readio_data_reg_7(.CP(n_62370), .D(n_5406), .SD(1'b1), .Q
		(readio_data[7]));
	notech_mux2 i_5336(.S(\nbus_11696[0] ), .A(readio_data[7]), .B(axi_io_R[
		7]), .Z(n_5406));
	notech_reg_set readio_data_reg_8(.CP(n_62370), .D(n_5412), .SD(1'b1), .Q
		(readio_data[8]));
	notech_mux2 i_5344(.S(\nbus_11696[0] ), .A(readio_data[8]), .B(axi_io_R[
		8]), .Z(n_5412));
	notech_reg_set readio_data_reg_9(.CP(n_62370), .D(n_5418), .SD(1'b1), .Q
		(readio_data[9]));
	notech_mux2 i_5352(.S(\nbus_11696[0] ), .A(readio_data[9]), .B(axi_io_R[
		9]), .Z(n_5418));
	notech_reg_set readio_data_reg_10(.CP(n_62370), .D(n_5424), .SD(1'b1), .Q
		(readio_data[10]));
	notech_mux2 i_5360(.S(\nbus_11696[0] ), .A(readio_data[10]), .B(axi_io_R
		[10]), .Z(n_5424));
	notech_reg_set readio_data_reg_11(.CP(n_62370), .D(n_5430), .SD(1'b1), .Q
		(readio_data[11]));
	notech_mux2 i_5368(.S(\nbus_11696[0] ), .A(readio_data[11]), .B(axi_io_R
		[11]), .Z(n_5430));
	notech_reg_set readio_data_reg_12(.CP(n_62396), .D(n_5436), .SD(1'b1), .Q
		(readio_data[12]));
	notech_mux2 i_5376(.S(\nbus_11696[0] ), .A(readio_data[12]), .B(axi_io_R
		[12]), .Z(n_5436));
	notech_reg_set readio_data_reg_13(.CP(n_62392), .D(n_5442), .SD(1'b1), .Q
		(readio_data[13]));
	notech_mux2 i_5384(.S(\nbus_11696[0] ), .A(readio_data[13]), .B(axi_io_R
		[13]), .Z(n_5442));
	notech_reg_set readio_data_reg_14(.CP(n_62368), .D(n_5448), .SD(1'b1), .Q
		(readio_data[14]));
	notech_mux2 i_5392(.S(\nbus_11696[0] ), .A(readio_data[14]), .B(axi_io_R
		[14]), .Z(n_5448));
	notech_reg_set readio_data_reg_15(.CP(n_62392), .D(n_5454), .SD(1'b1), .Q
		(readio_data[15]));
	notech_mux2 i_5400(.S(\nbus_11696[0] ), .A(readio_data[15]), .B(axi_io_R
		[15]), .Z(n_5454));
	notech_reg_set readio_data_reg_16(.CP(n_62392), .D(n_5460), .SD(1'b1), .Q
		(readio_data[16]));
	notech_mux2 i_5408(.S(n_54994), .A(readio_data[16]), .B(axi_io_R[16]), .Z
		(n_5460));
	notech_reg_set readio_data_reg_17(.CP(n_62392), .D(n_5466), .SD(1'b1), .Q
		(readio_data[17]));
	notech_mux2 i_5416(.S(n_54994), .A(readio_data[17]), .B(axi_io_R[17]), .Z
		(n_5466));
	notech_reg_set readio_data_reg_18(.CP(n_62392), .D(n_5472), .SD(1'b1), .Q
		(readio_data[18]));
	notech_mux2 i_5424(.S(n_54994), .A(readio_data[18]), .B(axi_io_R[18]), .Z
		(n_5472));
	notech_reg_set readio_data_reg_19(.CP(n_62392), .D(n_5478), .SD(1'b1), .Q
		(readio_data[19]));
	notech_mux2 i_5432(.S(n_54994), .A(readio_data[19]), .B(axi_io_R[19]), .Z
		(n_5478));
	notech_reg_set readio_data_reg_20(.CP(n_62392), .D(n_5484), .SD(1'b1), .Q
		(readio_data[20]));
	notech_mux2 i_5440(.S(n_54994), .A(readio_data[20]), .B(axi_io_R[20]), .Z
		(n_5484));
	notech_reg_set readio_data_reg_21(.CP(n_62392), .D(n_5490), .SD(1'b1), .Q
		(readio_data[21]));
	notech_mux2 i_5448(.S(n_54994), .A(readio_data[21]), .B(axi_io_R[21]), .Z
		(n_5490));
	notech_reg_set readio_data_reg_22(.CP(n_62392), .D(n_5496), .SD(1'b1), .Q
		(readio_data[22]));
	notech_mux2 i_5456(.S(n_54994), .A(readio_data[22]), .B(axi_io_R[22]), .Z
		(n_5496));
	notech_reg_set readio_data_reg_23(.CP(n_62392), .D(n_5502), .SD(1'b1), .Q
		(readio_data[23]));
	notech_mux2 i_5464(.S(n_54994), .A(readio_data[23]), .B(axi_io_R[23]), .Z
		(n_5502));
	notech_reg_set readio_data_reg_24(.CP(n_62392), .D(n_5508), .SD(1'b1), .Q
		(readio_data[24]));
	notech_mux2 i_5472(.S(n_54994), .A(readio_data[24]), .B(axi_io_R[24]), .Z
		(n_5508));
	notech_reg_set readio_data_reg_25(.CP(n_62392), .D(n_5514), .SD(1'b1), .Q
		(readio_data[25]));
	notech_mux2 i_5480(.S(n_54994), .A(readio_data[25]), .B(axi_io_R[25]), .Z
		(n_5514));
	notech_reg_set readio_data_reg_26(.CP(n_62392), .D(n_5520), .SD(1'b1), .Q
		(readio_data[26]));
	notech_mux2 i_5488(.S(n_54994), .A(readio_data[26]), .B(axi_io_R[26]), .Z
		(n_5520));
	notech_reg_set readio_data_reg_27(.CP(n_62392), .D(n_5526), .SD(1'b1), .Q
		(readio_data[27]));
	notech_mux2 i_5496(.S(n_54994), .A(readio_data[27]), .B(axi_io_R[27]), .Z
		(n_5526));
	notech_reg_set readio_data_reg_28(.CP(n_62392), .D(n_5532), .SD(1'b1), .Q
		(readio_data[28]));
	notech_mux2 i_5504(.S(n_54994), .A(readio_data[28]), .B(axi_io_R[28]), .Z
		(n_5532));
	notech_reg_set readio_data_reg_29(.CP(n_62392), .D(n_5538), .SD(1'b1), .Q
		(readio_data[29]));
	notech_mux2 i_5512(.S(n_54994), .A(readio_data[29]), .B(axi_io_R[29]), .Z
		(n_5538));
	notech_reg_set readio_data_reg_30(.CP(n_62414), .D(n_5544), .SD(1'b1), .Q
		(readio_data[30]));
	notech_mux2 i_5520(.S(n_54994), .A(readio_data[30]), .B(axi_io_R[30]), .Z
		(n_5544));
	notech_reg_set readio_data_reg_31(.CP(n_62414), .D(n_5550), .SD(1'b1), .Q
		(readio_data[31]));
	notech_mux2 i_5528(.S(n_54994), .A(readio_data[31]), .B(axi_io_R[31]), .Z
		(n_5550));
	notech_reg axi_AWLEN_reg_0(.CP(n_62414), .D(n_5559), .CD(n_61807), .Q(axi_AWLEN
		[0]));
	notech_and4 i_5538(.A(n_61959), .B(n_61873), .C(n_61888), .D(axi_AWLEN[0
		]), .Z(n_5559));
	notech_ao3 i_1016(.A(n_2020), .B(n_1711), .C(n_1742), .Z(n_221257049));
	notech_reg axi_AWLEN_reg_1(.CP(n_62414), .D(n_5565), .CD(n_61807), .Q(axi_AWLEN
		[1]));
	notech_and4 i_5546(.A(n_61959), .B(n_61873), .C(n_61888), .D(axi_AWLEN[1
		]), .Z(n_5565));
	notech_reg axi_AWLEN_reg_2(.CP(n_62414), .D(n_5571), .CD(n_61807), .Q(axi_AWLEN
		[2]));
	notech_and4 i_5554(.A(n_61959), .B(n_61873), .C(n_61888), .D(axi_AWLEN[2
		]), .Z(n_5571));
	notech_reg axi_AWLEN_reg_3(.CP(n_62414), .D(n_5577), .CD(n_61808), .Q(axi_AWLEN
		[3]));
	notech_and4 i_5562(.A(n_61959), .B(n_61873), .C(n_61888), .D(axi_AWLEN[3
		]), .Z(n_5577));
	notech_ao3 i_118(.A(n_1996), .B(n_972), .C(n_1742), .Z(n_221557052));
	notech_reg axi_AWLEN_reg_4(.CP(n_62414), .D(n_5583), .CD(n_61808), .Q(axi_AWLEN
		[4]));
	notech_and4 i_5570(.A(n_61959), .B(n_61873), .C(n_61888), .D(axi_AWLEN[4
		]), .Z(n_5583));
	notech_ao4 i_1058(.A(n_6675), .B(n_2033), .C(n_2017), .D(n_2012), .Z(n_221657053
		));
	notech_reg axi_AWLEN_reg_5(.CP(n_62414), .D(n_5589), .CD(n_61808), .Q(axi_AWLEN
		[5]));
	notech_and4 i_5578(.A(n_61959), .B(n_28023), .C(n_61888), .D(axi_AWLEN[5
		]), .Z(n_5589));
	notech_reg axi_AWLEN_reg_6(.CP(n_62414), .D(n_5595), .CD(n_61808), .Q(axi_AWLEN
		[6]));
	notech_and4 i_5586(.A(n_967), .B(n_61873), .C(n_61888), .D(axi_AWLEN[6])
		, .Z(n_5595));
	notech_reg axi_AWLEN_reg_7(.CP(n_62414), .D(n_5601), .CD(n_61808), .Q(axi_AWLEN
		[7]));
	notech_and4 i_5594(.A(n_61959), .B(n_61873), .C(n_61888), .D(axi_AWLEN[7
		]), .Z(n_5601));
	notech_ao4 i_1063(.A(n_2032), .B(n_6631), .C(n_2017), .D(n_2012), .Z(n_221957056
		));
	notech_reg_set axi_AWBURST_reg_0(.CP(n_62414), .D(n_5609), .SD(n_61809),
		 .Q(axi_AWBURST[0]));
	notech_nao3 i_5605(.A(n_61959), .B(1'b1), .C(axi_AWBURST[0]), .Z(n_5609)
		);
	notech_reg axi_AWBURST_reg_1(.CP(n_62414), .D(n_5613), .CD(n_61809), .Q(axi_AWBURST
		[1]));
	notech_and2 i_5610(.A(n_61959), .B(axi_AWBURST[1]), .Z(n_5613));
	notech_reg_set code_data_reg_0(.CP(n_62414), .D(n_5616), .SD(1'b1), .Q(\nbus_14527[0] 
		));
	notech_mux2 i_5616(.S(n_6743), .A(n_60807), .B(axi_R[0]), .Z(n_5616));
	notech_or2 i_57(.A(readio_ack), .B(writeio_ack), .Z(n_222257059));
	notech_reg_set code_data_reg_1(.CP(n_62414), .D(n_5622), .SD(1'b1), .Q(code_data
		[1]));
	notech_mux2 i_5624(.S(n_6743), .A(code_data[1]), .B(axi_R[1]), .Z(n_5622
		));
	notech_nao3 i_120(.A(n_6975), .B(n_6747), .C(readio_ack), .Z(n_222357060
		));
	notech_reg_set code_data_reg_2(.CP(n_62414), .D(n_5628), .SD(1'b1), .Q(code_data
		[2]));
	notech_mux2 i_5632(.S(n_6743), .A(code_data[2]), .B(axi_R[2]), .Z(n_5628
		));
	notech_nand2 i_124(.A(axi_io_WVALID), .B(axi_io_WREADY), .Z(n_222457061)
		);
	notech_reg_set code_data_reg_3(.CP(n_62414), .D(n_5634), .SD(1'b1), .Q(code_data
		[3]));
	notech_mux2 i_5640(.S(n_6743), .A(code_data[3]), .B(axi_R[3]), .Z(n_5634
		));
	notech_nao3 i_52(.A(n_222457061), .B(n_6747), .C(n_222257059), .Z(n_222557062
		));
	notech_reg_set code_data_reg_4(.CP(n_62414), .D(n_5640), .SD(1'b1), .Q(code_data
		[4]));
	notech_mux2 i_5648(.S(n_6743), .A(code_data[4]), .B(axi_R[4]), .Z(n_5640
		));
	notech_ao3 i_69(.A(n_222457061), .B(n_6740), .C(n_222357060), .Z(n_222657063
		));
	notech_reg_set code_data_reg_5(.CP(n_62414), .D(n_5646), .SD(1'b1), .Q(code_data
		[5]));
	notech_mux2 i_5656(.S(n_6743), .A(code_data[5]), .B(axi_R[5]), .Z(n_5646
		));
	notech_and2 i_80(.A(axi_io_RREADY), .B(axi_io_RVALID), .Z(n_222757064)
		);
	notech_reg_set code_data_reg_6(.CP(n_62392), .D(n_5652), .SD(1'b1), .Q(code_data
		[6]));
	notech_mux2 i_5664(.S(n_6743), .A(code_data[6]), .B(axi_R[6]), .Z(n_5652
		));
	notech_nao3 i_66(.A(n_6740), .B(n_6628), .C(n_222557062), .Z(n_222857065
		));
	notech_reg_set code_data_reg_7(.CP(n_62414), .D(n_5658), .SD(1'b1), .Q(code_data
		[7]));
	notech_mux2 i_5672(.S(n_6743), .A(code_data[7]), .B(axi_R[7]), .Z(n_5658
		));
	notech_nand2 i_19(.A(writeio_req), .B(n_6739), .Z(n_222957066));
	notech_reg_set code_data_reg_8(.CP(n_62394), .D(n_5664), .SD(1'b1), .Q(code_data
		[8]));
	notech_mux2 i_5680(.S(n_6743), .A(code_data[8]), .B(axi_R[8]), .Z(n_5664
		));
	notech_reg_set code_data_reg_9(.CP(n_62394), .D(n_5670), .SD(1'b1), .Q(code_data
		[9]));
	notech_mux2 i_5688(.S(n_6743), .A(code_data[9]), .B(axi_R[9]), .Z(n_5670
		));
	notech_nao3 i_1108(.A(readio_req), .B(n_222957066), .C(rf), .Z(n_223157068
		));
	notech_reg_set code_data_reg_10(.CP(n_62394), .D(n_5676), .SD(1'b1), .Q(code_data
		[10]));
	notech_mux2 i_5696(.S(n_6743), .A(code_data[10]), .B(axi_R[10]), .Z(n_5676
		));
	notech_reg_set code_data_reg_11(.CP(n_62394), .D(n_5682), .SD(1'b1), .Q(code_data
		[11]));
	notech_mux2 i_5704(.S(n_6743), .A(code_data[11]), .B(axi_R[11]), .Z(n_5682
		));
	notech_reg_set code_data_reg_12(.CP(n_62394), .D(n_5688), .SD(1'b1), .Q(code_data
		[12]));
	notech_mux2 i_5712(.S(n_6743), .A(code_data[12]), .B(axi_R[12]), .Z(n_5688
		));
	notech_reg_set code_data_reg_13(.CP(n_62394), .D(n_5694), .SD(1'b1), .Q(code_data
		[13]));
	notech_mux2 i_5720(.S(n_6743), .A(code_data[13]), .B(axi_R[13]), .Z(n_5694
		));
	notech_reg_set code_data_reg_14(.CP(n_62394), .D(n_5700), .SD(1'b1), .Q(code_data
		[14]));
	notech_mux2 i_5728(.S(n_6743), .A(code_data[14]), .B(axi_R[14]), .Z(n_5700
		));
	notech_and3 i_54(.A(n_2032), .B(n_1770), .C(n_6675), .Z(n_223657073));
	notech_reg_set code_data_reg_15(.CP(n_62394), .D(n_5706), .SD(1'b1), .Q(code_data
		[15]));
	notech_mux2 i_5736(.S(n_6743), .A(code_data[15]), .B(axi_R[15]), .Z(n_5706
		));
	notech_reg_set code_data_reg_16(.CP(n_62394), .D(n_5712), .SD(1'b1), .Q(code_data
		[16]));
	notech_mux2 i_5744(.S(n_57110), .A(code_data[16]), .B(axi_R[16]), .Z(n_5712
		));
	notech_nand3 i_38(.A(A4[1]), .B(n_1996), .C(n_59892), .Z(n_223857075));
	notech_reg_set code_data_reg_17(.CP(n_62394), .D(n_5718), .SD(1'b1), .Q(code_data
		[17]));
	notech_mux2 i_5752(.S(n_57110), .A(code_data[17]), .B(axi_R[17]), .Z(n_5718
		));
	notech_reg_set code_data_reg_18(.CP(n_62394), .D(n_5724), .SD(1'b1), .Q(code_data
		[18]));
	notech_mux2 i_5760(.S(n_57110), .A(code_data[18]), .B(axi_R[18]), .Z(n_5724
		));
	notech_nao3 i_39(.A(n_59892), .B(n_61972), .C(A4[1]), .Z(n_224057077));
	notech_reg_set code_data_reg_19(.CP(n_62394), .D(n_5730), .SD(1'b1), .Q(code_data
		[19]));
	notech_mux2 i_5768(.S(n_57110), .A(code_data[19]), .B(axi_R[19]), .Z(n_5730
		));
	notech_ao4 i_1166(.A(n_224057077), .B(n_6890), .C(n_223857075), .D(n_6922
		), .Z(n_224157078));
	notech_reg_set code_data_reg_20(.CP(n_62394), .D(n_5736), .SD(1'b1), .Q(code_data
		[20]));
	notech_mux2 i_5776(.S(n_57110), .A(code_data[20]), .B(axi_R[20]), .Z(n_5736
		));
	notech_reg_set code_data_reg_21(.CP(n_62394), .D(n_5742), .SD(1'b1), .Q(code_data
		[21]));
	notech_mux2 i_5784(.S(n_57110), .A(code_data[21]), .B(axi_R[21]), .Z(n_5742
		));
	notech_and3 i_37(.A(A4[1]), .B(n_61972), .C(n_6716), .Z(n_224357080));
	notech_reg_set code_data_reg_22(.CP(n_62394), .D(n_5748), .SD(1'b1), .Q(code_data
		[22]));
	notech_mux2 i_5792(.S(n_57110), .A(code_data[22]), .B(axi_R[22]), .Z(n_5748
		));
	notech_reg_set code_data_reg_23(.CP(n_62394), .D(n_5754), .SD(1'b1), .Q(code_data
		[23]));
	notech_mux2 i_5800(.S(n_57110), .A(code_data[23]), .B(axi_R[23]), .Z(n_5754
		));
	notech_nao3 i_36(.A(n_61972), .B(n_6716), .C(A4[1]), .Z(n_2245));
	notech_reg_set code_data_reg_24(.CP(n_62394), .D(n_5760), .SD(1'b1), .Q(code_data
		[24]));
	notech_mux2 i_5808(.S(n_57110), .A(code_data[24]), .B(axi_R[24]), .Z(n_5760
		));
	notech_ao4 i_1165(.A(n_61972), .B(n_6750), .C(n_2245), .D(n_6858), .Z(n_2246
		));
	notech_reg_set code_data_reg_25(.CP(n_62394), .D(n_5766), .SD(1'b1), .Q(code_data
		[25]));
	notech_mux2 i_5816(.S(n_57110), .A(code_data[25]), .B(axi_R[25]), .Z(n_5766
		));
	notech_reg_set code_data_reg_26(.CP(n_62394), .D(n_5772), .SD(1'b1), .Q(code_data
		[26]));
	notech_mux2 i_5824(.S(n_57110), .A(code_data[26]), .B(axi_R[26]), .Z(n_5772
		));
	notech_ao4 i_1175(.A(n_224057077), .B(n_6891), .C(n_223857075), .D(n_6923
		), .Z(n_2248));
	notech_reg_set code_data_reg_27(.CP(n_62368), .D(n_5778), .SD(1'b1), .Q(code_data
		[27]));
	notech_mux2 i_5832(.S(n_57110), .A(code_data[27]), .B(axi_R[27]), .Z(n_5778
		));
	notech_ao4 i_1174(.A(n_61972), .B(n_6751), .C(n_2245), .D(n_6859), .Z(n_2249
		));
	notech_reg_set code_data_reg_28(.CP(n_62368), .D(n_5784), .SD(1'b1), .Q(code_data
		[28]));
	notech_mux2 i_5840(.S(n_57110), .A(code_data[28]), .B(axi_R[28]), .Z(n_5784
		));
	notech_reg_set code_data_reg_29(.CP(n_62368), .D(n_5790), .SD(1'b1), .Q(code_data
		[29]));
	notech_mux2 i_5848(.S(n_57110), .A(code_data[29]), .B(axi_R[29]), .Z(n_5790
		));
	notech_ao4 i_1184(.A(n_224057077), .B(n_6892), .C(n_223857075), .D(n_6924
		), .Z(n_2251));
	notech_reg_set code_data_reg_30(.CP(n_62368), .D(n_5796), .SD(1'b1), .Q(code_data
		[30]));
	notech_mux2 i_5856(.S(n_57110), .A(code_data[30]), .B(axi_R[30]), .Z(n_5796
		));
	notech_ao4 i_1183(.A(n_1996), .B(n_6752), .C(n_2245), .D(n_6860), .Z(n_2252
		));
	notech_reg_set code_data_reg_31(.CP(n_62368), .D(n_5802), .SD(1'b1), .Q(code_data
		[31]));
	notech_mux2 i_5864(.S(n_57110), .A(code_data[31]), .B(axi_R[31]), .Z(n_5802
		));
	notech_reg_set code_data_reg_32(.CP(n_62368), .D(n_5808), .SD(1'b1), .Q(code_data
		[32]));
	notech_mux2 i_5872(.S(n_6744), .A(code_data[32]), .B(axi_R[0]), .Z(n_5808
		));
	notech_ao4 i_1193(.A(n_224057077), .B(n_6893), .C(n_223857075), .D(n_6925
		), .Z(n_2254));
	notech_reg_set code_data_reg_33(.CP(n_62352), .D(n_5814), .SD(1'b1), .Q(code_data
		[33]));
	notech_mux2 i_5880(.S(n_6744), .A(code_data[33]), .B(axi_R[1]), .Z(n_5814
		));
	notech_ao4 i_1192(.A(n_1996), .B(n_6753), .C(n_2245), .D(n_6861), .Z(n_2255
		));
	notech_reg_set code_data_reg_34(.CP(n_62368), .D(n_5820), .SD(1'b1), .Q(code_data
		[34]));
	notech_mux2 i_5888(.S(n_6744), .A(code_data[34]), .B(axi_R[2]), .Z(n_5820
		));
	notech_reg_set code_data_reg_35(.CP(n_62368), .D(n_5826), .SD(1'b1), .Q(code_data
		[35]));
	notech_mux2 i_5896(.S(n_6744), .A(code_data[35]), .B(axi_R[3]), .Z(n_5826
		));
	notech_ao4 i_1202(.A(n_224057077), .B(n_6894), .C(n_223857075), .D(n_6926
		), .Z(n_2257));
	notech_reg_set code_data_reg_36(.CP(n_62368), .D(n_5832), .SD(1'b1), .Q(code_data
		[36]));
	notech_mux2 i_5904(.S(n_6744), .A(code_data[36]), .B(axi_R[4]), .Z(n_5832
		));
	notech_ao4 i_1201(.A(n_1996), .B(n_6754), .C(n_2245), .D(n_6862), .Z(n_2258
		));
	notech_reg_set code_data_reg_37(.CP(n_62368), .D(n_5838), .SD(1'b1), .Q(code_data
		[37]));
	notech_mux2 i_5912(.S(n_6744), .A(code_data[37]), .B(axi_R[5]), .Z(n_5838
		));
	notech_reg_set code_data_reg_38(.CP(n_62368), .D(n_5844), .SD(1'b1), .Q(code_data
		[38]));
	notech_mux2 i_5920(.S(n_6744), .A(code_data[38]), .B(axi_R[6]), .Z(n_5844
		));
	notech_ao4 i_1211(.A(n_224057077), .B(n_6895), .C(n_223857075), .D(n_6927
		), .Z(n_2260));
	notech_reg_set code_data_reg_39(.CP(n_62368), .D(n_5850), .SD(1'b1), .Q(code_data
		[39]));
	notech_mux2 i_5928(.S(n_6744), .A(code_data[39]), .B(axi_R[7]), .Z(n_5850
		));
	notech_ao4 i_1210(.A(n_1996), .B(n_6755), .C(n_2245), .D(n_6863), .Z(n_2261
		));
	notech_reg_set code_data_reg_40(.CP(n_62368), .D(n_5856), .SD(1'b1), .Q(code_data
		[40]));
	notech_mux2 i_5936(.S(n_6744), .A(code_data[40]), .B(axi_R[8]), .Z(n_5856
		));
	notech_reg_set code_data_reg_41(.CP(n_62368), .D(n_5862), .SD(1'b1), .Q(code_data
		[41]));
	notech_mux2 i_5944(.S(n_6744), .A(code_data[41]), .B(axi_R[9]), .Z(n_5862
		));
	notech_ao4 i_1220(.A(n_224057077), .B(n_6896), .C(n_223857075), .D(n_6928
		), .Z(n_2263));
	notech_reg_set code_data_reg_42(.CP(n_62352), .D(n_5868), .SD(1'b1), .Q(code_data
		[42]));
	notech_mux2 i_5952(.S(n_6744), .A(code_data[42]), .B(axi_R[10]), .Z(n_5868
		));
	notech_ao4 i_1219(.A(n_1996), .B(n_6756), .C(n_2245), .D(n_6864), .Z(n_2264
		));
	notech_reg_set code_data_reg_43(.CP(n_62368), .D(n_5874), .SD(1'b1), .Q(code_data
		[43]));
	notech_mux2 i_5960(.S(n_6744), .A(code_data[43]), .B(axi_R[11]), .Z(n_5874
		));
	notech_reg_set code_data_reg_44(.CP(n_62374), .D(n_5880), .SD(1'b1), .Q(code_data
		[44]));
	notech_mux2 i_5968(.S(n_6744), .A(code_data[44]), .B(axi_R[12]), .Z(n_5880
		));
	notech_ao4 i_1229(.A(n_224057077), .B(n_6897), .C(n_223857075), .D(n_6929
		), .Z(n_2266));
	notech_reg_set code_data_reg_45(.CP(n_62354), .D(n_5886), .SD(1'b1), .Q(code_data
		[45]));
	notech_mux2 i_5976(.S(n_6744), .A(code_data[45]), .B(axi_R[13]), .Z(n_5886
		));
	notech_ao4 i_1228(.A(n_1996), .B(n_6757), .C(n_2245), .D(n_6865), .Z(n_2267
		));
	notech_reg_set code_data_reg_46(.CP(n_62354), .D(n_5892), .SD(1'b1), .Q(code_data
		[46]));
	notech_mux2 i_5984(.S(n_6744), .A(code_data[46]), .B(axi_R[14]), .Z(n_5892
		));
	notech_reg_set code_data_reg_47(.CP(n_62354), .D(n_5898), .SD(1'b1), .Q(code_data
		[47]));
	notech_mux2 i_5992(.S(n_6744), .A(code_data[47]), .B(axi_R[15]), .Z(n_5898
		));
	notech_ao4 i_1238(.A(n_224057077), .B(n_6898), .C(n_223857075), .D(n_6930
		), .Z(n_2269));
	notech_reg_set code_data_reg_48(.CP(n_62354), .D(n_5904), .SD(1'b1), .Q(code_data
		[48]));
	notech_mux2 i_6000(.S(n_54502), .A(code_data[48]), .B(axi_R[16]), .Z(n_5904
		));
	notech_ao4 i_1237(.A(n_1996), .B(n_6758), .C(n_2245), .D(n_6866), .Z(n_2270
		));
	notech_reg_set code_data_reg_49(.CP(n_62354), .D(n_5910), .SD(1'b1), .Q(code_data
		[49]));
	notech_mux2 i_6008(.S(n_54502), .A(code_data[49]), .B(axi_R[17]), .Z(n_5910
		));
	notech_reg_set code_data_reg_50(.CP(n_62354), .D(n_5916), .SD(1'b1), .Q(code_data
		[50]));
	notech_mux2 i_6016(.S(n_54502), .A(code_data[50]), .B(axi_R[18]), .Z(n_5916
		));
	notech_ao4 i_1247(.A(n_224057077), .B(n_6899), .C(n_223857075), .D(n_6931
		), .Z(n_2272));
	notech_reg_set code_data_reg_51(.CP(n_62354), .D(n_5922), .SD(1'b1), .Q(code_data
		[51]));
	notech_mux2 i_6024(.S(n_54502), .A(code_data[51]), .B(axi_R[19]), .Z(n_5922
		));
	notech_ao4 i_1246(.A(n_1996), .B(n_6759), .C(n_2245), .D(n_6867), .Z(n_2273
		));
	notech_reg_set code_data_reg_52(.CP(n_62354), .D(n_5928), .SD(1'b1), .Q(code_data
		[52]));
	notech_mux2 i_6032(.S(n_54502), .A(code_data[52]), .B(axi_R[20]), .Z(n_5928
		));
	notech_reg_set code_data_reg_53(.CP(n_62354), .D(n_5934), .SD(1'b1), .Q(code_data
		[53]));
	notech_mux2 i_6040(.S(n_54502), .A(code_data[53]), .B(axi_R[21]), .Z(n_5934
		));
	notech_ao4 i_1256(.A(n_224057077), .B(n_6900), .C(n_223857075), .D(n_6932
		), .Z(n_2275));
	notech_reg_set code_data_reg_54(.CP(n_62354), .D(n_5940), .SD(1'b1), .Q(code_data
		[54]));
	notech_mux2 i_6048(.S(n_54502), .A(code_data[54]), .B(axi_R[22]), .Z(n_5940
		));
	notech_ao4 i_1255(.A(n_1996), .B(n_6760), .C(n_2245), .D(n_6868), .Z(n_2276
		));
	notech_reg_set code_data_reg_55(.CP(n_62376), .D(n_5946), .SD(1'b1), .Q(code_data
		[55]));
	notech_mux2 i_6056(.S(n_54502), .A(code_data[55]), .B(axi_R[23]), .Z(n_5946
		));
	notech_reg_set code_data_reg_56(.CP(n_62376), .D(n_5952), .SD(1'b1), .Q(code_data
		[56]));
	notech_mux2 i_6064(.S(n_54502), .A(code_data[56]), .B(axi_R[24]), .Z(n_5952
		));
	notech_ao4 i_1265(.A(n_224057077), .B(n_6901), .C(n_223857075), .D(n_6933
		), .Z(n_2278));
	notech_reg_set code_data_reg_57(.CP(n_62376), .D(n_5958), .SD(1'b1), .Q(code_data
		[57]));
	notech_mux2 i_6072(.S(n_54502), .A(code_data[57]), .B(axi_R[25]), .Z(n_5958
		));
	notech_ao4 i_1264(.A(n_1996), .B(n_6761), .C(n_2245), .D(n_6869), .Z(n_2279
		));
	notech_reg_set code_data_reg_58(.CP(n_62376), .D(n_5964), .SD(1'b1), .Q(code_data
		[58]));
	notech_mux2 i_6080(.S(n_54502), .A(code_data[58]), .B(axi_R[26]), .Z(n_5964
		));
	notech_reg_set code_data_reg_59(.CP(n_62376), .D(n_5970), .SD(1'b1), .Q(code_data
		[59]));
	notech_mux2 i_6088(.S(n_54502), .A(code_data[59]), .B(axi_R[27]), .Z(n_5970
		));
	notech_ao4 i_1274(.A(n_224057077), .B(n_6902), .C(n_223857075), .D(n_6934
		), .Z(n_2281));
	notech_reg_set code_data_reg_60(.CP(n_62376), .D(n_5976), .SD(1'b1), .Q(code_data
		[60]));
	notech_mux2 i_6096(.S(n_54502), .A(code_data[60]), .B(axi_R[28]), .Z(n_5976
		));
	notech_ao4 i_1273(.A(n_1996), .B(n_6762), .C(n_2245), .D(n_6870), .Z(n_2282
		));
	notech_reg_set code_data_reg_61(.CP(n_62376), .D(n_5982), .SD(1'b1), .Q(code_data
		[61]));
	notech_mux2 i_6104(.S(n_54502), .A(code_data[61]), .B(axi_R[29]), .Z(n_5982
		));
	notech_reg_set code_data_reg_62(.CP(n_62376), .D(n_5988), .SD(1'b1), .Q(code_data
		[62]));
	notech_mux2 i_6112(.S(n_54502), .A(code_data[62]), .B(axi_R[30]), .Z(n_5988
		));
	notech_ao4 i_1283(.A(n_224057077), .B(n_6903), .C(n_223857075), .D(n_6935
		), .Z(n_2284));
	notech_reg_set code_data_reg_63(.CP(n_62376), .D(n_5994), .SD(1'b1), .Q(code_data
		[63]));
	notech_mux2 i_6120(.S(n_54502), .A(code_data[63]), .B(axi_R[31]), .Z(n_5994
		));
	notech_ao4 i_1282(.A(n_61972), .B(n_6763), .C(n_2245), .D(n_6871), .Z(n_2285
		));
	notech_reg_set code_data_reg_64(.CP(n_62376), .D(n_6000), .SD(1'b1), .Q(code_data
		[64]));
	notech_mux2 i_6128(.S(n_6745), .A(code_data[64]), .B(axi_R[0]), .Z(n_6000
		));
	notech_reg_set code_data_reg_65(.CP(n_62376), .D(n_6006), .SD(1'b1), .Q(code_data
		[65]));
	notech_mux2 i_6136(.S(n_6745), .A(code_data[65]), .B(axi_R[1]), .Z(n_6006
		));
	notech_ao4 i_1292(.A(n_224057077), .B(n_6904), .C(n_223857075), .D(n_6936
		), .Z(n_2287));
	notech_reg_set code_data_reg_66(.CP(n_62376), .D(n_6012), .SD(1'b1), .Q(code_data
		[66]));
	notech_mux2 i_6144(.S(n_6745), .A(code_data[66]), .B(axi_R[2]), .Z(n_6012
		));
	notech_ao4 i_1291(.A(n_61968), .B(n_6764), .C(n_2245), .D(n_6872), .Z(n_2288
		));
	notech_reg_set code_data_reg_67(.CP(n_62376), .D(n_6018), .SD(1'b1), .Q(code_data
		[67]));
	notech_mux2 i_6152(.S(n_6745), .A(code_data[67]), .B(axi_R[3]), .Z(n_6018
		));
	notech_reg_set code_data_reg_68(.CP(n_62376), .D(n_6024), .SD(1'b1), .Q(code_data
		[68]));
	notech_mux2 i_6160(.S(n_6745), .A(code_data[68]), .B(axi_R[4]), .Z(n_6024
		));
	notech_ao4 i_1301(.A(n_224057077), .B(n_6905), .C(n_223857075), .D(n_6937
		), .Z(n_2290));
	notech_reg_set code_data_reg_69(.CP(n_62376), .D(n_6030), .SD(1'b1), .Q(code_data
		[69]));
	notech_mux2 i_6168(.S(n_6745), .A(code_data[69]), .B(axi_R[5]), .Z(n_6030
		));
	notech_ao4 i_1300(.A(n_61968), .B(n_6765), .C(n_2245), .D(n_6873), .Z(n_2291
		));
	notech_reg_set code_data_reg_70(.CP(n_62376), .D(n_6036), .SD(1'b1), .Q(code_data
		[70]));
	notech_mux2 i_6176(.S(n_6745), .A(code_data[70]), .B(axi_R[6]), .Z(n_6036
		));
	notech_reg_set code_data_reg_71(.CP(n_62376), .D(n_6042), .SD(1'b1), .Q(code_data
		[71]));
	notech_mux2 i_6184(.S(n_6745), .A(code_data[71]), .B(axi_R[7]), .Z(n_6042
		));
	notech_ao4 i_1310(.A(n_54358), .B(n_6906), .C(n_54349), .D(n_6938), .Z(n_2293
		));
	notech_reg_set code_data_reg_72(.CP(n_62376), .D(n_6048), .SD(1'b1), .Q(code_data
		[72]));
	notech_mux2 i_6192(.S(n_6745), .A(code_data[72]), .B(axi_R[8]), .Z(n_6048
		));
	notech_ao4 i_1309(.A(n_61968), .B(n_6766), .C(n_54369), .D(n_6874), .Z(n_2294
		));
	notech_reg_set code_data_reg_73(.CP(n_62376), .D(n_6054), .SD(1'b1), .Q(code_data
		[73]));
	notech_mux2 i_6200(.S(n_6745), .A(code_data[73]), .B(axi_R[9]), .Z(n_6054
		));
	notech_reg_set code_data_reg_74(.CP(n_62398), .D(n_6060), .SD(1'b1), .Q(code_data
		[74]));
	notech_mux2 i_6208(.S(n_6745), .A(code_data[74]), .B(axi_R[10]), .Z(n_6060
		));
	notech_ao4 i_1319(.A(n_54358), .B(n_6907), .C(n_54349), .D(n_6939), .Z(n_2296
		));
	notech_reg_set code_data_reg_75(.CP(n_62374), .D(n_6066), .SD(1'b1), .Q(code_data
		[75]));
	notech_mux2 i_6216(.S(n_6745), .A(code_data[75]), .B(axi_R[11]), .Z(n_6066
		));
	notech_ao4 i_1318(.A(n_61972), .B(n_6767), .C(n_54369), .D(n_6875), .Z(n_2297
		));
	notech_reg_set code_data_reg_76(.CP(n_62398), .D(n_6072), .SD(1'b1), .Q(code_data
		[76]));
	notech_mux2 i_6224(.S(n_6745), .A(code_data[76]), .B(axi_R[12]), .Z(n_6072
		));
	notech_reg_set code_data_reg_77(.CP(n_62398), .D(n_6078), .SD(1'b1), .Q(code_data
		[77]));
	notech_mux2 i_6232(.S(n_6745), .A(code_data[77]), .B(axi_R[13]), .Z(n_6078
		));
	notech_ao4 i_1328(.A(n_54358), .B(n_6908), .C(n_54349), .D(n_6940), .Z(n_2299
		));
	notech_reg_set code_data_reg_78(.CP(n_62398), .D(n_6084), .SD(1'b1), .Q(code_data
		[78]));
	notech_mux2 i_6240(.S(n_6745), .A(code_data[78]), .B(axi_R[14]), .Z(n_6084
		));
	notech_ao4 i_1327(.A(n_61972), .B(n_6768), .C(n_54369), .D(n_6876), .Z(n_2300
		));
	notech_reg_set code_data_reg_79(.CP(n_62398), .D(n_6090), .SD(1'b1), .Q(code_data
		[79]));
	notech_mux2 i_6248(.S(n_6745), .A(code_data[79]), .B(axi_R[15]), .Z(n_6090
		));
	notech_reg_set code_data_reg_80(.CP(n_62398), .D(n_6096), .SD(1'b1), .Q(code_data
		[80]));
	notech_mux2 i_6256(.S(n_54513), .A(code_data[80]), .B(axi_R[16]), .Z(n_6096
		));
	notech_ao4 i_1337(.A(n_54358), .B(n_6909), .C(n_54349), .D(n_6941), .Z(n_2302
		));
	notech_reg_set code_data_reg_81(.CP(n_62398), .D(n_6102), .SD(1'b1), .Q(code_data
		[81]));
	notech_mux2 i_6264(.S(n_54513), .A(code_data[81]), .B(axi_R[17]), .Z(n_6102
		));
	notech_ao4 i_1336(.A(n_61968), .B(n_6769), .C(n_54369), .D(n_6877), .Z(n_2303
		));
	notech_reg_set code_data_reg_82(.CP(n_62398), .D(n_6108), .SD(1'b1), .Q(code_data
		[82]));
	notech_mux2 i_6272(.S(n_54513), .A(code_data[82]), .B(axi_R[18]), .Z(n_6108
		));
	notech_reg_set code_data_reg_83(.CP(n_62398), .D(n_6114), .SD(1'b1), .Q(code_data
		[83]));
	notech_mux2 i_6280(.S(n_54513), .A(code_data[83]), .B(axi_R[19]), .Z(n_6114
		));
	notech_ao4 i_1346(.A(n_54358), .B(n_6910), .C(n_54349), .D(n_6942), .Z(n_2305
		));
	notech_reg_set code_data_reg_84(.CP(n_62398), .D(n_6120), .SD(1'b1), .Q(code_data
		[84]));
	notech_mux2 i_6288(.S(n_54513), .A(code_data[84]), .B(axi_R[20]), .Z(n_6120
		));
	notech_ao4 i_1345(.A(n_61968), .B(n_6770), .C(n_54369), .D(n_6878), .Z(n_2306
		));
	notech_reg_set code_data_reg_85(.CP(n_62398), .D(n_6126), .SD(1'b1), .Q(code_data
		[85]));
	notech_mux2 i_6296(.S(n_54513), .A(code_data[85]), .B(axi_R[21]), .Z(n_6126
		));
	notech_reg_set code_data_reg_86(.CP(n_62398), .D(n_6132), .SD(1'b1), .Q(code_data
		[86]));
	notech_mux2 i_6304(.S(n_54513), .A(code_data[86]), .B(axi_R[22]), .Z(n_6132
		));
	notech_ao4 i_1355(.A(n_54358), .B(n_6911), .C(n_54349), .D(n_6943), .Z(n_2308
		));
	notech_reg_set code_data_reg_87(.CP(n_62398), .D(n_6138), .SD(1'b1), .Q(code_data
		[87]));
	notech_mux2 i_6312(.S(n_54513), .A(code_data[87]), .B(axi_R[23]), .Z(n_6138
		));
	notech_ao4 i_1354(.A(n_61968), .B(n_6771), .C(n_54369), .D(n_6879), .Z(n_2309
		));
	notech_reg_set code_data_reg_88(.CP(n_62398), .D(n_6144), .SD(1'b1), .Q(code_data
		[88]));
	notech_mux2 i_6320(.S(n_54513), .A(code_data[88]), .B(axi_R[24]), .Z(n_6144
		));
	notech_reg_set code_data_reg_89(.CP(n_62398), .D(n_6150), .SD(1'b1), .Q(code_data
		[89]));
	notech_mux2 i_6328(.S(n_54513), .A(code_data[89]), .B(axi_R[25]), .Z(n_6150
		));
	notech_ao4 i_1364(.A(n_54358), .B(n_6912), .C(n_54349), .D(n_6944), .Z(n_2311
		));
	notech_reg_set code_data_reg_90(.CP(n_62398), .D(n_6156), .SD(1'b1), .Q(code_data
		[90]));
	notech_mux2 i_6336(.S(n_54513), .A(code_data[90]), .B(axi_R[26]), .Z(n_6156
		));
	notech_ao4 i_1363(.A(n_61968), .B(n_6772), .C(n_54369), .D(n_6880), .Z(n_2312
		));
	notech_reg_set code_data_reg_91(.CP(n_62398), .D(n_6162), .SD(1'b1), .Q(code_data
		[91]));
	notech_mux2 i_6344(.S(n_54513), .A(code_data[91]), .B(axi_R[27]), .Z(n_6162
		));
	notech_reg_set code_data_reg_92(.CP(n_62398), .D(n_6168), .SD(1'b1), .Q(code_data
		[92]));
	notech_mux2 i_6352(.S(n_54513), .A(code_data[92]), .B(axi_R[28]), .Z(n_6168
		));
	notech_ao4 i_1373(.A(n_54358), .B(n_6913), .C(n_54349), .D(n_6945), .Z(n_2314
		));
	notech_reg_set code_data_reg_93(.CP(n_62398), .D(n_6174), .SD(1'b1), .Q(code_data
		[93]));
	notech_mux2 i_6360(.S(n_54513), .A(code_data[93]), .B(axi_R[29]), .Z(n_6174
		));
	notech_ao4 i_1372(.A(n_61968), .B(n_6773), .C(n_54369), .D(n_6881), .Z(n_2315
		));
	notech_reg_set code_data_reg_94(.CP(n_62374), .D(n_6180), .SD(1'b1), .Q(code_data
		[94]));
	notech_mux2 i_6368(.S(n_54513), .A(code_data[94]), .B(axi_R[30]), .Z(n_6180
		));
	notech_reg_set code_data_reg_95(.CP(n_62374), .D(n_6186), .SD(1'b1), .Q(code_data
		[95]));
	notech_mux2 i_6376(.S(n_54513), .A(code_data[95]), .B(axi_R[31]), .Z(n_6186
		));
	notech_ao4 i_1382(.A(n_54358), .B(n_6914), .C(n_54349), .D(n_6946), .Z(n_2317
		));
	notech_reg_set code_data_reg_96(.CP(n_62374), .D(n_6192), .SD(1'b1), .Q(code_data
		[96]));
	notech_mux2 i_6384(.S(n_6746), .A(code_data[96]), .B(axi_R[0]), .Z(n_6192
		));
	notech_ao4 i_1381(.A(n_61972), .B(n_6774), .C(n_54369), .D(n_6882), .Z(n_2318
		));
	notech_reg_set code_data_reg_97(.CP(n_62374), .D(n_6198), .SD(1'b1), .Q(code_data
		[97]));
	notech_mux2 i_6392(.S(n_6746), .A(code_data[97]), .B(axi_R[1]), .Z(n_6198
		));
	notech_reg_set code_data_reg_98(.CP(n_62374), .D(n_6204), .SD(1'b1), .Q(code_data
		[98]));
	notech_mux2 i_6400(.S(n_6746), .A(code_data[98]), .B(axi_R[2]), .Z(n_6204
		));
	notech_ao4 i_1391(.A(n_54358), .B(n_6915), .C(n_54349), .D(n_6947), .Z(n_2320
		));
	notech_reg_set code_data_reg_99(.CP(n_62374), .D(n_6210), .SD(1'b1), .Q(code_data
		[99]));
	notech_mux2 i_6408(.S(n_6746), .A(code_data[99]), .B(axi_R[3]), .Z(n_6210
		));
	notech_ao4 i_1390(.A(n_61972), .B(n_6775), .C(n_54369), .D(n_6883), .Z(n_2321
		));
	notech_reg_set code_data_reg_100(.CP(n_62374), .D(n_6216), .SD(1'b1), .Q
		(code_data[100]));
	notech_mux2 i_6416(.S(n_6746), .A(code_data[100]), .B(axi_R[4]), .Z(n_6216
		));
	notech_reg_set code_data_reg_101(.CP(n_62374), .D(n_6222), .SD(1'b1), .Q
		(code_data[101]));
	notech_mux2 i_6424(.S(n_6746), .A(code_data[101]), .B(axi_R[5]), .Z(n_6222
		));
	notech_ao4 i_1400(.A(n_54358), .B(n_6916), .C(n_223857075), .D(n_6948), 
		.Z(n_2323));
	notech_reg_set code_data_reg_102(.CP(n_62374), .D(n_6228), .SD(1'b1), .Q
		(code_data[102]));
	notech_mux2 i_6432(.S(n_6746), .A(code_data[102]), .B(axi_R[6]), .Z(n_6228
		));
	notech_ao4 i_1399(.A(n_61972), .B(n_6776), .C(n_2245), .D(n_6884), .Z(n_2324
		));
	notech_reg_set code_data_reg_103(.CP(n_62374), .D(n_6234), .SD(1'b1), .Q
		(code_data[103]));
	notech_mux2 i_6440(.S(n_6746), .A(code_data[103]), .B(axi_R[7]), .Z(n_6234
		));
	notech_reg_set code_data_reg_104(.CP(n_62354), .D(n_6240), .SD(1'b1), .Q
		(code_data[104]));
	notech_mux2 i_6448(.S(n_6746), .A(code_data[104]), .B(axi_R[8]), .Z(n_6240
		));
	notech_ao4 i_1409(.A(n_54358), .B(n_6917), .C(n_54349), .D(n_6949), .Z(n_2326
		));
	notech_reg_set code_data_reg_105(.CP(n_62354), .D(n_6246), .SD(1'b1), .Q
		(code_data[105]));
	notech_mux2 i_6456(.S(n_6746), .A(code_data[105]), .B(axi_R[9]), .Z(n_6246
		));
	notech_ao4 i_1408(.A(n_61972), .B(n_6777), .C(n_54369), .D(n_6885), .Z(n_2327
		));
	notech_reg_set code_data_reg_106(.CP(n_62378), .D(n_6252), .SD(1'b1), .Q
		(code_data[106]));
	notech_mux2 i_6464(.S(n_6746), .A(code_data[106]), .B(axi_R[10]), .Z(n_6252
		));
	notech_reg_set code_data_reg_107(.CP(n_62356), .D(n_6258), .SD(1'b1), .Q
		(code_data[107]));
	notech_mux2 i_6472(.S(n_6746), .A(code_data[107]), .B(axi_R[11]), .Z(n_6258
		));
	notech_ao4 i_1418(.A(n_54358), .B(n_6918), .C(n_54349), .D(n_6950), .Z(n_2329
		));
	notech_reg_set code_data_reg_108(.CP(n_62356), .D(n_6264), .SD(1'b1), .Q
		(code_data[108]));
	notech_mux2 i_6480(.S(n_6746), .A(code_data[108]), .B(axi_R[12]), .Z(n_6264
		));
	notech_ao4 i_1417(.A(n_61972), .B(n_6778), .C(n_54369), .D(n_6886), .Z(n_2330
		));
	notech_reg_set code_data_reg_109(.CP(n_62356), .D(n_6270), .SD(1'b1), .Q
		(code_data[109]));
	notech_mux2 i_6488(.S(n_6746), .A(code_data[109]), .B(axi_R[13]), .Z(n_6270
		));
	notech_reg_set code_data_reg_110(.CP(n_62356), .D(n_6276), .SD(1'b1), .Q
		(code_data[110]));
	notech_mux2 i_6496(.S(n_6746), .A(code_data[110]), .B(axi_R[14]), .Z(n_6276
		));
	notech_ao4 i_1427(.A(n_54358), .B(n_6919), .C(n_54349), .D(n_6951), .Z(n_2332
		));
	notech_reg_set code_data_reg_111(.CP(n_62356), .D(n_6282), .SD(1'b1), .Q
		(code_data[111]));
	notech_mux2 i_6504(.S(n_6746), .A(code_data[111]), .B(axi_R[15]), .Z(n_6282
		));
	notech_ao4 i_1426(.A(n_61972), .B(n_6779), .C(n_54369), .D(n_6887), .Z(n_2333
		));
	notech_reg_set code_data_reg_112(.CP(n_62356), .D(n_6288), .SD(1'b1), .Q
		(code_data[112]));
	notech_mux2 i_6512(.S(n_54524), .A(code_data[112]), .B(axi_R[16]), .Z(n_6288
		));
	notech_reg_set code_data_reg_113(.CP(n_62356), .D(n_6294), .SD(1'b1), .Q
		(code_data[113]));
	notech_mux2 i_6520(.S(n_54524), .A(code_data[113]), .B(axi_R[17]), .Z(n_6294
		));
	notech_ao4 i_1436(.A(n_54358), .B(n_6920), .C(n_54349), .D(n_6952), .Z(n_2335
		));
	notech_reg_set code_data_reg_114(.CP(n_62356), .D(n_6300), .SD(1'b1), .Q
		(code_data[114]));
	notech_mux2 i_6528(.S(n_54524), .A(code_data[114]), .B(axi_R[18]), .Z(n_6300
		));
	notech_ao4 i_1435(.A(n_61972), .B(n_6780), .C(n_54369), .D(n_6888), .Z(n_2336
		));
	notech_reg_set code_data_reg_115(.CP(n_62356), .D(n_6306), .SD(1'b1), .Q
		(code_data[115]));
	notech_mux2 i_6536(.S(n_54524), .A(code_data[115]), .B(axi_R[19]), .Z(n_6306
		));
	notech_reg_set code_data_reg_116(.CP(n_62356), .D(n_6312), .SD(1'b1), .Q
		(code_data[116]));
	notech_mux2 i_6544(.S(n_54524), .A(code_data[116]), .B(axi_R[20]), .Z(n_6312
		));
	notech_ao4 i_1445(.A(n_54358), .B(n_6921), .C(n_54349), .D(n_6953), .Z(n_2338
		));
	notech_reg_set code_data_reg_117(.CP(n_62378), .D(n_6318), .SD(1'b1), .Q
		(code_data[117]));
	notech_mux2 i_6552(.S(n_54524), .A(code_data[117]), .B(axi_R[21]), .Z(n_6318
		));
	notech_ao4 i_1444(.A(n_61972), .B(n_6781), .C(n_54369), .D(n_6889), .Z(n_2339
		));
	notech_reg_set code_data_reg_118(.CP(n_62378), .D(n_6324), .SD(1'b1), .Q
		(code_data[118]));
	notech_mux2 i_6560(.S(n_54524), .A(code_data[118]), .B(axi_R[22]), .Z(n_6324
		));
	notech_reg_set code_data_reg_119(.CP(n_62378), .D(n_6330), .SD(1'b1), .Q
		(code_data[119]));
	notech_mux2 i_6568(.S(n_54524), .A(code_data[119]), .B(axi_R[23]), .Z(n_6330
		));
	notech_and2 i_1096(.A(n_61808), .B(n_962), .Z(\nbus_11697[0] ));
	notech_reg_set code_data_reg_120(.CP(n_62378), .D(n_6336), .SD(1'b1), .Q
		(code_data[120]));
	notech_mux2 i_6576(.S(n_54524), .A(code_data[120]), .B(axi_R[24]), .Z(n_6336
		));
	notech_nor2 i_904(.A(n_222957066), .B(n_222857065), .Z(\nbus_11686[0] )
		);
	notech_reg_set code_data_reg_121(.CP(n_62378), .D(n_6342), .SD(1'b1), .Q
		(code_data[121]));
	notech_mux2 i_6584(.S(n_54524), .A(code_data[121]), .B(axi_R[25]), .Z(n_6342
		));
	notech_nor2 i_901(.A(n_223157068), .B(n_222857065), .Z(\nbus_11699[0] )
		);
	notech_reg_set code_data_reg_122(.CP(n_62378), .D(n_6348), .SD(1'b1), .Q
		(code_data[122]));
	notech_mux2 i_6592(.S(n_54524), .A(code_data[122]), .B(axi_R[26]), .Z(n_6348
		));
	notech_and4 i_900(.A(axi_io_RREADY), .B(axi_io_RVALID), .C(n_222657063),
		 .D(n_61809), .Z(\nbus_11696[0] ));
	notech_reg_set code_data_reg_123(.CP(n_62378), .D(n_6354), .SD(1'b1), .Q
		(code_data[123]));
	notech_mux2 i_6600(.S(n_54524), .A(code_data[123]), .B(axi_R[27]), .Z(n_6354
		));
	notech_or4 i_899(.A(n_2030), .B(n_2109), .C(n_1998), .D(n_2014), .Z(\nbus_11692[96] 
		));
	notech_reg_set code_data_reg_124(.CP(n_62378), .D(n_6360), .SD(1'b1), .Q
		(code_data[124]));
	notech_mux2 i_6608(.S(n_54524), .A(code_data[124]), .B(axi_R[28]), .Z(n_6360
		));
	notech_or4 i_898(.A(n_1998), .B(n_2014), .C(n_2030), .D(n_214256979), .Z
		(\nbus_11692[64] ));
	notech_reg_set code_data_reg_125(.CP(n_62378), .D(n_6366), .SD(1'b1), .Q
		(code_data[125]));
	notech_mux2 i_6616(.S(n_54524), .A(code_data[125]), .B(axi_R[29]), .Z(n_6366
		));
	notech_or4 i_897(.A(n_1998), .B(n_2014), .C(n_2030), .D(n_217757014), .Z
		(\nbus_11692[32] ));
	notech_reg_set code_data_reg_126(.CP(n_62378), .D(n_6372), .SD(1'b1), .Q
		(code_data[126]));
	notech_mux2 i_6624(.S(n_54524), .A(code_data[126]), .B(axi_R[30]), .Z(n_6372
		));
	notech_or4 i_896(.A(n_1998), .B(n_2014), .C(n_2030), .D(n_2038), .Z(\nbus_11692[0] 
		));
	notech_reg_set code_data_reg_127(.CP(n_62378), .D(n_6378), .SD(1'b1), .Q
		(code_data[127]));
	notech_mux2 i_6632(.S(n_54524), .A(code_data[127]), .B(axi_R[31]), .Z(n_6378
		));
	notech_or4 i_57456(.A(write_ack), .B(n_2001), .C(busy), .D(n_6982), .Z(n_28023
		));
	notech_reg axi_io_WLAST_reg(.CP(n_62378), .D(n_6384), .CD(n_61808), .Q(axi_io_WLAST
		));
	notech_mux2 i_6640(.S(n_1760), .A(n_27181), .B(axi_io_WLAST), .Z(n_6384)
		);
	notech_and2 i_29(.A(axi_io_ARVALID), .B(axi_io_ARREADY), .Z(n_28035));
	notech_reg_set axi_ARBURST_reg_0(.CP(n_62378), .D(n_6395), .SD(n_61808),
		 .Q(axi_ARBURST[0]));
	notech_and2 i_26(.A(axi_io_AWVALID), .B(axi_io_AWREADY), .Z(n_27181));
	notech_nao3 i_6653(.A(n_61959), .B(1'b1), .C(axi_ARBURST[0]), .Z(n_6395)
		);
	notech_reg axi_ARBURST_reg_1(.CP(n_62378), .D(n_6399), .CD(n_61808), .Q(axi_ARBURST
		[1]));
	notech_ao3 i_6658(.A(n_61972), .B(axi_ARBURST[1]), .C(n_1742), .Z(n_6399
		));
	notech_and2 i_916(.A(write_msk[1]), .B(n_6733), .Z(n_28066));
	notech_reg axi_AWSIZE_reg_0(.CP(n_62378), .D(n_6405), .CD(n_61808), .Q(axi_AWSIZE
		[0]));
	notech_ao3 i_6666(.A(n_61972), .B(axi_AWSIZE[0]), .C(n_1742), .Z(n_6405)
		);
	notech_and2 i_917(.A(write_msk[2]), .B(n_6733), .Z(n_28072));
	notech_reg_set axi_AWSIZE_reg_1(.CP(n_62378), .D(n_6413), .SD(n_61808), 
		.Q(axi_AWSIZE[1]));
	notech_and2 i_918(.A(write_msk[3]), .B(n_6733), .Z(n_28078));
	notech_nao3 i_6677(.A(n_61959), .B(1'b1), .C(axi_AWSIZE[1]), .Z(n_6413)
		);
	notech_reg axi_AWSIZE_reg_2(.CP(n_62378), .D(n_6417), .CD(n_61808), .Q(axi_AWSIZE
		[2]));
	notech_ao3 i_6682(.A(n_61972), .B(axi_AWSIZE[2]), .C(n_1742), .Z(n_6417)
		);
	notech_ao3 i_1048(.A(cacheQ[146]), .B(n_6977), .C(n_2032), .Z(n_27983)
		);
	notech_reg axi_WVALID_reg(.CP(n_62378), .D(n_6420), .CD(n_61808), .Q(axi_WVALID
		));
	notech_mux2 i_6688(.S(n_1221), .A(n_1767), .B(axi_WVALID), .Z(n_6420));
	notech_ao3 i_1049(.A(cacheQ[147]), .B(n_6977), .C(n_2032), .Z(n_27988)
		);
	notech_reg axi_io_W_reg_0(.CP(n_62356), .D(n_6426), .CD(n_61808), .Q(axi_io_W
		[0]));
	notech_mux2 i_6696(.S(\nbus_11686[0] ), .A(axi_io_W[0]), .B(writeio_data
		[0]), .Z(n_6426));
	notech_ao3 i_1050(.A(cacheQ[149]), .B(n_6977), .C(n_2032), .Z(n_27998)
		);
	notech_reg axi_io_W_reg_1(.CP(n_62356), .D(n_6432), .CD(n_61804), .Q(axi_io_W
		[1]));
	notech_mux2 i_6704(.S(\nbus_11686[0] ), .A(axi_io_W[1]), .B(writeio_data
		[1]), .Z(n_6432));
	notech_ao3 i_57501(.A(fsm[0]), .B(fsm[4]), .C(n_1998), .Z(n_27143));
	notech_reg axi_io_W_reg_2(.CP(n_62358), .D(n_6438), .CD(n_61804), .Q(axi_io_W
		[2]));
	notech_mux2 i_6712(.S(\nbus_11686[0] ), .A(axi_io_W[2]), .B(writeio_data
		[2]), .Z(n_6438));
	notech_and2 i_1072(.A(write_data[8]), .B(n_6629), .Z(n_29532));
	notech_reg axi_io_W_reg_3(.CP(n_62358), .D(n_6444), .CD(n_61804), .Q(axi_io_W
		[3]));
	notech_mux2 i_6720(.S(\nbus_11686[0] ), .A(axi_io_W[3]), .B(writeio_data
		[3]), .Z(n_6444));
	notech_and2 i_1073(.A(write_data[9]), .B(n_6629), .Z(n_29538));
	notech_reg axi_io_W_reg_4(.CP(n_62358), .D(n_6450), .CD(n_61804), .Q(axi_io_W
		[4]));
	notech_mux2 i_6728(.S(\nbus_11686[0] ), .A(axi_io_W[4]), .B(writeio_data
		[4]), .Z(n_6450));
	notech_and2 i_1074(.A(write_data[10]), .B(n_6629), .Z(n_29544));
	notech_reg axi_io_W_reg_5(.CP(n_62358), .D(n_6456), .CD(n_61804), .Q(axi_io_W
		[5]));
	notech_mux2 i_6736(.S(\nbus_11686[0] ), .A(axi_io_W[5]), .B(writeio_data
		[5]), .Z(n_6456));
	notech_and2 i_1075(.A(write_data[11]), .B(n_6629), .Z(n_29550));
	notech_reg axi_io_W_reg_6(.CP(n_62358), .D(n_6462), .CD(n_61804), .Q(axi_io_W
		[6]));
	notech_mux2 i_6744(.S(\nbus_11686[0] ), .A(axi_io_W[6]), .B(writeio_data
		[6]), .Z(n_6462));
	notech_and2 i_1076(.A(write_data[12]), .B(n_6629), .Z(n_29556));
	notech_reg axi_io_W_reg_7(.CP(n_62358), .D(n_6468), .CD(n_61804), .Q(axi_io_W
		[7]));
	notech_mux2 i_6752(.S(\nbus_11686[0] ), .A(axi_io_W[7]), .B(writeio_data
		[7]), .Z(n_6468));
	notech_and2 i_1077(.A(write_data[13]), .B(n_6629), .Z(n_29562));
	notech_reg axi_io_W_reg_8(.CP(n_62358), .D(n_6474), .CD(n_61804), .Q(axi_io_W
		[8]));
	notech_mux2 i_6760(.S(n_61206), .A(axi_io_W[8]), .B(writeio_data[8]), .Z
		(n_6474));
	notech_and2 i_1078(.A(write_data[14]), .B(n_6629), .Z(n_29568));
	notech_reg axi_io_W_reg_9(.CP(n_62358), .D(n_6480), .CD(n_61803), .Q(axi_io_W
		[9]));
	notech_mux2 i_6768(.S(n_61202), .A(axi_io_W[9]), .B(writeio_data[9]), .Z
		(n_6480));
	notech_and2 i_1079(.A(write_data[15]), .B(n_6629), .Z(n_29574));
	notech_reg axi_io_W_reg_10(.CP(n_62358), .D(n_6486), .CD(n_61803), .Q(axi_io_W
		[10]));
	notech_mux2 i_6776(.S(n_61202), .A(axi_io_W[10]), .B(writeio_data[10]), 
		.Z(n_6486));
	notech_and2 i_1080(.A(write_data[16]), .B(n_6629), .Z(n_29580));
	notech_reg axi_io_W_reg_11(.CP(n_62358), .D(n_6492), .CD(n_61803), .Q(axi_io_W
		[11]));
	notech_mux2 i_6784(.S(n_61202), .A(axi_io_W[11]), .B(writeio_data[11]), 
		.Z(n_6492));
	notech_and2 i_1081(.A(write_data[17]), .B(n_6629), .Z(n_29586));
	notech_reg axi_io_W_reg_12(.CP(n_62358), .D(n_6498), .CD(n_61803), .Q(axi_io_W
		[12]));
	notech_mux2 i_6792(.S(n_61202), .A(axi_io_W[12]), .B(writeio_data[12]), 
		.Z(n_6498));
	notech_and2 i_1082(.A(write_data[18]), .B(n_6629), .Z(n_29592));
	notech_reg axi_io_W_reg_13(.CP(n_62358), .D(n_6504), .CD(n_61804), .Q(axi_io_W
		[13]));
	notech_mux2 i_6800(.S(n_61202), .A(axi_io_W[13]), .B(writeio_data[13]), 
		.Z(n_6504));
	notech_and2 i_1083(.A(write_data[19]), .B(n_6629), .Z(n_29598));
	notech_reg axi_io_W_reg_14(.CP(n_62358), .D(n_6510), .CD(n_61804), .Q(axi_io_W
		[14]));
	notech_mux2 i_6808(.S(n_61202), .A(axi_io_W[14]), .B(writeio_data[14]), 
		.Z(n_6510));
	notech_and2 i_1084(.A(write_data[20]), .B(n_61215), .Z(n_29604));
	notech_reg axi_io_W_reg_15(.CP(n_62358), .D(n_6516), .CD(n_61803), .Q(axi_io_W
		[15]));
	notech_mux2 i_6816(.S(n_61202), .A(axi_io_W[15]), .B(writeio_data[15]), 
		.Z(n_6516));
	notech_and2 i_1085(.A(write_data[21]), .B(n_61215), .Z(n_29610));
	notech_reg axi_io_W_reg_16(.CP(n_62358), .D(n_6522), .CD(n_61804), .Q(axi_io_W
		[16]));
	notech_mux2 i_6824(.S(n_61202), .A(axi_io_W[16]), .B(writeio_data[16]), 
		.Z(n_6522));
	notech_and2 i_1086(.A(write_data[22]), .B(n_61215), .Z(n_29616));
	notech_reg axi_io_W_reg_17(.CP(n_62358), .D(n_6528), .CD(n_61804), .Q(axi_io_W
		[17]));
	notech_mux2 i_6832(.S(n_61202), .A(axi_io_W[17]), .B(writeio_data[17]), 
		.Z(n_6528));
	notech_and2 i_1087(.A(write_data[23]), .B(n_61215), .Z(n_29622));
	notech_reg axi_io_W_reg_18(.CP(n_62358), .D(n_6534), .CD(n_61806), .Q(axi_io_W
		[18]));
	notech_mux2 i_6840(.S(n_61202), .A(axi_io_W[18]), .B(writeio_data[18]), 
		.Z(n_6534));
	notech_and2 i_1088(.A(write_data[24]), .B(n_61215), .Z(n_29628));
	notech_reg axi_io_W_reg_19(.CP(n_62358), .D(n_6540), .CD(n_61806), .Q(axi_io_W
		[19]));
	notech_mux2 i_6848(.S(n_61202), .A(axi_io_W[19]), .B(writeio_data[19]), 
		.Z(n_6540));
	notech_and2 i_1089(.A(write_data[25]), .B(n_61215), .Z(n_29634));
	notech_reg axi_io_W_reg_20(.CP(n_62358), .D(n_6546), .CD(n_61806), .Q(axi_io_W
		[20]));
	notech_mux2 i_6856(.S(n_61202), .A(axi_io_W[20]), .B(writeio_data[20]), 
		.Z(n_6546));
	notech_and2 i_1090(.A(write_data[26]), .B(n_61215), .Z(n_29640));
	notech_reg axi_io_W_reg_21(.CP(clk), .D(n_6552), .CD(n_61806), .Q(axi_io_W
		[21]));
	notech_mux2 i_6864(.S(n_61206), .A(axi_io_W[21]), .B(writeio_data[21]), 
		.Z(n_6552));
	notech_and2 i_1091(.A(write_data[27]), .B(n_61215), .Z(n_29646));
	notech_reg axi_io_W_reg_22(.CP(clk), .D(n_6558), .CD(n_61806), .Q(axi_io_W
		[22]));
	notech_mux2 i_6872(.S(n_61206), .A(axi_io_W[22]), .B(writeio_data[22]), 
		.Z(n_6558));
	notech_and2 i_1092(.A(write_data[28]), .B(n_61215), .Z(n_29652));
	notech_reg axi_io_W_reg_23(.CP(clk), .D(n_6564), .CD(n_61806), .Q(axi_io_W
		[23]));
	notech_mux2 i_6880(.S(n_61206), .A(axi_io_W[23]), .B(writeio_data[23]), 
		.Z(n_6564));
	notech_and2 i_1093(.A(write_data[29]), .B(n_61215), .Z(n_29658));
	notech_reg axi_io_W_reg_24(.CP(clk), .D(n_6570), .CD(n_61806), .Q(axi_io_W
		[24]));
	notech_mux2 i_6888(.S(n_61206), .A(axi_io_W[24]), .B(writeio_data[24]), 
		.Z(n_6570));
	notech_and2 i_1094(.A(write_data[30]), .B(n_61215), .Z(n_29664));
	notech_reg axi_io_W_reg_25(.CP(clk), .D(n_6576), .CD(n_61806), .Q(axi_io_W
		[25]));
	notech_mux2 i_6896(.S(n_61206), .A(axi_io_W[25]), .B(writeio_data[25]), 
		.Z(n_6576));
	notech_and2 i_1095(.A(write_data[31]), .B(n_61215), .Z(n_29670));
	notech_reg axi_io_W_reg_26(.CP(clk), .D(n_6582), .CD(n_61804), .Q(axi_io_W
		[26]));
	notech_mux2 i_6904(.S(n_61206), .A(axi_io_W[26]), .B(writeio_data[26]), 
		.Z(n_6582));
	notech_and2 i_1101(.A(n_963), .B(n_6626), .Z(n_30150));
	notech_reg axi_io_W_reg_27(.CP(clk), .D(n_6588), .CD(n_61806), .Q(axi_io_W
		[27]));
	notech_mux2 i_6912(.S(n_61202), .A(axi_io_W[27]), .B(writeio_data[27]), 
		.Z(n_6588));
	notech_and2 i_1102(.A(n_964), .B(n_6626), .Z(n_30155));
	notech_reg axi_io_W_reg_28(.CP(clk), .D(n_6594), .CD(n_61804), .Q(axi_io_W
		[28]));
	notech_mux2 i_6920(.S(n_61202), .A(axi_io_W[28]), .B(writeio_data[28]), 
		.Z(n_6594));
	notech_and2 i_1103(.A(n_965), .B(n_6626), .Z(n_30160));
	notech_reg axi_io_W_reg_29(.CP(clk), .D(n_6600), .CD(n_61804), .Q(axi_io_W
		[29]));
	notech_mux2 i_6928(.S(n_61202), .A(axi_io_W[29]), .B(writeio_data[29]), 
		.Z(n_6600));
	notech_and2 i_1104(.A(n_966), .B(n_6626), .Z(n_30165));
	notech_reg axi_io_W_reg_30(.CP(clk), .D(n_6606), .CD(n_61806), .Q(axi_io_W
		[30]));
	notech_mux2 i_6936(.S(n_61206), .A(axi_io_W[30]), .B(writeio_data[30]), 
		.Z(n_6606));
	notech_ao3 i_57514(.A(fsm[4]), .B(n_6735), .C(n_2012), .Z(n_29767));
	notech_reg axi_io_W_reg_31(.CP(clk), .D(n_6612), .CD(n_61806), .Q(axi_io_W
		[31]));
	notech_mux2 i_6944(.S(n_61206), .A(axi_io_W[31]), .B(writeio_data[31]), 
		.Z(n_6612));
	notech_reg axi_AWVALID_reg(.CP(clk), .D(n_6618), .CD(n_61806), .Q(axi_AWVALID
		));
	notech_mux2 i_6952(.S(n_1769), .A(n_1767), .B(axi_AWVALID), .Z(n_6618)
		);
	notech_inv i_9032(.A(n_2053), .Z(n_6624));
	notech_inv i_9033(.A(n_2043), .Z(n_6625));
	notech_inv i_9034(.A(n_2025), .Z(n_6626));
	notech_inv i_9035(.A(n_222657063), .Z(n_6627));
	notech_inv i_9036(.A(n_222757064), .Z(n_6628));
	notech_inv i_9037(.A(n_61825), .Z(n_6629));
	notech_inv i_9038(.A(n_1999), .Z(n_6630));
	notech_inv i_9039(.A(n_2040), .Z(n_6631));
	notech_inv i_9040(.A(n_2015), .Z(n_6632));
	notech_inv i_9041(.A(n_59872), .Z(n_6633));
	notech_inv i_9042(.A(n_1993), .Z(n_6634));
	notech_inv i_9043(.A(n_2026), .Z(n_6635));
	notech_inv i_9044(.A(n_1742), .Z(n_6636));
	notech_inv i_9045(.A(n_971), .Z(n_6637));
	notech_inv i_9046(.A(n_978), .Z(n_6638));
	notech_inv i_9047(.A(n_981), .Z(n_6639));
	notech_inv i_9048(.A(n_984), .Z(n_6640));
	notech_inv i_9049(.A(n_987), .Z(n_6641));
	notech_inv i_9050(.A(n_2044), .Z(n_6642));
	notech_inv i_9051(.A(n_990), .Z(n_6643));
	notech_inv i_9052(.A(n_993), .Z(n_6644));
	notech_inv i_9053(.A(n_996), .Z(n_6645));
	notech_inv i_9054(.A(n_999), .Z(n_6646));
	notech_inv i_9055(.A(n_2046), .Z(n_6647));
	notech_inv i_9056(.A(n_1002), .Z(n_6648));
	notech_inv i_9057(.A(n_1005), .Z(n_6649));
	notech_inv i_9058(.A(n_1008), .Z(n_6650));
	notech_inv i_9059(.A(n_1011), .Z(n_6651));
	notech_inv i_9060(.A(n_1014), .Z(n_6652));
	notech_inv i_9061(.A(n_1017), .Z(n_6653));
	notech_inv i_9062(.A(n_1020), .Z(n_6654));
	notech_inv i_9063(.A(n_1023), .Z(n_6655));
	notech_inv i_9064(.A(n_1026), .Z(n_6656));
	notech_inv i_9065(.A(n_1029), .Z(n_6657));
	notech_inv i_9066(.A(n_1032), .Z(n_6658));
	notech_inv i_9067(.A(n_1035), .Z(n_6659));
	notech_inv i_9068(.A(n_1038), .Z(n_6660));
	notech_inv i_9069(.A(n_1041), .Z(n_6661));
	notech_inv i_9070(.A(n_1044), .Z(n_6662));
	notech_inv i_9071(.A(n_1047), .Z(n_6663));
	notech_inv i_9072(.A(n_1050), .Z(n_6664));
	notech_inv i_9073(.A(n_1053), .Z(n_6665));
	notech_inv i_9074(.A(n_1056), .Z(n_6666));
	notech_inv i_9075(.A(n_1060), .Z(n_6667));
	notech_inv i_9076(.A(n_1063), .Z(n_6668));
	notech_inv i_9077(.A(n_1068), .Z(n_6669));
	notech_inv i_9078(.A(n_1071), .Z(n_6670));
	notech_inv i_9079(.A(n_1074), .Z(n_6671));
	notech_inv i_9080(.A(n_1077), .Z(n_6672));
	notech_inv i_9081(.A(n_1080), .Z(n_6673));
	notech_inv i_9082(.A(n_1083), .Z(n_6674));
	notech_inv i_9083(.A(n_29767), .Z(n_6675));
	notech_inv i_9084(.A(n_1086), .Z(n_6676));
	notech_inv i_9085(.A(n_27143), .Z(n_6677));
	notech_inv i_9086(.A(n_1089), .Z(n_6678));
	notech_inv i_9087(.A(n_1092), .Z(n_6679));
	notech_inv i_9088(.A(n_1095), .Z(n_6680));
	notech_inv i_9089(.A(n_1098), .Z(n_6681));
	notech_inv i_9090(.A(n_1101), .Z(n_6682));
	notech_inv i_9091(.A(n_1104), .Z(n_6683));
	notech_inv i_9092(.A(n_1107), .Z(n_6684));
	notech_inv i_9093(.A(n_1110), .Z(n_6685));
	notech_inv i_9094(.A(n_1113), .Z(n_6686));
	notech_inv i_9095(.A(n_1116), .Z(n_6687));
	notech_inv i_9096(.A(n_1119), .Z(n_6688));
	notech_inv i_9097(.A(n_1122), .Z(n_6689));
	notech_inv i_9098(.A(n_1125), .Z(n_6690));
	notech_inv i_9099(.A(n_1128), .Z(n_6691));
	notech_inv i_9100(.A(n_1131), .Z(n_6692));
	notech_inv i_9101(.A(n_1134), .Z(n_6693));
	notech_inv i_9102(.A(n_1137), .Z(n_6694));
	notech_inv i_9103(.A(n_1140), .Z(n_6695));
	notech_inv i_9104(.A(n_1143), .Z(n_6696));
	notech_inv i_9105(.A(n_1146), .Z(n_6697));
	notech_inv i_9106(.A(n_1149), .Z(n_6698));
	notech_inv i_9107(.A(n_1152), .Z(n_6699));
	notech_inv i_9108(.A(n_1155), .Z(n_6700));
	notech_inv i_9109(.A(n_1158), .Z(n_6701));
	notech_inv i_9110(.A(n_1172), .Z(n_6702));
	notech_inv i_9111(.A(n_1175), .Z(n_6703));
	notech_inv i_9112(.A(n_1178), .Z(n_6704));
	notech_inv i_9113(.A(n_1181), .Z(n_6705));
	notech_inv i_9114(.A(n_1184), .Z(n_6706));
	notech_inv i_9115(.A(n_1187), .Z(n_6707));
	notech_inv i_9116(.A(n_1190), .Z(n_6708));
	notech_inv i_9117(.A(n_1193), .Z(n_6709));
	notech_inv i_9118(.A(n_1196), .Z(n_6710));
	notech_inv i_9119(.A(n_1216), .Z(n_6711));
	notech_inv i_9120(.A(burst_idx[0]), .Z(n_6712));
	notech_inv i_9121(.A(n_1223), .Z(n_6713));
	notech_inv i_9122(.A(burst_idx[1]), .Z(n_6714));
	notech_inv i_9123(.A(n_1227), .Z(n_6715));
	notech_inv i_9124(.A(n_59892), .Z(n_6716));
	notech_inv i_9125(.A(n_1230), .Z(n_6717));
	notech_inv i_9126(.A(n_1233), .Z(n_6718));
	notech_inv i_9127(.A(n_1236), .Z(n_6719));
	notech_inv i_9128(.A(n_1239), .Z(n_6720));
	notech_inv i_9129(.A(n_1242), .Z(n_6721));
	notech_inv i_9130(.A(n_1245), .Z(n_6722));
	notech_inv i_9131(.A(n_1248), .Z(n_6723));
	notech_inv i_9132(.A(n_1251), .Z(n_6724));
	notech_inv i_9133(.A(n_1254), .Z(n_6725));
	notech_inv i_9134(.A(n_1257), .Z(n_6726));
	notech_inv i_9135(.A(n_1260), .Z(n_6727));
	notech_inv i_9136(.A(n_1263), .Z(n_6728));
	notech_inv i_9137(.A(n_1266), .Z(n_6729));
	notech_inv i_9138(.A(n_1269), .Z(n_6730));
	notech_inv i_9139(.A(n_1272), .Z(n_6731));
	notech_inv i_9140(.A(n_1275), .Z(n_6732));
	notech_inv i_9141(.A(n_61873), .Z(n_6733));
	notech_inv i_9142(.A(n_1280), .Z(n_6734));
	notech_inv i_9143(.A(fsm[0]), .Z(n_6735));
	notech_inv i_9144(.A(fsm[1]), .Z(n_6736));
	notech_inv i_9145(.A(fsm[2]), .Z(n_6737));
	notech_inv i_9146(.A(fsm[4]), .Z(n_6738));
	notech_inv i_9147(.A(wf), .Z(n_6739));
	notech_inv i_9148(.A(n_28035), .Z(n_6740));
	notech_inv i_9149(.A(n_1710), .Z(n_6741));
	notech_inv i_9150(.A(\nbus_11699[0] ), .Z(n_6742));
	notech_inv i_9151(.A(\nbus_11692[0] ), .Z(n_6743));
	notech_inv i_9152(.A(\nbus_11692[32] ), .Z(n_6744));
	notech_inv i_9153(.A(\nbus_11692[64] ), .Z(n_6745));
	notech_inv i_9154(.A(\nbus_11692[96] ), .Z(n_6746));
	notech_inv i_9155(.A(n_27181), .Z(n_6747));
	notech_inv i_9156(.A(n_61206), .Z(n_6748));
	notech_inv i_9157(.A(axi_WSTRB[0]), .Z(n_6749));
	notech_inv i_9158(.A(axi_R[0]), .Z(n_6750));
	notech_inv i_9159(.A(axi_R[1]), .Z(n_6751));
	notech_inv i_9160(.A(axi_R[2]), .Z(n_6752));
	notech_inv i_9161(.A(axi_R[3]), .Z(n_6753));
	notech_inv i_9162(.A(axi_R[4]), .Z(n_6754));
	notech_inv i_9163(.A(axi_R[5]), .Z(n_6755));
	notech_inv i_9164(.A(axi_R[6]), .Z(n_6756));
	notech_inv i_9165(.A(axi_R[7]), .Z(n_6757));
	notech_inv i_9166(.A(axi_R[8]), .Z(n_6758));
	notech_inv i_9167(.A(axi_R[9]), .Z(n_6759));
	notech_inv i_9168(.A(axi_R[10]), .Z(n_6760));
	notech_inv i_9169(.A(axi_R[11]), .Z(n_6761));
	notech_inv i_9170(.A(axi_R[12]), .Z(n_6762));
	notech_inv i_9171(.A(axi_R[13]), .Z(n_6763));
	notech_inv i_9172(.A(axi_R[14]), .Z(n_6764));
	notech_inv i_9173(.A(axi_R[15]), .Z(n_6765));
	notech_inv i_9174(.A(axi_R[16]), .Z(n_6766));
	notech_inv i_9175(.A(axi_R[17]), .Z(n_6767));
	notech_inv i_9176(.A(axi_R[18]), .Z(n_6768));
	notech_inv i_9177(.A(axi_R[19]), .Z(n_6769));
	notech_inv i_9178(.A(axi_R[20]), .Z(n_6770));
	notech_inv i_9179(.A(axi_R[21]), .Z(n_6771));
	notech_inv i_9180(.A(axi_R[22]), .Z(n_6772));
	notech_inv i_9181(.A(axi_R[23]), .Z(n_6773));
	notech_inv i_9182(.A(axi_R[24]), .Z(n_6774));
	notech_inv i_9183(.A(axi_R[25]), .Z(n_6775));
	notech_inv i_9184(.A(axi_R[26]), .Z(n_6776));
	notech_inv i_9185(.A(axi_R[27]), .Z(n_6777));
	notech_inv i_9186(.A(axi_R[28]), .Z(n_6778));
	notech_inv i_9187(.A(axi_R[29]), .Z(n_6779));
	notech_inv i_9188(.A(axi_R[30]), .Z(n_6780));
	notech_inv i_9189(.A(axi_R[31]), .Z(n_6781));
	notech_inv i_9190(.A(Daddr[2]), .Z(n_6782));
	notech_inv i_9191(.A(Daddr[3]), .Z(n_6783));
	notech_inv i_9192(.A(Daddr[13]), .Z(n_6784));
	notech_inv i_9193(.A(Daddr[12]), .Z(n_6785));
	notech_inv i_9194(.A(Daddr[11]), .Z(n_6786));
	notech_inv i_9195(.A(Daddr[10]), .Z(n_6787));
	notech_inv i_9196(.A(Daddr[9]), .Z(n_6788));
	notech_inv i_9197(.A(Daddr[8]), .Z(n_6789));
	notech_inv i_9198(.A(Daddr[7]), .Z(n_6790));
	notech_inv i_9199(.A(Daddr[6]), .Z(n_6791));
	notech_inv i_9200(.A(Daddr[5]), .Z(n_6792));
	notech_inv i_9201(.A(Daddr[4]), .Z(n_6793));
	notech_inv i_9202(.A(Daddr[14]), .Z(n_6794));
	notech_inv i_9203(.A(Daddr[15]), .Z(n_6795));
	notech_inv i_9204(.A(Daddr[16]), .Z(n_6796));
	notech_inv i_9205(.A(Daddr[17]), .Z(n_6797));
	notech_inv i_9206(.A(Daddr[18]), .Z(n_6798));
	notech_inv i_9207(.A(Daddr[19]), .Z(n_6799));
	notech_inv i_9208(.A(Daddr[20]), .Z(n_6800));
	notech_inv i_9209(.A(Daddr[21]), .Z(n_6801));
	notech_inv i_9210(.A(Daddr[22]), .Z(n_6802));
	notech_inv i_9211(.A(Daddr[23]), .Z(n_6803));
	notech_inv i_9212(.A(Daddr[24]), .Z(n_6804));
	notech_inv i_9213(.A(Daddr[25]), .Z(n_6805));
	notech_inv i_9214(.A(Daddr[26]), .Z(n_6806));
	notech_inv i_9215(.A(Daddr[27]), .Z(n_6807));
	notech_inv i_9216(.A(Daddr[28]), .Z(n_6808));
	notech_inv i_9217(.A(Daddr[29]), .Z(n_6809));
	notech_inv i_9218(.A(Daddr[30]), .Z(n_6810));
	notech_inv i_9219(.A(Daddr[31]), .Z(n_6811));
	notech_inv i_9220(.A(code_wdata[0]), .Z(n_6812));
	notech_inv i_9221(.A(code_wdata[1]), .Z(n_6813));
	notech_inv i_9222(.A(code_wdata[2]), .Z(n_6814));
	notech_inv i_9223(.A(code_wdata[3]), .Z(n_6815));
	notech_inv i_9224(.A(code_wdata[4]), .Z(n_6816));
	notech_inv i_9225(.A(code_wdata[5]), .Z(n_6817));
	notech_inv i_9226(.A(code_wdata[6]), .Z(n_6818));
	notech_inv i_9227(.A(code_wdata[7]), .Z(n_6819));
	notech_inv i_9228(.A(code_addr[2]), .Z(n_6820));
	notech_inv i_9229(.A(code_addr[3]), .Z(n_6821));
	notech_inv i_9230(.A(code_addr[4]), .Z(n_6822));
	notech_inv i_9231(.A(code_addr[5]), .Z(n_6823));
	notech_inv i_9232(.A(code_addr[6]), .Z(n_6824));
	notech_inv i_9233(.A(code_addr[7]), .Z(n_6825));
	notech_inv i_9234(.A(code_addr[8]), .Z(n_6826));
	notech_inv i_9235(.A(code_addr[9]), .Z(n_6827));
	notech_inv i_9236(.A(code_addr[10]), .Z(n_6828));
	notech_inv i_9237(.A(code_addr[11]), .Z(n_6829));
	notech_inv i_9238(.A(code_addr[12]), .Z(n_6830));
	notech_inv i_9239(.A(code_addr[13]), .Z(n_6831));
	notech_inv i_9240(.A(code_addr[14]), .Z(n_6832));
	notech_inv i_9241(.A(code_addr[15]), .Z(n_6833));
	notech_inv i_9242(.A(code_addr[16]), .Z(n_6834));
	notech_inv i_9243(.A(code_addr[17]), .Z(n_6835));
	notech_inv i_9244(.A(code_addr[18]), .Z(n_6836));
	notech_inv i_9245(.A(code_addr[19]), .Z(n_6837));
	notech_inv i_9246(.A(code_addr[20]), .Z(n_6838));
	notech_inv i_9247(.A(code_addr[21]), .Z(n_6839));
	notech_inv i_9248(.A(code_addr[22]), .Z(n_6840));
	notech_inv i_9249(.A(code_addr[23]), .Z(n_6841));
	notech_inv i_9250(.A(code_addr[24]), .Z(n_6842));
	notech_inv i_9251(.A(code_addr[25]), .Z(n_6843));
	notech_inv i_9252(.A(code_addr[26]), .Z(n_6844));
	notech_inv i_9253(.A(code_addr[27]), .Z(n_6845));
	notech_inv i_9254(.A(code_addr[28]), .Z(n_6846));
	notech_inv i_9255(.A(code_addr[29]), .Z(n_6847));
	notech_inv i_9256(.A(code_addr[30]), .Z(n_6848));
	notech_inv i_9257(.A(code_addr[31]), .Z(n_6849));
	notech_inv i_9258(.A(write_data[0]), .Z(n_6850));
	notech_inv i_9259(.A(write_data[1]), .Z(n_6851));
	notech_inv i_9260(.A(write_data[2]), .Z(n_6852));
	notech_inv i_9261(.A(write_data[3]), .Z(n_6853));
	notech_inv i_9262(.A(write_data[4]), .Z(n_6854));
	notech_inv i_9263(.A(write_data[5]), .Z(n_6855));
	notech_inv i_9264(.A(write_data[6]), .Z(n_6856));
	notech_inv i_9265(.A(write_data[7]), .Z(n_6857));
	notech_inv i_9266(.A(cacheQ[0]), .Z(n_6858));
	notech_inv i_9267(.A(cacheQ[1]), .Z(n_6859));
	notech_inv i_9268(.A(cacheQ[2]), .Z(n_6860));
	notech_inv i_9269(.A(cacheQ[3]), .Z(n_6861));
	notech_inv i_9270(.A(cacheQ[4]), .Z(n_6862));
	notech_inv i_9271(.A(cacheQ[5]), .Z(n_6863));
	notech_inv i_9272(.A(cacheQ[6]), .Z(n_6864));
	notech_inv i_9273(.A(cacheQ[7]), .Z(n_6865));
	notech_inv i_9274(.A(cacheQ[8]), .Z(n_6866));
	notech_inv i_9275(.A(cacheQ[9]), .Z(n_6867));
	notech_inv i_9276(.A(cacheQ[10]), .Z(n_6868));
	notech_inv i_9277(.A(cacheQ[11]), .Z(n_6869));
	notech_inv i_9278(.A(cacheQ[12]), .Z(n_6870));
	notech_inv i_9279(.A(cacheQ[13]), .Z(n_6871));
	notech_inv i_9280(.A(cacheQ[14]), .Z(n_6872));
	notech_inv i_9281(.A(cacheQ[15]), .Z(n_6873));
	notech_inv i_9282(.A(cacheQ[16]), .Z(n_6874));
	notech_inv i_9283(.A(cacheQ[17]), .Z(n_6875));
	notech_inv i_9284(.A(cacheQ[18]), .Z(n_6876));
	notech_inv i_9285(.A(cacheQ[19]), .Z(n_6877));
	notech_inv i_9286(.A(cacheQ[20]), .Z(n_6878));
	notech_inv i_9287(.A(cacheQ[21]), .Z(n_6879));
	notech_inv i_9288(.A(cacheQ[22]), .Z(n_6880));
	notech_inv i_9289(.A(cacheQ[23]), .Z(n_6881));
	notech_inv i_9290(.A(cacheQ[24]), .Z(n_6882));
	notech_inv i_9291(.A(cacheQ[25]), .Z(n_6883));
	notech_inv i_9292(.A(cacheQ[26]), .Z(n_6884));
	notech_inv i_9293(.A(cacheQ[27]), .Z(n_6885));
	notech_inv i_9294(.A(cacheQ[28]), .Z(n_6886));
	notech_inv i_9295(.A(cacheQ[29]), .Z(n_6887));
	notech_inv i_9296(.A(cacheQ[30]), .Z(n_6888));
	notech_inv i_9297(.A(cacheQ[31]), .Z(n_6889));
	notech_inv i_9298(.A(cacheQ[32]), .Z(n_6890));
	notech_inv i_9299(.A(cacheQ[33]), .Z(n_6891));
	notech_inv i_9300(.A(cacheQ[34]), .Z(n_6892));
	notech_inv i_9301(.A(cacheQ[35]), .Z(n_6893));
	notech_inv i_9302(.A(cacheQ[36]), .Z(n_6894));
	notech_inv i_9303(.A(cacheQ[37]), .Z(n_6895));
	notech_inv i_9304(.A(cacheQ[38]), .Z(n_6896));
	notech_inv i_9305(.A(cacheQ[39]), .Z(n_6897));
	notech_inv i_9306(.A(cacheQ[40]), .Z(n_6898));
	notech_inv i_9307(.A(cacheQ[41]), .Z(n_6899));
	notech_inv i_9308(.A(cacheQ[42]), .Z(n_6900));
	notech_inv i_9309(.A(cacheQ[43]), .Z(n_6901));
	notech_inv i_9310(.A(cacheQ[44]), .Z(n_6902));
	notech_inv i_9311(.A(cacheQ[45]), .Z(n_6903));
	notech_inv i_9312(.A(cacheQ[46]), .Z(n_6904));
	notech_inv i_9313(.A(cacheQ[47]), .Z(n_6905));
	notech_inv i_9314(.A(cacheQ[48]), .Z(n_6906));
	notech_inv i_9315(.A(cacheQ[49]), .Z(n_6907));
	notech_inv i_9316(.A(cacheQ[50]), .Z(n_6908));
	notech_inv i_9317(.A(cacheQ[51]), .Z(n_6909));
	notech_inv i_9318(.A(cacheQ[52]), .Z(n_6910));
	notech_inv i_9319(.A(cacheQ[53]), .Z(n_6911));
	notech_inv i_9320(.A(cacheQ[54]), .Z(n_6912));
	notech_inv i_9321(.A(cacheQ[55]), .Z(n_6913));
	notech_inv i_9322(.A(cacheQ[56]), .Z(n_6914));
	notech_inv i_9323(.A(cacheQ[57]), .Z(n_6915));
	notech_inv i_9324(.A(cacheQ[58]), .Z(n_6916));
	notech_inv i_9325(.A(cacheQ[59]), .Z(n_6917));
	notech_inv i_9326(.A(cacheQ[60]), .Z(n_6918));
	notech_inv i_9327(.A(cacheQ[61]), .Z(n_6919));
	notech_inv i_9328(.A(cacheQ[62]), .Z(n_6920));
	notech_inv i_9329(.A(cacheQ[63]), .Z(n_6921));
	notech_inv i_9330(.A(cacheQ[96]), .Z(n_6922));
	notech_inv i_9331(.A(cacheQ[97]), .Z(n_6923));
	notech_inv i_9332(.A(cacheQ[98]), .Z(n_6924));
	notech_inv i_9333(.A(cacheQ[99]), .Z(n_6925));
	notech_inv i_9334(.A(cacheQ[100]), .Z(n_6926));
	notech_inv i_9335(.A(cacheQ[101]), .Z(n_6927));
	notech_inv i_9336(.A(cacheQ[102]), .Z(n_6928));
	notech_inv i_9337(.A(cacheQ[103]), .Z(n_6929));
	notech_inv i_9338(.A(cacheQ[104]), .Z(n_6930));
	notech_inv i_9339(.A(cacheQ[105]), .Z(n_6931));
	notech_inv i_9340(.A(cacheQ[106]), .Z(n_6932));
	notech_inv i_9341(.A(cacheQ[107]), .Z(n_6933));
	notech_inv i_9342(.A(cacheQ[108]), .Z(n_6934));
	notech_inv i_9343(.A(cacheQ[109]), .Z(n_6935));
	notech_inv i_9344(.A(cacheQ[110]), .Z(n_6936));
	notech_inv i_9345(.A(cacheQ[111]), .Z(n_6937));
	notech_inv i_9346(.A(cacheQ[112]), .Z(n_6938));
	notech_inv i_9347(.A(cacheQ[113]), .Z(n_6939));
	notech_inv i_9348(.A(cacheQ[114]), .Z(n_6940));
	notech_inv i_9349(.A(cacheQ[115]), .Z(n_6941));
	notech_inv i_9350(.A(cacheQ[116]), .Z(n_6942));
	notech_inv i_9351(.A(cacheQ[117]), .Z(n_6943));
	notech_inv i_9352(.A(cacheQ[118]), .Z(n_6944));
	notech_inv i_9353(.A(cacheQ[119]), .Z(n_6945));
	notech_inv i_9354(.A(cacheQ[120]), .Z(n_6946));
	notech_inv i_9355(.A(cacheQ[121]), .Z(n_6947));
	notech_inv i_9356(.A(cacheQ[122]), .Z(n_6948));
	notech_inv i_9357(.A(cacheQ[123]), .Z(n_6949));
	notech_inv i_9358(.A(cacheQ[124]), .Z(n_6950));
	notech_inv i_9359(.A(cacheQ[125]), .Z(n_6951));
	notech_inv i_9360(.A(cacheQ[126]), .Z(n_6952));
	notech_inv i_9361(.A(cacheQ[127]), .Z(n_6953));
	notech_inv i_9362(.A(cacheQ[128]), .Z(n_6954));
	notech_inv i_9363(.A(cacheQ[129]), .Z(n_6955));
	notech_inv i_9364(.A(cacheQ[130]), .Z(n_6956));
	notech_inv i_9365(.A(cacheQ[131]), .Z(n_6957));
	notech_inv i_9366(.A(cacheQ[132]), .Z(n_6958));
	notech_inv i_9367(.A(cacheQ[133]), .Z(n_6959));
	notech_inv i_9368(.A(cacheQ[134]), .Z(n_6960));
	notech_inv i_9369(.A(cacheQ[135]), .Z(n_6961));
	notech_inv i_9370(.A(cacheQ[136]), .Z(n_6962));
	notech_inv i_9371(.A(cacheQ[137]), .Z(n_6963));
	notech_inv i_9372(.A(cacheQ[138]), .Z(n_6964));
	notech_inv i_9373(.A(cacheQ[139]), .Z(n_6965));
	notech_inv i_9374(.A(cacheQ[140]), .Z(n_6966));
	notech_inv i_9375(.A(cacheQ[141]), .Z(n_6967));
	notech_inv i_9376(.A(cacheQ[142]), .Z(n_6968));
	notech_inv i_9377(.A(cacheQ[143]), .Z(n_6969));
	notech_inv i_9378(.A(cacheQ[144]), .Z(n_6970));
	notech_inv i_9379(.A(cacheQ[145]), .Z(n_6971));
	notech_inv i_9380(.A(cacheQ[148]), .Z(n_6972));
	notech_inv i_9381(.A(write_msk[0]), .Z(n_6973));
	notech_inv i_9382(.A(axi_AR[30]), .Z(n_6974));
	notech_inv i_9383(.A(writeio_ack), .Z(n_6975));
	notech_inv i_9384(.A(n_61806), .Z(n_6976));
	notech_inv i_9385(.A(n_26108), .Z(n_6977));
	notech_inv i_9386(.A(read_ack), .Z(n_6978));
	notech_inv i_9387(.A(code_req), .Z(n_6979));
	notech_inv i_9388(.A(read_req), .Z(n_6980));
	notech_inv i_9389(.A(code_wreq), .Z(n_6981));
	notech_inv i_9390(.A(write_req), .Z(n_6982));
	notech_inv i_9391(.A(axi_RLAST), .Z(n_6983));
	datacache datacache1(.A(cacheA), .D(cacheD), .Q(cacheQ), .M(cacheM), .WEN
		(cacheWEN), .clk(clk));
endmodule
module AWDP_INC_10(O0, fsm5_cnt);

	output [8:0] O0;
	input [8:0] fsm5_cnt;




	notech_ha2 i_8(.A(fsm5_cnt[8]), .B(n_86), .Z(O0[8]));
	notech_ha2 i_7(.A(fsm5_cnt[7]), .B(n_84), .Z(O0[7]), .CO(n_86));
	notech_ha2 i_6(.A(fsm5_cnt[6]), .B(n_82), .Z(O0[6]), .CO(n_84));
	notech_ha2 i_5(.A(fsm5_cnt[5]), .B(n_80), .Z(O0[5]), .CO(n_82));
	notech_ha2 i_4(.A(fsm5_cnt[4]), .B(n_78), .Z(O0[4]), .CO(n_80));
	notech_ha2 i_3(.A(fsm5_cnt[3]), .B(n_76), .Z(O0[3]), .CO(n_78));
	notech_ha2 i_2(.A(fsm5_cnt[2]), .B(n_74), .Z(O0[2]), .CO(n_76));
	notech_ha2 i_1(.A(fsm5_cnt[1]), .B(fsm5_cnt[0]), .Z(O0[1]), .CO(n_74));
	notech_inv i_0(.A(fsm5_cnt[0]), .Z(O0[0]));
endmodule
module cmp14_0(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_10(.A(inb[2]), .B(ina[2]), .Z(n_34));
	notech_xor2 i_9(.A(inb[4]), .B(ina[4]), .Z(n_33));
	notech_xor2 i_8(.A(inb[6]), .B(ina[6]), .Z(n_32));
	notech_xor2 i_6(.A(inb[3]), .B(ina[3]), .Z(n_31));
	notech_xor2 i_5(.A(inb[5]), .B(ina[5]), .Z(n_30));
	notech_xor2 i_4(.A(inb[7]), .B(ina[7]), .Z(n_29));
	notech_xor2 i_0(.A(inb[9]), .B(ina[9]), .Z(n_55));
	notech_xor2 i_1(.A(inb[8]), .B(ina[8]), .Z(n_56));
	notech_xor2 i_3(.A(inb[1]), .B(ina[1]), .Z(n_57));
	notech_xor2 i_7(.A(inb[0]), .B(ina[0]), .Z(n_58));
	notech_or4 i_38(.A(n_57), .B(n_56), .C(n_55), .D(ina[13]), .Z(n_61));
	notech_or4 i_37(.A(n_34), .B(n_31), .C(n_33), .D(n_30), .Z(n_66));
	notech_or4 i_39(.A(n_32), .B(n_29), .C(n_58), .D(n_66), .Z(n_67));
	notech_nor2 i_2(.A(n_67), .B(n_61), .Z(out));
endmodule
module cmp14_1(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_10(.A(inb[2]), .B(ina[2]), .Z(n_34));
	notech_xor2 i_9(.A(inb[4]), .B(ina[4]), .Z(n_33));
	notech_xor2 i_8(.A(inb[6]), .B(ina[6]), .Z(n_32));
	notech_xor2 i_6(.A(inb[3]), .B(ina[3]), .Z(n_31));
	notech_xor2 i_5(.A(inb[5]), .B(ina[5]), .Z(n_30));
	notech_xor2 i_4(.A(inb[7]), .B(ina[7]), .Z(n_29));
	notech_xor2 i_0(.A(inb[9]), .B(ina[9]), .Z(n_55));
	notech_xor2 i_1(.A(inb[8]), .B(ina[8]), .Z(n_56));
	notech_xor2 i_3(.A(inb[1]), .B(ina[1]), .Z(n_57));
	notech_xor2 i_7(.A(inb[0]), .B(ina[0]), .Z(n_58));
	notech_or4 i_38(.A(n_57), .B(n_56), .C(n_55), .D(ina[13]), .Z(n_61));
	notech_or4 i_37(.A(n_34), .B(n_31), .C(n_33), .D(n_30), .Z(n_66));
	notech_or4 i_39(.A(n_32), .B(n_29), .C(n_58), .D(n_66), .Z(n_67));
	notech_nor2 i_2(.A(n_67), .B(n_61), .Z(out));
endmodule
module cmp14_2(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_215(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100168)
		);
	notech_inv i_15298(.A(out2100168), .Z(out2));
endmodule
module cmp14_3(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_215(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100167)
		);
	notech_inv i_15279(.A(out2100167), .Z(out2));
endmodule
module cmp14_4(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_215(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100166)
		);
	notech_inv i_15260(.A(out2100166), .Z(out2));
endmodule
module cmp14_5(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_215(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100165)
		);
	notech_inv i_15241(.A(out2100165), .Z(out2));
endmodule
module cmp14_6(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_215(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100164)
		);
	notech_inv i_15222(.A(out2100164), .Z(out2));
endmodule
module cmp14_7(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_215(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100163)
		);
	notech_inv i_15203(.A(out2100163), .Z(out2));
endmodule
module cmp14_8(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_215(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100162)
		);
	notech_inv i_15184(.A(out2100162), .Z(out2));
endmodule
module cmp14_9(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_215(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out2100161)
		);
	notech_inv i_15165(.A(out2100161), .Z(out2));
endmodule
module Dtlb(clk, rstn, addr_phys, cr3, cr0, data_miss, iDaddr, pg_en, iwrite_data
		, owrite_data, iread_req, iread_ack, iwrite_req, iwrite_ack, iread_sz
		, oread_sz, iwrite_sz, owrite_sz, oread_req, oread_ack, owrite_req
		, owrite_ack, pg_fault, wr_fault, cr2, flush_tlb, cs, pt_fault, busy_ram
		, outstanding);

	input clk;
	input rstn;
	output [31:0] addr_phys;
	input [31:0] cr3;
	input [31:0] cr0;
	input [31:0] data_miss;
	input [31:0] iDaddr;
	input pg_en;
	input [31:0] iwrite_data;
	output [31:0] owrite_data;
	input iread_req;
	input iread_ack;
	input iwrite_req;
	input iwrite_ack;
	input [1:0] iread_sz;
	output [1:0] oread_sz;
	input [1:0] iwrite_sz;
	output [1:0] owrite_sz;
	output oread_req;
	output oread_ack;
	output owrite_req;
	output owrite_ack;
	output pg_fault;
	output wr_fault;
	output [31:0] cr2;
	input flush_tlb;
	input [31:0] cs;
	output pt_fault;
	input busy_ram;
	output outstanding;

	wire [3:0] fsm;
	wire [31:0] addr_miss;
	wire [31:0] wrA;
	wire [31:0] iDaddr_f;
	wire [31:0] wrD;
	wire [1:0] nx_dir;
	wire [8:0] fsm5_cnt_0;
	wire [8:0] fsm5_cnt;



	notech_inv i_15395(.A(n_62121), .Z(n_62148));
	notech_inv i_15394(.A(n_62121), .Z(n_62147));
	notech_inv i_15393(.A(n_62121), .Z(n_62146));
	notech_inv i_15391(.A(n_62121), .Z(n_62144));
	notech_inv i_15390(.A(n_62121), .Z(n_62143));
	notech_inv i_15389(.A(n_62121), .Z(n_62142));
	notech_inv i_15385(.A(n_62121), .Z(n_62139));
	notech_inv i_15384(.A(n_62121), .Z(n_62138));
	notech_inv i_15383(.A(n_62121), .Z(n_62137));
	notech_inv i_15381(.A(n_62121), .Z(n_62135));
	notech_inv i_15379(.A(n_62121), .Z(n_62134));
	notech_inv i_15378(.A(n_62121), .Z(n_62133));
	notech_inv i_15375(.A(n_62121), .Z(n_62130));
	notech_inv i_15374(.A(n_62121), .Z(n_62129));
	notech_inv i_15373(.A(n_62121), .Z(n_62128));
	notech_inv i_15370(.A(n_62121), .Z(n_62126));
	notech_inv i_15369(.A(n_62121), .Z(n_62125));
	notech_inv i_15368(.A(n_62121), .Z(n_62124));
	notech_inv i_15365(.A(clk), .Z(n_62121));
	notech_inv i_15363(.A(n_62093), .Z(n_62120));
	notech_inv i_15362(.A(n_62093), .Z(n_62119));
	notech_inv i_15361(.A(n_62093), .Z(n_62118));
	notech_inv i_15359(.A(n_62093), .Z(n_62116));
	notech_inv i_15358(.A(n_62093), .Z(n_62115));
	notech_inv i_15357(.A(n_62093), .Z(n_62114));
	notech_inv i_15353(.A(n_62093), .Z(n_62111));
	notech_inv i_15352(.A(n_62093), .Z(n_62110));
	notech_inv i_15351(.A(n_62093), .Z(n_62109));
	notech_inv i_15349(.A(n_62093), .Z(n_62107));
	notech_inv i_15347(.A(n_62093), .Z(n_62106));
	notech_inv i_15346(.A(n_62093), .Z(n_62105));
	notech_inv i_15343(.A(n_62093), .Z(n_62102));
	notech_inv i_15342(.A(n_62093), .Z(n_62101));
	notech_inv i_15341(.A(n_62093), .Z(n_62100));
	notech_inv i_15338(.A(n_62093), .Z(n_62098));
	notech_inv i_15337(.A(n_62093), .Z(n_62097));
	notech_inv i_15336(.A(n_62093), .Z(n_62096));
	notech_inv i_15333(.A(clk), .Z(n_62093));
	notech_inv i_15331(.A(n_62065), .Z(n_62092));
	notech_inv i_15330(.A(n_62065), .Z(n_62091));
	notech_inv i_15329(.A(n_62065), .Z(n_62090));
	notech_inv i_15327(.A(n_62065), .Z(n_62088));
	notech_inv i_15326(.A(n_62065), .Z(n_62087));
	notech_inv i_15325(.A(n_62065), .Z(n_62086));
	notech_inv i_15322(.A(n_62065), .Z(n_62083));
	notech_inv i_15321(.A(n_62065), .Z(n_62082));
	notech_inv i_15320(.A(n_62065), .Z(n_62081));
	notech_inv i_15318(.A(n_62065), .Z(n_62079));
	notech_inv i_15317(.A(n_62065), .Z(n_62078));
	notech_inv i_15316(.A(n_62065), .Z(n_62077));
	notech_inv i_15313(.A(n_62065), .Z(n_62074));
	notech_inv i_15311(.A(n_62065), .Z(n_62072));
	notech_inv i_15308(.A(n_62065), .Z(n_62069));
	notech_inv i_15307(.A(n_62065), .Z(n_62068));
	notech_inv i_15304(.A(clk), .Z(n_62065));
	notech_inv i_15197(.A(n_61945), .Z(n_61954));
	notech_inv i_15193(.A(n_61945), .Z(n_61950));
	notech_inv i_15189(.A(n_61945), .Z(n_61946));
	notech_inv i_15188(.A(pg_en), .Z(n_61945));
	notech_inv i_14412(.A(n_61437), .Z(n_61464));
	notech_inv i_14411(.A(n_61437), .Z(n_61463));
	notech_inv i_14410(.A(n_61437), .Z(n_61462));
	notech_inv i_14408(.A(n_61437), .Z(n_61460));
	notech_inv i_14407(.A(n_61437), .Z(n_61459));
	notech_inv i_14406(.A(n_61437), .Z(n_61458));
	notech_inv i_14403(.A(n_61437), .Z(n_61455));
	notech_inv i_14402(.A(n_61437), .Z(n_61454));
	notech_inv i_14401(.A(n_61437), .Z(n_61453));
	notech_inv i_14399(.A(n_61437), .Z(n_61451));
	notech_inv i_14398(.A(n_61437), .Z(n_61450));
	notech_inv i_14397(.A(n_61437), .Z(n_61449));
	notech_inv i_14394(.A(n_61437), .Z(n_61446));
	notech_inv i_14393(.A(n_61437), .Z(n_61445));
	notech_inv i_14392(.A(n_61437), .Z(n_61444));
	notech_inv i_14390(.A(n_61437), .Z(n_61442));
	notech_inv i_14389(.A(n_61437), .Z(n_61441));
	notech_inv i_14388(.A(n_61437), .Z(n_61440));
	notech_inv i_14385(.A(rstn), .Z(n_61437));
	notech_inv i_14384(.A(n_61409), .Z(n_61436));
	notech_inv i_14383(.A(n_61409), .Z(n_61435));
	notech_inv i_14382(.A(n_61409), .Z(n_61434));
	notech_inv i_14380(.A(n_61409), .Z(n_61432));
	notech_inv i_14379(.A(n_61409), .Z(n_61431));
	notech_inv i_14378(.A(n_61409), .Z(n_61430));
	notech_inv i_14375(.A(n_61409), .Z(n_61427));
	notech_inv i_14374(.A(n_61409), .Z(n_61426));
	notech_inv i_14373(.A(n_61409), .Z(n_61425));
	notech_inv i_14371(.A(n_61409), .Z(n_61423));
	notech_inv i_14370(.A(n_61409), .Z(n_61422));
	notech_inv i_14369(.A(n_61409), .Z(n_61421));
	notech_inv i_14366(.A(n_61409), .Z(n_61418));
	notech_inv i_14365(.A(n_61409), .Z(n_61417));
	notech_inv i_14364(.A(n_61409), .Z(n_61416));
	notech_inv i_14362(.A(n_61409), .Z(n_61414));
	notech_inv i_14361(.A(n_61409), .Z(n_61413));
	notech_inv i_14360(.A(n_61409), .Z(n_61412));
	notech_inv i_14357(.A(rstn), .Z(n_61409));
	notech_inv i_14356(.A(n_61381), .Z(n_61408));
	notech_inv i_14355(.A(n_61381), .Z(n_61407));
	notech_inv i_14354(.A(n_61381), .Z(n_61406));
	notech_inv i_14352(.A(n_61381), .Z(n_61404));
	notech_inv i_14351(.A(n_61381), .Z(n_61403));
	notech_inv i_14350(.A(n_61381), .Z(n_61402));
	notech_inv i_14347(.A(n_61381), .Z(n_61399));
	notech_inv i_14346(.A(n_61381), .Z(n_61398));
	notech_inv i_14345(.A(n_61381), .Z(n_61397));
	notech_inv i_14343(.A(n_61381), .Z(n_61395));
	notech_inv i_14342(.A(n_61381), .Z(n_61394));
	notech_inv i_14341(.A(n_61381), .Z(n_61393));
	notech_inv i_14338(.A(n_61381), .Z(n_61390));
	notech_inv i_14336(.A(n_61381), .Z(n_61388));
	notech_inv i_14333(.A(n_61381), .Z(n_61385));
	notech_inv i_14332(.A(n_61381), .Z(n_61384));
	notech_inv i_14329(.A(rstn), .Z(n_61381));
	notech_inv i_12361(.A(n_59312), .Z(n_59313));
	notech_inv i_12360(.A(n_951), .Z(n_59312));
	notech_inv i_12353(.A(n_59303), .Z(n_59304));
	notech_inv i_12352(.A(hit_tab21), .Z(n_59303));
	notech_inv i_12345(.A(n_59294), .Z(n_59295));
	notech_inv i_12344(.A(hit_tab11), .Z(n_59294));
	notech_inv i_8792(.A(n_55468), .Z(n_55469));
	notech_inv i_8791(.A(\nbus_14038[0] ), .Z(n_55468));
	notech_inv i_8784(.A(n_55459), .Z(n_55460));
	notech_inv i_8783(.A(n_1016), .Z(n_55459));
	notech_inv i_8774(.A(n_55448), .Z(n_55449));
	notech_inv i_8773(.A(n_1013), .Z(n_55448));
	notech_inv i_8679(.A(n_55355), .Z(n_55356));
	notech_inv i_8678(.A(\nbus_14029[0] ), .Z(n_55355));
	notech_inv i_8662(.A(n_55337), .Z(n_55338));
	notech_inv i_8661(.A(n_13470), .Z(n_55337));
	notech_inv i_8654(.A(n_55328), .Z(n_55329));
	notech_inv i_8653(.A(\nbus_14044[0] ), .Z(n_55328));
	notech_inv i_8649(.A(n_55317), .Z(n_55323));
	notech_inv i_8644(.A(n_55317), .Z(n_55318));
	notech_inv i_8643(.A(n_52360), .Z(n_55317));
	notech_inv i_8636(.A(n_55308), .Z(n_55309));
	notech_inv i_8635(.A(\nbus_14017[0] ), .Z(n_55308));
	notech_inv i_8628(.A(n_55299), .Z(n_55300));
	notech_inv i_8627(.A(\nbus_14036[0] ), .Z(n_55299));
	notech_inv i_8620(.A(n_55290), .Z(n_55291));
	notech_inv i_8619(.A(\nbus_14028[0] ), .Z(n_55290));
	notech_inv i_8610(.A(n_55279), .Z(n_55280));
	notech_inv i_8609(.A(\nbus_14041[0] ), .Z(n_55279));
	notech_inv i_8602(.A(n_55270), .Z(n_55271));
	notech_inv i_8601(.A(\nbus_14035[0] ), .Z(n_55270));
	notech_inv i_8594(.A(n_55259), .Z(n_55260));
	notech_inv i_8593(.A(\nbus_14034[0] ), .Z(n_55259));
	notech_inv i_8586(.A(n_55248), .Z(n_55249));
	notech_inv i_8585(.A(\nbus_14014[0] ), .Z(n_55248));
	notech_inv i_8578(.A(n_55237), .Z(n_55238));
	notech_inv i_8577(.A(\nbus_14016[0] ), .Z(n_55237));
	notech_inv i_7882(.A(n_54492), .Z(n_54493));
	notech_inv i_7881(.A(n_897), .Z(n_54492));
	notech_inv i_7764(.A(n_54280), .Z(n_54285));
	notech_inv i_7760(.A(n_54280), .Z(n_54281));
	notech_inv i_7759(.A(n_1015), .Z(n_54280));
	notech_inv i_7757(.A(n_1085), .Z(n_54277));
	notech_inv i_7756(.A(n_1085), .Z(n_54276));
	notech_inv i_7752(.A(n_1085), .Z(n_54272));
	notech_inv i_7744(.A(n_54260), .Z(n_54261));
	notech_inv i_7743(.A(n_1098), .Z(n_54260));
	notech_inv i_7736(.A(n_54251), .Z(n_54252));
	notech_inv i_7735(.A(n_1081), .Z(n_54251));
	notech_inv i_7733(.A(\nbus_14013[0] ), .Z(n_54168));
	notech_inv i_7732(.A(\nbus_14013[0] ), .Z(n_54167));
	notech_inv i_7728(.A(\nbus_14013[0] ), .Z(n_54162));
	notech_inv i_7725(.A(\nbus_14013[0] ), .Z(n_54159));
	notech_inv i_7724(.A(\nbus_14013[0] ), .Z(n_54158));
	notech_nor2 i_178(.A(hit_adr12), .B(n_576), .Z(n_574));
	notech_xor2 i_177(.A(n_13523), .B(\nnx_tab1[0] ), .Z(n_569));
	notech_or4 i_169(.A(hit_adr13), .B(hit_adr14), .C(hit_adr12), .D(hit_adr11
		), .Z(n_567));
	notech_or4 i_628(.A(n_1030), .B(n_1031), .C(\nx_tab2[1] ), .D(n_13572), 
		.Z(n_563));
	notech_or4 i_627(.A(n_1030), .B(n_1031), .C(n_13572), .D(n_13574), .Z(n_562
		));
	notech_xor2 i_176(.A(n_13569), .B(\nnx_tab2[0] ), .Z(n_558));
	notech_or4 i_170(.A(hit_adr23), .B(hit_adr24), .C(hit_adr22), .D(hit_adr21
		), .Z(n_556));
	notech_ao4 i_175(.A(hit_adr22), .B(n_1047), .C(n_13574), .D(n_1048), .Z(n_549
		));
	notech_nor2 i_127(.A(hit_adr24), .B(\nx_tab2[0] ), .Z(n_547));
	notech_nor2 i_615(.A(hit_adr23), .B(n_547), .Z(n_546));
	notech_nor2 i_174(.A(hit_adr22), .B(n_546), .Z(n_544));
	notech_or4 i_612(.A(n_1030), .B(n_1037), .C(\nx_tab1[1] ), .D(\nx_tab1[0] 
		), .Z(n_542));
	notech_or4 i_611(.A(n_1030), .B(n_1031), .C(n_13574), .D(\nx_tab2[0] ), 
		.Z(n_541));
	notech_nao3 i_173(.A(n_1016), .B(n_944), .C(n_943), .Z(n_538));
	notech_ao4 i_172(.A(iwrite_req), .B(n_61954), .C(n_943), .D(n_1052), .Z(n_536
		));
	notech_nand2 i_605(.A(\dir2[29] ), .B(n_1054), .Z(n_534));
	notech_nand2 i_602(.A(\dir2[28] ), .B(n_1054), .Z(n_533));
	notech_nand2 i_599(.A(\dir2[27] ), .B(n_1054), .Z(n_532));
	notech_nand2 i_596(.A(\dir2[26] ), .B(n_1054), .Z(n_531));
	notech_nand2 i_593(.A(\dir2[25] ), .B(n_1054), .Z(n_530));
	notech_nand2 i_590(.A(\dir2[24] ), .B(n_1054), .Z(n_529));
	notech_nand2 i_587(.A(\dir2[23] ), .B(n_1054), .Z(n_528));
	notech_nand2 i_584(.A(\dir2[22] ), .B(n_1054), .Z(n_527));
	notech_nand2 i_581(.A(\dir2[21] ), .B(n_1054), .Z(n_526));
	notech_nand2 i_578(.A(\dir2[20] ), .B(n_1054), .Z(n_525));
	notech_nand2 i_575(.A(\dir2[19] ), .B(n_1054), .Z(n_524));
	notech_nand2 i_572(.A(\dir2[18] ), .B(n_1054), .Z(n_523));
	notech_nand2 i_568(.A(\dir2[17] ), .B(n_1054), .Z(n_522));
	notech_nand2 i_565(.A(\dir2[16] ), .B(n_1054), .Z(n_521));
	notech_nand2 i_562(.A(\dir2[15] ), .B(n_1054), .Z(n_520));
	notech_nand2 i_559(.A(\dir2[14] ), .B(n_1054), .Z(n_519));
	notech_nand2 i_556(.A(\dir2[13] ), .B(n_1054), .Z(n_518));
	notech_nand2 i_553(.A(\dir2[12] ), .B(n_1054), .Z(n_517));
	notech_nand2 i_550(.A(\dir2[11] ), .B(n_1054), .Z(n_516));
	notech_nand2 i_547(.A(\dir2[10] ), .B(n_1054), .Z(n_515));
	notech_nand3 i_524(.A(n_52420), .B(iread_ack), .C(n_61954), .Z(n_494));
	notech_nao3 i_521(.A(n_406), .B(n_13438), .C(req_miss), .Z(n_491));
	notech_xor2 i_171(.A(iread_req), .B(iread_ack), .Z(n_490));
	notech_and4 i_518(.A(n_987), .B(n_13441), .C(iread_ack), .D(n_61950), .Z
		(n_489));
	notech_and4 i_517(.A(n_13440), .B(n_992), .C(n_987), .D(n_61954), .Z(n_488
		));
	notech_nao3 i_221(.A(n_61954), .B(wrA[11]), .C(n_1015), .Z(n_421));
	notech_and2 i_55(.A(n_61954), .B(n_1080), .Z(n_420));
	notech_nao3 i_218(.A(n_61950), .B(wrA[10]), .C(n_1015), .Z(n_419));
	notech_nao3 i_215(.A(n_61950), .B(wrA[9]), .C(n_1015), .Z(n_418));
	notech_nao3 i_212(.A(n_61950), .B(wrA[8]), .C(n_1015), .Z(n_417));
	notech_nao3 i_209(.A(n_61950), .B(wrA[7]), .C(n_1015), .Z(n_416));
	notech_nao3 i_206(.A(n_61950), .B(wrA[6]), .C(n_1015), .Z(n_415));
	notech_nao3 i_203(.A(n_61950), .B(wrA[5]), .C(n_54285), .Z(n_414));
	notech_nao3 i_200(.A(n_61954), .B(wrA[4]), .C(n_54285), .Z(n_413));
	notech_nao3 i_197(.A(n_61954), .B(wrA[3]), .C(n_54285), .Z(n_412));
	notech_nao3 i_194(.A(n_61954), .B(wrA[2]), .C(n_54285), .Z(n_411));
	notech_nao3 i_191(.A(n_61954), .B(wrA[1]), .C(n_54285), .Z(n_410));
	notech_nao3 i_188(.A(n_61954), .B(wrA[0]), .C(n_54285), .Z(n_409));
	notech_nand2 i_183(.A(n_994), .B(n_13447), .Z(n_408));
	notech_nand2 i_168(.A(n_984), .B(n_61954), .Z(n_407));
	notech_nand3 i_113(.A(n_981), .B(iread_req), .C(n_13473), .Z(n_406));
	notech_nor2 i_638(.A(hit_adr13), .B(n_577), .Z(n_576));
	notech_nor2 i_129(.A(hit_adr14), .B(\nx_tab1[0] ), .Z(n_577));
	notech_ao4 i_179(.A(hit_adr12), .B(n_1043), .C(n_13519), .D(n_1044), .Z(n_579
		));
	notech_or4 i_643(.A(n_1030), .B(n_1037), .C(n_13517), .D(n_13519), .Z(n_583
		));
	notech_or4 i_644(.A(n_1030), .B(n_1037), .C(n_13519), .D(\nx_tab1[0] ), 
		.Z(n_584));
	notech_or4 i_645(.A(n_1030), .B(n_1037), .C(\nx_tab1[1] ), .D(n_13517), 
		.Z(n_585));
	notech_or4 i_648(.A(n_1030), .B(n_1031), .C(\nx_tab2[1] ), .D(\nx_tab2[0] 
		), .Z(n_588));
	notech_or4 i_667(.A(data_miss[0]), .B(n_996), .C(n_13761), .D(n_13760), 
		.Z(n_607));
	notech_nor2 i_668(.A(n_609), .B(n_950), .Z(n_608));
	notech_nor2 i_101(.A(nx_dir[0]), .B(nx_dir[1]), .Z(n_609));
	notech_nand3 i_669(.A(flush_tlb), .B(n_61954), .C(n_13473), .Z(n_610));
	notech_nand2 i_673(.A(n_609), .B(n_13617), .Z(n_613));
	notech_xor2 i_180(.A(fsm[0]), .B(iwrite_ack), .Z(n_632));
	notech_or4 i_701(.A(fsm[2]), .B(fsm[1]), .C(n_986), .D(n_13760), .Z(n_636
		));
	notech_ao4 i_181(.A(n_13446), .B(n_13444), .C(fsm[0]), .D(n_13447), .Z(n_637
		));
	notech_or4 i_182(.A(hit_dir2), .B(hit_dir1), .C(n_963), .D(busy_ram), .Z
		(n_638));
	notech_nao3 i_710(.A(n_987), .B(n_13441), .C(n_641), .Z(n_640));
	notech_ao3 i_75689(.A(data_miss[5]), .B(n_964), .C(n_963), .Z(n_641));
	notech_nao3 i_712(.A(iwrite_req), .B(n_644), .C(data_miss[1]), .Z(n_643)
		);
	notech_nao3 i_123(.A(n_13733), .B(n_13734), .C(cs[0]), .Z(n_644));
	notech_or4 i_715(.A(fsm5_cnt[6]), .B(fsm5_cnt[7]), .C(fsm5_cnt[5]), .D(n_967
		), .Z(n_646));
	notech_and2 i_718(.A(hit_dir1), .B(n_650), .Z(n_649));
	notech_or4 i_184(.A(hit_tab12), .B(hit_tab11), .C(hit_tab13), .D(hit_tab14
		), .Z(n_650));
	notech_and2 i_719(.A(hit_dir2), .B(n_652), .Z(n_651));
	notech_or4 i_185(.A(hit_tab22), .B(hit_tab24), .C(hit_tab21), .D(hit_tab23
		), .Z(n_652));
	notech_nand3 i_230(.A(n_54277), .B(\tab13[10] ), .C(n_1096), .Z(n_681)
		);
	notech_nand3 i_227(.A(hit_tab11), .B(\tab11[10] ), .C(n_54276), .Z(n_684
		));
	notech_nao3 i_224(.A(hit_tab21), .B(\tab21[10] ), .C(n_1081), .Z(n_687)
		);
	notech_nand3 i_241(.A(n_54277), .B(n_1096), .C(\tab13[11] ), .Z(n_692)
		);
	notech_nand3 i_238(.A(hit_tab11), .B(n_54277), .C(\tab11[11] ), .Z(n_695
		));
	notech_nao3 i_235(.A(hit_tab21), .B(\tab21[11] ), .C(n_1081), .Z(n_698)
		);
	notech_nand3 i_252(.A(n_54277), .B(n_1096), .C(\tab13[12] ), .Z(n_703)
		);
	notech_nand3 i_249(.A(hit_tab11), .B(n_54276), .C(\tab11[12] ), .Z(n_706
		));
	notech_nao3 i_246(.A(hit_tab21), .B(\tab21[12] ), .C(n_1081), .Z(n_709)
		);
	notech_nand3 i_268(.A(n_54276), .B(n_1096), .C(\tab13[13] ), .Z(n_714)
		);
	notech_nand3 i_260(.A(hit_tab11), .B(n_54276), .C(\tab11[13] ), .Z(n_717
		));
	notech_nao3 i_257(.A(hit_tab21), .B(\tab21[13] ), .C(n_1081), .Z(n_720)
		);
	notech_nand3 i_283(.A(n_54276), .B(n_1096), .C(\tab13[14] ), .Z(n_725)
		);
	notech_nand3 i_280(.A(hit_tab11), .B(n_54276), .C(\tab11[14] ), .Z(n_728
		));
	notech_nao3 i_277(.A(hit_tab21), .B(\tab21[14] ), .C(n_1081), .Z(n_731)
		);
	notech_nand3 i_294(.A(n_54277), .B(n_1096), .C(\tab13[15] ), .Z(n_736)
		);
	notech_nand3 i_291(.A(hit_tab11), .B(n_54277), .C(\tab11[15] ), .Z(n_739
		));
	notech_nao3 i_288(.A(hit_tab21), .B(\tab21[15] ), .C(n_1081), .Z(n_742)
		);
	notech_nand3 i_305(.A(n_54277), .B(n_1096), .C(\tab13[16] ), .Z(n_747)
		);
	notech_nand3 i_302(.A(hit_tab11), .B(n_54277), .C(\tab11[16] ), .Z(n_750
		));
	notech_nao3 i_299(.A(hit_tab21), .B(\tab21[16] ), .C(n_1081), .Z(n_753)
		);
	notech_nand3 i_316(.A(n_54277), .B(n_1096), .C(\tab13[17] ), .Z(n_758)
		);
	notech_nand3 i_313(.A(hit_tab11), .B(n_54277), .C(\tab11[17] ), .Z(n_761
		));
	notech_nao3 i_310(.A(hit_tab21), .B(\tab21[17] ), .C(n_1081), .Z(n_764)
		);
	notech_nand3 i_327(.A(n_54277), .B(n_1096), .C(\tab13[18] ), .Z(n_769)
		);
	notech_nand3 i_324(.A(hit_tab11), .B(n_54277), .C(\tab11[18] ), .Z(n_772
		));
	notech_nao3 i_321(.A(hit_tab21), .B(\tab21[18] ), .C(n_1081), .Z(n_775)
		);
	notech_nand3 i_338(.A(n_54277), .B(n_1096), .C(\tab13[19] ), .Z(n_780)
		);
	notech_nand3 i_335(.A(hit_tab11), .B(n_54277), .C(\tab11[19] ), .Z(n_783
		));
	notech_nao3 i_332(.A(hit_tab21), .B(\tab21[19] ), .C(n_1081), .Z(n_786)
		);
	notech_nand3 i_349(.A(n_54276), .B(n_1096), .C(\tab13[20] ), .Z(n_791)
		);
	notech_nand3 i_346(.A(hit_tab11), .B(n_54272), .C(\tab11[20] ), .Z(n_794
		));
	notech_nao3 i_343(.A(hit_tab21), .B(\tab21[20] ), .C(n_1081), .Z(n_797)
		);
	notech_nand3 i_360(.A(n_54272), .B(n_1096), .C(\tab13[21] ), .Z(n_802)
		);
	notech_nand3 i_357(.A(n_59295), .B(n_54272), .C(\tab11[21] ), .Z(n_805)
		);
	notech_nao3 i_354(.A(n_59304), .B(\tab21[21] ), .C(n_1081), .Z(n_808));
	notech_nand3 i_371(.A(n_54272), .B(n_1096), .C(\tab13[22] ), .Z(n_813)
		);
	notech_nand3 i_368(.A(n_59295), .B(n_54272), .C(\tab11[22] ), .Z(n_816)
		);
	notech_nao3 i_365(.A(n_59304), .B(\tab21[22] ), .C(n_54252), .Z(n_819)
		);
	notech_nand3 i_382(.A(n_54272), .B(n_1096), .C(\tab13[23] ), .Z(n_824)
		);
	notech_nand3 i_379(.A(n_59295), .B(n_54272), .C(\tab11[23] ), .Z(n_827)
		);
	notech_nao3 i_376(.A(n_59304), .B(\tab21[23] ), .C(n_54252), .Z(n_830)
		);
	notech_nand3 i_393(.A(n_54272), .B(n_1096), .C(\tab13[24] ), .Z(n_835)
		);
	notech_nand3 i_390(.A(n_59295), .B(n_54272), .C(\tab11[24] ), .Z(n_838)
		);
	notech_nao3 i_387(.A(n_59304), .B(\tab21[24] ), .C(n_54252), .Z(n_841)
		);
	notech_nand3 i_404(.A(n_54272), .B(n_1096), .C(\tab13[25] ), .Z(n_846)
		);
	notech_nand3 i_401(.A(n_59295), .B(n_54276), .C(\tab11[25] ), .Z(n_849)
		);
	notech_nao3 i_398(.A(n_59304), .B(\tab21[25] ), .C(n_54252), .Z(n_852)
		);
	notech_nand3 i_415(.A(n_54276), .B(n_1096), .C(\tab13[26] ), .Z(n_857)
		);
	notech_nand3 i_412(.A(n_59295), .B(n_54276), .C(\tab11[26] ), .Z(n_860)
		);
	notech_nao3 i_409(.A(n_59304), .B(\tab21[26] ), .C(n_54252), .Z(n_863)
		);
	notech_nand3 i_426(.A(n_54276), .B(n_1096), .C(\tab13[27] ), .Z(n_868)
		);
	notech_nand3 i_423(.A(n_59295), .B(n_54276), .C(\tab11[27] ), .Z(n_871)
		);
	notech_nao3 i_420(.A(n_59304), .B(\tab21[27] ), .C(n_54252), .Z(n_874)
		);
	notech_nand3 i_437(.A(n_54272), .B(n_1096), .C(\tab13[28] ), .Z(n_879)
		);
	notech_nand3 i_434(.A(n_59295), .B(n_54272), .C(\tab11[28] ), .Z(n_882)
		);
	notech_nao3 i_431(.A(n_59304), .B(\tab21[28] ), .C(n_54252), .Z(n_885)
		);
	notech_nand3 i_448(.A(n_54272), .B(n_1096), .C(\tab13[29] ), .Z(n_890)
		);
	notech_nand3 i_445(.A(n_59295), .B(n_54276), .C(\tab11[29] ), .Z(n_893)
		);
	notech_nao3 i_442(.A(n_59304), .B(\tab21[29] ), .C(n_54252), .Z(n_896)
		);
	notech_nand3 i_121(.A(iread_ack), .B(n_61954), .C(n_13595), .Z(n_897));
	notech_ao3 i_1010(.A(n_947), .B(n_1003), .C(data_miss[1]), .Z(n_898));
	notech_and2 i_1012(.A(iwrite_sz[0]), .B(n_1015), .Z(n_899));
	notech_and2 i_1013(.A(iwrite_sz[1]), .B(n_1015), .Z(n_900));
	notech_nao3 i_519(.A(n_61954), .B(n_1076), .C(iread_ack), .Z(n_901));
	notech_nand2 i_520(.A(n_490), .B(n_13760), .Z(n_902));
	notech_and3 i_115(.A(n_981), .B(iwrite_req), .C(n_13473), .Z(n_943));
	notech_nand2 i_610(.A(iwrite_req), .B(n_1052), .Z(n_944));
	notech_or4 i_1071(.A(n_963), .B(n_989), .C(n_1034), .D(n_1008), .Z(n_945
		));
	notech_nor2 i_1059(.A(n_1004), .B(n_13750), .Z(n_946));
	notech_and3 i_166(.A(n_987), .B(iwrite_req), .C(n_13441), .Z(n_947));
	notech_and3 i_1061(.A(n_987), .B(data_miss[1]), .C(n_13441), .Z(n_948)
		);
	notech_and4 i_1062(.A(n_995), .B(data_miss[0]), .C(n_13441), .D(n_50873)
		, .Z(n_949));
	notech_nao3 i_125(.A(data_miss[0]), .B(n_13438), .C(n_996), .Z(n_950));
	notech_or4 i_122(.A(fsm[0]), .B(fsm[3]), .C(fsm[2]), .D(fsm[1]), .Z(n_951
		));
	notech_and4 i_695(.A(n_13441), .B(n_995), .C(data_miss[0]), .D(data_miss
		[5]), .Z(n_954));
	notech_or4 i_698(.A(n_957), .B(n_989), .C(n_963), .D(n_1017), .Z(n_955)
		);
	notech_or4 i_699(.A(fsm[2]), .B(fsm[1]), .C(n_13447), .D(n_13760), .Z(n_956
		));
	notech_ao4 i_98(.A(hit_dir2), .B(hit_dir1), .C(pg_fault), .D(n_981), .Z(n_957
		));
	notech_nao3 i_706(.A(n_638), .B(n_13441), .C(n_982), .Z(n_960));
	notech_nor2 i_36(.A(iwrite_req), .B(iread_req), .Z(n_963));
	notech_or2 i_713(.A(iread_req), .B(data_miss[6]), .Z(n_964));
	notech_and2 i_1087(.A(iwrite_ack), .B(n_408), .Z(n_965));
	notech_and4 i_1088(.A(fsm[0]), .B(n_987), .C(fsm5_cnt_0[0]), .D(n_13447)
		, .Z(n_966));
	notech_and2 i_111(.A(fsm5_cnt[3]), .B(fsm5_cnt[4]), .Z(n_967));
	notech_and4 i_1091(.A(fsm[0]), .B(n_987), .C(fsm5_cnt_0[1]), .D(n_13447)
		, .Z(n_968));
	notech_and4 i_1092(.A(fsm[0]), .B(n_987), .C(fsm5_cnt_0[2]), .D(n_13447)
		, .Z(n_969));
	notech_and4 i_1093(.A(fsm[0]), .B(n_987), .C(fsm5_cnt_0[3]), .D(n_13447)
		, .Z(n_970));
	notech_and4 i_1094(.A(fsm[0]), .B(n_987), .C(fsm5_cnt_0[4]), .D(n_13447)
		, .Z(n_971));
	notech_and4 i_1095(.A(fsm[0]), .B(n_987), .C(fsm5_cnt_0[5]), .D(n_13447)
		, .Z(n_972));
	notech_and4 i_1096(.A(fsm[0]), .B(n_987), .C(fsm5_cnt_0[6]), .D(n_13447)
		, .Z(n_973));
	notech_and4 i_1097(.A(fsm[0]), .B(n_987), .C(fsm5_cnt_0[7]), .D(n_13447)
		, .Z(n_974));
	notech_and4 i_1098(.A(fsm[0]), .B(n_987), .C(fsm5_cnt_0[8]), .D(n_13447)
		, .Z(n_975));
	notech_and2 i_1099(.A(iwrite_ack), .B(n_407), .Z(owrite_ack));
	notech_or2 i_75619(.A(n_651), .B(n_649), .Z(n_981));
	notech_reg fsm5_cnt_reg_0(.CP(n_62124), .D(n_10171), .CD(n_61440), .Q(fsm5_cnt
		[0]));
	notech_mux2 i_15332(.S(n_13442), .A(fsm5_cnt[0]), .B(n_966), .Z(n_10171)
		);
	notech_nand2 i_160(.A(n_13446), .B(n_13444), .Z(n_982));
	notech_reg fsm5_cnt_reg_1(.CP(n_62124), .D(n_10177), .CD(n_61440), .Q(fsm5_cnt
		[1]));
	notech_mux2 i_15340(.S(n_13442), .A(fsm5_cnt[1]), .B(n_968), .Z(n_10177)
		);
	notech_or2 i_161(.A(fsm[0]), .B(fsm[3]), .Z(n_983));
	notech_reg fsm5_cnt_reg_2(.CP(n_62124), .D(n_10183), .CD(n_61440), .Q(fsm5_cnt
		[2]));
	notech_mux2 i_15348(.S(n_13442), .A(fsm5_cnt[2]), .B(n_969), .Z(n_10183)
		);
	notech_nao3 i_38(.A(n_981), .B(n_13441), .C(n_982), .Z(n_984));
	notech_reg fsm5_cnt_reg_3(.CP(n_62124), .D(n_10189), .CD(n_61440), .Q(fsm5_cnt
		[3]));
	notech_mux2 i_15356(.S(n_13442), .A(fsm5_cnt[3]), .B(n_970), .Z(n_10189)
		);
	notech_nand2 i_47(.A(iread_ack), .B(n_61954), .Z(n_985));
	notech_reg fsm5_cnt_reg_4(.CP(n_62124), .D(n_10195), .CD(n_61440), .Q(fsm5_cnt
		[4]));
	notech_mux2 i_15364(.S(n_13442), .A(fsm5_cnt[4]), .B(n_971), .Z(n_10195)
		);
	notech_nand2 i_109(.A(fsm[0]), .B(n_13447), .Z(n_986));
	notech_reg fsm5_cnt_reg_5(.CP(n_62120), .D(n_10201), .CD(n_61436), .Q(fsm5_cnt
		[5]));
	notech_mux2 i_15372(.S(n_13442), .A(fsm5_cnt[5]), .B(n_972), .Z(n_10201)
		);
	notech_and2 i_998(.A(fsm[2]), .B(n_13444), .Z(n_987));
	notech_reg fsm5_cnt_reg_6(.CP(n_62120), .D(n_10207), .CD(n_61436), .Q(fsm5_cnt
		[6]));
	notech_mux2 i_15380(.S(n_13442), .A(fsm5_cnt[6]), .B(n_973), .Z(n_10207)
		);
	notech_reg fsm5_cnt_reg_7(.CP(n_62120), .D(n_10213), .CD(n_61436), .Q(fsm5_cnt
		[7]));
	notech_mux2 i_15388(.S(n_13442), .A(fsm5_cnt[7]), .B(n_974), .Z(n_10213)
		);
	notech_or4 i_103(.A(fsm[0]), .B(n_982), .C(fsm[3]), .D(n_13760), .Z(n_989
		));
	notech_reg fsm5_cnt_reg_8(.CP(n_62120), .D(n_10219), .CD(n_61436), .Q(fsm5_cnt
		[8]));
	notech_mux2 i_15396(.S(n_13442), .A(fsm5_cnt[8]), .B(n_975), .Z(n_10219)
		);
	notech_reg fsm_reg_0(.CP(n_62125), .D(n_10225), .CD(n_61441), .Q(fsm[0])
		);
	notech_mux2 i_15404(.S(\nbus_14033[0] ), .A(fsm[0]), .B(n_54349), .Z(n_10225
		));
	notech_reg fsm_reg_1(.CP(n_62124), .D(n_10231), .CD(n_61440), .Q(fsm[1])
		);
	notech_mux2 i_15412(.S(\nbus_14033[0] ), .A(fsm[1]), .B(n_13443), .Z(n_10231
		));
	notech_and2 i_50(.A(fsm5_cnt[8]), .B(n_646), .Z(n_992));
	notech_reg fsm_reg_2(.CP(n_62125), .D(n_10237), .CD(n_61441), .Q(fsm[2])
		);
	notech_mux2 i_15420(.S(\nbus_14033[0] ), .A(fsm[2]), .B(n_13445), .Z(n_10237
		));
	notech_nand3 i_167(.A(n_987), .B(n_13440), .C(n_61954), .Z(n_993));
	notech_reg fsm_reg_3(.CP(n_62125), .D(n_10243), .CD(n_61441), .Q(fsm[3])
		);
	notech_mux2 i_15428(.S(\nbus_14033[0] ), .A(fsm[3]), .B(n_965), .Z(n_10243
		));
	notech_nand2 i_100(.A(fsm[2]), .B(fsm[1]), .Z(n_994));
	notech_reg nx_dir_reg_0(.CP(n_62124), .D(n_10249), .CD(n_61440), .Q(nx_dir
		[0]));
	notech_mux2 i_15436(.S(n_950), .A(n_609), .B(nx_dir[0]), .Z(n_10249));
	notech_and2 i_985(.A(fsm[1]), .B(n_13446), .Z(n_995));
	notech_reg nx_dir_reg_1(.CP(n_62124), .D(n_10259), .CD(n_61440), .Q(nx_dir
		[1]));
	notech_or4 i_120(.A(fsm[0]), .B(fsm[3]), .C(n_13444), .D(fsm[2]), .Z(n_996
		));
	notech_ao3 i_15448(.A(nx_dir[1]), .B(1'b1), .C(n_13617), .Z(n_10259));
	notech_reg iDaddr_f_reg_0(.CP(n_62124), .D(n_10261), .CD(n_61440), .Q(iDaddr_f
		[0]));
	notech_mux2 i_15452(.S(n_951), .A(iDaddr[0]), .B(iDaddr_f[0]), .Z(n_10261
		));
	notech_nand3 i_44(.A(n_995), .B(data_miss[0]), .C(n_13441), .Z(n_997));
	notech_reg iDaddr_f_reg_1(.CP(n_62124), .D(n_10267), .CD(n_61440), .Q(iDaddr_f
		[1]));
	notech_mux2 i_15460(.S(n_951), .A(iDaddr[1]), .B(iDaddr_f[1]), .Z(n_10267
		));
	notech_ao4 i_980(.A(n_997), .B(data_miss[5]), .C(iwrite_ack), .D(n_994),
		 .Z(n_998));
	notech_reg iDaddr_f_reg_2(.CP(n_62124), .D(n_10273), .CD(n_61440), .Q(iDaddr_f
		[2]));
	notech_mux2 i_15468(.S(n_951), .A(iDaddr[2]), .B(iDaddr_f[2]), .Z(n_10273
		));
	notech_nand3 i_75725(.A(fsm[0]), .B(n_995), .C(n_13447), .Z(n_999));
	notech_reg iDaddr_f_reg_3(.CP(n_62119), .D(n_10279), .CD(n_61435), .Q(iDaddr_f
		[3]));
	notech_mux2 i_15476(.S(n_951), .A(iDaddr[3]), .B(iDaddr_f[3]), .Z(n_10279
		));
	notech_reg iDaddr_f_reg_4(.CP(n_62119), .D(n_10285), .CD(n_61435), .Q(iDaddr_f
		[4]));
	notech_mux2 i_15484(.S(n_951), .A(iDaddr[4]), .B(iDaddr_f[4]), .Z(n_10285
		));
	notech_reg iDaddr_f_reg_5(.CP(n_62119), .D(n_10291), .CD(n_61435), .Q(iDaddr_f
		[5]));
	notech_mux2 i_15492(.S(n_951), .A(iDaddr[5]), .B(iDaddr_f[5]), .Z(n_10291
		));
	notech_reg iDaddr_f_reg_6(.CP(n_62119), .D(n_10297), .CD(n_61435), .Q(iDaddr_f
		[6]));
	notech_mux2 i_15500(.S(n_951), .A(iDaddr[6]), .B(iDaddr_f[6]), .Z(n_10297
		));
	notech_nand2 i_75694(.A(data_miss[0]), .B(n_643), .Z(n_1003));
	notech_reg iDaddr_f_reg_7(.CP(n_62119), .D(n_10303), .CD(n_61435), .Q(iDaddr_f
		[7]));
	notech_mux2 i_15508(.S(n_951), .A(iDaddr[7]), .B(iDaddr_f[7]), .Z(n_10303
		));
	notech_or4 i_119(.A(fsm[0]), .B(fsm[3]), .C(n_13446), .D(fsm[1]), .Z(n_1004
		));
	notech_reg iDaddr_f_reg_8(.CP(n_62119), .D(n_10309), .CD(n_61435), .Q(iDaddr_f
		[8]));
	notech_mux2 i_15516(.S(n_951), .A(iDaddr[8]), .B(iDaddr_f[8]), .Z(n_10309
		));
	notech_reg iDaddr_f_reg_9(.CP(n_62119), .D(n_10315), .CD(n_61435), .Q(iDaddr_f
		[9]));
	notech_mux2 i_15524(.S(n_951), .A(iDaddr[9]), .B(iDaddr_f[9]), .Z(n_10315
		));
	notech_nand2 i_159(.A(n_640), .B(n_52377), .Z(n_1006));
	notech_reg iDaddr_f_reg_10(.CP(n_62119), .D(n_10321), .CD(n_61435), .Q(iDaddr_f
		[10]));
	notech_mux2 i_15532(.S(n_951), .A(iDaddr[10]), .B(iDaddr_f[10]), .Z(n_10321
		));
	notech_reg iDaddr_f_reg_11(.CP(n_62119), .D(n_10327), .CD(n_61435), .Q(iDaddr_f
		[11]));
	notech_mux2 i_15540(.S(n_951), .A(iDaddr[11]), .B(iDaddr_f[11]), .Z(n_10327
		));
	notech_nor2 i_37(.A(hit_dir2), .B(hit_dir1), .Z(n_1008));
	notech_reg iDaddr_f_reg_12(.CP(n_62120), .D(\addr_miss_0[2] ), .CD(n_61436
		), .Q(iDaddr_f[12]));
	notech_reg iDaddr_f_reg_13(.CP(n_62120), .D(\addr_miss_0[3] ), .CD(n_61436
		), .Q(iDaddr_f[13]));
	notech_nand3 i_978(.A(n_987), .B(n_13441), .C(n_13439), .Z(n_1010));
	notech_reg iDaddr_f_reg_14(.CP(n_62120), .D(\addr_miss_0[4] ), .CD(n_61436
		), .Q(iDaddr_f[14]));
	notech_ao4 i_975(.A(n_637), .B(iwrite_ack), .C(n_641), .D(n_1010), .Z(n_1011
		));
	notech_reg iDaddr_f_reg_15(.CP(n_62120), .D(\addr_miss_0[5] ), .CD(n_61436
		), .Q(iDaddr_f[15]));
	notech_reg iDaddr_f_reg_16(.CP(n_62120), .D(\addr_miss_0[6] ), .CD(n_61436
		), .Q(iDaddr_f[16]));
	notech_nand3 i_75718(.A(n_13446), .B(n_13444), .C(n_13440), .Z(n_1013)
		);
	notech_reg iDaddr_f_reg_17(.CP(n_62119), .D(\addr_miss_0[7] ), .CD(n_61435
		), .Q(iDaddr_f[17]));
	notech_reg iDaddr_f_reg_18(.CP(n_62119), .D(\addr_miss_0[8] ), .CD(n_61435
		), .Q(iDaddr_f[18]));
	notech_nand3 i_112(.A(fsm[2]), .B(fsm[1]), .C(n_13447), .Z(n_1015));
	notech_reg iDaddr_f_reg_19(.CP(n_62120), .D(\addr_miss_0[9] ), .CD(n_61436
		), .Q(iDaddr_f[19]));
	notech_or4 i_51(.A(n_13446), .B(n_13444), .C(fsm[3]), .D(n_13760), .Z(n_1016
		));
	notech_reg iDaddr_f_reg_20(.CP(n_62120), .D(\addr_miss_0[10] ), .CD(n_61436
		), .Q(iDaddr_f[20]));
	notech_or2 i_972(.A(busy_ram), .B(flush_tlb), .Z(n_1017));
	notech_reg iDaddr_f_reg_21(.CP(n_62125), .D(\addr_miss_0[11] ), .CD(n_61441
		), .Q(iDaddr_f[21]));
	notech_reg iDaddr_f_reg_22(.CP(n_62128), .D(n_50869), .CD(n_61444), .Q(iDaddr_f
		[22]));
	notech_reg iDaddr_f_reg_23(.CP(n_62128), .D(n_50870), .CD(n_61444), .Q(iDaddr_f
		[23]));
	notech_reg iDaddr_f_reg_24(.CP(n_62128), .D(n_50871), .CD(n_61444), .Q(iDaddr_f
		[24]));
	notech_reg iDaddr_f_reg_25(.CP(n_62128), .D(n_50872), .CD(n_61444), .Q(iDaddr_f
		[25]));
	notech_nand3 i_969(.A(n_955), .B(n_1016), .C(n_956), .Z(n_1022));
	notech_reg iDaddr_f_reg_26(.CP(n_62128), .D(n_50873), .CD(n_61444), .Q(iDaddr_f
		[26]));
	notech_nand3 i_40(.A(n_995), .B(n_13440), .C(n_61954), .Z(n_1023));
	notech_reg iDaddr_f_reg_27(.CP(n_62128), .D(n_50874), .CD(n_61444), .Q(iDaddr_f
		[27]));
	notech_reg iDaddr_f_reg_28(.CP(n_62128), .D(n_50875), .CD(n_61444), .Q(iDaddr_f
		[28]));
	notech_ao4 i_965(.A(n_994), .B(n_986), .C(n_632), .D(n_13447), .Z(n_1025
		));
	notech_reg iDaddr_f_reg_29(.CP(n_62128), .D(n_50876), .CD(n_61444), .Q(iDaddr_f
		[29]));
	notech_reg iDaddr_f_reg_30(.CP(n_62128), .D(n_50877), .CD(n_61444), .Q(iDaddr_f
		[30]));
	notech_reg iDaddr_f_reg_31(.CP(n_62129), .D(n_50878), .CD(n_61445), .Q(iDaddr_f
		[31]));
	notech_reg_set dir1_reg_0(.CP(n_62129), .D(n_10453), .SD(n_61445), .Q(\dir1[0] 
		));
	notech_mux2 i_15708(.S(\nbus_14041[0] ), .A(\dir1[0] ), .B(n_54025), .Z(n_10453
		));
	notech_reg_set dir1_reg_1(.CP(n_62129), .D(n_10459), .SD(n_61445), .Q(\dir1[1] 
		));
	notech_mux2 i_15716(.S(\nbus_14041[0] ), .A(\dir1[1] ), .B(n_54031), .Z(n_10459
		));
	notech_nao3 i_54(.A(iread_ack), .B(n_61954), .C(n_1010), .Z(n_1030));
	notech_reg_set dir1_reg_2(.CP(n_62129), .D(n_10465), .SD(n_61445), .Q(\dir1[2] 
		));
	notech_mux2 i_15724(.S(\nbus_14041[0] ), .A(\dir1[2] ), .B(n_54037), .Z(n_10465
		));
	notech_nand2 i_126(.A(hit_dir2), .B(n_13758), .Z(n_1031));
	notech_reg_set dir1_reg_3(.CP(n_62129), .D(n_10471), .SD(n_61445), .Q(\dir1[3] 
		));
	notech_mux2 i_15732(.S(\nbus_14041[0] ), .A(\dir1[3] ), .B(n_54043), .Z(n_10471
		));
	notech_or4 i_45(.A(n_1010), .B(n_1031), .C(n_13761), .D(n_13760), .Z(n_1032
		));
	notech_reg dir1_reg_4(.CP(n_62128), .D(n_10477), .CD(n_61444), .Q(\dir1[4] 
		));
	notech_mux2 i_15740(.S(\nbus_14041[0] ), .A(\dir1[4] ), .B(n_949), .Z(n_10477
		));
	notech_reg_set dir1_reg_5(.CP(n_62128), .D(n_10483), .SD(n_61444), .Q(\dir1[5] 
		));
	notech_mux2 i_15748(.S(\nbus_14041[0] ), .A(\dir1[5] ), .B(n_54055), .Z(n_10483
		));
	notech_or4 i_956(.A(pg_fault), .B(n_1017), .C(n_651), .D(n_649), .Z(n_1034
		));
	notech_reg_set dir1_reg_6(.CP(n_62129), .D(n_10489), .SD(n_61445), .Q(\dir1[6] 
		));
	notech_mux2 i_15756(.S(\nbus_14041[0] ), .A(\dir1[6] ), .B(n_54061), .Z(n_10489
		));
	notech_reg_set dir1_reg_7(.CP(n_62129), .D(n_10495), .SD(n_61445), .Q(\dir1[7] 
		));
	notech_mux2 i_15764(.S(\nbus_14041[0] ), .A(\dir1[7] ), .B(n_54067), .Z(n_10495
		));
	notech_reg_set dir1_reg_8(.CP(n_62125), .D(n_10501), .SD(n_61441), .Q(\dir1[8] 
		));
	notech_mux2 i_15772(.S(\nbus_14041[0] ), .A(\dir1[8] ), .B(n_54073), .Z(n_10501
		));
	notech_or2 i_128(.A(hit_dir2), .B(n_13758), .Z(n_1037));
	notech_reg_set dir1_reg_9(.CP(n_62125), .D(n_10507), .SD(n_61441), .Q(\dir1[9] 
		));
	notech_mux2 i_15780(.S(\nbus_14041[0] ), .A(\dir1[9] ), .B(n_54079), .Z(n_10507
		));
	notech_or4 i_48(.A(n_1010), .B(n_1037), .C(n_13761), .D(n_13760), .Z(n_1038
		));
	notech_reg_set dir1_reg_10(.CP(n_62126), .D(n_10513), .SD(n_61442), .Q(\dir1[10] 
		));
	notech_mux2 i_15788(.S(\nbus_14041[0] ), .A(\dir1[10] ), .B(n_54085), .Z
		(n_10513));
	notech_reg_set dir1_reg_11(.CP(n_62126), .D(n_10519), .SD(n_61442), .Q(\dir1[11] 
		));
	notech_mux2 i_15796(.S(\nbus_14041[0] ), .A(\dir1[11] ), .B(n_54091), .Z
		(n_10519));
	notech_reg_set dir1_reg_12(.CP(n_62125), .D(n_10525), .SD(n_61441), .Q(\dir1[12] 
		));
	notech_mux2 i_15804(.S(\nbus_14041[0] ), .A(\dir1[12] ), .B(n_54097), .Z
		(n_10525));
	notech_reg_set dir1_reg_13(.CP(n_62125), .D(n_10531), .SD(n_61441), .Q(\dir1[13] 
		));
	notech_mux2 i_15812(.S(\nbus_14041[0] ), .A(\dir1[13] ), .B(n_54103), .Z
		(n_10531));
	notech_nao3 i_102(.A(n_13440), .B(n_995), .C(hit_adr11), .Z(n_1042));
	notech_reg_set dir1_reg_14(.CP(n_62125), .D(n_10537), .SD(n_61441), .Q(\dir1[14] 
		));
	notech_mux2 i_15820(.S(\nbus_14041[0] ), .A(\dir1[14] ), .B(n_54109), .Z
		(n_10537));
	notech_nor2 i_49(.A(hit_adr13), .B(hit_adr14), .Z(n_1043));
	notech_reg_set dir1_reg_15(.CP(n_62125), .D(n_10543), .SD(n_61441), .Q(\dir1[15] 
		));
	notech_mux2 i_15828(.S(\nbus_14041[0] ), .A(\dir1[15] ), .B(n_54115), .Z
		(n_10543));
	notech_nand2 i_162(.A(n_1043), .B(n_13494), .Z(n_1044));
	notech_reg_set dir1_reg_16(.CP(n_62125), .D(n_10549), .SD(n_61441), .Q(\dir1[16] 
		));
	notech_mux2 i_15836(.S(n_55280), .A(\dir1[16] ), .B(n_54121), .Z(n_10549
		));
	notech_reg_set dir1_reg_17(.CP(n_62126), .D(n_10555), .SD(n_61442), .Q(\dir1[17] 
		));
	notech_mux2 i_15844(.S(n_55280), .A(\dir1[17] ), .B(n_54127), .Z(n_10555
		));
	notech_reg_set dir1_reg_18(.CP(n_62126), .D(n_10561), .SD(n_61442), .Q(\dir1[18] 
		));
	notech_mux2 i_15852(.S(n_55280), .A(\dir1[18] ), .B(n_54133), .Z(n_10561
		));
	notech_nor2 i_53(.A(hit_adr23), .B(hit_adr24), .Z(n_1047));
	notech_reg_set dir1_reg_19(.CP(n_62126), .D(n_10567), .SD(n_61442), .Q(\dir1[19] 
		));
	notech_mux2 i_15860(.S(n_55280), .A(\dir1[19] ), .B(n_54139), .Z(n_10567
		));
	notech_nand2 i_163(.A(n_1047), .B(n_13545), .Z(n_1048));
	notech_reg_set dir1_reg_20(.CP(n_62126), .D(n_10573), .SD(n_61442), .Q(\dir1[20] 
		));
	notech_mux2 i_15868(.S(n_55280), .A(\dir1[20] ), .B(n_54145), .Z(n_10573
		));
	notech_nao3 i_104(.A(n_13440), .B(n_995), .C(hit_adr21), .Z(n_1049));
	notech_reg_set dir1_reg_21(.CP(n_62126), .D(n_10579), .SD(n_61442), .Q(\dir1[21] 
		));
	notech_mux2 i_15876(.S(n_55280), .A(\dir1[21] ), .B(n_54151), .Z(n_10579
		));
	notech_reg_set dir1_reg_22(.CP(n_62126), .D(n_10585), .SD(n_61442), .Q(\dir1[22] 
		));
	notech_mux2 i_15884(.S(n_55280), .A(\dir1[22] ), .B(n_54157), .Z(n_10585
		));
	notech_reg_set dir1_reg_23(.CP(n_62126), .D(n_10591), .SD(n_61442), .Q(\dir1[23] 
		));
	notech_mux2 i_15892(.S(n_55280), .A(\dir1[23] ), .B(n_54163), .Z(n_10591
		));
	notech_nand2 i_68(.A(n_1015), .B(n_61946), .Z(n_1052));
	notech_reg_set dir1_reg_24(.CP(n_62126), .D(n_10597), .SD(n_61442), .Q(\dir1[24] 
		));
	notech_mux2 i_15900(.S(n_55280), .A(\dir1[24] ), .B(n_54169), .Z(n_10597
		));
	notech_reg_set dir1_reg_25(.CP(n_62126), .D(n_10603), .SD(n_61442), .Q(\dir1[25] 
		));
	notech_mux2 i_15908(.S(n_55280), .A(\dir1[25] ), .B(n_54175), .Z(n_10603
		));
	notech_ao3 i_58(.A(n_995), .B(n_13440), .C(hit_dir1), .Z(n_1054));
	notech_reg_set dir1_reg_26(.CP(n_62118), .D(n_10609), .SD(n_61434), .Q(\dir1[26] 
		));
	notech_mux2 i_15916(.S(n_55280), .A(\dir1[26] ), .B(n_54181), .Z(n_10609
		));
	notech_nand3 i_66(.A(n_995), .B(hit_dir1), .C(n_13440), .Z(n_1055));
	notech_reg_set dir1_reg_27(.CP(n_62111), .D(n_10615), .SD(n_61427), .Q(\dir1[27] 
		));
	notech_mux2 i_15924(.S(n_55280), .A(\dir1[27] ), .B(n_54187), .Z(n_10615
		));
	notech_ao4 i_942(.A(n_1055), .B(n_13468), .C(n_1013), .D(n_13681), .Z(n_1056
		));
	notech_reg_set dir1_reg_28(.CP(n_62111), .D(n_10621), .SD(n_61427), .Q(\dir1[28] 
		));
	notech_mux2 i_15932(.S(n_55280), .A(\dir1[28] ), .B(n_54193), .Z(n_10621
		));
	notech_ao4 i_941(.A(n_1055), .B(n_13467), .C(n_1013), .D(n_13682), .Z(n_1057
		));
	notech_reg_set dir1_reg_29(.CP(n_62111), .D(n_10627), .SD(n_61427), .Q(\dir1[29] 
		));
	notech_mux2 i_15940(.S(n_55280), .A(\dir1[29] ), .B(n_54199), .Z(n_10627
		));
	notech_ao4 i_940(.A(n_1055), .B(n_13466), .C(n_1013), .D(n_13683), .Z(n_1058
		));
	notech_reg_set dir1_reg_33(.CP(n_62111), .D(n_10633), .SD(n_61427), .Q(\dir1[33] 
		));
	notech_mux2 i_15948(.S(n_55280), .A(\dir1[33] ), .B(n_13470), .Z(n_10633
		));
	notech_ao4 i_939(.A(n_1055), .B(n_13465), .C(n_1013), .D(n_13684), .Z(n_1059
		));
	notech_reg_set dir2_reg_0(.CP(n_62111), .D(n_10639), .SD(n_61427), .Q(\dir2[0] 
		));
	notech_mux2 i_15956(.S(\nbus_14029[0] ), .A(\dir2[0] ), .B(n_54025), .Z(n_10639
		));
	notech_ao4 i_938(.A(n_1055), .B(n_13464), .C(n_1013), .D(n_13685), .Z(n_1060
		));
	notech_reg_set dir2_reg_1(.CP(n_62111), .D(n_10645), .SD(n_61427), .Q(\dir2[1] 
		));
	notech_mux2 i_15964(.S(\nbus_14029[0] ), .A(\dir2[1] ), .B(n_54031), .Z(n_10645
		));
	notech_ao4 i_937(.A(n_1055), .B(n_13463), .C(n_1013), .D(n_13686), .Z(n_1061
		));
	notech_reg_set dir2_reg_2(.CP(n_62110), .D(n_10651), .SD(n_61426), .Q(\dir2[2] 
		));
	notech_mux2 i_15972(.S(\nbus_14029[0] ), .A(\dir2[2] ), .B(n_54037), .Z(n_10651
		));
	notech_ao4 i_936(.A(n_1055), .B(n_13462), .C(n_1013), .D(n_13687), .Z(n_1062
		));
	notech_reg_set dir2_reg_3(.CP(n_62111), .D(n_10657), .SD(n_61427), .Q(\dir2[3] 
		));
	notech_mux2 i_15980(.S(\nbus_14029[0] ), .A(\dir2[3] ), .B(n_54043), .Z(n_10657
		));
	notech_ao4 i_935(.A(n_1055), .B(n_13461), .C(n_1013), .D(n_13688), .Z(n_1063
		));
	notech_reg dir2_reg_4(.CP(n_62111), .D(n_10663), .CD(n_61427), .Q(\dir2[4] 
		));
	notech_mux2 i_15988(.S(\nbus_14029[0] ), .A(\dir2[4] ), .B(n_949), .Z(n_10663
		));
	notech_ao4 i_934(.A(n_1055), .B(n_13460), .C(n_1013), .D(n_13689), .Z(n_1064
		));
	notech_reg_set dir2_reg_5(.CP(n_62114), .D(n_10669), .SD(n_61430), .Q(\dir2[5] 
		));
	notech_mux2 i_15996(.S(\nbus_14029[0] ), .A(\dir2[5] ), .B(n_54055), .Z(n_10669
		));
	notech_ao4 i_933(.A(n_1055), .B(n_13459), .C(n_1013), .D(n_13690), .Z(n_1065
		));
	notech_reg_set dir2_reg_6(.CP(n_62114), .D(n_10675), .SD(n_61430), .Q(\dir2[6] 
		));
	notech_mux2 i_16004(.S(\nbus_14029[0] ), .A(\dir2[6] ), .B(n_54061), .Z(n_10675
		));
	notech_ao4 i_932(.A(n_1055), .B(n_13458), .C(n_1013), .D(n_13691), .Z(n_1066
		));
	notech_reg_set dir2_reg_7(.CP(n_62114), .D(n_10681), .SD(n_61430), .Q(\dir2[7] 
		));
	notech_mux2 i_16012(.S(\nbus_14029[0] ), .A(\dir2[7] ), .B(n_54067), .Z(n_10681
		));
	notech_ao4 i_931(.A(n_1055), .B(n_13457), .C(n_1013), .D(n_13692), .Z(n_1067
		));
	notech_reg_set dir2_reg_8(.CP(n_62114), .D(n_10687), .SD(n_61430), .Q(\dir2[8] 
		));
	notech_mux2 i_16020(.S(\nbus_14029[0] ), .A(\dir2[8] ), .B(n_54073), .Z(n_10687
		));
	notech_ao4 i_930(.A(n_1055), .B(n_13456), .C(n_1013), .D(n_13693), .Z(n_1068
		));
	notech_reg_set dir2_reg_9(.CP(n_62114), .D(n_10693), .SD(n_61430), .Q(\dir2[9] 
		));
	notech_mux2 i_16028(.S(\nbus_14029[0] ), .A(\dir2[9] ), .B(n_54079), .Z(n_10693
		));
	notech_ao4 i_929(.A(n_1055), .B(n_13455), .C(n_1013), .D(n_13694), .Z(n_1069
		));
	notech_reg_set dir2_reg_10(.CP(n_62111), .D(n_10699), .SD(n_61427), .Q(\dir2[10] 
		));
	notech_mux2 i_16036(.S(\nbus_14029[0] ), .A(\dir2[10] ), .B(n_54085), .Z
		(n_10699));
	notech_ao4 i_928(.A(n_1055), .B(n_13454), .C(n_1013), .D(n_13695), .Z(n_1070
		));
	notech_reg_set dir2_reg_11(.CP(n_62111), .D(n_10705), .SD(n_61427), .Q(\dir2[11] 
		));
	notech_mux2 i_16044(.S(\nbus_14029[0] ), .A(\dir2[11] ), .B(n_54091), .Z
		(n_10705));
	notech_ao4 i_927(.A(n_1055), .B(n_13453), .C(n_1013), .D(n_13696), .Z(n_1071
		));
	notech_reg_set dir2_reg_12(.CP(n_62114), .D(n_10711), .SD(n_61430), .Q(\dir2[12] 
		));
	notech_mux2 i_16052(.S(\nbus_14029[0] ), .A(\dir2[12] ), .B(n_54097), .Z
		(n_10711));
	notech_ao4 i_926(.A(n_1055), .B(n_13452), .C(n_55449), .D(n_13697), .Z(n_1072
		));
	notech_reg_set dir2_reg_13(.CP(n_62111), .D(n_10717), .SD(n_61427), .Q(\dir2[13] 
		));
	notech_mux2 i_16060(.S(\nbus_14029[0] ), .A(\dir2[13] ), .B(n_54103), .Z
		(n_10717));
	notech_ao4 i_925(.A(n_1055), .B(n_13451), .C(n_55449), .D(n_13698), .Z(n_1073
		));
	notech_reg_set dir2_reg_14(.CP(n_62109), .D(n_10723), .SD(n_61425), .Q(\dir2[14] 
		));
	notech_mux2 i_16068(.S(\nbus_14029[0] ), .A(\dir2[14] ), .B(n_54109), .Z
		(n_10723));
	notech_ao4 i_924(.A(n_1055), .B(n_13450), .C(n_55449), .D(n_13699), .Z(n_1074
		));
	notech_reg_set dir2_reg_15(.CP(n_62109), .D(n_10729), .SD(n_61425), .Q(\dir2[15] 
		));
	notech_mux2 i_16076(.S(\nbus_14029[0] ), .A(\dir2[15] ), .B(n_54115), .Z
		(n_10729));
	notech_ao4 i_923(.A(n_1055), .B(n_13449), .C(n_55449), .D(n_13700), .Z(n_1075
		));
	notech_reg_set dir2_reg_16(.CP(n_62110), .D(n_10735), .SD(n_61426), .Q(\dir2[16] 
		));
	notech_mux2 i_16084(.S(n_55356), .A(\dir2[16] ), .B(n_54121), .Z(n_10735
		));
	notech_nand2 i_114(.A(n_406), .B(n_13606), .Z(n_1076));
	notech_reg_set dir2_reg_17(.CP(n_62109), .D(n_10741), .SD(n_61425), .Q(\dir2[17] 
		));
	notech_mux2 i_16092(.S(n_55356), .A(\dir2[17] ), .B(n_54127), .Z(n_10741
		));
	notech_reg_set dir2_reg_18(.CP(n_62109), .D(n_10747), .SD(n_61425), .Q(\dir2[18] 
		));
	notech_mux2 i_16100(.S(n_55356), .A(\dir2[18] ), .B(n_54133), .Z(n_10747
		));
	notech_reg_set dir2_reg_19(.CP(n_62109), .D(n_10753), .SD(n_61425), .Q(\dir2[19] 
		));
	notech_mux2 i_16108(.S(n_55356), .A(\dir2[19] ), .B(n_54139), .Z(n_10753
		));
	notech_reg_set dir2_reg_20(.CP(n_62109), .D(n_10759), .SD(n_61425), .Q(\dir2[20] 
		));
	notech_mux2 i_16116(.S(n_55356), .A(\dir2[20] ), .B(n_54145), .Z(n_10759
		));
	notech_nand3 i_33(.A(n_1015), .B(n_981), .C(n_61946), .Z(n_1080));
	notech_reg_set dir2_reg_21(.CP(n_62109), .D(n_10765), .SD(n_61425), .Q(\dir2[21] 
		));
	notech_mux2 i_16124(.S(n_55356), .A(\dir2[21] ), .B(n_54151), .Z(n_10765
		));
	notech_nao3 i_108(.A(n_981), .B(n_13434), .C(hit_dir1), .Z(n_1081));
	notech_reg_set dir2_reg_22(.CP(n_62109), .D(n_10771), .SD(n_61425), .Q(\dir2[22] 
		));
	notech_mux2 i_16132(.S(n_55356), .A(\dir2[22] ), .B(n_54157), .Z(n_10771
		));
	notech_reg_set dir2_reg_23(.CP(n_62110), .D(n_10777), .SD(n_61426), .Q(\dir2[23] 
		));
	notech_mux2 i_16140(.S(n_55356), .A(\dir2[23] ), .B(n_54163), .Z(n_10777
		));
	notech_reg_set dir2_reg_24(.CP(n_62110), .D(n_10783), .SD(n_61426), .Q(\dir2[24] 
		));
	notech_mux2 i_16148(.S(n_55356), .A(\dir2[24] ), .B(n_54169), .Z(n_10783
		));
	notech_nao3 i_64(.A(hit_tab22), .B(n_13759), .C(n_54252), .Z(n_1084));
	notech_reg_set dir2_reg_25(.CP(n_62110), .D(n_10789), .SD(n_61426), .Q(\dir2[25] 
		));
	notech_mux2 i_16156(.S(n_55356), .A(\dir2[25] ), .B(n_54175), .Z(n_10789
		));
	notech_nand3 i_106(.A(n_981), .B(hit_dir1), .C(n_13434), .Z(n_1085));
	notech_reg_set dir2_reg_26(.CP(n_62110), .D(n_10795), .SD(n_61426), .Q(\dir2[26] 
		));
	notech_mux2 i_16164(.S(n_55356), .A(\dir2[26] ), .B(n_54181), .Z(n_10795
		));
	notech_or4 i_67(.A(hit_tab12), .B(n_59295), .C(hit_tab13), .D(n_1085), .Z
		(n_1086));
	notech_reg_set dir2_reg_27(.CP(n_62110), .D(n_10801), .SD(n_61426), .Q(\dir2[27] 
		));
	notech_mux2 i_16172(.S(n_55356), .A(\dir2[27] ), .B(n_54187), .Z(n_10801
		));
	notech_ao4 i_909(.A(n_1086), .B(n_13515), .C(n_1084), .D(n_13544), .Z(n_1087
		));
	notech_reg_set dir2_reg_28(.CP(n_62110), .D(n_10807), .SD(n_61426), .Q(\dir2[28] 
		));
	notech_mux2 i_16180(.S(n_55356), .A(\dir2[28] ), .B(n_54193), .Z(n_10807
		));
	notech_reg_set dir2_reg_29(.CP(n_62110), .D(n_10813), .SD(n_61426), .Q(\dir2[29] 
		));
	notech_mux2 i_16188(.S(n_55356), .A(\dir2[29] ), .B(n_54199), .Z(n_10813
		));
	notech_reg_set dir2_reg_33(.CP(n_62110), .D(n_10819), .SD(n_61426), .Q(\dir2[33] 
		));
	notech_mux2 i_16196(.S(n_55356), .A(\dir2[33] ), .B(n_13470), .Z(n_10819
		));
	notech_or4 i_61(.A(hit_tab22), .B(n_59304), .C(n_54252), .D(hit_tab23), 
		.Z(n_1090));
	notech_reg_set tab21_reg_0(.CP(n_62110), .D(n_10825), .SD(n_61426), .Q(\tab21[0] 
		));
	notech_mux2 i_16204(.S(\nbus_14036[0] ), .A(\tab21[0] ), .B(n_52162), .Z
		(n_10825));
	notech_reg_set tab21_reg_1(.CP(n_62114), .D(n_10831), .SD(n_61430), .Q(\tab21[1] 
		));
	notech_mux2 i_16212(.S(\nbus_14036[0] ), .A(\tab21[1] ), .B(n_52168), .Z
		(n_10831));
	notech_or4 i_63(.A(hit_tab22), .B(n_59304), .C(n_54252), .D(n_13757), .Z
		(n_1092));
	notech_reg_set tab21_reg_2(.CP(n_62116), .D(n_10837), .SD(n_61432), .Q(\tab21[2] 
		));
	notech_mux2 i_16220(.S(\nbus_14036[0] ), .A(\tab21[2] ), .B(n_52174), .Z
		(n_10837));
	notech_ao4 i_907(.A(n_1092), .B(n_13594), .C(n_1090), .D(n_13565), .Z(n_1093
		));
	notech_reg_set tab21_reg_3(.CP(n_62116), .D(n_10843), .SD(n_61432), .Q(\tab21[3] 
		));
	notech_mux2 i_16228(.S(\nbus_14036[0] ), .A(\tab21[3] ), .B(n_52180), .Z
		(n_10843));
	notech_reg tab21_reg_4(.CP(n_62118), .D(n_10849), .CD(n_61434), .Q(\tab21[4] 
		));
	notech_mux2 i_16236(.S(\nbus_14036[0] ), .A(\tab21[4] ), .B(n_946), .Z(n_10849
		));
	notech_and4 i_911(.A(n_1093), .B(n_1087), .C(n_893), .D(n_896), .Z(n_1095
		));
	notech_reg_set tab21_reg_5(.CP(n_62116), .D(n_10855), .SD(n_61432), .Q(\tab21[5] 
		));
	notech_mux2 i_16244(.S(\nbus_14036[0] ), .A(\tab21[5] ), .B(n_52192), .Z
		(n_10855));
	notech_ao3 i_912(.A(hit_tab13), .B(n_13756), .C(n_59295), .Z(n_1096));
	notech_reg_set tab21_reg_6(.CP(n_62116), .D(n_10861), .SD(n_61432), .Q(\tab21[6] 
		));
	notech_mux2 i_16252(.S(\nbus_14036[0] ), .A(\tab21[6] ), .B(n_52198), .Z
		(n_10861));
	notech_reg_set tab21_reg_7(.CP(n_62116), .D(n_10867), .SD(n_61432), .Q(\tab21[7] 
		));
	notech_mux2 i_16260(.S(\nbus_14036[0] ), .A(\tab21[7] ), .B(n_52204), .Z
		(n_10867));
	notech_nao3 i_52(.A(n_1015), .B(n_61946), .C(n_981), .Z(n_1098));
	notech_reg_set tab21_reg_8(.CP(n_62116), .D(n_10873), .SD(n_61432), .Q(\tab21[8] 
		));
	notech_mux2 i_16268(.S(\nbus_14036[0] ), .A(\tab21[8] ), .B(n_52210), .Z
		(n_10873));
	notech_reg_set tab21_reg_9(.CP(n_62116), .D(n_10879), .SD(n_61432), .Q(\tab21[9] 
		));
	notech_mux2 i_16276(.S(\nbus_14036[0] ), .A(\tab21[9] ), .B(n_52216), .Z
		(n_10879));
	notech_nao3 i_60(.A(hit_tab12), .B(n_54276), .C(n_59295), .Z(n_1100));
	notech_reg_set tab21_reg_10(.CP(n_62116), .D(n_10885), .SD(n_61432), .Q(\tab21[10] 
		));
	notech_mux2 i_16284(.S(\nbus_14036[0] ), .A(\tab21[10] ), .B(n_52222), .Z
		(n_10885));
	notech_ao4 i_904(.A(n_1100), .B(n_13493), .C(n_1098), .D(n_13658), .Z(n_1101
		));
	notech_reg_set tab21_reg_11(.CP(n_62118), .D(n_10891), .SD(n_61434), .Q(\tab21[11] 
		));
	notech_mux2 i_16292(.S(\nbus_14036[0] ), .A(\tab21[11] ), .B(n_52228), .Z
		(n_10891));
	notech_reg_set tab21_reg_12(.CP(n_62118), .D(n_10897), .SD(n_61434), .Q(\tab21[12] 
		));
	notech_mux2 i_16300(.S(\nbus_14036[0] ), .A(\tab21[12] ), .B(n_52234), .Z
		(n_10897));
	notech_ao4 i_903(.A(n_61946), .B(n_13732), .C(n_1016), .D(n_13659), .Z(n_1103
		));
	notech_reg_set tab21_reg_13(.CP(n_62118), .D(n_10903), .SD(n_61434), .Q(\tab21[13] 
		));
	notech_mux2 i_16308(.S(\nbus_14036[0] ), .A(\tab21[13] ), .B(n_52240), .Z
		(n_10903));
	notech_reg_set tab21_reg_14(.CP(n_62118), .D(n_10909), .SD(n_61434), .Q(\tab21[14] 
		));
	notech_mux2 i_16316(.S(\nbus_14036[0] ), .A(\tab21[14] ), .B(n_52246), .Z
		(n_10909));
	notech_ao4 i_900(.A(n_1086), .B(n_13514), .C(n_1084), .D(n_13543), .Z(n_1105
		));
	notech_reg_set tab21_reg_15(.CP(n_62118), .D(n_10915), .SD(n_61434), .Q(\tab21[15] 
		));
	notech_mux2 i_16324(.S(\nbus_14036[0] ), .A(\tab21[15] ), .B(n_52252), .Z
		(n_10915));
	notech_reg_set tab21_reg_16(.CP(n_62118), .D(n_10921), .SD(n_61434), .Q(\tab21[16] 
		));
	notech_mux2 i_16332(.S(\nbus_14036[0] ), .A(\tab21[16] ), .B(n_52258), .Z
		(n_10921));
	notech_ao4 i_898(.A(n_1092), .B(n_13593), .C(n_1090), .D(n_13564), .Z(n_1107
		));
	notech_reg_set tab21_reg_17(.CP(n_62118), .D(n_10927), .SD(n_61434), .Q(\tab21[17] 
		));
	notech_mux2 i_16340(.S(n_55300), .A(\tab21[17] ), .B(n_52264), .Z(n_10927
		));
	notech_reg_set tab21_reg_18(.CP(n_62118), .D(n_10933), .SD(n_61434), .Q(\tab21[18] 
		));
	notech_mux2 i_16348(.S(n_55300), .A(\tab21[18] ), .B(n_52270), .Z(n_10933
		));
	notech_and4 i_902(.A(n_1107), .B(n_1105), .C(n_882), .D(n_885), .Z(n_1109
		));
	notech_reg_set tab21_reg_19(.CP(n_62118), .D(n_10939), .SD(n_61434), .Q(\tab21[19] 
		));
	notech_mux2 i_16356(.S(n_55300), .A(\tab21[19] ), .B(n_52276), .Z(n_10939
		));
	notech_ao4 i_895(.A(n_1100), .B(n_13492), .C(n_1098), .D(n_13656), .Z(n_1110
		));
	notech_reg_set tab21_reg_20(.CP(n_62115), .D(n_10945), .SD(n_61431), .Q(\tab21[20] 
		));
	notech_mux2 i_16364(.S(n_55300), .A(\tab21[20] ), .B(n_52282), .Z(n_10945
		));
	notech_reg_set tab21_reg_21(.CP(n_62115), .D(n_10951), .SD(n_61431), .Q(\tab21[21] 
		));
	notech_mux2 i_16372(.S(n_55300), .A(\tab21[21] ), .B(n_52288), .Z(n_10951
		));
	notech_ao4 i_894(.A(n_61946), .B(n_13731), .C(n_1016), .D(n_13657), .Z(n_1112
		));
	notech_reg_set tab21_reg_22(.CP(n_62115), .D(n_10957), .SD(n_61431), .Q(\tab21[22] 
		));
	notech_mux2 i_16380(.S(n_55300), .A(\tab21[22] ), .B(n_52294), .Z(n_10957
		));
	notech_reg_set tab21_reg_23(.CP(n_62115), .D(n_10963), .SD(n_61431), .Q(\tab21[23] 
		));
	notech_mux2 i_16388(.S(n_55300), .A(\tab21[23] ), .B(n_52300), .Z(n_10963
		));
	notech_ao4 i_891(.A(n_1086), .B(n_13513), .C(n_1084), .D(n_13542), .Z(n_1114
		));
	notech_reg_set tab21_reg_24(.CP(n_62115), .D(n_10969), .SD(n_61431), .Q(\tab21[24] 
		));
	notech_mux2 i_16396(.S(n_55300), .A(\tab21[24] ), .B(n_52306), .Z(n_10969
		));
	notech_reg_set tab21_reg_25(.CP(n_62114), .D(n_10975), .SD(n_61430), .Q(\tab21[25] 
		));
	notech_mux2 i_16404(.S(n_55300), .A(\tab21[25] ), .B(n_52312), .Z(n_10975
		));
	notech_ao4 i_889(.A(n_1092), .B(n_13592), .C(n_1090), .D(n_13563), .Z(n_1116
		));
	notech_reg_set tab21_reg_26(.CP(n_62114), .D(n_10981), .SD(n_61430), .Q(\tab21[26] 
		));
	notech_mux2 i_16412(.S(n_55300), .A(\tab21[26] ), .B(n_52318), .Z(n_10981
		));
	notech_reg_set tab21_reg_27(.CP(n_62114), .D(n_10987), .SD(n_61430), .Q(\tab21[27] 
		));
	notech_mux2 i_16420(.S(\nbus_14036[0] ), .A(\tab21[27] ), .B(n_52324), .Z
		(n_10987));
	notech_and4 i_893(.A(n_1116), .B(n_1114), .C(n_871), .D(n_874), .Z(n_1118
		));
	notech_reg_set tab21_reg_28(.CP(n_62114), .D(n_10993), .SD(n_61430), .Q(\tab21[28] 
		));
	notech_mux2 i_16428(.S(n_55300), .A(\tab21[28] ), .B(n_52330), .Z(n_10993
		));
	notech_ao4 i_886(.A(n_1100), .B(n_13491), .C(n_1098), .D(n_13654), .Z(n_1119
		));
	notech_reg_set tab21_reg_29(.CP(n_62116), .D(n_10999), .SD(n_61432), .Q(\tab21[29] 
		));
	notech_mux2 i_16436(.S(n_55300), .A(\tab21[29] ), .B(n_52336), .Z(n_10999
		));
	notech_reg tab21_reg_30(.CP(n_62115), .D(n_11005), .CD(n_61431), .Q(\tab21[30] 
		));
	notech_mux2 i_16444(.S(n_55300), .A(\tab21[30] ), .B(n_947), .Z(n_11005)
		);
	notech_ao4 i_885(.A(n_61946), .B(n_13730), .C(n_1016), .D(n_13655), .Z(n_1121
		));
	notech_reg tab21_reg_32(.CP(n_62116), .D(n_11011), .CD(n_61432), .Q(\tab21[32] 
		));
	notech_mux2 i_16452(.S(n_55300), .A(\tab21[32] ), .B(n_948), .Z(n_11011)
		);
	notech_reg_set tab21_reg_33(.CP(n_62116), .D(n_11017), .SD(n_61432), .Q(\tab21[33] 
		));
	notech_mux2 i_16460(.S(n_55300), .A(\tab21[33] ), .B(n_55323), .Z(n_11017
		));
	notech_ao4 i_882(.A(n_1086), .B(n_13512), .C(n_1084), .D(n_13541), .Z(n_1123
		));
	notech_reg hit_adr11_reg(.CP(n_62115), .D(n_11023), .CD(n_61431), .Q(hit_adr11
		));
	notech_mux2 i_16468(.S(n_945), .A(hit_add11), .B(hit_adr11), .Z(n_11023)
		);
	notech_reg_set tab12_reg_0(.CP(n_62115), .D(n_11029), .SD(n_61431), .Q(\tab12[0] 
		));
	notech_mux2 i_16476(.S(\nbus_14035[0] ), .A(\tab12[0] ), .B(n_52162), .Z
		(n_11029));
	notech_ao4 i_880(.A(n_1092), .B(n_13591), .C(n_1090), .D(n_13562), .Z(n_1125
		));
	notech_reg_set tab12_reg_1(.CP(n_62115), .D(n_11035), .SD(n_61431), .Q(\tab12[1] 
		));
	notech_mux2 i_16484(.S(\nbus_14035[0] ), .A(\tab12[1] ), .B(n_52168), .Z
		(n_11035));
	notech_reg_set tab12_reg_2(.CP(n_62115), .D(n_11041), .SD(n_61431), .Q(\tab12[2] 
		));
	notech_mux2 i_16492(.S(\nbus_14035[0] ), .A(\tab12[2] ), .B(n_52174), .Z
		(n_11041));
	notech_and4 i_884(.A(n_1125), .B(n_1123), .C(n_860), .D(n_863), .Z(n_1127
		));
	notech_reg_set tab12_reg_3(.CP(n_62115), .D(n_11047), .SD(n_61431), .Q(\tab12[3] 
		));
	notech_mux2 i_16500(.S(\nbus_14035[0] ), .A(\tab12[3] ), .B(n_52180), .Z
		(n_11047));
	notech_ao4 i_877(.A(n_1100), .B(n_13490), .C(n_1098), .D(n_13652), .Z(n_1128
		));
	notech_reg tab12_reg_4(.CP(n_62143), .D(n_11053), .CD(n_61459), .Q(\tab12[4] 
		));
	notech_mux2 i_16508(.S(\nbus_14035[0] ), .A(\tab12[4] ), .B(n_946), .Z(n_11053
		));
	notech_reg_set tab12_reg_5(.CP(n_62143), .D(n_11059), .SD(n_61459), .Q(\tab12[5] 
		));
	notech_mux2 i_16516(.S(\nbus_14035[0] ), .A(\tab12[5] ), .B(n_52192), .Z
		(n_11059));
	notech_ao4 i_876(.A(n_61946), .B(n_13729), .C(n_1016), .D(n_13653), .Z(n_1130
		));
	notech_reg_set tab12_reg_6(.CP(n_62143), .D(n_11065), .SD(n_61459), .Q(\tab12[6] 
		));
	notech_mux2 i_16524(.S(\nbus_14035[0] ), .A(\tab12[6] ), .B(n_52198), .Z
		(n_11065));
	notech_reg_set tab12_reg_7(.CP(n_62143), .D(n_11071), .SD(n_61459), .Q(\tab12[7] 
		));
	notech_mux2 i_16532(.S(\nbus_14035[0] ), .A(\tab12[7] ), .B(n_52204), .Z
		(n_11071));
	notech_ao4 i_873(.A(n_1086), .B(n_13511), .C(n_1084), .D(n_13540), .Z(n_1132
		));
	notech_reg_set tab12_reg_8(.CP(n_62143), .D(n_11077), .SD(n_61459), .Q(\tab12[8] 
		));
	notech_mux2 i_16540(.S(\nbus_14035[0] ), .A(\tab12[8] ), .B(n_52210), .Z
		(n_11077));
	notech_reg_set tab12_reg_9(.CP(n_62143), .D(n_11083), .SD(n_61459), .Q(\tab12[9] 
		));
	notech_mux2 i_16548(.S(\nbus_14035[0] ), .A(\tab12[9] ), .B(n_52216), .Z
		(n_11083));
	notech_ao4 i_871(.A(n_1092), .B(n_13590), .C(n_1090), .D(n_13561), .Z(n_1134
		));
	notech_reg_set tab12_reg_10(.CP(n_62143), .D(n_11089), .SD(n_61459), .Q(\tab12[10] 
		));
	notech_mux2 i_16556(.S(\nbus_14035[0] ), .A(\tab12[10] ), .B(n_52222), .Z
		(n_11089));
	notech_reg_set tab12_reg_11(.CP(n_62143), .D(n_11095), .SD(n_61459), .Q(\tab12[11] 
		));
	notech_mux2 i_16564(.S(\nbus_14035[0] ), .A(\tab12[11] ), .B(n_52228), .Z
		(n_11095));
	notech_and4 i_875(.A(n_1134), .B(n_1132), .C(n_849), .D(n_852), .Z(n_1136
		));
	notech_reg_set tab12_reg_12(.CP(n_62143), .D(n_11101), .SD(n_61459), .Q(\tab12[12] 
		));
	notech_mux2 i_16572(.S(\nbus_14035[0] ), .A(\tab12[12] ), .B(n_52234), .Z
		(n_11101));
	notech_ao4 i_868(.A(n_1100), .B(n_13489), .C(n_1098), .D(n_13650), .Z(n_1137
		));
	notech_reg_set tab12_reg_13(.CP(n_62144), .D(n_11107), .SD(n_61460), .Q(\tab12[13] 
		));
	notech_mux2 i_16580(.S(\nbus_14035[0] ), .A(\tab12[13] ), .B(n_52240), .Z
		(n_11107));
	notech_reg_set tab12_reg_14(.CP(n_62144), .D(n_11113), .SD(n_61460), .Q(\tab12[14] 
		));
	notech_mux2 i_16588(.S(\nbus_14035[0] ), .A(\tab12[14] ), .B(n_52246), .Z
		(n_11113));
	notech_ao4 i_867(.A(n_61946), .B(n_13728), .C(n_1016), .D(n_13651), .Z(n_1139
		));
	notech_reg_set tab12_reg_15(.CP(n_62144), .D(n_11119), .SD(n_61460), .Q(\tab12[15] 
		));
	notech_mux2 i_16596(.S(\nbus_14035[0] ), .A(\tab12[15] ), .B(n_52252), .Z
		(n_11119));
	notech_reg_set tab12_reg_16(.CP(n_62144), .D(n_11125), .SD(n_61460), .Q(\tab12[16] 
		));
	notech_mux2 i_16604(.S(\nbus_14035[0] ), .A(\tab12[16] ), .B(n_52258), .Z
		(n_11125));
	notech_ao4 i_864(.A(n_1086), .B(n_13510), .C(n_1084), .D(n_13539), .Z(n_1141
		));
	notech_reg_set tab12_reg_17(.CP(n_62144), .D(n_11131), .SD(n_61460), .Q(\tab12[17] 
		));
	notech_mux2 i_16612(.S(n_55271), .A(\tab12[17] ), .B(n_52264), .Z(n_11131
		));
	notech_reg_set tab12_reg_18(.CP(n_62143), .D(n_11137), .SD(n_61459), .Q(\tab12[18] 
		));
	notech_mux2 i_16620(.S(n_55271), .A(\tab12[18] ), .B(n_52270), .Z(n_11137
		));
	notech_ao4 i_862(.A(n_1092), .B(n_13589), .C(n_1090), .D(n_13560), .Z(n_1143
		));
	notech_reg_set tab12_reg_19(.CP(n_62143), .D(n_11143), .SD(n_61459), .Q(\tab12[19] 
		));
	notech_mux2 i_16628(.S(n_55271), .A(\tab12[19] ), .B(n_52276), .Z(n_11143
		));
	notech_reg_set tab12_reg_20(.CP(n_62144), .D(n_11149), .SD(n_61460), .Q(\tab12[20] 
		));
	notech_mux2 i_16636(.S(n_55271), .A(\tab12[20] ), .B(n_52282), .Z(n_11149
		));
	notech_and4 i_866(.A(n_1143), .B(n_1141), .C(n_838), .D(n_841), .Z(n_1145
		));
	notech_reg_set tab12_reg_21(.CP(n_62144), .D(n_11155), .SD(n_61460), .Q(\tab12[21] 
		));
	notech_mux2 i_16644(.S(n_55271), .A(\tab12[21] ), .B(n_52288), .Z(n_11155
		));
	notech_ao4 i_859(.A(n_1100), .B(n_13488), .C(n_1098), .D(n_13648), .Z(n_1146
		));
	notech_reg_set tab12_reg_22(.CP(n_62139), .D(n_11161), .SD(n_61455), .Q(\tab12[22] 
		));
	notech_mux2 i_16652(.S(n_55271), .A(\tab12[22] ), .B(n_52294), .Z(n_11161
		));
	notech_reg_set tab12_reg_23(.CP(n_62139), .D(n_11167), .SD(n_61455), .Q(\tab12[23] 
		));
	notech_mux2 i_16660(.S(n_55271), .A(\tab12[23] ), .B(n_52300), .Z(n_11167
		));
	notech_ao4 i_858(.A(n_61946), .B(n_13727), .C(n_1016), .D(n_13649), .Z(n_1148
		));
	notech_reg_set tab12_reg_24(.CP(n_62142), .D(n_11173), .SD(n_61458), .Q(\tab12[24] 
		));
	notech_mux2 i_16668(.S(n_55271), .A(\tab12[24] ), .B(n_52306), .Z(n_11173
		));
	notech_reg_set tab12_reg_25(.CP(n_62142), .D(n_11179), .SD(n_61458), .Q(\tab12[25] 
		));
	notech_mux2 i_16676(.S(n_55271), .A(\tab12[25] ), .B(n_52312), .Z(n_11179
		));
	notech_ao4 i_855(.A(n_1086), .B(n_13509), .C(n_1084), .D(n_13538), .Z(n_1150
		));
	notech_reg_set tab12_reg_26(.CP(n_62139), .D(n_11185), .SD(n_61455), .Q(\tab12[26] 
		));
	notech_mux2 i_16684(.S(n_55271), .A(\tab12[26] ), .B(n_52318), .Z(n_11185
		));
	notech_reg_set tab12_reg_27(.CP(n_62139), .D(n_11191), .SD(n_61455), .Q(\tab12[27] 
		));
	notech_mux2 i_16692(.S(\nbus_14035[0] ), .A(\tab12[27] ), .B(n_52324), .Z
		(n_11191));
	notech_ao4 i_853(.A(n_1092), .B(n_13588), .C(n_1090), .D(n_13559), .Z(n_1152
		));
	notech_reg_set tab12_reg_28(.CP(n_62139), .D(n_11197), .SD(n_61455), .Q(\tab12[28] 
		));
	notech_mux2 i_16700(.S(n_55271), .A(\tab12[28] ), .B(n_52330), .Z(n_11197
		));
	notech_reg_set tab12_reg_29(.CP(n_62139), .D(n_11203), .SD(n_61455), .Q(\tab12[29] 
		));
	notech_mux2 i_16708(.S(n_55271), .A(\tab12[29] ), .B(n_52336), .Z(n_11203
		));
	notech_and4 i_857(.A(n_1152), .B(n_1150), .C(n_827), .D(n_830), .Z(n_1154
		));
	notech_reg tab12_reg_30(.CP(n_62139), .D(n_11209), .CD(n_61455), .Q(\tab12[30] 
		));
	notech_mux2 i_16716(.S(n_55271), .A(\tab12[30] ), .B(n_947), .Z(n_11209)
		);
	notech_ao4 i_850(.A(n_1100), .B(n_13487), .C(n_1098), .D(n_13646), .Z(n_1155
		));
	notech_reg tab12_reg_32(.CP(n_62142), .D(n_11215), .CD(n_61458), .Q(\tab12[32] 
		));
	notech_mux2 i_16724(.S(n_55271), .A(\tab12[32] ), .B(n_948), .Z(n_11215)
		);
	notech_reg_set tab12_reg_33(.CP(n_62142), .D(n_11221), .SD(n_61458), .Q(\tab12[33] 
		));
	notech_mux2 i_16732(.S(n_55271), .A(\tab12[33] ), .B(n_55323), .Z(n_11221
		));
	notech_ao4 i_849(.A(n_61946), .B(n_13726), .C(n_1016), .D(n_13647), .Z(n_1157
		));
	notech_reg hit_adr12_reg(.CP(n_62142), .D(n_11227), .CD(n_61458), .Q(hit_adr12
		));
	notech_mux2 i_16740(.S(n_945), .A(hit_add12), .B(hit_adr12), .Z(n_11227)
		);
	notech_reg_set tab13_reg_0(.CP(n_62142), .D(n_11233), .SD(n_61458), .Q(\tab13[0] 
		));
	notech_mux2 i_16748(.S(\nbus_14014[0] ), .A(\tab13[0] ), .B(n_52162), .Z
		(n_11233));
	notech_ao4 i_846(.A(n_1086), .B(n_13508), .C(n_1084), .D(n_13537), .Z(n_1159
		));
	notech_reg_set tab13_reg_1(.CP(n_62142), .D(n_11239), .SD(n_61458), .Q(\tab13[1] 
		));
	notech_mux2 i_16756(.S(\nbus_14014[0] ), .A(\tab13[1] ), .B(n_52168), .Z
		(n_11239));
	notech_reg_set tab13_reg_2(.CP(n_62142), .D(n_11245), .SD(n_61458), .Q(\tab13[2] 
		));
	notech_mux2 i_16764(.S(\nbus_14014[0] ), .A(\tab13[2] ), .B(n_52174), .Z
		(n_11245));
	notech_ao4 i_844(.A(n_1092), .B(n_13587), .C(n_1090), .D(n_13558), .Z(n_1161
		));
	notech_reg_set tab13_reg_3(.CP(n_62142), .D(n_11251), .SD(n_61458), .Q(\tab13[3] 
		));
	notech_mux2 i_16772(.S(\nbus_14014[0] ), .A(\tab13[3] ), .B(n_52180), .Z
		(n_11251));
	notech_reg tab13_reg_4(.CP(n_62142), .D(n_11257), .CD(n_61458), .Q(\tab13[4] 
		));
	notech_mux2 i_16780(.S(\nbus_14014[0] ), .A(\tab13[4] ), .B(n_946), .Z(n_11257
		));
	notech_and4 i_848(.A(n_1161), .B(n_1159), .C(n_816), .D(n_819), .Z(n_1163
		));
	notech_reg_set tab13_reg_5(.CP(n_62142), .D(n_11263), .SD(n_61458), .Q(\tab13[5] 
		));
	notech_mux2 i_16788(.S(\nbus_14014[0] ), .A(\tab13[5] ), .B(n_52192), .Z
		(n_11263));
	notech_ao4 i_841(.A(n_1100), .B(n_13486), .C(n_1098), .D(n_13644), .Z(n_1164
		));
	notech_reg_set tab13_reg_6(.CP(n_62144), .D(n_11269), .SD(n_61460), .Q(\tab13[6] 
		));
	notech_mux2 i_16796(.S(\nbus_14014[0] ), .A(\tab13[6] ), .B(n_52198), .Z
		(n_11269));
	notech_reg_set tab13_reg_7(.CP(n_62147), .D(n_11275), .SD(n_61463), .Q(\tab13[7] 
		));
	notech_mux2 i_16804(.S(\nbus_14014[0] ), .A(\tab13[7] ), .B(n_52204), .Z
		(n_11275));
	notech_ao4 i_840(.A(n_61946), .B(n_13725), .C(n_1016), .D(n_13645), .Z(n_1166
		));
	notech_reg_set tab13_reg_8(.CP(n_62147), .D(n_11281), .SD(n_61463), .Q(\tab13[8] 
		));
	notech_mux2 i_16812(.S(\nbus_14014[0] ), .A(\tab13[8] ), .B(n_52210), .Z
		(n_11281));
	notech_reg_set tab13_reg_9(.CP(n_62148), .D(n_11287), .SD(n_61464), .Q(\tab13[9] 
		));
	notech_mux2 i_16820(.S(\nbus_14014[0] ), .A(\tab13[9] ), .B(n_52216), .Z
		(n_11287));
	notech_ao4 i_837(.A(n_1086), .B(n_13507), .C(n_1084), .D(n_13536), .Z(n_1168
		));
	notech_reg_set tab13_reg_10(.CP(n_62148), .D(n_11293), .SD(n_61464), .Q(\tab13[10] 
		));
	notech_mux2 i_16828(.S(\nbus_14014[0] ), .A(\tab13[10] ), .B(n_52222), .Z
		(n_11293));
	notech_reg_set tab13_reg_11(.CP(n_62147), .D(n_11299), .SD(n_61463), .Q(\tab13[11] 
		));
	notech_mux2 i_16836(.S(\nbus_14014[0] ), .A(\tab13[11] ), .B(n_52228), .Z
		(n_11299));
	notech_ao4 i_835(.A(n_1092), .B(n_13586), .C(n_1090), .D(n_13557), .Z(n_1170
		));
	notech_reg_set tab13_reg_12(.CP(n_62147), .D(n_11305), .SD(n_61463), .Q(\tab13[12] 
		));
	notech_mux2 i_16844(.S(\nbus_14014[0] ), .A(\tab13[12] ), .B(n_52234), .Z
		(n_11305));
	notech_reg_set tab13_reg_13(.CP(n_62147), .D(n_11311), .SD(n_61463), .Q(\tab13[13] 
		));
	notech_mux2 i_16852(.S(\nbus_14014[0] ), .A(\tab13[13] ), .B(n_52240), .Z
		(n_11311));
	notech_and4 i_839(.A(n_1170), .B(n_1168), .C(n_805), .D(n_808), .Z(n_1172
		));
	notech_reg_set tab13_reg_14(.CP(n_62147), .D(n_11317), .SD(n_61463), .Q(\tab13[14] 
		));
	notech_mux2 i_16860(.S(\nbus_14014[0] ), .A(\tab13[14] ), .B(n_52246), .Z
		(n_11317));
	notech_ao4 i_832(.A(n_1100), .B(n_13485), .C(n_1098), .D(n_13642), .Z(n_1173
		));
	notech_reg_set tab13_reg_15(.CP(n_62147), .D(n_11323), .SD(n_61463), .Q(\tab13[15] 
		));
	notech_mux2 i_16868(.S(\nbus_14014[0] ), .A(\tab13[15] ), .B(n_52252), .Z
		(n_11323));
	notech_reg_set tab13_reg_16(.CP(n_62148), .D(n_11329), .SD(n_61464), .Q(\tab13[16] 
		));
	notech_mux2 i_16876(.S(\nbus_14014[0] ), .A(\tab13[16] ), .B(n_52258), .Z
		(n_11329));
	notech_ao4 i_831(.A(n_61946), .B(n_13724), .C(n_1016), .D(n_13643), .Z(n_1175
		));
	notech_reg_set tab13_reg_17(.CP(n_62148), .D(n_11335), .SD(n_61464), .Q(\tab13[17] 
		));
	notech_mux2 i_16884(.S(n_55249), .A(\tab13[17] ), .B(n_52264), .Z(n_11335
		));
	notech_reg_set tab13_reg_18(.CP(n_62148), .D(n_11341), .SD(n_61464), .Q(\tab13[18] 
		));
	notech_mux2 i_16892(.S(n_55249), .A(\tab13[18] ), .B(n_52270), .Z(n_11341
		));
	notech_ao4 i_828(.A(n_1086), .B(n_13506), .C(n_1084), .D(n_13535), .Z(n_1177
		));
	notech_reg_set tab13_reg_19(.CP(n_62148), .D(n_11347), .SD(n_61464), .Q(\tab13[19] 
		));
	notech_mux2 i_16900(.S(n_55249), .A(\tab13[19] ), .B(n_52276), .Z(n_11347
		));
	notech_reg_set tab13_reg_20(.CP(n_62148), .D(n_11353), .SD(n_61464), .Q(\tab13[20] 
		));
	notech_mux2 i_16908(.S(n_55249), .A(\tab13[20] ), .B(n_52282), .Z(n_11353
		));
	notech_ao4 i_826(.A(n_1092), .B(n_13585), .C(n_1090), .D(n_13556), .Z(n_1179
		));
	notech_reg_set tab13_reg_21(.CP(n_62148), .D(n_11359), .SD(n_61464), .Q(\tab13[21] 
		));
	notech_mux2 i_16916(.S(n_55249), .A(\tab13[21] ), .B(n_52288), .Z(n_11359
		));
	notech_reg_set tab13_reg_22(.CP(n_62148), .D(n_11365), .SD(n_61464), .Q(\tab13[22] 
		));
	notech_mux2 i_16924(.S(n_55249), .A(\tab13[22] ), .B(n_52294), .Z(n_11365
		));
	notech_and4 i_830(.A(n_1179), .B(n_1177), .C(n_794), .D(n_797), .Z(n_1181
		));
	notech_reg_set tab13_reg_23(.CP(n_62148), .D(n_11371), .SD(n_61464), .Q(\tab13[23] 
		));
	notech_mux2 i_16932(.S(n_55249), .A(\tab13[23] ), .B(n_52300), .Z(n_11371
		));
	notech_ao4 i_823(.A(n_1100), .B(n_13484), .C(n_1098), .D(n_13640), .Z(n_1182
		));
	notech_reg_set tab13_reg_24(.CP(n_62148), .D(n_11377), .SD(n_61464), .Q(\tab13[24] 
		));
	notech_mux2 i_16940(.S(n_55249), .A(\tab13[24] ), .B(n_52306), .Z(n_11377
		));
	notech_reg_set tab13_reg_25(.CP(n_62146), .D(n_11383), .SD(n_61462), .Q(\tab13[25] 
		));
	notech_mux2 i_16948(.S(n_55249), .A(\tab13[25] ), .B(n_52312), .Z(n_11383
		));
	notech_ao4 i_822(.A(n_61946), .B(n_13723), .C(n_55460), .D(n_13641), .Z(n_1184
		));
	notech_reg_set tab13_reg_26(.CP(n_62146), .D(n_11389), .SD(n_61462), .Q(\tab13[26] 
		));
	notech_mux2 i_16956(.S(n_55249), .A(\tab13[26] ), .B(n_52318), .Z(n_11389
		));
	notech_reg_set tab13_reg_27(.CP(n_62146), .D(n_11395), .SD(n_61462), .Q(\tab13[27] 
		));
	notech_mux2 i_16964(.S(\nbus_14014[0] ), .A(\tab13[27] ), .B(n_52324), .Z
		(n_11395));
	notech_ao4 i_819(.A(n_1086), .B(n_13505), .C(n_1084), .D(n_13534), .Z(n_1186
		));
	notech_reg_set tab13_reg_28(.CP(n_62146), .D(n_11401), .SD(n_61462), .Q(\tab13[28] 
		));
	notech_mux2 i_16972(.S(n_55249), .A(\tab13[28] ), .B(n_52330), .Z(n_11401
		));
	notech_reg_set tab13_reg_29(.CP(n_62146), .D(n_11407), .SD(n_61462), .Q(\tab13[29] 
		));
	notech_mux2 i_16980(.S(n_55249), .A(\tab13[29] ), .B(n_52336), .Z(n_11407
		));
	notech_ao4 i_817(.A(n_1092), .B(n_13584), .C(n_1090), .D(n_13555), .Z(n_1188
		));
	notech_reg tab13_reg_30(.CP(n_62144), .D(n_11413), .CD(n_61460), .Q(\tab13[30] 
		));
	notech_mux2 i_16988(.S(n_55249), .A(\tab13[30] ), .B(n_947), .Z(n_11413)
		);
	notech_reg tab13_reg_32(.CP(n_62144), .D(n_11419), .CD(n_61460), .Q(\tab13[32] 
		));
	notech_mux2 i_16996(.S(n_55249), .A(\tab13[32] ), .B(n_948), .Z(n_11419)
		);
	notech_and4 i_821(.A(n_1188), .B(n_1186), .C(n_783), .D(n_786), .Z(n_1190
		));
	notech_reg_set tab13_reg_33(.CP(n_62146), .D(n_11425), .SD(n_61462), .Q(\tab13[33] 
		));
	notech_mux2 i_17004(.S(n_55249), .A(\tab13[33] ), .B(n_55323), .Z(n_11425
		));
	notech_ao4 i_814(.A(n_1100), .B(n_13483), .C(n_1098), .D(n_13638), .Z(n_1191
		));
	notech_reg hit_adr13_reg(.CP(n_62144), .D(n_11431), .CD(n_61460), .Q(hit_adr13
		));
	notech_mux2 i_17012(.S(n_945), .A(hit_add13), .B(hit_adr13), .Z(n_11431)
		);
	notech_reg_set tab14_reg_0(.CP(n_62147), .D(n_11437), .SD(n_61463), .Q(\tab14[0] 
		));
	notech_mux2 i_17020(.S(\nbus_14016[0] ), .A(\tab14[0] ), .B(n_52162), .Z
		(n_11437));
	notech_ao4 i_813(.A(n_61950), .B(n_13722), .C(n_55460), .D(n_13639), .Z(n_1193
		));
	notech_reg_set tab14_reg_1(.CP(n_62147), .D(n_11443), .SD(n_61463), .Q(\tab14[1] 
		));
	notech_mux2 i_17028(.S(\nbus_14016[0] ), .A(\tab14[1] ), .B(n_52168), .Z
		(n_11443));
	notech_reg_set tab14_reg_2(.CP(n_62147), .D(n_11449), .SD(n_61463), .Q(\tab14[2] 
		));
	notech_mux2 i_17036(.S(\nbus_14016[0] ), .A(\tab14[2] ), .B(n_52174), .Z
		(n_11449));
	notech_ao4 i_810(.A(n_1086), .B(n_13504), .C(n_1084), .D(n_13533), .Z(n_1195
		));
	notech_reg_set tab14_reg_3(.CP(n_62147), .D(n_11455), .SD(n_61463), .Q(\tab14[3] 
		));
	notech_mux2 i_17044(.S(\nbus_14016[0] ), .A(\tab14[3] ), .B(n_52180), .Z
		(n_11455));
	notech_reg tab14_reg_4(.CP(n_62146), .D(n_11461), .CD(n_61462), .Q(\tab14[4] 
		));
	notech_mux2 i_17052(.S(\nbus_14016[0] ), .A(\tab14[4] ), .B(n_946), .Z(n_11461
		));
	notech_ao4 i_808(.A(n_1092), .B(n_13583), .C(n_1090), .D(n_13554), .Z(n_1197
		));
	notech_reg_set tab14_reg_5(.CP(n_62146), .D(n_11467), .SD(n_61462), .Q(\tab14[5] 
		));
	notech_mux2 i_17060(.S(\nbus_14016[0] ), .A(\tab14[5] ), .B(n_52192), .Z
		(n_11467));
	notech_reg_set tab14_reg_6(.CP(n_62146), .D(n_11473), .SD(n_61462), .Q(\tab14[6] 
		));
	notech_mux2 i_17068(.S(\nbus_14016[0] ), .A(\tab14[6] ), .B(n_52198), .Z
		(n_11473));
	notech_and4 i_812(.A(n_1197), .B(n_1195), .C(n_772), .D(n_775), .Z(n_1199
		));
	notech_reg_set tab14_reg_7(.CP(n_62146), .D(n_11479), .SD(n_61462), .Q(\tab14[7] 
		));
	notech_mux2 i_17076(.S(\nbus_14016[0] ), .A(\tab14[7] ), .B(n_52204), .Z
		(n_11479));
	notech_ao4 i_805(.A(n_1100), .B(n_13482), .C(n_1098), .D(n_13636), .Z(n_1200
		));
	notech_reg_set tab14_reg_8(.CP(n_62146), .D(n_11485), .SD(n_61462), .Q(\tab14[8] 
		));
	notech_mux2 i_17084(.S(\nbus_14016[0] ), .A(\tab14[8] ), .B(n_52210), .Z
		(n_11485));
	notech_reg_set tab14_reg_9(.CP(n_62139), .D(n_11491), .SD(n_61455), .Q(\tab14[9] 
		));
	notech_mux2 i_17092(.S(\nbus_14016[0] ), .A(\tab14[9] ), .B(n_52216), .Z
		(n_11491));
	notech_ao4 i_804(.A(n_61950), .B(n_13721), .C(n_55460), .D(n_13637), .Z(n_1202
		));
	notech_reg_set tab14_reg_10(.CP(n_62133), .D(n_11497), .SD(n_61449), .Q(\tab14[10] 
		));
	notech_mux2 i_17100(.S(\nbus_14016[0] ), .A(\tab14[10] ), .B(n_52222), .Z
		(n_11497));
	notech_reg_set tab14_reg_11(.CP(n_62133), .D(n_11503), .SD(n_61449), .Q(\tab14[11] 
		));
	notech_mux2 i_17108(.S(\nbus_14016[0] ), .A(\tab14[11] ), .B(n_52228), .Z
		(n_11503));
	notech_ao4 i_801(.A(n_1086), .B(n_13503), .C(n_1084), .D(n_13532), .Z(n_1204
		));
	notech_reg_set tab14_reg_12(.CP(n_62134), .D(n_11509), .SD(n_61450), .Q(\tab14[12] 
		));
	notech_mux2 i_17116(.S(\nbus_14016[0] ), .A(\tab14[12] ), .B(n_52234), .Z
		(n_11509));
	notech_reg_set tab14_reg_13(.CP(n_62133), .D(n_11515), .SD(n_61449), .Q(\tab14[13] 
		));
	notech_mux2 i_17124(.S(\nbus_14016[0] ), .A(\tab14[13] ), .B(n_52240), .Z
		(n_11515));
	notech_ao4 i_799(.A(n_1092), .B(n_13582), .C(n_1090), .D(n_13553), .Z(n_1206
		));
	notech_reg_set tab14_reg_14(.CP(n_62133), .D(n_11521), .SD(n_61449), .Q(\tab14[14] 
		));
	notech_mux2 i_17132(.S(\nbus_14016[0] ), .A(\tab14[14] ), .B(n_52246), .Z
		(n_11521));
	notech_reg_set tab14_reg_15(.CP(n_62133), .D(n_11527), .SD(n_61449), .Q(\tab14[15] 
		));
	notech_mux2 i_17140(.S(\nbus_14016[0] ), .A(\tab14[15] ), .B(n_52252), .Z
		(n_11527));
	notech_and4 i_803(.A(n_1206), .B(n_1204), .C(n_761), .D(n_764), .Z(n_1208
		));
	notech_reg_set tab14_reg_16(.CP(n_62133), .D(n_11533), .SD(n_61449), .Q(\tab14[16] 
		));
	notech_mux2 i_17148(.S(\nbus_14016[0] ), .A(\tab14[16] ), .B(n_52258), .Z
		(n_11533));
	notech_ao4 i_796(.A(n_1100), .B(n_13481), .C(n_1098), .D(n_13634), .Z(n_1209
		));
	notech_reg_set tab14_reg_17(.CP(n_62133), .D(n_11539), .SD(n_61449), .Q(\tab14[17] 
		));
	notech_mux2 i_17156(.S(n_55238), .A(\tab14[17] ), .B(n_52264), .Z(n_11539
		));
	notech_reg_set tab14_reg_18(.CP(n_62133), .D(n_11545), .SD(n_61449), .Q(\tab14[18] 
		));
	notech_mux2 i_17164(.S(n_55238), .A(\tab14[18] ), .B(n_52270), .Z(n_11545
		));
	notech_ao4 i_795(.A(n_61950), .B(n_13720), .C(n_55460), .D(n_13635), .Z(n_1211
		));
	notech_reg_set tab14_reg_19(.CP(n_62134), .D(n_11551), .SD(n_61450), .Q(\tab14[19] 
		));
	notech_mux2 i_17172(.S(n_55238), .A(\tab14[19] ), .B(n_52276), .Z(n_11551
		));
	notech_reg_set tab14_reg_20(.CP(n_62134), .D(n_11557), .SD(n_61450), .Q(\tab14[20] 
		));
	notech_mux2 i_17180(.S(n_55238), .A(\tab14[20] ), .B(n_52282), .Z(n_11557
		));
	notech_ao4 i_792(.A(n_1086), .B(n_13502), .C(n_1084), .D(n_13531), .Z(n_1213
		));
	notech_reg_set tab14_reg_21(.CP(n_62134), .D(n_11563), .SD(n_61450), .Q(\tab14[21] 
		));
	notech_mux2 i_17188(.S(n_55238), .A(\tab14[21] ), .B(n_52288), .Z(n_11563
		));
	notech_reg_set tab14_reg_22(.CP(n_62134), .D(n_11569), .SD(n_61450), .Q(\tab14[22] 
		));
	notech_mux2 i_17196(.S(n_55238), .A(\tab14[22] ), .B(n_52294), .Z(n_11569
		));
	notech_ao4 i_790(.A(n_1092), .B(n_13581), .C(n_1090), .D(n_13552), .Z(n_1215
		));
	notech_reg_set tab14_reg_23(.CP(n_62134), .D(n_11575), .SD(n_61450), .Q(\tab14[23] 
		));
	notech_mux2 i_17204(.S(n_55238), .A(\tab14[23] ), .B(n_52300), .Z(n_11575
		));
	notech_reg_set tab14_reg_24(.CP(n_62134), .D(n_11581), .SD(n_61450), .Q(\tab14[24] 
		));
	notech_mux2 i_17212(.S(n_55238), .A(\tab14[24] ), .B(n_52306), .Z(n_11581
		));
	notech_and4 i_794(.A(n_1215), .B(n_1213), .C(n_750), .D(n_753), .Z(n_1217
		));
	notech_reg_set tab14_reg_25(.CP(n_62134), .D(n_11587), .SD(n_61450), .Q(\tab14[25] 
		));
	notech_mux2 i_17220(.S(n_55238), .A(\tab14[25] ), .B(n_52312), .Z(n_11587
		));
	notech_ao4 i_787(.A(n_1100), .B(n_13480), .C(n_1098), .D(n_13632), .Z(n_1218
		));
	notech_reg_set tab14_reg_26(.CP(n_62134), .D(n_11593), .SD(n_61450), .Q(\tab14[26] 
		));
	notech_mux2 i_17228(.S(n_55238), .A(\tab14[26] ), .B(n_52318), .Z(n_11593
		));
	notech_reg_set tab14_reg_27(.CP(n_62134), .D(n_11599), .SD(n_61450), .Q(\tab14[27] 
		));
	notech_mux2 i_17236(.S(\nbus_14016[0] ), .A(\tab14[27] ), .B(n_52324), .Z
		(n_11599));
	notech_ao4 i_786(.A(n_61950), .B(n_13719), .C(n_55460), .D(n_13633), .Z(n_1220
		));
	notech_reg_set tab14_reg_28(.CP(n_62130), .D(n_11605), .SD(n_61446), .Q(\tab14[28] 
		));
	notech_mux2 i_17244(.S(n_55238), .A(\tab14[28] ), .B(n_52330), .Z(n_11605
		));
	notech_reg_set tab14_reg_29(.CP(n_62130), .D(n_11611), .SD(n_61446), .Q(\tab14[29] 
		));
	notech_mux2 i_17252(.S(n_55238), .A(\tab14[29] ), .B(n_52336), .Z(n_11611
		));
	notech_ao4 i_783(.A(n_1086), .B(n_13501), .C(n_1084), .D(n_13530), .Z(n_1222
		));
	notech_reg tab14_reg_30(.CP(n_62130), .D(n_11617), .CD(n_61446), .Q(\tab14[30] 
		));
	notech_mux2 i_17260(.S(n_55238), .A(\tab14[30] ), .B(n_947), .Z(n_11617)
		);
	notech_reg tab14_reg_32(.CP(n_62130), .D(n_11623), .CD(n_61446), .Q(\tab14[32] 
		));
	notech_mux2 i_17268(.S(n_55238), .A(\tab14[32] ), .B(n_948), .Z(n_11623)
		);
	notech_ao4 i_781(.A(n_1092), .B(n_13580), .C(n_1090), .D(n_13551), .Z(n_1224
		));
	notech_reg_set tab14_reg_33(.CP(n_62130), .D(n_11629), .SD(n_61446), .Q(\tab14[33] 
		));
	notech_mux2 i_17276(.S(n_55238), .A(\tab14[33] ), .B(n_55323), .Z(n_11629
		));
	notech_reg hit_adr14_reg(.CP(n_62129), .D(n_11635), .CD(n_61445), .Q(hit_adr14
		));
	notech_mux2 i_17284(.S(n_945), .A(hit_add14), .B(hit_adr14), .Z(n_11635)
		);
	notech_and4 i_785(.A(n_1224), .B(n_1222), .C(n_739), .D(n_742), .Z(n_1226
		));
	notech_reg nx_tab1_reg_0(.CP(n_62129), .D(n_11641), .CD(n_61445), .Q(\nx_tab1[0] 
		));
	notech_mux2 i_17292(.S(\nbus_14037[0] ), .A(\nx_tab1[0] ), .B(n_13516), 
		.Z(n_11641));
	notech_ao4 i_778(.A(n_1100), .B(n_13479), .C(n_1098), .D(n_13630), .Z(n_1227
		));
	notech_reg nx_tab1_reg_1(.CP(n_62129), .D(n_11647), .CD(n_61445), .Q(\nx_tab1[1] 
		));
	notech_mux2 i_17300(.S(\nbus_14037[0] ), .A(\nx_tab1[1] ), .B(n_13518), 
		.Z(n_11647));
	notech_reg_set nnx_tab1_reg_0(.CP(n_62129), .D(n_11653), .SD(n_61445), .Q
		(\nnx_tab1[0] ));
	notech_mux2 i_17308(.S(n_13524), .A(\nnx_tab1[0] ), .B(n_13520), .Z(n_11653
		));
	notech_ao4 i_777(.A(n_61950), .B(n_13718), .C(n_55460), .D(n_13631), .Z(n_1229
		));
	notech_reg nnx_tab1_reg_1(.CP(n_62133), .D(n_11659), .CD(n_61449), .Q(\nnx_tab1[1] 
		));
	notech_mux2 i_17316(.S(n_13524), .A(\nnx_tab1[1] ), .B(n_13522), .Z(n_11659
		));
	notech_reg hit_adr21_reg(.CP(n_62130), .D(n_11665), .CD(n_61446), .Q(hit_adr21
		));
	notech_mux2 i_17324(.S(n_945), .A(hit_add21), .B(hit_adr21), .Z(n_11665)
		);
	notech_ao4 i_774(.A(n_1086), .B(n_13500), .C(n_1084), .D(n_13529), .Z(n_1231
		));
	notech_reg_set tab22_reg_0(.CP(n_62133), .D(n_11671), .SD(n_61449), .Q(\tab22[0] 
		));
	notech_mux2 i_17332(.S(\nbus_14044[0] ), .A(\tab22[0] ), .B(n_52162), .Z
		(n_11671));
	notech_reg_set tab22_reg_1(.CP(n_62133), .D(n_11677), .SD(n_61449), .Q(\tab22[1] 
		));
	notech_mux2 i_17340(.S(\nbus_14044[0] ), .A(\tab22[1] ), .B(n_52168), .Z
		(n_11677));
	notech_ao4 i_772(.A(n_1092), .B(n_13579), .C(n_1090), .D(n_13550), .Z(n_1233
		));
	notech_reg_set tab22_reg_2(.CP(n_62130), .D(n_11683), .SD(n_61446), .Q(\tab22[2] 
		));
	notech_mux2 i_17348(.S(\nbus_14044[0] ), .A(\tab22[2] ), .B(n_52174), .Z
		(n_11683));
	notech_reg_set tab22_reg_3(.CP(n_62130), .D(n_11689), .SD(n_61446), .Q(\tab22[3] 
		));
	notech_mux2 i_17356(.S(\nbus_14044[0] ), .A(\tab22[3] ), .B(n_52180), .Z
		(n_11689));
	notech_and4 i_776(.A(n_1233), .B(n_1231), .C(n_728), .D(n_731), .Z(n_1235
		));
	notech_reg tab22_reg_4(.CP(n_62130), .D(n_11695), .CD(n_61446), .Q(\tab22[4] 
		));
	notech_mux2 i_17364(.S(\nbus_14044[0] ), .A(\tab22[4] ), .B(n_946), .Z(n_11695
		));
	notech_ao4 i_769(.A(n_1100), .B(n_13478), .C(n_1098), .D(n_13628), .Z(n_1236
		));
	notech_reg_set tab22_reg_5(.CP(n_62130), .D(n_11701), .SD(n_61446), .Q(\tab22[5] 
		));
	notech_mux2 i_17372(.S(\nbus_14044[0] ), .A(\tab22[5] ), .B(n_52192), .Z
		(n_11701));
	notech_reg_set tab22_reg_6(.CP(n_62130), .D(n_11707), .SD(n_61446), .Q(\tab22[6] 
		));
	notech_mux2 i_17380(.S(\nbus_14044[0] ), .A(\tab22[6] ), .B(n_52198), .Z
		(n_11707));
	notech_ao4 i_768(.A(n_61950), .B(n_13717), .C(n_55460), .D(n_13629), .Z(n_1238
		));
	notech_reg_set tab22_reg_7(.CP(n_62134), .D(n_11713), .SD(n_61450), .Q(\tab22[7] 
		));
	notech_mux2 i_17388(.S(\nbus_14044[0] ), .A(\tab22[7] ), .B(n_52204), .Z
		(n_11713));
	notech_reg_set tab22_reg_8(.CP(n_62138), .D(n_11719), .SD(n_61454), .Q(\tab22[8] 
		));
	notech_mux2 i_17396(.S(\nbus_14044[0] ), .A(\tab22[8] ), .B(n_52210), .Z
		(n_11719));
	notech_ao4 i_765(.A(n_1086), .B(n_13499), .C(n_1084), .D(n_13528), .Z(n_1240
		));
	notech_reg_set tab22_reg_9(.CP(n_62138), .D(n_11725), .SD(n_61454), .Q(\tab22[9] 
		));
	notech_mux2 i_17404(.S(\nbus_14044[0] ), .A(\tab22[9] ), .B(n_52216), .Z
		(n_11725));
	notech_reg_set tab22_reg_10(.CP(n_62138), .D(n_11731), .SD(n_61454), .Q(\tab22[10] 
		));
	notech_mux2 i_17412(.S(\nbus_14044[0] ), .A(\tab22[10] ), .B(n_52222), .Z
		(n_11731));
	notech_ao4 i_763(.A(n_1092), .B(n_13578), .C(n_1090), .D(n_13549), .Z(n_1242
		));
	notech_reg_set tab22_reg_11(.CP(n_62138), .D(n_11737), .SD(n_61454), .Q(\tab22[11] 
		));
	notech_mux2 i_17420(.S(\nbus_14044[0] ), .A(\tab22[11] ), .B(n_52228), .Z
		(n_11737));
	notech_reg_set tab22_reg_12(.CP(n_62138), .D(n_11743), .SD(n_61454), .Q(\tab22[12] 
		));
	notech_mux2 i_17428(.S(\nbus_14044[0] ), .A(\tab22[12] ), .B(n_52234), .Z
		(n_11743));
	notech_and4 i_767(.A(n_1242), .B(n_1240), .C(n_717), .D(n_720), .Z(n_1244
		));
	notech_reg_set tab22_reg_13(.CP(n_62137), .D(n_11749), .SD(n_61453), .Q(\tab22[13] 
		));
	notech_mux2 i_17436(.S(\nbus_14044[0] ), .A(\tab22[13] ), .B(n_52240), .Z
		(n_11749));
	notech_ao4 i_760(.A(n_1100), .B(n_13477), .C(n_54261), .D(n_13626), .Z(n_1245
		));
	notech_reg_set tab22_reg_14(.CP(n_62137), .D(n_11755), .SD(n_61453), .Q(\tab22[14] 
		));
	notech_mux2 i_17444(.S(\nbus_14044[0] ), .A(\tab22[14] ), .B(n_52246), .Z
		(n_11755));
	notech_reg_set tab22_reg_15(.CP(n_62137), .D(n_11761), .SD(n_61453), .Q(\tab22[15] 
		));
	notech_mux2 i_17452(.S(\nbus_14044[0] ), .A(\tab22[15] ), .B(n_52252), .Z
		(n_11761));
	notech_ao4 i_759(.A(n_61950), .B(n_13716), .C(n_1016), .D(n_13627), .Z(n_1247
		));
	notech_reg_set tab22_reg_16(.CP(n_62137), .D(n_11767), .SD(n_61453), .Q(\tab22[16] 
		));
	notech_mux2 i_17460(.S(\nbus_14044[0] ), .A(\tab22[16] ), .B(n_52258), .Z
		(n_11767));
	notech_reg_set tab22_reg_17(.CP(n_62139), .D(n_11773), .SD(n_61455), .Q(\tab22[17] 
		));
	notech_mux2 i_17468(.S(n_55329), .A(\tab22[17] ), .B(n_52264), .Z(n_11773
		));
	notech_ao4 i_756(.A(n_1086), .B(n_13498), .C(n_1084), .D(n_13527), .Z(n_1249
		));
	notech_reg_set tab22_reg_18(.CP(n_62138), .D(n_11779), .SD(n_61454), .Q(\tab22[18] 
		));
	notech_mux2 i_17476(.S(n_55329), .A(\tab22[18] ), .B(n_52270), .Z(n_11779
		));
	notech_reg_set tab22_reg_19(.CP(n_62139), .D(n_11785), .SD(n_61455), .Q(\tab22[19] 
		));
	notech_mux2 i_17484(.S(n_55329), .A(\tab22[19] ), .B(n_52276), .Z(n_11785
		));
	notech_ao4 i_754(.A(n_1092), .B(n_13577), .C(n_1090), .D(n_13548), .Z(n_1251
		));
	notech_reg_set tab22_reg_20(.CP(n_62139), .D(n_11791), .SD(n_61455), .Q(\tab22[20] 
		));
	notech_mux2 i_17492(.S(n_55329), .A(\tab22[20] ), .B(n_52282), .Z(n_11791
		));
	notech_reg_set tab22_reg_21(.CP(n_62138), .D(n_11797), .SD(n_61454), .Q(\tab22[21] 
		));
	notech_mux2 i_17500(.S(n_55329), .A(\tab22[21] ), .B(n_52288), .Z(n_11797
		));
	notech_and4 i_758(.A(n_1251), .B(n_1249), .C(n_706), .D(n_709), .Z(n_1253
		));
	notech_reg_set tab22_reg_22(.CP(n_62138), .D(n_11803), .SD(n_61454), .Q(\tab22[22] 
		));
	notech_mux2 i_17508(.S(n_55329), .A(\tab22[22] ), .B(n_52294), .Z(n_11803
		));
	notech_ao4 i_751(.A(n_1100), .B(n_13476), .C(n_54261), .D(n_13624), .Z(n_1254
		));
	notech_reg_set tab22_reg_23(.CP(n_62138), .D(n_11809), .SD(n_61454), .Q(\tab22[23] 
		));
	notech_mux2 i_17516(.S(n_55329), .A(\tab22[23] ), .B(n_52300), .Z(n_11809
		));
	notech_reg_set tab22_reg_24(.CP(n_62138), .D(n_11815), .SD(n_61454), .Q(\tab22[24] 
		));
	notech_mux2 i_17524(.S(n_55329), .A(\tab22[24] ), .B(n_52306), .Z(n_11815
		));
	notech_ao4 i_750(.A(n_61946), .B(n_13715), .C(n_55460), .D(n_13625), .Z(n_1256
		));
	notech_reg_set tab22_reg_25(.CP(n_62138), .D(n_11821), .SD(n_61454), .Q(\tab22[25] 
		));
	notech_mux2 i_17532(.S(n_55329), .A(\tab22[25] ), .B(n_52312), .Z(n_11821
		));
	notech_reg_set tab22_reg_26(.CP(n_62135), .D(n_11827), .SD(n_61451), .Q(\tab22[26] 
		));
	notech_mux2 i_17540(.S(n_55329), .A(\tab22[26] ), .B(n_52318), .Z(n_11827
		));
	notech_ao4 i_747(.A(n_1086), .B(n_13497), .C(n_1084), .D(n_13526), .Z(n_1258
		));
	notech_reg_set tab22_reg_27(.CP(n_62135), .D(n_11833), .SD(n_61451), .Q(\tab22[27] 
		));
	notech_mux2 i_17548(.S(\nbus_14044[0] ), .A(\tab22[27] ), .B(n_52324), .Z
		(n_11833));
	notech_reg_set tab22_reg_28(.CP(n_62135), .D(n_11839), .SD(n_61451), .Q(\tab22[28] 
		));
	notech_mux2 i_17556(.S(n_55329), .A(\tab22[28] ), .B(n_52330), .Z(n_11839
		));
	notech_ao4 i_745(.A(n_1092), .B(n_13576), .C(n_1090), .D(n_13547), .Z(n_1260
		));
	notech_reg_set tab22_reg_29(.CP(n_62135), .D(n_11845), .SD(n_61451), .Q(\tab22[29] 
		));
	notech_mux2 i_17564(.S(n_55329), .A(\tab22[29] ), .B(n_52336), .Z(n_11845
		));
	notech_reg tab22_reg_30(.CP(n_62135), .D(n_11851), .CD(n_61451), .Q(\tab22[30] 
		));
	notech_mux2 i_17572(.S(n_55329), .A(\tab22[30] ), .B(n_947), .Z(n_11851)
		);
	notech_and4 i_749(.A(n_1260), .B(n_1258), .C(n_695), .D(n_698), .Z(n_1262
		));
	notech_reg tab22_reg_32(.CP(n_62135), .D(n_11857), .CD(n_61451), .Q(\tab22[32] 
		));
	notech_mux2 i_17580(.S(n_55329), .A(\tab22[32] ), .B(n_948), .Z(n_11857)
		);
	notech_ao4 i_742(.A(n_1100), .B(n_13475), .C(n_54261), .D(n_13622), .Z(n_1263
		));
	notech_reg_set tab22_reg_33(.CP(n_62135), .D(n_11863), .SD(n_61451), .Q(\tab22[33] 
		));
	notech_mux2 i_17588(.S(n_55329), .A(\tab22[33] ), .B(n_55323), .Z(n_11863
		));
	notech_reg hit_adr22_reg(.CP(n_62135), .D(n_11869), .CD(n_61451), .Q(hit_adr22
		));
	notech_mux2 i_17596(.S(n_945), .A(hit_add22), .B(hit_adr22), .Z(n_11869)
		);
	notech_ao4 i_741(.A(n_61946), .B(n_13714), .C(n_55460), .D(n_13623), .Z(n_1265
		));
	notech_reg_set tab24_reg_0(.CP(n_62135), .D(n_11875), .SD(n_61451), .Q(\tab24[0] 
		));
	notech_mux2 i_17604(.S(\nbus_14017[0] ), .A(\tab24[0] ), .B(n_52162), .Z
		(n_11875));
	notech_reg_set tab24_reg_1(.CP(n_62137), .D(n_11881), .SD(n_61453), .Q(\tab24[1] 
		));
	notech_mux2 i_17612(.S(\nbus_14017[0] ), .A(\tab24[1] ), .B(n_52168), .Z
		(n_11881));
	notech_ao4 i_738(.A(n_1086), .B(n_13496), .C(n_1084), .D(n_13525), .Z(n_1267
		));
	notech_reg_set tab24_reg_2(.CP(n_62137), .D(n_11887), .SD(n_61453), .Q(\tab24[2] 
		));
	notech_mux2 i_17620(.S(\nbus_14017[0] ), .A(\tab24[2] ), .B(n_52174), .Z
		(n_11887));
	notech_reg_set tab24_reg_3(.CP(n_62137), .D(n_11893), .SD(n_61453), .Q(\tab24[3] 
		));
	notech_mux2 i_17628(.S(\nbus_14017[0] ), .A(\tab24[3] ), .B(n_52180), .Z
		(n_11893));
	notech_ao4 i_736(.A(n_1092), .B(n_13575), .C(n_1090), .D(n_13546), .Z(n_1269
		));
	notech_reg tab24_reg_4(.CP(n_62137), .D(n_11899), .CD(n_61453), .Q(\tab24[4] 
		));
	notech_mux2 i_17636(.S(\nbus_14017[0] ), .A(\tab24[4] ), .B(n_946), .Z(n_11899
		));
	notech_reg_set tab24_reg_5(.CP(n_62137), .D(n_11905), .SD(n_61453), .Q(\tab24[5] 
		));
	notech_mux2 i_17644(.S(\nbus_14017[0] ), .A(\tab24[5] ), .B(n_52192), .Z
		(n_11905));
	notech_and4 i_740(.A(n_1269), .B(n_1267), .C(n_687), .D(n_684), .Z(n_1271
		));
	notech_reg_set tab24_reg_6(.CP(n_62135), .D(n_11911), .SD(n_61451), .Q(\tab24[6] 
		));
	notech_mux2 i_17652(.S(\nbus_14017[0] ), .A(\tab24[6] ), .B(n_52198), .Z
		(n_11911));
	notech_ao4 i_733(.A(n_1100), .B(n_13474), .C(n_54261), .D(n_13620), .Z(n_1272
		));
	notech_reg_set tab24_reg_7(.CP(n_62135), .D(n_11917), .SD(n_61451), .Q(\tab24[7] 
		));
	notech_mux2 i_17660(.S(\nbus_14017[0] ), .A(\tab24[7] ), .B(n_52204), .Z
		(n_11917));
	notech_reg_set tab24_reg_8(.CP(n_62137), .D(n_11923), .SD(n_61453), .Q(\tab24[8] 
		));
	notech_mux2 i_17668(.S(\nbus_14017[0] ), .A(\tab24[8] ), .B(n_52210), .Z
		(n_11923));
	notech_ao4 i_732(.A(n_61950), .B(n_13713), .C(n_55460), .D(n_13621), .Z(n_1274
		));
	notech_reg_set tab24_reg_9(.CP(n_62137), .D(n_11929), .SD(n_61453), .Q(\tab24[9] 
		));
	notech_mux2 i_17676(.S(\nbus_14017[0] ), .A(\tab24[9] ), .B(n_52216), .Z
		(n_11929));
	notech_reg_set tab24_reg_10(.CP(n_62109), .D(n_11935), .SD(n_61425), .Q(\tab24[10] 
		));
	notech_mux2 i_17684(.S(\nbus_14017[0] ), .A(\tab24[10] ), .B(n_52222), .Z
		(n_11935));
	notech_ao4 i_731(.A(n_54261), .B(n_13619), .C(n_420), .D(n_13712), .Z(n_1276
		));
	notech_reg_set tab24_reg_11(.CP(n_62081), .D(n_11941), .SD(n_61397), .Q(\tab24[11] 
		));
	notech_mux2 i_17692(.S(\nbus_14017[0] ), .A(\tab24[11] ), .B(n_52228), .Z
		(n_11941));
	notech_ao4 i_730(.A(n_54261), .B(n_13618), .C(n_420), .D(n_13711), .Z(n_1277
		));
	notech_reg_set tab24_reg_12(.CP(n_62081), .D(n_11947), .SD(n_61397), .Q(\tab24[12] 
		));
	notech_mux2 i_17700(.S(\nbus_14017[0] ), .A(\tab24[12] ), .B(n_52234), .Z
		(n_11947));
	notech_ao4 i_729(.A(n_54261), .B(n_13616), .C(n_420), .D(n_13710), .Z(n_1278
		));
	notech_reg_set tab24_reg_13(.CP(n_62081), .D(n_11953), .SD(n_61397), .Q(\tab24[13] 
		));
	notech_mux2 i_17708(.S(\nbus_14017[0] ), .A(\tab24[13] ), .B(n_52240), .Z
		(n_11953));
	notech_ao4 i_728(.A(n_54261), .B(n_13615), .C(n_420), .D(n_13709), .Z(n_1279
		));
	notech_reg_set tab24_reg_14(.CP(n_62081), .D(n_11959), .SD(n_61397), .Q(\tab24[14] 
		));
	notech_mux2 i_17716(.S(\nbus_14017[0] ), .A(\tab24[14] ), .B(n_52246), .Z
		(n_11959));
	notech_ao4 i_727(.A(n_54261), .B(n_13614), .C(n_420), .D(n_13708), .Z(n_1280
		));
	notech_reg_set tab24_reg_15(.CP(n_62081), .D(n_11965), .SD(n_61397), .Q(\tab24[15] 
		));
	notech_mux2 i_17724(.S(\nbus_14017[0] ), .A(\tab24[15] ), .B(n_52252), .Z
		(n_11965));
	notech_ao4 i_726(.A(n_54261), .B(n_13613), .C(n_420), .D(n_13707), .Z(n_1281
		));
	notech_reg_set tab24_reg_16(.CP(n_62079), .D(n_11971), .SD(n_61395), .Q(\tab24[16] 
		));
	notech_mux2 i_17732(.S(\nbus_14017[0] ), .A(\tab24[16] ), .B(n_52258), .Z
		(n_11971));
	notech_ao4 i_725(.A(n_1098), .B(n_13612), .C(n_420), .D(n_13706), .Z(n_1282
		));
	notech_reg_set tab24_reg_17(.CP(n_62079), .D(n_11977), .SD(n_61395), .Q(\tab24[17] 
		));
	notech_mux2 i_17740(.S(n_55309), .A(\tab24[17] ), .B(n_52264), .Z(n_11977
		));
	notech_ao4 i_724(.A(n_54261), .B(n_13611), .C(n_420), .D(n_13705), .Z(n_1283
		));
	notech_reg_set tab24_reg_18(.CP(n_62081), .D(n_11983), .SD(n_61397), .Q(\tab24[18] 
		));
	notech_mux2 i_17748(.S(n_55309), .A(\tab24[18] ), .B(n_52270), .Z(n_11983
		));
	notech_ao4 i_723(.A(n_54261), .B(n_13610), .C(n_420), .D(n_13704), .Z(n_1284
		));
	notech_reg_set tab24_reg_19(.CP(n_62081), .D(n_11989), .SD(n_61397), .Q(\tab24[19] 
		));
	notech_mux2 i_17756(.S(n_55309), .A(\tab24[19] ), .B(n_52276), .Z(n_11989
		));
	notech_ao4 i_722(.A(n_54261), .B(n_13609), .C(n_420), .D(n_13703), .Z(n_1285
		));
	notech_reg_set tab24_reg_20(.CP(n_62082), .D(n_11995), .SD(n_61398), .Q(\tab24[20] 
		));
	notech_mux2 i_17764(.S(n_55309), .A(\tab24[20] ), .B(n_52282), .Z(n_11995
		));
	notech_ao4 i_721(.A(n_54261), .B(n_13608), .C(n_420), .D(n_13702), .Z(n_1286
		));
	notech_reg_set tab24_reg_21(.CP(n_62082), .D(n_12001), .SD(n_61398), .Q(\tab24[21] 
		));
	notech_mux2 i_17772(.S(n_55309), .A(\tab24[21] ), .B(n_52288), .Z(n_12001
		));
	notech_ao4 i_720(.A(n_54261), .B(n_13607), .C(n_420), .D(n_13701), .Z(n_1287
		));
	notech_reg_set tab24_reg_22(.CP(n_62082), .D(n_12007), .SD(n_61398), .Q(\tab24[22] 
		));
	notech_mux2 i_17780(.S(n_55309), .A(\tab24[22] ), .B(n_52294), .Z(n_12007
		));
	notech_ao4 i_75908(.A(n_61950), .B(n_13761), .C(n_984), .D(n_985), .Z(oread_ack100169
		));
	notech_reg_set tab24_reg_23(.CP(n_62082), .D(n_12013), .SD(n_61398), .Q(\tab24[23] 
		));
	notech_mux2 i_17788(.S(n_55309), .A(\tab24[23] ), .B(n_52300), .Z(n_12013
		));
	notech_ao4 i_77497(.A(n_951), .B(n_13760), .C(n_992), .D(n_993), .Z(\nbus_14018[0] 
		));
	notech_reg_set tab24_reg_24(.CP(n_62082), .D(n_12019), .SD(n_61398), .Q(\tab24[24] 
		));
	notech_mux2 i_17796(.S(n_55309), .A(\tab24[24] ), .B(n_52306), .Z(n_12019
		));
	notech_or4 i_78139(.A(n_488), .B(\nbus_14038[0] ), .C(n_1022), .D(n_13448
		), .Z(\nbus_14033[0] ));
	notech_reg_set tab24_reg_25(.CP(n_62081), .D(n_12025), .SD(n_61397), .Q(\tab24[25] 
		));
	notech_mux2 i_17804(.S(n_55309), .A(\tab24[25] ), .B(n_52312), .Z(n_12025
		));
	notech_nand3 i_78746(.A(n_613), .B(n_610), .C(n_607), .Z(\nbus_14041[0] 
		));
	notech_reg_set tab24_reg_26(.CP(n_62081), .D(n_12031), .SD(n_61397), .Q(\tab24[26] 
		));
	notech_mux2 i_17812(.S(n_55309), .A(\tab24[26] ), .B(n_52318), .Z(n_12031
		));
	notech_nao3 i_77955(.A(n_610), .B(n_607), .C(n_608), .Z(\nbus_14029[0] )
		);
	notech_reg_set tab24_reg_27(.CP(n_62081), .D(n_12037), .SD(n_61397), .Q(\tab24[27] 
		));
	notech_mux2 i_17820(.S(\nbus_14017[0] ), .A(\tab24[27] ), .B(n_52324), .Z
		(n_12037));
	notech_nao3 i_78395(.A(n_610), .B(n_588), .C(n_608), .Z(\nbus_14036[0] )
		);
	notech_reg_set tab24_reg_28(.CP(n_62081), .D(n_12043), .SD(n_61397), .Q(\tab24[28] 
		));
	notech_mux2 i_17828(.S(n_55309), .A(\tab24[28] ), .B(n_52330), .Z(n_12043
		));
	notech_nand3 i_78283(.A(n_613), .B(n_610), .C(n_585), .Z(\nbus_14035[0] 
		));
	notech_reg_set tab24_reg_29(.CP(n_62078), .D(n_12049), .SD(n_61394), .Q(\tab24[29] 
		));
	notech_mux2 i_17836(.S(n_55309), .A(\tab24[29] ), .B(n_52336), .Z(n_12049
		));
	notech_nand3 i_76910(.A(n_613), .B(n_610), .C(n_584), .Z(\nbus_14014[0] 
		));
	notech_reg tab24_reg_30(.CP(n_62078), .D(n_12055), .CD(n_61394), .Q(\tab24[30] 
		));
	notech_mux2 i_17844(.S(n_55309), .A(\tab24[30] ), .B(n_947), .Z(n_12055)
		);
	notech_nand3 i_77183(.A(n_613), .B(n_610), .C(n_583), .Z(\nbus_14016[0] 
		));
	notech_reg tab24_reg_32(.CP(n_62078), .D(n_12061), .CD(n_61394), .Q(\tab24[32] 
		));
	notech_mux2 i_17852(.S(n_55309), .A(\tab24[32] ), .B(n_948), .Z(n_12061)
		);
	notech_nand2 i_78505(.A(n_1023), .B(n_1038), .Z(\nbus_14037[0] ));
	notech_reg_set tab24_reg_33(.CP(n_62078), .D(n_12067), .SD(n_61394), .Q(\tab24[33] 
		));
	notech_mux2 i_17860(.S(n_55309), .A(\tab24[33] ), .B(n_55323), .Z(n_12067
		));
	notech_ao4 i_78107(.A(n_1030), .B(n_1037), .C(n_1023), .D(n_13472), .Z(\nbus_14032[0] 
		));
	notech_reg hit_adr24_reg(.CP(n_62078), .D(n_12073), .CD(n_61394), .Q(hit_adr24
		));
	notech_mux2 i_17868(.S(n_945), .A(hit_add24), .B(hit_adr24), .Z(n_12073)
		);
	notech_nao3 i_78858(.A(n_610), .B(n_563), .C(n_608), .Z(\nbus_14044[0] )
		);
	notech_reg_set nnx_tab2_reg_0(.CP(n_62078), .D(n_12079), .SD(n_61394), .Q
		(\nnx_tab2[0] ));
	notech_mux2 i_17876(.S(n_13570), .A(\nnx_tab2[0] ), .B(n_13566), .Z(n_12079
		));
	notech_nao3 i_77295(.A(n_610), .B(n_562), .C(n_608), .Z(\nbus_14017[0] )
		);
	notech_reg nnx_tab2_reg_1(.CP(n_62078), .D(n_12085), .CD(n_61394), .Q(\nnx_tab2[1] 
		));
	notech_mux2 i_17884(.S(n_13570), .A(\nnx_tab2[1] ), .B(n_13568), .Z(n_12085
		));
	notech_ao4 i_78083(.A(n_1031), .B(n_1030), .C(n_1023), .D(n_13471), .Z(\nbus_14031[0] 
		));
	notech_reg nx_tab2_reg_0(.CP(n_62078), .D(n_12091), .CD(n_61394), .Q(\nx_tab2[0] 
		));
	notech_mux2 i_17892(.S(\nbus_14040[0] ), .A(\nx_tab2[0] ), .B(n_13571), 
		.Z(n_12091));
	notech_nand2 i_78723(.A(n_1023), .B(n_1032), .Z(\nbus_14040[0] ));
	notech_reg nx_tab2_reg_1(.CP(n_62078), .D(n_12097), .CD(n_61394), .Q(\nx_tab2[1] 
		));
	notech_mux2 i_17900(.S(\nbus_14040[0] ), .A(\nx_tab2[1] ), .B(n_13573), 
		.Z(n_12097));
	notech_nand3 i_78171(.A(n_613), .B(n_610), .C(n_542), .Z(\nbus_14034[0] 
		));
	notech_reg_set tab11_reg_0(.CP(n_62079), .D(n_12103), .SD(n_61395), .Q(\tab11[0] 
		));
	notech_mux2 i_17908(.S(\nbus_14034[0] ), .A(\tab11[0] ), .B(n_52162), .Z
		(n_12103));
	notech_nao3 i_77774(.A(n_610), .B(n_541), .C(n_608), .Z(\nbus_14028[0] )
		);
	notech_reg_set tab11_reg_1(.CP(n_62079), .D(n_12109), .SD(n_61395), .Q(\tab11[1] 
		));
	notech_mux2 i_17916(.S(\nbus_14034[0] ), .A(\tab11[1] ), .B(n_52168), .Z
		(n_12109));
	notech_or2 i_116(.A(n_488), .B(n_13448), .Z(n_52374));
	notech_reg_set tab11_reg_2(.CP(n_62079), .D(n_12115), .SD(n_61395), .Q(\tab11[2] 
		));
	notech_mux2 i_17924(.S(\nbus_14034[0] ), .A(\tab11[2] ), .B(n_52174), .Z
		(n_12115));
	notech_nand2 i_118(.A(n_1023), .B(n_636), .Z(\nbus_14038[0] ));
	notech_reg_set tab11_reg_3(.CP(n_62079), .D(n_12121), .SD(n_61395), .Q(\tab11[3] 
		));
	notech_mux2 i_17932(.S(\nbus_14034[0] ), .A(\tab11[3] ), .B(n_52180), .Z
		(n_12121));
	notech_reg tab11_reg_4(.CP(n_62079), .D(n_12127), .CD(n_61395), .Q(\tab11[4] 
		));
	notech_mux2 i_17940(.S(\nbus_14034[0] ), .A(\tab11[4] ), .B(n_946), .Z(n_12127
		));
	notech_or2 i_77919(.A(n_488), .B(n_489), .Z(n_53974));
	notech_reg_set tab11_reg_5(.CP(n_62079), .D(n_12133), .SD(n_61395), .Q(\tab11[5] 
		));
	notech_mux2 i_17948(.S(\nbus_14034[0] ), .A(\tab11[5] ), .B(n_52192), .Z
		(n_12133));
	notech_ao4 i_117(.A(n_1030), .B(n_641), .C(data_miss[5]), .D(n_950), .Z(\nbus_14013[0] 
		));
	notech_reg_set tab11_reg_6(.CP(n_62079), .D(n_12139), .SD(n_61395), .Q(\tab11[6] 
		));
	notech_mux2 i_17956(.S(\nbus_14034[0] ), .A(\tab11[6] ), .B(n_52198), .Z
		(n_12139));
	notech_ao4 i_99(.A(data_miss[0]), .B(n_996), .C(n_1004), .D(n_13439), .Z
		(n_52377));
	notech_reg_set tab11_reg_7(.CP(n_62079), .D(n_12145), .SD(n_61395), .Q(\tab11[7] 
		));
	notech_mux2 i_17964(.S(\nbus_14034[0] ), .A(\tab11[7] ), .B(n_52204), .Z
		(n_12145));
	notech_mux2 i_122740(.S(n_951), .A(iDaddr[12]), .B(iDaddr_f[12]), .Z(\addr_miss_0[2] 
		));
	notech_reg_set tab11_reg_8(.CP(n_62079), .D(n_12151), .SD(n_61395), .Q(\tab11[8] 
		));
	notech_mux2 i_17972(.S(\nbus_14034[0] ), .A(\tab11[8] ), .B(n_52210), .Z
		(n_12151));
	notech_mux2 i_222741(.S(n_951), .A(iDaddr[13]), .B(iDaddr_f[13]), .Z(\addr_miss_0[3] 
		));
	notech_reg_set tab11_reg_9(.CP(n_62082), .D(n_12157), .SD(n_61398), .Q(\tab11[9] 
		));
	notech_mux2 i_17980(.S(\nbus_14034[0] ), .A(\tab11[9] ), .B(n_52216), .Z
		(n_12157));
	notech_mux2 i_322742(.S(n_951), .A(iDaddr[14]), .B(iDaddr_f[14]), .Z(\addr_miss_0[4] 
		));
	notech_reg_set tab11_reg_10(.CP(n_62086), .D(n_12163), .SD(n_61402), .Q(\tab11[10] 
		));
	notech_mux2 i_17988(.S(\nbus_14034[0] ), .A(\tab11[10] ), .B(n_52222), .Z
		(n_12163));
	notech_mux2 i_422743(.S(n_951), .A(iDaddr[15]), .B(iDaddr_f[15]), .Z(\addr_miss_0[5] 
		));
	notech_reg_set tab11_reg_11(.CP(n_62086), .D(n_12169), .SD(n_61402), .Q(\tab11[11] 
		));
	notech_mux2 i_17996(.S(\nbus_14034[0] ), .A(\tab11[11] ), .B(n_52228), .Z
		(n_12169));
	notech_mux2 i_522744(.S(n_951), .A(iDaddr[16]), .B(iDaddr_f[16]), .Z(\addr_miss_0[6] 
		));
	notech_reg_set tab11_reg_12(.CP(n_62086), .D(n_12175), .SD(n_61402), .Q(\tab11[12] 
		));
	notech_mux2 i_18004(.S(\nbus_14034[0] ), .A(\tab11[12] ), .B(n_52234), .Z
		(n_12175));
	notech_mux2 i_622745(.S(n_59313), .A(iDaddr[17]), .B(iDaddr_f[17]), .Z(\addr_miss_0[7] 
		));
	notech_reg_set tab11_reg_13(.CP(n_62086), .D(n_12181), .SD(n_61402), .Q(\tab11[13] 
		));
	notech_mux2 i_18012(.S(\nbus_14034[0] ), .A(\tab11[13] ), .B(n_52240), .Z
		(n_12181));
	notech_mux2 i_722746(.S(n_59313), .A(iDaddr[18]), .B(iDaddr_f[18]), .Z(\addr_miss_0[8] 
		));
	notech_reg_set tab11_reg_14(.CP(n_62086), .D(n_12187), .SD(n_61402), .Q(\tab11[14] 
		));
	notech_mux2 i_18020(.S(\nbus_14034[0] ), .A(\tab11[14] ), .B(n_52246), .Z
		(n_12187));
	notech_mux2 i_822747(.S(n_59313), .A(iDaddr[19]), .B(iDaddr_f[19]), .Z(\addr_miss_0[9] 
		));
	notech_reg_set tab11_reg_15(.CP(n_62086), .D(n_12193), .SD(n_61402), .Q(\tab11[15] 
		));
	notech_mux2 i_18028(.S(\nbus_14034[0] ), .A(\tab11[15] ), .B(n_52252), .Z
		(n_12193));
	notech_mux2 i_922748(.S(n_59313), .A(iDaddr[20]), .B(iDaddr_f[20]), .Z(\addr_miss_0[10] 
		));
	notech_reg_set tab11_reg_16(.CP(n_62086), .D(n_12199), .SD(n_61402), .Q(\tab11[16] 
		));
	notech_mux2 i_18036(.S(\nbus_14034[0] ), .A(\tab11[16] ), .B(n_52258), .Z
		(n_12199));
	notech_mux2 i_1022749(.S(n_59313), .A(iDaddr[21]), .B(iDaddr_f[21]), .Z(\addr_miss_0[11] 
		));
	notech_reg_set tab11_reg_17(.CP(n_62086), .D(n_12205), .SD(n_61402), .Q(\tab11[17] 
		));
	notech_mux2 i_18044(.S(n_55260), .A(\tab11[17] ), .B(n_52264), .Z(n_12205
		));
	notech_mux2 i_1122750(.S(n_59313), .A(iDaddr[22]), .B(iDaddr_f[22]), .Z(n_50869
		));
	notech_reg_set tab11_reg_18(.CP(n_62086), .D(n_12211), .SD(n_61402), .Q(\tab11[18] 
		));
	notech_mux2 i_18052(.S(n_55260), .A(\tab11[18] ), .B(n_52270), .Z(n_12211
		));
	notech_mux2 i_1222751(.S(n_59313), .A(iDaddr[23]), .B(iDaddr_f[23]), .Z(n_50870
		));
	notech_reg_set tab11_reg_19(.CP(n_62087), .D(n_12217), .SD(n_61403), .Q(\tab11[19] 
		));
	notech_mux2 i_18060(.S(n_55260), .A(\tab11[19] ), .B(n_52276), .Z(n_12217
		));
	notech_mux2 i_1322752(.S(n_59313), .A(iDaddr[24]), .B(iDaddr_f[24]), .Z(n_50871
		));
	notech_reg_set tab11_reg_20(.CP(n_62087), .D(n_12223), .SD(n_61403), .Q(\tab11[20] 
		));
	notech_mux2 i_18068(.S(n_55260), .A(\tab11[20] ), .B(n_52282), .Z(n_12223
		));
	notech_mux2 i_1422753(.S(n_59313), .A(iDaddr[25]), .B(iDaddr_f[25]), .Z(n_50872
		));
	notech_reg_set tab11_reg_21(.CP(n_62087), .D(n_12229), .SD(n_61403), .Q(\tab11[21] 
		));
	notech_mux2 i_18076(.S(n_55260), .A(\tab11[21] ), .B(n_52288), .Z(n_12229
		));
	notech_mux2 i_1522754(.S(n_59313), .A(iDaddr[26]), .B(iDaddr_f[26]), .Z(n_50873
		));
	notech_reg_set tab11_reg_22(.CP(n_62087), .D(n_12235), .SD(n_61403), .Q(\tab11[22] 
		));
	notech_mux2 i_18084(.S(n_55260), .A(\tab11[22] ), .B(n_52294), .Z(n_12235
		));
	notech_mux2 i_1622755(.S(n_59313), .A(iDaddr[27]), .B(iDaddr_f[27]), .Z(n_50874
		));
	notech_reg_set tab11_reg_23(.CP(n_62087), .D(n_12241), .SD(n_61403), .Q(\tab11[23] 
		));
	notech_mux2 i_18092(.S(n_55260), .A(\tab11[23] ), .B(n_52300), .Z(n_12241
		));
	notech_mux2 i_1722756(.S(n_59313), .A(iDaddr[28]), .B(iDaddr_f[28]), .Z(n_50875
		));
	notech_reg_set tab11_reg_24(.CP(n_62087), .D(n_12247), .SD(n_61403), .Q(\tab11[24] 
		));
	notech_mux2 i_18100(.S(n_55260), .A(\tab11[24] ), .B(n_52306), .Z(n_12247
		));
	notech_mux2 i_1822757(.S(n_59313), .A(iDaddr[29]), .B(iDaddr_f[29]), .Z(n_50876
		));
	notech_reg_set tab11_reg_25(.CP(n_62087), .D(n_12253), .SD(n_61403), .Q(\tab11[25] 
		));
	notech_mux2 i_18108(.S(n_55260), .A(\tab11[25] ), .B(n_52312), .Z(n_12253
		));
	notech_mux2 i_1922758(.S(n_59313), .A(iDaddr[30]), .B(iDaddr_f[30]), .Z(n_50877
		));
	notech_reg_set tab11_reg_26(.CP(n_62087), .D(n_12259), .SD(n_61403), .Q(\tab11[26] 
		));
	notech_mux2 i_18116(.S(n_55260), .A(\tab11[26] ), .B(n_52318), .Z(n_12259
		));
	notech_mux2 i_2022759(.S(n_59313), .A(iDaddr[31]), .B(iDaddr_f[31]), .Z(n_50878
		));
	notech_reg_set tab11_reg_27(.CP(n_62087), .D(n_12265), .SD(n_61403), .Q(\tab11[27] 
		));
	notech_mux2 i_18124(.S(\nbus_14034[0] ), .A(\tab11[27] ), .B(n_52324), .Z
		(n_12265));
	notech_nand2 i_122216(.A(n_1287), .B(n_409), .Z(n_53038));
	notech_reg_set tab11_reg_28(.CP(n_62083), .D(n_12271), .SD(n_61399), .Q(\tab11[28] 
		));
	notech_mux2 i_18132(.S(n_55260), .A(\tab11[28] ), .B(n_52330), .Z(n_12271
		));
	notech_nand2 i_222217(.A(n_1286), .B(n_410), .Z(n_53045));
	notech_reg_set tab11_reg_29(.CP(n_62083), .D(n_12277), .SD(n_61399), .Q(\tab11[29] 
		));
	notech_mux2 i_18140(.S(n_55260), .A(\tab11[29] ), .B(n_52336), .Z(n_12277
		));
	notech_nand2 i_322218(.A(n_1285), .B(n_411), .Z(n_53052));
	notech_reg tab11_reg_30(.CP(n_62083), .D(n_12283), .CD(n_61399), .Q(\tab11[30] 
		));
	notech_mux2 i_18148(.S(n_55260), .A(\tab11[30] ), .B(n_947), .Z(n_12283)
		);
	notech_nand2 i_422219(.A(n_1284), .B(n_412), .Z(n_53059));
	notech_reg tab11_reg_32(.CP(n_62083), .D(n_12289), .CD(n_61399), .Q(\tab11[32] 
		));
	notech_mux2 i_18156(.S(n_55260), .A(\tab11[32] ), .B(n_948), .Z(n_12289)
		);
	notech_nand2 i_522220(.A(n_1283), .B(n_413), .Z(n_53066));
	notech_reg_set tab11_reg_33(.CP(n_62082), .D(n_12295), .SD(n_61398), .Q(\tab11[33] 
		));
	notech_mux2 i_18164(.S(n_55260), .A(\tab11[33] ), .B(n_55323), .Z(n_12295
		));
	notech_nand2 i_622221(.A(n_1282), .B(n_414), .Z(n_53073));
	notech_reg_set tab23_reg_0(.CP(n_62082), .D(n_12301), .SD(n_61398), .Q(\tab23[0] 
		));
	notech_mux2 i_18172(.S(\nbus_14028[0] ), .A(\tab23[0] ), .B(n_52162), .Z
		(n_12301));
	notech_nand2 i_722222(.A(n_1281), .B(n_415), .Z(n_53080));
	notech_reg_set tab23_reg_1(.CP(n_62082), .D(n_12307), .SD(n_61398), .Q(\tab23[1] 
		));
	notech_mux2 i_18180(.S(\nbus_14028[0] ), .A(\tab23[1] ), .B(n_52168), .Z
		(n_12307));
	notech_nand2 i_822223(.A(n_1280), .B(n_416), .Z(n_53087));
	notech_reg_set tab23_reg_2(.CP(n_62082), .D(n_12313), .SD(n_61398), .Q(\tab23[2] 
		));
	notech_mux2 i_18188(.S(\nbus_14028[0] ), .A(\tab23[2] ), .B(n_52174), .Z
		(n_12313));
	notech_nand2 i_922224(.A(n_1279), .B(n_417), .Z(n_53094));
	notech_reg_set tab23_reg_3(.CP(n_62082), .D(n_12319), .SD(n_61398), .Q(\tab23[3] 
		));
	notech_mux2 i_18196(.S(\nbus_14028[0] ), .A(\tab23[3] ), .B(n_52180), .Z
		(n_12319));
	notech_nand2 i_1022225(.A(n_1278), .B(n_418), .Z(n_53101));
	notech_reg tab23_reg_4(.CP(n_62083), .D(n_12325), .CD(n_61399), .Q(\tab23[4] 
		));
	notech_mux2 i_18204(.S(\nbus_14028[0] ), .A(\tab23[4] ), .B(n_946), .Z(n_12325
		));
	notech_nand2 i_1122226(.A(n_1277), .B(n_419), .Z(n_53108));
	notech_reg_set tab23_reg_5(.CP(n_62083), .D(n_12331), .SD(n_61399), .Q(\tab23[5] 
		));
	notech_mux2 i_18212(.S(\nbus_14028[0] ), .A(\tab23[5] ), .B(n_52192), .Z
		(n_12331));
	notech_nand2 i_1222227(.A(n_1276), .B(n_421), .Z(n_53115));
	notech_reg_set tab23_reg_6(.CP(n_62086), .D(n_12337), .SD(n_61402), .Q(\tab23[6] 
		));
	notech_mux2 i_18220(.S(\nbus_14028[0] ), .A(\tab23[6] ), .B(n_52198), .Z
		(n_12337));
	notech_and4 i_1322228(.A(n_1272), .B(n_1274), .C(n_1271), .D(n_681), .Z(n_53122
		));
	notech_reg_set tab23_reg_7(.CP(n_62086), .D(n_12343), .SD(n_61402), .Q(\tab23[7] 
		));
	notech_mux2 i_18228(.S(\nbus_14028[0] ), .A(\tab23[7] ), .B(n_52204), .Z
		(n_12343));
	notech_and4 i_1422229(.A(n_1263), .B(n_1265), .C(n_1262), .D(n_692), .Z(n_53129
		));
	notech_reg_set tab23_reg_8(.CP(n_62083), .D(n_12349), .SD(n_61399), .Q(\tab23[8] 
		));
	notech_mux2 i_18236(.S(\nbus_14028[0] ), .A(\tab23[8] ), .B(n_52210), .Z
		(n_12349));
	notech_and4 i_1522230(.A(n_1254), .B(n_1256), .C(n_1253), .D(n_703), .Z(n_53136
		));
	notech_reg_set tab23_reg_9(.CP(n_62083), .D(n_12355), .SD(n_61399), .Q(\tab23[9] 
		));
	notech_mux2 i_18244(.S(\nbus_14028[0] ), .A(\tab23[9] ), .B(n_52216), .Z
		(n_12355));
	notech_and4 i_1622231(.A(n_1245), .B(n_1247), .C(n_1244), .D(n_714), .Z(n_53143
		));
	notech_reg_set tab23_reg_10(.CP(n_62083), .D(n_12361), .SD(n_61399), .Q(\tab23[10] 
		));
	notech_mux2 i_18252(.S(\nbus_14028[0] ), .A(\tab23[10] ), .B(n_52222), .Z
		(n_12361));
	notech_and4 i_1722232(.A(n_1236), .B(n_1238), .C(n_1235), .D(n_725), .Z(n_53150
		));
	notech_reg_set tab23_reg_11(.CP(n_62083), .D(n_12367), .SD(n_61399), .Q(\tab23[11] 
		));
	notech_mux2 i_18260(.S(\nbus_14028[0] ), .A(\tab23[11] ), .B(n_52228), .Z
		(n_12367));
	notech_and4 i_1822233(.A(n_1227), .B(n_1229), .C(n_1226), .D(n_736), .Z(n_53157
		));
	notech_reg_set tab23_reg_12(.CP(n_62083), .D(n_12373), .SD(n_61399), .Q(\tab23[12] 
		));
	notech_mux2 i_18268(.S(\nbus_14028[0] ), .A(\tab23[12] ), .B(n_52234), .Z
		(n_12373));
	notech_and4 i_1922234(.A(n_1218), .B(n_1220), .C(n_1217), .D(n_747), .Z(n_53164
		));
	notech_reg_set tab23_reg_13(.CP(n_62078), .D(n_12379), .SD(n_61394), .Q(\tab23[13] 
		));
	notech_mux2 i_18276(.S(\nbus_14028[0] ), .A(\tab23[13] ), .B(n_52240), .Z
		(n_12379));
	notech_and4 i_2022235(.A(n_1209), .B(n_1211), .C(n_1208), .D(n_758), .Z(n_53171
		));
	notech_reg_set tab23_reg_14(.CP(n_62069), .D(n_12385), .SD(n_61385), .Q(\tab23[14] 
		));
	notech_mux2 i_18284(.S(\nbus_14028[0] ), .A(\tab23[14] ), .B(n_52246), .Z
		(n_12385));
	notech_and4 i_2122236(.A(n_1200), .B(n_1202), .C(n_1199), .D(n_769), .Z(n_53178
		));
	notech_reg_set tab23_reg_15(.CP(n_62069), .D(n_12391), .SD(n_61385), .Q(\tab23[15] 
		));
	notech_mux2 i_18292(.S(\nbus_14028[0] ), .A(\tab23[15] ), .B(n_52252), .Z
		(n_12391));
	notech_and4 i_2222237(.A(n_1191), .B(n_1193), .C(n_1190), .D(n_780), .Z(n_53185
		));
	notech_reg_set tab23_reg_16(.CP(n_62069), .D(n_12397), .SD(n_61385), .Q(\tab23[16] 
		));
	notech_mux2 i_18300(.S(\nbus_14028[0] ), .A(\tab23[16] ), .B(n_52258), .Z
		(n_12397));
	notech_and4 i_2322238(.A(n_1182), .B(n_1184), .C(n_1181), .D(n_791), .Z(n_53192
		));
	notech_reg_set tab23_reg_17(.CP(n_62069), .D(n_12403), .SD(n_61385), .Q(\tab23[17] 
		));
	notech_mux2 i_18308(.S(n_55291), .A(\tab23[17] ), .B(n_52264), .Z(n_12403
		));
	notech_and4 i_2422239(.A(n_1173), .B(n_1175), .C(n_1172), .D(n_802), .Z(n_53199
		));
	notech_reg_set tab23_reg_18(.CP(n_62069), .D(n_12409), .SD(n_61385), .Q(\tab23[18] 
		));
	notech_mux2 i_18316(.S(n_55291), .A(\tab23[18] ), .B(n_52270), .Z(n_12409
		));
	notech_and4 i_2522240(.A(n_1164), .B(n_1166), .C(n_1163), .D(n_813), .Z(n_53206
		));
	notech_reg_set tab23_reg_19(.CP(n_62069), .D(n_12415), .SD(n_61385), .Q(\tab23[19] 
		));
	notech_mux2 i_18324(.S(n_55291), .A(\tab23[19] ), .B(n_52276), .Z(n_12415
		));
	notech_and4 i_2622241(.A(n_1155), .B(n_1157), .C(n_1154), .D(n_824), .Z(n_53213
		));
	notech_reg_set tab23_reg_20(.CP(n_62069), .D(n_12421), .SD(n_61385), .Q(\tab23[20] 
		));
	notech_mux2 i_18332(.S(n_55291), .A(\tab23[20] ), .B(n_52282), .Z(n_12421
		));
	notech_and4 i_2722242(.A(n_1146), .B(n_1148), .C(n_1145), .D(n_835), .Z(n_53220
		));
	notech_reg_set tab23_reg_21(.CP(n_62069), .D(n_12427), .SD(n_61385), .Q(\tab23[21] 
		));
	notech_mux2 i_18340(.S(n_55291), .A(\tab23[21] ), .B(n_52288), .Z(n_12427
		));
	notech_and4 i_2822243(.A(n_1137), .B(n_1139), .C(n_1136), .D(n_846), .Z(n_53227
		));
	notech_reg_set tab23_reg_22(.CP(n_62069), .D(n_12433), .SD(n_61385), .Q(\tab23[22] 
		));
	notech_mux2 i_18348(.S(n_55291), .A(\tab23[22] ), .B(n_52294), .Z(n_12433
		));
	notech_and4 i_2922244(.A(n_1128), .B(n_1130), .C(n_1127), .D(n_857), .Z(n_53234
		));
	notech_reg_set tab23_reg_23(.CP(n_62072), .D(n_12439), .SD(n_61388), .Q(\tab23[23] 
		));
	notech_mux2 i_18356(.S(n_55291), .A(\tab23[23] ), .B(n_52300), .Z(n_12439
		));
	notech_and4 i_3022245(.A(n_1119), .B(n_1121), .C(n_1118), .D(n_868), .Z(n_53241
		));
	notech_reg_set tab23_reg_24(.CP(n_62072), .D(n_12445), .SD(n_61388), .Q(\tab23[24] 
		));
	notech_mux2 i_18364(.S(n_55291), .A(\tab23[24] ), .B(n_52306), .Z(n_12445
		));
	notech_and4 i_3122246(.A(n_1110), .B(n_1112), .C(n_1109), .D(n_879), .Z(n_53248
		));
	notech_reg_set tab23_reg_25(.CP(n_62072), .D(n_12451), .SD(n_61388), .Q(\tab23[25] 
		));
	notech_mux2 i_18372(.S(n_55291), .A(\tab23[25] ), .B(n_52312), .Z(n_12451
		));
	notech_and4 i_3222247(.A(n_1101), .B(n_1103), .C(n_1095), .D(n_890), .Z(n_53255
		));
	notech_reg_set tab23_reg_26(.CP(n_62072), .D(n_12457), .SD(n_61388), .Q(\tab23[26] 
		));
	notech_mux2 i_18380(.S(n_55291), .A(\tab23[26] ), .B(n_52318), .Z(n_12457
		));
	notech_mux2 i_1(.S(n_1015), .A(wrD[0]), .B(iwrite_data[0]), .Z(n_53527)
		);
	notech_reg_set tab23_reg_27(.CP(n_62072), .D(n_12463), .SD(n_61388), .Q(\tab23[27] 
		));
	notech_mux2 i_18388(.S(\nbus_14028[0] ), .A(\tab23[27] ), .B(n_52324), .Z
		(n_12463));
	notech_mux2 i_222150(.S(n_1015), .A(wrD[1]), .B(iwrite_data[1]), .Z(n_53534
		));
	notech_reg_set tab23_reg_28(.CP(n_62069), .D(n_12469), .SD(n_61385), .Q(\tab23[28] 
		));
	notech_mux2 i_18396(.S(n_55291), .A(\tab23[28] ), .B(n_52330), .Z(n_12469
		));
	notech_mux2 i_3(.S(n_1015), .A(wrD[2]), .B(iwrite_data[2]), .Z(n_53541)
		);
	notech_reg_set tab23_reg_29(.CP(n_62069), .D(n_12475), .SD(n_61385), .Q(\tab23[29] 
		));
	notech_mux2 i_18404(.S(n_55291), .A(\tab23[29] ), .B(n_52336), .Z(n_12475
		));
	notech_mux2 i_4(.S(n_1015), .A(wrD[3]), .B(iwrite_data[3]), .Z(n_53548)
		);
	notech_reg tab23_reg_30(.CP(n_62072), .D(n_12481), .CD(n_61388), .Q(\tab23[30] 
		));
	notech_mux2 i_18412(.S(n_55291), .A(\tab23[30] ), .B(n_947), .Z(n_12481)
		);
	notech_mux2 i_522151(.S(n_1015), .A(wrD[4]), .B(iwrite_data[4]), .Z(n_53555
		));
	notech_reg tab23_reg_32(.CP(n_62069), .D(n_12487), .CD(n_61385), .Q(\tab23[32] 
		));
	notech_mux2 i_18420(.S(n_55291), .A(\tab23[32] ), .B(n_948), .Z(n_12487)
		);
	notech_mux2 i_6(.S(n_1015), .A(wrD[5]), .B(iwrite_data[5]), .Z(n_53562)
		);
	notech_reg_set tab23_reg_33(.CP(n_62068), .D(n_12493), .SD(n_61384), .Q(\tab23[33] 
		));
	notech_mux2 i_18428(.S(n_55291), .A(\tab23[33] ), .B(n_55323), .Z(n_12493
		));
	notech_mux2 i_7(.S(n_1015), .A(wrD[6]), .B(iwrite_data[6]), .Z(n_53569)
		);
	notech_reg pg_fault_reg(.CP(n_62068), .D(n_12499), .CD(n_61384), .Q(pg_fault
		));
	notech_mux2 i_18436(.S(n_52374), .A(pg_fault), .B(n_13595), .Z(n_12499)
		);
	notech_mux2 i_8(.S(n_54285), .A(wrD[7]), .B(iwrite_data[7]), .Z(n_53576)
		);
	notech_reg hit_adr23_reg(.CP(n_62068), .D(n_12505), .CD(n_61384), .Q(hit_adr23
		));
	notech_mux2 i_18444(.S(n_945), .A(hit_add23), .B(hit_adr23), .Z(n_12505)
		);
	notech_mux2 i_9(.S(n_54281), .A(wrD[8]), .B(iwrite_data[8]), .Z(n_53583)
		);
	notech_reg owrite_req_reg(.CP(n_62068), .D(n_55935), .CD(n_61384), .Q(owrite_req
		));
	notech_reg addr_miss_reg_0(.CP(n_62068), .D(n_12516), .CD(n_61384), .Q(addr_miss
		[0]));
	notech_and3 i_18458(.A(n_1023), .B(n_636), .C(addr_miss[0]), .Z(n_12516)
		);
	notech_mux2 i_10(.S(n_54281), .A(wrD[9]), .B(iwrite_data[9]), .Z(n_53590
		));
	notech_reg addr_miss_reg_1(.CP(n_62068), .D(n_12522), .CD(n_61384), .Q(addr_miss
		[1]));
	notech_and3 i_18466(.A(n_1023), .B(n_636), .C(addr_miss[1]), .Z(n_12522)
		);
	notech_mux2 i_11(.S(n_54281), .A(wrD[10]), .B(iwrite_data[10]), .Z(n_53597
		));
	notech_reg addr_miss_reg_2(.CP(n_62068), .D(n_12525), .CD(n_61384), .Q(addr_miss
		[2]));
	notech_mux2 i_18472(.S(\nbus_14038[0] ), .A(addr_miss[2]), .B(n_13596), 
		.Z(n_12525));
	notech_mux2 i_12(.S(n_54281), .A(wrD[11]), .B(iwrite_data[11]), .Z(n_53604
		));
	notech_reg addr_miss_reg_3(.CP(n_62068), .D(n_12531), .CD(n_61384), .Q(addr_miss
		[3]));
	notech_mux2 i_18480(.S(\nbus_14038[0] ), .A(addr_miss[3]), .B(n_13597), 
		.Z(n_12531));
	notech_mux2 i_13(.S(n_54281), .A(wrD[12]), .B(iwrite_data[12]), .Z(n_53611
		));
	notech_reg addr_miss_reg_4(.CP(n_62068), .D(n_12537), .CD(n_61384), .Q(addr_miss
		[4]));
	notech_mux2 i_18488(.S(\nbus_14038[0] ), .A(addr_miss[4]), .B(n_13598), 
		.Z(n_12537));
	notech_mux2 i_14(.S(n_54281), .A(wrD[13]), .B(iwrite_data[13]), .Z(n_53618
		));
	notech_reg addr_miss_reg_5(.CP(n_62069), .D(n_12543), .CD(n_61385), .Q(addr_miss
		[5]));
	notech_mux2 i_18496(.S(\nbus_14038[0] ), .A(addr_miss[5]), .B(n_13599), 
		.Z(n_12543));
	notech_mux2 i_15(.S(n_54281), .A(wrD[14]), .B(iwrite_data[14]), .Z(n_53625
		));
	notech_reg addr_miss_reg_6(.CP(n_62069), .D(n_12549), .CD(n_61385), .Q(addr_miss
		[6]));
	notech_mux2 i_18504(.S(\nbus_14038[0] ), .A(addr_miss[6]), .B(n_13600), 
		.Z(n_12549));
	notech_mux2 i_16(.S(n_54281), .A(wrD[15]), .B(iwrite_data[15]), .Z(n_53632
		));
	notech_reg addr_miss_reg_7(.CP(n_62069), .D(n_12555), .CD(n_61385), .Q(addr_miss
		[7]));
	notech_mux2 i_18512(.S(\nbus_14038[0] ), .A(addr_miss[7]), .B(n_13601), 
		.Z(n_12555));
	notech_mux2 i_17(.S(n_54281), .A(wrD[16]), .B(iwrite_data[16]), .Z(n_53639
		));
	notech_reg addr_miss_reg_8(.CP(n_62069), .D(n_12561), .CD(n_61385), .Q(addr_miss
		[8]));
	notech_mux2 i_18520(.S(\nbus_14038[0] ), .A(addr_miss[8]), .B(n_13602), 
		.Z(n_12561));
	notech_mux2 i_18(.S(n_54281), .A(wrD[17]), .B(iwrite_data[17]), .Z(n_53646
		));
	notech_reg addr_miss_reg_9(.CP(n_62069), .D(n_12567), .CD(n_61385), .Q(addr_miss
		[9]));
	notech_mux2 i_18528(.S(\nbus_14038[0] ), .A(addr_miss[9]), .B(n_13603), 
		.Z(n_12567));
	notech_mux2 i_19(.S(n_54281), .A(wrD[18]), .B(iwrite_data[18]), .Z(n_53653
		));
	notech_reg addr_miss_reg_10(.CP(n_62069), .D(n_12573), .CD(n_61385), .Q(addr_miss
		[10]));
	notech_mux2 i_18536(.S(\nbus_14038[0] ), .A(addr_miss[10]), .B(n_13604),
		 .Z(n_12573));
	notech_mux2 i_20(.S(n_54281), .A(wrD[19]), .B(iwrite_data[19]), .Z(n_53660
		));
	notech_reg addr_miss_reg_11(.CP(n_62068), .D(n_12579), .CD(n_61384), .Q(addr_miss
		[11]));
	notech_mux2 i_18544(.S(\nbus_14038[0] ), .A(addr_miss[11]), .B(n_13605),
		 .Z(n_12579));
	notech_mux2 i_21(.S(n_54285), .A(wrD[20]), .B(iwrite_data[20]), .Z(n_53667
		));
	notech_reg addr_miss_reg_12(.CP(n_62069), .D(n_12585), .CD(n_61385), .Q(addr_miss
		[12]));
	notech_mux2 i_18552(.S(\nbus_14038[0] ), .A(addr_miss[12]), .B(n_55155),
		 .Z(n_12585));
	notech_mux2 i_22(.S(n_54285), .A(wrD[21]), .B(iwrite_data[21]), .Z(n_53674
		));
	notech_reg addr_miss_reg_13(.CP(n_62069), .D(n_12591), .CD(n_61385), .Q(addr_miss
		[13]));
	notech_mux2 i_18560(.S(\nbus_14038[0] ), .A(addr_miss[13]), .B(n_55161),
		 .Z(n_12591));
	notech_mux2 i_23(.S(n_54285), .A(wrD[22]), .B(iwrite_data[22]), .Z(n_53681
		));
	notech_reg addr_miss_reg_14(.CP(n_62072), .D(n_12597), .CD(n_61388), .Q(addr_miss
		[14]));
	notech_mux2 i_18568(.S(\nbus_14038[0] ), .A(addr_miss[14]), .B(n_55167),
		 .Z(n_12597));
	notech_mux2 i_24(.S(n_54285), .A(wrD[23]), .B(iwrite_data[23]), .Z(n_53688
		));
	notech_reg addr_miss_reg_15(.CP(n_62077), .D(n_12603), .CD(n_61393), .Q(addr_miss
		[15]));
	notech_mux2 i_18576(.S(\nbus_14038[0] ), .A(addr_miss[15]), .B(n_55173),
		 .Z(n_12603));
	notech_mux2 i_25(.S(n_54285), .A(wrD[24]), .B(iwrite_data[24]), .Z(n_53695
		));
	notech_reg addr_miss_reg_16(.CP(n_62074), .D(n_12609), .CD(n_61390), .Q(addr_miss
		[16]));
	notech_mux2 i_18584(.S(\nbus_14038[0] ), .A(addr_miss[16]), .B(n_55179),
		 .Z(n_12609));
	notech_mux2 i_26(.S(n_54285), .A(wrD[25]), .B(iwrite_data[25]), .Z(n_53702
		));
	notech_reg addr_miss_reg_17(.CP(n_62077), .D(n_12615), .CD(n_61393), .Q(addr_miss
		[17]));
	notech_mux2 i_18592(.S(n_55469), .A(addr_miss[17]), .B(n_55185), .Z(n_12615
		));
	notech_mux2 i_27(.S(n_54281), .A(wrD[26]), .B(iwrite_data[26]), .Z(n_53709
		));
	notech_reg addr_miss_reg_18(.CP(n_62077), .D(n_12621), .CD(n_61393), .Q(addr_miss
		[18]));
	notech_mux2 i_18600(.S(n_55469), .A(addr_miss[18]), .B(n_55191), .Z(n_12621
		));
	notech_mux2 i_28(.S(n_54281), .A(wrD[27]), .B(iwrite_data[27]), .Z(n_53716
		));
	notech_reg addr_miss_reg_19(.CP(n_62074), .D(n_12627), .CD(n_61390), .Q(addr_miss
		[19]));
	notech_mux2 i_18608(.S(n_55469), .A(addr_miss[19]), .B(n_55197), .Z(n_12627
		));
	notech_mux2 i_29(.S(n_54281), .A(wrD[28]), .B(iwrite_data[28]), .Z(n_53723
		));
	notech_reg addr_miss_reg_20(.CP(n_62074), .D(n_12633), .CD(n_61390), .Q(addr_miss
		[20]));
	notech_mux2 i_18616(.S(n_55469), .A(addr_miss[20]), .B(n_55203), .Z(n_12633
		));
	notech_mux2 i_30(.S(n_54285), .A(wrD[29]), .B(iwrite_data[29]), .Z(n_53730
		));
	notech_reg addr_miss_reg_21(.CP(n_62074), .D(n_12639), .CD(n_61390), .Q(addr_miss
		[21]));
	notech_mux2 i_18624(.S(n_55469), .A(addr_miss[21]), .B(n_55209), .Z(n_12639
		));
	notech_mux2 i_31(.S(n_54285), .A(wrD[30]), .B(iwrite_data[30]), .Z(n_53737
		));
	notech_reg addr_miss_reg_22(.CP(n_62074), .D(n_12645), .CD(n_61390), .Q(addr_miss
		[22]));
	notech_mux2 i_18632(.S(n_55469), .A(addr_miss[22]), .B(n_55215), .Z(n_12645
		));
	notech_mux2 i_32(.S(n_54285), .A(wrD[31]), .B(iwrite_data[31]), .Z(n_53744
		));
	notech_reg addr_miss_reg_23(.CP(n_62074), .D(n_12651), .CD(n_61390), .Q(addr_miss
		[23]));
	notech_mux2 i_18640(.S(n_55469), .A(addr_miss[23]), .B(n_55221), .Z(n_12651
		));
	notech_nand2 i_39(.A(n_1004), .B(n_996), .Z(n_52420));
	notech_reg addr_miss_reg_24(.CP(n_62077), .D(n_12657), .CD(n_61393), .Q(addr_miss
		[24]));
	notech_mux2 i_18648(.S(n_55469), .A(addr_miss[24]), .B(n_55227), .Z(n_12657
		));
	notech_or2 i_76273(.A(n_947), .B(data_miss[6]), .Z(n_52426));
	notech_reg addr_miss_reg_25(.CP(n_62077), .D(n_12663), .CD(n_61393), .Q(addr_miss
		[25]));
	notech_mux2 i_18656(.S(n_55469), .A(addr_miss[25]), .B(n_55233), .Z(n_12663
		));
	notech_nand3 i_75871(.A(n_902), .B(n_901), .C(n_491), .Z(n_54378));
	notech_reg addr_miss_reg_26(.CP(n_62078), .D(n_12669), .CD(n_61394), .Q(addr_miss
		[26]));
	notech_mux2 i_18664(.S(n_55469), .A(addr_miss[26]), .B(n_55239), .Z(n_12669
		));
	notech_reg addr_miss_reg_27(.CP(n_62077), .D(n_12675), .CD(n_61393), .Q(addr_miss
		[27]));
	notech_mux2 i_18672(.S(n_55469), .A(addr_miss[27]), .B(n_55245), .Z(n_12675
		));
	notech_ao4 i_75774(.A(n_55449), .B(n_13744), .C(n_999), .D(n_13754), .Z(n_55095
		));
	notech_reg addr_miss_reg_28(.CP(n_62077), .D(n_12681), .CD(n_61393), .Q(addr_miss
		[28]));
	notech_mux2 i_18680(.S(n_55469), .A(addr_miss[28]), .B(n_55251), .Z(n_12681
		));
	notech_ao4 i_75777(.A(n_55449), .B(n_13743), .C(n_999), .D(n_13753), .Z(n_55101
		));
	notech_reg addr_miss_reg_29(.CP(n_62077), .D(n_12687), .CD(n_61393), .Q(addr_miss
		[29]));
	notech_mux2 i_18688(.S(n_55469), .A(addr_miss[29]), .B(n_55257), .Z(n_12687
		));
	notech_ao4 i_75780(.A(n_55449), .B(n_13742), .C(n_999), .D(n_13752), .Z(n_55107
		));
	notech_reg addr_miss_reg_30(.CP(n_62077), .D(n_12693), .CD(n_61393), .Q(addr_miss
		[30]));
	notech_mux2 i_18696(.S(n_55469), .A(addr_miss[30]), .B(n_55263), .Z(n_12693
		));
	notech_ao4 i_75783(.A(n_55449), .B(n_13741), .C(n_999), .D(n_13751), .Z(n_55113
		));
	notech_reg addr_miss_reg_31(.CP(n_62077), .D(n_12699), .CD(n_61393), .Q(addr_miss
		[31]));
	notech_mux2 i_18704(.S(n_55469), .A(addr_miss[31]), .B(n_55269), .Z(n_12699
		));
	notech_ao4 i_75786(.A(n_55449), .B(n_13740), .C(n_999), .D(n_13750), .Z(n_55119
		));
	notech_reg req_miss_reg(.CP(n_62077), .D(n_12705), .CD(n_61393), .Q(req_miss
		));
	notech_or2 i_18712(.A(n_12707), .B(n_12708), .Z(n_12705));
	notech_ao4 i_18713(.A(n_13436), .B(n_13437), .C(n_55469), .D(n_13448), .Z
		(n_12707));
	notech_and4 i_18714(.A(req_miss), .B(n_1023), .C(n_636), .D(n_494), .Z(n_12708
		));
	notech_ao4 i_75789(.A(n_55449), .B(n_13739), .C(n_999), .D(n_13749), .Z(n_55125
		));
	notech_reg oread_req_reg(.CP(n_62072), .D(n_54378), .CD(n_61388), .Q(oread_req
		));
	notech_reg owrite_sz_reg_0(.CP(n_62072), .D(n_899), .CD(n_61388), .Q(owrite_sz
		[0]));
	notech_reg owrite_sz_reg_1(.CP(n_62072), .D(n_900), .CD(n_61388), .Q(owrite_sz
		[1]));
	notech_reg wr_fault_reg(.CP(n_62072), .D(n_12717), .CD(n_61388), .Q(wr_fault
		));
	notech_mux2 i_18732(.S(n_53974), .A(wr_fault), .B(n_898), .Z(n_12717));
	notech_ao4 i_75792(.A(n_55449), .B(n_13738), .C(n_999), .D(n_13748), .Z(n_55131
		));
	notech_reg wrD_reg_0(.CP(n_62072), .D(n_12728), .CD(n_61388), .Q(wrD[0])
		);
	notech_ao4 i_75795(.A(n_55449), .B(n_13737), .C(n_999), .D(n_13747), .Z(n_55137
		));
	notech_nao3 i_18745(.A(\nbus_14013[0] ), .B(1'b1), .C(wrD[0]), .Z(n_12728
		));
	notech_reg wrD_reg_1(.CP(n_62072), .D(n_12729), .CD(n_61388), .Q(wrD[1])
		);
	notech_mux2 i_18748(.S(n_54167), .A(wrD[1]), .B(data_miss[1]), .Z(n_12729
		));
	notech_ao4 i_75798(.A(n_55449), .B(n_13736), .C(n_999), .D(n_13746), .Z(n_55143
		));
	notech_reg wrD_reg_2(.CP(n_62072), .D(n_12735), .CD(n_61388), .Q(wrD[2])
		);
	notech_mux2 i_18756(.S(n_54167), .A(wrD[2]), .B(data_miss[2]), .Z(n_12735
		));
	notech_ao4 i_75801(.A(n_55449), .B(n_13735), .C(n_999), .D(n_13745), .Z(n_55149
		));
	notech_reg wrD_reg_3(.CP(n_62072), .D(n_12741), .CD(n_61388), .Q(wrD[3])
		);
	notech_mux2 i_18764(.S(n_54167), .A(wrD[3]), .B(data_miss[3]), .Z(n_12741
		));
	notech_nand2 i_75804(.A(n_1075), .B(n_515), .Z(n_55155));
	notech_reg wrD_reg_4(.CP(n_62072), .D(n_12747), .CD(n_61388), .Q(wrD[4])
		);
	notech_mux2 i_18772(.S(n_54167), .A(wrD[4]), .B(data_miss[4]), .Z(n_12747
		));
	notech_nand2 i_75807(.A(n_1074), .B(n_516), .Z(n_55161));
	notech_reg wrD_reg_5(.CP(n_62074), .D(n_12753), .CD(n_61390), .Q(wrD[5])
		);
	notech_mux2 i_18780(.S(n_54167), .A(wrD[5]), .B(n_52420), .Z(n_12753));
	notech_nand2 i_75810(.A(n_1073), .B(n_517), .Z(n_55167));
	notech_reg wrD_reg_6(.CP(n_62074), .D(n_12759), .CD(n_61390), .Q(wrD[6])
		);
	notech_mux2 i_18788(.S(n_54167), .A(wrD[6]), .B(n_52426), .Z(n_12759));
	notech_nand2 i_75813(.A(n_1072), .B(n_518), .Z(n_55173));
	notech_reg wrD_reg_7(.CP(n_62074), .D(n_12765), .CD(n_61390), .Q(wrD[7])
		);
	notech_mux2 i_18796(.S(n_54167), .A(wrD[7]), .B(data_miss[7]), .Z(n_12765
		));
	notech_nand2 i_75816(.A(n_1071), .B(n_519), .Z(n_55179));
	notech_reg wrD_reg_8(.CP(n_62074), .D(n_12771), .CD(n_61390), .Q(wrD[8])
		);
	notech_mux2 i_18804(.S(n_54167), .A(wrD[8]), .B(data_miss[8]), .Z(n_12771
		));
	notech_nand2 i_75819(.A(n_1070), .B(n_520), .Z(n_55185));
	notech_reg wrD_reg_9(.CP(n_62074), .D(n_12777), .CD(n_61390), .Q(wrD[9])
		);
	notech_mux2 i_18812(.S(n_54162), .A(wrD[9]), .B(data_miss[9]), .Z(n_12777
		));
	notech_nand2 i_75822(.A(n_1069), .B(n_521), .Z(n_55191));
	notech_reg wrD_reg_10(.CP(n_62072), .D(n_12783), .CD(n_61388), .Q(wrD[10
		]));
	notech_mux2 i_18820(.S(n_54162), .A(wrD[10]), .B(data_miss[10]), .Z(n_12783
		));
	notech_nand2 i_75825(.A(n_1068), .B(n_522), .Z(n_55197));
	notech_reg wrD_reg_11(.CP(n_62072), .D(n_12789), .CD(n_61388), .Q(wrD[11
		]));
	notech_mux2 i_18828(.S(n_54162), .A(wrD[11]), .B(data_miss[11]), .Z(n_12789
		));
	notech_nand2 i_75828(.A(n_1067), .B(n_523), .Z(n_55203));
	notech_reg wrD_reg_12(.CP(n_62072), .D(n_12795), .CD(n_61388), .Q(wrD[12
		]));
	notech_mux2 i_18836(.S(n_54167), .A(wrD[12]), .B(data_miss[12]), .Z(n_12795
		));
	notech_nand2 i_75831(.A(n_1066), .B(n_524), .Z(n_55209));
	notech_reg wrD_reg_13(.CP(n_62072), .D(n_12801), .CD(n_61388), .Q(wrD[13
		]));
	notech_mux2 i_18844(.S(n_54167), .A(wrD[13]), .B(data_miss[13]), .Z(n_12801
		));
	notech_nand2 i_75834(.A(n_1065), .B(n_525), .Z(n_55215));
	notech_reg wrD_reg_14(.CP(n_62101), .D(n_12807), .CD(n_61417), .Q(wrD[14
		]));
	notech_mux2 i_18852(.S(n_54167), .A(wrD[14]), .B(data_miss[14]), .Z(n_12807
		));
	notech_nand2 i_75837(.A(n_1064), .B(n_526), .Z(n_55221));
	notech_reg wrD_reg_15(.CP(n_62101), .D(n_12813), .CD(n_61417), .Q(wrD[15
		]));
	notech_mux2 i_18860(.S(n_54167), .A(wrD[15]), .B(data_miss[15]), .Z(n_12813
		));
	notech_nand2 i_75840(.A(n_1063), .B(n_527), .Z(n_55227));
	notech_reg wrD_reg_16(.CP(n_62101), .D(n_12819), .CD(n_61417), .Q(wrD[16
		]));
	notech_mux2 i_18868(.S(n_54167), .A(wrD[16]), .B(data_miss[16]), .Z(n_12819
		));
	notech_nand2 i_75843(.A(n_1062), .B(n_528), .Z(n_55233));
	notech_reg wrD_reg_17(.CP(n_62101), .D(n_12825), .CD(n_61417), .Q(wrD[17
		]));
	notech_mux2 i_18876(.S(n_54168), .A(wrD[17]), .B(data_miss[17]), .Z(n_12825
		));
	notech_nand2 i_75846(.A(n_1061), .B(n_529), .Z(n_55239));
	notech_reg wrD_reg_18(.CP(n_62101), .D(n_12831), .CD(n_61417), .Q(wrD[18
		]));
	notech_mux2 i_18884(.S(n_54168), .A(wrD[18]), .B(data_miss[18]), .Z(n_12831
		));
	notech_nand2 i_75849(.A(n_1060), .B(n_530), .Z(n_55245));
	notech_reg wrD_reg_19(.CP(n_62101), .D(n_12837), .CD(n_61417), .Q(wrD[19
		]));
	notech_mux2 i_18892(.S(n_54168), .A(wrD[19]), .B(data_miss[19]), .Z(n_12837
		));
	notech_nand2 i_75852(.A(n_1059), .B(n_531), .Z(n_55251));
	notech_reg wrD_reg_20(.CP(n_62101), .D(n_12843), .CD(n_61417), .Q(wrD[20
		]));
	notech_mux2 i_18900(.S(n_54168), .A(wrD[20]), .B(data_miss[20]), .Z(n_12843
		));
	notech_nand2 i_75855(.A(n_1058), .B(n_532), .Z(n_55257));
	notech_reg wrD_reg_21(.CP(n_62101), .D(n_12849), .CD(n_61417), .Q(wrD[21
		]));
	notech_mux2 i_18908(.S(n_54168), .A(wrD[21]), .B(data_miss[21]), .Z(n_12849
		));
	notech_nand2 i_75858(.A(n_1057), .B(n_533), .Z(n_55263));
	notech_reg wrD_reg_22(.CP(n_62101), .D(n_12855), .CD(n_61417), .Q(wrD[22
		]));
	notech_mux2 i_18916(.S(n_54168), .A(wrD[22]), .B(data_miss[22]), .Z(n_12855
		));
	notech_nand2 i_75861(.A(n_1056), .B(n_534), .Z(n_55269));
	notech_reg wrD_reg_23(.CP(n_62102), .D(n_12861), .CD(n_61418), .Q(wrD[23
		]));
	notech_mux2 i_18924(.S(n_54168), .A(wrD[23]), .B(data_miss[23]), .Z(n_12861
		));
	notech_mux2 i_75768(.S(iwrite_ack), .A(n_538), .B(n_13469), .Z(n_55935)
		);
	notech_reg wrD_reg_24(.CP(n_62102), .D(n_12867), .CD(n_61418), .Q(wrD[24
		]));
	notech_mux2 i_18932(.S(n_54168), .A(wrD[24]), .B(data_miss[24]), .Z(n_12867
		));
	notech_or2 i_69(.A(n_55323), .B(\addr_miss_0[2] ), .Z(n_52162));
	notech_reg wrD_reg_25(.CP(n_62102), .D(n_12873), .CD(n_61418), .Q(wrD[25
		]));
	notech_mux2 i_18940(.S(n_54168), .A(wrD[25]), .B(data_miss[25]), .Z(n_12873
		));
	notech_or2 i_70(.A(n_55323), .B(\addr_miss_0[3] ), .Z(n_52168));
	notech_reg wrD_reg_26(.CP(n_62102), .D(n_12879), .CD(n_61418), .Q(wrD[26
		]));
	notech_mux2 i_18948(.S(n_54168), .A(wrD[26]), .B(data_miss[26]), .Z(n_12879
		));
	notech_or2 i_71(.A(n_55323), .B(\addr_miss_0[4] ), .Z(n_52174));
	notech_reg wrD_reg_27(.CP(n_62102), .D(n_12885), .CD(n_61418), .Q(wrD[27
		]));
	notech_mux2 i_18956(.S(n_54167), .A(wrD[27]), .B(data_miss[27]), .Z(n_12885
		));
	notech_or2 i_72(.A(n_55323), .B(\addr_miss_0[5] ), .Z(n_52180));
	notech_reg wrD_reg_28(.CP(n_62102), .D(n_12891), .CD(n_61418), .Q(wrD[28
		]));
	notech_mux2 i_18964(.S(n_54168), .A(wrD[28]), .B(data_miss[28]), .Z(n_12891
		));
	notech_or2 i_73(.A(n_55323), .B(\addr_miss_0[7] ), .Z(n_52192));
	notech_reg wrD_reg_29(.CP(n_62102), .D(n_12897), .CD(n_61418), .Q(wrD[29
		]));
	notech_mux2 i_18972(.S(n_54168), .A(wrD[29]), .B(data_miss[29]), .Z(n_12897
		));
	notech_or2 i_74(.A(n_55323), .B(\addr_miss_0[8] ), .Z(n_52198));
	notech_reg wrD_reg_30(.CP(n_62102), .D(n_12903), .CD(n_61418), .Q(wrD[30
		]));
	notech_mux2 i_18980(.S(n_54168), .A(wrD[30]), .B(data_miss[30]), .Z(n_12903
		));
	notech_or2 i_75(.A(n_55323), .B(\addr_miss_0[9] ), .Z(n_52204));
	notech_reg wrD_reg_31(.CP(n_62102), .D(n_12909), .CD(n_61418), .Q(wrD[31
		]));
	notech_mux2 i_18988(.S(n_54168), .A(wrD[31]), .B(data_miss[31]), .Z(n_12909
		));
	notech_or2 i_76(.A(n_55323), .B(\addr_miss_0[10] ), .Z(n_52210));
	notech_reg owrite_data_reg_0(.CP(n_62100), .D(n_53527), .CD(n_61416), .Q
		(owrite_data[0]));
	notech_reg owrite_data_reg_1(.CP(n_62100), .D(n_53534), .CD(n_61416), .Q
		(owrite_data[1]));
	notech_reg owrite_data_reg_2(.CP(n_62100), .D(n_53541), .CD(n_61416), .Q
		(owrite_data[2]));
	notech_reg owrite_data_reg_3(.CP(n_62100), .D(n_53548), .CD(n_61416), .Q
		(owrite_data[3]));
	notech_reg owrite_data_reg_4(.CP(n_62098), .D(n_53555), .CD(n_61414), .Q
		(owrite_data[4]));
	notech_reg owrite_data_reg_5(.CP(n_62098), .D(n_53562), .CD(n_61414), .Q
		(owrite_data[5]));
	notech_reg owrite_data_reg_6(.CP(n_62098), .D(n_53569), .CD(n_61414), .Q
		(owrite_data[6]));
	notech_reg owrite_data_reg_7(.CP(n_62098), .D(n_53576), .CD(n_61414), .Q
		(owrite_data[7]));
	notech_reg owrite_data_reg_8(.CP(n_62098), .D(n_53583), .CD(n_61414), .Q
		(owrite_data[8]));
	notech_reg owrite_data_reg_9(.CP(n_62100), .D(n_53590), .CD(n_61416), .Q
		(owrite_data[9]));
	notech_reg owrite_data_reg_10(.CP(n_62100), .D(n_53597), .CD(n_61416), .Q
		(owrite_data[10]));
	notech_reg owrite_data_reg_11(.CP(n_62101), .D(n_53604), .CD(n_61417), .Q
		(owrite_data[11]));
	notech_reg owrite_data_reg_12(.CP(n_62101), .D(n_53611), .CD(n_61417), .Q
		(owrite_data[12]));
	notech_reg owrite_data_reg_13(.CP(n_62100), .D(n_53618), .CD(n_61416), .Q
		(owrite_data[13]));
	notech_reg owrite_data_reg_14(.CP(n_62100), .D(n_53625), .CD(n_61416), .Q
		(owrite_data[14]));
	notech_reg owrite_data_reg_15(.CP(n_62100), .D(n_53632), .CD(n_61416), .Q
		(owrite_data[15]));
	notech_reg owrite_data_reg_16(.CP(n_62100), .D(n_53639), .CD(n_61416), .Q
		(owrite_data[16]));
	notech_reg owrite_data_reg_17(.CP(n_62100), .D(n_53646), .CD(n_61416), .Q
		(owrite_data[17]));
	notech_reg owrite_data_reg_18(.CP(n_62102), .D(n_53653), .CD(n_61418), .Q
		(owrite_data[18]));
	notech_reg owrite_data_reg_19(.CP(n_62107), .D(n_53660), .CD(n_61423), .Q
		(owrite_data[19]));
	notech_reg owrite_data_reg_20(.CP(n_62107), .D(n_53667), .CD(n_61423), .Q
		(owrite_data[20]));
	notech_reg owrite_data_reg_21(.CP(n_62107), .D(n_53674), .CD(n_61423), .Q
		(owrite_data[21]));
	notech_reg owrite_data_reg_22(.CP(n_62107), .D(n_53681), .CD(n_61423), .Q
		(owrite_data[22]));
	notech_reg owrite_data_reg_23(.CP(n_62106), .D(n_53688), .CD(n_61422), .Q
		(owrite_data[23]));
	notech_reg owrite_data_reg_24(.CP(n_62106), .D(n_53695), .CD(n_61422), .Q
		(owrite_data[24]));
	notech_reg owrite_data_reg_25(.CP(n_62106), .D(n_53702), .CD(n_61422), .Q
		(owrite_data[25]));
	notech_reg owrite_data_reg_26(.CP(n_62106), .D(n_53709), .CD(n_61422), .Q
		(owrite_data[26]));
	notech_reg owrite_data_reg_27(.CP(n_62106), .D(n_53716), .CD(n_61422), .Q
		(owrite_data[27]));
	notech_reg owrite_data_reg_28(.CP(n_62107), .D(n_53723), .CD(n_61423), .Q
		(owrite_data[28]));
	notech_reg owrite_data_reg_29(.CP(n_62107), .D(n_53730), .CD(n_61423), .Q
		(owrite_data[29]));
	notech_reg owrite_data_reg_30(.CP(n_62109), .D(n_53737), .CD(n_61425), .Q
		(owrite_data[30]));
	notech_reg owrite_data_reg_31(.CP(n_62109), .D(n_53744), .CD(n_61425), .Q
		(owrite_data[31]));
	notech_reg pt_fault_reg(.CP(n_62107), .D(n_12979), .CD(n_61423), .Q(pt_fault
		));
	notech_mux2 i_19124(.S(n_897), .A(data_miss[0]), .B(pt_fault), .Z(n_12979
		));
	notech_or2 i_77(.A(n_55323), .B(\addr_miss_0[11] ), .Z(n_52216));
	notech_reg cr2_reg_0(.CP(n_62107), .D(n_12985), .CD(n_61423), .Q(cr2[0])
		);
	notech_mux2 i_19132(.S(n_897), .A(iDaddr_f[0]), .B(cr2[0]), .Z(n_12985)
		);
	notech_or2 i_78(.A(data_miss[12]), .B(n_55323), .Z(n_52222));
	notech_reg cr2_reg_1(.CP(n_62107), .D(n_12991), .CD(n_61423), .Q(cr2[1])
		);
	notech_mux2 i_19140(.S(n_897), .A(iDaddr_f[1]), .B(cr2[1]), .Z(n_12991)
		);
	notech_or2 i_79(.A(data_miss[13]), .B(n_55323), .Z(n_52228));
	notech_reg cr2_reg_2(.CP(n_62107), .D(n_12997), .CD(n_61423), .Q(cr2[2])
		);
	notech_mux2 i_19148(.S(n_897), .A(iDaddr_f[2]), .B(cr2[2]), .Z(n_12997)
		);
	notech_or2 i_80(.A(data_miss[14]), .B(n_55318), .Z(n_52234));
	notech_reg cr2_reg_3(.CP(n_62107), .D(n_13003), .CD(n_61423), .Q(cr2[3])
		);
	notech_mux2 i_19156(.S(n_897), .A(iDaddr_f[3]), .B(cr2[3]), .Z(n_13003)
		);
	notech_or2 i_81(.A(data_miss[15]), .B(n_55318), .Z(n_52240));
	notech_reg cr2_reg_4(.CP(n_62105), .D(n_13009), .CD(n_61421), .Q(cr2[4])
		);
	notech_mux2 i_19164(.S(n_897), .A(iDaddr_f[4]), .B(cr2[4]), .Z(n_13009)
		);
	notech_or2 i_82(.A(data_miss[16]), .B(n_55318), .Z(n_52246));
	notech_reg cr2_reg_5(.CP(n_62105), .D(n_13015), .CD(n_61421), .Q(cr2[5])
		);
	notech_mux2 i_19172(.S(n_897), .A(iDaddr_f[5]), .B(cr2[5]), .Z(n_13015)
		);
	notech_or2 i_83(.A(data_miss[17]), .B(n_55318), .Z(n_52252));
	notech_reg cr2_reg_6(.CP(n_62105), .D(n_13021), .CD(n_61421), .Q(cr2[6])
		);
	notech_mux2 i_19180(.S(n_897), .A(iDaddr_f[6]), .B(cr2[6]), .Z(n_13021)
		);
	notech_or2 i_84(.A(data_miss[18]), .B(n_55318), .Z(n_52258));
	notech_reg cr2_reg_7(.CP(n_62105), .D(n_13027), .CD(n_61421), .Q(cr2[7])
		);
	notech_mux2 i_19188(.S(n_897), .A(iDaddr_f[7]), .B(cr2[7]), .Z(n_13027)
		);
	notech_or2 i_85(.A(data_miss[19]), .B(n_55318), .Z(n_52264));
	notech_reg cr2_reg_8(.CP(n_62105), .D(n_13033), .CD(n_61421), .Q(cr2[8])
		);
	notech_mux2 i_19196(.S(n_897), .A(iDaddr_f[8]), .B(cr2[8]), .Z(n_13033)
		);
	notech_or2 i_86(.A(data_miss[20]), .B(n_55318), .Z(n_52270));
	notech_reg cr2_reg_9(.CP(n_62105), .D(n_13039), .CD(n_61421), .Q(cr2[9])
		);
	notech_mux2 i_19204(.S(n_897), .A(iDaddr_f[9]), .B(cr2[9]), .Z(n_13039)
		);
	notech_or2 i_87(.A(data_miss[21]), .B(n_55318), .Z(n_52276));
	notech_reg cr2_reg_10(.CP(n_62102), .D(n_13045), .CD(n_61418), .Q(cr2[10
		]));
	notech_mux2 i_19212(.S(n_897), .A(iDaddr_f[10]), .B(cr2[10]), .Z(n_13045
		));
	notech_or2 i_88(.A(data_miss[22]), .B(n_55318), .Z(n_52282));
	notech_reg cr2_reg_11(.CP(n_62105), .D(n_13051), .CD(n_61421), .Q(cr2[11
		]));
	notech_mux2 i_19220(.S(n_897), .A(iDaddr_f[11]), .B(cr2[11]), .Z(n_13051
		));
	notech_or2 i_89(.A(data_miss[23]), .B(n_55318), .Z(n_52288));
	notech_reg cr2_reg_12(.CP(n_62105), .D(n_13057), .CD(n_61421), .Q(cr2[12
		]));
	notech_mux2 i_19228(.S(n_897), .A(iDaddr_f[12]), .B(cr2[12]), .Z(n_13057
		));
	notech_or2 i_90(.A(data_miss[24]), .B(n_55318), .Z(n_52294));
	notech_reg cr2_reg_13(.CP(n_62106), .D(n_13063), .CD(n_61422), .Q(cr2[13
		]));
	notech_mux2 i_19236(.S(n_897), .A(iDaddr_f[13]), .B(cr2[13]), .Z(n_13063
		));
	notech_or2 i_91(.A(data_miss[25]), .B(n_55323), .Z(n_52300));
	notech_reg cr2_reg_14(.CP(n_62106), .D(n_13069), .CD(n_61422), .Q(cr2[14
		]));
	notech_mux2 i_19244(.S(n_897), .A(iDaddr_f[14]), .B(cr2[14]), .Z(n_13069
		));
	notech_or2 i_92(.A(data_miss[26]), .B(n_55318), .Z(n_52306));
	notech_reg cr2_reg_15(.CP(n_62106), .D(n_13075), .CD(n_61422), .Q(cr2[15
		]));
	notech_mux2 i_19252(.S(n_897), .A(iDaddr_f[15]), .B(cr2[15]), .Z(n_13075
		));
	notech_or2 i_93(.A(data_miss[27]), .B(n_55318), .Z(n_52312));
	notech_reg cr2_reg_16(.CP(n_62106), .D(n_13081), .CD(n_61422), .Q(cr2[16
		]));
	notech_mux2 i_19260(.S(n_54493), .A(iDaddr_f[16]), .B(cr2[16]), .Z(n_13081
		));
	notech_or2 i_94(.A(data_miss[28]), .B(n_55318), .Z(n_52318));
	notech_reg cr2_reg_17(.CP(n_62106), .D(n_13087), .CD(n_61422), .Q(cr2[17
		]));
	notech_mux2 i_19268(.S(n_54493), .A(iDaddr_f[17]), .B(cr2[17]), .Z(n_13087
		));
	notech_or2 i_95(.A(data_miss[29]), .B(n_55318), .Z(n_52324));
	notech_reg cr2_reg_18(.CP(n_62105), .D(n_13093), .CD(n_61421), .Q(cr2[18
		]));
	notech_mux2 i_19276(.S(n_54493), .A(iDaddr_f[18]), .B(cr2[18]), .Z(n_13093
		));
	notech_or2 i_96(.A(data_miss[30]), .B(n_55318), .Z(n_52330));
	notech_reg cr2_reg_19(.CP(n_62105), .D(n_13099), .CD(n_61421), .Q(cr2[19
		]));
	notech_mux2 i_19284(.S(n_54493), .A(iDaddr_f[19]), .B(cr2[19]), .Z(n_13099
		));
	notech_or2 i_97(.A(data_miss[31]), .B(n_55318), .Z(n_52336));
	notech_reg cr2_reg_20(.CP(n_62106), .D(n_13105), .CD(n_61422), .Q(cr2[20
		]));
	notech_mux2 i_19292(.S(n_54493), .A(iDaddr_f[20]), .B(cr2[20]), .Z(n_13105
		));
	notech_nand2 i_030892(.A(n_996), .B(n_59313), .Z(n_52360));
	notech_reg cr2_reg_21(.CP(n_62105), .D(n_13111), .CD(n_61421), .Q(cr2[21
		]));
	notech_mux2 i_19300(.S(n_54493), .A(iDaddr_f[21]), .B(cr2[21]), .Z(n_13111
		));
	notech_ao4 i_76779(.A(n_1004), .B(n_13567), .C(n_544), .D(n_1049), .Z(n_55480
		));
	notech_reg cr2_reg_22(.CP(n_62098), .D(n_13117), .CD(n_61414), .Q(cr2[22
		]));
	notech_mux2 i_19308(.S(n_54493), .A(iDaddr_f[22]), .B(cr2[22]), .Z(n_13117
		));
	notech_ao4 i_76782(.A(n_1004), .B(n_13569), .C(n_549), .D(n_1049), .Z(n_55486
		));
	notech_reg cr2_reg_23(.CP(n_62091), .D(n_13123), .CD(n_61407), .Q(cr2[23
		]));
	notech_mux2 i_19316(.S(n_54493), .A(iDaddr_f[23]), .B(cr2[23]), .Z(n_13123
		));
	notech_ao4 i_76769(.A(n_1004), .B(\nnx_tab2[0] ), .C(n_999), .D(n_13572)
		, .Z(n_54264));
	notech_reg cr2_reg_24(.CP(n_62090), .D(n_13129), .CD(n_61406), .Q(cr2[24
		]));
	notech_mux2 i_19324(.S(n_54493), .A(iDaddr_f[24]), .B(cr2[24]), .Z(n_13129
		));
	notech_ao4 i_76772(.A(n_999), .B(n_13574), .C(n_1004), .D(n_558), .Z(n_54270
		));
	notech_reg cr2_reg_25(.CP(n_62091), .D(n_13135), .CD(n_61407), .Q(cr2[25
		]));
	notech_mux2 i_19332(.S(n_54493), .A(iDaddr_f[25]), .B(cr2[25]), .Z(n_13135
		));
	notech_ao4 i_76625(.A(n_1004), .B(\nnx_tab1[0] ), .C(n_999), .D(n_13517)
		, .Z(n_54299));
	notech_reg cr2_reg_26(.CP(n_62091), .D(n_13141), .CD(n_61407), .Q(cr2[26
		]));
	notech_mux2 i_19340(.S(n_897), .A(iDaddr_f[26]), .B(cr2[26]), .Z(n_13141
		));
	notech_ao4 i_76628(.A(n_999), .B(n_13519), .C(n_1004), .D(n_569), .Z(n_54305
		));
	notech_reg cr2_reg_27(.CP(n_62090), .D(n_13147), .CD(n_61406), .Q(cr2[27
		]));
	notech_mux2 i_19348(.S(n_54493), .A(iDaddr_f[27]), .B(cr2[27]), .Z(n_13147
		));
	notech_ao4 i_76789(.A(n_1004), .B(n_13521), .C(n_574), .D(n_1042), .Z(n_55041
		));
	notech_reg cr2_reg_28(.CP(n_62090), .D(n_13153), .CD(n_61406), .Q(cr2[28
		]));
	notech_mux2 i_19356(.S(n_54493), .A(iDaddr_f[28]), .B(cr2[28]), .Z(n_13153
		));
	notech_ao4 i_76792(.A(n_1004), .B(n_13523), .C(n_579), .D(n_1042), .Z(n_55047
		));
	notech_reg cr2_reg_29(.CP(n_62090), .D(n_13159), .CD(n_61406), .Q(cr2[29
		]));
	notech_mux2 i_19364(.S(n_54493), .A(iDaddr_f[29]), .B(cr2[29]), .Z(n_13159
		));
	notech_nand2 i_130(.A(n_54224), .B(n_13744), .Z(n_54025));
	notech_reg cr2_reg_30(.CP(n_62090), .D(n_13165), .CD(n_61406), .Q(cr2[30
		]));
	notech_mux2 i_19372(.S(n_54493), .A(iDaddr_f[30]), .B(cr2[30]), .Z(n_13165
		));
	notech_nand2 i_131(.A(n_54224), .B(n_13743), .Z(n_54031));
	notech_reg cr2_reg_31(.CP(n_62090), .D(n_13171), .CD(n_61406), .Q(cr2[31
		]));
	notech_mux2 i_19380(.S(n_54493), .A(iDaddr_f[31]), .B(cr2[31]), .Z(n_13171
		));
	notech_nand2 i_132(.A(n_54224), .B(n_13742), .Z(n_54037));
	notech_reg wrA_reg_0(.CP(n_62091), .D(n_13177), .CD(n_61407), .Q(wrA[0])
		);
	notech_mux2 i_19388(.S(n_54162), .A(wrA[0]), .B(addr_miss[0]), .Z(n_13177
		));
	notech_nand2 i_133(.A(n_54224), .B(n_13741), .Z(n_54043));
	notech_reg wrA_reg_1(.CP(n_62091), .D(n_13183), .CD(n_61407), .Q(wrA[1])
		);
	notech_mux2 i_19396(.S(n_54159), .A(wrA[1]), .B(addr_miss[1]), .Z(n_13183
		));
	notech_nand2 i_134(.A(n_54224), .B(n_13739), .Z(n_54055));
	notech_reg wrA_reg_2(.CP(n_62092), .D(n_13189), .CD(n_61408), .Q(wrA[2])
		);
	notech_mux2 i_19404(.S(n_54159), .A(wrA[2]), .B(addr_miss[2]), .Z(n_13189
		));
	notech_nand2 i_135(.A(n_54224), .B(n_13738), .Z(n_54061));
	notech_reg wrA_reg_3(.CP(n_62091), .D(n_13195), .CD(n_61407), .Q(wrA[3])
		);
	notech_mux2 i_19412(.S(n_54159), .A(wrA[3]), .B(addr_miss[3]), .Z(n_13195
		));
	notech_nand2 i_136(.A(n_54224), .B(n_13737), .Z(n_54067));
	notech_reg wrA_reg_4(.CP(n_62091), .D(n_13201), .CD(n_61407), .Q(wrA[4])
		);
	notech_mux2 i_19420(.S(n_54159), .A(wrA[4]), .B(addr_miss[4]), .Z(n_13201
		));
	notech_nand2 i_137(.A(n_54224), .B(n_13736), .Z(n_54073));
	notech_reg wrA_reg_5(.CP(n_62091), .D(n_13207), .CD(n_61407), .Q(wrA[5])
		);
	notech_mux2 i_19428(.S(n_54159), .A(wrA[5]), .B(addr_miss[5]), .Z(n_13207
		));
	notech_nand2 i_138(.A(n_54224), .B(n_13735), .Z(n_54079));
	notech_reg wrA_reg_6(.CP(n_62091), .D(n_13213), .CD(n_61407), .Q(wrA[6])
		);
	notech_mux2 i_19436(.S(n_54159), .A(wrA[6]), .B(addr_miss[6]), .Z(n_13213
		));
	notech_or2 i_139(.A(data_miss[12]), .B(n_13470), .Z(n_54085));
	notech_reg wrA_reg_7(.CP(n_62091), .D(n_13219), .CD(n_61407), .Q(wrA[7])
		);
	notech_mux2 i_19444(.S(n_54159), .A(wrA[7]), .B(addr_miss[7]), .Z(n_13219
		));
	notech_or2 i_140(.A(data_miss[13]), .B(n_13470), .Z(n_54091));
	notech_reg wrA_reg_8(.CP(n_62091), .D(n_13225), .CD(n_61407), .Q(wrA[8])
		);
	notech_mux2 i_19452(.S(n_54159), .A(wrA[8]), .B(addr_miss[8]), .Z(n_13225
		));
	notech_or2 i_141(.A(data_miss[14]), .B(n_13470), .Z(n_54097));
	notech_reg wrA_reg_9(.CP(n_62088), .D(n_13231), .CD(n_61404), .Q(wrA[9])
		);
	notech_mux2 i_19460(.S(n_54158), .A(wrA[9]), .B(addr_miss[9]), .Z(n_13231
		));
	notech_or2 i_142(.A(data_miss[15]), .B(n_13470), .Z(n_54103));
	notech_reg wrA_reg_10(.CP(n_62088), .D(n_13237), .CD(n_61404), .Q(wrA[10
		]));
	notech_mux2 i_19468(.S(n_54158), .A(wrA[10]), .B(addr_miss[10]), .Z(n_13237
		));
	notech_or2 i_143(.A(data_miss[16]), .B(n_13470), .Z(n_54109));
	notech_reg wrA_reg_11(.CP(n_62088), .D(n_13243), .CD(n_61404), .Q(wrA[11
		]));
	notech_mux2 i_19476(.S(n_54158), .A(wrA[11]), .B(addr_miss[11]), .Z(n_13243
		));
	notech_or2 i_144(.A(data_miss[17]), .B(n_13470), .Z(n_54115));
	notech_reg wrA_reg_12(.CP(n_62088), .D(n_13249), .CD(n_61404), .Q(wrA[12
		]));
	notech_mux2 i_19484(.S(n_54158), .A(wrA[12]), .B(addr_miss[12]), .Z(n_13249
		));
	notech_or2 i_145(.A(data_miss[18]), .B(n_13470), .Z(n_54121));
	notech_reg wrA_reg_13(.CP(n_62088), .D(n_13255), .CD(n_61404), .Q(wrA[13
		]));
	notech_mux2 i_19492(.S(n_54158), .A(wrA[13]), .B(addr_miss[13]), .Z(n_13255
		));
	notech_or2 i_146(.A(data_miss[19]), .B(n_13470), .Z(n_54127));
	notech_reg wrA_reg_14(.CP(n_62087), .D(n_13261), .CD(n_61403), .Q(wrA[14
		]));
	notech_mux2 i_19500(.S(n_54158), .A(wrA[14]), .B(addr_miss[14]), .Z(n_13261
		));
	notech_or2 i_147(.A(data_miss[20]), .B(n_13470), .Z(n_54133));
	notech_reg wrA_reg_15(.CP(n_62087), .D(n_13267), .CD(n_61403), .Q(wrA[15
		]));
	notech_mux2 i_19508(.S(n_54158), .A(wrA[15]), .B(addr_miss[15]), .Z(n_13267
		));
	notech_or2 i_148(.A(data_miss[21]), .B(n_55338), .Z(n_54139));
	notech_reg wrA_reg_16(.CP(n_62088), .D(n_13273), .CD(n_61404), .Q(wrA[16
		]));
	notech_mux2 i_19516(.S(n_54159), .A(wrA[16]), .B(addr_miss[16]), .Z(n_13273
		));
	notech_or2 i_149(.A(data_miss[22]), .B(n_55338), .Z(n_54145));
	notech_reg wrA_reg_17(.CP(n_62088), .D(n_13279), .CD(n_61404), .Q(wrA[17
		]));
	notech_mux2 i_19524(.S(n_54162), .A(wrA[17]), .B(addr_miss[17]), .Z(n_13279
		));
	notech_or2 i_150(.A(data_miss[23]), .B(n_55338), .Z(n_54151));
	notech_reg wrA_reg_18(.CP(n_62090), .D(n_13285), .CD(n_61406), .Q(wrA[18
		]));
	notech_mux2 i_19532(.S(n_54162), .A(wrA[18]), .B(addr_miss[18]), .Z(n_13285
		));
	notech_or2 i_151(.A(data_miss[24]), .B(n_55338), .Z(n_54157));
	notech_reg wrA_reg_19(.CP(n_62090), .D(n_13291), .CD(n_61406), .Q(wrA[19
		]));
	notech_mux2 i_19540(.S(n_54162), .A(wrA[19]), .B(addr_miss[19]), .Z(n_13291
		));
	notech_or2 i_152(.A(data_miss[25]), .B(n_55338), .Z(n_54163));
	notech_reg wrA_reg_20(.CP(n_62090), .D(n_13297), .CD(n_61406), .Q(wrA[20
		]));
	notech_mux2 i_19548(.S(n_54162), .A(wrA[20]), .B(addr_miss[20]), .Z(n_13297
		));
	notech_or2 i_153(.A(data_miss[26]), .B(n_55338), .Z(n_54169));
	notech_reg wrA_reg_21(.CP(n_62090), .D(n_13303), .CD(n_61406), .Q(wrA[21
		]));
	notech_mux2 i_19556(.S(n_54162), .A(wrA[21]), .B(addr_miss[21]), .Z(n_13303
		));
	notech_or2 i_154(.A(data_miss[27]), .B(n_55338), .Z(n_54175));
	notech_reg wrA_reg_22(.CP(n_62090), .D(n_13309), .CD(n_61406), .Q(wrA[22
		]));
	notech_mux2 i_19564(.S(n_54162), .A(wrA[22]), .B(addr_miss[22]), .Z(n_13309
		));
	notech_or2 i_155(.A(data_miss[28]), .B(n_13470), .Z(n_54181));
	notech_reg wrA_reg_23(.CP(n_62088), .D(n_13315), .CD(n_61404), .Q(wrA[23
		]));
	notech_mux2 i_19572(.S(n_54162), .A(wrA[23]), .B(addr_miss[23]), .Z(n_13315
		));
	notech_or2 i_156(.A(data_miss[29]), .B(n_55338), .Z(n_54187));
	notech_reg wrA_reg_24(.CP(n_62088), .D(n_13321), .CD(n_61404), .Q(wrA[24
		]));
	notech_mux2 i_19580(.S(n_54162), .A(wrA[24]), .B(addr_miss[24]), .Z(n_13321
		));
	notech_or2 i_157(.A(data_miss[30]), .B(n_55338), .Z(n_54193));
	notech_reg wrA_reg_25(.CP(n_62088), .D(n_13327), .CD(n_61404), .Q(wrA[25
		]));
	notech_mux2 i_19588(.S(n_54159), .A(wrA[25]), .B(addr_miss[25]), .Z(n_13327
		));
	notech_or2 i_158(.A(data_miss[31]), .B(n_55338), .Z(n_54199));
	notech_reg wrA_reg_26(.CP(n_62088), .D(n_13333), .CD(n_61404), .Q(wrA[26
		]));
	notech_mux2 i_19596(.S(n_54159), .A(wrA[26]), .B(addr_miss[26]), .Z(n_13333
		));
	notech_ao4 i_34(.A(data_miss[0]), .B(n_996), .C(n_982), .D(n_983), .Z(n_54224
		));
	notech_reg wrA_reg_27(.CP(n_62092), .D(n_13339), .CD(n_61408), .Q(wrA[27
		]));
	notech_mux2 i_19604(.S(n_54159), .A(wrA[27]), .B(addr_miss[27]), .Z(n_13339
		));
	notech_or4 i_41(.A(n_954), .B(n_1006), .C(n_13473), .D(n_13435), .Z(n_54349
		));
	notech_reg wrA_reg_28(.CP(n_62097), .D(n_13345), .CD(n_61413), .Q(wrA[28
		]));
	notech_mux2 i_19612(.S(n_54159), .A(wrA[28]), .B(addr_miss[28]), .Z(n_13345
		));
	notech_and4 i_42(.A(n_55449), .B(n_1011), .C(n_997), .D(n_960), .Z(n_54355
		));
	notech_reg wrA_reg_29(.CP(n_62097), .D(n_13351), .CD(n_61413), .Q(wrA[29
		]));
	notech_mux2 i_19620(.S(n_54162), .A(wrA[29]), .B(addr_miss[29]), .Z(n_13351
		));
	notech_and4 i_43(.A(n_999), .B(n_998), .C(n_640), .D(n_52377), .Z(n_54361
		));
	notech_reg wrA_reg_30(.CP(n_62097), .D(n_13357), .CD(n_61413), .Q(wrA[30
		]));
	notech_mux2 i_19628(.S(n_54162), .A(wrA[30]), .B(addr_miss[30]), .Z(n_13357
		));
	notech_reg wrA_reg_31(.CP(n_62097), .D(n_13363), .CD(n_61413), .Q(wrA[31
		]));
	notech_mux2 i_19636(.S(n_54159), .A(wrA[31]), .B(addr_miss[31]), .Z(n_13363
		));
	notech_reg addr_phys_reg_0(.CP(n_62097), .D(n_53038), .CD(n_61413), .Q(addr_phys
		[0]));
	notech_reg addr_phys_reg_1(.CP(n_62096), .D(n_53045), .CD(n_61412), .Q(addr_phys
		[1]));
	notech_reg addr_phys_reg_2(.CP(n_62096), .D(n_53052), .CD(n_61412), .Q(addr_phys
		[2]));
	notech_reg addr_phys_reg_3(.CP(n_62097), .D(n_53059), .CD(n_61413), .Q(addr_phys
		[3]));
	notech_reg addr_phys_reg_4(.CP(n_62097), .D(n_53066), .CD(n_61413), .Q(addr_phys
		[4]));
	notech_reg addr_phys_reg_5(.CP(n_62098), .D(n_53073), .CD(n_61414), .Q(addr_phys
		[5]));
	notech_reg addr_phys_reg_6(.CP(n_62098), .D(n_53080), .CD(n_61414), .Q(addr_phys
		[6]));
	notech_reg addr_phys_reg_7(.CP(n_62098), .D(n_53087), .CD(n_61414), .Q(addr_phys
		[7]));
	notech_reg addr_phys_reg_8(.CP(n_62098), .D(n_53094), .CD(n_61414), .Q(addr_phys
		[8]));
	notech_reg addr_phys_reg_9(.CP(n_62098), .D(n_53101), .CD(n_61414), .Q(addr_phys
		[9]));
	notech_reg addr_phys_reg_10(.CP(n_62097), .D(n_53108), .CD(n_61413), .Q(addr_phys
		[10]));
	notech_reg addr_phys_reg_11(.CP(n_62097), .D(n_53115), .CD(n_61413), .Q(addr_phys
		[11]));
	notech_reg addr_phys_reg_12(.CP(n_62097), .D(n_13661), .CD(n_61413), .Q(addr_phys
		[12]));
	notech_reg addr_phys_reg_13(.CP(n_62097), .D(n_13662), .CD(n_61413), .Q(addr_phys
		[13]));
	notech_reg addr_phys_reg_14(.CP(n_62092), .D(n_13663), .CD(n_61408), .Q(addr_phys
		[14]));
	notech_reg addr_phys_reg_15(.CP(n_62092), .D(n_13664), .CD(n_61408), .Q(addr_phys
		[15]));
	notech_reg addr_phys_reg_16(.CP(n_62092), .D(n_13665), .CD(n_61408), .Q(addr_phys
		[16]));
	notech_reg addr_phys_reg_17(.CP(n_62092), .D(n_13666), .CD(n_61408), .Q(addr_phys
		[17]));
	notech_reg addr_phys_reg_18(.CP(n_62092), .D(n_13667), .CD(n_61408), .Q(addr_phys
		[18]));
	notech_reg addr_phys_reg_19(.CP(n_62092), .D(n_13668), .CD(n_61408), .Q(addr_phys
		[19]));
	notech_reg addr_phys_reg_20(.CP(n_62092), .D(n_13669), .CD(n_61408), .Q(addr_phys
		[20]));
	notech_reg addr_phys_reg_21(.CP(n_62092), .D(n_13670), .CD(n_61408), .Q(addr_phys
		[21]));
	notech_reg addr_phys_reg_22(.CP(n_62092), .D(n_13671), .CD(n_61408), .Q(addr_phys
		[22]));
	notech_reg addr_phys_reg_23(.CP(n_62096), .D(n_13672), .CD(n_61412), .Q(addr_phys
		[23]));
	notech_reg addr_phys_reg_24(.CP(n_62096), .D(n_13673), .CD(n_61412), .Q(addr_phys
		[24]));
	notech_reg addr_phys_reg_25(.CP(n_62096), .D(n_13674), .CD(n_61412), .Q(addr_phys
		[25]));
	notech_reg addr_phys_reg_26(.CP(n_62096), .D(n_13675), .CD(n_61412), .Q(addr_phys
		[26]));
	notech_reg addr_phys_reg_27(.CP(n_62096), .D(n_13676), .CD(n_61412), .Q(addr_phys
		[27]));
	notech_reg addr_phys_reg_28(.CP(n_62096), .D(n_13677), .CD(n_61412), .Q(addr_phys
		[28]));
	notech_reg addr_phys_reg_29(.CP(n_62096), .D(n_13678), .CD(n_61412), .Q(addr_phys
		[29]));
	notech_reg addr_phys_reg_30(.CP(n_62096), .D(n_13679), .CD(n_61412), .Q(addr_phys
		[30]));
	notech_reg addr_phys_reg_31(.CP(n_62096), .D(n_13680), .CD(n_61412), .Q(addr_phys
		[31]));
	notech_inv i_21458(.A(n_1052), .Z(n_13434));
	notech_inv i_21459(.A(n_1025), .Z(n_13435));
	notech_inv i_21460(.A(n_55449), .Z(n_13436));
	notech_inv i_21461(.A(n_999), .Z(n_13437));
	notech_inv i_21462(.A(n_985), .Z(n_13438));
	notech_inv i_21463(.A(n_1003), .Z(n_13439));
	notech_inv i_21464(.A(n_986), .Z(n_13440));
	notech_inv i_21465(.A(n_983), .Z(n_13441));
	notech_inv i_21466(.A(\nbus_14018[0] ), .Z(n_13442));
	notech_inv i_21467(.A(n_54355), .Z(n_13443));
	notech_inv i_21468(.A(fsm[1]), .Z(n_13444));
	notech_inv i_21469(.A(n_54361), .Z(n_13445));
	notech_inv i_21470(.A(fsm[2]), .Z(n_13446));
	notech_inv i_21471(.A(fsm[3]), .Z(n_13447));
	notech_inv i_21472(.A(n_494), .Z(n_13448));
	notech_inv i_21473(.A(\dir1[10] ), .Z(n_13449));
	notech_inv i_21474(.A(\dir1[11] ), .Z(n_13450));
	notech_inv i_21475(.A(\dir1[12] ), .Z(n_13451));
	notech_inv i_21476(.A(\dir1[13] ), .Z(n_13452));
	notech_inv i_21477(.A(\dir1[14] ), .Z(n_13453));
	notech_inv i_21478(.A(\dir1[15] ), .Z(n_13454));
	notech_inv i_21479(.A(\dir1[16] ), .Z(n_13455));
	notech_inv i_21480(.A(\dir1[17] ), .Z(n_13456));
	notech_inv i_21481(.A(\dir1[18] ), .Z(n_13457));
	notech_inv i_21482(.A(\dir1[19] ), .Z(n_13458));
	notech_inv i_21483(.A(\dir1[20] ), .Z(n_13459));
	notech_inv i_21484(.A(\dir1[21] ), .Z(n_13460));
	notech_inv i_21485(.A(\dir1[22] ), .Z(n_13461));
	notech_inv i_21486(.A(\dir1[23] ), .Z(n_13462));
	notech_inv i_21487(.A(\dir1[24] ), .Z(n_13463));
	notech_inv i_21488(.A(\dir1[25] ), .Z(n_13464));
	notech_inv i_21489(.A(\dir1[26] ), .Z(n_13465));
	notech_inv i_21490(.A(\dir1[27] ), .Z(n_13466));
	notech_inv i_21491(.A(\dir1[28] ), .Z(n_13467));
	notech_inv i_21492(.A(\dir1[29] ), .Z(n_13468));
	notech_inv i_21493(.A(n_536), .Z(n_13469));
	notech_inv i_21494(.A(n_54224), .Z(n_13470));
	notech_inv i_21495(.A(n_556), .Z(n_13471));
	notech_inv i_21496(.A(n_567), .Z(n_13472));
	notech_inv i_21497(.A(n_59313), .Z(n_13473));
	notech_inv i_21498(.A(\tab12[10] ), .Z(n_13474));
	notech_inv i_21499(.A(\tab12[11] ), .Z(n_13475));
	notech_inv i_21500(.A(\tab12[12] ), .Z(n_13476));
	notech_inv i_21501(.A(\tab12[13] ), .Z(n_13477));
	notech_inv i_21502(.A(\tab12[14] ), .Z(n_13478));
	notech_inv i_21503(.A(\tab12[15] ), .Z(n_13479));
	notech_inv i_21504(.A(\tab12[16] ), .Z(n_13480));
	notech_inv i_21505(.A(\tab12[17] ), .Z(n_13481));
	notech_inv i_21506(.A(\tab12[18] ), .Z(n_13482));
	notech_inv i_21507(.A(\tab12[19] ), .Z(n_13483));
	notech_inv i_21508(.A(\tab12[20] ), .Z(n_13484));
	notech_inv i_21509(.A(\tab12[21] ), .Z(n_13485));
	notech_inv i_21510(.A(\tab12[22] ), .Z(n_13486));
	notech_inv i_21511(.A(\tab12[23] ), .Z(n_13487));
	notech_inv i_21512(.A(\tab12[24] ), .Z(n_13488));
	notech_inv i_21513(.A(\tab12[25] ), .Z(n_13489));
	notech_inv i_21514(.A(\tab12[26] ), .Z(n_13490));
	notech_inv i_21515(.A(\tab12[27] ), .Z(n_13491));
	notech_inv i_21516(.A(\tab12[28] ), .Z(n_13492));
	notech_inv i_21517(.A(\tab12[29] ), .Z(n_13493));
	notech_inv i_21518(.A(hit_adr12), .Z(n_13494));
	notech_inv i_21519(.A(n_644), .Z(n_50854));
	notech_inv i_21520(.A(\tab14[10] ), .Z(n_13496));
	notech_inv i_21521(.A(\tab14[11] ), .Z(n_13497));
	notech_inv i_21522(.A(\tab14[12] ), .Z(n_13498));
	notech_inv i_21523(.A(\tab14[13] ), .Z(n_13499));
	notech_inv i_21524(.A(\tab14[14] ), .Z(n_13500));
	notech_inv i_21525(.A(\tab14[15] ), .Z(n_13501));
	notech_inv i_21526(.A(\tab14[16] ), .Z(n_13502));
	notech_inv i_21527(.A(\tab14[17] ), .Z(n_13503));
	notech_inv i_21528(.A(\tab14[18] ), .Z(n_13504));
	notech_inv i_21529(.A(\tab14[19] ), .Z(n_13505));
	notech_inv i_21530(.A(\tab14[20] ), .Z(n_13506));
	notech_inv i_21531(.A(\tab14[21] ), .Z(n_13507));
	notech_inv i_21532(.A(\tab14[22] ), .Z(n_13508));
	notech_inv i_21533(.A(\tab14[23] ), .Z(n_13509));
	notech_inv i_21534(.A(\tab14[24] ), .Z(n_13510));
	notech_inv i_21535(.A(\tab14[25] ), .Z(n_13511));
	notech_inv i_21536(.A(\tab14[26] ), .Z(n_13512));
	notech_inv i_21537(.A(\tab14[27] ), .Z(n_13513));
	notech_inv i_21538(.A(\tab14[28] ), .Z(n_13514));
	notech_inv i_21539(.A(\tab14[29] ), .Z(n_13515));
	notech_inv i_21540(.A(n_55041), .Z(n_13516));
	notech_inv i_21541(.A(\nx_tab1[0] ), .Z(n_13517));
	notech_inv i_21542(.A(n_55047), .Z(n_13518));
	notech_inv i_21543(.A(\nx_tab1[1] ), .Z(n_13519));
	notech_inv i_21544(.A(n_54299), .Z(n_13520));
	notech_inv i_21545(.A(\nnx_tab1[0] ), .Z(n_13521));
	notech_inv i_21546(.A(n_54305), .Z(n_13522));
	notech_inv i_21547(.A(\nnx_tab1[1] ), .Z(n_13523));
	notech_inv i_21548(.A(\nbus_14032[0] ), .Z(n_13524));
	notech_inv i_21549(.A(\tab22[10] ), .Z(n_13525));
	notech_inv i_21550(.A(\tab22[11] ), .Z(n_13526));
	notech_inv i_21551(.A(\tab22[12] ), .Z(n_13527));
	notech_inv i_21552(.A(\tab22[13] ), .Z(n_13528));
	notech_inv i_21553(.A(\tab22[14] ), .Z(n_13529));
	notech_inv i_21554(.A(\tab22[15] ), .Z(n_13530));
	notech_inv i_21555(.A(\tab22[16] ), .Z(n_13531));
	notech_inv i_21556(.A(\tab22[17] ), .Z(n_13532));
	notech_inv i_21557(.A(\tab22[18] ), .Z(n_13533));
	notech_inv i_21558(.A(\tab22[19] ), .Z(n_13534));
	notech_inv i_21559(.A(\tab22[20] ), .Z(n_13535));
	notech_inv i_21560(.A(\tab22[21] ), .Z(n_13536));
	notech_inv i_21561(.A(\tab22[22] ), .Z(n_13537));
	notech_inv i_21562(.A(\tab22[23] ), .Z(n_13538));
	notech_inv i_21563(.A(\tab22[24] ), .Z(n_13539));
	notech_inv i_21564(.A(\tab22[25] ), .Z(n_13540));
	notech_inv i_21565(.A(\tab22[26] ), .Z(n_13541));
	notech_inv i_21566(.A(\tab22[27] ), .Z(n_13542));
	notech_inv i_21567(.A(\tab22[28] ), .Z(n_13543));
	notech_inv i_21568(.A(\tab22[29] ), .Z(n_13544));
	notech_inv i_21569(.A(hit_adr22), .Z(n_13545));
	notech_inv i_21570(.A(\tab24[10] ), .Z(n_13546));
	notech_inv i_21571(.A(\tab24[11] ), .Z(n_13547));
	notech_inv i_21572(.A(\tab24[12] ), .Z(n_13548));
	notech_inv i_21573(.A(\tab24[13] ), .Z(n_13549));
	notech_inv i_21574(.A(\tab24[14] ), .Z(n_13550));
	notech_inv i_21575(.A(\tab24[15] ), .Z(n_13551));
	notech_inv i_21576(.A(\tab24[16] ), .Z(n_13552));
	notech_inv i_21577(.A(\tab24[17] ), .Z(n_13553));
	notech_inv i_21578(.A(\tab24[18] ), .Z(n_13554));
	notech_inv i_21579(.A(\tab24[19] ), .Z(n_13555));
	notech_inv i_21580(.A(\tab24[20] ), .Z(n_13556));
	notech_inv i_21581(.A(\tab24[21] ), .Z(n_13557));
	notech_inv i_21582(.A(\tab24[22] ), .Z(n_13558));
	notech_inv i_21583(.A(\tab24[23] ), .Z(n_13559));
	notech_inv i_21584(.A(\tab24[24] ), .Z(n_13560));
	notech_inv i_21585(.A(\tab24[25] ), .Z(n_13561));
	notech_inv i_21586(.A(\tab24[26] ), .Z(n_13562));
	notech_inv i_21587(.A(\tab24[27] ), .Z(n_13563));
	notech_inv i_21588(.A(\tab24[28] ), .Z(n_13564));
	notech_inv i_21589(.A(\tab24[29] ), .Z(n_13565));
	notech_inv i_21590(.A(n_54264), .Z(n_13566));
	notech_inv i_21591(.A(\nnx_tab2[0] ), .Z(n_13567));
	notech_inv i_21592(.A(n_54270), .Z(n_13568));
	notech_inv i_21593(.A(\nnx_tab2[1] ), .Z(n_13569));
	notech_inv i_21594(.A(\nbus_14031[0] ), .Z(n_13570));
	notech_inv i_21595(.A(n_55480), .Z(n_13571));
	notech_inv i_21596(.A(\nx_tab2[0] ), .Z(n_13572));
	notech_inv i_21597(.A(n_55486), .Z(n_13573));
	notech_inv i_21598(.A(\nx_tab2[1] ), .Z(n_13574));
	notech_inv i_21599(.A(\tab23[10] ), .Z(n_13575));
	notech_inv i_21600(.A(\tab23[11] ), .Z(n_13576));
	notech_inv i_21601(.A(\tab23[12] ), .Z(n_13577));
	notech_inv i_21602(.A(\tab23[13] ), .Z(n_13578));
	notech_inv i_21603(.A(\tab23[14] ), .Z(n_13579));
	notech_inv i_21604(.A(\tab23[15] ), .Z(n_13580));
	notech_inv i_21605(.A(\tab23[16] ), .Z(n_13581));
	notech_inv i_21606(.A(\tab23[17] ), .Z(n_13582));
	notech_inv i_21607(.A(\tab23[18] ), .Z(n_13583));
	notech_inv i_21608(.A(\tab23[19] ), .Z(n_13584));
	notech_inv i_21609(.A(\tab23[20] ), .Z(n_13585));
	notech_inv i_21610(.A(\tab23[21] ), .Z(n_13586));
	notech_inv i_21611(.A(\tab23[22] ), .Z(n_13587));
	notech_inv i_21612(.A(\tab23[23] ), .Z(n_13588));
	notech_inv i_21613(.A(\tab23[24] ), .Z(n_13589));
	notech_inv i_21614(.A(\tab23[25] ), .Z(n_13590));
	notech_inv i_21615(.A(\tab23[26] ), .Z(n_13591));
	notech_inv i_21616(.A(\tab23[27] ), .Z(n_13592));
	notech_inv i_21617(.A(\tab23[28] ), .Z(n_13593));
	notech_inv i_21618(.A(\tab23[29] ), .Z(n_13594));
	notech_inv i_21619(.A(n_52377), .Z(n_13595));
	notech_inv i_21620(.A(n_55095), .Z(n_13596));
	notech_inv i_21621(.A(n_55101), .Z(n_13597));
	notech_inv i_21622(.A(n_55107), .Z(n_13598));
	notech_inv i_21623(.A(n_55113), .Z(n_13599));
	notech_inv i_21624(.A(n_55119), .Z(n_13600));
	notech_inv i_21625(.A(n_55125), .Z(n_13601));
	notech_inv i_21626(.A(n_55131), .Z(n_13602));
	notech_inv i_21627(.A(n_55137), .Z(n_13603));
	notech_inv i_21628(.A(n_55143), .Z(n_13604));
	notech_inv i_21629(.A(n_55149), .Z(n_13605));
	notech_inv i_21630(.A(req_miss), .Z(n_13606));
	notech_inv i_21631(.A(addr_miss[0]), .Z(n_13607));
	notech_inv i_21632(.A(addr_miss[1]), .Z(n_13608));
	notech_inv i_21633(.A(addr_miss[2]), .Z(n_13609));
	notech_inv i_21634(.A(addr_miss[3]), .Z(n_13610));
	notech_inv i_21635(.A(addr_miss[4]), .Z(n_13611));
	notech_inv i_21636(.A(addr_miss[5]), .Z(n_13612));
	notech_inv i_21637(.A(addr_miss[6]), .Z(n_13613));
	notech_inv i_21638(.A(addr_miss[7]), .Z(n_13614));
	notech_inv i_21639(.A(addr_miss[8]), .Z(n_13615));
	notech_inv i_21640(.A(addr_miss[9]), .Z(n_13616));
	notech_inv i_21641(.A(n_950), .Z(n_13617));
	notech_inv i_21642(.A(addr_miss[10]), .Z(n_13618));
	notech_inv i_21643(.A(addr_miss[11]), .Z(n_13619));
	notech_inv i_21644(.A(addr_miss[12]), .Z(n_13620));
	notech_inv i_21645(.A(wrA[12]), .Z(n_13621));
	notech_inv i_21646(.A(addr_miss[13]), .Z(n_13622));
	notech_inv i_21647(.A(wrA[13]), .Z(n_13623));
	notech_inv i_21648(.A(addr_miss[14]), .Z(n_13624));
	notech_inv i_21649(.A(wrA[14]), .Z(n_13625));
	notech_inv i_21650(.A(addr_miss[15]), .Z(n_13626));
	notech_inv i_21651(.A(wrA[15]), .Z(n_13627));
	notech_inv i_21652(.A(addr_miss[16]), .Z(n_13628));
	notech_inv i_21653(.A(wrA[16]), .Z(n_13629));
	notech_inv i_21654(.A(addr_miss[17]), .Z(n_13630));
	notech_inv i_21655(.A(wrA[17]), .Z(n_13631));
	notech_inv i_21656(.A(addr_miss[18]), .Z(n_13632));
	notech_inv i_21657(.A(wrA[18]), .Z(n_13633));
	notech_inv i_21658(.A(addr_miss[19]), .Z(n_13634));
	notech_inv i_21659(.A(wrA[19]), .Z(n_13635));
	notech_inv i_21660(.A(addr_miss[20]), .Z(n_13636));
	notech_inv i_21661(.A(wrA[20]), .Z(n_13637));
	notech_inv i_21662(.A(addr_miss[21]), .Z(n_13638));
	notech_inv i_21663(.A(wrA[21]), .Z(n_13639));
	notech_inv i_21664(.A(addr_miss[22]), .Z(n_13640));
	notech_inv i_21665(.A(wrA[22]), .Z(n_13641));
	notech_inv i_21666(.A(addr_miss[23]), .Z(n_13642));
	notech_inv i_21667(.A(wrA[23]), .Z(n_13643));
	notech_inv i_21668(.A(addr_miss[24]), .Z(n_13644));
	notech_inv i_21669(.A(wrA[24]), .Z(n_13645));
	notech_inv i_21670(.A(addr_miss[25]), .Z(n_13646));
	notech_inv i_21671(.A(wrA[25]), .Z(n_13647));
	notech_inv i_21672(.A(addr_miss[26]), .Z(n_13648));
	notech_inv i_21673(.A(wrA[26]), .Z(n_13649));
	notech_inv i_21674(.A(addr_miss[27]), .Z(n_13650));
	notech_inv i_21675(.A(wrA[27]), .Z(n_13651));
	notech_inv i_21676(.A(addr_miss[28]), .Z(n_13652));
	notech_inv i_21677(.A(wrA[28]), .Z(n_13653));
	notech_inv i_21678(.A(addr_miss[29]), .Z(n_13654));
	notech_inv i_21679(.A(wrA[29]), .Z(n_13655));
	notech_inv i_21680(.A(addr_miss[30]), .Z(n_13656));
	notech_inv i_21681(.A(wrA[30]), .Z(n_13657));
	notech_inv i_21682(.A(addr_miss[31]), .Z(n_13658));
	notech_inv i_21683(.A(wrA[31]), .Z(n_13659));
	notech_inv i_21685(.A(n_53122), .Z(n_13661));
	notech_inv i_21686(.A(n_53129), .Z(n_13662));
	notech_inv i_21687(.A(n_53136), .Z(n_13663));
	notech_inv i_21688(.A(n_53143), .Z(n_13664));
	notech_inv i_21689(.A(n_53150), .Z(n_13665));
	notech_inv i_21690(.A(n_53157), .Z(n_13666));
	notech_inv i_21691(.A(n_53164), .Z(n_13667));
	notech_inv i_21692(.A(n_53171), .Z(n_13668));
	notech_inv i_21693(.A(n_53178), .Z(n_13669));
	notech_inv i_21694(.A(n_53185), .Z(n_13670));
	notech_inv i_21695(.A(n_53192), .Z(n_13671));
	notech_inv i_21696(.A(n_53199), .Z(n_13672));
	notech_inv i_21697(.A(n_53206), .Z(n_13673));
	notech_inv i_21698(.A(n_53213), .Z(n_13674));
	notech_inv i_21699(.A(n_53220), .Z(n_13675));
	notech_inv i_21700(.A(n_53227), .Z(n_13676));
	notech_inv i_21701(.A(n_53234), .Z(n_13677));
	notech_inv i_21702(.A(n_53241), .Z(n_13678));
	notech_inv i_21703(.A(n_53248), .Z(n_13679));
	notech_inv i_21704(.A(n_53255), .Z(n_13680));
	notech_inv i_21705(.A(cr3[31]), .Z(n_13681));
	notech_inv i_21706(.A(cr3[30]), .Z(n_13682));
	notech_inv i_21707(.A(cr3[29]), .Z(n_13683));
	notech_inv i_21708(.A(cr3[28]), .Z(n_13684));
	notech_inv i_21709(.A(cr3[27]), .Z(n_13685));
	notech_inv i_21710(.A(cr3[26]), .Z(n_13686));
	notech_inv i_21711(.A(cr3[25]), .Z(n_13687));
	notech_inv i_21712(.A(cr3[24]), .Z(n_13688));
	notech_inv i_21713(.A(cr3[23]), .Z(n_13689));
	notech_inv i_21714(.A(cr3[22]), .Z(n_13690));
	notech_inv i_21715(.A(cr3[21]), .Z(n_13691));
	notech_inv i_21716(.A(cr3[20]), .Z(n_13692));
	notech_inv i_21717(.A(cr3[19]), .Z(n_13693));
	notech_inv i_21718(.A(cr3[18]), .Z(n_13694));
	notech_inv i_21719(.A(cr3[17]), .Z(n_13695));
	notech_inv i_21720(.A(cr3[16]), .Z(n_13696));
	notech_inv i_21721(.A(cr3[15]), .Z(n_13697));
	notech_inv i_21722(.A(cr3[14]), .Z(n_13698));
	notech_inv i_21723(.A(cr3[13]), .Z(n_13699));
	notech_inv i_21724(.A(cr3[12]), .Z(n_13700));
	notech_inv i_21725(.A(iDaddr[0]), .Z(n_13701));
	notech_inv i_21726(.A(iDaddr[1]), .Z(n_13702));
	notech_inv i_21727(.A(iDaddr[2]), .Z(n_13703));
	notech_inv i_21728(.A(iDaddr[3]), .Z(n_13704));
	notech_inv i_21729(.A(iDaddr[4]), .Z(n_13705));
	notech_inv i_21730(.A(iDaddr[5]), .Z(n_13706));
	notech_inv i_21731(.A(iDaddr[6]), .Z(n_13707));
	notech_inv i_21732(.A(iDaddr[7]), .Z(n_13708));
	notech_inv i_21733(.A(iDaddr[8]), .Z(n_13709));
	notech_inv i_21734(.A(iDaddr[9]), .Z(n_13710));
	notech_inv i_21735(.A(iDaddr[10]), .Z(n_13711));
	notech_inv i_21736(.A(iDaddr[11]), .Z(n_13712));
	notech_inv i_21737(.A(iDaddr[12]), .Z(n_13713));
	notech_inv i_21738(.A(iDaddr[13]), .Z(n_13714));
	notech_inv i_21739(.A(iDaddr[14]), .Z(n_13715));
	notech_inv i_21740(.A(iDaddr[15]), .Z(n_13716));
	notech_inv i_21741(.A(iDaddr[16]), .Z(n_13717));
	notech_inv i_21742(.A(iDaddr[17]), .Z(n_13718));
	notech_inv i_21743(.A(iDaddr[18]), .Z(n_13719));
	notech_inv i_21744(.A(iDaddr[19]), .Z(n_13720));
	notech_inv i_21745(.A(iDaddr[20]), .Z(n_13721));
	notech_inv i_21746(.A(iDaddr[21]), .Z(n_13722));
	notech_inv i_21747(.A(iDaddr[22]), .Z(n_13723));
	notech_inv i_21748(.A(iDaddr[23]), .Z(n_13724));
	notech_inv i_21749(.A(iDaddr[24]), .Z(n_13725));
	notech_inv i_21750(.A(iDaddr[25]), .Z(n_13726));
	notech_inv i_21751(.A(iDaddr[26]), .Z(n_13727));
	notech_inv i_21752(.A(iDaddr[27]), .Z(n_13728));
	notech_inv i_21753(.A(iDaddr[28]), .Z(n_13729));
	notech_inv i_21754(.A(iDaddr[29]), .Z(n_13730));
	notech_inv i_21755(.A(iDaddr[30]), .Z(n_13731));
	notech_inv i_21756(.A(iDaddr[31]), .Z(n_13732));
	notech_inv i_21757(.A(cs[1]), .Z(n_13733));
	notech_inv i_21758(.A(cr0[16]), .Z(n_13734));
	notech_inv i_21759(.A(n_50878), .Z(n_13735));
	notech_inv i_21760(.A(n_50877), .Z(n_13736));
	notech_inv i_21761(.A(n_50876), .Z(n_13737));
	notech_inv i_21762(.A(n_50875), .Z(n_13738));
	notech_inv i_21763(.A(n_50874), .Z(n_13739));
	notech_inv i_21764(.A(n_50873), .Z(n_13740));
	notech_inv i_21765(.A(n_50872), .Z(n_13741));
	notech_inv i_21766(.A(n_50871), .Z(n_13742));
	notech_inv i_21767(.A(n_50870), .Z(n_13743));
	notech_inv i_21768(.A(n_50869), .Z(n_13744));
	notech_inv i_21769(.A(\addr_miss_0[11] ), .Z(n_13745));
	notech_inv i_21770(.A(\addr_miss_0[10] ), .Z(n_13746));
	notech_inv i_21771(.A(\addr_miss_0[9] ), .Z(n_13747));
	notech_inv i_21772(.A(\addr_miss_0[8] ), .Z(n_13748));
	notech_inv i_21773(.A(\addr_miss_0[7] ), .Z(n_13749));
	notech_inv i_21774(.A(\addr_miss_0[6] ), .Z(n_13750));
	notech_inv i_21775(.A(\addr_miss_0[5] ), .Z(n_13751));
	notech_inv i_21776(.A(\addr_miss_0[4] ), .Z(n_13752));
	notech_inv i_21777(.A(\addr_miss_0[3] ), .Z(n_13753));
	notech_inv i_21778(.A(\addr_miss_0[2] ), .Z(n_13754));
	notech_inv i_21779(.A(oread_ack100169), .Z(oread_ack));
	notech_inv i_21780(.A(hit_tab12), .Z(n_13756));
	notech_inv i_21781(.A(hit_tab23), .Z(n_13757));
	notech_inv i_21782(.A(hit_dir1), .Z(n_13758));
	notech_inv i_21783(.A(n_59304), .Z(n_13759));
	notech_inv i_21784(.A(n_61950), .Z(n_13760));
	notech_inv i_21785(.A(iread_ack), .Z(n_13761));
	cmp14_9 t23(.ina({\tab23[33] , \tab23[32] , UNCONNECTED_000, \tab23[30] 
		, \tab23[9] , \tab23[8] , \tab23[7] , \tab23[6] , \tab23[5] , \tab23[4] 
		, \tab23[3] , \tab23[2] , \tab23[1] , \tab23[0] }), .inb({
		UNCONNECTED_001, n_50854, UNCONNECTED_002, iwrite_req, \addr_miss_0[11] 
		, \addr_miss_0[10] , \addr_miss_0[9] , \addr_miss_0[8] , \addr_miss_0[7] 
		, \addr_miss_0[6] , \addr_miss_0[5] , \addr_miss_0[4] , \addr_miss_0[3] 
		, \addr_miss_0[2] }), .out(hit_tab23), .out2(hit_add23));
	cmp14_8 t11(.ina({\tab11[33] , \tab11[32] , UNCONNECTED_003, \tab11[30] 
		, \tab11[9] , \tab11[8] , \tab11[7] , \tab11[6] , \tab11[5] , \tab11[4] 
		, \tab11[3] , \tab11[2] , \tab11[1] , \tab11[0] }), .inb({
		UNCONNECTED_004, n_50854, UNCONNECTED_005, iwrite_req, \addr_miss_0[11] 
		, \addr_miss_0[10] , \addr_miss_0[9] , \addr_miss_0[8] , \addr_miss_0[7] 
		, \addr_miss_0[6] , \addr_miss_0[5] , \addr_miss_0[4] , \addr_miss_0[3] 
		, \addr_miss_0[2] }), .out(hit_tab11), .out2(hit_add11));
	cmp14_7 t24(.ina({\tab24[33] , \tab24[32] , UNCONNECTED_006, \tab24[30] 
		, \tab24[9] , \tab24[8] , \tab24[7] , \tab24[6] , \tab24[5] , \tab24[4] 
		, \tab24[3] , \tab24[2] , \tab24[1] , \tab24[0] }), .inb({
		UNCONNECTED_007, n_50854, UNCONNECTED_008, iwrite_req, \addr_miss_0[11] 
		, \addr_miss_0[10] , \addr_miss_0[9] , \addr_miss_0[8] , \addr_miss_0[7] 
		, \addr_miss_0[6] , \addr_miss_0[5] , \addr_miss_0[4] , \addr_miss_0[3] 
		, \addr_miss_0[2] }), .out(hit_tab24), .out2(hit_add24));
	cmp14_6 t22(.ina({\tab22[33] , \tab22[32] , UNCONNECTED_009, \tab22[30] 
		, \tab22[9] , \tab22[8] , \tab22[7] , \tab22[6] , \tab22[5] , \tab22[4] 
		, \tab22[3] , \tab22[2] , \tab22[1] , \tab22[0] }), .inb({
		UNCONNECTED_010, n_50854, UNCONNECTED_011, iwrite_req, \addr_miss_0[11] 
		, \addr_miss_0[10] , \addr_miss_0[9] , \addr_miss_0[8] , \addr_miss_0[7] 
		, \addr_miss_0[6] , \addr_miss_0[5] , \addr_miss_0[4] , \addr_miss_0[3] 
		, \addr_miss_0[2] }), .out(hit_tab22), .out2(hit_add22));
	cmp14_5 t21(.ina({\tab21[33] , \tab21[32] , UNCONNECTED_012, \tab21[30] 
		, \tab21[9] , \tab21[8] , \tab21[7] , \tab21[6] , \tab21[5] , \tab21[4] 
		, \tab21[3] , \tab21[2] , \tab21[1] , \tab21[0] }), .inb({
		UNCONNECTED_013, n_50854, UNCONNECTED_014, iwrite_req, \addr_miss_0[11] 
		, \addr_miss_0[10] , \addr_miss_0[9] , \addr_miss_0[8] , \addr_miss_0[7] 
		, \addr_miss_0[6] , \addr_miss_0[5] , \addr_miss_0[4] , \addr_miss_0[3] 
		, \addr_miss_0[2] }), .out(hit_tab21), .out2(hit_add21));
	cmp14_4 t14(.ina({\tab14[33] , \tab14[32] , UNCONNECTED_015, \tab14[30] 
		, \tab14[9] , \tab14[8] , \tab14[7] , \tab14[6] , \tab14[5] , \tab14[4] 
		, \tab14[3] , \tab14[2] , \tab14[1] , \tab14[0] }), .inb({
		UNCONNECTED_016, n_50854, UNCONNECTED_017, iwrite_req, \addr_miss_0[11] 
		, \addr_miss_0[10] , \addr_miss_0[9] , \addr_miss_0[8] , \addr_miss_0[7] 
		, \addr_miss_0[6] , \addr_miss_0[5] , \addr_miss_0[4] , \addr_miss_0[3] 
		, \addr_miss_0[2] }), .out(hit_tab14), .out2(hit_add14));
	cmp14_3 t13(.ina({\tab13[33] , \tab13[32] , UNCONNECTED_018, \tab13[30] 
		, \tab13[9] , \tab13[8] , \tab13[7] , \tab13[6] , \tab13[5] , \tab13[4] 
		, \tab13[3] , \tab13[2] , \tab13[1] , \tab13[0] }), .inb({
		UNCONNECTED_019, n_50854, UNCONNECTED_020, iwrite_req, \addr_miss_0[11] 
		, \addr_miss_0[10] , \addr_miss_0[9] , \addr_miss_0[8] , \addr_miss_0[7] 
		, \addr_miss_0[6] , \addr_miss_0[5] , \addr_miss_0[4] , \addr_miss_0[3] 
		, \addr_miss_0[2] }), .out(hit_tab13), .out2(hit_add13));
	cmp14_2 t12(.ina({\tab12[33] , \tab12[32] , UNCONNECTED_021, \tab12[30] 
		, \tab12[9] , \tab12[8] , \tab12[7] , \tab12[6] , \tab12[5] , \tab12[4] 
		, \tab12[3] , \tab12[2] , \tab12[1] , \tab12[0] }), .inb({
		UNCONNECTED_022, n_50854, UNCONNECTED_023, iwrite_req, \addr_miss_0[11] 
		, \addr_miss_0[10] , \addr_miss_0[9] , \addr_miss_0[8] , \addr_miss_0[7] 
		, \addr_miss_0[6] , \addr_miss_0[5] , \addr_miss_0[4] , \addr_miss_0[3] 
		, \addr_miss_0[2] }), .out(hit_tab12), .out2(hit_add12));
	cmp14_1 d2(.ina({\dir2[33] , UNCONNECTED_024, UNCONNECTED_025, 
		UNCONNECTED_026, \dir2[9] , \dir2[8] , \dir2[7] , \dir2[6] , \dir2[5] 
		, \dir2[4] , \dir2[3] , \dir2[2] , \dir2[1] , \dir2[0] }), .inb(
		{UNCONNECTED_027, UNCONNECTED_028, UNCONNECTED_029, 
		UNCONNECTED_030, n_50878, n_50877, n_50876, n_50875, n_50874, n_50873
		, n_50872, n_50871, n_50870, n_50869}), .out(hit_dir2));
	cmp14_0 d1(.ina({\dir1[33] , UNCONNECTED_031, UNCONNECTED_032, 
		UNCONNECTED_033, \dir1[9] , \dir1[8] , \dir1[7] , \dir1[6] , \dir1[5] 
		, \dir1[4] , \dir1[3] , \dir1[2] , \dir1[1] , \dir1[0] }), .inb(
		{UNCONNECTED_034, UNCONNECTED_035, UNCONNECTED_036, 
		UNCONNECTED_037, n_50878, n_50877, n_50876, n_50875, n_50874, n_50873
		, n_50872, n_50871, n_50870, n_50869}), .out(hit_dir1));
	AWDP_INC_10 i_75688(.O0(fsm5_cnt_0), .fsm5_cnt(fsm5_cnt));
endmodule
module AWDP_INC_26(O0, fsm5_cnt);

	output [8:0] O0;
	input [8:0] fsm5_cnt;




	notech_ha2 i_8(.A(fsm5_cnt[8]), .B(n_86), .Z(O0[8]));
	notech_ha2 i_7(.A(fsm5_cnt[7]), .B(n_84), .Z(O0[7]), .CO(n_86));
	notech_ha2 i_6(.A(fsm5_cnt[6]), .B(n_82), .Z(O0[6]), .CO(n_84));
	notech_ha2 i_5(.A(fsm5_cnt[5]), .B(n_80), .Z(O0[5]), .CO(n_82));
	notech_ha2 i_4(.A(fsm5_cnt[4]), .B(n_78), .Z(O0[4]), .CO(n_80));
	notech_ha2 i_3(.A(fsm5_cnt[3]), .B(n_76), .Z(O0[3]), .CO(n_78));
	notech_ha2 i_2(.A(fsm5_cnt[2]), .B(n_74), .Z(O0[2]), .CO(n_76));
	notech_ha2 i_1(.A(fsm5_cnt[1]), .B(fsm5_cnt[0]), .Z(O0[1]), .CO(n_74));
	notech_inv i_0(.A(fsm5_cnt[0]), .Z(O0[0]));
endmodule
module cmp14_10(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_10(.A(inb[2]), .B(ina[2]), .Z(n_34));
	notech_xor2 i_9(.A(inb[4]), .B(ina[4]), .Z(n_33));
	notech_xor2 i_8(.A(inb[6]), .B(ina[6]), .Z(n_32));
	notech_xor2 i_6(.A(inb[3]), .B(ina[3]), .Z(n_31));
	notech_xor2 i_5(.A(inb[5]), .B(ina[5]), .Z(n_30));
	notech_xor2 i_4(.A(inb[7]), .B(ina[7]), .Z(n_29));
	notech_xor2 i_0(.A(inb[9]), .B(ina[9]), .Z(n_55));
	notech_xor2 i_1(.A(inb[8]), .B(ina[8]), .Z(n_56));
	notech_xor2 i_3(.A(inb[1]), .B(ina[1]), .Z(n_57));
	notech_xor2 i_7(.A(inb[0]), .B(ina[0]), .Z(n_58));
	notech_or4 i_38(.A(n_57), .B(n_56), .C(n_55), .D(ina[13]), .Z(n_61));
	notech_or4 i_37(.A(n_34), .B(n_31), .C(n_33), .D(n_30), .Z(n_66));
	notech_or4 i_39(.A(n_32), .B(n_29), .C(n_58), .D(n_66), .Z(n_67));
	notech_nor2 i_2(.A(n_67), .B(n_61), .Z(out));
endmodule
module cmp14_11(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_10(.A(inb[2]), .B(ina[2]), .Z(n_34));
	notech_xor2 i_9(.A(inb[4]), .B(ina[4]), .Z(n_33));
	notech_xor2 i_8(.A(inb[6]), .B(ina[6]), .Z(n_32));
	notech_xor2 i_6(.A(inb[3]), .B(ina[3]), .Z(n_31));
	notech_xor2 i_5(.A(inb[5]), .B(ina[5]), .Z(n_30));
	notech_xor2 i_4(.A(inb[7]), .B(ina[7]), .Z(n_29));
	notech_xor2 i_0(.A(inb[9]), .B(ina[9]), .Z(n_55));
	notech_xor2 i_1(.A(inb[8]), .B(ina[8]), .Z(n_56));
	notech_xor2 i_3(.A(inb[1]), .B(ina[1]), .Z(n_57));
	notech_xor2 i_7(.A(inb[0]), .B(ina[0]), .Z(n_58));
	notech_or4 i_38(.A(n_57), .B(n_56), .C(n_55), .D(ina[13]), .Z(n_61));
	notech_or4 i_37(.A(n_34), .B(n_31), .C(n_33), .D(n_30), .Z(n_66));
	notech_or4 i_39(.A(n_32), .B(n_29), .C(n_58), .D(n_66), .Z(n_67));
	notech_nor2 i_2(.A(n_67), .B(n_61), .Z(out));
endmodule
module cmp14_12(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2100139), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2100139)
		);
	notech_inv i_9520(.A(out2100139), .Z(out2));
endmodule
module cmp14_13(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2100138), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2100138)
		);
	notech_inv i_9504(.A(out2100138), .Z(out2));
endmodule
module cmp14_14(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2100137), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2100137)
		);
	notech_inv i_9488(.A(out2100137), .Z(out2));
endmodule
module cmp14_15(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2100136), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2100136)
		);
	notech_inv i_9472(.A(out2100136), .Z(out2));
endmodule
module cmp14_16(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2100135), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2100135)
		);
	notech_inv i_9456(.A(out2100135), .Z(out2));
endmodule
module cmp14_17(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2100134), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2100134)
		);
	notech_inv i_9440(.A(out2100134), .Z(out2));
endmodule
module cmp14_18(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2100133), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2100133)
		);
	notech_inv i_9424(.A(out2100133), .Z(out2));
endmodule
module cmp14_19(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out2100132), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out2100132)
		);
	notech_inv i_9408(.A(out2100132), .Z(out2));
endmodule
module Itlb(clk, rstn, addr_phys, cr3, cr0, data_miss, iDaddr, pg_en, iwrite_data
		, owrite_data, iread_req, iread_ack, iwrite_req, iwrite_ack, iread_sz
		, oread_sz, oread_req, oread_ack, owrite_req, owrite_ack, pg_fault
		, wr_fault, cr2, flush_tlb, cs, pt_fault, busy_ram);

	input clk;
	input rstn;
	output [31:0] addr_phys;
	input [31:0] cr3;
	input [31:0] cr0;
	input [31:0] data_miss;
	input [31:0] iDaddr;
	input pg_en;
	input [31:0] iwrite_data;
	output [31:0] owrite_data;
	input iread_req;
	input iread_ack;
	input iwrite_req;
	input iwrite_ack;
	input [1:0] iread_sz;
	output [1:0] oread_sz;
	output oread_req;
	output oread_ack;
	output owrite_req;
	output owrite_ack;
	output pg_fault;
	output wr_fault;
	output [31:0] cr2;
	input flush_tlb;
	input [31:0] cs;
	output pt_fault;
	input busy_ram;

	wire [3:0] fsm;
	wire [31:0] iDaddr_f;
	wire [1:0] nx_dir;
	wire [8:0] fsm5_cnt_0;
	wire [8:0] fsm5_cnt;



	notech_inv i_15302(.A(n_62008), .Z(n_62062));
	notech_inv i_15301(.A(n_62008), .Z(n_62061));
	notech_inv i_15297(.A(n_62008), .Z(n_62057));
	notech_inv i_15293(.A(n_62008), .Z(n_62053));
	notech_inv i_15292(.A(n_62008), .Z(n_62052));
	notech_inv i_15288(.A(n_62008), .Z(n_62048));
	notech_inv i_15284(.A(n_62008), .Z(n_62044));
	notech_inv i_15283(.A(n_62008), .Z(n_62043));
	notech_inv i_15279(.A(n_62008), .Z(n_62039));
	notech_inv i_15274(.A(n_62008), .Z(n_62034));
	notech_inv i_15273(.A(n_62008), .Z(n_62033));
	notech_inv i_15269(.A(n_62008), .Z(n_62029));
	notech_inv i_15265(.A(n_62008), .Z(n_62025));
	notech_inv i_15264(.A(n_62008), .Z(n_62024));
	notech_inv i_15260(.A(n_62008), .Z(n_62020));
	notech_inv i_15256(.A(n_62008), .Z(n_62016));
	notech_inv i_15255(.A(n_62008), .Z(n_62015));
	notech_inv i_15251(.A(n_62008), .Z(n_62011));
	notech_inv i_15248(.A(clk), .Z(n_62008));
	notech_inv i_15246(.A(n_61980), .Z(n_62006));
	notech_inv i_15245(.A(n_61980), .Z(n_62005));
	notech_inv i_15241(.A(n_61980), .Z(n_62001));
	notech_inv i_15237(.A(n_61980), .Z(n_61997));
	notech_inv i_15236(.A(n_61980), .Z(n_61996));
	notech_inv i_15232(.A(n_61980), .Z(n_61992));
	notech_inv i_15228(.A(n_61980), .Z(n_61988));
	notech_inv i_15227(.A(n_61980), .Z(n_61987));
	notech_inv i_15223(.A(n_61980), .Z(n_61983));
	notech_inv i_15220(.A(clk), .Z(n_61980));
	notech_inv i_15186(.A(n_61936), .Z(n_61942));
	notech_inv i_15185(.A(n_61936), .Z(n_61941));
	notech_inv i_15181(.A(n_61936), .Z(n_61937));
	notech_inv i_15180(.A(pg_en), .Z(n_61936));
	notech_inv i_15176(.A(n_61925), .Z(n_61931));
	notech_inv i_15171(.A(n_61925), .Z(n_61926));
	notech_inv i_15170(.A(fsm[0]), .Z(n_61925));
	notech_inv i_15168(.A(n_61909), .Z(n_61922));
	notech_inv i_15166(.A(n_61909), .Z(n_61920));
	notech_inv i_15163(.A(n_61909), .Z(n_61917));
	notech_inv i_15161(.A(n_61909), .Z(n_61915));
	notech_inv i_15158(.A(n_61909), .Z(n_61912));
	notech_inv i_15156(.A(n_61909), .Z(n_61910));
	notech_inv i_15155(.A(n_551), .Z(n_61909));
	notech_inv i_15148(.A(n_61900), .Z(n_61901));
	notech_inv i_15147(.A(n_878), .Z(n_61900));
	notech_inv i_14795(.A(n_61847), .Z(n_61853));
	notech_inv i_14794(.A(n_61847), .Z(n_61852));
	notech_inv i_14790(.A(n_61847), .Z(n_61848));
	notech_inv i_14789(.A(n_886), .Z(n_61847));
	notech_inv i_14782(.A(n_61838), .Z(n_61839));
	notech_inv i_14781(.A(n_993), .Z(n_61838));
	notech_inv i_14774(.A(n_61829), .Z(n_61830));
	notech_inv i_14773(.A(n_9843), .Z(n_61829));
	notech_inv i_14297(.A(n_61293), .Z(n_61347));
	notech_inv i_14296(.A(n_61293), .Z(n_61346));
	notech_inv i_14292(.A(n_61293), .Z(n_61342));
	notech_inv i_14288(.A(n_61293), .Z(n_61338));
	notech_inv i_14287(.A(n_61293), .Z(n_61337));
	notech_inv i_14283(.A(n_61293), .Z(n_61333));
	notech_inv i_14279(.A(n_61293), .Z(n_61329));
	notech_inv i_14278(.A(n_61293), .Z(n_61328));
	notech_inv i_14274(.A(n_61293), .Z(n_61324));
	notech_inv i_14269(.A(n_61293), .Z(n_61319));
	notech_inv i_14268(.A(n_61293), .Z(n_61318));
	notech_inv i_14264(.A(n_61293), .Z(n_61314));
	notech_inv i_14260(.A(n_61293), .Z(n_61310));
	notech_inv i_14259(.A(n_61293), .Z(n_61309));
	notech_inv i_14255(.A(n_61293), .Z(n_61305));
	notech_inv i_14251(.A(n_61293), .Z(n_61301));
	notech_inv i_14250(.A(n_61293), .Z(n_61300));
	notech_inv i_14246(.A(n_61293), .Z(n_61296));
	notech_inv i_14243(.A(rstn), .Z(n_61293));
	notech_inv i_14241(.A(n_61265), .Z(n_61291));
	notech_inv i_14240(.A(n_61265), .Z(n_61290));
	notech_inv i_14236(.A(n_61265), .Z(n_61286));
	notech_inv i_14232(.A(n_61265), .Z(n_61282));
	notech_inv i_14231(.A(n_61265), .Z(n_61281));
	notech_inv i_14227(.A(n_61265), .Z(n_61277));
	notech_inv i_14223(.A(n_61265), .Z(n_61273));
	notech_inv i_14222(.A(n_61265), .Z(n_61272));
	notech_inv i_14218(.A(n_61265), .Z(n_61268));
	notech_inv i_14215(.A(rstn), .Z(n_61265));
	notech_inv i_14150(.A(n_61192), .Z(n_61193));
	notech_inv i_14149(.A(n_885), .Z(n_61192));
	notech_inv i_14142(.A(n_61183), .Z(n_61184));
	notech_inv i_14141(.A(n_890), .Z(n_61183));
	notech_inv i_13770(.A(n_60818), .Z(n_60819));
	notech_inv i_13769(.A(n_853), .Z(n_60818));
	notech_inv i_13766(.A(n_60809), .Z(n_60814));
	notech_inv i_13762(.A(n_60809), .Z(n_60810));
	notech_inv i_13761(.A(data_miss[0]), .Z(n_60809));
	notech_inv i_13577(.A(n_60524), .Z(n_60525));
	notech_inv i_13576(.A(\nbus_14490[0] ), .Z(n_60524));
	notech_inv i_13567(.A(n_60513), .Z(n_60514));
	notech_inv i_13566(.A(\nbus_14498[0] ), .Z(n_60513));
	notech_inv i_13557(.A(n_60502), .Z(n_60503));
	notech_inv i_13556(.A(\nbus_14491[0] ), .Z(n_60502));
	notech_inv i_13547(.A(n_60491), .Z(n_60492));
	notech_inv i_13546(.A(\nbus_14513[0] ), .Z(n_60491));
	notech_inv i_13537(.A(n_60480), .Z(n_60481));
	notech_inv i_13536(.A(\nbus_14502[0] ), .Z(n_60480));
	notech_inv i_13527(.A(n_60469), .Z(n_60470));
	notech_inv i_13526(.A(\nbus_14501[0] ), .Z(n_60469));
	notech_inv i_13517(.A(n_60458), .Z(n_60459));
	notech_inv i_13516(.A(\nbus_14500[0] ), .Z(n_60458));
	notech_inv i_13507(.A(n_60447), .Z(n_60448));
	notech_inv i_13506(.A(\nbus_14492[0] ), .Z(n_60447));
	notech_inv i_13497(.A(n_60436), .Z(n_60437));
	notech_inv i_13496(.A(\nbus_14503[0] ), .Z(n_60436));
	notech_inv i_13487(.A(n_60425), .Z(n_60426));
	notech_inv i_13486(.A(\nbus_14514[0] ), .Z(n_60425));
	notech_inv i_13464(.A(\nbus_14497[0] ), .Z(n_60401));
	notech_inv i_13459(.A(\nbus_14497[0] ), .Z(n_60396));
	notech_inv i_7872(.A(n_54439), .Z(n_54440));
	notech_inv i_7871(.A(n_808), .Z(n_54439));
	notech_xor2 i_77(.A(n_9961), .B(\nnx_tab1[0] ), .Z(n_490));
	notech_or4 i_72(.A(hit_adr13), .B(hit_adr14), .C(hit_adr12), .D(hit_adr11
		), .Z(n_488));
	notech_nand3 i_464(.A(\nx_tab2[0] ), .B(n_10012), .C(n_9844), .Z(n_484)
		);
	notech_nand3 i_463(.A(n_9844), .B(\nx_tab2[1] ), .C(n_10010), .Z(n_483)
		);
	notech_nand3 i_462(.A(n_9844), .B(\nx_tab2[1] ), .C(\nx_tab2[0] ), .Z(n_482
		));
	notech_xor2 i_78(.A(\nnx_tab2[1] ), .B(n_10005), .Z(n_478));
	notech_or4 i_73(.A(hit_adr23), .B(hit_adr24), .C(hit_adr22), .D(hit_adr21
		), .Z(n_476));
	notech_ao3 i_69(.A(n_10012), .B(n_9983), .C(hit_adr24), .Z(n_471));
	notech_nor2 i_66(.A(hit_adr24), .B(\nx_tab2[0] ), .Z(n_469));
	notech_nor2 i_452(.A(hit_adr23), .B(n_469), .Z(n_468));
	notech_nor2 i_79(.A(hit_adr22), .B(n_468), .Z(n_466));
	notech_or4 i_449(.A(n_899), .B(n_910), .C(\nx_tab1[1] ), .D(\nx_tab1[0] 
		), .Z(n_464));
	notech_and2 i_61(.A(fsm5_cnt[7]), .B(n_387), .Z(n_463));
	notech_or4 i_448(.A(fsm5_cnt[8]), .B(n_10158), .C(n_930), .D(n_463), .Z(n_462
		));
	notech_nor2 i_74(.A(n_463), .B(fsm5_cnt[8]), .Z(n_461));
	notech_nand2 i_445(.A(fsm[2]), .B(fsm[1]), .Z(n_459));
	notech_and3 i_51(.A(data_miss[5]), .B(iread_req), .C(n_60814), .Z(n_458)
		);
	notech_and2 i_82(.A(data_miss[5]), .B(n_60814), .Z(n_457));
	notech_ao3 i_85(.A(n_905), .B(iread_req), .C(busy_ram), .Z(n_454));
	notech_mux2 i_84(.S(fsm[3]), .A(n_459), .B(n_61931), .Z(n_453));
	notech_ao4 i_83(.A(n_61931), .B(n_889), .C(n_934), .D(n_896), .Z(n_452)
		);
	notech_or2 i_433(.A(iwrite_ack), .B(n_10035), .Z(n_450));
	notech_nor2 i_58(.A(data_miss[5]), .B(n_10101), .Z(n_449));
	notech_nand2 i_87(.A(n_948), .B(n_450), .Z(n_447));
	notech_mux2 i_86(.S(fsm[3]), .A(n_9845), .B(iwrite_ack), .Z(n_445));
	notech_nand3 i_427(.A(n_61931), .B(cr3[31]), .C(n_885), .Z(n_443));
	notech_nand3 i_424(.A(n_61931), .B(n_885), .C(cr3[30]), .Z(n_442));
	notech_nand3 i_421(.A(n_61931), .B(n_885), .C(cr3[29]), .Z(n_441));
	notech_nand3 i_418(.A(n_61931), .B(n_885), .C(cr3[28]), .Z(n_440));
	notech_nand3 i_415(.A(n_61931), .B(n_885), .C(cr3[27]), .Z(n_439));
	notech_nand3 i_412(.A(n_61931), .B(n_885), .C(cr3[26]), .Z(n_438));
	notech_nand3 i_409(.A(n_61931), .B(n_885), .C(cr3[25]), .Z(n_437));
	notech_nand3 i_406(.A(n_61931), .B(n_885), .C(cr3[24]), .Z(n_436));
	notech_nand3 i_403(.A(n_61931), .B(n_885), .C(cr3[23]), .Z(n_435));
	notech_nand3 i_400(.A(n_61931), .B(n_885), .C(cr3[22]), .Z(n_434));
	notech_nand3 i_397(.A(n_61931), .B(n_885), .C(cr3[21]), .Z(n_433));
	notech_nand3 i_394(.A(n_61931), .B(n_61193), .C(cr3[20]), .Z(n_432));
	notech_nand3 i_391(.A(n_61931), .B(n_61193), .C(cr3[19]), .Z(n_431));
	notech_nand3 i_388(.A(n_61931), .B(n_61193), .C(cr3[18]), .Z(n_430));
	notech_nand3 i_385(.A(n_61931), .B(n_61193), .C(cr3[17]), .Z(n_429));
	notech_nand3 i_382(.A(n_61931), .B(n_61193), .C(cr3[16]), .Z(n_428));
	notech_nand3 i_379(.A(n_61931), .B(n_61193), .C(cr3[15]), .Z(n_427));
	notech_nand3 i_376(.A(n_61926), .B(n_885), .C(cr3[14]), .Z(n_426));
	notech_nand3 i_373(.A(n_61926), .B(n_61193), .C(cr3[13]), .Z(n_425));
	notech_nand3 i_370(.A(n_61926), .B(n_61193), .C(cr3[12]), .Z(n_424));
	notech_nand3 i_344(.A(n_61941), .B(\wrA[2] ), .C(n_61853), .Z(n_400));
	notech_nor2 i_27(.A(n_972), .B(n_10158), .Z(n_399));
	notech_nand3 i_341(.A(n_61941), .B(n_61852), .C(\wrA[3] ), .Z(n_398));
	notech_nand3 i_338(.A(n_61942), .B(n_61853), .C(\wrA[4] ), .Z(n_397));
	notech_nand3 i_335(.A(n_61942), .B(n_61853), .C(\wrA[5] ), .Z(n_396));
	notech_nand3 i_332(.A(n_61942), .B(n_61853), .C(\wrA[6] ), .Z(n_395));
	notech_nand3 i_329(.A(n_61941), .B(n_61852), .C(\wrA[7] ), .Z(n_394));
	notech_nand3 i_326(.A(n_61941), .B(n_61852), .C(\wrA[8] ), .Z(n_393));
	notech_nand3 i_323(.A(n_61941), .B(n_61852), .C(\wrA[9] ), .Z(n_392));
	notech_nand3 i_320(.A(n_61941), .B(n_61852), .C(\wrA[10] ), .Z(n_391));
	notech_nand3 i_317(.A(n_61941), .B(n_61852), .C(\wrA[11] ), .Z(n_390));
	notech_nand2 i_81(.A(n_459), .B(n_10035), .Z(n_389));
	notech_nao3 i_21(.A(flush_tlb), .B(n_61942), .C(n_61920), .Z(n_388));
	notech_or2 i_60(.A(fsm5_cnt[6]), .B(n_386), .Z(n_387));
	notech_and3 i_52(.A(fsm5_cnt[4]), .B(fsm5_cnt[5]), .C(n_385), .Z(n_386)
		);
	notech_or2 i_48(.A(fsm5_cnt[2]), .B(fsm5_cnt[3]), .Z(n_385));
	notech_nor2 i_80(.A(hit_adr12), .B(n_497), .Z(n_495));
	notech_nor2 i_474(.A(hit_adr13), .B(n_498), .Z(n_497));
	notech_nor2 i_67(.A(hit_adr14), .B(\nx_tab1[0] ), .Z(n_498));
	notech_ao3 i_68(.A(n_9957), .B(n_9933), .C(hit_adr14), .Z(n_500));
	notech_or4 i_477(.A(n_899), .B(n_910), .C(n_9957), .D(n_9955), .Z(n_502)
		);
	notech_or4 i_478(.A(n_899), .B(n_910), .C(n_9957), .D(\nx_tab1[0] ), .Z(n_503
		));
	notech_or4 i_479(.A(n_899), .B(n_910), .C(n_9955), .D(\nx_tab1[1] ), .Z(n_504
		));
	notech_nand3 i_480(.A(n_60814), .B(n_875), .C(n_891), .Z(n_505));
	notech_nand3 i_483(.A(n_9844), .B(n_10012), .C(n_10010), .Z(n_508));
	notech_or2 i_484(.A(n_876), .B(n_875), .Z(n_509));
	notech_or4 i_503(.A(n_61926), .B(n_875), .C(n_889), .D(n_887), .Z(n_528)
		);
	notech_or4 i_506(.A(nx_dir[0]), .B(nx_dir[1]), .C(n_887), .D(n_890), .Z(n_531
		));
	notech_or4 i_507(.A(n_61926), .B(n_889), .C(n_887), .D(n_60814), .Z(n_532
		));
	notech_or4 i_829694(.A(fsm[1]), .B(fsm[3]), .C(fsm[2]), .D(n_61926), .Z(n_551
		));
	notech_nand2 i_47(.A(n_61942), .B(n_555), .Z(n_553));
	notech_or4 i_528(.A(fsm[2]), .B(n_884), .C(n_61926), .D(n_883), .Z(n_555
		));
	notech_or4 i_75(.A(hit_tab12), .B(hit_tab11), .C(hit_tab13), .D(hit_tab14
		), .Z(n_557));
	notech_or4 i_76(.A(hit_tab22), .B(hit_tab21), .C(hit_tab24), .D(hit_tab23
		), .Z(n_559));
	notech_nao3 i_96(.A(n_973), .B(\addr_miss[31] ), .C(n_61853), .Z(n_564)
		);
	notech_nao3 i_93(.A(n_994), .B(\tab22[29] ), .C(n_993), .Z(n_567));
	notech_nand3 i_90(.A(n_9843), .B(n_986), .C(\tab13[29] ), .Z(n_570));
	notech_nao3 i_107(.A(n_973), .B(\addr_miss[30] ), .C(n_61853), .Z(n_575)
		);
	notech_nao3 i_104(.A(n_994), .B(\tab22[28] ), .C(n_993), .Z(n_578));
	notech_nand3 i_101(.A(n_9843), .B(n_986), .C(\tab13[28] ), .Z(n_581));
	notech_nao3 i_118(.A(n_973), .B(\addr_miss[29] ), .C(n_61853), .Z(n_586)
		);
	notech_nao3 i_115(.A(n_994), .B(\tab22[27] ), .C(n_993), .Z(n_589));
	notech_nand3 i_112(.A(n_9843), .B(n_986), .C(\tab13[27] ), .Z(n_592));
	notech_nao3 i_129(.A(n_973), .B(\addr_miss[28] ), .C(n_61853), .Z(n_597)
		);
	notech_nao3 i_126(.A(n_994), .B(\tab22[26] ), .C(n_993), .Z(n_600));
	notech_nand3 i_123(.A(n_9843), .B(n_986), .C(\tab13[26] ), .Z(n_603));
	notech_nao3 i_140(.A(n_973), .B(\addr_miss[27] ), .C(n_61853), .Z(n_608)
		);
	notech_nao3 i_137(.A(n_994), .B(\tab22[25] ), .C(n_993), .Z(n_611));
	notech_nand3 i_134(.A(n_9843), .B(n_986), .C(\tab13[25] ), .Z(n_614));
	notech_nao3 i_151(.A(n_973), .B(\addr_miss[26] ), .C(n_61853), .Z(n_619)
		);
	notech_nao3 i_148(.A(n_994), .B(\tab22[24] ), .C(n_993), .Z(n_622));
	notech_nand3 i_145(.A(n_9843), .B(n_986), .C(\tab13[24] ), .Z(n_625));
	notech_nao3 i_162(.A(n_973), .B(\addr_miss[25] ), .C(n_61853), .Z(n_630)
		);
	notech_nao3 i_159(.A(n_994), .B(\tab22[23] ), .C(n_993), .Z(n_633));
	notech_nand3 i_156(.A(n_9843), .B(n_986), .C(\tab13[23] ), .Z(n_636));
	notech_nao3 i_173(.A(n_973), .B(\addr_miss[24] ), .C(n_61853), .Z(n_641)
		);
	notech_nao3 i_170(.A(n_994), .B(\tab22[22] ), .C(n_993), .Z(n_644));
	notech_nand3 i_167(.A(n_9843), .B(n_986), .C(\tab13[22] ), .Z(n_647));
	notech_nao3 i_184(.A(n_973), .B(\addr_miss[23] ), .C(n_61853), .Z(n_652)
		);
	notech_nao3 i_181(.A(n_994), .B(\tab22[21] ), .C(n_993), .Z(n_655));
	notech_nand3 i_178(.A(n_9843), .B(n_986), .C(\tab13[21] ), .Z(n_658));
	notech_nao3 i_195(.A(n_973), .B(\addr_miss[22] ), .C(n_61853), .Z(n_663)
		);
	notech_nao3 i_192(.A(n_994), .B(\tab22[20] ), .C(n_993), .Z(n_666));
	notech_nand3 i_189(.A(n_9843), .B(n_986), .C(\tab13[20] ), .Z(n_669));
	notech_nao3 i_206(.A(n_973), .B(\addr_miss[21] ), .C(n_61852), .Z(n_674)
		);
	notech_nao3 i_203(.A(n_994), .B(\tab22[19] ), .C(n_993), .Z(n_677));
	notech_nand3 i_200(.A(n_9843), .B(n_986), .C(\tab13[19] ), .Z(n_680));
	notech_nao3 i_219(.A(n_973), .B(\addr_miss[20] ), .C(n_61848), .Z(n_685)
		);
	notech_nao3 i_214(.A(n_994), .B(\tab22[18] ), .C(n_61839), .Z(n_688));
	notech_nand3 i_211(.A(n_61830), .B(n_986), .C(\tab13[18] ), .Z(n_691));
	notech_nao3 i_235(.A(n_973), .B(\addr_miss[19] ), .C(n_61848), .Z(n_696)
		);
	notech_nao3 i_232(.A(n_994), .B(\tab22[17] ), .C(n_61839), .Z(n_699));
	notech_nand3 i_229(.A(n_61830), .B(n_986), .C(\tab13[17] ), .Z(n_702));
	notech_nao3 i_246(.A(n_973), .B(\addr_miss[18] ), .C(n_61848), .Z(n_707)
		);
	notech_nao3 i_243(.A(n_994), .B(\tab22[16] ), .C(n_61839), .Z(n_710));
	notech_nand3 i_240(.A(n_61830), .B(n_986), .C(\tab13[16] ), .Z(n_713));
	notech_nao3 i_257(.A(n_973), .B(\addr_miss[17] ), .C(n_61848), .Z(n_718)
		);
	notech_nao3 i_254(.A(n_994), .B(\tab22[15] ), .C(n_61839), .Z(n_721));
	notech_nand3 i_251(.A(n_61830), .B(n_986), .C(\tab13[15] ), .Z(n_724));
	notech_nao3 i_268(.A(n_973), .B(\addr_miss[16] ), .C(n_61848), .Z(n_729)
		);
	notech_nao3 i_265(.A(n_994), .B(\tab22[14] ), .C(n_61839), .Z(n_732));
	notech_nand3 i_262(.A(n_61830), .B(n_986), .C(\tab13[14] ), .Z(n_735));
	notech_nao3 i_279(.A(n_973), .B(\addr_miss[15] ), .C(n_61848), .Z(n_740)
		);
	notech_nao3 i_276(.A(n_994), .B(\tab22[13] ), .C(n_61839), .Z(n_743));
	notech_nand3 i_273(.A(n_61830), .B(n_986), .C(\tab13[13] ), .Z(n_746));
	notech_nao3 i_290(.A(n_973), .B(\addr_miss[14] ), .C(n_61848), .Z(n_751)
		);
	notech_nao3 i_287(.A(n_994), .B(\tab22[12] ), .C(n_61839), .Z(n_754));
	notech_nand3 i_284(.A(n_61830), .B(n_986), .C(\tab13[12] ), .Z(n_757));
	notech_nao3 i_301(.A(n_973), .B(\addr_miss[13] ), .C(n_61848), .Z(n_762)
		);
	notech_nao3 i_298(.A(n_994), .B(\tab22[11] ), .C(n_993), .Z(n_765));
	notech_nand3 i_295(.A(n_9843), .B(n_986), .C(\tab13[11] ), .Z(n_768));
	notech_nao3 i_312(.A(\addr_miss[12] ), .B(n_973), .C(n_61848), .Z(n_773)
		);
	notech_nao3 i_309(.A(\tab22[10] ), .B(n_994), .C(n_61839), .Z(n_776));
	notech_nand3 i_306(.A(n_61830), .B(\tab13[10] ), .C(n_986), .Z(n_779));
	notech_and2 i_8(.A(\wrD[7] ), .B(n_61848), .Z(owrite_data[7]));
	notech_and2 i_7(.A(\wrD[6] ), .B(n_61852), .Z(owrite_data[6]));
	notech_and2 i_6(.A(\wrD[5] ), .B(n_61852), .Z(owrite_data[5]));
	notech_and2 i_522313(.A(\wrD[4] ), .B(n_61852), .Z(owrite_data[4]));
	notech_and2 i_4(.A(\wrD[3] ), .B(n_61852), .Z(owrite_data[3]));
	notech_and2 i_3(.A(\wrD[2] ), .B(n_61852), .Z(owrite_data[2]));
	notech_and2 i_222312(.A(\wrD[1] ), .B(n_61848), .Z(owrite_data[1]));
	notech_and2 i_1(.A(\wrD[0] ), .B(n_61848), .Z(owrite_data[0]));
	notech_nao3 i_80198(.A(n_58203), .B(n_10101), .C(n_887), .Z(n_808));
	notech_or4 i_434(.A(n_854), .B(flush_tlb), .C(n_893), .D(n_906), .Z(n_851
		));
	notech_or4 i_435(.A(fsm[2]), .B(fsm[1]), .C(n_10158), .D(n_10035), .Z(n_852
		));
	notech_nand2 i_81549(.A(n_61942), .B(n_58109), .Z(n_853));
	notech_ao4 i_49(.A(hit_dir2), .B(\hit_dir1[7] ), .C(pg_fault), .D(n_9847
		), .Z(n_854));
	notech_or4 i_439(.A(fsm[1]), .B(fsm[3]), .C(fsm[2]), .D(n_454), .Z(n_855
		));
	notech_nao3 i_444(.A(n_10035), .B(n_9845), .C(iwrite_ack), .Z(n_858));
	notech_and2 i_44(.A(iwrite_ack), .B(n_389), .Z(n_861));
	notech_and2 i_79451(.A(n_58203), .B(n_10101), .Z(n_862));
	notech_ao3 i_79439(.A(fsm5_cnt_0[0]), .B(n_929), .C(n_884), .Z(n_863));
	notech_ao3 i_79440(.A(n_929), .B(fsm5_cnt_0[1]), .C(n_884), .Z(n_864));
	notech_ao3 i_79441(.A(n_929), .B(fsm5_cnt_0[2]), .C(n_884), .Z(n_865));
	notech_ao3 i_79442(.A(n_929), .B(fsm5_cnt_0[3]), .C(n_884), .Z(n_866));
	notech_ao3 i_79443(.A(n_929), .B(fsm5_cnt_0[4]), .C(n_884), .Z(n_867));
	notech_ao3 i_79444(.A(n_929), .B(fsm5_cnt_0[5]), .C(n_884), .Z(n_868));
	notech_ao3 i_79445(.A(n_929), .B(fsm5_cnt_0[6]), .C(n_884), .Z(n_869));
	notech_ao3 i_79446(.A(n_929), .B(fsm5_cnt_0[7]), .C(n_884), .Z(n_870));
	notech_ao3 i_79447(.A(n_929), .B(fsm5_cnt_0[8]), .C(n_884), .Z(n_871));
	notech_or4 i_80182(.A(n_906), .B(n_893), .C(n_904), .D(n_905), .Z(n_872)
		);
	notech_nor2 i_80085(.A(n_896), .B(n_10148), .Z(n_873));
	notech_ao3 i_79278(.A(n_60814), .B(\dir1_0[4] ), .C(n_890), .Z(n_874));
	notech_nor2 i_329692(.A(nx_dir[0]), .B(nx_dir[1]), .Z(n_875));
	notech_or4 i_80843(.A(n_61926), .B(n_889), .C(n_887), .D(n_10101), .Z(n_876
		));
	notech_and2 i_79195(.A(iread_ack), .B(n_553), .Z(oread_ack));
	notech_reg nx_dir_reg_0(.CP(n_62039), .D(n_6993), .CD(n_61324), .Q(nx_dir
		[0]));
	notech_mux2 i_9554(.S(n_876), .A(n_875), .B(nx_dir[0]), .Z(n_6993));
	notech_nand3 i_79167(.A(n_10035), .B(n_9845), .C(n_61942), .Z(n_878));
	notech_reg nx_dir_reg_1(.CP(n_62039), .D(n_7002), .CD(n_61324), .Q(nx_dir
		[1]));
	notech_and2 i_9564(.A(n_876), .B(nx_dir[1]), .Z(n_7002));
	notech_reg iDaddr_f_reg_0(.CP(n_62039), .D(n_7005), .CD(n_61324), .Q(iDaddr_f
		[0]));
	notech_mux2 i_9570(.S(n_61920), .A(iDaddr[0]), .B(iDaddr_f[0]), .Z(n_7005
		));
	notech_reg iDaddr_f_reg_1(.CP(n_62039), .D(n_7011), .CD(n_61324), .Q(iDaddr_f
		[1]));
	notech_mux2 i_9578(.S(n_61920), .A(iDaddr[1]), .B(iDaddr_f[1]), .Z(n_7011
		));
	notech_reg iDaddr_f_reg_2(.CP(n_62034), .D(n_7017), .CD(n_61319), .Q(iDaddr_f
		[2]));
	notech_mux2 i_9586(.S(n_61917), .A(iDaddr[2]), .B(iDaddr_f[2]), .Z(n_7017
		));
	notech_reg iDaddr_f_reg_3(.CP(n_62039), .D(n_7023), .CD(n_61324), .Q(iDaddr_f
		[3]));
	notech_mux2 i_9594(.S(n_61917), .A(iDaddr[3]), .B(iDaddr_f[3]), .Z(n_7023
		));
	notech_ao4 i_79025(.A(n_10160), .B(n_9932), .C(n_10157), .D(n_9931), .Z(n_883
		));
	notech_reg iDaddr_f_reg_4(.CP(n_62039), .D(n_7029), .CD(n_61324), .Q(iDaddr_f
		[4]));
	notech_mux2 i_9602(.S(n_61920), .A(iDaddr[4]), .B(iDaddr_f[4]), .Z(n_7029
		));
	notech_or2 i_30(.A(fsm[1]), .B(fsm[3]), .Z(n_884));
	notech_reg iDaddr_f_reg_5(.CP(n_62039), .D(n_7035), .CD(n_61324), .Q(iDaddr_f
		[5]));
	notech_mux2 i_9610(.S(n_61920), .A(iDaddr[5]), .B(iDaddr_f[5]), .Z(n_7035
		));
	notech_nor2 i_59(.A(fsm[2]), .B(n_884), .Z(n_885));
	notech_reg iDaddr_f_reg_6(.CP(n_62039), .D(n_7041), .CD(n_61324), .Q(iDaddr_f
		[6]));
	notech_mux2 i_9618(.S(n_61920), .A(iDaddr[6]), .B(iDaddr_f[6]), .Z(n_7041
		));
	notech_and3 i_20(.A(fsm[2]), .B(fsm[1]), .C(n_10035), .Z(n_886));
	notech_reg iDaddr_f_reg_7(.CP(n_62039), .D(n_7047), .CD(n_61324), .Q(iDaddr_f
		[7]));
	notech_mux2 i_9626(.S(n_61920), .A(iDaddr[7]), .B(iDaddr_f[7]), .Z(n_7047
		));
	notech_nand2 i_31(.A(iread_ack), .B(n_61942), .Z(n_887));
	notech_reg iDaddr_f_reg_8(.CP(n_62039), .D(n_7053), .CD(n_61324), .Q(iDaddr_f
		[8]));
	notech_mux2 i_9634(.S(n_61920), .A(iDaddr[8]), .B(iDaddr_f[8]), .Z(n_7053
		));
	notech_reg iDaddr_f_reg_9(.CP(n_62039), .D(n_7059), .CD(n_61324), .Q(iDaddr_f
		[9]));
	notech_mux2 i_9642(.S(n_61920), .A(iDaddr[9]), .B(iDaddr_f[9]), .Z(n_7059
		));
	notech_nao3 i_18(.A(fsm[1]), .B(n_10035), .C(fsm[2]), .Z(n_889));
	notech_reg iDaddr_f_reg_10(.CP(n_62039), .D(n_7065), .CD(n_61324), .Q(iDaddr_f
		[10]));
	notech_mux2 i_9650(.S(n_61917), .A(iDaddr[10]), .B(iDaddr_f[10]), .Z(n_7065
		));
	notech_nand2 i_32(.A(n_10034), .B(n_9846), .Z(n_890));
	notech_reg iDaddr_f_reg_11(.CP(n_62039), .D(n_7071), .CD(n_61324), .Q(iDaddr_f
		[11]));
	notech_mux2 i_9658(.S(n_61917), .A(iDaddr[11]), .B(iDaddr_f[11]), .Z(n_7071
		));
	notech_ao3 i_55(.A(iread_ack), .B(n_61942), .C(n_890), .Z(n_891));
	notech_reg iDaddr_f_reg_12(.CP(n_62034), .D(\tab11_0[0] ), .CD(n_61319),
		 .Q(iDaddr_f[12]));
	notech_reg iDaddr_f_reg_13(.CP(n_62034), .D(\tab11_0[1] ), .CD(n_61319),
		 .Q(iDaddr_f[13]));
	notech_or4 i_64(.A(fsm[2]), .B(n_884), .C(n_61926), .D(n_10158), .Z(n_893
		));
	notech_reg iDaddr_f_reg_14(.CP(n_62034), .D(\tab11_0[2] ), .CD(n_61319),
		 .Q(iDaddr_f[14]));
	notech_reg iDaddr_f_reg_15(.CP(n_62034), .D(\tab11_0[3] ), .CD(n_61319),
		 .Q(iDaddr_f[15]));
	notech_nand2 i_802(.A(fsm[2]), .B(n_10034), .Z(n_895));
	notech_reg iDaddr_f_reg_16(.CP(n_62034), .D(\tab11_0[4] ), .CD(n_61319),
		 .Q(iDaddr_f[16]));
	notech_or2 i_79143(.A(n_884), .B(n_895), .Z(n_896));
	notech_reg iDaddr_f_reg_17(.CP(n_62034), .D(\tab11_0[5] ), .CD(n_61319),
		 .Q(iDaddr_f[17]));
	notech_reg iDaddr_f_reg_18(.CP(n_62034), .D(\tab11_0[6] ), .CD(n_61319),
		 .Q(iDaddr_f[18]));
	notech_reg iDaddr_f_reg_19(.CP(n_62034), .D(\tab11_0[7] ), .CD(n_61319),
		 .Q(iDaddr_f[19]));
	notech_or4 i_10(.A(n_887), .B(n_884), .C(n_895), .D(n_10101), .Z(n_899)
		);
	notech_reg iDaddr_f_reg_20(.CP(n_62034), .D(\tab11_0[8] ), .CD(n_61319),
		 .Q(iDaddr_f[20]));
	notech_nand2 i_19(.A(hit_dir2), .B(n_10157), .Z(n_900));
	notech_reg iDaddr_f_reg_21(.CP(n_62034), .D(\tab11_0[9] ), .CD(n_61319),
		 .Q(iDaddr_f[21]));
	notech_or4 i_33(.A(n_896), .B(n_887), .C(n_900), .D(n_10101), .Z(n_901)
		);
	notech_reg iDaddr_f_reg_22(.CP(n_62034), .D(\dir1_0[0] ), .CD(n_61319), 
		.Q(iDaddr_f[22]));
	notech_reg iDaddr_f_reg_23(.CP(n_62034), .D(\dir1_0[1] ), .CD(n_61319), 
		.Q(iDaddr_f[23]));
	notech_reg iDaddr_f_reg_24(.CP(n_62034), .D(\dir1_0[2] ), .CD(n_61319), 
		.Q(iDaddr_f[24]));
	notech_nao3 i_798(.A(n_883), .B(n_10161), .C(flush_tlb), .Z(n_904));
	notech_reg iDaddr_f_reg_25(.CP(n_62034), .D(\dir1_0[3] ), .CD(n_61319), 
		.Q(iDaddr_f[25]));
	notech_and2 i_26(.A(n_10160), .B(n_10157), .Z(n_905));
	notech_reg iDaddr_f_reg_26(.CP(n_62034), .D(\dir1_0[4] ), .CD(n_61319), 
		.Q(iDaddr_f[26]));
	notech_or2 i_45(.A(busy_ram), .B(n_10159), .Z(n_906));
	notech_reg iDaddr_f_reg_27(.CP(n_62039), .D(\dir1_0[5] ), .CD(n_61324), 
		.Q(iDaddr_f[27]));
	notech_reg iDaddr_f_reg_28(.CP(n_62043), .D(\dir1_0[6] ), .CD(n_61328), 
		.Q(iDaddr_f[28]));
	notech_reg iDaddr_f_reg_29(.CP(n_62043), .D(\dir1_0[7] ), .CD(n_61328), 
		.Q(iDaddr_f[29]));
	notech_reg iDaddr_f_reg_30(.CP(n_62043), .D(\dir1_0[8] ), .CD(n_61328), 
		.Q(iDaddr_f[30]));
	notech_nand2 i_17(.A(\hit_dir1[7] ), .B(n_10160), .Z(n_910));
	notech_reg iDaddr_f_reg_31(.CP(n_62043), .D(\dir1_0[9] ), .CD(n_61328), 
		.Q(iDaddr_f[31]));
	notech_or4 i_34(.A(n_896), .B(n_887), .C(n_910), .D(n_10101), .Z(n_911)
		);
	notech_reg_set dir1_reg_0(.CP(n_62043), .D(n_7197), .SD(n_61328), .Q(\dir1[0] 
		));
	notech_mux2 i_9826(.S(\nbus_14501[0] ), .A(\dir1[0] ), .B(n_57422), .Z(n_7197
		));
	notech_reg_set dir1_reg_1(.CP(n_62043), .D(n_7203), .SD(n_61328), .Q(\dir1[1] 
		));
	notech_mux2 i_9834(.S(\nbus_14501[0] ), .A(\dir1[1] ), .B(n_57428), .Z(n_7203
		));
	notech_reg_set dir1_reg_2(.CP(n_62043), .D(n_7209), .SD(n_61328), .Q(\dir1[2] 
		));
	notech_mux2 i_9842(.S(\nbus_14501[0] ), .A(\dir1[2] ), .B(n_57434), .Z(n_7209
		));
	notech_reg_set dir1_reg_3(.CP(n_62044), .D(n_7215), .SD(n_61329), .Q(\dir1[3] 
		));
	notech_mux2 i_9850(.S(\nbus_14501[0] ), .A(\dir1[3] ), .B(n_57440), .Z(n_7215
		));
	notech_reg dir1_reg_4(.CP(n_62044), .D(n_7221), .CD(n_61329), .Q(\dir1[4] 
		));
	notech_mux2 i_9858(.S(\nbus_14501[0] ), .A(\dir1[4] ), .B(n_874), .Z(n_7221
		));
	notech_nand2 i_79139(.A(n_61926), .B(n_9846), .Z(n_916));
	notech_reg_set dir1_reg_5(.CP(n_62044), .D(n_7227), .SD(n_61329), .Q(\dir1[5] 
		));
	notech_mux2 i_9866(.S(\nbus_14501[0] ), .A(\dir1[5] ), .B(n_57452), .Z(n_7227
		));
	notech_or2 i_53(.A(n_916), .B(hit_adr11), .Z(n_917));
	notech_reg_set dir1_reg_6(.CP(n_62044), .D(n_7233), .SD(n_61329), .Q(\dir1[6] 
		));
	notech_mux2 i_9874(.S(\nbus_14501[0] ), .A(\dir1[6] ), .B(n_57458), .Z(n_7233
		));
	notech_or2 i_790(.A(hit_adr12), .B(n_917), .Z(n_918));
	notech_reg_set dir1_reg_7(.CP(n_62044), .D(n_7239), .SD(n_61329), .Q(\dir1[7] 
		));
	notech_mux2 i_9882(.S(\nbus_14501[0] ), .A(\dir1[7] ), .B(n_57464), .Z(n_7239
		));
	notech_nao3 i_29(.A(n_61926), .B(n_61942), .C(n_889), .Z(n_919));
	notech_reg_set dir1_reg_8(.CP(n_62044), .D(n_7245), .SD(n_61329), .Q(\dir1[8] 
		));
	notech_mux2 i_9890(.S(\nbus_14501[0] ), .A(\dir1[8] ), .B(n_57470), .Z(n_7245
		));
	notech_reg_set dir1_reg_9(.CP(n_62044), .D(n_7251), .SD(n_61329), .Q(\dir1[9] 
		));
	notech_mux2 i_9898(.S(\nbus_14501[0] ), .A(\dir1[9] ), .B(n_57476), .Z(n_7251
		));
	notech_reg_set dir1_reg_10(.CP(n_62043), .D(n_7257), .SD(n_61328), .Q(\dir1[10] 
		));
	notech_mux2 i_9906(.S(\nbus_14501[0] ), .A(\dir1[10] ), .B(n_57482), .Z(n_7257
		));
	notech_reg_set dir1_reg_11(.CP(n_62043), .D(n_7263), .SD(n_61328), .Q(\dir1[11] 
		));
	notech_mux2 i_9914(.S(\nbus_14501[0] ), .A(\dir1[11] ), .B(n_57488), .Z(n_7263
		));
	notech_reg_set dir1_reg_12(.CP(n_62043), .D(n_7269), .SD(n_61328), .Q(\dir1[12] 
		));
	notech_mux2 i_9922(.S(\nbus_14501[0] ), .A(\dir1[12] ), .B(n_57494), .Z(n_7269
		));
	notech_reg_set dir1_reg_13(.CP(n_62043), .D(n_7275), .SD(n_61328), .Q(\dir1[13] 
		));
	notech_mux2 i_9930(.S(\nbus_14501[0] ), .A(\dir1[13] ), .B(n_57500), .Z(n_7275
		));
	notech_reg_set dir1_reg_14(.CP(n_62039), .D(n_7281), .SD(n_61324), .Q(\dir1[14] 
		));
	notech_mux2 i_9938(.S(\nbus_14501[0] ), .A(\dir1[14] ), .B(n_57506), .Z(n_7281
		));
	notech_or2 i_54(.A(n_916), .B(hit_adr21), .Z(n_926));
	notech_reg_set dir1_reg_15(.CP(n_62039), .D(n_7287), .SD(n_61324), .Q(\dir1[15] 
		));
	notech_mux2 i_9946(.S(\nbus_14501[0] ), .A(\dir1[15] ), .B(n_57512), .Z(n_7287
		));
	notech_or2 i_784(.A(hit_adr22), .B(n_926), .Z(n_927));
	notech_reg_set dir1_reg_16(.CP(n_62039), .D(n_7293), .SD(n_61324), .Q(\dir1[16] 
		));
	notech_mux2 i_9954(.S(n_60470), .A(\dir1[16] ), .B(n_57518), .Z(n_7293)
		);
	notech_reg_set dir1_reg_17(.CP(n_62039), .D(n_7299), .SD(n_61324), .Q(\dir1[17] 
		));
	notech_mux2 i_9962(.S(n_60470), .A(\dir1[17] ), .B(n_57524), .Z(n_7299)
		);
	notech_and2 i_782(.A(fsm[2]), .B(n_61931), .Z(n_929));
	notech_reg_set dir1_reg_18(.CP(n_62043), .D(n_7305), .SD(n_61328), .Q(\dir1[18] 
		));
	notech_mux2 i_9970(.S(n_60470), .A(\dir1[18] ), .B(n_57530), .Z(n_7305)
		);
	notech_nao3 i_79146(.A(fsm[2]), .B(n_61926), .C(n_884), .Z(n_930));
	notech_reg_set dir1_reg_19(.CP(n_62043), .D(n_7311), .SD(n_61328), .Q(\dir1[19] 
		));
	notech_mux2 i_9978(.S(n_60470), .A(\dir1[19] ), .B(n_57536), .Z(n_7311)
		);
	notech_reg_set dir1_reg_20(.CP(n_62043), .D(n_7317), .SD(n_61328), .Q(\dir1[20] 
		));
	notech_mux2 i_9986(.S(n_60470), .A(\dir1[20] ), .B(n_57542), .Z(n_7317)
		);
	notech_nao3 i_35(.A(n_929), .B(n_61942), .C(n_884), .Z(n_932));
	notech_reg_set dir1_reg_21(.CP(n_62043), .D(n_7323), .SD(n_61328), .Q(\dir1[21] 
		));
	notech_mux2 i_9994(.S(n_60470), .A(\dir1[21] ), .B(n_57548), .Z(n_7323)
		);
	notech_reg_set dir1_reg_22(.CP(n_62043), .D(n_7329), .SD(n_61328), .Q(\dir1[22] 
		));
	notech_mux2 i_10002(.S(n_60470), .A(\dir1[22] ), .B(n_57554), .Z(n_7329)
		);
	notech_and2 i_28(.A(data_miss[5]), .B(iread_req), .Z(n_934));
	notech_reg_set dir1_reg_23(.CP(n_62043), .D(n_7335), .SD(n_61328), .Q(\dir1[23] 
		));
	notech_mux2 i_10010(.S(n_60470), .A(\dir1[23] ), .B(n_57560), .Z(n_7335)
		);
	notech_ao4 i_769(.A(n_896), .B(n_458), .C(n_889), .D(n_457), .Z(n_935)
		);
	notech_reg_set dir1_reg_24(.CP(n_62043), .D(n_7341), .SD(n_61328), .Q(\dir1[24] 
		));
	notech_mux2 i_10018(.S(n_60470), .A(\dir1[24] ), .B(n_57566), .Z(n_7341)
		);
	notech_reg_set dir1_reg_25(.CP(n_62025), .D(n_7347), .SD(n_61310), .Q(\dir1[25] 
		));
	notech_mux2 i_10026(.S(n_60470), .A(\dir1[25] ), .B(n_57572), .Z(n_7347)
		);
	notech_ao4 i_767(.A(n_453), .B(iwrite_ack), .C(n_452), .D(n_10101), .Z(n_937
		));
	notech_reg_set dir1_reg_26(.CP(n_62025), .D(n_7353), .SD(n_61310), .Q(\dir1[26] 
		));
	notech_mux2 i_10034(.S(n_60470), .A(\dir1[26] ), .B(n_57578), .Z(n_7353)
		);
	notech_nand2 i_79132(.A(n_61926), .B(n_61193), .Z(n_938));
	notech_reg_set dir1_reg_27(.CP(n_62029), .D(n_7359), .SD(n_61314), .Q(\dir1[27] 
		));
	notech_mux2 i_10042(.S(n_60470), .A(\dir1[27] ), .B(n_57584), .Z(n_7359)
		);
	notech_reg_set dir1_reg_28(.CP(n_62025), .D(n_7365), .SD(n_61310), .Q(\dir1[28] 
		));
	notech_mux2 i_10050(.S(n_60470), .A(\dir1[28] ), .B(n_57590), .Z(n_7365)
		);
	notech_reg_set dir1_reg_29(.CP(n_62025), .D(n_7371), .SD(n_61310), .Q(\dir1[29] 
		));
	notech_mux2 i_10058(.S(n_60470), .A(\dir1[29] ), .B(n_57596), .Z(n_7371)
		);
	notech_reg_set dir1_reg_33(.CP(n_62025), .D(n_7377), .SD(n_61310), .Q(\dir1[33] 
		));
	notech_mux2 i_10066(.S(n_60470), .A(\dir1[33] ), .B(n_57621), .Z(n_7377)
		);
	notech_reg_set dir2_reg_0(.CP(n_62025), .D(n_7383), .SD(n_61310), .Q(\dir2[0] 
		));
	notech_mux2 i_10074(.S(\nbus_14490[0] ), .A(\dir2[0] ), .B(n_57422), .Z(n_7383
		));
	notech_reg_set dir2_reg_1(.CP(n_62029), .D(n_7389), .SD(n_61314), .Q(\dir2[1] 
		));
	notech_mux2 i_10082(.S(\nbus_14490[0] ), .A(\dir2[1] ), .B(n_57428), .Z(n_7389
		));
	notech_reg_set dir2_reg_2(.CP(n_62029), .D(n_7395), .SD(n_61314), .Q(\dir2[2] 
		));
	notech_mux2 i_10090(.S(\nbus_14490[0] ), .A(\dir2[2] ), .B(n_57434), .Z(n_7395
		));
	notech_and3 i_760(.A(n_852), .B(n_851), .C(n_853), .Z(n_945));
	notech_reg_set dir2_reg_3(.CP(n_62029), .D(n_7401), .SD(n_61314), .Q(\dir2[3] 
		));
	notech_mux2 i_10098(.S(\nbus_14490[0] ), .A(\dir2[3] ), .B(n_57440), .Z(n_7401
		));
	notech_reg dir2_reg_4(.CP(n_62029), .D(n_7407), .CD(n_61314), .Q(\dir2[4] 
		));
	notech_mux2 i_10106(.S(\nbus_14490[0] ), .A(\dir2[4] ), .B(n_874), .Z(n_7407
		));
	notech_or2 i_757(.A(fsm[2]), .B(fsm[3]), .Z(n_947));
	notech_reg_set dir2_reg_5(.CP(n_62029), .D(n_7413), .SD(n_61314), .Q(\dir2[5] 
		));
	notech_mux2 i_10114(.S(\nbus_14490[0] ), .A(\dir2[5] ), .B(n_57452), .Z(n_7413
		));
	notech_ao4 i_756(.A(n_458), .B(n_884), .C(n_449), .D(n_947), .Z(n_948)
		);
	notech_reg_set dir2_reg_6(.CP(n_62029), .D(n_7419), .SD(n_61314), .Q(\dir2[6] 
		));
	notech_mux2 i_10122(.S(\nbus_14490[0] ), .A(\dir2[6] ), .B(n_57458), .Z(n_7419
		));
	notech_or2 i_15(.A(\hit_dir1[7] ), .B(n_916), .Z(n_949));
	notech_reg_set dir2_reg_7(.CP(n_62029), .D(n_7425), .SD(n_61314), .Q(\dir2[7] 
		));
	notech_mux2 i_10130(.S(\nbus_14490[0] ), .A(\dir2[7] ), .B(n_57464), .Z(n_7425
		));
	notech_nao3 i_11(.A(n_61926), .B(\hit_dir1[7] ), .C(n_889), .Z(n_950));
	notech_reg_set dir2_reg_8(.CP(n_62025), .D(n_7431), .SD(n_61310), .Q(\dir2[8] 
		));
	notech_mux2 i_10138(.S(\nbus_14490[0] ), .A(\dir2[8] ), .B(n_57470), .Z(n_7431
		));
	notech_ao4 i_755(.A(n_950), .B(n_9867), .C(n_949), .D(n_9887), .Z(n_951)
		);
	notech_reg_set dir2_reg_9(.CP(n_62025), .D(n_7437), .SD(n_61310), .Q(\dir2[9] 
		));
	notech_mux2 i_10146(.S(\nbus_14490[0] ), .A(\dir2[9] ), .B(n_57476), .Z(n_7437
		));
	notech_ao4 i_754(.A(n_950), .B(n_9866), .C(n_949), .D(n_9886), .Z(n_952)
		);
	notech_reg_set dir2_reg_10(.CP(n_62025), .D(n_7443), .SD(n_61310), .Q(\dir2[10] 
		));
	notech_mux2 i_10154(.S(\nbus_14490[0] ), .A(\dir2[10] ), .B(n_57482), .Z
		(n_7443));
	notech_ao4 i_753(.A(n_950), .B(n_9865), .C(n_949), .D(n_9885), .Z(n_953)
		);
	notech_reg_set dir2_reg_11(.CP(n_62025), .D(n_7449), .SD(n_61310), .Q(\dir2[11] 
		));
	notech_mux2 i_10162(.S(\nbus_14490[0] ), .A(\dir2[11] ), .B(n_57488), .Z
		(n_7449));
	notech_ao4 i_752(.A(n_950), .B(n_9864), .C(n_949), .D(n_9884), .Z(n_954)
		);
	notech_reg_set dir2_reg_12(.CP(n_62025), .D(n_7455), .SD(n_61310), .Q(\dir2[12] 
		));
	notech_mux2 i_10170(.S(\nbus_14490[0] ), .A(\dir2[12] ), .B(n_57494), .Z
		(n_7455));
	notech_ao4 i_751(.A(n_950), .B(n_9863), .C(n_949), .D(n_9883), .Z(n_955)
		);
	notech_reg_set dir2_reg_13(.CP(n_62024), .D(n_7461), .SD(n_61309), .Q(\dir2[13] 
		));
	notech_mux2 i_10178(.S(\nbus_14490[0] ), .A(\dir2[13] ), .B(n_57500), .Z
		(n_7461));
	notech_ao4 i_750(.A(n_950), .B(n_9862), .C(n_949), .D(n_9882), .Z(n_956)
		);
	notech_reg_set dir2_reg_14(.CP(n_62024), .D(n_7467), .SD(n_61309), .Q(\dir2[14] 
		));
	notech_mux2 i_10186(.S(\nbus_14490[0] ), .A(\dir2[14] ), .B(n_57506), .Z
		(n_7467));
	notech_ao4 i_749(.A(n_950), .B(n_9861), .C(n_949), .D(n_9881), .Z(n_957)
		);
	notech_reg_set dir2_reg_15(.CP(n_62024), .D(n_7473), .SD(n_61309), .Q(\dir2[15] 
		));
	notech_mux2 i_10194(.S(\nbus_14490[0] ), .A(\dir2[15] ), .B(n_57512), .Z
		(n_7473));
	notech_ao4 i_748(.A(n_950), .B(n_9860), .C(n_949), .D(n_9880), .Z(n_958)
		);
	notech_reg_set dir2_reg_16(.CP(n_62025), .D(n_7479), .SD(n_61310), .Q(\dir2[16] 
		));
	notech_mux2 i_10202(.S(n_60525), .A(\dir2[16] ), .B(n_57518), .Z(n_7479)
		);
	notech_ao4 i_747(.A(n_950), .B(n_9859), .C(n_949), .D(n_9879), .Z(n_959)
		);
	notech_reg_set dir2_reg_17(.CP(n_62025), .D(n_7485), .SD(n_61310), .Q(\dir2[17] 
		));
	notech_mux2 i_10210(.S(n_60525), .A(\dir2[17] ), .B(n_57524), .Z(n_7485)
		);
	notech_ao4 i_746(.A(n_950), .B(n_9858), .C(n_949), .D(n_9878), .Z(n_960)
		);
	notech_reg_set dir2_reg_18(.CP(n_62025), .D(n_7491), .SD(n_61310), .Q(\dir2[18] 
		));
	notech_mux2 i_10218(.S(n_60525), .A(\dir2[18] ), .B(n_57530), .Z(n_7491)
		);
	notech_ao4 i_745(.A(n_950), .B(n_9857), .C(n_949), .D(n_9877), .Z(n_961)
		);
	notech_reg_set dir2_reg_19(.CP(n_62025), .D(n_7497), .SD(n_61310), .Q(\dir2[19] 
		));
	notech_mux2 i_10226(.S(n_60525), .A(\dir2[19] ), .B(n_57536), .Z(n_7497)
		);
	notech_ao4 i_744(.A(n_950), .B(n_9856), .C(n_949), .D(n_9876), .Z(n_962)
		);
	notech_reg_set dir2_reg_20(.CP(n_62025), .D(n_7503), .SD(n_61310), .Q(\dir2[20] 
		));
	notech_mux2 i_10234(.S(n_60525), .A(\dir2[20] ), .B(n_57542), .Z(n_7503)
		);
	notech_ao4 i_743(.A(n_950), .B(n_9855), .C(n_949), .D(n_9875), .Z(n_963)
		);
	notech_reg_set dir2_reg_21(.CP(n_62025), .D(n_7509), .SD(n_61310), .Q(\dir2[21] 
		));
	notech_mux2 i_10242(.S(n_60525), .A(\dir2[21] ), .B(n_57548), .Z(n_7509)
		);
	notech_ao4 i_742(.A(n_950), .B(n_9854), .C(n_949), .D(n_9874), .Z(n_964)
		);
	notech_reg_set dir2_reg_22(.CP(n_62025), .D(n_7515), .SD(n_61310), .Q(\dir2[22] 
		));
	notech_mux2 i_10250(.S(n_60525), .A(\dir2[22] ), .B(n_57554), .Z(n_7515)
		);
	notech_ao4 i_741(.A(n_950), .B(n_9853), .C(n_949), .D(n_9873), .Z(n_965)
		);
	notech_reg_set dir2_reg_23(.CP(n_62029), .D(n_7521), .SD(n_61314), .Q(\dir2[23] 
		));
	notech_mux2 i_10258(.S(n_60525), .A(\dir2[23] ), .B(n_57560), .Z(n_7521)
		);
	notech_ao4 i_740(.A(n_950), .B(n_9852), .C(n_949), .D(n_9872), .Z(n_966)
		);
	notech_reg_set dir2_reg_24(.CP(n_62033), .D(n_7527), .SD(n_61318), .Q(\dir2[24] 
		));
	notech_mux2 i_10266(.S(n_60525), .A(\dir2[24] ), .B(n_57566), .Z(n_7527)
		);
	notech_ao4 i_739(.A(n_950), .B(n_9851), .C(n_949), .D(n_9871), .Z(n_967)
		);
	notech_reg_set dir2_reg_25(.CP(n_62033), .D(n_7533), .SD(n_61318), .Q(\dir2[25] 
		));
	notech_mux2 i_10274(.S(n_60525), .A(\dir2[25] ), .B(n_57572), .Z(n_7533)
		);
	notech_ao4 i_738(.A(n_950), .B(n_9850), .C(n_949), .D(n_9870), .Z(n_968)
		);
	notech_reg_set dir2_reg_26(.CP(n_62033), .D(n_7539), .SD(n_61318), .Q(\dir2[26] 
		));
	notech_mux2 i_10282(.S(n_60525), .A(\dir2[26] ), .B(n_57578), .Z(n_7539)
		);
	notech_ao4 i_737(.A(n_950), .B(n_9849), .C(n_949), .D(n_9869), .Z(n_969)
		);
	notech_reg_set dir2_reg_27(.CP(n_62033), .D(n_7545), .SD(n_61318), .Q(\dir2[27] 
		));
	notech_mux2 i_10290(.S(n_60525), .A(\dir2[27] ), .B(n_57584), .Z(n_7545)
		);
	notech_ao4 i_736(.A(n_950), .B(n_9848), .C(n_949), .D(n_9868), .Z(n_970)
		);
	notech_reg_set dir2_reg_28(.CP(n_62033), .D(n_7551), .SD(n_61318), .Q(\dir2[28] 
		));
	notech_mux2 i_10298(.S(n_60525), .A(\dir2[28] ), .B(n_57590), .Z(n_7551)
		);
	notech_reg_set dir2_reg_29(.CP(n_62033), .D(n_7557), .SD(n_61318), .Q(\dir2[29] 
		));
	notech_mux2 i_10306(.S(n_60525), .A(\dir2[29] ), .B(n_57596), .Z(n_7557)
		);
	notech_ao3 i_030881(.A(n_61942), .B(n_9847), .C(n_61848), .Z(n_972));
	notech_reg_set dir2_reg_33(.CP(n_62033), .D(n_7563), .SD(n_61318), .Q(\dir2[33] 
		));
	notech_mux2 i_10314(.S(n_60525), .A(\dir2[33] ), .B(n_57621), .Z(n_7563)
		);
	notech_and2 i_725(.A(n_61942), .B(n_883), .Z(n_973));
	notech_reg_set tab21_reg_0(.CP(n_62033), .D(n_7569), .SD(n_61318), .Q(\tab21[0] 
		));
	notech_mux2 i_10322(.S(\nbus_14491[0] ), .A(\tab21[0] ), .B(n_57646), .Z
		(n_7569));
	notech_nao3 i_9(.A(n_61942), .B(n_883), .C(n_61852), .Z(n_974));
	notech_reg_set tab21_reg_1(.CP(n_62034), .D(n_7575), .SD(n_61319), .Q(\tab21[1] 
		));
	notech_mux2 i_10330(.S(\nbus_14491[0] ), .A(\tab21[1] ), .B(n_57652), .Z
		(n_7575));
	notech_ao4 i_724(.A(n_974), .B(n_10046), .C(n_399), .D(n_10102), .Z(n_975
		));
	notech_reg_set tab21_reg_2(.CP(n_62034), .D(n_7581), .SD(n_61319), .Q(\tab21[2] 
		));
	notech_mux2 i_10338(.S(\nbus_14491[0] ), .A(\tab21[2] ), .B(n_57658), .Z
		(n_7581));
	notech_ao4 i_723(.A(n_974), .B(n_10047), .C(n_399), .D(n_10103), .Z(n_976
		));
	notech_reg_set tab21_reg_3(.CP(n_62033), .D(n_7587), .SD(n_61318), .Q(\tab21[3] 
		));
	notech_mux2 i_10346(.S(\nbus_14491[0] ), .A(\tab21[3] ), .B(n_57664), .Z
		(n_7587));
	notech_ao4 i_722(.A(n_974), .B(n_10048), .C(n_399), .D(n_10104), .Z(n_977
		));
	notech_reg tab21_reg_4(.CP(n_62033), .D(n_7593), .CD(n_61318), .Q(\tab21[4] 
		));
	notech_mux2 i_10354(.S(\nbus_14491[0] ), .A(\tab21[4] ), .B(n_873), .Z(n_7593
		));
	notech_ao4 i_721(.A(n_974), .B(n_10049), .C(n_399), .D(n_10105), .Z(n_978
		));
	notech_reg_set tab21_reg_5(.CP(n_62033), .D(n_7599), .SD(n_61318), .Q(\tab21[5] 
		));
	notech_mux2 i_10362(.S(\nbus_14491[0] ), .A(\tab21[5] ), .B(n_57676), .Z
		(n_7599));
	notech_ao4 i_720(.A(n_974), .B(n_10050), .C(n_399), .D(n_10106), .Z(n_979
		));
	notech_reg_set tab21_reg_6(.CP(n_62033), .D(n_7605), .SD(n_61318), .Q(\tab21[6] 
		));
	notech_mux2 i_10370(.S(\nbus_14491[0] ), .A(\tab21[6] ), .B(n_57682), .Z
		(n_7605));
	notech_ao4 i_719(.A(n_974), .B(n_10051), .C(n_399), .D(n_10107), .Z(n_980
		));
	notech_reg_set tab21_reg_7(.CP(n_62033), .D(n_7611), .SD(n_61318), .Q(\tab21[7] 
		));
	notech_mux2 i_10378(.S(\nbus_14491[0] ), .A(\tab21[7] ), .B(n_57688), .Z
		(n_7611));
	notech_ao4 i_718(.A(n_974), .B(n_10052), .C(n_399), .D(n_10108), .Z(n_981
		));
	notech_reg_set tab21_reg_8(.CP(n_62029), .D(n_7617), .SD(n_61314), .Q(\tab21[8] 
		));
	notech_mux2 i_10386(.S(\nbus_14491[0] ), .A(\tab21[8] ), .B(n_57694), .Z
		(n_7617));
	notech_ao4 i_717(.A(n_974), .B(n_10053), .C(n_399), .D(n_10109), .Z(n_982
		));
	notech_reg_set tab21_reg_9(.CP(n_62029), .D(n_7623), .SD(n_61314), .Q(\tab21[9] 
		));
	notech_mux2 i_10394(.S(\nbus_14491[0] ), .A(\tab21[9] ), .B(n_57700), .Z
		(n_7623));
	notech_ao4 i_716(.A(n_974), .B(n_10054), .C(n_399), .D(n_10110), .Z(n_983
		));
	notech_reg_set tab21_reg_10(.CP(n_62029), .D(n_7629), .SD(n_61314), .Q(\tab21[10] 
		));
	notech_mux2 i_10402(.S(\nbus_14491[0] ), .A(\tab21[10] ), .B(n_57706), .Z
		(n_7629));
	notech_ao4 i_715(.A(n_974), .B(n_10055), .C(n_399), .D(n_10111), .Z(n_984
		));
	notech_reg_set tab21_reg_11(.CP(n_62029), .D(n_7635), .SD(n_61314), .Q(\tab21[11] 
		));
	notech_mux2 i_10410(.S(\nbus_14491[0] ), .A(\tab21[11] ), .B(n_57712), .Z
		(n_7635));
	notech_nand2 i_63(.A(\hit_dir1[7] ), .B(n_972), .Z(n_985));
	notech_reg_set tab21_reg_12(.CP(n_62029), .D(n_7641), .SD(n_61314), .Q(\tab21[12] 
		));
	notech_mux2 i_10418(.S(\nbus_14491[0] ), .A(\tab21[12] ), .B(n_57718), .Z
		(n_7641));
	notech_ao3 i_713(.A(hit_tab13), .B(n_10156), .C(hit_tab11), .Z(n_986));
	notech_reg_set tab21_reg_13(.CP(n_62029), .D(n_7647), .SD(n_61314), .Q(\tab21[13] 
		));
	notech_mux2 i_10426(.S(\nbus_14491[0] ), .A(\tab21[13] ), .B(n_57724), .Z
		(n_7647));
	notech_reg_set tab21_reg_14(.CP(n_62029), .D(n_7653), .SD(n_61314), .Q(\tab21[14] 
		));
	notech_mux2 i_10434(.S(\nbus_14491[0] ), .A(\tab21[14] ), .B(n_57730), .Z
		(n_7653));
	notech_or4 i_25(.A(hit_tab12), .B(hit_tab11), .C(hit_tab13), .D(n_985), 
		.Z(n_988));
	notech_reg_set tab21_reg_15(.CP(n_62033), .D(n_7659), .SD(n_61318), .Q(\tab21[15] 
		));
	notech_mux2 i_10442(.S(\nbus_14491[0] ), .A(\tab21[15] ), .B(n_57736), .Z
		(n_7659));
	notech_reg_set tab21_reg_16(.CP(n_62033), .D(n_7665), .SD(n_61318), .Q(\tab21[16] 
		));
	notech_mux2 i_10450(.S(n_60503), .A(\tab21[16] ), .B(n_57742), .Z(n_7665
		));
	notech_nao3 i_24(.A(hit_tab12), .B(n_61830), .C(hit_tab11), .Z(n_990));
	notech_reg_set tab21_reg_17(.CP(n_62033), .D(n_7671), .SD(n_61318), .Q(\tab21[17] 
		));
	notech_mux2 i_10458(.S(n_60503), .A(\tab21[17] ), .B(n_57748), .Z(n_7671
		));
	notech_ao4 i_708(.A(n_9910), .B(n_990), .C(n_988), .D(n_9934), .Z(n_991)
		);
	notech_reg_set tab21_reg_18(.CP(n_62033), .D(n_7677), .SD(n_61318), .Q(\tab21[18] 
		));
	notech_mux2 i_10466(.S(n_60503), .A(\tab21[18] ), .B(n_57754), .Z(n_7677
		));
	notech_reg_set tab21_reg_19(.CP(n_62029), .D(n_7683), .SD(n_61314), .Q(\tab21[19] 
		));
	notech_mux2 i_10474(.S(n_60503), .A(\tab21[19] ), .B(n_57760), .Z(n_7683
		));
	notech_or4 i_62(.A(n_61852), .B(\hit_dir1[7] ), .C(n_10158), .D(n_883), 
		.Z(n_993));
	notech_reg_set tab21_reg_20(.CP(n_62029), .D(n_7689), .SD(n_61314), .Q(\tab21[20] 
		));
	notech_mux2 i_10482(.S(n_60503), .A(\tab21[20] ), .B(n_57766), .Z(n_7689
		));
	notech_and2 i_711(.A(hit_tab22), .B(n_10154), .Z(n_994));
	notech_reg_set tab21_reg_21(.CP(n_62033), .D(n_7695), .SD(n_61318), .Q(\tab21[21] 
		));
	notech_mux2 i_10490(.S(n_60503), .A(\tab21[21] ), .B(n_57772), .Z(n_7695
		));
	notech_reg_set tab21_reg_22(.CP(n_62044), .D(n_7701), .SD(n_61329), .Q(\tab21[22] 
		));
	notech_mux2 i_10498(.S(n_60503), .A(\tab21[22] ), .B(n_57778), .Z(n_7701
		));
	notech_nand2 i_22(.A(hit_tab11), .B(n_61830), .Z(n_996));
	notech_reg_set tab21_reg_23(.CP(n_62057), .D(n_7707), .SD(n_61342), .Q(\tab21[23] 
		));
	notech_mux2 i_10506(.S(n_60503), .A(\tab21[23] ), .B(n_57784), .Z(n_7707
		));
	notech_reg_set tab21_reg_24(.CP(n_62057), .D(n_7713), .SD(n_61342), .Q(\tab21[24] 
		));
	notech_mux2 i_10514(.S(n_60503), .A(\tab21[24] ), .B(n_57790), .Z(n_7713
		));
	notech_or4 i_16(.A(hit_tab22), .B(hit_tab21), .C(n_61839), .D(n_10155), 
		.Z(n_998));
	notech_reg_set tab21_reg_25(.CP(n_62057), .D(n_7719), .SD(n_61342), .Q(\tab21[25] 
		));
	notech_mux2 i_10522(.S(n_60503), .A(\tab21[25] ), .B(n_57796), .Z(n_7719
		));
	notech_ao4 i_706(.A(n_998), .B(n_9963), .C(n_996), .D(n_10013), .Z(n_999
		));
	notech_reg_set tab21_reg_26(.CP(n_62057), .D(n_7725), .SD(n_61342), .Q(\tab21[26] 
		));
	notech_mux2 i_10530(.S(n_60503), .A(\tab21[26] ), .B(n_57802), .Z(n_7725
		));
	notech_reg_set tab21_reg_27(.CP(n_62057), .D(n_7731), .SD(n_61342), .Q(\tab21[27] 
		));
	notech_mux2 i_10538(.S(n_60503), .A(\tab21[27] ), .B(n_57808), .Z(n_7731
		));
	notech_and4 i_710(.A(n_999), .B(n_991), .C(n_776), .D(n_779), .Z(n_1001)
		);
	notech_reg_set tab21_reg_28(.CP(n_62057), .D(n_7737), .SD(n_61342), .Q(\tab21[28] 
		));
	notech_mux2 i_10546(.S(n_60503), .A(\tab21[28] ), .B(n_57814), .Z(n_7737
		));
	notech_nao3 i_13(.A(hit_tab21), .B(n_972), .C(\hit_dir1[7] ), .Z(n_1002)
		);
	notech_reg_set tab21_reg_29(.CP(n_62057), .D(n_7743), .SD(n_61342), .Q(\tab21[29] 
		));
	notech_mux2 i_10554(.S(n_60503), .A(\tab21[29] ), .B(n_57820), .Z(n_7743
		));
	notech_or4 i_12(.A(hit_tab22), .B(hit_tab21), .C(hit_tab23), .D(n_61839)
		, .Z(n_1003));
	notech_reg_set tab21_reg_33(.CP(n_62061), .D(n_7749), .SD(n_61346), .Q(\tab21[33] 
		));
	notech_mux2 i_10562(.S(n_60503), .A(\tab21[33] ), .B(n_57844), .Z(n_7749
		));
	notech_ao4 i_703(.A(n_1003), .B(n_9984), .C(n_1002), .D(n_9889), .Z(n_1004
		));
	notech_reg hit_adr11_reg(.CP(n_62061), .D(n_7755), .CD(n_61346), .Q(hit_adr11
		));
	notech_mux2 i_10570(.S(n_872), .A(hit_add11), .B(hit_adr11), .Z(n_7755)
		);
	notech_reg_set tab12_reg_0(.CP(n_62061), .D(n_7761), .SD(n_61346), .Q(\tab12[0] 
		));
	notech_mux2 i_10578(.S(\nbus_14500[0] ), .A(\tab12[0] ), .B(n_57646), .Z
		(n_7761));
	notech_ao4 i_702(.A(n_61937), .B(n_10112), .C(n_878), .D(n_10056), .Z(n_1006
		));
	notech_reg_set tab12_reg_1(.CP(n_62061), .D(n_7767), .SD(n_61346), .Q(\tab12[1] 
		));
	notech_mux2 i_10586(.S(\nbus_14500[0] ), .A(\tab12[1] ), .B(n_57652), .Z
		(n_7767));
	notech_reg_set tab12_reg_2(.CP(n_62057), .D(n_7773), .SD(n_61342), .Q(\tab12[2] 
		));
	notech_mux2 i_10594(.S(\nbus_14500[0] ), .A(\tab12[2] ), .B(n_57658), .Z
		(n_7773));
	notech_ao4 i_699(.A(n_990), .B(n_9911), .C(n_988), .D(n_9935), .Z(n_1008
		));
	notech_reg_set tab12_reg_3(.CP(n_62061), .D(n_7779), .SD(n_61346), .Q(\tab12[3] 
		));
	notech_mux2 i_10602(.S(\nbus_14500[0] ), .A(\tab12[3] ), .B(n_57664), .Z
		(n_7779));
	notech_reg tab12_reg_4(.CP(n_62061), .D(n_7785), .CD(n_61346), .Q(\tab12[4] 
		));
	notech_mux2 i_10610(.S(\nbus_14500[0] ), .A(\tab12[4] ), .B(n_873), .Z(n_7785
		));
	notech_ao4 i_697(.A(n_998), .B(n_9964), .C(n_996), .D(n_10014), .Z(n_1010
		));
	notech_reg_set tab12_reg_5(.CP(n_62057), .D(n_7791), .SD(n_61342), .Q(\tab12[5] 
		));
	notech_mux2 i_10618(.S(\nbus_14500[0] ), .A(\tab12[5] ), .B(n_57676), .Z
		(n_7791));
	notech_reg_set tab12_reg_6(.CP(n_62053), .D(n_7797), .SD(n_61338), .Q(\tab12[6] 
		));
	notech_mux2 i_10626(.S(\nbus_14500[0] ), .A(\tab12[6] ), .B(n_57682), .Z
		(n_7797));
	notech_and4 i_701(.A(n_1010), .B(n_1008), .C(n_765), .D(n_768), .Z(n_1012
		));
	notech_reg_set tab12_reg_7(.CP(n_62057), .D(n_7803), .SD(n_61342), .Q(\tab12[7] 
		));
	notech_mux2 i_10634(.S(\nbus_14500[0] ), .A(\tab12[7] ), .B(n_57688), .Z
		(n_7803));
	notech_ao4 i_694(.A(n_1003), .B(n_9985), .C(n_1002), .D(n_9890), .Z(n_1013
		));
	notech_reg_set tab12_reg_8(.CP(n_62057), .D(n_7809), .SD(n_61342), .Q(\tab12[8] 
		));
	notech_mux2 i_10642(.S(\nbus_14500[0] ), .A(\tab12[8] ), .B(n_57694), .Z
		(n_7809));
	notech_reg_set tab12_reg_9(.CP(n_62053), .D(n_7815), .SD(n_61338), .Q(\tab12[9] 
		));
	notech_mux2 i_10650(.S(\nbus_14500[0] ), .A(\tab12[9] ), .B(n_57700), .Z
		(n_7815));
	notech_ao4 i_693(.A(n_61937), .B(n_10113), .C(n_878), .D(n_10057), .Z(n_1015
		));
	notech_reg_set tab12_reg_10(.CP(n_62053), .D(n_7821), .SD(n_61338), .Q(\tab12[10] 
		));
	notech_mux2 i_10658(.S(\nbus_14500[0] ), .A(\tab12[10] ), .B(n_57706), .Z
		(n_7821));
	notech_reg_set tab12_reg_11(.CP(n_62053), .D(n_7827), .SD(n_61338), .Q(\tab12[11] 
		));
	notech_mux2 i_10666(.S(\nbus_14500[0] ), .A(\tab12[11] ), .B(n_57712), .Z
		(n_7827));
	notech_ao4 i_690(.A(n_990), .B(n_9912), .C(n_988), .D(n_9936), .Z(n_1017
		));
	notech_reg_set tab12_reg_12(.CP(n_62053), .D(n_7833), .SD(n_61338), .Q(\tab12[12] 
		));
	notech_mux2 i_10674(.S(\nbus_14500[0] ), .A(\tab12[12] ), .B(n_57718), .Z
		(n_7833));
	notech_reg_set tab12_reg_13(.CP(n_62057), .D(n_7839), .SD(n_61342), .Q(\tab12[13] 
		));
	notech_mux2 i_10682(.S(\nbus_14500[0] ), .A(\tab12[13] ), .B(n_57724), .Z
		(n_7839));
	notech_ao4 i_688(.A(n_998), .B(n_9965), .C(n_996), .D(n_10015), .Z(n_1019
		));
	notech_reg_set tab12_reg_14(.CP(n_62057), .D(n_7845), .SD(n_61342), .Q(\tab12[14] 
		));
	notech_mux2 i_10690(.S(\nbus_14500[0] ), .A(\tab12[14] ), .B(n_57730), .Z
		(n_7845));
	notech_reg_set tab12_reg_15(.CP(n_62057), .D(n_7851), .SD(n_61342), .Q(\tab12[15] 
		));
	notech_mux2 i_10698(.S(\nbus_14500[0] ), .A(\tab12[15] ), .B(n_57736), .Z
		(n_7851));
	notech_and4 i_692(.A(n_1019), .B(n_1017), .C(n_754), .D(n_757), .Z(n_1021
		));
	notech_reg_set tab12_reg_16(.CP(n_62057), .D(n_7857), .SD(n_61342), .Q(\tab12[16] 
		));
	notech_mux2 i_10706(.S(n_60459), .A(\tab12[16] ), .B(n_57742), .Z(n_7857
		));
	notech_ao4 i_685(.A(n_1003), .B(n_9986), .C(n_1002), .D(n_9891), .Z(n_1022
		));
	notech_reg_set tab12_reg_17(.CP(n_62057), .D(n_7863), .SD(n_61342), .Q(\tab12[17] 
		));
	notech_mux2 i_10714(.S(n_60459), .A(\tab12[17] ), .B(n_57748), .Z(n_7863
		));
	notech_reg_set tab12_reg_18(.CP(n_62057), .D(n_7869), .SD(n_61342), .Q(\tab12[18] 
		));
	notech_mux2 i_10722(.S(n_60459), .A(\tab12[18] ), .B(n_57754), .Z(n_7869
		));
	notech_ao4 i_684(.A(n_61937), .B(n_10114), .C(n_878), .D(n_10058), .Z(n_1024
		));
	notech_reg_set tab12_reg_19(.CP(n_62057), .D(n_7875), .SD(n_61342), .Q(\tab12[19] 
		));
	notech_mux2 i_10730(.S(n_60459), .A(\tab12[19] ), .B(n_57760), .Z(n_7875
		));
	notech_reg_set tab12_reg_20(.CP(n_62061), .D(n_7881), .SD(n_61346), .Q(\tab12[20] 
		));
	notech_mux2 i_10738(.S(n_60459), .A(\tab12[20] ), .B(n_57766), .Z(n_7881
		));
	notech_ao4 i_681(.A(n_990), .B(n_9913), .C(n_988), .D(n_9937), .Z(n_1026
		));
	notech_reg_set tab12_reg_21(.CP(n_62062), .D(n_7887), .SD(n_61347), .Q(\tab12[21] 
		));
	notech_mux2 i_10746(.S(n_60459), .A(\tab12[21] ), .B(n_57772), .Z(n_7887
		));
	notech_reg_set tab12_reg_22(.CP(n_62062), .D(n_7893), .SD(n_61347), .Q(\tab12[22] 
		));
	notech_mux2 i_10754(.S(n_60459), .A(\tab12[22] ), .B(n_57778), .Z(n_7893
		));
	notech_ao4 i_679(.A(n_998), .B(n_9966), .C(n_996), .D(n_10016), .Z(n_1028
		));
	notech_reg_set tab12_reg_23(.CP(n_62062), .D(n_7899), .SD(n_61347), .Q(\tab12[23] 
		));
	notech_mux2 i_10762(.S(n_60459), .A(\tab12[23] ), .B(n_57784), .Z(n_7899
		));
	notech_reg_set tab12_reg_24(.CP(n_62062), .D(n_7905), .SD(n_61347), .Q(\tab12[24] 
		));
	notech_mux2 i_10770(.S(n_60459), .A(\tab12[24] ), .B(n_57790), .Z(n_7905
		));
	notech_and4 i_683(.A(n_1028), .B(n_1026), .C(n_743), .D(n_746), .Z(n_1030
		));
	notech_reg_set tab12_reg_25(.CP(n_62062), .D(n_7911), .SD(n_61347), .Q(\tab12[25] 
		));
	notech_mux2 i_10778(.S(n_60459), .A(\tab12[25] ), .B(n_57796), .Z(n_7911
		));
	notech_ao4 i_676(.A(n_1003), .B(n_9987), .C(n_1002), .D(n_9892), .Z(n_1031
		));
	notech_reg_set tab12_reg_26(.CP(n_62062), .D(n_7917), .SD(n_61347), .Q(\tab12[26] 
		));
	notech_mux2 i_10786(.S(n_60459), .A(\tab12[26] ), .B(n_57802), .Z(n_7917
		));
	notech_reg_set tab12_reg_27(.CP(n_62062), .D(n_7923), .SD(n_61347), .Q(\tab12[27] 
		));
	notech_mux2 i_10794(.S(n_60459), .A(\tab12[27] ), .B(n_57808), .Z(n_7923
		));
	notech_ao4 i_675(.A(n_61937), .B(n_10115), .C(n_878), .D(n_10059), .Z(n_1033
		));
	notech_reg_set tab12_reg_28(.CP(n_62062), .D(n_7929), .SD(n_61347), .Q(\tab12[28] 
		));
	notech_mux2 i_10802(.S(n_60459), .A(\tab12[28] ), .B(n_57814), .Z(n_7929
		));
	notech_reg_set tab12_reg_29(.CP(n_62062), .D(n_7935), .SD(n_61347), .Q(\tab12[29] 
		));
	notech_mux2 i_10810(.S(n_60459), .A(\tab12[29] ), .B(n_57820), .Z(n_7935
		));
	notech_ao4 i_672(.A(n_990), .B(n_9914), .C(n_988), .D(n_9938), .Z(n_1035
		));
	notech_reg_set tab12_reg_33(.CP(n_62062), .D(n_7941), .SD(n_61347), .Q(\tab12[33] 
		));
	notech_mux2 i_10818(.S(n_60459), .A(\tab12[33] ), .B(n_57844), .Z(n_7941
		));
	notech_reg hit_adr12_reg(.CP(n_62062), .D(n_7947), .CD(n_61347), .Q(hit_adr12
		));
	notech_mux2 i_10826(.S(n_872), .A(hit_add12), .B(hit_adr12), .Z(n_7947)
		);
	notech_ao4 i_670(.A(n_998), .B(n_9967), .C(n_996), .D(n_10017), .Z(n_1037
		));
	notech_reg_set tab13_reg_0(.CP(n_62062), .D(n_7953), .SD(n_61347), .Q(\tab13[0] 
		));
	notech_mux2 i_10834(.S(\nbus_14503[0] ), .A(\tab13[0] ), .B(n_57646), .Z
		(n_7953));
	notech_reg_set tab13_reg_1(.CP(n_62062), .D(n_7959), .SD(n_61347), .Q(\tab13[1] 
		));
	notech_mux2 i_10842(.S(\nbus_14503[0] ), .A(\tab13[1] ), .B(n_57652), .Z
		(n_7959));
	notech_and4 i_674(.A(n_1037), .B(n_1035), .C(n_732), .D(n_735), .Z(n_1039
		));
	notech_reg_set tab13_reg_2(.CP(n_62062), .D(n_7965), .SD(n_61347), .Q(\tab13[2] 
		));
	notech_mux2 i_10850(.S(\nbus_14503[0] ), .A(\tab13[2] ), .B(n_57658), .Z
		(n_7965));
	notech_ao4 i_667(.A(n_1003), .B(n_9988), .C(n_1002), .D(n_9893), .Z(n_1040
		));
	notech_reg_set tab13_reg_3(.CP(n_62062), .D(n_7971), .SD(n_61347), .Q(\tab13[3] 
		));
	notech_mux2 i_10858(.S(\nbus_14503[0] ), .A(\tab13[3] ), .B(n_57664), .Z
		(n_7971));
	notech_reg tab13_reg_4(.CP(n_62061), .D(n_7977), .CD(n_61346), .Q(\tab13[4] 
		));
	notech_mux2 i_10866(.S(\nbus_14503[0] ), .A(\tab13[4] ), .B(n_873), .Z(n_7977
		));
	notech_ao4 i_666(.A(n_61937), .B(n_10116), .C(n_878), .D(n_10060), .Z(n_1042
		));
	notech_reg_set tab13_reg_5(.CP(n_62061), .D(n_7983), .SD(n_61346), .Q(\tab13[5] 
		));
	notech_mux2 i_10874(.S(\nbus_14503[0] ), .A(\tab13[5] ), .B(n_57676), .Z
		(n_7983));
	notech_reg_set tab13_reg_6(.CP(n_62061), .D(n_7989), .SD(n_61346), .Q(\tab13[6] 
		));
	notech_mux2 i_10882(.S(\nbus_14503[0] ), .A(\tab13[6] ), .B(n_57682), .Z
		(n_7989));
	notech_ao4 i_663(.A(n_990), .B(n_9915), .C(n_988), .D(n_9939), .Z(n_1044
		));
	notech_reg_set tab13_reg_7(.CP(n_62061), .D(n_7995), .SD(n_61346), .Q(\tab13[7] 
		));
	notech_mux2 i_10890(.S(\nbus_14503[0] ), .A(\tab13[7] ), .B(n_57688), .Z
		(n_7995));
	notech_reg_set tab13_reg_8(.CP(n_62061), .D(n_8001), .SD(n_61346), .Q(\tab13[8] 
		));
	notech_mux2 i_10898(.S(\nbus_14503[0] ), .A(\tab13[8] ), .B(n_57694), .Z
		(n_8001));
	notech_ao4 i_661(.A(n_998), .B(n_9968), .C(n_996), .D(n_10018), .Z(n_1046
		));
	notech_reg_set tab13_reg_9(.CP(n_62061), .D(n_8007), .SD(n_61346), .Q(\tab13[9] 
		));
	notech_mux2 i_10906(.S(\nbus_14503[0] ), .A(\tab13[9] ), .B(n_57700), .Z
		(n_8007));
	notech_reg_set tab13_reg_10(.CP(n_62061), .D(n_8013), .SD(n_61346), .Q(\tab13[10] 
		));
	notech_mux2 i_10914(.S(\nbus_14503[0] ), .A(\tab13[10] ), .B(n_57706), .Z
		(n_8013));
	notech_and4 i_665(.A(n_1046), .B(n_1044), .C(n_721), .D(n_724), .Z(n_1048
		));
	notech_reg_set tab13_reg_11(.CP(n_62062), .D(n_8019), .SD(n_61347), .Q(\tab13[11] 
		));
	notech_mux2 i_10922(.S(\nbus_14503[0] ), .A(\tab13[11] ), .B(n_57712), .Z
		(n_8019));
	notech_ao4 i_658(.A(n_1003), .B(n_9989), .C(n_1002), .D(n_9895), .Z(n_1049
		));
	notech_reg_set tab13_reg_12(.CP(n_62062), .D(n_8025), .SD(n_61347), .Q(\tab13[12] 
		));
	notech_mux2 i_10930(.S(\nbus_14503[0] ), .A(\tab13[12] ), .B(n_57718), .Z
		(n_8025));
	notech_reg_set tab13_reg_13(.CP(n_62062), .D(n_8031), .SD(n_61347), .Q(\tab13[13] 
		));
	notech_mux2 i_10938(.S(\nbus_14503[0] ), .A(\tab13[13] ), .B(n_57724), .Z
		(n_8031));
	notech_ao4 i_657(.A(n_61937), .B(n_10117), .C(n_878), .D(n_10061), .Z(n_1051
		));
	notech_reg_set tab13_reg_14(.CP(n_62061), .D(n_8037), .SD(n_61346), .Q(\tab13[14] 
		));
	notech_mux2 i_10946(.S(\nbus_14503[0] ), .A(\tab13[14] ), .B(n_57730), .Z
		(n_8037));
	notech_reg_set tab13_reg_15(.CP(n_62061), .D(n_8043), .SD(n_61346), .Q(\tab13[15] 
		));
	notech_mux2 i_10954(.S(\nbus_14503[0] ), .A(\tab13[15] ), .B(n_57736), .Z
		(n_8043));
	notech_ao4 i_654(.A(n_990), .B(n_9916), .C(n_988), .D(n_9940), .Z(n_1053
		));
	notech_reg_set tab13_reg_16(.CP(n_62061), .D(n_8049), .SD(n_61346), .Q(\tab13[16] 
		));
	notech_mux2 i_10962(.S(n_60437), .A(\tab13[16] ), .B(n_57742), .Z(n_8049
		));
	notech_reg_set tab13_reg_17(.CP(n_62061), .D(n_8055), .SD(n_61346), .Q(\tab13[17] 
		));
	notech_mux2 i_10970(.S(n_60437), .A(\tab13[17] ), .B(n_57748), .Z(n_8055
		));
	notech_ao4 i_652(.A(n_998), .B(n_9969), .C(n_996), .D(n_10019), .Z(n_1055
		));
	notech_reg_set tab13_reg_18(.CP(n_62048), .D(n_8061), .SD(n_61333), .Q(\tab13[18] 
		));
	notech_mux2 i_10978(.S(n_60437), .A(\tab13[18] ), .B(n_57754), .Z(n_8061
		));
	notech_reg_set tab13_reg_19(.CP(n_62048), .D(n_8067), .SD(n_61333), .Q(\tab13[19] 
		));
	notech_mux2 i_10986(.S(n_60437), .A(\tab13[19] ), .B(n_57760), .Z(n_8067
		));
	notech_and4 i_656(.A(n_1055), .B(n_1053), .C(n_710), .D(n_713), .Z(n_1057
		));
	notech_reg_set tab13_reg_20(.CP(n_62048), .D(n_8073), .SD(n_61333), .Q(\tab13[20] 
		));
	notech_mux2 i_10994(.S(n_60437), .A(\tab13[20] ), .B(n_57766), .Z(n_8073
		));
	notech_ao4 i_649(.A(n_1003), .B(n_9990), .C(n_1002), .D(n_9896), .Z(n_1058
		));
	notech_reg_set tab13_reg_21(.CP(n_62048), .D(n_8079), .SD(n_61333), .Q(\tab13[21] 
		));
	notech_mux2 i_11002(.S(n_60437), .A(\tab13[21] ), .B(n_57772), .Z(n_8079
		));
	notech_reg_set tab13_reg_22(.CP(n_62048), .D(n_8085), .SD(n_61333), .Q(\tab13[22] 
		));
	notech_mux2 i_11010(.S(n_60437), .A(\tab13[22] ), .B(n_57778), .Z(n_8085
		));
	notech_ao4 i_648(.A(n_61937), .B(n_10118), .C(n_878), .D(n_10062), .Z(n_1060
		));
	notech_reg_set tab13_reg_23(.CP(n_62048), .D(n_8091), .SD(n_61333), .Q(\tab13[23] 
		));
	notech_mux2 i_11018(.S(n_60437), .A(\tab13[23] ), .B(n_57784), .Z(n_8091
		));
	notech_reg_set tab13_reg_24(.CP(n_62048), .D(n_8097), .SD(n_61333), .Q(\tab13[24] 
		));
	notech_mux2 i_11026(.S(n_60437), .A(\tab13[24] ), .B(n_57790), .Z(n_8097
		));
	notech_ao4 i_645(.A(n_990), .B(n_9917), .C(n_988), .D(n_9941), .Z(n_1062
		));
	notech_reg_set tab13_reg_25(.CP(n_62048), .D(n_8103), .SD(n_61333), .Q(\tab13[25] 
		));
	notech_mux2 i_11034(.S(n_60437), .A(\tab13[25] ), .B(n_57796), .Z(n_8103
		));
	notech_reg_set tab13_reg_26(.CP(n_62048), .D(n_8109), .SD(n_61333), .Q(\tab13[26] 
		));
	notech_mux2 i_11042(.S(n_60437), .A(\tab13[26] ), .B(n_57802), .Z(n_8109
		));
	notech_ao4 i_643(.A(n_998), .B(n_9970), .C(n_996), .D(n_10020), .Z(n_1064
		));
	notech_reg_set tab13_reg_27(.CP(n_62052), .D(n_8115), .SD(n_61337), .Q(\tab13[27] 
		));
	notech_mux2 i_11050(.S(n_60437), .A(\tab13[27] ), .B(n_57808), .Z(n_8115
		));
	notech_reg_set tab13_reg_28(.CP(n_62048), .D(n_8121), .SD(n_61333), .Q(\tab13[28] 
		));
	notech_mux2 i_11058(.S(n_60437), .A(\tab13[28] ), .B(n_57814), .Z(n_8121
		));
	notech_and4 i_647(.A(n_1064), .B(n_1062), .C(n_699), .D(n_702), .Z(n_1066
		));
	notech_reg_set tab13_reg_29(.CP(n_62048), .D(n_8127), .SD(n_61333), .Q(\tab13[29] 
		));
	notech_mux2 i_11066(.S(n_60437), .A(\tab13[29] ), .B(n_57820), .Z(n_8127
		));
	notech_ao4 i_640(.A(n_1003), .B(n_9991), .C(n_1002), .D(n_9897), .Z(n_1067
		));
	notech_reg_set tab13_reg_33(.CP(n_62048), .D(n_8133), .SD(n_61333), .Q(\tab13[33] 
		));
	notech_mux2 i_11074(.S(n_60437), .A(\tab13[33] ), .B(n_57844), .Z(n_8133
		));
	notech_reg hit_adr13_reg(.CP(n_62048), .D(n_8139), .CD(n_61333), .Q(hit_adr13
		));
	notech_mux2 i_11082(.S(n_872), .A(hit_add13), .B(hit_adr13), .Z(n_8139)
		);
	notech_ao4 i_639(.A(n_61937), .B(n_10119), .C(n_878), .D(n_10063), .Z(n_1069
		));
	notech_reg_set tab14_reg_0(.CP(n_62048), .D(n_8145), .SD(n_61333), .Q(\tab14[0] 
		));
	notech_mux2 i_11090(.S(\nbus_14514[0] ), .A(\tab14[0] ), .B(n_57646), .Z
		(n_8145));
	notech_reg_set tab14_reg_1(.CP(n_62044), .D(n_8151), .SD(n_61329), .Q(\tab14[1] 
		));
	notech_mux2 i_11098(.S(\nbus_14514[0] ), .A(\tab14[1] ), .B(n_57652), .Z
		(n_8151));
	notech_ao4 i_636(.A(n_990), .B(n_9918), .C(n_988), .D(n_9942), .Z(n_1071
		));
	notech_reg_set tab14_reg_2(.CP(n_62044), .D(n_8157), .SD(n_61329), .Q(\tab14[2] 
		));
	notech_mux2 i_11106(.S(\nbus_14514[0] ), .A(\tab14[2] ), .B(n_57658), .Z
		(n_8157));
	notech_reg_set tab14_reg_3(.CP(n_62044), .D(n_8163), .SD(n_61329), .Q(\tab14[3] 
		));
	notech_mux2 i_11114(.S(\nbus_14514[0] ), .A(\tab14[3] ), .B(n_57664), .Z
		(n_8163));
	notech_ao4 i_634(.A(n_998), .B(n_9971), .C(n_996), .D(n_10021), .Z(n_1073
		));
	notech_reg tab14_reg_4(.CP(n_62044), .D(n_8169), .CD(n_61329), .Q(\tab14[4] 
		));
	notech_mux2 i_11122(.S(\nbus_14514[0] ), .A(\tab14[4] ), .B(n_873), .Z(n_8169
		));
	notech_reg_set tab14_reg_5(.CP(n_62044), .D(n_8175), .SD(n_61329), .Q(\tab14[5] 
		));
	notech_mux2 i_11130(.S(\nbus_14514[0] ), .A(\tab14[5] ), .B(n_57676), .Z
		(n_8175));
	notech_and4 i_638(.A(n_1073), .B(n_1071), .C(n_688), .D(n_691), .Z(n_1075
		));
	notech_reg_set tab14_reg_6(.CP(n_62044), .D(n_8181), .SD(n_61329), .Q(\tab14[6] 
		));
	notech_mux2 i_11138(.S(\nbus_14514[0] ), .A(\tab14[6] ), .B(n_57682), .Z
		(n_8181));
	notech_ao4 i_631(.A(n_1003), .B(n_9992), .C(n_1002), .D(n_9898), .Z(n_1076
		));
	notech_reg_set tab14_reg_7(.CP(n_62044), .D(n_8187), .SD(n_61329), .Q(\tab14[7] 
		));
	notech_mux2 i_11146(.S(\nbus_14514[0] ), .A(\tab14[7] ), .B(n_57688), .Z
		(n_8187));
	notech_reg_set tab14_reg_8(.CP(n_62048), .D(n_8193), .SD(n_61333), .Q(\tab14[8] 
		));
	notech_mux2 i_11154(.S(\nbus_14514[0] ), .A(\tab14[8] ), .B(n_57694), .Z
		(n_8193));
	notech_ao4 i_630(.A(n_61937), .B(n_10120), .C(n_878), .D(n_10064), .Z(n_1078
		));
	notech_reg_set tab14_reg_9(.CP(n_62048), .D(n_8199), .SD(n_61333), .Q(\tab14[9] 
		));
	notech_mux2 i_11162(.S(\nbus_14514[0] ), .A(\tab14[9] ), .B(n_57700), .Z
		(n_8199));
	notech_reg_set tab14_reg_10(.CP(n_62048), .D(n_8205), .SD(n_61333), .Q(\tab14[10] 
		));
	notech_mux2 i_11170(.S(\nbus_14514[0] ), .A(\tab14[10] ), .B(n_57706), .Z
		(n_8205));
	notech_ao4 i_627(.A(n_990), .B(n_9919), .C(n_988), .D(n_9943), .Z(n_1080
		));
	notech_reg_set tab14_reg_11(.CP(n_62048), .D(n_8211), .SD(n_61333), .Q(\tab14[11] 
		));
	notech_mux2 i_11178(.S(\nbus_14514[0] ), .A(\tab14[11] ), .B(n_57712), .Z
		(n_8211));
	notech_reg_set tab14_reg_12(.CP(n_62044), .D(n_8217), .SD(n_61329), .Q(\tab14[12] 
		));
	notech_mux2 i_11186(.S(\nbus_14514[0] ), .A(\tab14[12] ), .B(n_57718), .Z
		(n_8217));
	notech_ao4 i_625(.A(n_998), .B(n_9972), .C(n_996), .D(n_10022), .Z(n_1082
		));
	notech_reg_set tab14_reg_13(.CP(n_62044), .D(n_8223), .SD(n_61329), .Q(\tab14[13] 
		));
	notech_mux2 i_11194(.S(\nbus_14514[0] ), .A(\tab14[13] ), .B(n_57724), .Z
		(n_8223));
	notech_reg_set tab14_reg_14(.CP(n_62044), .D(n_8229), .SD(n_61329), .Q(\tab14[14] 
		));
	notech_mux2 i_11202(.S(\nbus_14514[0] ), .A(\tab14[14] ), .B(n_57730), .Z
		(n_8229));
	notech_and4 i_629(.A(n_1082), .B(n_1080), .C(n_677), .D(n_680), .Z(n_1084
		));
	notech_reg_set tab14_reg_15(.CP(n_62052), .D(n_8235), .SD(n_61337), .Q(\tab14[15] 
		));
	notech_mux2 i_11210(.S(\nbus_14514[0] ), .A(\tab14[15] ), .B(n_57736), .Z
		(n_8235));
	notech_ao4 i_622(.A(n_1003), .B(n_9993), .C(n_1002), .D(n_9899), .Z(n_1085
		));
	notech_reg_set tab14_reg_16(.CP(n_62053), .D(n_8241), .SD(n_61338), .Q(\tab14[16] 
		));
	notech_mux2 i_11218(.S(n_60426), .A(\tab14[16] ), .B(n_57742), .Z(n_8241
		));
	notech_reg_set tab14_reg_17(.CP(n_62053), .D(n_8247), .SD(n_61338), .Q(\tab14[17] 
		));
	notech_mux2 i_11226(.S(n_60426), .A(\tab14[17] ), .B(n_57748), .Z(n_8247
		));
	notech_ao4 i_621(.A(n_61937), .B(n_10121), .C(n_878), .D(n_10065), .Z(n_1087
		));
	notech_reg_set tab14_reg_18(.CP(n_62053), .D(n_8253), .SD(n_61338), .Q(\tab14[18] 
		));
	notech_mux2 i_11234(.S(n_60426), .A(\tab14[18] ), .B(n_57754), .Z(n_8253
		));
	notech_reg_set tab14_reg_19(.CP(n_62053), .D(n_8259), .SD(n_61338), .Q(\tab14[19] 
		));
	notech_mux2 i_11242(.S(n_60426), .A(\tab14[19] ), .B(n_57760), .Z(n_8259
		));
	notech_ao4 i_618(.A(n_990), .B(n_9920), .C(n_988), .D(n_9944), .Z(n_1089
		));
	notech_reg_set tab14_reg_20(.CP(n_62052), .D(n_8265), .SD(n_61337), .Q(\tab14[20] 
		));
	notech_mux2 i_11250(.S(n_60426), .A(\tab14[20] ), .B(n_57766), .Z(n_8265
		));
	notech_reg_set tab14_reg_21(.CP(n_62053), .D(n_8271), .SD(n_61338), .Q(\tab14[21] 
		));
	notech_mux2 i_11258(.S(n_60426), .A(\tab14[21] ), .B(n_57772), .Z(n_8271
		));
	notech_ao4 i_616(.A(n_998), .B(n_9973), .C(n_996), .D(n_10023), .Z(n_1091
		));
	notech_reg_set tab14_reg_22(.CP(n_62053), .D(n_8277), .SD(n_61338), .Q(\tab14[22] 
		));
	notech_mux2 i_11266(.S(n_60426), .A(\tab14[22] ), .B(n_57778), .Z(n_8277
		));
	notech_reg_set tab14_reg_23(.CP(n_62053), .D(n_8283), .SD(n_61338), .Q(\tab14[23] 
		));
	notech_mux2 i_11274(.S(n_60426), .A(\tab14[23] ), .B(n_57784), .Z(n_8283
		));
	notech_and4 i_620(.A(n_1091), .B(n_1089), .C(n_666), .D(n_669), .Z(n_1093
		));
	notech_reg_set tab14_reg_24(.CP(n_62053), .D(n_8289), .SD(n_61338), .Q(\tab14[24] 
		));
	notech_mux2 i_11282(.S(n_60426), .A(\tab14[24] ), .B(n_57790), .Z(n_8289
		));
	notech_ao4 i_613(.A(n_1003), .B(n_9994), .C(n_1002), .D(n_9900), .Z(n_1094
		));
	notech_reg_set tab14_reg_25(.CP(n_62053), .D(n_8295), .SD(n_61338), .Q(\tab14[25] 
		));
	notech_mux2 i_11290(.S(n_60426), .A(\tab14[25] ), .B(n_57796), .Z(n_8295
		));
	notech_reg_set tab14_reg_26(.CP(n_62053), .D(n_8301), .SD(n_61338), .Q(\tab14[26] 
		));
	notech_mux2 i_11298(.S(n_60426), .A(\tab14[26] ), .B(n_57802), .Z(n_8301
		));
	notech_ao4 i_612(.A(n_61937), .B(n_10122), .C(n_878), .D(n_10066), .Z(n_1096
		));
	notech_reg_set tab14_reg_27(.CP(n_62053), .D(n_8307), .SD(n_61338), .Q(\tab14[27] 
		));
	notech_mux2 i_11306(.S(n_60426), .A(\tab14[27] ), .B(n_57808), .Z(n_8307
		));
	notech_reg_set tab14_reg_28(.CP(n_62053), .D(n_8313), .SD(n_61338), .Q(\tab14[28] 
		));
	notech_mux2 i_11314(.S(n_60426), .A(\tab14[28] ), .B(n_57814), .Z(n_8313
		));
	notech_ao4 i_609(.A(n_990), .B(n_9921), .C(n_988), .D(n_9945), .Z(n_1098
		));
	notech_reg_set tab14_reg_29(.CP(n_62053), .D(n_8319), .SD(n_61338), .Q(\tab14[29] 
		));
	notech_mux2 i_11322(.S(n_60426), .A(\tab14[29] ), .B(n_57820), .Z(n_8319
		));
	notech_reg_set tab14_reg_33(.CP(n_62052), .D(n_8325), .SD(n_61337), .Q(\tab14[33] 
		));
	notech_mux2 i_11330(.S(n_60426), .A(\tab14[33] ), .B(n_57844), .Z(n_8325
		));
	notech_ao4 i_607(.A(n_998), .B(n_9974), .C(n_996), .D(n_10024), .Z(n_1100
		));
	notech_reg hit_adr14_reg(.CP(n_62052), .D(n_8331), .CD(n_61337), .Q(hit_adr14
		));
	notech_mux2 i_11338(.S(n_872), .A(hit_add14), .B(hit_adr14), .Z(n_8331)
		);
	notech_reg nx_tab1_reg_0(.CP(n_62052), .D(n_8337), .CD(n_61337), .Q(\nx_tab1[0] 
		));
	notech_mux2 i_11346(.S(\nbus_14495[0] ), .A(\nx_tab1[0] ), .B(n_9954), .Z
		(n_8337));
	notech_and4 i_611(.A(n_1100), .B(n_1098), .C(n_655), .D(n_658), .Z(n_1102
		));
	notech_reg nx_tab1_reg_1(.CP(n_62052), .D(n_8343), .CD(n_61337), .Q(\nx_tab1[1] 
		));
	notech_mux2 i_11354(.S(\nbus_14495[0] ), .A(\nx_tab1[1] ), .B(n_9956), .Z
		(n_8343));
	notech_ao4 i_604(.A(n_1003), .B(n_9995), .C(n_1002), .D(n_9901), .Z(n_1103
		));
	notech_reg_set nnx_tab1_reg_0(.CP(n_62052), .D(n_8349), .SD(n_61337), .Q
		(\nnx_tab1[0] ));
	notech_mux2 i_11362(.S(n_9962), .A(\nnx_tab1[0] ), .B(n_9958), .Z(n_8349
		));
	notech_reg nnx_tab1_reg_1(.CP(n_62052), .D(n_8355), .CD(n_61337), .Q(\nnx_tab1[1] 
		));
	notech_mux2 i_11370(.S(n_9962), .A(\nnx_tab1[1] ), .B(n_9960), .Z(n_8355
		));
	notech_ao4 i_603(.A(n_61941), .B(n_10123), .C(n_61901), .D(n_10067), .Z(n_1105
		));
	notech_reg hit_adr21_reg(.CP(n_62052), .D(n_8361), .CD(n_61337), .Q(hit_adr21
		));
	notech_mux2 i_11378(.S(n_872), .A(hit_add21), .B(hit_adr21), .Z(n_8361)
		);
	notech_reg_set tab22_reg_0(.CP(n_62052), .D(n_8367), .SD(n_61337), .Q(\tab22[0] 
		));
	notech_mux2 i_11386(.S(\nbus_14498[0] ), .A(\tab22[0] ), .B(n_57646), .Z
		(n_8367));
	notech_ao4 i_600(.A(n_990), .B(n_9922), .C(n_988), .D(n_9946), .Z(n_1107
		));
	notech_reg_set tab22_reg_1(.CP(n_62052), .D(n_8373), .SD(n_61337), .Q(\tab22[1] 
		));
	notech_mux2 i_11394(.S(\nbus_14498[0] ), .A(\tab22[1] ), .B(n_57652), .Z
		(n_8373));
	notech_reg_set tab22_reg_2(.CP(n_62052), .D(n_8379), .SD(n_61337), .Q(\tab22[2] 
		));
	notech_mux2 i_11402(.S(\nbus_14498[0] ), .A(\tab22[2] ), .B(n_57658), .Z
		(n_8379));
	notech_ao4 i_598(.A(n_998), .B(n_9975), .C(n_996), .D(n_10025), .Z(n_1109
		));
	notech_reg_set tab22_reg_3(.CP(n_62052), .D(n_8385), .SD(n_61337), .Q(\tab22[3] 
		));
	notech_mux2 i_11410(.S(\nbus_14498[0] ), .A(\tab22[3] ), .B(n_57664), .Z
		(n_8385));
	notech_reg tab22_reg_4(.CP(n_62052), .D(n_8391), .CD(n_61337), .Q(\tab22[4] 
		));
	notech_mux2 i_11418(.S(\nbus_14498[0] ), .A(\tab22[4] ), .B(n_873), .Z(n_8391
		));
	notech_and4 i_602(.A(n_1109), .B(n_1107), .C(n_644), .D(n_647), .Z(n_1111
		));
	notech_reg_set tab22_reg_5(.CP(n_62052), .D(n_8397), .SD(n_61337), .Q(\tab22[5] 
		));
	notech_mux2 i_11426(.S(\nbus_14498[0] ), .A(\tab22[5] ), .B(n_57676), .Z
		(n_8397));
	notech_ao4 i_595(.A(n_1003), .B(n_9996), .C(n_1002), .D(n_9902), .Z(n_1112
		));
	notech_reg_set tab22_reg_6(.CP(n_62052), .D(n_8403), .SD(n_61337), .Q(\tab22[6] 
		));
	notech_mux2 i_11434(.S(\nbus_14498[0] ), .A(\tab22[6] ), .B(n_57682), .Z
		(n_8403));
	notech_reg_set tab22_reg_7(.CP(n_62052), .D(n_8409), .SD(n_61337), .Q(\tab22[7] 
		));
	notech_mux2 i_11442(.S(\nbus_14498[0] ), .A(\tab22[7] ), .B(n_57688), .Z
		(n_8409));
	notech_ao4 i_594(.A(n_61941), .B(n_10124), .C(n_61901), .D(n_10068), .Z(n_1114
		));
	notech_reg_set tab22_reg_8(.CP(n_62024), .D(n_8415), .SD(n_61309), .Q(\tab22[8] 
		));
	notech_mux2 i_11450(.S(\nbus_14498[0] ), .A(\tab22[8] ), .B(n_57694), .Z
		(n_8415));
	notech_reg_set tab22_reg_9(.CP(n_61996), .D(n_8421), .SD(n_61281), .Q(\tab22[9] 
		));
	notech_mux2 i_11458(.S(\nbus_14498[0] ), .A(\tab22[9] ), .B(n_57700), .Z
		(n_8421));
	notech_ao4 i_591(.A(n_990), .B(n_9923), .C(n_988), .D(n_9947), .Z(n_1116
		));
	notech_reg_set tab22_reg_10(.CP(n_61996), .D(n_8427), .SD(n_61281), .Q(\tab22[10] 
		));
	notech_mux2 i_11466(.S(\nbus_14498[0] ), .A(\tab22[10] ), .B(n_57706), .Z
		(n_8427));
	notech_reg_set tab22_reg_11(.CP(n_61997), .D(n_8433), .SD(n_61282), .Q(\tab22[11] 
		));
	notech_mux2 i_11474(.S(\nbus_14498[0] ), .A(\tab22[11] ), .B(n_57712), .Z
		(n_8433));
	notech_ao4 i_589(.A(n_998), .B(n_9976), .C(n_996), .D(n_10026), .Z(n_1118
		));
	notech_reg_set tab22_reg_12(.CP(n_61996), .D(n_8439), .SD(n_61281), .Q(\tab22[12] 
		));
	notech_mux2 i_11482(.S(\nbus_14498[0] ), .A(\tab22[12] ), .B(n_57718), .Z
		(n_8439));
	notech_reg_set tab22_reg_13(.CP(n_61996), .D(n_8445), .SD(n_61281), .Q(\tab22[13] 
		));
	notech_mux2 i_11490(.S(\nbus_14498[0] ), .A(\tab22[13] ), .B(n_57724), .Z
		(n_8445));
	notech_and4 i_593(.A(n_1118), .B(n_1116), .C(n_633), .D(n_636), .Z(n_1120
		));
	notech_reg_set tab22_reg_14(.CP(n_61996), .D(n_8451), .SD(n_61281), .Q(\tab22[14] 
		));
	notech_mux2 i_11498(.S(\nbus_14498[0] ), .A(\tab22[14] ), .B(n_57730), .Z
		(n_8451));
	notech_ao4 i_586(.A(n_1003), .B(n_9997), .C(n_1002), .D(n_9903), .Z(n_1121
		));
	notech_reg_set tab22_reg_15(.CP(n_61996), .D(n_8457), .SD(n_61281), .Q(\tab22[15] 
		));
	notech_mux2 i_11506(.S(\nbus_14498[0] ), .A(\tab22[15] ), .B(n_57736), .Z
		(n_8457));
	notech_reg_set tab22_reg_16(.CP(n_61997), .D(n_8463), .SD(n_61282), .Q(\tab22[16] 
		));
	notech_mux2 i_11514(.S(n_60514), .A(\tab22[16] ), .B(n_57742), .Z(n_8463
		));
	notech_ao4 i_585(.A(n_61941), .B(n_10125), .C(n_61901), .D(n_10069), .Z(n_1123
		));
	notech_reg_set tab22_reg_17(.CP(n_61997), .D(n_8469), .SD(n_61282), .Q(\tab22[17] 
		));
	notech_mux2 i_11522(.S(n_60514), .A(\tab22[17] ), .B(n_57748), .Z(n_8469
		));
	notech_reg_set tab22_reg_18(.CP(n_61997), .D(n_8475), .SD(n_61282), .Q(\tab22[18] 
		));
	notech_mux2 i_11530(.S(n_60514), .A(\tab22[18] ), .B(n_57754), .Z(n_8475
		));
	notech_ao4 i_582(.A(n_990), .B(n_9924), .C(n_988), .D(n_9948), .Z(n_1125
		));
	notech_reg_set tab22_reg_19(.CP(n_61997), .D(n_8481), .SD(n_61282), .Q(\tab22[19] 
		));
	notech_mux2 i_11538(.S(n_60514), .A(\tab22[19] ), .B(n_57760), .Z(n_8481
		));
	notech_reg_set tab22_reg_20(.CP(n_61997), .D(n_8487), .SD(n_61282), .Q(\tab22[20] 
		));
	notech_mux2 i_11546(.S(n_60514), .A(\tab22[20] ), .B(n_57766), .Z(n_8487
		));
	notech_ao4 i_580(.A(n_998), .B(n_9977), .C(n_996), .D(n_10027), .Z(n_1127
		));
	notech_reg_set tab22_reg_21(.CP(n_61997), .D(n_8493), .SD(n_61282), .Q(\tab22[21] 
		));
	notech_mux2 i_11554(.S(n_60514), .A(\tab22[21] ), .B(n_57772), .Z(n_8493
		));
	notech_reg_set tab22_reg_22(.CP(n_61997), .D(n_8499), .SD(n_61282), .Q(\tab22[22] 
		));
	notech_mux2 i_11562(.S(n_60514), .A(\tab22[22] ), .B(n_57778), .Z(n_8499
		));
	notech_and4 i_584(.A(n_1127), .B(n_1125), .C(n_622), .D(n_625), .Z(n_1129
		));
	notech_reg_set tab22_reg_23(.CP(n_61996), .D(n_8505), .SD(n_61281), .Q(\tab22[23] 
		));
	notech_mux2 i_11570(.S(n_60514), .A(\tab22[23] ), .B(n_57784), .Z(n_8505
		));
	notech_ao4 i_577(.A(n_1003), .B(n_9998), .C(n_1002), .D(n_9904), .Z(n_1130
		));
	notech_reg_set tab22_reg_24(.CP(n_61992), .D(n_8511), .SD(n_61277), .Q(\tab22[24] 
		));
	notech_mux2 i_11578(.S(n_60514), .A(\tab22[24] ), .B(n_57790), .Z(n_8511
		));
	notech_reg_set tab22_reg_25(.CP(n_61996), .D(n_8517), .SD(n_61281), .Q(\tab22[25] 
		));
	notech_mux2 i_11586(.S(n_60514), .A(\tab22[25] ), .B(n_57796), .Z(n_8517
		));
	notech_ao4 i_576(.A(n_61941), .B(n_10126), .C(n_61901), .D(n_10070), .Z(n_1132
		));
	notech_reg_set tab22_reg_26(.CP(n_61996), .D(n_8523), .SD(n_61281), .Q(\tab22[26] 
		));
	notech_mux2 i_11594(.S(n_60514), .A(\tab22[26] ), .B(n_57802), .Z(n_8523
		));
	notech_reg_set tab22_reg_27(.CP(n_61992), .D(n_8529), .SD(n_61277), .Q(\tab22[27] 
		));
	notech_mux2 i_11602(.S(n_60514), .A(\tab22[27] ), .B(n_57808), .Z(n_8529
		));
	notech_ao4 i_573(.A(n_990), .B(n_9925), .C(n_988), .D(n_9949), .Z(n_1134
		));
	notech_reg_set tab22_reg_28(.CP(n_61992), .D(n_8535), .SD(n_61277), .Q(\tab22[28] 
		));
	notech_mux2 i_11610(.S(n_60514), .A(\tab22[28] ), .B(n_57814), .Z(n_8535
		));
	notech_reg_set tab22_reg_29(.CP(n_61992), .D(n_8541), .SD(n_61277), .Q(\tab22[29] 
		));
	notech_mux2 i_11618(.S(n_60514), .A(\tab22[29] ), .B(n_57820), .Z(n_8541
		));
	notech_ao4 i_571(.A(n_998), .B(n_9978), .C(n_996), .D(n_10028), .Z(n_1136
		));
	notech_reg_set tab22_reg_33(.CP(n_61992), .D(n_8547), .SD(n_61277), .Q(\tab22[33] 
		));
	notech_mux2 i_11626(.S(n_60514), .A(\tab22[33] ), .B(n_57844), .Z(n_8547
		));
	notech_reg hit_adr22_reg(.CP(n_61996), .D(n_8553), .CD(n_61281), .Q(hit_adr22
		));
	notech_mux2 i_11634(.S(n_872), .A(hit_add22), .B(hit_adr22), .Z(n_8553)
		);
	notech_and4 i_575(.A(n_1136), .B(n_1134), .C(n_611), .D(n_614), .Z(n_1138
		));
	notech_reg_set tab23_reg_0(.CP(n_61996), .D(n_8559), .SD(n_61281), .Q(\tab23[0] 
		));
	notech_mux2 i_11642(.S(\nbus_14502[0] ), .A(\tab23[0] ), .B(n_57646), .Z
		(n_8559));
	notech_ao4 i_568(.A(n_1003), .B(n_9999), .C(n_1002), .D(n_9905), .Z(n_1139
		));
	notech_reg_set tab23_reg_1(.CP(n_61996), .D(n_8565), .SD(n_61281), .Q(\tab23[1] 
		));
	notech_mux2 i_11650(.S(\nbus_14502[0] ), .A(\tab23[1] ), .B(n_57652), .Z
		(n_8565));
	notech_reg_set tab23_reg_2(.CP(n_61996), .D(n_8571), .SD(n_61281), .Q(\tab23[2] 
		));
	notech_mux2 i_11658(.S(\nbus_14502[0] ), .A(\tab23[2] ), .B(n_57658), .Z
		(n_8571));
	notech_ao4 i_567(.A(n_61941), .B(n_10127), .C(n_61901), .D(n_10071), .Z(n_1141
		));
	notech_reg_set tab23_reg_3(.CP(n_61996), .D(n_8577), .SD(n_61281), .Q(\tab23[3] 
		));
	notech_mux2 i_11666(.S(\nbus_14502[0] ), .A(\tab23[3] ), .B(n_57664), .Z
		(n_8577));
	notech_reg tab23_reg_4(.CP(n_61996), .D(n_8583), .CD(n_61281), .Q(\tab23[4] 
		));
	notech_mux2 i_11674(.S(\nbus_14502[0] ), .A(\tab23[4] ), .B(n_873), .Z(n_8583
		));
	notech_ao4 i_564(.A(n_990), .B(n_9926), .C(n_988), .D(n_9950), .Z(n_1143
		));
	notech_reg_set tab23_reg_5(.CP(n_61996), .D(n_8589), .SD(n_61281), .Q(\tab23[5] 
		));
	notech_mux2 i_11682(.S(\nbus_14502[0] ), .A(\tab23[5] ), .B(n_57676), .Z
		(n_8589));
	notech_reg_set tab23_reg_6(.CP(n_61997), .D(n_8595), .SD(n_61282), .Q(\tab23[6] 
		));
	notech_mux2 i_11690(.S(\nbus_14502[0] ), .A(\tab23[6] ), .B(n_57682), .Z
		(n_8595));
	notech_ao4 i_562(.A(n_998), .B(n_9979), .C(n_996), .D(n_10029), .Z(n_1145
		));
	notech_reg_set tab23_reg_7(.CP(n_62001), .D(n_8601), .SD(n_61286), .Q(\tab23[7] 
		));
	notech_mux2 i_11698(.S(\nbus_14502[0] ), .A(\tab23[7] ), .B(n_57688), .Z
		(n_8601));
	notech_reg_set tab23_reg_8(.CP(n_62001), .D(n_8607), .SD(n_61286), .Q(\tab23[8] 
		));
	notech_mux2 i_11706(.S(\nbus_14502[0] ), .A(\tab23[8] ), .B(n_57694), .Z
		(n_8607));
	notech_and4 i_566(.A(n_1145), .B(n_1143), .C(n_600), .D(n_603), .Z(n_1147
		));
	notech_reg_set tab23_reg_9(.CP(n_62001), .D(n_8613), .SD(n_61286), .Q(\tab23[9] 
		));
	notech_mux2 i_11714(.S(\nbus_14502[0] ), .A(\tab23[9] ), .B(n_57700), .Z
		(n_8613));
	notech_ao4 i_559(.A(n_1003), .B(n_10000), .C(n_1002), .D(n_9906), .Z(n_1148
		));
	notech_reg_set tab23_reg_10(.CP(n_62001), .D(n_8619), .SD(n_61286), .Q(\tab23[10] 
		));
	notech_mux2 i_11722(.S(\nbus_14502[0] ), .A(\tab23[10] ), .B(n_57706), .Z
		(n_8619));
	notech_reg_set tab23_reg_11(.CP(n_62001), .D(n_8625), .SD(n_61286), .Q(\tab23[11] 
		));
	notech_mux2 i_11730(.S(\nbus_14502[0] ), .A(\tab23[11] ), .B(n_57712), .Z
		(n_8625));
	notech_ao4 i_558(.A(n_61937), .B(n_10128), .C(n_61901), .D(n_10072), .Z(n_1150
		));
	notech_reg_set tab23_reg_12(.CP(n_62001), .D(n_8631), .SD(n_61286), .Q(\tab23[12] 
		));
	notech_mux2 i_11738(.S(\nbus_14502[0] ), .A(\tab23[12] ), .B(n_57718), .Z
		(n_8631));
	notech_reg_set tab23_reg_13(.CP(n_62001), .D(n_8637), .SD(n_61286), .Q(\tab23[13] 
		));
	notech_mux2 i_11746(.S(\nbus_14502[0] ), .A(\tab23[13] ), .B(n_57724), .Z
		(n_8637));
	notech_ao4 i_555(.A(n_990), .B(n_9927), .C(n_988), .D(n_9951), .Z(n_1152
		));
	notech_reg_set tab23_reg_14(.CP(n_62005), .D(n_8643), .SD(n_61290), .Q(\tab23[14] 
		));
	notech_mux2 i_11754(.S(\nbus_14502[0] ), .A(\tab23[14] ), .B(n_57730), .Z
		(n_8643));
	notech_reg_set tab23_reg_15(.CP(n_62005), .D(n_8649), .SD(n_61290), .Q(\tab23[15] 
		));
	notech_mux2 i_11762(.S(\nbus_14502[0] ), .A(\tab23[15] ), .B(n_57736), .Z
		(n_8649));
	notech_ao4 i_553(.A(n_998), .B(n_9980), .C(n_996), .D(n_10030), .Z(n_1154
		));
	notech_reg_set tab23_reg_16(.CP(n_62005), .D(n_8655), .SD(n_61290), .Q(\tab23[16] 
		));
	notech_mux2 i_11770(.S(n_60481), .A(\tab23[16] ), .B(n_57742), .Z(n_8655
		));
	notech_reg_set tab23_reg_17(.CP(n_62001), .D(n_8661), .SD(n_61286), .Q(\tab23[17] 
		));
	notech_mux2 i_11778(.S(n_60481), .A(\tab23[17] ), .B(n_57748), .Z(n_8661
		));
	notech_and4 i_557(.A(n_1154), .B(n_1152), .C(n_589), .D(n_592), .Z(n_1156
		));
	notech_reg_set tab23_reg_18(.CP(n_62001), .D(n_8667), .SD(n_61286), .Q(\tab23[18] 
		));
	notech_mux2 i_11786(.S(n_60481), .A(\tab23[18] ), .B(n_57754), .Z(n_8667
		));
	notech_ao4 i_550(.A(n_1003), .B(n_10001), .C(n_1002), .D(n_9907), .Z(n_1157
		));
	notech_reg_set tab23_reg_19(.CP(n_62001), .D(n_8673), .SD(n_61286), .Q(\tab23[19] 
		));
	notech_mux2 i_11794(.S(n_60481), .A(\tab23[19] ), .B(n_57760), .Z(n_8673
		));
	notech_reg_set tab23_reg_20(.CP(n_62001), .D(n_8679), .SD(n_61286), .Q(\tab23[20] 
		));
	notech_mux2 i_11802(.S(n_60481), .A(\tab23[20] ), .B(n_57766), .Z(n_8679
		));
	notech_ao4 i_549(.A(n_61937), .B(n_10129), .C(n_61901), .D(n_10073), .Z(n_1159
		));
	notech_reg_set tab23_reg_21(.CP(n_62001), .D(n_8685), .SD(n_61286), .Q(\tab23[21] 
		));
	notech_mux2 i_11810(.S(n_60481), .A(\tab23[21] ), .B(n_57772), .Z(n_8685
		));
	notech_reg_set tab23_reg_22(.CP(n_61997), .D(n_8691), .SD(n_61282), .Q(\tab23[22] 
		));
	notech_mux2 i_11818(.S(n_60481), .A(\tab23[22] ), .B(n_57778), .Z(n_8691
		));
	notech_ao4 i_546(.A(n_990), .B(n_9928), .C(n_988), .D(n_9952), .Z(n_1161
		));
	notech_reg_set tab23_reg_23(.CP(n_61997), .D(n_8697), .SD(n_61282), .Q(\tab23[23] 
		));
	notech_mux2 i_11826(.S(n_60481), .A(\tab23[23] ), .B(n_57784), .Z(n_8697
		));
	notech_reg_set tab23_reg_24(.CP(n_61997), .D(n_8703), .SD(n_61282), .Q(\tab23[24] 
		));
	notech_mux2 i_11834(.S(n_60481), .A(\tab23[24] ), .B(n_57790), .Z(n_8703
		));
	notech_ao4 i_544(.A(n_998), .B(n_9981), .C(n_996), .D(n_10031), .Z(n_1163
		));
	notech_reg_set tab23_reg_25(.CP(n_61997), .D(n_8709), .SD(n_61282), .Q(\tab23[25] 
		));
	notech_mux2 i_11842(.S(n_60481), .A(\tab23[25] ), .B(n_57796), .Z(n_8709
		));
	notech_reg_set tab23_reg_26(.CP(n_61997), .D(n_8715), .SD(n_61282), .Q(\tab23[26] 
		));
	notech_mux2 i_11850(.S(n_60481), .A(\tab23[26] ), .B(n_57802), .Z(n_8715
		));
	notech_and4 i_548(.A(n_1163), .B(n_1161), .C(n_578), .D(n_581), .Z(n_1165
		));
	notech_reg_set tab23_reg_27(.CP(n_61997), .D(n_8721), .SD(n_61282), .Q(\tab23[27] 
		));
	notech_mux2 i_11858(.S(n_60481), .A(\tab23[27] ), .B(n_57808), .Z(n_8721
		));
	notech_ao4 i_541(.A(n_1003), .B(n_10002), .C(n_1002), .D(n_9908), .Z(n_1166
		));
	notech_reg_set tab23_reg_28(.CP(n_61997), .D(n_8727), .SD(n_61282), .Q(\tab23[28] 
		));
	notech_mux2 i_11866(.S(n_60481), .A(\tab23[28] ), .B(n_57814), .Z(n_8727
		));
	notech_reg_set tab23_reg_29(.CP(n_62001), .D(n_8733), .SD(n_61286), .Q(\tab23[29] 
		));
	notech_mux2 i_11874(.S(n_60481), .A(\tab23[29] ), .B(n_57820), .Z(n_8733
		));
	notech_ao4 i_540(.A(n_61937), .B(n_10130), .C(n_878), .D(n_10074), .Z(n_1168
		));
	notech_reg_set tab23_reg_33(.CP(n_62001), .D(n_8739), .SD(n_61286), .Q(\tab23[33] 
		));
	notech_mux2 i_11882(.S(n_60481), .A(\tab23[33] ), .B(n_57844), .Z(n_8739
		));
	notech_reg hit_adr23_reg(.CP(n_62001), .D(n_8745), .CD(n_61286), .Q(hit_adr23
		));
	notech_mux2 i_11890(.S(n_872), .A(hit_add23), .B(hit_adr23), .Z(n_8745)
		);
	notech_ao4 i_537(.A(n_990), .B(n_9929), .C(n_988), .D(n_9953), .Z(n_1170
		));
	notech_reg_set tab24_reg_0(.CP(n_62001), .D(n_8751), .SD(n_61286), .Q(\tab24[0] 
		));
	notech_mux2 i_11898(.S(\nbus_14513[0] ), .A(\tab24[0] ), .B(n_57646), .Z
		(n_8751));
	notech_reg_set tab24_reg_1(.CP(n_61997), .D(n_8757), .SD(n_61282), .Q(\tab24[1] 
		));
	notech_mux2 i_11906(.S(\nbus_14513[0] ), .A(\tab24[1] ), .B(n_57652), .Z
		(n_8757));
	notech_ao4 i_535(.A(n_998), .B(n_9982), .C(n_996), .D(n_10032), .Z(n_1172
		));
	notech_reg_set tab24_reg_2(.CP(n_62001), .D(n_8763), .SD(n_61286), .Q(\tab24[2] 
		));
	notech_mux2 i_11914(.S(\nbus_14513[0] ), .A(\tab24[2] ), .B(n_57658), .Z
		(n_8763));
	notech_reg_set tab24_reg_3(.CP(n_62001), .D(n_8769), .SD(n_61286), .Q(\tab24[3] 
		));
	notech_mux2 i_11922(.S(\nbus_14513[0] ), .A(\tab24[3] ), .B(n_57664), .Z
		(n_8769));
	notech_and4 i_539(.A(n_1172), .B(n_1170), .C(n_567), .D(n_570), .Z(n_1174
		));
	notech_reg tab24_reg_4(.CP(n_61987), .D(n_8775), .CD(n_61272), .Q(\tab24[4] 
		));
	notech_mux2 i_11930(.S(\nbus_14513[0] ), .A(\tab24[4] ), .B(n_873), .Z(n_8775
		));
	notech_ao4 i_532(.A(n_1003), .B(n_10003), .C(n_1002), .D(n_9909), .Z(n_1175
		));
	notech_reg_set tab24_reg_5(.CP(n_61987), .D(n_8781), .SD(n_61272), .Q(\tab24[5] 
		));
	notech_mux2 i_11938(.S(\nbus_14513[0] ), .A(\tab24[5] ), .B(n_57676), .Z
		(n_8781));
	notech_reg_set tab24_reg_6(.CP(n_61987), .D(n_8787), .SD(n_61272), .Q(\tab24[6] 
		));
	notech_mux2 i_11946(.S(\nbus_14513[0] ), .A(\tab24[6] ), .B(n_57682), .Z
		(n_8787));
	notech_ao4 i_531(.A(n_61941), .B(n_10131), .C(n_61901), .D(n_10075), .Z(n_1177
		));
	notech_reg_set tab24_reg_7(.CP(n_61987), .D(n_8793), .SD(n_61272), .Q(\tab24[7] 
		));
	notech_mux2 i_11954(.S(\nbus_14513[0] ), .A(\tab24[7] ), .B(n_57688), .Z
		(n_8793));
	notech_reg_set tab24_reg_8(.CP(n_61983), .D(n_8799), .SD(n_61268), .Q(\tab24[8] 
		));
	notech_mux2 i_11962(.S(\nbus_14513[0] ), .A(\tab24[8] ), .B(n_57694), .Z
		(n_8799));
	notech_ao4 i_79165(.A(n_10079), .B(n_10158), .C(n_9930), .D(n_10159), .Z
		(oread_req100140));
	notech_reg_set tab24_reg_9(.CP(n_61987), .D(n_8805), .SD(n_61272), .Q(\tab24[9] 
		));
	notech_mux2 i_11970(.S(\nbus_14513[0] ), .A(\tab24[9] ), .B(n_57700), .Z
		(n_8805));
	notech_nand3 i_81221(.A(n_532), .B(n_388), .C(n_531), .Z(\nbus_14501[0] 
		));
	notech_reg_set tab24_reg_10(.CP(n_61987), .D(n_8811), .SD(n_61272), .Q(\tab24[10] 
		));
	notech_mux2 i_11978(.S(\nbus_14513[0] ), .A(\tab24[10] ), .B(n_57706), .Z
		(n_8811));
	notech_nand3 i_80438(.A(n_532), .B(n_388), .C(n_528), .Z(\nbus_14490[0] 
		));
	notech_reg_set tab24_reg_11(.CP(n_61987), .D(n_8817), .SD(n_61272), .Q(\tab24[11] 
		));
	notech_mux2 i_11986(.S(\nbus_14513[0] ), .A(\tab24[11] ), .B(n_57712), .Z
		(n_8817));
	notech_nand3 i_80557(.A(n_509), .B(n_388), .C(n_508), .Z(\nbus_14491[0] 
		));
	notech_reg_set tab24_reg_12(.CP(n_61987), .D(n_8823), .SD(n_61272), .Q(\tab24[12] 
		));
	notech_mux2 i_11994(.S(\nbus_14513[0] ), .A(\tab24[12] ), .B(n_57718), .Z
		(n_8823));
	notech_nand3 i_81112(.A(n_505), .B(n_388), .C(n_504), .Z(\nbus_14500[0] 
		));
	notech_reg_set tab24_reg_13(.CP(n_61987), .D(n_8829), .SD(n_61272), .Q(\tab24[13] 
		));
	notech_mux2 i_12002(.S(\nbus_14513[0] ), .A(\tab24[13] ), .B(n_57724), .Z
		(n_8829));
	notech_nand3 i_81445(.A(n_505), .B(n_388), .C(n_503), .Z(\nbus_14503[0] 
		));
	notech_reg_set tab24_reg_14(.CP(n_61987), .D(n_8835), .SD(n_61272), .Q(\tab24[14] 
		));
	notech_mux2 i_12010(.S(\nbus_14513[0] ), .A(\tab24[14] ), .B(n_57730), .Z
		(n_8835));
	notech_nand3 i_81823(.A(n_505), .B(n_388), .C(n_502), .Z(\nbus_14514[0] 
		));
	notech_reg_set tab24_reg_15(.CP(n_61987), .D(n_8841), .SD(n_61272), .Q(\tab24[15] 
		));
	notech_mux2 i_12018(.S(\nbus_14513[0] ), .A(\tab24[15] ), .B(n_57736), .Z
		(n_8841));
	notech_nand2 i_80831(.A(n_919), .B(n_911), .Z(\nbus_14495[0] ));
	notech_reg_set tab24_reg_16(.CP(n_61987), .D(n_8847), .SD(n_61272), .Q(\tab24[16] 
		));
	notech_mux2 i_12026(.S(n_60492), .A(\tab24[16] ), .B(n_57742), .Z(n_8847
		));
	notech_ao4 i_80309(.A(n_899), .B(n_910), .C(n_919), .D(n_9894), .Z(\nbus_14489[0] 
		));
	notech_reg_set tab24_reg_17(.CP(n_61987), .D(n_8853), .SD(n_61272), .Q(\tab24[17] 
		));
	notech_mux2 i_12034(.S(n_60492), .A(\tab24[17] ), .B(n_57748), .Z(n_8853
		));
	notech_nand3 i_80970(.A(n_509), .B(n_388), .C(n_484), .Z(\nbus_14498[0] 
		));
	notech_reg_set tab24_reg_18(.CP(n_61983), .D(n_8859), .SD(n_61268), .Q(\tab24[18] 
		));
	notech_mux2 i_12042(.S(n_60492), .A(\tab24[18] ), .B(n_57754), .Z(n_8859
		));
	notech_nand3 i_81333(.A(n_509), .B(n_388), .C(n_483), .Z(\nbus_14502[0] 
		));
	notech_reg_set tab24_reg_19(.CP(n_61983), .D(n_8865), .SD(n_61268), .Q(\tab24[19] 
		));
	notech_mux2 i_12050(.S(n_60492), .A(\tab24[19] ), .B(n_57760), .Z(n_8865
		));
	notech_nand3 i_81670(.A(n_509), .B(n_388), .C(n_482), .Z(\nbus_14513[0] 
		));
	notech_reg_set tab24_reg_20(.CP(n_61983), .D(n_8871), .SD(n_61268), .Q(\tab24[20] 
		));
	notech_mux2 i_12058(.S(n_60492), .A(\tab24[20] ), .B(n_57766), .Z(n_8871
		));
	notech_ao4 i_81940(.A(n_899), .B(n_900), .C(n_919), .D(n_9888), .Z(\nbus_14515[0] 
		));
	notech_reg_set tab24_reg_21(.CP(n_61983), .D(n_8877), .SD(n_61268), .Q(\tab24[21] 
		));
	notech_mux2 i_12066(.S(n_60492), .A(\tab24[21] ), .B(n_57772), .Z(n_8877
		));
	notech_nand2 i_81957(.A(n_919), .B(n_901), .Z(\nbus_14516[0] ));
	notech_reg_set tab24_reg_22(.CP(n_61983), .D(n_8883), .SD(n_61268), .Q(\tab24[22] 
		));
	notech_mux2 i_12074(.S(n_60492), .A(\tab24[22] ), .B(n_57778), .Z(n_8883
		));
	notech_nand3 i_80669(.A(n_505), .B(n_388), .C(n_464), .Z(\nbus_14492[0] 
		));
	notech_reg_set tab24_reg_23(.CP(n_61983), .D(n_8889), .SD(n_61268), .Q(\tab24[23] 
		));
	notech_mux2 i_12082(.S(n_60492), .A(\tab24[23] ), .B(n_57784), .Z(n_8889
		));
	notech_nand2 i_81075(.A(n_893), .B(n_462), .Z(\nbus_14499[0] ));
	notech_reg_set tab24_reg_24(.CP(n_61983), .D(n_8895), .SD(n_61268), .Q(\tab24[24] 
		));
	notech_mux2 i_12090(.S(n_60492), .A(\tab24[24] ), .B(n_57790), .Z(n_8895
		));
	notech_ao4 i_81810(.A(n_461), .B(n_932), .C(n_887), .D(n_10076), .Z(n_59947
		));
	notech_reg_set tab24_reg_25(.CP(n_61983), .D(n_8901), .SD(n_61268), .Q(\tab24[25] 
		));
	notech_mux2 i_12098(.S(n_60492), .A(\tab24[25] ), .B(n_57796), .Z(n_8901
		));
	notech_nand3 i_80788(.A(n_61901), .B(n_59947), .C(n_945), .Z(\nbus_14493[0] 
		));
	notech_reg_set tab24_reg_26(.CP(n_61983), .D(n_8907), .SD(n_61268), .Q(\tab24[26] 
		));
	notech_mux2 i_12106(.S(n_60492), .A(\tab24[26] ), .B(n_57802), .Z(n_8907
		));
	notech_nand2 i_79652(.A(n_938), .B(n_916), .Z(n_58109));
	notech_reg_set tab24_reg_27(.CP(n_61983), .D(n_8913), .SD(n_61268), .Q(\tab24[27] 
		));
	notech_mux2 i_12114(.S(n_60492), .A(\tab24[27] ), .B(n_57808), .Z(n_8913
		));
	notech_ao4 i_80864(.A(n_876), .B(data_miss[5]), .C(n_899), .D(n_934), .Z
		(\nbus_14497[0] ));
	notech_reg_set tab24_reg_28(.CP(n_61983), .D(n_8919), .SD(n_61268), .Q(\tab24[28] 
		));
	notech_mux2 i_12122(.S(n_60492), .A(\tab24[28] ), .B(n_57814), .Z(n_8919
		));
	notech_ao4 i_80806(.A(n_10158), .B(n_10078), .C(n_887), .D(n_10076), .Z(n_58106
		));
	notech_reg_set tab24_reg_29(.CP(n_61983), .D(n_8925), .SD(n_61268), .Q(\tab24[29] 
		));
	notech_mux2 i_12130(.S(n_60492), .A(\tab24[29] ), .B(n_57820), .Z(n_8925
		));
	notech_nand2 i_322380(.A(n_975), .B(n_400), .Z(addr_phys[2]));
	notech_reg_set tab24_reg_33(.CP(n_61983), .D(n_8931), .SD(n_61268), .Q(\tab24[33] 
		));
	notech_mux2 i_12138(.S(n_60492), .A(\tab24[33] ), .B(n_57844), .Z(n_8931
		));
	notech_nand2 i_422381(.A(n_976), .B(n_398), .Z(addr_phys[3]));
	notech_reg hit_adr24_reg(.CP(n_61983), .D(n_8937), .CD(n_61268), .Q(hit_adr24
		));
	notech_mux2 i_12146(.S(n_872), .A(hit_add24), .B(hit_adr24), .Z(n_8937)
		);
	notech_nand2 i_522382(.A(n_977), .B(n_397), .Z(addr_phys[4]));
	notech_reg_set nnx_tab2_reg_0(.CP(n_61983), .D(n_8943), .SD(n_61268), .Q
		(\nnx_tab2[0] ));
	notech_mux2 i_12154(.S(n_10008), .A(\nnx_tab2[0] ), .B(n_10004), .Z(n_8943
		));
	notech_nand2 i_622383(.A(n_978), .B(n_396), .Z(addr_phys[5]));
	notech_reg nnx_tab2_reg_1(.CP(n_61987), .D(n_8949), .CD(n_61272), .Q(\nnx_tab2[1] 
		));
	notech_mux2 i_12162(.S(n_10008), .A(\nnx_tab2[1] ), .B(n_10006), .Z(n_8949
		));
	notech_nand2 i_722384(.A(n_979), .B(n_395), .Z(addr_phys[6]));
	notech_reg nx_tab2_reg_0(.CP(n_61992), .D(n_8955), .CD(n_61277), .Q(\nx_tab2[0] 
		));
	notech_mux2 i_12170(.S(\nbus_14516[0] ), .A(\nx_tab2[0] ), .B(n_10009), 
		.Z(n_8955));
	notech_nand2 i_822385(.A(n_980), .B(n_394), .Z(addr_phys[7]));
	notech_reg nx_tab2_reg_1(.CP(n_61992), .D(n_8961), .CD(n_61277), .Q(\nx_tab2[1] 
		));
	notech_mux2 i_12178(.S(\nbus_14516[0] ), .A(\nx_tab2[1] ), .B(n_10011), 
		.Z(n_8961));
	notech_nand2 i_922386(.A(n_981), .B(n_393), .Z(addr_phys[8]));
	notech_reg_set tab11_reg_0(.CP(n_61992), .D(n_8967), .SD(n_61277), .Q(\tab11[0] 
		));
	notech_mux2 i_12186(.S(\nbus_14492[0] ), .A(\tab11[0] ), .B(n_57646), .Z
		(n_8967));
	notech_nand2 i_1022387(.A(n_982), .B(n_392), .Z(addr_phys[9]));
	notech_reg_set tab11_reg_1(.CP(n_61992), .D(n_8973), .SD(n_61277), .Q(\tab11[1] 
		));
	notech_mux2 i_12194(.S(\nbus_14492[0] ), .A(\tab11[1] ), .B(n_57652), .Z
		(n_8973));
	notech_nand2 i_1122388(.A(n_983), .B(n_391), .Z(addr_phys[10]));
	notech_reg_set tab11_reg_2(.CP(n_61988), .D(n_8979), .SD(n_61273), .Q(\tab11[2] 
		));
	notech_mux2 i_12202(.S(\nbus_14492[0] ), .A(\tab11[2] ), .B(n_57658), .Z
		(n_8979));
	notech_nand2 i_1222389(.A(n_984), .B(n_390), .Z(addr_phys[11]));
	notech_reg_set tab11_reg_3(.CP(n_61988), .D(n_8985), .SD(n_61273), .Q(\tab11[3] 
		));
	notech_mux2 i_12210(.S(\nbus_14492[0] ), .A(\tab11[3] ), .B(n_57664), .Z
		(n_8985));
	notech_and4 i_1322390(.A(n_1004), .B(n_1006), .C(n_1001), .D(n_773), .Z(addr_phys_12100141
		));
	notech_reg tab11_reg_4(.CP(n_61988), .D(n_8991), .CD(n_61273), .Q(\tab11[4] 
		));
	notech_mux2 i_12218(.S(\nbus_14492[0] ), .A(\tab11[4] ), .B(n_873), .Z(n_8991
		));
	notech_and4 i_1422391(.A(n_1013), .B(n_1015), .C(n_1012), .D(n_762), .Z(addr_phys_13100142
		));
	notech_reg_set tab11_reg_5(.CP(n_61992), .D(n_8997), .SD(n_61277), .Q(\tab11[5] 
		));
	notech_mux2 i_12226(.S(\nbus_14492[0] ), .A(\tab11[5] ), .B(n_57676), .Z
		(n_8997));
	notech_and4 i_1522392(.A(n_1022), .B(n_1024), .C(n_1021), .D(n_751), .Z(addr_phys_14100143
		));
	notech_reg_set tab11_reg_6(.CP(n_61992), .D(n_9003), .SD(n_61277), .Q(\tab11[6] 
		));
	notech_mux2 i_12234(.S(\nbus_14492[0] ), .A(\tab11[6] ), .B(n_57682), .Z
		(n_9003));
	notech_and4 i_1622393(.A(n_1031), .B(n_1033), .C(n_1030), .D(n_740), .Z(addr_phys_15100144
		));
	notech_reg_set tab11_reg_7(.CP(n_61992), .D(n_9009), .SD(n_61277), .Q(\tab11[7] 
		));
	notech_mux2 i_12242(.S(\nbus_14492[0] ), .A(\tab11[7] ), .B(n_57688), .Z
		(n_9009));
	notech_and4 i_1722394(.A(n_1040), .B(n_1042), .C(n_1039), .D(n_729), .Z(addr_phys_16100145
		));
	notech_reg_set tab11_reg_8(.CP(n_61992), .D(n_9015), .SD(n_61277), .Q(\tab11[8] 
		));
	notech_mux2 i_12250(.S(\nbus_14492[0] ), .A(\tab11[8] ), .B(n_57694), .Z
		(n_9015));
	notech_and4 i_1822395(.A(n_1049), .B(n_1051), .C(n_1048), .D(n_718), .Z(addr_phys_17100146
		));
	notech_reg_set tab11_reg_9(.CP(n_61992), .D(n_9021), .SD(n_61277), .Q(\tab11[9] 
		));
	notech_mux2 i_12258(.S(\nbus_14492[0] ), .A(\tab11[9] ), .B(n_57700), .Z
		(n_9021));
	notech_and4 i_1922396(.A(n_1058), .B(n_1060), .C(n_1057), .D(n_707), .Z(addr_phys_18100147
		));
	notech_reg_set tab11_reg_10(.CP(n_61992), .D(n_9027), .SD(n_61277), .Q(\tab11[10] 
		));
	notech_mux2 i_12266(.S(\nbus_14492[0] ), .A(\tab11[10] ), .B(n_57706), .Z
		(n_9027));
	notech_and4 i_2022397(.A(n_1067), .B(n_1069), .C(n_1066), .D(n_696), .Z(addr_phys_19100148
		));
	notech_reg_set tab11_reg_11(.CP(n_61992), .D(n_9033), .SD(n_61277), .Q(\tab11[11] 
		));
	notech_mux2 i_12274(.S(\nbus_14492[0] ), .A(\tab11[11] ), .B(n_57712), .Z
		(n_9033));
	notech_and4 i_2122398(.A(n_1076), .B(n_1078), .C(n_1075), .D(n_685), .Z(addr_phys_20100149
		));
	notech_reg_set tab11_reg_12(.CP(n_61988), .D(n_9039), .SD(n_61273), .Q(\tab11[12] 
		));
	notech_mux2 i_12282(.S(\nbus_14492[0] ), .A(\tab11[12] ), .B(n_57718), .Z
		(n_9039));
	notech_and4 i_2222399(.A(n_1085), .B(n_1087), .C(n_1084), .D(n_674), .Z(addr_phys_21100150
		));
	notech_reg_set tab11_reg_13(.CP(n_61988), .D(n_9045), .SD(n_61273), .Q(\tab11[13] 
		));
	notech_mux2 i_12290(.S(\nbus_14492[0] ), .A(\tab11[13] ), .B(n_57724), .Z
		(n_9045));
	notech_and4 i_2322400(.A(n_1094), .B(n_1096), .C(n_1093), .D(n_663), .Z(addr_phys_22100151
		));
	notech_reg_set tab11_reg_14(.CP(n_61988), .D(n_9051), .SD(n_61273), .Q(\tab11[14] 
		));
	notech_mux2 i_12298(.S(\nbus_14492[0] ), .A(\tab11[14] ), .B(n_57730), .Z
		(n_9051));
	notech_and4 i_2422401(.A(n_1103), .B(n_1105), .C(n_1102), .D(n_652), .Z(addr_phys_23100152
		));
	notech_reg_set tab11_reg_15(.CP(n_61988), .D(n_9057), .SD(n_61273), .Q(\tab11[15] 
		));
	notech_mux2 i_12306(.S(\nbus_14492[0] ), .A(\tab11[15] ), .B(n_57736), .Z
		(n_9057));
	notech_and4 i_2522402(.A(n_1112), .B(n_1114), .C(n_1111), .D(n_641), .Z(addr_phys_24100153
		));
	notech_reg_set tab11_reg_16(.CP(n_61988), .D(n_9063), .SD(n_61273), .Q(\tab11[16] 
		));
	notech_mux2 i_12314(.S(n_60448), .A(\tab11[16] ), .B(n_57742), .Z(n_9063
		));
	notech_and4 i_2622403(.A(n_1121), .B(n_1123), .C(n_1120), .D(n_630), .Z(addr_phys_25100154
		));
	notech_reg_set tab11_reg_17(.CP(n_61987), .D(n_9069), .SD(n_61272), .Q(\tab11[17] 
		));
	notech_mux2 i_12322(.S(n_60448), .A(\tab11[17] ), .B(n_57748), .Z(n_9069
		));
	notech_and4 i_2722404(.A(n_1130), .B(n_1132), .C(n_1129), .D(n_619), .Z(addr_phys_26100155
		));
	notech_reg_set tab11_reg_18(.CP(n_61987), .D(n_9075), .SD(n_61272), .Q(\tab11[18] 
		));
	notech_mux2 i_12330(.S(n_60448), .A(\tab11[18] ), .B(n_57754), .Z(n_9075
		));
	notech_and4 i_2822405(.A(n_1139), .B(n_1141), .C(n_1138), .D(n_608), .Z(addr_phys_27100156
		));
	notech_reg_set tab11_reg_19(.CP(n_61988), .D(n_9081), .SD(n_61273), .Q(\tab11[19] 
		));
	notech_mux2 i_12338(.S(n_60448), .A(\tab11[19] ), .B(n_57760), .Z(n_9081
		));
	notech_and4 i_2922406(.A(n_1148), .B(n_1150), .C(n_1147), .D(n_597), .Z(addr_phys_28100157
		));
	notech_reg_set tab11_reg_20(.CP(n_61988), .D(n_9087), .SD(n_61273), .Q(\tab11[20] 
		));
	notech_mux2 i_12346(.S(n_60448), .A(\tab11[20] ), .B(n_57766), .Z(n_9087
		));
	notech_and4 i_3022407(.A(n_1157), .B(n_1159), .C(n_1156), .D(n_586), .Z(addr_phys_29100158
		));
	notech_reg_set tab11_reg_21(.CP(n_61988), .D(n_9093), .SD(n_61273), .Q(\tab11[21] 
		));
	notech_mux2 i_12354(.S(n_60448), .A(\tab11[21] ), .B(n_57772), .Z(n_9093
		));
	notech_and4 i_3122408(.A(n_1166), .B(n_1168), .C(n_1165), .D(n_575), .Z(addr_phys_30100159
		));
	notech_reg_set tab11_reg_22(.CP(n_61988), .D(n_9099), .SD(n_61273), .Q(\tab11[22] 
		));
	notech_mux2 i_12362(.S(n_60448), .A(\tab11[22] ), .B(n_57778), .Z(n_9099
		));
	notech_and4 i_3222409(.A(n_1175), .B(n_1177), .C(n_1174), .D(n_564), .Z(addr_phys_31100160
		));
	notech_reg_set tab11_reg_23(.CP(n_61988), .D(n_9105), .SD(n_61273), .Q(\tab11[23] 
		));
	notech_mux2 i_12370(.S(n_60448), .A(\tab11[23] ), .B(n_57784), .Z(n_9105
		));
	notech_mux2 i_122920(.S(n_61917), .A(iDaddr[12]), .B(iDaddr_f[12]), .Z(\tab11_0[0] 
		));
	notech_reg_set tab11_reg_24(.CP(n_61988), .D(n_9111), .SD(n_61273), .Q(\tab11[24] 
		));
	notech_mux2 i_12378(.S(n_60448), .A(\tab11[24] ), .B(n_57790), .Z(n_9111
		));
	notech_mux2 i_222921(.S(n_61917), .A(iDaddr[13]), .B(iDaddr_f[13]), .Z(\tab11_0[1] 
		));
	notech_reg_set tab11_reg_25(.CP(n_61988), .D(n_9117), .SD(n_61273), .Q(\tab11[25] 
		));
	notech_mux2 i_12386(.S(n_60448), .A(\tab11[25] ), .B(n_57796), .Z(n_9117
		));
	notech_mux2 i_322922(.S(n_61917), .A(iDaddr[14]), .B(iDaddr_f[14]), .Z(\tab11_0[2] 
		));
	notech_reg_set tab11_reg_26(.CP(n_61988), .D(n_9123), .SD(n_61273), .Q(\tab11[26] 
		));
	notech_mux2 i_12394(.S(n_60448), .A(\tab11[26] ), .B(n_57802), .Z(n_9123
		));
	notech_mux2 i_422923(.S(n_61917), .A(iDaddr[15]), .B(iDaddr_f[15]), .Z(\tab11_0[3] 
		));
	notech_reg_set tab11_reg_27(.CP(n_62005), .D(n_9129), .SD(n_61290), .Q(\tab11[27] 
		));
	notech_mux2 i_12402(.S(n_60448), .A(\tab11[27] ), .B(n_57808), .Z(n_9129
		));
	notech_mux2 i_522924(.S(n_61917), .A(iDaddr[16]), .B(iDaddr_f[16]), .Z(\tab11_0[4] 
		));
	notech_reg_set tab11_reg_28(.CP(n_62016), .D(n_9135), .SD(n_61301), .Q(\tab11[28] 
		));
	notech_mux2 i_12410(.S(n_60448), .A(\tab11[28] ), .B(n_57814), .Z(n_9135
		));
	notech_mux2 i_622925(.S(n_61917), .A(iDaddr[17]), .B(iDaddr_f[17]), .Z(\tab11_0[5] 
		));
	notech_reg_set tab11_reg_29(.CP(n_62016), .D(n_9141), .SD(n_61301), .Q(\tab11[29] 
		));
	notech_mux2 i_12418(.S(n_60448), .A(\tab11[29] ), .B(n_57820), .Z(n_9141
		));
	notech_mux2 i_722926(.S(n_61917), .A(iDaddr[18]), .B(iDaddr_f[18]), .Z(\tab11_0[6] 
		));
	notech_reg_set tab11_reg_33(.CP(n_62016), .D(n_9147), .SD(n_61301), .Q(\tab11[33] 
		));
	notech_mux2 i_12426(.S(n_60448), .A(\tab11[33] ), .B(n_57844), .Z(n_9147
		));
	notech_mux2 i_822927(.S(n_61917), .A(iDaddr[19]), .B(iDaddr_f[19]), .Z(\tab11_0[7] 
		));
	notech_reg fsm5_cnt_reg_0(.CP(n_62016), .D(n_9153), .CD(n_61301), .Q(fsm5_cnt
		[0]));
	notech_mux2 i_12434(.S(\nbus_14499[0] ), .A(fsm5_cnt[0]), .B(n_863), .Z(n_9153
		));
	notech_mux2 i_922928(.S(n_61917), .A(iDaddr[20]), .B(iDaddr_f[20]), .Z(\tab11_0[8] 
		));
	notech_reg fsm5_cnt_reg_1(.CP(n_62016), .D(n_9159), .CD(n_61301), .Q(fsm5_cnt
		[1]));
	notech_mux2 i_12442(.S(\nbus_14499[0] ), .A(fsm5_cnt[1]), .B(n_864), .Z(n_9159
		));
	notech_mux2 i_1022929(.S(n_61917), .A(iDaddr[21]), .B(iDaddr_f[21]), .Z(\tab11_0[9] 
		));
	notech_reg fsm5_cnt_reg_2(.CP(n_62016), .D(n_9165), .CD(n_61301), .Q(fsm5_cnt
		[2]));
	notech_mux2 i_12450(.S(\nbus_14499[0] ), .A(fsm5_cnt[2]), .B(n_865), .Z(n_9165
		));
	notech_mux2 i_1122930(.S(n_61922), .A(iDaddr[22]), .B(iDaddr_f[22]), .Z(\dir1_0[0] 
		));
	notech_reg fsm5_cnt_reg_3(.CP(n_62016), .D(n_9171), .CD(n_61301), .Q(fsm5_cnt
		[3]));
	notech_mux2 i_12458(.S(\nbus_14499[0] ), .A(fsm5_cnt[3]), .B(n_866), .Z(n_9171
		));
	notech_mux2 i_1222931(.S(n_61922), .A(iDaddr[23]), .B(iDaddr_f[23]), .Z(\dir1_0[1] 
		));
	notech_reg fsm5_cnt_reg_4(.CP(n_62016), .D(n_9177), .CD(n_61301), .Q(fsm5_cnt
		[4]));
	notech_mux2 i_12466(.S(\nbus_14499[0] ), .A(fsm5_cnt[4]), .B(n_867), .Z(n_9177
		));
	notech_mux2 i_1322932(.S(n_61922), .A(iDaddr[24]), .B(iDaddr_f[24]), .Z(\dir1_0[2] 
		));
	notech_reg fsm5_cnt_reg_5(.CP(n_62020), .D(n_9183), .CD(n_61305), .Q(fsm5_cnt
		[5]));
	notech_mux2 i_12474(.S(\nbus_14499[0] ), .A(fsm5_cnt[5]), .B(n_868), .Z(n_9183
		));
	notech_mux2 i_1422933(.S(n_61922), .A(iDaddr[25]), .B(iDaddr_f[25]), .Z(\dir1_0[3] 
		));
	notech_reg fsm5_cnt_reg_6(.CP(n_62020), .D(n_9189), .CD(n_61305), .Q(fsm5_cnt
		[6]));
	notech_mux2 i_12482(.S(\nbus_14499[0] ), .A(fsm5_cnt[6]), .B(n_869), .Z(n_9189
		));
	notech_mux2 i_1522934(.S(n_61922), .A(iDaddr[26]), .B(iDaddr_f[26]), .Z(\dir1_0[4] 
		));
	notech_reg fsm5_cnt_reg_7(.CP(n_62016), .D(n_9195), .CD(n_61301), .Q(fsm5_cnt
		[7]));
	notech_mux2 i_12490(.S(\nbus_14499[0] ), .A(fsm5_cnt[7]), .B(n_870), .Z(n_9195
		));
	notech_mux2 i_1622935(.S(n_61922), .A(iDaddr[27]), .B(iDaddr_f[27]), .Z(\dir1_0[5] 
		));
	notech_reg fsm5_cnt_reg_8(.CP(n_62016), .D(n_9201), .CD(n_61301), .Q(fsm5_cnt
		[8]));
	notech_mux2 i_12498(.S(\nbus_14499[0] ), .A(fsm5_cnt[8]), .B(n_871), .Z(n_9201
		));
	notech_mux2 i_1722936(.S(n_61922), .A(iDaddr[28]), .B(iDaddr_f[28]), .Z(\dir1_0[6] 
		));
	notech_reg pg_fault_reg(.CP(n_62016), .D(n_9207), .CD(n_61301), .Q(pg_fault
		));
	notech_mux2 i_12506(.S(n_10033), .A(pg_fault), .B(n_862), .Z(n_9207));
	notech_mux2 i_1822937(.S(n_61922), .A(iDaddr[29]), .B(iDaddr_f[29]), .Z(\dir1_0[7] 
		));
	notech_reg fsm_reg_0(.CP(n_62016), .D(n_9213), .CD(n_61301), .Q(fsm[0])
		);
	notech_mux2 i_12514(.S(\nbus_14493[0] ), .A(n_61926), .B(n_58079), .Z(n_9213
		));
	notech_mux2 i_1922938(.S(n_61922), .A(iDaddr[30]), .B(iDaddr_f[30]), .Z(\dir1_0[8] 
		));
	notech_reg fsm_reg_1(.CP(n_62016), .D(n_9219), .CD(n_61301), .Q(fsm[1])
		);
	notech_mux2 i_12522(.S(\nbus_14493[0] ), .A(fsm[1]), .B(n_58085), .Z(n_9219
		));
	notech_mux2 i_2022939(.S(n_61922), .A(iDaddr[31]), .B(iDaddr_f[31]), .Z(\dir1_0[9] 
		));
	notech_reg fsm_reg_2(.CP(n_62015), .D(n_9225), .CD(n_61300), .Q(fsm[2])
		);
	notech_mux2 i_12530(.S(\nbus_14493[0] ), .A(fsm[2]), .B(n_58091), .Z(n_9225
		));
	notech_nand3 i_79271(.A(n_60814), .B(n_61922), .C(n_10142), .Z(n_57422)
		);
	notech_reg fsm_reg_3(.CP(n_62015), .D(n_9231), .CD(n_61300), .Q(fsm[3])
		);
	notech_mux2 i_12538(.S(\nbus_14493[0] ), .A(fsm[3]), .B(n_861), .Z(n_9231
		));
	notech_nand3 i_79273(.A(n_60814), .B(n_61922), .C(n_10141), .Z(n_57428)
		);
	notech_reg addr_miss_reg_2(.CP(n_62015), .D(n_9237), .CD(n_61300), .Q(\addr_miss[2] 
		));
	notech_mux2 i_12546(.S(n_853), .A(n_10036), .B(\addr_miss[2] ), .Z(n_9237
		));
	notech_nand3 i_79275(.A(n_60814), .B(n_61920), .C(n_10140), .Z(n_57434)
		);
	notech_reg addr_miss_reg_3(.CP(n_62015), .D(n_9243), .CD(n_61300), .Q(\addr_miss[3] 
		));
	notech_mux2 i_12554(.S(n_853), .A(n_10037), .B(\addr_miss[3] ), .Z(n_9243
		));
	notech_nand3 i_79277(.A(n_60814), .B(n_61920), .C(n_10139), .Z(n_57440)
		);
	notech_reg addr_miss_reg_4(.CP(n_62015), .D(n_9249), .CD(n_61300), .Q(\addr_miss[4] 
		));
	notech_mux2 i_12562(.S(n_853), .A(n_10038), .B(\addr_miss[4] ), .Z(n_9249
		));
	notech_nand3 i_79281(.A(n_60814), .B(n_61920), .C(n_10137), .Z(n_57452)
		);
	notech_reg addr_miss_reg_5(.CP(n_62015), .D(n_9255), .CD(n_61300), .Q(\addr_miss[5] 
		));
	notech_mux2 i_12570(.S(n_853), .A(n_10039), .B(\addr_miss[5] ), .Z(n_9255
		));
	notech_nand3 i_79283(.A(n_60814), .B(n_61920), .C(n_10136), .Z(n_57458)
		);
	notech_reg addr_miss_reg_6(.CP(n_62015), .D(n_9261), .CD(n_61300), .Q(\addr_miss[6] 
		));
	notech_mux2 i_12578(.S(n_853), .A(n_10040), .B(\addr_miss[6] ), .Z(n_9261
		));
	notech_nand3 i_79285(.A(n_60814), .B(n_61920), .C(n_10135), .Z(n_57464)
		);
	notech_reg addr_miss_reg_7(.CP(n_62016), .D(n_9267), .CD(n_61301), .Q(\addr_miss[7] 
		));
	notech_mux2 i_12586(.S(n_853), .A(n_10041), .B(\addr_miss[7] ), .Z(n_9267
		));
	notech_nand3 i_79287(.A(n_60814), .B(n_61920), .C(n_10134), .Z(n_57470)
		);
	notech_reg addr_miss_reg_8(.CP(n_62016), .D(n_9273), .CD(n_61301), .Q(\addr_miss[8] 
		));
	notech_mux2 i_12594(.S(n_853), .A(n_10042), .B(\addr_miss[8] ), .Z(n_9273
		));
	notech_nand3 i_79289(.A(n_60814), .B(n_61922), .C(n_10133), .Z(n_57476)
		);
	notech_reg addr_miss_reg_9(.CP(n_62016), .D(n_9279), .CD(n_61301), .Q(\addr_miss[9] 
		));
	notech_mux2 i_12602(.S(n_853), .A(n_10043), .B(\addr_miss[9] ), .Z(n_9279
		));
	notech_nao3 i_79291(.A(n_61922), .B(n_60814), .C(data_miss[12]), .Z(n_57482
		));
	notech_reg addr_miss_reg_10(.CP(n_62016), .D(n_9285), .CD(n_61301), .Q(\addr_miss[10] 
		));
	notech_mux2 i_12610(.S(n_853), .A(n_10044), .B(\addr_miss[10] ), .Z(n_9285
		));
	notech_nao3 i_79293(.A(n_61922), .B(n_60814), .C(data_miss[13]), .Z(n_57488
		));
	notech_reg addr_miss_reg_11(.CP(n_62015), .D(n_9291), .CD(n_61300), .Q(\addr_miss[11] 
		));
	notech_mux2 i_12618(.S(n_853), .A(n_10045), .B(\addr_miss[11] ), .Z(n_9291
		));
	notech_nao3 i_79295(.A(n_61920), .B(n_60814), .C(data_miss[14]), .Z(n_57494
		));
	notech_reg addr_miss_reg_12(.CP(n_62015), .D(n_9297), .CD(n_61300), .Q(\addr_miss[12] 
		));
	notech_mux2 i_12626(.S(n_853), .A(n_59590), .B(\addr_miss[12] ), .Z(n_9297
		));
	notech_nao3 i_79297(.A(n_61922), .B(n_60814), .C(data_miss[15]), .Z(n_57500
		));
	notech_reg addr_miss_reg_13(.CP(n_62016), .D(n_9303), .CD(n_61301), .Q(\addr_miss[13] 
		));
	notech_mux2 i_12634(.S(n_853), .A(n_59596), .B(\addr_miss[13] ), .Z(n_9303
		));
	notech_nao3 i_79299(.A(n_61917), .B(n_60810), .C(data_miss[16]), .Z(n_57506
		));
	notech_reg addr_miss_reg_14(.CP(n_62020), .D(n_9309), .CD(n_61305), .Q(\addr_miss[14] 
		));
	notech_mux2 i_12642(.S(n_853), .A(n_59602), .B(\addr_miss[14] ), .Z(n_9309
		));
	notech_nao3 i_79301(.A(n_61912), .B(n_60810), .C(data_miss[17]), .Z(n_57512
		));
	notech_reg addr_miss_reg_15(.CP(n_62024), .D(n_9315), .CD(n_61309), .Q(\addr_miss[15] 
		));
	notech_mux2 i_12650(.S(n_853), .A(n_59608), .B(\addr_miss[15] ), .Z(n_9315
		));
	notech_nao3 i_79303(.A(n_61912), .B(n_60810), .C(data_miss[18]), .Z(n_57518
		));
	notech_reg addr_miss_reg_16(.CP(n_62024), .D(n_9321), .CD(n_61309), .Q(\addr_miss[16] 
		));
	notech_mux2 i_12658(.S(n_853), .A(n_59614), .B(\addr_miss[16] ), .Z(n_9321
		));
	notech_nao3 i_79305(.A(n_61912), .B(n_60810), .C(data_miss[19]), .Z(n_57524
		));
	notech_reg addr_miss_reg_17(.CP(n_62024), .D(n_9327), .CD(n_61309), .Q(\addr_miss[17] 
		));
	notech_mux2 i_12666(.S(n_60819), .A(n_59620), .B(\addr_miss[17] ), .Z(n_9327
		));
	notech_nao3 i_79307(.A(n_61910), .B(n_60810), .C(data_miss[20]), .Z(n_57530
		));
	notech_reg addr_miss_reg_18(.CP(n_62024), .D(n_9333), .CD(n_61309), .Q(\addr_miss[18] 
		));
	notech_mux2 i_12674(.S(n_60819), .A(n_59626), .B(\addr_miss[18] ), .Z(n_9333
		));
	notech_nao3 i_79309(.A(n_61910), .B(n_60810), .C(data_miss[21]), .Z(n_57536
		));
	notech_reg addr_miss_reg_19(.CP(n_62024), .D(n_9339), .CD(n_61309), .Q(\addr_miss[19] 
		));
	notech_mux2 i_12682(.S(n_60819), .A(n_59632), .B(\addr_miss[19] ), .Z(n_9339
		));
	notech_nao3 i_79311(.A(n_61912), .B(n_60810), .C(data_miss[22]), .Z(n_57542
		));
	notech_reg addr_miss_reg_20(.CP(n_62024), .D(n_9345), .CD(n_61309), .Q(\addr_miss[20] 
		));
	notech_mux2 i_12690(.S(n_60819), .A(n_59638), .B(\addr_miss[20] ), .Z(n_9345
		));
	notech_nao3 i_79313(.A(n_61912), .B(n_60810), .C(data_miss[23]), .Z(n_57548
		));
	notech_reg addr_miss_reg_21(.CP(n_62024), .D(n_9351), .CD(n_61309), .Q(\addr_miss[21] 
		));
	notech_mux2 i_12698(.S(n_60819), .A(n_59644), .B(\addr_miss[21] ), .Z(n_9351
		));
	notech_nao3 i_79315(.A(n_61912), .B(n_60810), .C(data_miss[24]), .Z(n_57554
		));
	notech_reg addr_miss_reg_22(.CP(n_62024), .D(n_9357), .CD(n_61309), .Q(\addr_miss[22] 
		));
	notech_mux2 i_12706(.S(n_60819), .A(n_59650), .B(\addr_miss[22] ), .Z(n_9357
		));
	notech_nao3 i_79317(.A(n_61912), .B(n_60810), .C(data_miss[25]), .Z(n_57560
		));
	notech_reg addr_miss_reg_23(.CP(n_62024), .D(n_9363), .CD(n_61309), .Q(\addr_miss[23] 
		));
	notech_mux2 i_12714(.S(n_60819), .A(n_59656), .B(\addr_miss[23] ), .Z(n_9363
		));
	notech_nao3 i_79319(.A(n_61912), .B(n_60810), .C(data_miss[26]), .Z(n_57566
		));
	notech_reg addr_miss_reg_24(.CP(n_62024), .D(n_9369), .CD(n_61309), .Q(\addr_miss[24] 
		));
	notech_mux2 i_12722(.S(n_60819), .A(n_59662), .B(\addr_miss[24] ), .Z(n_9369
		));
	notech_nao3 i_79321(.A(n_61912), .B(n_60810), .C(data_miss[27]), .Z(n_57572
		));
	notech_reg addr_miss_reg_25(.CP(n_62024), .D(n_9375), .CD(n_61309), .Q(\addr_miss[25] 
		));
	notech_mux2 i_12730(.S(n_60819), .A(n_59668), .B(\addr_miss[25] ), .Z(n_9375
		));
	notech_nao3 i_79323(.A(n_61910), .B(n_60810), .C(data_miss[28]), .Z(n_57578
		));
	notech_reg addr_miss_reg_26(.CP(n_62024), .D(n_9381), .CD(n_61309), .Q(\addr_miss[26] 
		));
	notech_mux2 i_12738(.S(n_60819), .A(n_59674), .B(\addr_miss[26] ), .Z(n_9381
		));
	notech_nao3 i_79325(.A(n_61910), .B(n_60810), .C(data_miss[29]), .Z(n_57584
		));
	notech_reg addr_miss_reg_27(.CP(n_62024), .D(n_9387), .CD(n_61309), .Q(\addr_miss[27] 
		));
	notech_mux2 i_12746(.S(n_60819), .A(n_59680), .B(\addr_miss[27] ), .Z(n_9387
		));
	notech_nao3 i_79327(.A(n_61910), .B(n_60810), .C(data_miss[30]), .Z(n_57590
		));
	notech_reg addr_miss_reg_28(.CP(n_62024), .D(n_9393), .CD(n_61309), .Q(\addr_miss[28] 
		));
	notech_mux2 i_12754(.S(n_60819), .A(n_59686), .B(\addr_miss[28] ), .Z(n_9393
		));
	notech_nao3 i_79329(.A(n_61910), .B(n_60810), .C(data_miss[31]), .Z(n_57596
		));
	notech_reg addr_miss_reg_29(.CP(n_62020), .D(n_9399), .CD(n_61305), .Q(\addr_miss[29] 
		));
	notech_mux2 i_12762(.S(n_60819), .A(n_59692), .B(\addr_miss[29] ), .Z(n_9399
		));
	notech_nand2 i_79335(.A(n_61910), .B(n_60810), .Z(n_57621));
	notech_reg addr_miss_reg_30(.CP(n_62020), .D(n_9405), .CD(n_61305), .Q(\addr_miss[30] 
		));
	notech_mux2 i_12770(.S(n_60819), .A(n_59698), .B(\addr_miss[30] ), .Z(n_9405
		));
	notech_nand2 i_79572(.A(n_896), .B(n_890), .Z(n_58203));
	notech_reg addr_miss_reg_31(.CP(n_62020), .D(n_9411), .CD(n_61305), .Q(\addr_miss[31] 
		));
	notech_mux2 i_12778(.S(n_60819), .A(n_59704), .B(\addr_miss[31] ), .Z(n_9411
		));
	notech_ao4 i_79465(.A(n_938), .B(n_10142), .C(n_916), .D(n_10152), .Z(n_59530
		));
	notech_reg wrA_reg_2(.CP(n_62020), .D(n_9417), .CD(n_61305), .Q(\wrA[2] 
		));
	notech_mux2 i_12786(.S(n_60401), .A(\wrA[2] ), .B(\addr_miss[2] ), .Z(n_9417
		));
	notech_ao4 i_79468(.A(n_938), .B(n_10141), .C(n_916), .D(n_10151), .Z(n_59536
		));
	notech_reg wrA_reg_3(.CP(n_62020), .D(n_9423), .CD(n_61305), .Q(\wrA[3] 
		));
	notech_mux2 i_12794(.S(n_60401), .A(\wrA[3] ), .B(\addr_miss[3] ), .Z(n_9423
		));
	notech_ao4 i_79471(.A(n_938), .B(n_10140), .C(n_916), .D(n_10150), .Z(n_59542
		));
	notech_reg wrA_reg_4(.CP(n_62020), .D(n_9429), .CD(n_61305), .Q(\wrA[4] 
		));
	notech_mux2 i_12802(.S(n_60401), .A(\wrA[4] ), .B(\addr_miss[4] ), .Z(n_9429
		));
	notech_ao4 i_79474(.A(n_938), .B(n_10139), .C(n_916), .D(n_10149), .Z(n_59548
		));
	notech_reg wrA_reg_5(.CP(n_62020), .D(n_9435), .CD(n_61305), .Q(\wrA[5] 
		));
	notech_mux2 i_12810(.S(n_60401), .A(\wrA[5] ), .B(\addr_miss[5] ), .Z(n_9435
		));
	notech_ao4 i_79477(.A(n_938), .B(n_10138), .C(n_916), .D(n_10148), .Z(n_59554
		));
	notech_reg wrA_reg_6(.CP(n_62020), .D(n_9441), .CD(n_61305), .Q(\wrA[6] 
		));
	notech_mux2 i_12818(.S(n_60401), .A(\wrA[6] ), .B(\addr_miss[6] ), .Z(n_9441
		));
	notech_ao4 i_79480(.A(n_938), .B(n_10137), .C(n_916), .D(n_10147), .Z(n_59560
		));
	notech_reg wrA_reg_7(.CP(n_62020), .D(n_9447), .CD(n_61305), .Q(\wrA[7] 
		));
	notech_mux2 i_12826(.S(n_60401), .A(\wrA[7] ), .B(\addr_miss[7] ), .Z(n_9447
		));
	notech_ao4 i_79483(.A(n_938), .B(n_10136), .C(n_916), .D(n_10146), .Z(n_59566
		));
	notech_reg wrA_reg_8(.CP(n_62020), .D(n_9453), .CD(n_61305), .Q(\wrA[8] 
		));
	notech_mux2 i_12834(.S(n_60401), .A(\wrA[8] ), .B(\addr_miss[8] ), .Z(n_9453
		));
	notech_ao4 i_79486(.A(n_938), .B(n_10135), .C(n_916), .D(n_10145), .Z(n_59572
		));
	notech_reg wrA_reg_9(.CP(n_62020), .D(n_9459), .CD(n_61305), .Q(\wrA[9] 
		));
	notech_mux2 i_12842(.S(n_60401), .A(\wrA[9] ), .B(\addr_miss[9] ), .Z(n_9459
		));
	notech_ao4 i_79489(.A(n_938), .B(n_10134), .C(n_916), .D(n_10144), .Z(n_59578
		));
	notech_reg wrA_reg_10(.CP(n_62020), .D(n_9465), .CD(n_61305), .Q(\wrA[10] 
		));
	notech_mux2 i_12850(.S(n_60401), .A(\wrA[10] ), .B(\addr_miss[10] ), .Z(n_9465
		));
	notech_ao4 i_79492(.A(n_938), .B(n_10133), .C(n_916), .D(n_10143), .Z(n_59584
		));
	notech_reg wrA_reg_11(.CP(n_62020), .D(n_9471), .CD(n_61305), .Q(\wrA[11] 
		));
	notech_mux2 i_12858(.S(n_60401), .A(\wrA[11] ), .B(\addr_miss[11] ), .Z(n_9471
		));
	notech_nand2 i_79495(.A(n_970), .B(n_424), .Z(n_59590));
	notech_reg wrA_reg_12(.CP(n_62020), .D(n_9477), .CD(n_61305), .Q(\wrA[12] 
		));
	notech_mux2 i_12866(.S(n_60401), .A(\wrA[12] ), .B(\addr_miss[12] ), .Z(n_9477
		));
	notech_nand2 i_79498(.A(n_969), .B(n_425), .Z(n_59596));
	notech_reg wrA_reg_13(.CP(n_62020), .D(n_9483), .CD(n_61305), .Q(\wrA[13] 
		));
	notech_mux2 i_12874(.S(n_60401), .A(\wrA[13] ), .B(\addr_miss[13] ), .Z(n_9483
		));
	notech_nand2 i_79501(.A(n_968), .B(n_426), .Z(n_59602));
	notech_reg wrA_reg_14(.CP(n_62006), .D(n_9489), .CD(n_61291), .Q(\wrA[14] 
		));
	notech_mux2 i_12882(.S(n_60401), .A(\wrA[14] ), .B(\addr_miss[14] ), .Z(n_9489
		));
	notech_nand2 i_79504(.A(n_967), .B(n_427), .Z(n_59608));
	notech_reg wrA_reg_15(.CP(n_62006), .D(n_9495), .CD(n_61291), .Q(\wrA[15] 
		));
	notech_mux2 i_12890(.S(n_60401), .A(\wrA[15] ), .B(\addr_miss[15] ), .Z(n_9495
		));
	notech_nand2 i_79507(.A(n_966), .B(n_428), .Z(n_59614));
	notech_reg wrA_reg_16(.CP(n_62006), .D(n_9501), .CD(n_61291), .Q(\wrA[16] 
		));
	notech_mux2 i_12898(.S(n_60401), .A(\wrA[16] ), .B(\addr_miss[16] ), .Z(n_9501
		));
	notech_nand2 i_79510(.A(n_965), .B(n_429), .Z(n_59620));
	notech_reg wrA_reg_17(.CP(n_62006), .D(n_9507), .CD(n_61291), .Q(\wrA[17] 
		));
	notech_mux2 i_12906(.S(n_60401), .A(\wrA[17] ), .B(\addr_miss[17] ), .Z(n_9507
		));
	notech_nand2 i_79513(.A(n_964), .B(n_430), .Z(n_59626));
	notech_reg wrA_reg_18(.CP(n_62006), .D(n_9513), .CD(n_61291), .Q(\wrA[18] 
		));
	notech_mux2 i_12914(.S(n_60401), .A(\wrA[18] ), .B(\addr_miss[18] ), .Z(n_9513
		));
	notech_nand2 i_79516(.A(n_963), .B(n_431), .Z(n_59632));
	notech_reg wrA_reg_19(.CP(n_62006), .D(n_9519), .CD(n_61291), .Q(\wrA[19] 
		));
	notech_mux2 i_12922(.S(n_60401), .A(\wrA[19] ), .B(\addr_miss[19] ), .Z(n_9519
		));
	notech_nand2 i_79519(.A(n_962), .B(n_432), .Z(n_59638));
	notech_reg wrA_reg_20(.CP(n_62006), .D(n_9525), .CD(n_61291), .Q(\wrA[20] 
		));
	notech_mux2 i_12930(.S(n_60401), .A(\wrA[20] ), .B(\addr_miss[20] ), .Z(n_9525
		));
	notech_nand2 i_79522(.A(n_961), .B(n_433), .Z(n_59644));
	notech_reg wrA_reg_21(.CP(n_62006), .D(n_9531), .CD(n_61291), .Q(\wrA[21] 
		));
	notech_mux2 i_12938(.S(n_60396), .A(\wrA[21] ), .B(\addr_miss[21] ), .Z(n_9531
		));
	notech_nand2 i_79525(.A(n_960), .B(n_434), .Z(n_59650));
	notech_reg wrA_reg_22(.CP(n_62006), .D(n_9537), .CD(n_61291), .Q(\wrA[22] 
		));
	notech_mux2 i_12946(.S(n_60396), .A(\wrA[22] ), .B(\addr_miss[22] ), .Z(n_9537
		));
	notech_nand2 i_79528(.A(n_959), .B(n_435), .Z(n_59656));
	notech_reg wrA_reg_23(.CP(n_62006), .D(n_9543), .CD(n_61291), .Q(\wrA[23] 
		));
	notech_mux2 i_12954(.S(n_60396), .A(\wrA[23] ), .B(\addr_miss[23] ), .Z(n_9543
		));
	notech_nand2 i_79531(.A(n_958), .B(n_436), .Z(n_59662));
	notech_reg wrA_reg_24(.CP(n_62006), .D(n_9549), .CD(n_61291), .Q(\wrA[24] 
		));
	notech_mux2 i_12962(.S(n_60396), .A(\wrA[24] ), .B(\addr_miss[24] ), .Z(n_9549
		));
	notech_nand2 i_79534(.A(n_957), .B(n_437), .Z(n_59668));
	notech_reg wrA_reg_25(.CP(n_62006), .D(n_9555), .CD(n_61291), .Q(\wrA[25] 
		));
	notech_mux2 i_12970(.S(n_60396), .A(\wrA[25] ), .B(\addr_miss[25] ), .Z(n_9555
		));
	notech_nand2 i_79537(.A(n_956), .B(n_438), .Z(n_59674));
	notech_reg wrA_reg_26(.CP(n_62006), .D(n_9561), .CD(n_61291), .Q(\wrA[26] 
		));
	notech_mux2 i_12978(.S(n_60396), .A(\wrA[26] ), .B(\addr_miss[26] ), .Z(n_9561
		));
	notech_nand2 i_79540(.A(n_955), .B(n_439), .Z(n_59680));
	notech_reg wrA_reg_27(.CP(n_62006), .D(n_9567), .CD(n_61291), .Q(\wrA[27] 
		));
	notech_mux2 i_12986(.S(n_60396), .A(\wrA[27] ), .B(\addr_miss[27] ), .Z(n_9567
		));
	notech_nand2 i_79543(.A(n_954), .B(n_440), .Z(n_59686));
	notech_reg wrA_reg_28(.CP(n_62006), .D(n_9573), .CD(n_61291), .Q(\wrA[28] 
		));
	notech_mux2 i_12994(.S(n_60396), .A(\wrA[28] ), .B(\addr_miss[28] ), .Z(n_9573
		));
	notech_nand2 i_79546(.A(n_953), .B(n_441), .Z(n_59692));
	notech_reg wrA_reg_29(.CP(n_62005), .D(n_9579), .CD(n_61290), .Q(\wrA[29] 
		));
	notech_mux2 i_13002(.S(n_60396), .A(\wrA[29] ), .B(\addr_miss[29] ), .Z(n_9579
		));
	notech_nand2 i_79549(.A(n_952), .B(n_442), .Z(n_59698));
	notech_reg wrA_reg_30(.CP(n_62005), .D(n_9585), .CD(n_61290), .Q(\wrA[30] 
		));
	notech_mux2 i_13010(.S(n_60396), .A(\wrA[30] ), .B(\addr_miss[30] ), .Z(n_9585
		));
	notech_nand2 i_79552(.A(n_951), .B(n_443), .Z(n_59704));
	notech_reg wrA_reg_31(.CP(n_62005), .D(n_9591), .CD(n_61290), .Q(\wrA[31] 
		));
	notech_mux2 i_13018(.S(n_60396), .A(\wrA[31] ), .B(\addr_miss[31] ), .Z(n_9591
		));
	notech_ao4 i_79935(.A(n_916), .B(n_9955), .C(n_896), .D(\nnx_tab1[0] ), 
		.Z(n_57173));
	notech_reg wrD_reg_0(.CP(n_62005), .D(n_9597), .CD(n_61290), .Q(\wrD[0] 
		));
	notech_mux2 i_13026(.S(n_60396), .A(\wrD[0] ), .B(n_58203), .Z(n_9597)
		);
	notech_ao4 i_79938(.A(n_916), .B(n_9957), .C(n_896), .D(n_490), .Z(n_57179
		));
	notech_reg wrD_reg_1(.CP(n_62005), .D(n_9603), .CD(n_61290), .Q(\wrD[1] 
		));
	notech_mux2 i_13034(.S(n_60401), .A(\wrD[1] ), .B(data_miss[1]), .Z(n_9603
		));
	notech_nand3 i_80078(.A(n_890), .B(n_61910), .C(n_10152), .Z(n_57646));
	notech_reg wrD_reg_2(.CP(n_62005), .D(n_9609), .CD(n_61290), .Q(\wrD[2] 
		));
	notech_mux2 i_13042(.S(n_60396), .A(\wrD[2] ), .B(data_miss[2]), .Z(n_9609
		));
	notech_nand3 i_80080(.A(n_890), .B(n_61910), .C(n_10151), .Z(n_57652));
	notech_reg wrD_reg_3(.CP(n_62005), .D(n_9615), .CD(n_61290), .Q(\wrD[3] 
		));
	notech_mux2 i_13050(.S(n_60396), .A(\wrD[3] ), .B(data_miss[3]), .Z(n_9615
		));
	notech_nand3 i_80082(.A(n_890), .B(n_61910), .C(n_10150), .Z(n_57658));
	notech_reg wrD_reg_4(.CP(n_62005), .D(n_9621), .CD(n_61290), .Q(\wrD[4] 
		));
	notech_mux2 i_13058(.S(n_60396), .A(\wrD[4] ), .B(data_miss[4]), .Z(n_9621
		));
	notech_nand3 i_80084(.A(n_890), .B(n_61910), .C(n_10149), .Z(n_57664));
	notech_reg wrD_reg_5(.CP(n_62005), .D(n_9627), .CD(n_61290), .Q(\wrD[5] 
		));
	notech_mux2 i_13066(.S(n_60396), .A(\wrD[5] ), .B(n_58203), .Z(n_9627)
		);
	notech_nand3 i_80088(.A(n_890), .B(n_61910), .C(n_10147), .Z(n_57676));
	notech_reg wrD_reg_6(.CP(n_62005), .D(n_9633), .CD(n_61290), .Q(\wrD[6] 
		));
	notech_mux2 i_13074(.S(n_60396), .A(\wrD[6] ), .B(data_miss[6]), .Z(n_9633
		));
	notech_nand3 i_80090(.A(n_890), .B(n_61910), .C(n_10146), .Z(n_57682));
	notech_reg wrD_reg_7(.CP(n_62005), .D(n_9639), .CD(n_61290), .Q(\wrD[7] 
		));
	notech_mux2 i_13082(.S(n_60396), .A(\wrD[7] ), .B(data_miss[7]), .Z(n_9639
		));
	notech_nand3 i_80092(.A(n_890), .B(n_61910), .C(n_10145), .Z(n_57688));
	notech_reg req_miss_reg(.CP(n_62005), .D(n_9645), .CD(n_61290), .Q(req_miss
		));
	notech_mux2 i_13090(.S(n_10080), .A(req_miss), .B(n_58109), .Z(n_9645)
		);
	notech_nand3 i_80094(.A(n_890), .B(n_61915), .C(n_10144), .Z(n_57694));
	notech_reg cr2_reg_0(.CP(n_62005), .D(n_9651), .CD(n_61290), .Q(cr2[0])
		);
	notech_mux2 i_13098(.S(n_808), .A(iDaddr_f[0]), .B(cr2[0]), .Z(n_9651)
		);
	notech_nand3 i_80096(.A(n_890), .B(n_61915), .C(n_10143), .Z(n_57700));
	notech_reg cr2_reg_1(.CP(n_62005), .D(n_9657), .CD(n_61290), .Q(cr2[1])
		);
	notech_mux2 i_13106(.S(n_808), .A(iDaddr_f[1]), .B(cr2[1]), .Z(n_9657)
		);
	notech_nao3 i_80098(.A(n_890), .B(n_61915), .C(data_miss[12]), .Z(n_57706
		));
	notech_reg cr2_reg_2(.CP(n_62006), .D(n_9663), .CD(n_61291), .Q(cr2[2])
		);
	notech_mux2 i_13114(.S(n_808), .A(iDaddr_f[2]), .B(cr2[2]), .Z(n_9663)
		);
	notech_nao3 i_80100(.A(n_890), .B(n_61915), .C(data_miss[13]), .Z(n_57712
		));
	notech_reg cr2_reg_3(.CP(n_62011), .D(n_9669), .CD(n_61296), .Q(cr2[3])
		);
	notech_mux2 i_13122(.S(n_808), .A(iDaddr_f[3]), .B(cr2[3]), .Z(n_9669)
		);
	notech_nao3 i_80102(.A(n_890), .B(n_61915), .C(data_miss[14]), .Z(n_57718
		));
	notech_reg cr2_reg_4(.CP(n_62015), .D(n_9675), .CD(n_61300), .Q(cr2[4])
		);
	notech_mux2 i_13130(.S(n_808), .A(iDaddr_f[4]), .B(cr2[4]), .Z(n_9675)
		);
	notech_nao3 i_80104(.A(n_890), .B(n_61915), .C(data_miss[15]), .Z(n_57724
		));
	notech_reg cr2_reg_5(.CP(n_62015), .D(n_9681), .CD(n_61300), .Q(cr2[5])
		);
	notech_mux2 i_13138(.S(n_808), .A(iDaddr_f[5]), .B(cr2[5]), .Z(n_9681)
		);
	notech_nao3 i_80106(.A(n_61184), .B(n_61915), .C(data_miss[16]), .Z(n_57730
		));
	notech_reg cr2_reg_6(.CP(n_62011), .D(n_9687), .CD(n_61296), .Q(cr2[6])
		);
	notech_mux2 i_13146(.S(n_808), .A(iDaddr_f[6]), .B(cr2[6]), .Z(n_9687)
		);
	notech_nao3 i_80108(.A(n_61184), .B(n_61917), .C(data_miss[17]), .Z(n_57736
		));
	notech_reg cr2_reg_7(.CP(n_62011), .D(n_9693), .CD(n_61296), .Q(cr2[7])
		);
	notech_mux2 i_13154(.S(n_808), .A(iDaddr_f[7]), .B(cr2[7]), .Z(n_9693)
		);
	notech_nao3 i_80110(.A(n_61184), .B(n_61915), .C(data_miss[18]), .Z(n_57742
		));
	notech_reg cr2_reg_8(.CP(n_62011), .D(n_9699), .CD(n_61296), .Q(cr2[8])
		);
	notech_mux2 i_13162(.S(n_808), .A(iDaddr_f[8]), .B(cr2[8]), .Z(n_9699)
		);
	notech_nao3 i_80112(.A(n_61184), .B(n_61915), .C(data_miss[19]), .Z(n_57748
		));
	notech_reg cr2_reg_9(.CP(n_62011), .D(n_9705), .CD(n_61296), .Q(cr2[9])
		);
	notech_mux2 i_13170(.S(n_808), .A(iDaddr_f[9]), .B(cr2[9]), .Z(n_9705)
		);
	notech_nao3 i_80114(.A(n_61184), .B(n_61915), .C(data_miss[20]), .Z(n_57754
		));
	notech_reg cr2_reg_10(.CP(n_62015), .D(n_9711), .CD(n_61300), .Q(cr2[10]
		));
	notech_mux2 i_13178(.S(n_808), .A(iDaddr_f[10]), .B(cr2[10]), .Z(n_9711)
		);
	notech_nao3 i_80116(.A(n_61184), .B(n_61915), .C(data_miss[21]), .Z(n_57760
		));
	notech_reg cr2_reg_11(.CP(n_62015), .D(n_9717), .CD(n_61300), .Q(cr2[11]
		));
	notech_mux2 i_13186(.S(n_808), .A(iDaddr_f[11]), .B(cr2[11]), .Z(n_9717)
		);
	notech_nao3 i_80118(.A(n_61184), .B(n_61912), .C(data_miss[22]), .Z(n_57766
		));
	notech_reg cr2_reg_12(.CP(n_62015), .D(n_9723), .CD(n_61300), .Q(cr2[12]
		));
	notech_mux2 i_13194(.S(n_808), .A(iDaddr_f[12]), .B(cr2[12]), .Z(n_9723)
		);
	notech_nao3 i_80120(.A(n_61184), .B(n_61912), .C(data_miss[23]), .Z(n_57772
		));
	notech_reg cr2_reg_13(.CP(n_62015), .D(n_9729), .CD(n_61300), .Q(cr2[13]
		));
	notech_mux2 i_13202(.S(n_808), .A(iDaddr_f[13]), .B(cr2[13]), .Z(n_9729)
		);
	notech_nao3 i_80122(.A(n_61184), .B(n_61912), .C(data_miss[24]), .Z(n_57778
		));
	notech_reg cr2_reg_14(.CP(n_62015), .D(n_9735), .CD(n_61300), .Q(cr2[14]
		));
	notech_mux2 i_13210(.S(n_808), .A(iDaddr_f[14]), .B(cr2[14]), .Z(n_9735)
		);
	notech_nao3 i_80124(.A(n_61184), .B(n_61912), .C(data_miss[25]), .Z(n_57784
		));
	notech_reg cr2_reg_15(.CP(n_62015), .D(n_9741), .CD(n_61300), .Q(cr2[15]
		));
	notech_mux2 i_13218(.S(n_808), .A(iDaddr_f[15]), .B(cr2[15]), .Z(n_9741)
		);
	notech_nao3 i_80126(.A(n_61184), .B(n_61912), .C(data_miss[26]), .Z(n_57790
		));
	notech_reg cr2_reg_16(.CP(n_62015), .D(n_9747), .CD(n_61300), .Q(cr2[16]
		));
	notech_mux2 i_13226(.S(n_54440), .A(iDaddr_f[16]), .B(cr2[16]), .Z(n_9747
		));
	notech_nao3 i_80128(.A(n_890), .B(n_61912), .C(data_miss[27]), .Z(n_57796
		));
	notech_reg cr2_reg_17(.CP(n_62011), .D(n_9753), .CD(n_61296), .Q(cr2[17]
		));
	notech_mux2 i_13234(.S(n_54440), .A(iDaddr_f[17]), .B(cr2[17]), .Z(n_9753
		));
	notech_nao3 i_80130(.A(n_61184), .B(n_61915), .C(data_miss[28]), .Z(n_57802
		));
	notech_reg cr2_reg_18(.CP(n_62011), .D(n_9759), .CD(n_61296), .Q(cr2[18]
		));
	notech_mux2 i_13242(.S(n_54440), .A(iDaddr_f[18]), .B(cr2[18]), .Z(n_9759
		));
	notech_nao3 i_80132(.A(n_61184), .B(n_61915), .C(data_miss[29]), .Z(n_57808
		));
	notech_reg cr2_reg_19(.CP(n_62011), .D(n_9765), .CD(n_61296), .Q(cr2[19]
		));
	notech_mux2 i_13250(.S(n_54440), .A(iDaddr_f[19]), .B(cr2[19]), .Z(n_9765
		));
	notech_nao3 i_80134(.A(n_61184), .B(n_61915), .C(data_miss[30]), .Z(n_57814
		));
	notech_reg cr2_reg_20(.CP(n_62011), .D(n_9771), .CD(n_61296), .Q(cr2[20]
		));
	notech_mux2 i_13258(.S(n_54440), .A(iDaddr_f[20]), .B(cr2[20]), .Z(n_9771
		));
	notech_nao3 i_80136(.A(n_61184), .B(n_61915), .C(data_miss[31]), .Z(n_57820
		));
	notech_reg cr2_reg_21(.CP(n_62011), .D(n_9777), .CD(n_61296), .Q(cr2[21]
		));
	notech_mux2 i_13266(.S(n_54440), .A(iDaddr_f[21]), .B(cr2[21]), .Z(n_9777
		));
	notech_nand2 i_80142(.A(n_61184), .B(n_61915), .Z(n_57844));
	notech_reg cr2_reg_22(.CP(n_62006), .D(n_9783), .CD(n_61291), .Q(cr2[22]
		));
	notech_mux2 i_13274(.S(n_54440), .A(iDaddr_f[22]), .B(cr2[22]), .Z(n_9783
		));
	notech_ao4 i_80150(.A(n_916), .B(n_10010), .C(n_896), .D(\nnx_tab2[0] ),
		 .Z(n_60188));
	notech_reg cr2_reg_23(.CP(n_62006), .D(n_9789), .CD(n_61291), .Q(cr2[23]
		));
	notech_mux2 i_13282(.S(n_54440), .A(iDaddr_f[23]), .B(cr2[23]), .Z(n_9789
		));
	notech_ao4 i_80153(.A(n_916), .B(n_10012), .C(n_896), .D(n_478), .Z(n_60194
		));
	notech_reg cr2_reg_24(.CP(n_62011), .D(n_9795), .CD(n_61296), .Q(cr2[24]
		));
	notech_mux2 i_13290(.S(n_54440), .A(iDaddr_f[24]), .B(cr2[24]), .Z(n_9795
		));
	notech_ao4 i_80160(.A(n_896), .B(n_10005), .C(n_466), .D(n_926), .Z(n_60215
		));
	notech_reg cr2_reg_25(.CP(n_62011), .D(n_9801), .CD(n_61296), .Q(cr2[25]
		));
	notech_mux2 i_13298(.S(n_54440), .A(iDaddr_f[25]), .B(cr2[25]), .Z(n_9801
		));
	notech_ao4 i_80163(.A(n_896), .B(n_10007), .C(n_471), .D(n_927), .Z(n_60221
		));
	notech_reg cr2_reg_26(.CP(n_62011), .D(n_9807), .CD(n_61296), .Q(cr2[26]
		));
	notech_mux2 i_13306(.S(n_54440), .A(iDaddr_f[26]), .B(cr2[26]), .Z(n_9807
		));
	notech_ao4 i_80170(.A(n_896), .B(n_9959), .C(n_495), .D(n_917), .Z(n_58149
		));
	notech_reg cr2_reg_27(.CP(n_62011), .D(n_9813), .CD(n_61296), .Q(cr2[27]
		));
	notech_mux2 i_13314(.S(n_54440), .A(iDaddr_f[27]), .B(cr2[27]), .Z(n_9813
		));
	notech_ao4 i_80173(.A(n_896), .B(n_9961), .C(n_500), .D(n_918), .Z(n_58155
		));
	notech_reg cr2_reg_28(.CP(n_62011), .D(n_9819), .CD(n_61296), .Q(cr2[28]
		));
	notech_mux2 i_13322(.S(n_54440), .A(iDaddr_f[28]), .B(cr2[28]), .Z(n_9819
		));
	notech_nand3 i_43(.A(n_916), .B(n_935), .C(n_858), .Z(n_58091));
	notech_reg cr2_reg_29(.CP(n_62011), .D(n_9825), .CD(n_61296), .Q(cr2[29]
		));
	notech_mux2 i_13330(.S(n_54440), .A(iDaddr_f[29]), .B(cr2[29]), .Z(n_9825
		));
	notech_nand3 i_42(.A(n_938), .B(n_855), .C(n_937), .Z(n_58085));
	notech_reg cr2_reg_30(.CP(n_62011), .D(n_9831), .CD(n_61296), .Q(cr2[30]
		));
	notech_mux2 i_13338(.S(n_54440), .A(iDaddr_f[30]), .B(cr2[30]), .Z(n_9831
		));
	notech_mux2 i_41(.S(n_61926), .A(n_447), .B(n_445), .Z(n_58079));
	notech_reg cr2_reg_31(.CP(n_62011), .D(n_9837), .CD(n_61296), .Q(cr2[31]
		));
	notech_mux2 i_13346(.S(n_54440), .A(iDaddr_f[31]), .B(cr2[31]), .Z(n_9837
		));
	notech_inv i_14828(.A(n_985), .Z(n_9843));
	notech_inv i_14829(.A(n_901), .Z(n_9844));
	notech_inv i_14830(.A(n_459), .Z(n_9845));
	notech_inv i_14831(.A(n_889), .Z(n_9846));
	notech_inv i_14832(.A(n_883), .Z(n_9847));
	notech_inv i_14833(.A(\dir1[10] ), .Z(n_9848));
	notech_inv i_14834(.A(\dir1[11] ), .Z(n_9849));
	notech_inv i_14835(.A(\dir1[12] ), .Z(n_9850));
	notech_inv i_14836(.A(\dir1[13] ), .Z(n_9851));
	notech_inv i_14837(.A(\dir1[14] ), .Z(n_9852));
	notech_inv i_14838(.A(\dir1[15] ), .Z(n_9853));
	notech_inv i_14839(.A(\dir1[16] ), .Z(n_9854));
	notech_inv i_14840(.A(\dir1[17] ), .Z(n_9855));
	notech_inv i_14841(.A(\dir1[18] ), .Z(n_9856));
	notech_inv i_14842(.A(\dir1[19] ), .Z(n_9857));
	notech_inv i_14843(.A(\dir1[20] ), .Z(n_9858));
	notech_inv i_14844(.A(\dir1[21] ), .Z(n_9859));
	notech_inv i_14845(.A(\dir1[22] ), .Z(n_9860));
	notech_inv i_14846(.A(\dir1[23] ), .Z(n_9861));
	notech_inv i_14847(.A(\dir1[24] ), .Z(n_9862));
	notech_inv i_14848(.A(\dir1[25] ), .Z(n_9863));
	notech_inv i_14849(.A(\dir1[26] ), .Z(n_9864));
	notech_inv i_14850(.A(\dir1[27] ), .Z(n_9865));
	notech_inv i_14851(.A(\dir1[28] ), .Z(n_9866));
	notech_inv i_14852(.A(\dir1[29] ), .Z(n_9867));
	notech_inv i_14853(.A(\dir2[10] ), .Z(n_9868));
	notech_inv i_14854(.A(\dir2[11] ), .Z(n_9869));
	notech_inv i_14855(.A(\dir2[12] ), .Z(n_9870));
	notech_inv i_14856(.A(\dir2[13] ), .Z(n_9871));
	notech_inv i_14857(.A(\dir2[14] ), .Z(n_9872));
	notech_inv i_14858(.A(\dir2[15] ), .Z(n_9873));
	notech_inv i_14859(.A(\dir2[16] ), .Z(n_9874));
	notech_inv i_14860(.A(\dir2[17] ), .Z(n_9875));
	notech_inv i_14861(.A(\dir2[18] ), .Z(n_9876));
	notech_inv i_14862(.A(\dir2[19] ), .Z(n_9877));
	notech_inv i_14863(.A(\dir2[20] ), .Z(n_9878));
	notech_inv i_14864(.A(\dir2[21] ), .Z(n_9879));
	notech_inv i_14865(.A(\dir2[22] ), .Z(n_9880));
	notech_inv i_14866(.A(\dir2[23] ), .Z(n_9881));
	notech_inv i_14867(.A(\dir2[24] ), .Z(n_9882));
	notech_inv i_14868(.A(\dir2[25] ), .Z(n_9883));
	notech_inv i_14869(.A(\dir2[26] ), .Z(n_9884));
	notech_inv i_14870(.A(\dir2[27] ), .Z(n_9885));
	notech_inv i_14871(.A(\dir2[28] ), .Z(n_9886));
	notech_inv i_14872(.A(\dir2[29] ), .Z(n_9887));
	notech_inv i_14873(.A(n_476), .Z(n_9888));
	notech_inv i_14874(.A(\tab21[10] ), .Z(n_9889));
	notech_inv i_14875(.A(\tab21[11] ), .Z(n_9890));
	notech_inv i_14876(.A(\tab21[12] ), .Z(n_9891));
	notech_inv i_14877(.A(\tab21[13] ), .Z(n_9892));
	notech_inv i_14878(.A(\tab21[14] ), .Z(n_9893));
	notech_inv i_14879(.A(n_488), .Z(n_9894));
	notech_inv i_14880(.A(\tab21[15] ), .Z(n_9895));
	notech_inv i_14881(.A(\tab21[16] ), .Z(n_9896));
	notech_inv i_14882(.A(\tab21[17] ), .Z(n_9897));
	notech_inv i_14883(.A(\tab21[18] ), .Z(n_9898));
	notech_inv i_14884(.A(\tab21[19] ), .Z(n_9899));
	notech_inv i_14885(.A(\tab21[20] ), .Z(n_9900));
	notech_inv i_14886(.A(\tab21[21] ), .Z(n_9901));
	notech_inv i_14887(.A(\tab21[22] ), .Z(n_9902));
	notech_inv i_14888(.A(\tab21[23] ), .Z(n_9903));
	notech_inv i_14889(.A(\tab21[24] ), .Z(n_9904));
	notech_inv i_14890(.A(\tab21[25] ), .Z(n_9905));
	notech_inv i_14891(.A(\tab21[26] ), .Z(n_9906));
	notech_inv i_14892(.A(\tab21[27] ), .Z(n_9907));
	notech_inv i_14893(.A(\tab21[28] ), .Z(n_9908));
	notech_inv i_14894(.A(\tab21[29] ), .Z(n_9909));
	notech_inv i_14895(.A(\tab12[10] ), .Z(n_9910));
	notech_inv i_14896(.A(\tab12[11] ), .Z(n_9911));
	notech_inv i_14897(.A(\tab12[12] ), .Z(n_9912));
	notech_inv i_14898(.A(\tab12[13] ), .Z(n_9913));
	notech_inv i_14899(.A(\tab12[14] ), .Z(n_9914));
	notech_inv i_14900(.A(\tab12[15] ), .Z(n_9915));
	notech_inv i_14901(.A(\tab12[16] ), .Z(n_9916));
	notech_inv i_14902(.A(\tab12[17] ), .Z(n_9917));
	notech_inv i_14903(.A(\tab12[18] ), .Z(n_9918));
	notech_inv i_14904(.A(\tab12[19] ), .Z(n_9919));
	notech_inv i_14905(.A(\tab12[20] ), .Z(n_9920));
	notech_inv i_14906(.A(\tab12[21] ), .Z(n_9921));
	notech_inv i_14907(.A(\tab12[22] ), .Z(n_9922));
	notech_inv i_14908(.A(\tab12[23] ), .Z(n_9923));
	notech_inv i_14909(.A(\tab12[24] ), .Z(n_9924));
	notech_inv i_14910(.A(\tab12[25] ), .Z(n_9925));
	notech_inv i_14911(.A(\tab12[26] ), .Z(n_9926));
	notech_inv i_14912(.A(\tab12[27] ), .Z(n_9927));
	notech_inv i_14913(.A(\tab12[28] ), .Z(n_9928));
	notech_inv i_14914(.A(\tab12[29] ), .Z(n_9929));
	notech_inv i_14915(.A(n_553), .Z(n_9930));
	notech_inv i_14916(.A(n_557), .Z(n_9931));
	notech_inv i_14917(.A(n_559), .Z(n_9932));
	notech_inv i_14918(.A(hit_adr13), .Z(n_9933));
	notech_inv i_14919(.A(\tab14[10] ), .Z(n_9934));
	notech_inv i_14920(.A(\tab14[11] ), .Z(n_9935));
	notech_inv i_14921(.A(\tab14[12] ), .Z(n_9936));
	notech_inv i_14922(.A(\tab14[13] ), .Z(n_9937));
	notech_inv i_14923(.A(\tab14[14] ), .Z(n_9938));
	notech_inv i_14924(.A(\tab14[15] ), .Z(n_9939));
	notech_inv i_14925(.A(\tab14[16] ), .Z(n_9940));
	notech_inv i_14926(.A(\tab14[17] ), .Z(n_9941));
	notech_inv i_14927(.A(\tab14[18] ), .Z(n_9942));
	notech_inv i_14928(.A(\tab14[19] ), .Z(n_9943));
	notech_inv i_14929(.A(\tab14[20] ), .Z(n_9944));
	notech_inv i_14930(.A(\tab14[21] ), .Z(n_9945));
	notech_inv i_14931(.A(\tab14[22] ), .Z(n_9946));
	notech_inv i_14932(.A(\tab14[23] ), .Z(n_9947));
	notech_inv i_14933(.A(\tab14[24] ), .Z(n_9948));
	notech_inv i_14934(.A(\tab14[25] ), .Z(n_9949));
	notech_inv i_14935(.A(\tab14[26] ), .Z(n_9950));
	notech_inv i_14936(.A(\tab14[27] ), .Z(n_9951));
	notech_inv i_14937(.A(\tab14[28] ), .Z(n_9952));
	notech_inv i_14938(.A(\tab14[29] ), .Z(n_9953));
	notech_inv i_14939(.A(n_58149), .Z(n_9954));
	notech_inv i_14940(.A(\nx_tab1[0] ), .Z(n_9955));
	notech_inv i_14941(.A(n_58155), .Z(n_9956));
	notech_inv i_14942(.A(\nx_tab1[1] ), .Z(n_9957));
	notech_inv i_14943(.A(n_57173), .Z(n_9958));
	notech_inv i_14944(.A(\nnx_tab1[0] ), .Z(n_9959));
	notech_inv i_14945(.A(n_57179), .Z(n_9960));
	notech_inv i_14946(.A(\nnx_tab1[1] ), .Z(n_9961));
	notech_inv i_14947(.A(\nbus_14489[0] ), .Z(n_9962));
	notech_inv i_14948(.A(\tab23[10] ), .Z(n_9963));
	notech_inv i_14949(.A(\tab23[11] ), .Z(n_9964));
	notech_inv i_14950(.A(\tab23[12] ), .Z(n_9965));
	notech_inv i_14951(.A(\tab23[13] ), .Z(n_9966));
	notech_inv i_14952(.A(\tab23[14] ), .Z(n_9967));
	notech_inv i_14953(.A(\tab23[15] ), .Z(n_9968));
	notech_inv i_14954(.A(\tab23[16] ), .Z(n_9969));
	notech_inv i_14955(.A(\tab23[17] ), .Z(n_9970));
	notech_inv i_14956(.A(\tab23[18] ), .Z(n_9971));
	notech_inv i_14957(.A(\tab23[19] ), .Z(n_9972));
	notech_inv i_14958(.A(\tab23[20] ), .Z(n_9973));
	notech_inv i_14959(.A(\tab23[21] ), .Z(n_9974));
	notech_inv i_14960(.A(\tab23[22] ), .Z(n_9975));
	notech_inv i_14961(.A(\tab23[23] ), .Z(n_9976));
	notech_inv i_14962(.A(\tab23[24] ), .Z(n_9977));
	notech_inv i_14963(.A(\tab23[25] ), .Z(n_9978));
	notech_inv i_14964(.A(\tab23[26] ), .Z(n_9979));
	notech_inv i_14965(.A(\tab23[27] ), .Z(n_9980));
	notech_inv i_14966(.A(\tab23[28] ), .Z(n_9981));
	notech_inv i_14967(.A(\tab23[29] ), .Z(n_9982));
	notech_inv i_14968(.A(hit_adr23), .Z(n_9983));
	notech_inv i_14969(.A(\tab24[10] ), .Z(n_9984));
	notech_inv i_14970(.A(\tab24[11] ), .Z(n_9985));
	notech_inv i_14971(.A(\tab24[12] ), .Z(n_9986));
	notech_inv i_14972(.A(\tab24[13] ), .Z(n_9987));
	notech_inv i_14973(.A(\tab24[14] ), .Z(n_9988));
	notech_inv i_14974(.A(\tab24[15] ), .Z(n_9989));
	notech_inv i_14975(.A(\tab24[16] ), .Z(n_9990));
	notech_inv i_14976(.A(\tab24[17] ), .Z(n_9991));
	notech_inv i_14977(.A(\tab24[18] ), .Z(n_9992));
	notech_inv i_14978(.A(\tab24[19] ), .Z(n_9993));
	notech_inv i_14979(.A(\tab24[20] ), .Z(n_9994));
	notech_inv i_14980(.A(\tab24[21] ), .Z(n_9995));
	notech_inv i_14981(.A(\tab24[22] ), .Z(n_9996));
	notech_inv i_14982(.A(\tab24[23] ), .Z(n_9997));
	notech_inv i_14983(.A(\tab24[24] ), .Z(n_9998));
	notech_inv i_14984(.A(\tab24[25] ), .Z(n_9999));
	notech_inv i_14985(.A(\tab24[26] ), .Z(n_10000));
	notech_inv i_14986(.A(\tab24[27] ), .Z(n_10001));
	notech_inv i_14987(.A(\tab24[28] ), .Z(n_10002));
	notech_inv i_14988(.A(\tab24[29] ), .Z(n_10003));
	notech_inv i_14989(.A(n_60188), .Z(n_10004));
	notech_inv i_14990(.A(\nnx_tab2[0] ), .Z(n_10005));
	notech_inv i_14991(.A(n_60194), .Z(n_10006));
	notech_inv i_14992(.A(\nnx_tab2[1] ), .Z(n_10007));
	notech_inv i_14993(.A(\nbus_14515[0] ), .Z(n_10008));
	notech_inv i_14994(.A(n_60215), .Z(n_10009));
	notech_inv i_14995(.A(\nx_tab2[0] ), .Z(n_10010));
	notech_inv i_14996(.A(n_60221), .Z(n_10011));
	notech_inv i_14997(.A(\nx_tab2[1] ), .Z(n_10012));
	notech_inv i_14998(.A(\tab11[10] ), .Z(n_10013));
	notech_inv i_14999(.A(\tab11[11] ), .Z(n_10014));
	notech_inv i_15000(.A(\tab11[12] ), .Z(n_10015));
	notech_inv i_15001(.A(\tab11[13] ), .Z(n_10016));
	notech_inv i_15002(.A(\tab11[14] ), .Z(n_10017));
	notech_inv i_15003(.A(\tab11[15] ), .Z(n_10018));
	notech_inv i_15004(.A(\tab11[16] ), .Z(n_10019));
	notech_inv i_15005(.A(\tab11[17] ), .Z(n_10020));
	notech_inv i_15006(.A(\tab11[18] ), .Z(n_10021));
	notech_inv i_15007(.A(\tab11[19] ), .Z(n_10022));
	notech_inv i_15008(.A(\tab11[20] ), .Z(n_10023));
	notech_inv i_15009(.A(\tab11[21] ), .Z(n_10024));
	notech_inv i_15010(.A(\tab11[22] ), .Z(n_10025));
	notech_inv i_15011(.A(\tab11[23] ), .Z(n_10026));
	notech_inv i_15012(.A(\tab11[24] ), .Z(n_10027));
	notech_inv i_15013(.A(\tab11[25] ), .Z(n_10028));
	notech_inv i_15014(.A(\tab11[26] ), .Z(n_10029));
	notech_inv i_15015(.A(\tab11[27] ), .Z(n_10030));
	notech_inv i_15016(.A(\tab11[28] ), .Z(n_10031));
	notech_inv i_15017(.A(\tab11[29] ), .Z(n_10032));
	notech_inv i_15018(.A(n_59947), .Z(n_10033));
	notech_inv i_15019(.A(n_61926), .Z(n_10034));
	notech_inv i_15020(.A(fsm[3]), .Z(n_10035));
	notech_inv i_15021(.A(n_59530), .Z(n_10036));
	notech_inv i_15022(.A(n_59536), .Z(n_10037));
	notech_inv i_15023(.A(n_59542), .Z(n_10038));
	notech_inv i_15024(.A(n_59548), .Z(n_10039));
	notech_inv i_15025(.A(n_59554), .Z(n_10040));
	notech_inv i_15026(.A(n_59560), .Z(n_10041));
	notech_inv i_15027(.A(n_59566), .Z(n_10042));
	notech_inv i_15028(.A(n_59572), .Z(n_10043));
	notech_inv i_15029(.A(n_59578), .Z(n_10044));
	notech_inv i_15030(.A(n_59584), .Z(n_10045));
	notech_inv i_15031(.A(\addr_miss[2] ), .Z(n_10046));
	notech_inv i_15032(.A(\addr_miss[3] ), .Z(n_10047));
	notech_inv i_15033(.A(\addr_miss[4] ), .Z(n_10048));
	notech_inv i_15034(.A(\addr_miss[5] ), .Z(n_10049));
	notech_inv i_15035(.A(\addr_miss[6] ), .Z(n_10050));
	notech_inv i_15036(.A(\addr_miss[7] ), .Z(n_10051));
	notech_inv i_15037(.A(\addr_miss[8] ), .Z(n_10052));
	notech_inv i_15038(.A(\addr_miss[9] ), .Z(n_10053));
	notech_inv i_15039(.A(\addr_miss[10] ), .Z(n_10054));
	notech_inv i_15040(.A(\addr_miss[11] ), .Z(n_10055));
	notech_inv i_15041(.A(\wrA[12] ), .Z(n_10056));
	notech_inv i_15042(.A(\wrA[13] ), .Z(n_10057));
	notech_inv i_15043(.A(\wrA[14] ), .Z(n_10058));
	notech_inv i_15044(.A(\wrA[15] ), .Z(n_10059));
	notech_inv i_15045(.A(\wrA[16] ), .Z(n_10060));
	notech_inv i_15046(.A(\wrA[17] ), .Z(n_10061));
	notech_inv i_15047(.A(\wrA[18] ), .Z(n_10062));
	notech_inv i_15048(.A(\wrA[19] ), .Z(n_10063));
	notech_inv i_15049(.A(\wrA[20] ), .Z(n_10064));
	notech_inv i_15050(.A(\wrA[21] ), .Z(n_10065));
	notech_inv i_15051(.A(\wrA[22] ), .Z(n_10066));
	notech_inv i_15052(.A(\wrA[23] ), .Z(n_10067));
	notech_inv i_15053(.A(\wrA[24] ), .Z(n_10068));
	notech_inv i_15054(.A(\wrA[25] ), .Z(n_10069));
	notech_inv i_15055(.A(\wrA[26] ), .Z(n_10070));
	notech_inv i_15056(.A(\wrA[27] ), .Z(n_10071));
	notech_inv i_15057(.A(\wrA[28] ), .Z(n_10072));
	notech_inv i_15058(.A(\wrA[29] ), .Z(n_10073));
	notech_inv i_15059(.A(\wrA[30] ), .Z(n_10074));
	notech_inv i_15060(.A(\wrA[31] ), .Z(n_10075));
	notech_inv i_15061(.A(n_58203), .Z(n_10076));
	notech_inv i_15063(.A(n_58109), .Z(n_10078));
	notech_inv i_15064(.A(req_miss), .Z(n_10079));
	notech_inv i_15065(.A(n_58106), .Z(n_10080));
	notech_inv i_15066(.A(addr_phys_31100160), .Z(addr_phys[31]));
	notech_inv i_15067(.A(addr_phys_30100159), .Z(addr_phys[30]));
	notech_inv i_15068(.A(addr_phys_29100158), .Z(addr_phys[29]));
	notech_inv i_15069(.A(addr_phys_28100157), .Z(addr_phys[28]));
	notech_inv i_15070(.A(addr_phys_27100156), .Z(addr_phys[27]));
	notech_inv i_15071(.A(addr_phys_26100155), .Z(addr_phys[26]));
	notech_inv i_15072(.A(addr_phys_25100154), .Z(addr_phys[25]));
	notech_inv i_15073(.A(addr_phys_24100153), .Z(addr_phys[24]));
	notech_inv i_15074(.A(addr_phys_23100152), .Z(addr_phys[23]));
	notech_inv i_15075(.A(addr_phys_22100151), .Z(addr_phys[22]));
	notech_inv i_15076(.A(addr_phys_21100150), .Z(addr_phys[21]));
	notech_inv i_15077(.A(addr_phys_20100149), .Z(addr_phys[20]));
	notech_inv i_15078(.A(addr_phys_19100148), .Z(addr_phys[19]));
	notech_inv i_15079(.A(addr_phys_18100147), .Z(addr_phys[18]));
	notech_inv i_15080(.A(addr_phys_17100146), .Z(addr_phys[17]));
	notech_inv i_15081(.A(addr_phys_16100145), .Z(addr_phys[16]));
	notech_inv i_15082(.A(addr_phys_15100144), .Z(addr_phys[15]));
	notech_inv i_15083(.A(addr_phys_14100143), .Z(addr_phys[14]));
	notech_inv i_15084(.A(addr_phys_13100142), .Z(addr_phys[13]));
	notech_inv i_15085(.A(addr_phys_12100141), .Z(addr_phys[12]));
	notech_inv i_15086(.A(n_60810), .Z(n_10101));
	notech_inv i_15087(.A(iDaddr[2]), .Z(n_10102));
	notech_inv i_15088(.A(iDaddr[3]), .Z(n_10103));
	notech_inv i_15089(.A(iDaddr[4]), .Z(n_10104));
	notech_inv i_15090(.A(iDaddr[5]), .Z(n_10105));
	notech_inv i_15091(.A(iDaddr[6]), .Z(n_10106));
	notech_inv i_15092(.A(iDaddr[7]), .Z(n_10107));
	notech_inv i_15093(.A(iDaddr[8]), .Z(n_10108));
	notech_inv i_15094(.A(iDaddr[9]), .Z(n_10109));
	notech_inv i_15095(.A(iDaddr[10]), .Z(n_10110));
	notech_inv i_15096(.A(iDaddr[11]), .Z(n_10111));
	notech_inv i_15097(.A(iDaddr[12]), .Z(n_10112));
	notech_inv i_15098(.A(iDaddr[13]), .Z(n_10113));
	notech_inv i_15099(.A(iDaddr[14]), .Z(n_10114));
	notech_inv i_15100(.A(iDaddr[15]), .Z(n_10115));
	notech_inv i_15101(.A(iDaddr[16]), .Z(n_10116));
	notech_inv i_15102(.A(iDaddr[17]), .Z(n_10117));
	notech_inv i_15103(.A(iDaddr[18]), .Z(n_10118));
	notech_inv i_15104(.A(iDaddr[19]), .Z(n_10119));
	notech_inv i_15105(.A(iDaddr[20]), .Z(n_10120));
	notech_inv i_15106(.A(iDaddr[21]), .Z(n_10121));
	notech_inv i_15107(.A(iDaddr[22]), .Z(n_10122));
	notech_inv i_15108(.A(iDaddr[23]), .Z(n_10123));
	notech_inv i_15109(.A(iDaddr[24]), .Z(n_10124));
	notech_inv i_15110(.A(iDaddr[25]), .Z(n_10125));
	notech_inv i_15111(.A(iDaddr[26]), .Z(n_10126));
	notech_inv i_15112(.A(iDaddr[27]), .Z(n_10127));
	notech_inv i_15113(.A(iDaddr[28]), .Z(n_10128));
	notech_inv i_15114(.A(iDaddr[29]), .Z(n_10129));
	notech_inv i_15115(.A(iDaddr[30]), .Z(n_10130));
	notech_inv i_15116(.A(iDaddr[31]), .Z(n_10131));
	notech_inv i_15117(.A(n_61901), .Z(owrite_req));
	notech_inv i_15118(.A(\dir1_0[9] ), .Z(n_10133));
	notech_inv i_15119(.A(\dir1_0[8] ), .Z(n_10134));
	notech_inv i_15120(.A(\dir1_0[7] ), .Z(n_10135));
	notech_inv i_15121(.A(\dir1_0[6] ), .Z(n_10136));
	notech_inv i_15122(.A(\dir1_0[5] ), .Z(n_10137));
	notech_inv i_15123(.A(\dir1_0[4] ), .Z(n_10138));
	notech_inv i_15124(.A(\dir1_0[3] ), .Z(n_10139));
	notech_inv i_15125(.A(\dir1_0[2] ), .Z(n_10140));
	notech_inv i_15126(.A(\dir1_0[1] ), .Z(n_10141));
	notech_inv i_15127(.A(\dir1_0[0] ), .Z(n_10142));
	notech_inv i_15128(.A(\tab11_0[9] ), .Z(n_10143));
	notech_inv i_15129(.A(\tab11_0[8] ), .Z(n_10144));
	notech_inv i_15130(.A(\tab11_0[7] ), .Z(n_10145));
	notech_inv i_15131(.A(\tab11_0[6] ), .Z(n_10146));
	notech_inv i_15132(.A(\tab11_0[5] ), .Z(n_10147));
	notech_inv i_15133(.A(\tab11_0[4] ), .Z(n_10148));
	notech_inv i_15134(.A(\tab11_0[3] ), .Z(n_10149));
	notech_inv i_15135(.A(\tab11_0[2] ), .Z(n_10150));
	notech_inv i_15136(.A(\tab11_0[1] ), .Z(n_10151));
	notech_inv i_15137(.A(\tab11_0[0] ), .Z(n_10152));
	notech_inv i_15138(.A(oread_req100140), .Z(oread_req));
	notech_inv i_15139(.A(hit_tab21), .Z(n_10154));
	notech_inv i_15140(.A(hit_tab23), .Z(n_10155));
	notech_inv i_15141(.A(hit_tab12), .Z(n_10156));
	notech_inv i_15142(.A(\hit_dir1[7] ), .Z(n_10157));
	notech_inv i_15143(.A(n_61941), .Z(n_10158));
	notech_inv i_15144(.A(iread_req), .Z(n_10159));
	notech_inv i_15145(.A(hit_dir2), .Z(n_10160));
	notech_inv i_15146(.A(pg_fault), .Z(n_10161));
	cmp14_19 t11(.ina({\tab11[33] , UNCONNECTED_000, UNCONNECTED_001, 
		UNCONNECTED_002, \tab11[9] , \tab11[8] , \tab11[7] , \tab11[6] ,
		 \tab11[5] , \tab11[4] , \tab11[3] , \tab11[2] , \tab11[1] , \tab11[0] 
		}), .inb({UNCONNECTED_003, UNCONNECTED_004, UNCONNECTED_005, 
		UNCONNECTED_006, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab11), .out2(hit_add11));
	cmp14_18 t24(.ina({\tab24[33] , UNCONNECTED_007, UNCONNECTED_008, 
		UNCONNECTED_009, \tab24[9] , \tab24[8] , \tab24[7] , \tab24[6] ,
		 \tab24[5] , \tab24[4] , \tab24[3] , \tab24[2] , \tab24[1] , \tab24[0] 
		}), .inb({UNCONNECTED_010, UNCONNECTED_011, UNCONNECTED_012, 
		UNCONNECTED_013, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab24), .out2(hit_add24));
	cmp14_17 t23(.ina({\tab23[33] , UNCONNECTED_014, UNCONNECTED_015, 
		UNCONNECTED_016, \tab23[9] , \tab23[8] , \tab23[7] , \tab23[6] ,
		 \tab23[5] , \tab23[4] , \tab23[3] , \tab23[2] , \tab23[1] , \tab23[0] 
		}), .inb({UNCONNECTED_017, UNCONNECTED_018, UNCONNECTED_019, 
		UNCONNECTED_020, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab23), .out2(hit_add23));
	cmp14_16 t22(.ina({\tab22[33] , UNCONNECTED_021, UNCONNECTED_022, 
		UNCONNECTED_023, \tab22[9] , \tab22[8] , \tab22[7] , \tab22[6] ,
		 \tab22[5] , \tab22[4] , \tab22[3] , \tab22[2] , \tab22[1] , \tab22[0] 
		}), .inb({UNCONNECTED_024, UNCONNECTED_025, UNCONNECTED_026, 
		UNCONNECTED_027, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab22), .out2(hit_add22));
	cmp14_15 t21(.ina({\tab21[33] , UNCONNECTED_028, UNCONNECTED_029, 
		UNCONNECTED_030, \tab21[9] , \tab21[8] , \tab21[7] , \tab21[6] ,
		 \tab21[5] , \tab21[4] , \tab21[3] , \tab21[2] , \tab21[1] , \tab21[0] 
		}), .inb({UNCONNECTED_031, UNCONNECTED_032, UNCONNECTED_033, 
		UNCONNECTED_034, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab21), .out2(hit_add21));
	cmp14_14 t14(.ina({\tab14[33] , UNCONNECTED_035, UNCONNECTED_036, 
		UNCONNECTED_037, \tab14[9] , \tab14[8] , \tab14[7] , \tab14[6] ,
		 \tab14[5] , \tab14[4] , \tab14[3] , \tab14[2] , \tab14[1] , \tab14[0] 
		}), .inb({UNCONNECTED_038, UNCONNECTED_039, UNCONNECTED_040, 
		UNCONNECTED_041, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab14), .out2(hit_add14));
	cmp14_13 t13(.ina({\tab13[33] , UNCONNECTED_042, UNCONNECTED_043, 
		UNCONNECTED_044, \tab13[9] , \tab13[8] , \tab13[7] , \tab13[6] ,
		 \tab13[5] , \tab13[4] , \tab13[3] , \tab13[2] , \tab13[1] , \tab13[0] 
		}), .inb({UNCONNECTED_045, UNCONNECTED_046, UNCONNECTED_047, 
		UNCONNECTED_048, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab13), .out2(hit_add13));
	cmp14_12 t12(.ina({\tab12[33] , UNCONNECTED_049, UNCONNECTED_050, 
		UNCONNECTED_051, \tab12[9] , \tab12[8] , \tab12[7] , \tab12[6] ,
		 \tab12[5] , \tab12[4] , \tab12[3] , \tab12[2] , \tab12[1] , \tab12[0] 
		}), .inb({UNCONNECTED_052, UNCONNECTED_053, UNCONNECTED_054, 
		UNCONNECTED_055, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab12), .out2(hit_add12));
	cmp14_11 d2(.ina({\dir2[33] , UNCONNECTED_056, UNCONNECTED_057, 
		UNCONNECTED_058, \dir2[9] , \dir2[8] , \dir2[7] , \dir2[6] , \dir2[5] 
		, \dir2[4] , \dir2[3] , \dir2[2] , \dir2[1] , \dir2[0] }), .inb(
		{UNCONNECTED_059, UNCONNECTED_060, UNCONNECTED_061, 
		UNCONNECTED_062, \dir1_0[9] , \dir1_0[8] , \dir1_0[7] , \dir1_0[6] 
		, \dir1_0[5] , \dir1_0[4] , \dir1_0[3] , \dir1_0[2] , \dir1_0[1] 
		, \dir1_0[0] }), .out(hit_dir2));
	cmp14_10 d1(.ina({\dir1[33] , UNCONNECTED_063, UNCONNECTED_064, 
		UNCONNECTED_065, \dir1[9] , \dir1[8] , \dir1[7] , \dir1[6] , \dir1[5] 
		, \dir1[4] , \dir1[3] , \dir1[2] , \dir1[1] , \dir1[0] }), .inb(
		{UNCONNECTED_066, UNCONNECTED_067, UNCONNECTED_068, 
		UNCONNECTED_069, \dir1_0[9] , \dir1_0[8] , \dir1_0[7] , \dir1_0[6] 
		, \dir1_0[5] , \dir1_0[4] , \dir1_0[3] , \dir1_0[2] , \dir1_0[1] 
		, \dir1_0[0] }), .out(\hit_dir1[7] ));
	AWDP_INC_26 i_79019(.O0(fsm5_cnt_0), .fsm5_cnt(fsm5_cnt));
endmodule
module AWDP_partition_33(O0, mod_dec, sib_dec, displc, imm_sz, pfx_sz, twobyte, fpu);
    output [5:0] O0;
    input  mod_dec;
    input  sib_dec;
    input [2:0] displc;
    input [2:0] imm_sz;
    input [4:0] pfx_sz;
    input  twobyte;
    input  fpu;
    // Line 404
    wire [5:0] N20;
    // Line 404
    wire [6:0] N26;
    // Line 211
    wire [5:0] O0;
    // Line 405
    wire [5:0] N36;
    // Line 404
    wire [7:0] N17;

    // Line 404
    assign N20 = N17 + imm_sz;
    // Line 404
    assign N26 = mod_dec + 7'h1 + N36;
    // Line 211
    assign O0 = N20;
    // Line 405
    assign N36 = pfx_sz + twobyte + fpu;
    // Line 404
    assign N17 = N26 + displc + sib_dec;
endmodule

module deco8(in8, indic);

	input [7:0] in8;
	output [72:0] indic;

	wire \indic[10] ;
	wire \indic[14] ;
	wire \indic[15] ;
	wire \indic[22] ;
	wire \indic[0] ;
	wire \indic[1] ;
	wire \indic[2] ;
	wire \indic[3] ;
	wire \indic[4] ;
	wire \indic[5] ;
	wire \indic[6] ;
	wire \indic[7] ;
	wire \indic[8] ;
	wire \indic[9] ;
	wire \indic[11] ;
	wire \indic[12] ;
	wire \indic[13] ;
	wire \indic[16] ;
	wire \indic[17] ;
	wire \indic[18] ;
	wire \indic[19] ;
	wire \indic[20] ;
	wire \indic[21] ;
	wire \indic[23] ;
	wire \indic[24] ;
	wire \indic[25] ;
	wire \indic[26] ;
	wire \indic[27] ;
	wire \indic[28] ;
	wire \indic[29] ;
	wire \indic[30] ;
	wire \indic[32] ;
	wire \indic[33] ;
	wire \indic[34] ;
	wire \indic[35] ;
	wire \indic[36] ;
	wire \indic[37] ;
	wire \indic[38] ;
	wire \indic[39] ;
	wire \indic[40] ;
	wire \indic[41] ;
	wire \indic[42] ;
	wire \indic[43] ;
	wire \indic[44] ;
	wire \indic[45] ;
	wire \indic[46] ;
	wire \indic[47] ;
	wire \indic[48] ;
	wire \indic[49] ;
	wire \indic[50] ;
	wire \indic[51] ;
	wire \indic[53] ;
	wire \indic[54] ;
	wire \indic[55] ;
	wire \indic[56] ;
	wire \indic[57] ;
	wire \indic[58] ;
	wire \indic[59] ;
	wire \indic[60] ;
	wire \indic[61] ;
	wire \indic[62] ;
	wire \indic[63] ;
	wire \indic[64] ;
	wire \indic[67] ;
	wire \indic[68] ;
	wire \indic[69] ;
	wire \indic[70] ;
	wire \indic[71] ;
	wire \indic[72] ;


	assign indic[10] = \indic[10] ;
	assign indic[14] = \indic[14] ;
	assign indic[15] = \indic[15] ;
	assign indic[22] = \indic[22] ;
	assign indic[0] = \indic[0] ;
	assign indic[1] = \indic[1] ;
	assign indic[2] = \indic[2] ;
	assign indic[3] = \indic[3] ;
	assign indic[4] = \indic[4] ;
	assign indic[5] = \indic[5] ;
	assign indic[6] = \indic[6] ;
	assign indic[7] = \indic[7] ;
	assign indic[8] = \indic[8] ;
	assign indic[9] = \indic[9] ;
	assign indic[11] = \indic[11] ;
	assign indic[12] = \indic[12] ;
	assign indic[13] = \indic[13] ;
	assign indic[16] = \indic[16] ;
	assign indic[17] = \indic[17] ;
	assign indic[18] = \indic[18] ;
	assign indic[19] = \indic[19] ;
	assign indic[20] = \indic[20] ;
	assign indic[21] = \indic[21] ;
	assign indic[23] = \indic[23] ;
	assign indic[24] = \indic[24] ;
	assign indic[25] = \indic[25] ;
	assign indic[26] = \indic[26] ;
	assign indic[27] = \indic[27] ;
	assign indic[28] = \indic[28] ;
	assign indic[29] = \indic[29] ;
	assign indic[30] = \indic[30] ;
	assign indic[32] = \indic[32] ;
	assign indic[33] = \indic[33] ;
	assign indic[34] = \indic[34] ;
	assign indic[66] = \indic[35] ;
	assign indic[35] = \indic[35] ;
	assign indic[36] = \indic[36] ;
	assign indic[37] = \indic[37] ;
	assign indic[38] = \indic[38] ;
	assign indic[39] = \indic[39] ;
	assign indic[40] = \indic[40] ;
	assign indic[52] = \indic[41] ;
	assign indic[41] = \indic[41] ;
	assign indic[42] = \indic[42] ;
	assign indic[43] = \indic[43] ;
	assign indic[44] = \indic[44] ;
	assign indic[45] = \indic[45] ;
	assign indic[46] = \indic[46] ;
	assign indic[47] = \indic[47] ;
	assign indic[48] = \indic[48] ;
	assign indic[49] = \indic[49] ;
	assign indic[65] = \indic[50] ;
	assign indic[50] = \indic[50] ;
	assign indic[51] = \indic[51] ;
	assign indic[53] = \indic[53] ;
	assign indic[54] = \indic[54] ;
	assign indic[55] = \indic[55] ;
	assign indic[56] = \indic[56] ;
	assign indic[57] = \indic[57] ;
	assign indic[58] = \indic[58] ;
	assign indic[59] = \indic[59] ;
	assign indic[60] = \indic[60] ;
	assign indic[61] = \indic[61] ;
	assign indic[62] = \indic[62] ;
	assign indic[63] = \indic[63] ;
	assign indic[64] = \indic[64] ;
	assign indic[67] = \indic[67] ;
	assign indic[68] = \indic[68] ;
	assign indic[69] = \indic[69] ;
	assign indic[70] = \indic[70] ;
	assign indic[71] = \indic[71] ;
	assign indic[72] = \indic[72] ;

	notech_and3 i_79(.A(in8[6]), .B(in8[7]), .C(n_75), .Z(n_102));
	notech_and3 i_77(.A(n_30638), .B(n_30639), .C(in8[3]), .Z(n_96));
	notech_and2 i_80(.A(n_30638), .B(n_30637), .Z(n_93));
	notech_and2 i_97(.A(n_30639), .B(n_30637), .Z(n_92));
	notech_and2 i_96(.A(in8[0]), .B(in8[2]), .Z(n_90));
	notech_and4 i_72(.A(in8[6]), .B(in8[7]), .C(in8[4]), .D(n_30641), .Z(n_88
		));
	notech_and3 i_69(.A(in8[6]), .B(in8[7]), .C(n_85), .Z(n_86));
	notech_nor2 i_78(.A(in8[4]), .B(in8[5]), .Z(n_85));
	notech_and2 i_86(.A(n_30637), .B(in8[2]), .Z(n_80));
	notech_and2 i_88(.A(n_78), .B(in8[1]), .Z(n_79));
	notech_nor2 i_71(.A(in8[7]), .B(in8[6]), .Z(n_78));
	notech_nor2 i_70(.A(in8[4]), .B(n_30641), .Z(n_75));
	notech_and3 i_15(.A(in8[0]), .B(in8[3]), .C(in8[2]), .Z(n_73));
	notech_and3 i_10(.A(n_30640), .B(in8[1]), .C(n_30639), .Z(n_72));
	notech_and2 i_23(.A(in8[6]), .B(in8[7]), .Z(n_71));
	notech_and2 i_14(.A(n_30640), .B(n_30639), .Z(n_70));
	notech_and4 i_116(.A(n_92), .B(in8[1]), .C(n_30641), .D(in8[3]), .Z(n_113
		));
	notech_nand3 i_119(.A(\indic[4] ), .B(n_30640), .C(in8[0]), .Z(n_116));
	notech_and4 i_071110(.A(n_71), .B(\indic[41] ), .C(n_30640), .D(n_30639)
		, .Z(\indic[0] ));
	notech_and4 i_1(.A(n_75), .B(\indic[24] ), .C(n_30640), .D(in8[2]), .Z(\indic[1] 
		));
	notech_and4 i_2(.A(n_80), .B(in8[3]), .C(in8[5]), .D(n_79), .Z(\indic[2] 
		));
	notech_and4 i_3(.A(\indic[6] ), .B(n_80), .C(n_78), .D(in8[5]), .Z(\indic[3] 
		));
	notech_and2 i_4(.A(n_78), .B(n_30639), .Z(\indic[4] ));
	notech_and3 i_5(.A(n_75), .B(\indic[24] ), .C(n_30639), .Z(\indic[5] )
		);
	notech_and2 i_6(.A(n_30640), .B(in8[1]), .Z(\indic[6] ));
	notech_and2 i_7(.A(in8[0]), .B(in8[3]), .Z(\indic[7] ));
	notech_ao3 i_8(.A(in8[7]), .B(n_85), .C(in8[6]), .Z(\indic[8] ));
	notech_and4 i_9(.A(in8[6]), .B(in8[7]), .C(n_85), .D(n_30640), .Z(\indic[9] 
		));
	notech_and4 i_11(.A(in8[4]), .B(n_71), .C(n_70), .D(n_30641), .Z(\indic[11] 
		));
	notech_and4 i_12(.A(n_71), .B(\indic[41] ), .C(in8[2]), .D(in8[1]), .Z(\indic[12] 
		));
	notech_ao3 i_13(.A(n_78), .B(n_30641), .C(in8[4]), .Z(\indic[13] ));
	notech_and3 i_16(.A(in8[4]), .B(n_78), .C(in8[5]), .Z(\indic[16] ));
	notech_and4 i_17(.A(n_90), .B(\indic[28] ), .C(n_30640), .D(in8[1]), .Z(\indic[17] 
		));
	notech_ao3 i_18(.A(in8[7]), .B(n_75), .C(in8[6]), .Z(\indic[18] ));
	notech_and2 i_19(.A(n_30638), .B(n_30639), .Z(\indic[19] ));
	notech_and3 i_20(.A(n_30639), .B(n_30637), .C(in8[1]), .Z(\indic[60] )
		);
	notech_and4 i_21(.A(in8[6]), .B(in8[7]), .C(n_85), .D(in8[3]), .Z(\indic[20] 
		));
	notech_and3 i_22(.A(n_30638), .B(n_30637), .C(in8[2]), .Z(\indic[21] )
		);
	notech_and3 i_24(.A(n_78), .B(in8[0]), .C(in8[2]), .Z(\indic[23] ));
	notech_and2 i_25(.A(in8[6]), .B(n_30642), .Z(\indic[24] ));
	notech_nor2 i_26(.A(in8[6]), .B(n_30642), .Z(\indic[25] ));
	notech_and4 i_27(.A(n_78), .B(n_30638), .C(n_30637), .D(in8[2]), .Z(\indic[26] 
		));
	notech_and3 i_28(.A(in8[3]), .B(\indic[5] ), .C(in8[1]), .Z(\indic[27] )
		);
	notech_and3 i_29(.A(in8[4]), .B(\indic[24] ), .C(in8[5]), .Z(\indic[28] 
		));
	notech_ao3 i_30(.A(\indic[43] ), .B(n_30638), .C(in8[0]), .Z(\indic[29] 
		));
	notech_and4 i_31(.A(n_85), .B(in8[0]), .C(\indic[25] ), .D(n_72), .Z(\indic[30] 
		));
	notech_ao3 i_32(.A(\indic[18] ), .B(n_96), .C(in8[0]), .Z(\indic[32] )
		);
	notech_and4 i_33(.A(in8[4]), .B(\indic[25] ), .C(in8[5]), .D(n_30640), .Z
		(\indic[33] ));
	notech_and4 i_34(.A(n_71), .B(n_85), .C(n_70), .D(n_30638), .Z(\indic[34] 
		));
	notech_and3 i_35(.A(n_73), .B(n_86), .C(n_30638), .Z(\indic[36] ));
	notech_and4 i_36(.A(in8[2]), .B(n_30638), .C(n_88), .D(n_30640), .Z(\indic[37] 
		));
	notech_ao3 i_37(.A(n_71), .B(n_75), .C(in8[3]), .Z(\indic[38] ));
	notech_and4 i_38(.A(n_102), .B(in8[1]), .C(\indic[7] ), .D(n_30639), .Z(\indic[39] 
		));
	notech_and4 i_39(.A(\indic[6] ), .B(n_71), .C(\indic[41] ), .D(n_80), .Z
		(\indic[40] ));
	notech_and4 i_40(.A(n_86), .B(n_30639), .C(n_30637), .D(in8[1]), .Z(\indic[42] 
		));
	notech_and4 i_41(.A(\indic[25] ), .B(n_85), .C(n_30640), .D(n_30639), .Z
		(\indic[43] ));
	notech_and4 i_42(.A(n_78), .B(in8[0]), .C(in8[2]), .D(n_30638), .Z(\indic[44] 
		));
	notech_and4 i_43(.A(in8[4]), .B(\indic[25] ), .C(in8[5]), .D(in8[3]), .Z
		(\indic[45] ));
	notech_and4 i_44(.A(in8[6]), .B(in8[7]), .C(n_75), .D(n_96), .Z(\indic[46] 
		));
	notech_and3 i_45(.A(n_75), .B(\indic[24] ), .C(n_96), .Z(\indic[47] ));
	notech_and4 i_46(.A(\indic[25] ), .B(n_75), .C(n_30640), .D(n_30639), .Z
		(\indic[48] ));
	notech_and3 i_47(.A(\indic[25] ), .B(n_96), .C(in8[5]), .Z(\indic[49] )
		);
	notech_and4 i_48(.A(\indic[6] ), .B(n_71), .C(\indic[41] ), .D(n_90), .Z
		(\indic[51] ));
	notech_and2 i_49(.A(in8[4]), .B(in8[5]), .Z(\indic[41] ));
	notech_and3 i_50(.A(\indic[45] ), .B(in8[1]), .C(n_92), .Z(\indic[53] )
		);
	notech_and4 i_51(.A(n_85), .B(n_78), .C(in8[1]), .D(n_73), .Z(\indic[54] 
		));
	notech_and4 i_52(.A(n_93), .B(\indic[41] ), .C(\indic[24] ), .D(n_70), .Z
		(\indic[55] ));
	notech_ao3 i_53(.A(\indic[18] ), .B(\indic[21] ), .C(in8[3]), .Z(\indic[56] 
		));
	notech_ao3 i_54(.A(n_72), .B(n_86), .C(in8[0]), .Z(\indic[57] ));
	notech_and3 i_55(.A(in8[2]), .B(\indic[9] ), .C(n_93), .Z(\indic[58] )
		);
	notech_and4 i_56(.A(in8[0]), .B(in8[2]), .C(\indic[9] ), .D(n_30638), .Z
		(\indic[59] ));
	notech_and4 i_57(.A(in8[4]), .B(n_71), .C(in8[3]), .D(n_30641), .Z(\indic[61] 
		));
	notech_and4 i_58(.A(n_75), .B(\indic[24] ), .C(\indic[6] ), .D(n_80), .Z
		(\indic[62] ));
	notech_and4 i_59(.A(\indic[6] ), .B(n_71), .C(\indic[41] ), .D(n_30639),
		 .Z(\indic[63] ));
	notech_and4 i_60(.A(n_92), .B(in8[3]), .C(n_102), .D(in8[1]), .Z(\indic[64] 
		));
	notech_and4 i_61(.A(\indic[6] ), .B(n_86), .C(in8[0]), .D(in8[2]), .Z(\indic[50] 
		));
	notech_and4 i_62(.A(n_86), .B(n_30637), .C(in8[2]), .D(\indic[6] ), .Z(\indic[35] 
		));
	notech_and4 i_63(.A(\indic[6] ), .B(n_90), .C(n_75), .D(\indic[24] ), .Z
		(\indic[67] ));
	notech_and3 i_64(.A(in8[4]), .B(\indic[25] ), .C(n_113), .Z(\indic[68] )
		);
	notech_ao3 i_65(.A(n_85), .B(n_30638), .C(n_116), .Z(\indic[69] ));
	notech_and4 i_66(.A(\indic[18] ), .B(n_30638), .C(n_30637), .D(in8[2]), 
		.Z(\indic[70] ));
	notech_and4 i_67(.A(n_72), .B(\indic[25] ), .C(n_85), .D(n_30637), .Z(\indic[71] 
		));
	notech_and4 i_68(.A(n_72), .B(\indic[41] ), .C(\indic[25] ), .D(n_30637)
		, .Z(\indic[72] ));
	notech_inv i_34617(.A(in8[0]), .Z(n_30637));
	notech_inv i_34618(.A(in8[1]), .Z(n_30638));
	notech_inv i_34619(.A(in8[2]), .Z(n_30639));
	notech_inv i_34620(.A(in8[3]), .Z(n_30640));
	notech_inv i_34621(.A(in8[5]), .Z(n_30641));
	notech_inv i_34622(.A(in8[7]), .Z(n_30642));
	notech_inv i_34623(.A(n_70), .Z(\indic[14] ));
	notech_inv i_34624(.A(n_71), .Z(\indic[22] ));
	notech_inv i_34625(.A(n_72), .Z(\indic[10] ));
	notech_inv i_34626(.A(n_73), .Z(\indic[15] ));
endmodule
module deco_rm(in8, indic);

	input [7:0] in8;
	output [7:0] indic;




	notech_nand2 i_1(.A(in8[7]), .B(in8[6]), .Z(indic[1]));
	notech_and3 i_071111(.A(in8[2]), .B(n_30649), .C(n_30648), .Z(indic[0])
		);
	notech_and4 i_2(.A(in8[2]), .B(in8[0]), .C(indic[7]), .D(n_30648), .Z(indic
		[2]));
	notech_and2 i_3(.A(in8[7]), .B(n_30647), .Z(indic[3]));
	notech_nor2 i_4(.A(in8[7]), .B(n_30647), .Z(indic[4]));
	notech_nor2 i_5(.A(in8[5]), .B(in8[4]), .Z(indic[5]));
	notech_and4 i_6(.A(indic[7]), .B(in8[2]), .C(in8[1]), .D(n_30649), .Z(indic
		[6]));
	notech_nor2 i_7(.A(in8[7]), .B(in8[6]), .Z(indic[7]));
	notech_inv i_34636(.A(in8[6]), .Z(n_30647));
	notech_inv i_34637(.A(in8[1]), .Z(n_30648));
	notech_inv i_34638(.A(in8[0]), .Z(n_30649));
endmodule
module udecox(op, modrm, twobyte, cpl, adz, opz, jsz, udeco, fpu, emul, ipg_fault
		);

	input [7:0] op;
	input [7:0] modrm;
	input twobyte;
	input [1:0] cpl;
	input adz;
	input [2:0] opz;
	input [3:0] jsz;
	output [127:0] udeco;
	input fpu;
	input emul;
	input ipg_fault;

	wire n_4024;
	wire \udeco[0] ;
	wire \udeco[1] ;
	wire \udeco[2] ;
	wire \udeco[3] ;
	wire \udeco[4] ;
	wire \udeco[5] ;
	wire \udeco[6] ;
	wire \udeco[8] ;
	wire \udeco[9] ;
	wire \udeco[10] ;
	wire \udeco[11] ;
	wire \udeco[12] ;
	wire \udeco[13] ;
	wire \udeco[14] ;
	wire \udeco[15] ;
	wire \udeco[16] ;
	wire \udeco[17] ;
	wire \udeco[18] ;
	wire \udeco[19] ;
	wire \udeco[20] ;
	wire \udeco[21] ;
	wire \udeco[22] ;
	wire \udeco[23] ;
	wire \udeco[24] ;
	wire \udeco[25] ;
	wire \udeco[26] ;
	wire \udeco[27] ;
	wire \udeco[28] ;
	wire \udeco[29] ;
	wire \udeco[30] ;
	wire \udeco[31] ;
	wire \udeco[32] ;
	wire \udeco[33] ;
	wire \udeco[34] ;
	wire \udeco[35] ;
	wire \udeco[36] ;
	wire \udeco[37] ;
	wire \udeco[38] ;
	wire \udeco[39] ;
	wire \udeco[40] ;
	wire \udeco[41] ;
	wire \udeco[42] ;
	wire \udeco[43] ;
	wire \udeco[44] ;
	wire \udeco[45] ;
	wire \udeco[46] ;
	wire \udeco[47] ;
	wire \udeco[48] ;
	wire \udeco[49] ;
	wire \udeco[50] ;
	wire \udeco[51] ;
	wire \udeco[52] ;
	wire \udeco[53] ;
	wire \udeco[54] ;
	wire \udeco[55] ;
	wire \udeco[56] ;
	wire \udeco[57] ;
	wire \udeco[58] ;
	wire \udeco[59] ;
	wire \udeco[60] ;
	wire \udeco[61] ;
	wire \udeco[62] ;
	wire \udeco[63] ;
	wire \udeco[64] ;
	wire \udeco[65] ;
	wire \udeco[66] ;
	wire \udeco[67] ;
	wire \udeco[68] ;
	wire \udeco[69] ;
	wire \udeco[70] ;
	wire \udeco[71] ;
	wire \udeco[72] ;
	wire \udeco[73] ;
	wire \udeco[74] ;
	wire \udeco[75] ;
	wire \udeco[77] ;
	wire \udeco[78] ;
	wire \udeco[80] ;
	wire \udeco[81] ;
	wire \udeco[82] ;
	wire \udeco[83] ;
	wire \udeco[84] ;
	wire \udeco[85] ;
	wire \udeco[86] ;
	wire \udeco[87] ;
	wire \udeco[88] ;
	wire \udeco[89] ;
	wire \udeco[90] ;
	wire \udeco[91] ;
	wire \udeco[92] ;
	wire \udeco[93] ;
	wire \udeco[95] ;
	wire \udeco[96] ;
	wire \udeco[98] ;
	wire \udeco[99] ;
	wire \udeco[100] ;
	wire \udeco[101] ;
	wire \udeco[102] ;
	wire \udeco[103] ;
	wire \udeco[104] ;
	wire \udeco[105] ;
	wire \udeco[106] ;
	wire \udeco[107] ;
	wire \udeco[108] ;
	wire \udeco[109] ;
	wire \udeco[110] ;
	wire \udeco[112] ;
	wire \udeco[113] ;
	wire \udeco[114] ;
	wire \udeco[115] ;
	wire \udeco[116] ;
	wire \udeco[117] ;
	wire \udeco[118] ;
	wire \udeco[119] ;
	wire \udeco[120] ;
	wire \udeco[121] ;
	wire \udeco[122] ;
	wire \udeco[123] ;
	wire \udeco[124] ;
	wire \udeco[125] ;
	wire \udeco[126] ;
	wire \udeco[127] ;


	assign udeco[111] = n_4024;
	assign udeco[0] = \udeco[0] ;
	assign udeco[1] = \udeco[1] ;
	assign udeco[2] = \udeco[2] ;
	assign udeco[3] = \udeco[3] ;
	assign udeco[4] = \udeco[4] ;
	assign udeco[5] = \udeco[5] ;
	assign udeco[7] = \udeco[6] ;
	assign udeco[6] = \udeco[6] ;
	assign udeco[8] = \udeco[8] ;
	assign udeco[9] = \udeco[9] ;
	assign udeco[10] = \udeco[10] ;
	assign udeco[11] = \udeco[11] ;
	assign udeco[12] = \udeco[12] ;
	assign udeco[13] = \udeco[13] ;
	assign udeco[14] = \udeco[14] ;
	assign udeco[15] = \udeco[15] ;
	assign udeco[16] = \udeco[16] ;
	assign udeco[17] = \udeco[17] ;
	assign udeco[18] = \udeco[18] ;
	assign udeco[19] = \udeco[19] ;
	assign udeco[20] = \udeco[20] ;
	assign udeco[21] = \udeco[21] ;
	assign udeco[22] = \udeco[22] ;
	assign udeco[23] = \udeco[23] ;
	assign udeco[24] = \udeco[24] ;
	assign udeco[25] = \udeco[25] ;
	assign udeco[26] = \udeco[26] ;
	assign udeco[27] = \udeco[27] ;
	assign udeco[28] = \udeco[28] ;
	assign udeco[29] = \udeco[29] ;
	assign udeco[30] = \udeco[30] ;
	assign udeco[31] = \udeco[31] ;
	assign udeco[32] = \udeco[32] ;
	assign udeco[33] = \udeco[33] ;
	assign udeco[34] = \udeco[34] ;
	assign udeco[35] = \udeco[35] ;
	assign udeco[36] = \udeco[36] ;
	assign udeco[37] = \udeco[37] ;
	assign udeco[38] = \udeco[38] ;
	assign udeco[39] = \udeco[39] ;
	assign udeco[40] = \udeco[40] ;
	assign udeco[41] = \udeco[41] ;
	assign udeco[42] = \udeco[42] ;
	assign udeco[43] = \udeco[43] ;
	assign udeco[44] = \udeco[44] ;
	assign udeco[45] = \udeco[45] ;
	assign udeco[46] = \udeco[46] ;
	assign udeco[47] = \udeco[47] ;
	assign udeco[48] = \udeco[48] ;
	assign udeco[49] = \udeco[49] ;
	assign udeco[50] = \udeco[50] ;
	assign udeco[51] = \udeco[51] ;
	assign udeco[52] = \udeco[52] ;
	assign udeco[53] = \udeco[53] ;
	assign udeco[54] = \udeco[54] ;
	assign udeco[55] = \udeco[55] ;
	assign udeco[56] = \udeco[56] ;
	assign udeco[57] = \udeco[57] ;
	assign udeco[58] = \udeco[58] ;
	assign udeco[59] = \udeco[59] ;
	assign udeco[60] = \udeco[60] ;
	assign udeco[61] = \udeco[61] ;
	assign udeco[62] = \udeco[62] ;
	assign udeco[63] = \udeco[63] ;
	assign udeco[64] = \udeco[64] ;
	assign udeco[65] = \udeco[65] ;
	assign udeco[66] = \udeco[66] ;
	assign udeco[67] = \udeco[67] ;
	assign udeco[68] = \udeco[68] ;
	assign udeco[69] = \udeco[69] ;
	assign udeco[70] = \udeco[70] ;
	assign udeco[71] = \udeco[71] ;
	assign udeco[72] = \udeco[72] ;
	assign udeco[73] = \udeco[73] ;
	assign udeco[76] = \udeco[74] ;
	assign udeco[74] = \udeco[74] ;
	assign udeco[75] = \udeco[75] ;
	assign udeco[77] = \udeco[77] ;
	assign udeco[79] = \udeco[78] ;
	assign udeco[78] = \udeco[78] ;
	assign udeco[80] = \udeco[80] ;
	assign udeco[81] = \udeco[81] ;
	assign udeco[82] = \udeco[82] ;
	assign udeco[83] = \udeco[83] ;
	assign udeco[84] = \udeco[84] ;
	assign udeco[85] = \udeco[85] ;
	assign udeco[86] = \udeco[86] ;
	assign udeco[87] = \udeco[87] ;
	assign udeco[88] = \udeco[88] ;
	assign udeco[89] = \udeco[89] ;
	assign udeco[90] = \udeco[90] ;
	assign udeco[91] = \udeco[91] ;
	assign udeco[92] = \udeco[92] ;
	assign udeco[94] = \udeco[93] ;
	assign udeco[93] = \udeco[93] ;
	assign udeco[95] = \udeco[95] ;
	assign udeco[96] = \udeco[96] ;
	assign udeco[98] = \udeco[98] ;
	assign udeco[99] = \udeco[99] ;
	assign udeco[97] = \udeco[100] ;
	assign udeco[100] = \udeco[100] ;
	assign udeco[101] = \udeco[101] ;
	assign udeco[102] = \udeco[102] ;
	assign udeco[103] = \udeco[103] ;
	assign udeco[104] = \udeco[104] ;
	assign udeco[105] = \udeco[105] ;
	assign udeco[106] = \udeco[106] ;
	assign udeco[107] = \udeco[107] ;
	assign udeco[108] = \udeco[108] ;
	assign udeco[109] = \udeco[109] ;
	assign udeco[110] = \udeco[110] ;
	assign udeco[112] = \udeco[112] ;
	assign udeco[113] = \udeco[113] ;
	assign udeco[114] = \udeco[114] ;
	assign udeco[115] = \udeco[115] ;
	assign udeco[116] = \udeco[116] ;
	assign udeco[117] = \udeco[117] ;
	assign udeco[118] = \udeco[118] ;
	assign udeco[119] = \udeco[119] ;
	assign udeco[120] = \udeco[120] ;
	assign udeco[121] = \udeco[121] ;
	assign udeco[122] = \udeco[122] ;
	assign udeco[123] = \udeco[123] ;
	assign udeco[124] = \udeco[124] ;
	assign udeco[125] = \udeco[125] ;
	assign udeco[126] = \udeco[126] ;
	assign udeco[127] = \udeco[127] ;

	notech_inv i_11674(.A(n_58596), .Z(n_58601));
	notech_inv i_11670(.A(n_58596), .Z(n_58597));
	notech_inv i_11669(.A(op[0]), .Z(n_58596));
	notech_inv i_11666(.A(n_58585), .Z(n_58592));
	notech_inv i_11665(.A(n_58585), .Z(n_58591));
	notech_inv i_11660(.A(n_58585), .Z(n_58586));
	notech_inv i_11659(.A(op[3]), .Z(n_58585));
	notech_inv i_11656(.A(n_58572), .Z(n_58581));
	notech_inv i_11652(.A(n_58572), .Z(n_58577));
	notech_inv i_11648(.A(n_58572), .Z(n_58573));
	notech_inv i_11647(.A(op[6]), .Z(n_58572));
	notech_inv i_11644(.A(n_58563), .Z(n_58568));
	notech_inv i_11640(.A(n_58563), .Z(n_58564));
	notech_inv i_11639(.A(op[5]), .Z(n_58563));
	notech_inv i_11632(.A(n_58554), .Z(n_58555));
	notech_inv i_11631(.A(n_30845), .Z(n_58554));
	notech_inv i_11628(.A(n_58545), .Z(n_58550));
	notech_inv i_11624(.A(n_58545), .Z(n_58546));
	notech_inv i_11623(.A(op[4]), .Z(n_58545));
	notech_inv i_11616(.A(n_58536), .Z(n_58537));
	notech_inv i_11615(.A(n_30844), .Z(n_58536));
	notech_inv i_11612(.A(n_58527), .Z(n_58532));
	notech_inv i_11608(.A(n_58527), .Z(n_58528));
	notech_inv i_11607(.A(op[1]), .Z(n_58527));
	notech_inv i_11600(.A(n_58518), .Z(n_58519));
	notech_inv i_11599(.A(n_30841), .Z(n_58518));
	notech_inv i_11596(.A(n_58509), .Z(n_58514));
	notech_inv i_11592(.A(n_58509), .Z(n_58510));
	notech_inv i_11591(.A(op[2]), .Z(n_58509));
	notech_inv i_11582(.A(n_58486), .Z(n_58498));
	notech_inv i_11581(.A(n_58486), .Z(n_58497));
	notech_inv i_11576(.A(n_58486), .Z(n_58492));
	notech_inv i_11571(.A(n_58486), .Z(n_58487));
	notech_inv i_11570(.A(n_2328), .Z(n_58486));
	notech_inv i_11567(.A(n_58597), .Z(n_58482));
	notech_inv i_11566(.A(n_58597), .Z(n_58481));
	notech_inv i_11561(.A(n_58597), .Z(n_58476));
	notech_inv i_11556(.A(n_58591), .Z(n_58470));
	notech_inv i_11551(.A(n_58591), .Z(n_58465));
	notech_inv i_11543(.A(n_58455), .Z(n_58456));
	notech_inv i_11542(.A(n_30842), .Z(n_58455));
	notech_inv i_11516(.A(n_58425), .Z(n_58426));
	notech_inv i_11515(.A(modrm[5]), .Z(n_58425));
	notech_inv i_11508(.A(n_58416), .Z(n_58417));
	notech_inv i_11507(.A(n_2271), .Z(n_58416));
	notech_inv i_11500(.A(n_58407), .Z(n_58408));
	notech_inv i_11499(.A(n_2360), .Z(n_58407));
	notech_inv i_11492(.A(n_58398), .Z(n_58399));
	notech_inv i_11491(.A(n_30659), .Z(n_58398));
	notech_inv i_11484(.A(n_58389), .Z(n_58390));
	notech_inv i_11483(.A(n_30851), .Z(n_58389));
	notech_inv i_11476(.A(n_58380), .Z(n_58381));
	notech_inv i_11475(.A(n_2325), .Z(n_58380));
	notech_inv i_11468(.A(n_58371), .Z(n_58372));
	notech_inv i_11467(.A(n_2286), .Z(n_58371));
	notech_inv i_11460(.A(n_58362), .Z(n_58363));
	notech_inv i_11459(.A(n_2282), .Z(n_58362));
	notech_inv i_11452(.A(n_58353), .Z(n_58354));
	notech_inv i_11451(.A(n_2410), .Z(n_58353));
	notech_and4 i_1531(.A(n_2839), .B(n_1543), .C(n_2931), .D(n_2924), .Z(n_2934
		));
	notech_ao3 i_1534(.A(n_2934), .B(n_2904), .C(n_30759), .Z(n_2936));
	notech_and2 i_793(.A(n_2179), .B(n_1603), .Z(n_2937));
	notech_and4 i_1535(.A(n_2663), .B(n_2352), .C(n_2937), .D(n_2567), .Z(n_2939
		));
	notech_and4 i_1546(.A(n_3993), .B(n_4040), .C(n_3733), .D(n_1907), .Z(n_2942
		));
	notech_and4 i_306(.A(n_2137), .B(n_2942), .C(n_2026), .D(n_3984), .Z(n_2945
		));
	notech_and3 i_770(.A(n_2638), .B(n_2014), .C(n_1896), .Z(n_2946));
	notech_and4 i_1552(.A(n_4019), .B(n_2080), .C(n_2945), .D(n_2946), .Z(n_2949
		));
	notech_and4 i_1557(.A(n_2189), .B(n_2206), .C(n_2028), .D(n_2457), .Z(n_2953
		));
	notech_and4 i_245(.A(n_2611), .B(n_2949), .C(n_2953), .D(n_2484), .Z(n_2955
		));
	notech_and4 i_1561(.A(n_2435), .B(n_2631), .C(n_1953), .D(n_2030), .Z(n_2958
		));
	notech_and4 i_303(.A(n_2141), .B(n_4013), .C(n_2058), .D(n_2958), .Z(n_2959
		));
	notech_and3 i_1569(.A(n_2033), .B(n_2032), .C(n_4020), .Z(n_2961));
	notech_and4 i_1572(.A(n_2176), .B(n_1837), .C(n_2034), .D(n_2961), .Z(n_2964
		));
	notech_and4 i_724(.A(n_2332), .B(n_2964), .C(n_2091), .D(n_3972), .Z(n_2967
		));
	notech_and4 i_521(.A(n_30726), .B(n_30691), .C(n_30725), .D(n_2031), .Z(n_2969
		));
	notech_ao4 i_1576(.A(n_3963), .B(n_2574), .C(n_2362), .D(n_2331), .Z(n_2970
		));
	notech_and4 i_1578(.A(n_3992), .B(n_1895), .C(n_2970), .D(n_3672), .Z(n_2972
		));
	notech_and4 i_1581(.A(n_2972), .B(n_2406), .C(n_2969), .D(n_2967), .Z(n_2975
		));
	notech_ao3 i_653(.A(n_2668), .B(n_3777), .C(n_30663), .Z(n_2978));
	notech_and4 i_1607(.A(n_843), .B(n_1332), .C(n_2494), .D(n_2046), .Z(n_2983
		));
	notech_and3 i_1611(.A(n_3994), .B(n_2983), .C(n_1340), .Z(n_2985));
	notech_and4 i_1615(.A(n_1329), .B(n_2021), .C(n_2562), .D(n_2985), .Z(n_2987
		));
	notech_ao4 i_510(.A(n_2098), .B(n_2101), .C(n_4065), .D(n_2027), .Z(n_2988
		));
	notech_ao4 i_1598(.A(n_30729), .B(n_30776), .C(adz), .D(n_2305), .Z(n_2989
		));
	notech_and4 i_1596(.A(n_2040), .B(n_2219), .C(n_30713), .D(n_2041), .Z(n_2992
		));
	notech_and4 i_1600(.A(n_2042), .B(n_2045), .C(n_2989), .D(n_2992), .Z(n_2995
		));
	notech_and4 i_1603(.A(n_2195), .B(n_4022), .C(n_2995), .D(n_1346), .Z(n_2999
		));
	notech_and4 i_1610(.A(n_2050), .B(n_2999), .C(n_2051), .D(n_2053), .Z(n_3002
		));
	notech_and4 i_1616(.A(n_3002), .B(n_1728), .C(n_2665), .D(n_2246), .Z(n_3005
		));
	notech_ao4 i_1633(.A(n_30729), .B(n_2574), .C(n_30787), .D(n_2355), .Z(n_3008
		));
	notech_ao3 i_1635(.A(n_2829), .B(n_3008), .C(n_3820), .Z(n_3010));
	notech_and4 i_244(.A(n_2392), .B(n_2967), .C(n_3955), .D(n_3010), .Z(n_3013
		));
	notech_and4 i_1640(.A(n_2435), .B(n_2631), .C(n_1526), .D(n_4025), .Z(n_3015
		));
	notech_and4 i_1643(.A(n_3015), .B(n_2379), .C(n_2852), .D(n_1905), .Z(n_3018
		));
	notech_and2 i_726(.A(n_3890), .B(n_2238), .Z(n_3021));
	notech_and4 i_1656(.A(n_1855), .B(n_1854), .C(n_4028), .D(n_2071), .Z(n_3023
		));
	notech_and4 i_1662(.A(n_2073), .B(n_3023), .C(n_1656), .D(n_2076), .Z(n_3026
		));
	notech_ao3 i_1669(.A(n_3026), .B(n_3021), .C(n_2077), .Z(n_3028));
	notech_and3 i_176(.A(n_4026), .B(n_1284), .C(n_4027), .Z(n_3030));
	notech_and4 i_1672(.A(n_3977), .B(n_1306), .C(n_3030), .D(n_3028), .Z(n_3033
		));
	notech_and4 i_1653(.A(n_2252), .B(n_222294221), .C(n_2188), .D(n_2070), 
		.Z(n_3039));
	notech_and4 i_1659(.A(n_2190), .B(n_3039), .C(n_2709), .D(n_2072), .Z(n_3042
		));
	notech_and4 i_1668(.A(n_3042), .B(n_4029), .C(n_2074), .D(n_1290), .Z(n_3045
		));
	notech_and4 i_1671(.A(n_3045), .B(n_2075), .C(n_2598), .D(n_4005), .Z(n_3046
		));
	notech_and4 i_1675(.A(n_4055), .B(n_1857), .C(n_3046), .D(n_3033), .Z(n_3048
		));
	notech_and2 i_549(.A(n_2264), .B(n_1911), .Z(n_3049));
	notech_and4 i_1677(.A(n_3049), .B(n_3048), .C(n_2789), .D(n_30664), .Z(n_3052
		));
	notech_and4 i_1679(.A(n_1329), .B(n_2021), .C(n_2826), .D(n_3052), .Z(n_3054
		));
	notech_and3 i_210(.A(n_4027), .B(n_4036), .C(n_4076), .Z(n_3056));
	notech_and4 i_1720(.A(n_2151), .B(n_3992), .C(n_3977), .D(n_30699), .Z(n_3059
		));
	notech_and2 i_624(.A(n_4017), .B(n_4019), .Z(n_3061));
	notech_and3 i_556(.A(n_2192), .B(n_4017), .C(n_3981), .Z(n_3062));
	notech_and4 i_1527(.A(n_1434), .B(n_2928), .C(n_30693), .D(n_4016), .Z(n_2931
		));
	notech_and3 i_206(.A(n_30712), .B(n_1958), .C(n_2377), .Z(n_3064));
	notech_ao4 i_1780(.A(n_30792), .B(n_58482), .C(n_30834), .D(n_30849), .Z
		(n_3067));
	notech_and3 i_1782(.A(n_3067), .B(n_2086), .C(n_3980), .Z(n_3069));
	notech_and4 i_1787(.A(n_4047), .B(n_223492236), .C(n_3069), .D(n_2305), 
		.Z(n_3072));
	notech_ao4 i_1788(.A(n_2124), .B(n_58470), .C(n_2333), .D(n_2359), .Z(n_3073
		));
	notech_and4 i_1792(.A(n_4017), .B(n_3073), .C(n_3072), .D(n_4019), .Z(n_3075
		));
	notech_and4 i_1799(.A(n_3075), .B(n_3967), .C(n_2090), .D(n_3064), .Z(n_3078
		));
	notech_and2 i_4702(.A(n_30695), .B(n_4082), .Z(n_3079));
	notech_and4 i_1789(.A(n_3079), .B(n_2087), .C(n_2089), .D(n_1624), .Z(n_3083
		));
	notech_and4 i_1795(.A(n_3083), .B(n_2579), .C(n_2609), .D(n_3981), .Z(n_3086
		));
	notech_and4 i_1800(.A(n_2663), .B(n_3086), .C(n_2978), .D(n_2091), .Z(n_3089
		));
	notech_and4 i_1803(.A(n_3089), .B(n_3078), .C(n_5254), .D(n_30720), .Z(n_3091
		));
	notech_and2 i_1808(.A(n_4040), .B(n_733), .Z(n_3095));
	notech_and4 i_258(.A(n_4002), .B(n_1332), .C(n_1329), .D(n_3095), .Z(n_3098
		));
	notech_ao3 i_809(.A(n_4055), .B(n_2097), .C(n_2100), .Z(n_3102));
	notech_ao4 i_560(.A(n_2499), .B(n_2485), .C(n_2596), .D(n_2302), .Z(n_3103
		));
	notech_and4 i_1821(.A(n_1984), .B(n_1801), .C(n_2159), .D(n_2104), .Z(n_3105
		));
	notech_and3 i_20373078(.A(n_2206), .B(n_4028), .C(n_2790), .Z(n_3107));
	notech_and3 i_296(.A(n_3965), .B(n_2579), .C(n_30723), .Z(n_2928));
	notech_and3 i_64773048(.A(n_2238), .B(n_4053), .C(n_2159), .Z(n_3109));
	notech_and4 i_1864(.A(n_3109), .B(n_222194220), .C(n_3107), .D(n_30728),
		 .Z(n_3111));
	notech_and4 i_1869(.A(n_3111), .B(n_2327), .C(n_2103), .D(n_30695), .Z(n_3114
		));
	notech_and4 i_1874(.A(n_30712), .B(n_4044), .C(n_3114), .D(n_4027), .Z(n_3117
		));
	notech_and4 i_1877(.A(n_2057), .B(n_1794), .C(n_2105), .D(n_3117), .Z(n_3119
		));
	notech_and4 i_1884(.A(n_3119), .B(n_2480), .C(n_2108), .D(n_2572), .Z(n_3122
		));
	notech_and2 i_719(.A(n_2218), .B(n_3970), .Z(n_3124));
	notech_and4 i_1887(.A(n_3970), .B(n_3122), .C(n_2218), .D(n_2116), .Z(n_3126
		));
	notech_ao3 i_317(.A(n_2609), .B(n_1792), .C(n_1795), .Z(n_3128));
	notech_and4 i_1871(.A(n_1932), .B(n_2123), .C(n_4041), .D(n_4043), .Z(n_3131
		));
	notech_and4 i_1879(.A(n_3131), .B(n_2107), .C(n_2104), .D(n_2106), .Z(n_3134
		));
	notech_and4 i_1883(.A(n_2176), .B(n_2195), .C(n_1970), .D(n_3134), .Z(n_3136
		));
	notech_and4 i_1888(.A(n_30797), .B(n_3128), .C(n_3136), .D(n_30693), .Z(n_3138
		));
	notech_and4 i_1891(.A(n_3098), .B(n_3126), .C(n_2109), .D(n_3138), .Z(n_3141
		));
	notech_and2 i_4754(.A(n_2688), .B(n_3739), .Z(n_3143));
	notech_and4 i_1924(.A(n_2579), .B(n_1970), .C(n_222894227), .D(n_2125), 
		.Z(n_3145));
	notech_and4 i_1917(.A(n_3061), .B(n_4032), .C(n_3981), .D(n_2122), .Z(n_3150
		));
	notech_and4 i_1919(.A(n_574), .B(n_4046), .C(n_2121), .D(n_3150), .Z(n_3151
		));
	notech_ao4 i_746(.A(n_2297), .B(n_2118), .C(n_2382), .D(n_2325), .Z(n_3152
		));
	notech_and4 i_444(.A(n_1855), .B(n_1854), .C(n_2111), .D(n_2255), .Z(n_3154
		));
	notech_and3 i_1904(.A(n_2119), .B(n_223492236), .C(n_30834), .Z(n_3157)
		);
	notech_and4 i_1908(.A(n_2627), .B(n_30695), .C(n_2364), .D(n_3157), .Z(n_3160
		));
	notech_and4 i_1910(.A(n_3154), .B(n_3160), .C(n_3992), .D(n_2120), .Z(n_3162
		));
	notech_and4 i_1918(.A(n_3152), .B(n_709), .C(n_3162), .D(n_2465), .Z(n_3165
		));
	notech_and4 i_1923(.A(n_673), .B(n_3165), .C(n_3151), .D(n_960), .Z(n_3168
		));
	notech_and4 i_1927(.A(n_3168), .B(n_703), .C(n_2126), .D(n_3145), .Z(n_3171
		));
	notech_nand2 i_441(.A(n_2625), .B(n_3779), .Z(n_3174));
	notech_and4 i_817(.A(n_2631), .B(n_1780), .C(n_2137), .D(n_30665), .Z(n_3177
		));
	notech_and3 i_811(.A(n_4058), .B(n_2049), .C(n_2129), .Z(n_3178));
	notech_and2 i_234(.A(n_3178), .B(n_2130), .Z(n_3179));
	notech_and3 i_1937(.A(n_2141), .B(n_2131), .C(n_30706), .Z(n_3181));
	notech_and4 i_1940(.A(n_2258), .B(n_3975), .C(n_3181), .D(n_30680), .Z(n_3184
		));
	notech_and3 i_1988(.A(n_3982), .B(n_30692), .C(n_455), .Z(n_3187));
	notech_and4 i_1981(.A(n_3977), .B(n_2377), .C(n_2134), .D(n_2978), .Z(n_3193
		));
	notech_and4 i_1986(.A(n_2218), .B(n_3970), .C(n_3193), .D(n_444), .Z(n_3195
		));
	notech_and3 i_37473064(.A(n_2104), .B(n_3154), .C(n_4046), .Z(n_3197));
	notech_ao4 i_1972(.A(n_2400), .B(n_2497), .C(n_2278), .D(n_2339), .Z(n_3200
		));
	notech_and4 i_1974(.A(n_3197), .B(n_2216), .C(n_4051), .D(n_3200), .Z(n_3201
		));
	notech_and4 i_1976(.A(n_30712), .B(n_4019), .C(n_3201), .D(n_1923), .Z(n_3204
		));
	notech_and4 i_1983(.A(n_3204), .B(n_2579), .C(n_2395), .D(n_3021), .Z(n_3207
		));
	notech_and4 i_1985(.A(n_4002), .B(n_1526), .C(n_3207), .D(n_2166), .Z(n_3208
		));
	notech_and4 i_1991(.A(n_2522), .B(n_3208), .C(n_3195), .D(n_2352), .Z(n_3211
		));
	notech_and4 i_1993(.A(n_3177), .B(n_3187), .C(n_3211), .D(n_2893), .Z(n_3213
		));
	notech_and4 i_2032(.A(n_2555), .B(n_1873), .C(n_3102), .D(n_3178), .Z(n_3217
		));
	notech_and4 i_2039(.A(n_3217), .B(n_2352), .C(n_2308), .D(n_2294), .Z(n_3219
		));
	notech_and4 i_2030(.A(n_3021), .B(n_2513), .C(n_3972), .D(n_2144), .Z(n_3223
		));
	notech_ao3 i_2013(.A(n_4028), .B(n_1829), .C(n_2142), .Z(n_3225));
	notech_and4 i_2007(.A(n_2433), .B(n_4048), .C(n_1263), .D(n_696), .Z(n_3227
		));
	notech_and4 i_2010(.A(n_2140), .B(n_4014), .C(n_2141), .D(n_3227), .Z(n_3230
		));
	notech_and4 i_2015(.A(n_3230), .B(n_4051), .C(n_3225), .D(n_30706), .Z(n_3233
		));
	notech_and4 i_2019(.A(n_1656), .B(n_4007), .C(n_3233), .D(n_30689), .Z(n_3236
		));
	notech_and3 i_2020(.A(n_1958), .B(n_4022), .C(n_30680), .Z(n_3240));
	notech_and4 i_2026(.A(n_3103), .B(n_3240), .C(n_2143), .D(n_30696), .Z(n_3243
		));
	notech_and4 i_2028(.A(n_3236), .B(n_3243), .C(n_3697), .D(n_2614), .Z(n_3244
		));
	notech_and4 i_2037(.A(n_3244), .B(n_466), .C(n_2854), .D(n_3223), .Z(n_3247
		));
	notech_and4 i_259(.A(n_3970), .B(n_2136), .C(n_2137), .D(n_1332), .Z(n_3250
		));
	notech_ao4 i_571(.A(n_2139), .B(n_30791), .C(n_2458), .D(n_2275), .Z(n_3252
		));
	notech_and4 i_2038(.A(n_3252), .B(n_3250), .C(n_2145), .D(n_455), .Z(n_3254
		));
	notech_and4 i_2042(.A(n_3254), .B(n_3247), .C(n_3219), .D(n_2834), .Z(n_3257
		));
	notech_ao4 i_171(.A(n_2278), .B(n_2154), .C(n_2318), .D(n_2161), .Z(n_3261
		));
	notech_and3 i_2073(.A(n_3970), .B(n_2166), .C(n_2168), .Z(n_3263));
	notech_and4 i_2082(.A(n_2065), .B(n_3261), .C(n_3263), .D(n_1623), .Z(n_3266
		));
	notech_and4 i_2091(.A(n_2538), .B(n_2663), .C(n_2173), .D(n_3266), .Z(n_3269
		));
	notech_and4 i_2097(.A(n_3979), .B(n_3269), .C(n_4032), .D(n_3984), .Z(n_3271
		));
	notech_and4 i_2105(.A(n_3271), .B(n_2526), .C(n_3179), .D(n_2175), .Z(n_3273
		));
	notech_and4 i_764(.A(n_2234), .B(n_4005), .C(n_2159), .D(n_4004), .Z(n_3275
		));
	notech_ao4 i_627(.A(n_30785), .B(n_2517), .C(n_3963), .D(n_2407), .Z(n_3276
		));
	notech_or4 i_98(.A(n_2403), .B(n_2311), .C(n_58514), .D(n_30841), .Z(n_3277
		));
	notech_and2 i_360473097(.A(n_1797), .B(n_2106), .Z(n_3279));
	notech_ao4 i_1502(.A(n_2140), .B(n_58601), .C(n_2433), .D(n_58592), .Z(n_2925
		));
	notech_and3 i_38273063(.A(n_1993), .B(n_2665), .C(n_3143), .Z(n_3280));
	notech_ao3 i_2067(.A(n_3280), .B(n_3279), .C(n_30825), .Z(n_3282));
	notech_and3 i_2068(.A(n_1925), .B(n_3107), .C(n_3282), .Z(n_3283));
	notech_and4 i_2072(.A(n_2516), .B(n_3283), .C(n_2163), .D(n_1828), .Z(n_3286
		));
	notech_and4 i_2079(.A(n_3286), .B(n_2170), .C(n_3276), .D(n_2169), .Z(n_3289
		));
	notech_ao4 i_777(.A(n_2495), .B(n_2376), .C(n_2337), .D(n_30702), .Z(n_3290
		));
	notech_and4 i_2083(.A(n_3290), .B(n_2076), .C(n_3289), .D(n_3890), .Z(n_3293
		));
	notech_and4 i_2087(.A(n_3975), .B(n_4037), .C(n_2172), .D(n_2174), .Z(n_3297
		));
	notech_and4 i_2092(.A(n_3293), .B(n_1526), .C(n_2639), .D(n_3297), .Z(n_3299
		));
	notech_and4 i_2103(.A(n_673), .B(n_3299), .C(n_3275), .D(n_3177), .Z(n_3302
		));
	notech_and4 i_2096(.A(n_3987), .B(n_2029), .C(n_3128), .D(n_1712), .Z(n_3307
		));
	notech_and4 i_2104(.A(n_3252), .B(n_3307), .C(n_2563), .D(n_497), .Z(n_3309
		));
	notech_ao4 i_2112(.A(n_2329), .B(n_2448), .C(n_2407), .D(n_2408), .Z(n_3312
		));
	notech_and2 i_2127(.A(n_2188), .B(n_4013), .Z(n_3316));
	notech_and4 i_2130(.A(n_2189), .B(n_2234), .C(n_2190), .D(n_3316), .Z(n_3319
		));
	notech_and4 i_2139(.A(n_2192), .B(n_3319), .C(n_4051), .D(n_3290), .Z(n_3322
		));
	notech_ao4 i_2131(.A(n_2278), .B(n_30800), .C(n_30777), .D(n_2531), .Z(n_3323
		));
	notech_and4 i_2140(.A(n_3323), .B(n_2631), .C(n_3276), .D(n_30686), .Z(n_3326
		));
	notech_and4 i_2150(.A(n_3326), .B(n_3322), .C(n_2196), .D(n_30723), .Z(n_3329
		));
	notech_and4 i_2138(.A(n_2193), .B(n_223492236), .C(n_2327), .D(n_30688),
		 .Z(n_3333));
	notech_and4 i_2147(.A(n_3333), .B(n_1892), .C(n_3672), .D(n_1806), .Z(n_3336
		));
	notech_and4 i_2154(.A(n_3329), .B(n_2380), .C(n_2377), .D(n_3336), .Z(n_3338
		));
	notech_and4 i_2162(.A(n_2198), .B(n_3056), .C(n_1970), .D(n_3338), .Z(n_3340
		));
	notech_and4 i_2172(.A(n_3340), .B(n_3728), .C(n_493), .D(n_2200), .Z(n_3343
		));
	notech_ao4 i_2144(.A(n_2186), .B(n_58470), .C(n_1819), .D(n_2285), .Z(n_3347
		));
	notech_and4 i_2152(.A(n_3347), .B(n_2195), .C(n_2639), .D(n_2565), .Z(n_3349
		));
	notech_and4 i_2160(.A(n_2723), .B(n_3349), .C(n_2533), .D(n_2197), .Z(n_3351
		));
	notech_and4 i_2167(.A(n_2663), .B(n_3351), .C(n_2945), .D(n_2183), .Z(n_3353
		));
	notech_and3 i_453(.A(n_4032), .B(n_2365), .C(n_2181), .Z(n_3355));
	notech_and4 i_2161(.A(n_4034), .B(n_2465), .C(n_4053), .D(n_1924), .Z(n_3358
		));
	notech_and4 i_1529(.A(n_2921), .B(n_2534), .C(n_2620), .D(n_2656), .Z(n_2924
		));
	notech_and3 i_3668(.A(n_4031), .B(n_4056), .C(n_30720), .Z(n_3360));
	notech_and4 i_2168(.A(n_497), .B(n_3358), .C(n_3360), .D(n_2199), .Z(n_3362
		));
	notech_and4 i_2173(.A(n_3362), .B(n_533), .C(n_3353), .D(n_3355), .Z(n_3364
		));
	notech_and3 i_2177(.A(n_2258), .B(n_3739), .C(n_2202), .Z(n_3367));
	notech_and4 i_375(.A(n_3049), .B(n_2790), .C(n_3367), .D(n_1905), .Z(n_3370
		));
	notech_and4 i_2203(.A(n_4005), .B(n_2532), .C(n_2218), .D(n_3779), .Z(n_3373
		));
	notech_ao4 i_488(.A(n_2412), .B(n_30801), .C(n_2455), .D(n_2297), .Z(n_3374
		));
	notech_and4 i_2195(.A(n_2637), .B(n_3374), .C(n_3965), .D(n_2207), .Z(n_3377
		));
	notech_and4 i_2186(.A(n_4048), .B(n_3109), .C(n_2516), .D(n_2206), .Z(n_3381
		));
	notech_and4 i_2189(.A(n_1855), .B(n_3381), .C(n_1854), .D(n_30688), .Z(n_3383
		));
	notech_and4 i_2192(.A(n_2668), .B(n_3383), .C(n_3973), .D(n_30685), .Z(n_3385
		));
	notech_and4 i_2199(.A(n_3385), .B(n_3377), .C(n_2305), .D(n_4056), .Z(n_3388
		));
	notech_ao4 i_815(.A(n_2205), .B(n_2285), .C(n_2331), .D(n_2586), .Z(n_3389
		));
	notech_and4 i_2202(.A(n_3777), .B(n_4055), .C(n_3389), .D(n_3388), .Z(n_3392
		));
	notech_and4 i_2205(.A(n_1796), .B(n_3392), .C(n_3373), .D(n_4029), .Z(n_3394
		));
	notech_and4 i_2208(.A(n_3250), .B(n_3394), .C(n_960), .D(n_3370), .Z(n_3397
		));
	notech_and2 i_408973096(.A(n_4079), .B(n_1984), .Z(n_3402));
	notech_and4 i_59973055(.A(n_2192), .B(n_2305), .C(n_30706), .D(n_30685),
		 .Z(n_3403));
	notech_and4 i_2219(.A(n_3403), .B(n_3402), .C(n_4048), .D(n_2668), .Z(n_3406
		));
	notech_and4 i_2222(.A(n_4058), .B(n_3406), .C(n_3838), .D(n_2216), .Z(n_3408
		));
	notech_and4 i_2225(.A(n_3408), .B(n_4029), .C(n_2217), .D(n_730), .Z(n_3411
		));
	notech_and4 i_2228(.A(n_2218), .B(n_3411), .C(n_3030), .D(n_3981), .Z(n_3413
		));
	notech_and4 i_2232(.A(n_3413), .B(n_2538), .C(n_2111), .D(n_30693), .Z(n_3415
		));
	notech_and4 i_2233(.A(n_2395), .B(n_218), .C(n_4049), .D(n_2411), .Z(n_3419
		));
	notech_and4 i_2236(.A(n_2534), .B(n_3415), .C(n_3250), .D(n_3419), .Z(n_3421
		));
	notech_ao4 i_2214(.A(n_30785), .B(n_2594), .C(n_2391), .D(n_30702), .Z(n_3422
		));
	notech_and4 i_2239(.A(n_204), .B(n_3421), .C(n_3370), .D(n_2379), .Z(n_3425
		));
	notech_and4 i_2281(.A(n_3994), .B(n_204), .C(n_3370), .D(n_4085), .Z(n_3429
		));
	notech_ao4 i_2258(.A(n_2678), .B(n_30845), .C(n_2485), .D(n_2689), .Z(n_3430
		));
	notech_and4 i_2261(.A(n_2631), .B(n_3374), .C(n_3430), .D(n_2222), .Z(n_3433
		));
	notech_and4 i_2253(.A(n_3998), .B(n_2220), .C(n_3402), .D(n_30724), .Z(n_3437
		));
	notech_and4 i_2257(.A(n_2221), .B(n_2130), .C(n_2223), .D(n_3437), .Z(n_3440
		));
	notech_and4 i_2264(.A(n_3975), .B(n_3103), .C(n_3389), .D(n_3440), .Z(n_3443
		));
	notech_and4 i_2268(.A(n_3433), .B(n_3443), .C(n_2116), .D(n_30699), .Z(n_3445
		));
	notech_and4 i_2269(.A(n_3030), .B(n_1130), .C(n_2695), .D(n_2854), .Z(n_3449
		));
	notech_and4 i_2274(.A(n_2675), .B(n_3449), .C(n_3445), .D(n_30694), .Z(n_3451
		));
	notech_and4 i_2272(.A(n_2076), .B(n_2080), .C(n_3275), .D(n_30680), .Z(n_3452
		));
	notech_and4 i_2278(.A(n_444), .B(n_960), .C(n_2722), .D(n_2226), .Z(n_3457
		));
	notech_and4 i_2280(.A(n_2534), .B(n_3452), .C(n_3451), .D(n_3457), .Z(n_3458
		));
	notech_and4 i_2326(.A(n_2294), .B(n_2587), .C(n_1340), .D(n_2228), .Z(n_3463
		));
	notech_and4 i_2330(.A(n_3994), .B(n_3463), .C(n_30694), .D(n_2850), .Z(n_3465
		));
	notech_ao4 i_2300(.A(n_2363), .B(n_2412), .C(n_2065), .D(n_30841), .Z(n_3466
		));
	notech_and4 i_2308(.A(n_3466), .B(n_3154), .C(n_2598), .D(n_4037), .Z(n_3469
		));
	notech_and4 i_2318(.A(n_3469), .B(n_2614), .C(n_1332), .D(n_30678), .Z(n_3472
		));
	notech_and4 i_2312(.A(n_2238), .B(n_4031), .C(n_2239), .D(n_2099), .Z(n_3475
		));
	notech_and4 i_2321(.A(n_4034), .B(n_3475), .C(n_3062), .D(n_3472), .Z(n_3478
		));
	notech_and2 i_631(.A(n_2229), .B(n_3965), .Z(n_3481));
	notech_and4 i_2297(.A(n_2231), .B(n_3279), .C(n_2232), .D(n_2233), .Z(n_3485
		));
	notech_and4 i_2301(.A(n_4028), .B(n_3485), .C(n_223492236), .D(n_4044), 
		.Z(n_3488));
	notech_and4 i_2307(.A(n_3488), .B(n_2394), .C(n_2237), .D(n_4084), .Z(n_3490
		));
	notech_and4 i_2310(.A(n_4007), .B(n_30685), .C(n_1936), .D(n_3490), .Z(n_3491
		));
	notech_and4 i_2317(.A(n_2572), .B(n_30692), .C(n_3481), .D(n_3491), .Z(n_3494
		));
	notech_and4 i_2322(.A(n_4076), .B(n_3494), .C(n_2615), .D(n_3128), .Z(n_3496
		));
	notech_and4 i_2327(.A(n_3496), .B(n_3252), .C(n_2240), .D(n_3478), .Z(n_3498
		));
	notech_and4 i_2331(.A(n_1329), .B(n_2021), .C(n_3498), .D(n_2898), .Z(n_3500
		));
	notech_and2 i_2381(.A(n_2723), .B(n_2946), .Z(n_3507));
	notech_ao4 i_2368(.A(n_58482), .B(n_2250), .C(n_2285), .D(n_2245), .Z(n_3508
		));
	notech_and2 i_21973077(.A(n_4007), .B(n_4047), .Z(n_3510));
	notech_and4 i_2356(.A(n_1193), .B(n_1833), .C(n_3510), .D(n_30681), .Z(n_3513
		));
	notech_and4 i_2359(.A(n_2252), .B(n_3513), .C(n_2253), .D(n_2254), .Z(n_3516
		));
	notech_ao3 i_2361(.A(n_3516), .B(n_2255), .C(n_1807), .Z(n_3518));
	notech_and4 i_2364(.A(n_4058), .B(n_2256), .C(n_2257), .D(n_3518), .Z(n_3521
		));
	notech_and4 i_2367(.A(n_2233), .B(n_1938), .C(n_3521), .D(n_2571), .Z(n_3523
		));
	notech_and4 i_2374(.A(n_2263), .B(n_3523), .C(n_3508), .D(n_2262), .Z(n_3525
		));
	notech_and4 i_2375(.A(n_4017), .B(n_4019), .C(n_4022), .D(n_2264), .Z(n_3528
		));
	notech_and4 i_2379(.A(n_2206), .B(n_733), .C(n_2265), .D(n_3528), .Z(n_3530
		));
	notech_and4 i_2384(.A(n_3525), .B(n_3530), .C(n_3507), .D(n_2266), .Z(n_3532
		));
	notech_ao4 i_2366(.A(n_30785), .B(n_30776), .C(n_2285), .D(n_2288), .Z(n_3534
		));
	notech_and4 i_2377(.A(n_3534), .B(n_3261), .C(n_2532), .D(n_3481), .Z(n_3537
		));
	notech_and4 i_2385(.A(n_4046), .B(n_3537), .C(n_3967), .D(n_30720), .Z(n_3540
		));
	notech_and4 i_2390(.A(n_3540), .B(n_3532), .C(n_466), .D(n_2790), .Z(n_3542
		));
	notech_and4 i_2391(.A(n_2304), .B(n_960), .C(n_3542), .D(n_2267), .Z(n_3543
		));
	notech_and3 i_3610(.A(n_223492236), .B(n_1792), .C(n_3355), .Z(n_3545)
		);
	notech_and4 i_2394(.A(n_68), .B(n_901), .C(n_3543), .D(n_3545), .Z(n_3548
		));
	notech_ao3 i_2425(.A(n_894), .B(n_2620), .C(n_30754), .Z(n_3552));
	notech_and4 i_2431(.A(n_2826), .B(n_3452), .C(n_2157), .D(n_3552), .Z(n_3553
		));
	notech_and4 i_2432(.A(n_2884), .B(n_1728), .C(n_2379), .D(n_2850), .Z(n_3556
		));
	notech_and3 i_2433(.A(n_4016), .B(n_2498), .C(n_3972), .Z(n_3558));
	notech_and4 i_2440(.A(n_3556), .B(n_3553), .C(n_3558), .D(n_2937), .Z(n_3560
		));
	notech_and4 i_2416(.A(n_3062), .B(n_2560), .C(n_2610), .D(n_2829), .Z(n_3564
		));
	notech_and4 i_2400(.A(n_3107), .B(n_2614), .C(n_2269), .D(n_30724), .Z(n_3567
		));
	notech_and4 i_2404(.A(n_2516), .B(n_2638), .C(n_3567), .D(n_1985), .Z(n_3570
		));
	notech_and4 i_2407(.A(n_3570), .B(n_2709), .C(n_2631), .D(n_3834), .Z(n_3572
		));
	notech_and4 i_2411(.A(n_4058), .B(n_2049), .C(n_2457), .D(n_3572), .Z(n_3574
		));
	notech_and4 i_2408(.A(n_2678), .B(n_2791), .C(n_730), .D(n_1958), .Z(n_3576
		));
	notech_and4 i_2415(.A(n_3576), .B(n_3779), .C(n_3574), .D(n_2099), .Z(n_3579
		));
	notech_and4 i_2420(.A(n_2555), .B(n_3579), .C(n_3564), .D(n_2557), .Z(n_3581
		));
	notech_and4 i_2423(.A(n_2686), .B(n_2675), .C(n_2526), .D(n_3581), .Z(n_3584
		));
	notech_and4 i_2434(.A(n_2903), .B(n_3584), .C(n_2654), .D(n_2702), .Z(n_3586
		));
	notech_and4 i_2435(.A(n_2572), .B(n_2415), .C(n_2309), .D(n_1969), .Z(n_3588
		));
	notech_and4 i_2441(.A(n_2904), .B(n_3588), .C(n_3586), .D(n_2664), .Z(n_3591
		));
	notech_and4 i_1522(.A(n_2572), .B(n_2906), .C(n_2513), .D(n_2918), .Z(n_2921
		));
	notech_or2 i_104573104(.A(n_3957), .B(n_2401), .Z(n_208149924));
	notech_and2 i_186(.A(n_2689), .B(n_2501), .Z(n_3957));
	notech_ao3 i_117073103(.A(n_30658), .B(n_30655), .C(n_3277), .Z(n_207949923
		));
	notech_nao3 i_23111411(.A(n_58592), .B(n_2397), .C(n_2282), .Z(n_1984)
		);
	notech_or4 i_860(.A(n_2282), .B(n_2407), .C(n_58514), .D(n_30841), .Z(n_4079
		));
	notech_and2 i_5673091(.A(n_30696), .B(n_30856), .Z(n_1960));
	notech_and4 i_63865(.A(n_2688), .B(n_2684), .C(n_2662), .D(n_1996), .Z(n_4024
		));
	notech_nor2 i_14(.A(n_2182), .B(n_2185), .Z(n_3971));
	notech_nao3 i_448(.A(modrm[5]), .B(n_30656), .C(n_2325), .Z(n_4027));
	notech_or4 i_23110640(.A(n_2311), .B(n_58592), .C(n_58482), .D(n_30785),
		 .Z(n_4047));
	notech_or2 i_462(.A(n_3957), .B(n_2355), .Z(n_4007));
	notech_or4 i_23111096(.A(n_2383), .B(n_2486), .C(n_2290), .D(n_2292), .Z
		(n_4055));
	notech_and2 i_28473072(.A(n_4022), .B(n_30721), .Z(n_1114));
	notech_or4 i_409(.A(n_2292), .B(n_58601), .C(n_58592), .D(n_30800), .Z(n_4022
		));
	notech_nor2 i_23111399(.A(n_2299), .B(n_2339), .Z(n_4088));
	notech_nor2 i_67173070(.A(n_2101), .B(n_2485), .Z(n_204849898));
	notech_or4 i_359(.A(n_58497), .B(n_2313), .C(n_2389), .D(n_2303), .Z(n_4046
		));
	notech_ao4 i_45773061(.A(n_2118), .B(n_2363), .C(n_2278), .D(n_2339), .Z
		(n_1193));
	notech_or4 i_23111396(.A(n_2339), .B(n_58592), .C(n_58482), .D(n_2271), 
		.Z(n_4044));
	notech_or4 i_8(.A(n_2360), .B(n_2280), .C(n_2282), .D(n_2363), .Z(n_4056
		));
	notech_and4 i_1518(.A(n_4017), .B(n_2915), .C(n_2628), .D(n_3996), .Z(n_2918
		));
	notech_and3 i_55873057(.A(n_4031), .B(n_4036), .C(n_1637), .Z(n_696));
	notech_ao3 i_188(.A(n_30658), .B(n_30690), .C(n_2297), .Z(n_4050));
	notech_nand2 i_63973050(.A(n_3107), .B(n_2614), .Z(n_1086));
	notech_and2 i_68873045(.A(n_4048), .B(n_2195), .Z(n_1925));
	notech_or4 i_23110877(.A(n_58497), .B(n_30844), .C(n_30806), .D(n_58592)
		, .Z(n_4048));
	notech_or4 i_853(.A(n_2311), .B(n_58601), .C(n_58470), .D(n_30729), .Z(n_2305
		));
	notech_or4 i_23110865(.A(n_2286), .B(n_2383), .C(n_30844), .D(n_30806), 
		.Z(n_3993));
	notech_ao3 i_23110757(.A(n_58482), .B(n_58470), .C(n_2464), .Z(n_3969)
		);
	notech_and3 i_79573034(.A(n_4064), .B(n_2377), .C(n_4040), .Z(n_1263));
	notech_or4 i_23110871(.A(n_58497), .B(n_2428), .C(n_58514), .D(n_58532),
		 .Z(n_4040));
	notech_and3 i_816(.A(n_2707), .B(n_2598), .C(n_2704), .Z(n_4071));
	notech_and2 i_541(.A(n_2516), .B(n_3733), .Z(n_4070));
	notech_or4 i_38(.A(n_2410), .B(n_2372), .C(n_4090), .D(n_30851), .Z(n_3984
		));
	notech_and4 i_1515(.A(n_2912), .B(n_2709), .C(n_3980), .D(n_3931), .Z(n_2915
		));
	notech_and4 i_337(.A(n_2310), .B(n_30660), .C(n_58568), .D(n_30653), .Z(n_3974
		));
	notech_or2 i_685(.A(n_2400), .B(n_4072), .Z(n_4030));
	notech_or4 i_23110610(.A(n_2286), .B(n_2311), .C(n_30785), .D(n_30855), 
		.Z(n_4093));
	notech_and4 i_1511(.A(n_2285), .B(n_4014), .C(n_3838), .D(n_2909), .Z(n_2912
		));
	notech_nand3 i_1279(.A(n_58482), .B(n_58591), .C(n_30690), .Z(n_4064));
	notech_or4 i_1053(.A(n_58581), .B(n_58568), .C(n_58550), .D(n_2355), .Z(n_4076
		));
	notech_or4 i_23110880(.A(n_58581), .B(n_2382), .C(n_58568), .D(n_58550),
		 .Z(n_4002));
	notech_or4 i_670(.A(n_2214), .B(n_2497), .C(n_30849), .D(n_30850), .Z(n_4086
		));
	notech_nor2 i_10(.A(n_3935), .B(n_2577), .Z(n_3978));
	notech_or4 i_23111093(.A(n_2360), .B(n_58497), .C(n_2333), .D(n_30702), 
		.Z(n_4026));
	notech_or4 i_11(.A(n_2360), .B(n_2280), .C(n_2282), .D(n_1818), .Z(n_4031
		));
	notech_nor2 i_19(.A(n_4090), .B(n_30791), .Z(n_3986));
	notech_ao3 i_255(.A(n_30658), .B(n_30793), .C(n_2101), .Z(n_4060));
	notech_and4 i_1508(.A(n_4013), .B(n_2255), .C(n_30707), .D(n_30682), .Z(n_2909
		));
	notech_and4 i_1519(.A(n_2162), .B(n_2623), .C(n_4082), .D(n_2019), .Z(n_2906
		));
	notech_or4 i_447(.A(n_58498), .B(n_2519), .C(n_58514), .D(n_30841), .Z(n_4014
		));
	notech_and2 i_412(.A(n_2206), .B(n_4028), .Z(n_2124));
	notech_and2 i_330(.A(n_2359), .B(n_2355), .Z(n_4072));
	notech_and4 i_155(.A(n_3967), .B(n_2171), .C(n_2479), .D(n_2014), .Z(n_2904
		));
	notech_and2 i_613(.A(n_3965), .B(n_3994), .Z(n_2903));
	notech_nao3 i_466(.A(n_30851), .B(n_30656), .C(n_2325), .Z(n_4036));
	notech_ao3 i_93(.A(n_3895), .B(adz), .C(n_2348), .Z(n_4001));
	notech_nor2 i_843(.A(n_2382), .B(n_30791), .Z(n_4080));
	notech_or4 i_139(.A(n_2360), .B(n_58498), .C(n_30738), .D(n_1802), .Z(n_4017
		));
	notech_and3 i_1429(.A(n_2516), .B(n_1890), .C(n_2264), .Z(n_2900));
	notech_or4 i_660(.A(n_2410), .B(n_2037), .C(n_3954), .D(modrm[5]), .Z(n_4053
		));
	notech_and2 i_272(.A(n_2400), .B(n_30787), .Z(n_3958));
	notech_nao3 i_526(.A(n_2397), .B(n_30659), .C(n_2276), .Z(n_4013));
	notech_and2 i_17(.A(n_4067), .B(n_30713), .Z(n_2151));
	notech_or2 i_248(.A(n_3836), .B(n_3957), .Z(n_3994));
	notech_and2 i_772(.A(n_2557), .B(n_2555), .Z(n_2899));
	notech_and4 i_177(.A(n_4008), .B(n_2894), .C(n_30680), .D(n_2895), .Z(n_2898
		));
	notech_ao4 i_239(.A(n_2410), .B(n_2403), .C(n_2325), .D(n_2282), .Z(n_2398
		));
	notech_ao3 i_243(.A(n_2380), .B(n_1951), .C(n_30781), .Z(n_1942));
	notech_and3 i_654(.A(n_2709), .B(n_2071), .C(n_2587), .Z(n_1856));
	notech_and4 i_304(.A(n_2379), .B(n_2699), .C(n_2483), .D(n_1870), .Z(n_1865
		));
	notech_and3 i_260(.A(n_30724), .B(n_1921), .C(n_30696), .Z(n_1834));
	notech_nor2 i_481(.A(n_4057), .B(n_30757), .Z(n_1950));
	notech_and2 i_4450(.A(n_3803), .B(n_3982), .Z(n_1014));
	notech_and2 i_4611(.A(n_4031), .B(n_4036), .Z(n_853));
	notech_and4 i_166(.A(n_4055), .B(n_2538), .C(n_2663), .D(n_3059), .Z(n_872
		));
	notech_and3 i_268(.A(n_2216), .B(n_4037), .C(n_4038), .Z(n_738));
	notech_ao4 i_744(.A(n_3957), .B(n_2485), .C(n_30785), .D(n_2519), .Z(n_811
		));
	notech_and2 i_1433(.A(n_2014), .B(n_2305), .Z(n_2895));
	notech_and4 i_3961(.A(n_3838), .B(n_3973), .C(n_3987), .D(n_4029), .Z(n_2894
		));
	notech_and4 i_162(.A(n_3665), .B(n_1915), .C(n_2212), .D(n_1728), .Z(n_2893
		));
	notech_ao3 i_23111288(.A(n_30849), .B(n_30850), .C(n_2113), .Z(n_4091)
		);
	notech_and4 i_384(.A(n_2654), .B(n_2887), .C(n_1951), .D(n_2619), .Z(n_2890
		));
	notech_and2 i_420(.A(n_2384), .B(n_2382), .Z(n_4090));
	notech_ao3 i_136(.A(n_58601), .B(n_58591), .C(n_2464), .Z(n_4089));
	notech_or4 i_15(.A(n_2315), .B(n_2330), .C(n_2214), .D(n_1900), .Z(n_4087
		));
	notech_or4 i_23111405(.A(n_2289), .B(n_2280), .C(n_2338), .D(n_30659), .Z
		(n_4085));
	notech_nand3 i_274(.A(n_2037), .B(n_2287), .C(n_2375), .Z(n_4084));
	notech_or4 i_33(.A(n_2360), .B(n_58497), .C(n_3935), .D(n_30855), .Z(n_4082
		));
	notech_and2 i_238(.A(n_2517), .B(n_2407), .Z(n_3935));
	notech_and4 i_1439(.A(n_2049), .B(n_2500), .C(n_2510), .D(n_30720), .Z(n_2887
		));
	notech_nao3 i_2969(.A(n_58581), .B(n_2272), .C(n_2403), .Z(n_3733));
	notech_or4 i_1256(.A(n_2282), .B(n_2300), .C(n_30844), .D(n_30806), .Z(n_4067
		));
	notech_or4 i_1265(.A(n_2346), .B(n_2302), .C(n_30851), .D(n_2374), .Z(n_4066
		));
	notech_and2 i_331(.A(n_3277), .B(n_2318), .Z(n_4065));
	notech_or4 i_1294(.A(n_2286), .B(n_2311), .C(n_30785), .D(adz), .Z(n_4062
		));
	notech_or2 i_1295(.A(n_2410), .B(n_2403), .Z(n_4061));
	notech_nor2 i_586(.A(n_3836), .B(n_2101), .Z(n_4059));
	notech_and2 i_207(.A(n_2497), .B(n_2359), .Z(n_3836));
	notech_or4 i_62(.A(n_2276), .B(n_1902), .C(n_2316), .D(n_2289), .Z(n_4058
		));
	notech_ao3 i_23110703(.A(n_58581), .B(n_2272), .C(n_2330), .Z(n_4057));
	notech_ao3 i_201(.A(n_30658), .B(n_30690), .C(n_2275), .Z(n_4054));
	notech_and3 i_355(.A(n_3777), .B(n_4046), .C(n_4034), .Z(n_2884));
	notech_and2 i_332(.A(n_2485), .B(n_2401), .Z(n_3954));
	notech_ao3 i_848(.A(n_30659), .B(n_2296), .C(n_2393), .Z(n_4052));
	notech_or4 i_235(.A(n_2289), .B(n_2338), .C(n_2271), .D(n_2280), .Z(n_4051
		));
	notech_and2 i_487(.A(n_3777), .B(n_4046), .Z(n_2883));
	notech_or2 i_368(.A(n_2285), .B(n_2128), .Z(n_4049));
	notech_ao3 i_23110868(.A(n_58550), .B(n_2324), .C(n_2368), .Z(n_4045));
	notech_or2 i_859(.A(n_2278), .B(n_2337), .Z(n_4043));
	notech_or4 i_669(.A(n_2360), .B(n_58497), .C(n_2486), .D(n_30702), .Z(n_4041
		));
	notech_or2 i_1025(.A(n_2285), .B(n_2095), .Z(n_4038));
	notech_or2 i_35(.A(n_1819), .B(n_2285), .Z(n_4037));
	notech_nor2 i_216(.A(n_2485), .B(n_2215), .Z(n_4035));
	notech_or4 i_25(.A(n_58497), .B(n_2313), .C(n_2389), .D(n_2291), .Z(n_4034
		));
	notech_ao3 i_31(.A(n_30658), .B(n_2349), .C(n_2297), .Z(n_4033));
	notech_or4 i_36(.A(n_2348), .B(n_2360), .C(n_2282), .D(n_1812), .Z(n_4032
		));
	notech_or4 i_23110664(.A(n_2292), .B(n_58601), .C(n_58591), .D(n_30703),
		 .Z(n_4029));
	notech_nand3 i_212(.A(n_30659), .B(n_2530), .C(n_30841), .Z(n_4028));
	notech_or4 i_123(.A(n_2469), .B(n_30794), .C(n_30855), .D(n_30779), .Z(n_4025
		));
	notech_ao3 i_680(.A(modrm[2]), .B(n_2271), .C(n_2564), .Z(n_4023));
	notech_or4 i_1109(.A(n_2347), .B(n_2289), .C(n_3963), .D(n_30845), .Z(n_4020
		));
	notech_and2 i_343(.A(n_30785), .B(n_30729), .Z(n_3963));
	notech_or4 i_23111423(.A(n_2289), .B(n_30738), .C(n_2284), .D(n_2271), .Z
		(n_4019));
	notech_and4 i_23011455(.A(emul), .B(fpu), .C(n_30853), .D(n_2469), .Z(n_4018
		));
	notech_nao3 i_318(.A(n_30658), .B(n_30662), .C(n_2101), .Z(n_4016));
	notech_nor2 i_388(.A(n_3958), .B(n_4072), .Z(n_4015));
	notech_and4 i_1404(.A(n_2834), .B(n_2880), .C(n_2009), .D(n_2010), .Z(n_2881
		));
	notech_and4 i_1403(.A(n_1920), .B(n_2847), .C(n_1870), .D(n_30747), .Z(n_2880
		));
	notech_and4 i_27(.A(emul), .B(fpu), .C(n_30853), .D(n_30657), .Z(n_4011)
		);
	notech_and3 i_23011467(.A(cpl[1]), .B(cpl[0]), .C(ipg_fault), .Z(n_4010)
		);
	notech_and2 i_20(.A(n_30657), .B(ipg_fault), .Z(n_4009));
	notech_or4 i_1117(.A(n_2410), .B(n_2037), .C(n_30851), .D(n_2401), .Z(n_4008
		));
	notech_ao3 i_249(.A(n_58581), .B(n_2272), .C(n_2381), .Z(n_4006));
	notech_nand3 i_133(.A(n_3895), .B(n_58550), .C(n_2324), .Z(n_4005));
	notech_nand2 i_407(.A(n_2330), .B(n_2381), .Z(n_3895));
	notech_or4 i_464(.A(n_58497), .B(n_2519), .C(n_58514), .D(n_58532), .Z(n_4004
		));
	notech_nor2 i_141(.A(n_2244), .B(n_2523), .Z(n_4003));
	notech_and2 i_411(.A(n_2485), .B(n_2497), .Z(n_3845));
	notech_or4 i_217(.A(n_2403), .B(n_2316), .C(n_2311), .D(n_2290), .Z(n_3998
		));
	notech_nao3 i_668(.A(n_30660), .B(adz), .C(n_2519), .Z(n_3996));
	notech_or4 i_1399(.A(n_30809), .B(n_30759), .C(n_2875), .D(n_30763), .Z(n_2878
		));
	notech_or4 i_23111108(.A(n_2289), .B(n_2325), .C(n_2271), .D(n_30785), .Z
		(n_3992));
	notech_or4 i_229(.A(n_2348), .B(n_2360), .C(n_2282), .D(n_2331), .Z(n_3991
		));
	notech_nor2 i_538(.A(n_2278), .B(n_2393), .Z(n_3990));
	notech_or4 i_231(.A(n_58497), .B(n_2316), .C(n_2389), .D(n_2291), .Z(n_3987
		));
	notech_ao3 i_23111162(.A(n_58470), .B(n_58601), .C(n_2318), .Z(n_3985)
		);
	notech_nao3 i_285(.A(n_30658), .B(n_30790), .C(n_2101), .Z(n_3982));
	notech_or4 i_42(.A(n_2311), .B(n_3963), .C(n_58481), .D(n_58470), .Z(n_3981
		));
	notech_or4 i_16(.A(n_58497), .B(n_3935), .C(n_2283), .D(n_30855), .Z(n_3980
		));
	notech_or4 i_125(.A(n_2360), .B(n_58497), .C(n_3935), .D(adz), .Z(n_3979
		));
	notech_or4 i_370(.A(n_2290), .B(n_2292), .C(n_2383), .D(n_2333), .Z(n_3977
		));
	notech_or4 i_498(.A(n_2360), .B(n_58497), .C(n_2325), .D(n_2299), .Z(n_3975
		));
	notech_nao3 i_2992(.A(modrm[2]), .B(n_2530), .C(n_30659), .Z(n_3973));
	notech_or4 i_51(.A(n_2410), .B(n_2373), .C(n_4090), .D(n_30851), .Z(n_3972
		));
	notech_or4 i_23110592(.A(n_2360), .B(n_58497), .C(n_2289), .D(n_2410), .Z
		(n_3970));
	notech_ao3 i_23110727(.A(n_58581), .B(n_2272), .C(n_2368), .Z(n_3968));
	notech_or4 i_338(.A(n_58497), .B(n_2316), .C(n_30738), .D(n_2303), .Z(n_3967
		));
	notech_or4 i_128(.A(n_30738), .B(n_58481), .C(n_58470), .D(n_30729), .Z(n_3965
		));
	notech_or4 i_23110595(.A(n_58498), .B(n_2621), .C(n_58532), .D(n_30842),
		 .Z(n_3964));
	notech_and2 i_147(.A(n_3867), .B(n_1875), .Z(n_2380));
	notech_or4 i_1297(.A(n_58481), .B(n_58470), .C(adz), .D(n_30794), .Z(n_3867
		));
	notech_and2 i_3098(.A(n_4062), .B(n_4093), .Z(n_2366));
	notech_ao3 i_30(.A(n_30842), .B(n_30841), .C(n_58498), .Z(n_2354));
	notech_ao3 i_37(.A(n_30842), .B(n_58532), .C(n_58498), .Z(n_2369));
	notech_nand2 i_3157(.A(n_2327), .B(n_30692), .Z(n_2307));
	notech_or4 i_1392(.A(n_30775), .B(n_30805), .C(n_2873), .D(n_30749), .Z(n_2875
		));
	notech_and2 i_415(.A(n_2286), .B(n_2290), .Z(n_3961));
	notech_ao3 i_256(.A(n_2385), .B(n_30851), .C(n_2410), .Z(n_3959));
	notech_ao3 i_89(.A(n_30849), .B(modrm[4]), .C(n_2214), .Z(n_2210));
	notech_or4 i_3282(.A(n_2386), .B(n_58601), .C(n_58470), .D(n_30844), .Z(n_2182
		));
	notech_or4 i_3297(.A(n_2386), .B(n_58481), .C(n_58470), .D(n_30844), .Z(n_2167
		));
	notech_nand2 i_3299(.A(n_30726), .B(n_30691), .Z(n_2165));
	notech_nand3 i_1388(.A(n_2538), .B(n_2111), .C(n_2872), .Z(n_2873));
	notech_or4 i_110(.A(n_2280), .B(n_2282), .C(n_58532), .D(n_30842), .Z(n_2118
		));
	notech_or4 i_3446(.A(n_58481), .B(n_58470), .C(n_2271), .D(n_30807), .Z(n_2018
		));
	notech_and4 i_1384(.A(n_1815), .B(n_4005), .C(n_2870), .D(n_2789), .Z(n_2872
		));
	notech_nor2 i_23111378(.A(n_2564), .B(n_2271), .Z(n_1987));
	notech_and2 i_12(.A(n_4025), .B(n_30723), .Z(n_1953));
	notech_and4 i_23110715(.A(adz), .B(n_2296), .C(n_2469), .D(n_2466), .Z(n_3950
		));
	notech_and4 i_1381(.A(n_2171), .B(n_2867), .C(n_2857), .D(n_2022), .Z(n_2870
		));
	notech_and3 i_3727(.A(n_3996), .B(n_2579), .C(n_4082), .Z(n_1737));
	notech_and4 i_1377(.A(n_1656), .B(n_2627), .C(n_2863), .D(n_1623), .Z(n_2867
		));
	notech_nand3 i_699(.A(n_4031), .B(n_4056), .C(n_2611), .Z(n_3956));
	notech_and2 i_3849(.A(n_3838), .B(n_4028), .Z(n_1615));
	notech_nand3 i_198(.A(n_30659), .B(n_30841), .C(n_2536), .Z(n_3838));
	notech_and4 i_3919(.A(n_2579), .B(n_1970), .C(n_3998), .D(n_30724), .Z(n_1545
		));
	notech_and2 i_72(.A(n_2063), .B(n_2969), .Z(n_3955));
	notech_or4 i_861(.A(n_58498), .B(n_2865), .C(n_58532), .D(n_30842), .Z(n_3803
		));
	notech_and2 i_4744(.A(n_3739), .B(n_2195), .Z(n_720));
	notech_or4 i_467(.A(n_58577), .B(n_58568), .C(n_58550), .D(n_2401), .Z(n_3739
		));
	notech_or2 i_273(.A(n_1858), .B(n_3963), .Z(n_3880));
	notech_and3 i_5210(.A(n_1829), .B(n_1828), .C(n_4084), .Z(n_254));
	notech_nand3 i_4(.A(n_58577), .B(n_58568), .C(n_58550), .Z(n_2410));
	notech_or4 i_1350(.A(n_2347), .B(n_2244), .C(n_30845), .D(adz), .Z(n_2865
		));
	notech_nand3 i_60(.A(n_58482), .B(n_58591), .C(n_30659), .Z(n_2302));
	notech_nand3 i_65(.A(n_58601), .B(n_58591), .C(n_30659), .Z(n_2275));
	notech_nao3 i_23(.A(n_30841), .B(n_58514), .C(n_58498), .Z(n_2383));
	notech_or4 i_18(.A(n_2372), .B(n_2214), .C(n_2330), .D(n_2504), .Z(n_3931
		));
	notech_and2 i_21(.A(n_30856), .B(n_1919), .Z(n_1951));
	notech_and2 i_22(.A(n_223492236), .B(n_1792), .Z(n_2017));
	notech_and3 i_24(.A(n_58581), .B(n_30845), .C(n_30844), .Z(n_2397));
	notech_nand3 i_61(.A(n_58470), .B(n_58601), .C(n_30659), .Z(n_2278));
	notech_and3 i_76(.A(n_58482), .B(n_58470), .C(n_30659), .Z(n_3908));
	notech_ao4 i_26(.A(n_2278), .B(n_2458), .C(n_2455), .D(n_30702), .Z(n_2123
		));
	notech_and2 i_29(.A(n_2141), .B(n_4013), .Z(n_2065));
	notech_nand2 i_74(.A(opz[1]), .B(n_2322), .Z(n_2320));
	notech_and2 i_34(.A(n_4031), .B(n_4056), .Z(n_2116));
	notech_and4 i_1374(.A(n_3964), .B(n_4004), .C(n_2860), .D(n_2676), .Z(n_2863
		));
	notech_and2 i_53(.A(n_2192), .B(n_4017), .Z(n_2176));
	notech_and2 i_57(.A(n_2071), .B(n_1835), .Z(n_2171));
	notech_and3 i_58(.A(n_2233), .B(n_1938), .C(n_4079), .Z(n_2049));
	notech_and3 i_80(.A(n_2629), .B(n_30709), .C(n_30707), .Z(n_2357));
	notech_and4 i_1371(.A(n_2435), .B(n_3998), .C(n_2008), .D(n_2630), .Z(n_2860
		));
	notech_nand3 i_97(.A(n_2062), .B(adz), .C(n_30660), .Z(n_3890));
	notech_nand3 i_122(.A(n_30726), .B(n_30691), .C(n_30725), .Z(n_2164));
	notech_or4 i_167(.A(n_58498), .B(n_2316), .C(n_30738), .D(n_2291), .Z(n_3876
		));
	notech_ao4 i_130(.A(n_2278), .B(n_2346), .C(n_2275), .D(n_2393), .Z(n_1958
		));
	notech_or4 i_131(.A(fpu), .B(twobyte), .C(ipg_fault), .D(op[7]), .Z(n_2403
		));
	notech_and4 i_135(.A(n_2623), .B(n_3964), .C(n_3965), .D(n_2380), .Z(n_2332
		));
	notech_and3 i_146(.A(n_2327), .B(n_30692), .C(n_2305), .Z(n_2304));
	notech_and2 i_160(.A(n_1918), .B(n_1794), .Z(n_1978));
	notech_ao3 i_704(.A(n_4014), .B(n_1921), .C(n_30661), .Z(n_2857));
	notech_and4 i_170(.A(n_3876), .B(n_2609), .C(n_2663), .D(n_2500), .Z(n_901
		));
	notech_and4 i_175(.A(n_1874), .B(n_2702), .C(n_2900), .D(n_30665), .Z(n_1504
		));
	notech_nand2 i_182(.A(n_30850), .B(modrm[3]), .Z(n_2315));
	notech_and4 i_191(.A(n_58581), .B(n_30845), .C(n_58550), .D(n_2369), .Z(n_3846
		));
	notech_and2 i_204(.A(n_3994), .B(n_30694), .Z(n_1999));
	notech_ao4 i_208(.A(n_2290), .B(n_2447), .C(n_30729), .D(n_2448), .Z(n_2327
		));
	notech_and2 i_211(.A(n_2308), .B(n_2294), .Z(n_2058));
	notech_or4 i_469(.A(n_2410), .B(n_2315), .C(n_2382), .D(n_30851), .Z(n_3834
		));
	notech_and2 i_214(.A(n_3996), .B(n_4082), .Z(n_1972));
	notech_and3 i_220(.A(n_4002), .B(n_1797), .C(n_4017), .Z(n_1777));
	notech_and4 i_309(.A(n_2638), .B(n_2014), .C(n_2192), .D(n_30678), .Z(n_2854
		));
	notech_ao4 i_225(.A(n_1879), .B(n_2488), .C(n_2037), .D(n_2489), .Z(n_2024
		));
	notech_and2 i_240(.A(n_4014), .B(n_2005), .Z(n_1624));
	notech_and2 i_241(.A(n_2057), .B(n_1794), .Z(n_1290));
	notech_nor2 i_862(.A(n_2400), .B(n_2098), .Z(n_3820));
	notech_and2 i_252(.A(n_1985), .B(n_30711), .Z(n_1678));
	notech_and4 i_364(.A(n_2394), .B(n_1958), .C(n_2065), .D(n_2285), .Z(n_2852
		));
	notech_and4 i_261(.A(n_2094), .B(n_4026), .C(n_2155), .D(n_1825), .Z(n_497
		));
	notech_and4 i_263(.A(n_2394), .B(n_1958), .C(n_2026), .D(n_2925), .Z(n_1434
		));
	notech_and4 i_265(.A(n_2179), .B(n_3312), .C(n_3179), .D(n_2180), .Z(n_493
		));
	notech_and4 i_267(.A(n_2398), .B(n_1545), .C(n_30706), .D(n_30685), .Z(n_68
		));
	notech_and4 i_270(.A(n_2639), .B(n_3184), .C(n_3179), .D(n_2937), .Z(n_537
		));
	notech_and2 i_271(.A(n_30689), .B(n_30688), .Z(n_2099));
	notech_ao4 i_278(.A(n_2244), .B(n_2523), .C(n_30787), .D(n_2485), .Z(n_2212
		));
	notech_and2 i_279(.A(n_4041), .B(n_1896), .Z(n_2094));
	notech_and3 i_280(.A(n_1993), .B(n_2665), .C(n_2688), .Z(n_1718));
	notech_and3 i_289(.A(n_2046), .B(n_1912), .C(n_1914), .Z(n_1993));
	notech_and2 i_295(.A(n_2136), .B(n_2978), .Z(n_1329));
	notech_and2 i_299(.A(n_3803), .B(n_30722), .Z(n_1623));
	notech_and4 i_477(.A(n_2151), .B(n_2166), .C(n_2588), .D(n_1890), .Z(n_2850
		));
	notech_and4 i_305(.A(n_2678), .B(n_2791), .C(n_1857), .D(n_533), .Z(n_530
		));
	notech_and4 i_1396(.A(n_2707), .B(n_2352), .C(n_2839), .D(n_2844), .Z(n_2847
		));
	notech_and2 i_314(.A(n_3977), .B(n_4086), .Z(n_1332));
	notech_and4 i_323(.A(n_208149924), .B(n_4049), .C(n_30689), .D(n_3981), 
		.Z(n_444));
	notech_and3 i_324(.A(n_2663), .B(n_2183), .C(n_3422), .Z(n_204));
	notech_and2 i_333(.A(n_4032), .B(n_2365), .Z(n_1905));
	notech_ao4 i_341(.A(n_2400), .B(n_3845), .C(n_3958), .D(n_2401), .Z(n_2157
		));
	notech_and4 i_357(.A(n_3996), .B(n_4014), .C(n_4082), .D(n_3980), .Z(n_1970
		));
	notech_or4 i_360(.A(n_58498), .B(n_2316), .C(n_2389), .D(n_2303), .Z(n_3779
		));
	notech_or4 i_406(.A(n_2389), .B(n_2290), .C(n_2292), .D(n_30729), .Z(n_3777
		));
	notech_and4 i_1391(.A(n_2465), .B(n_2198), .C(n_2842), .D(n_2831), .Z(n_2844
		));
	notech_or4 i_367(.A(n_3956), .B(n_30778), .C(n_30746), .D(n_30772), .Z(n_3773
		));
	notech_and3 i_371(.A(n_2157), .B(n_1930), .C(n_2625), .Z(n_1870));
	notech_and4 i_1386(.A(n_4084), .B(n_2377), .C(n_2827), .D(n_1712), .Z(n_2842
		));
	notech_and3 i_379(.A(n_2231), .B(n_1833), .C(n_1936), .Z(n_1780));
	notech_and4 i_381(.A(n_3739), .B(n_2195), .C(n_2264), .D(n_719), .Z(n_717
		));
	notech_mux2 i_391(.S(n_58532), .A(modrm[0]), .B(modrm[3]), .Z(n_3763));
	notech_nor2 i_395(.A(n_2301), .B(n_3908), .Z(n_3761));
	notech_mux2 i_397(.S(n_58532), .A(n_30849), .B(n_30847), .Z(n_3760));
	notech_nao3 i_401(.A(n_58550), .B(n_30851), .C(n_2386), .Z(n_2214));
	notech_and3 i_402(.A(n_223492236), .B(n_1792), .C(n_30699), .Z(n_2015)
		);
	notech_and2 i_413(.A(n_3838), .B(n_3973), .Z(n_2076));
	notech_and3 i_421(.A(n_4062), .B(n_4093), .C(n_30695), .Z(n_2022));
	notech_nao3 i_852(.A(n_2385), .B(n_30790), .C(n_2214), .Z(n_3751));
	notech_and2 i_425(.A(n_3751), .B(n_30723), .Z(n_1526));
	notech_and2 i_428(.A(n_4055), .B(n_1857), .Z(n_2029));
	notech_and2 i_437(.A(n_30714), .B(n_30694), .Z(n_1728));
	notech_ao4 i_440(.A(n_2501), .B(n_2382), .C(n_58498), .D(n_2646), .Z(n_733
		));
	notech_and4 i_310(.A(n_4002), .B(n_2195), .C(n_2414), .D(n_2597), .Z(n_2839
		));
	notech_and2 i_454(.A(n_2073), .B(n_2202), .Z(n_2162));
	notech_and4 i_455(.A(n_3979), .B(n_1970), .C(n_30722), .D(n_1978), .Z(n_1969
		));
	notech_and2 i_474(.A(n_3979), .B(n_3980), .Z(n_1816));
	notech_or4 i_835(.A(n_2214), .B(n_2384), .C(modrm[3]), .D(n_30850), .Z(n_3736
		));
	notech_and2 i_476(.A(n_2587), .B(n_1851), .Z(n_1603));
	notech_nand2 i_479(.A(n_3998), .B(n_30724), .Z(n_1967));
	notech_and4 i_492(.A(n_3967), .B(n_3987), .C(n_1796), .D(n_4029), .Z(n_3728
		));
	notech_or4 i_493(.A(n_58498), .B(n_2286), .C(n_58514), .D(n_30841), .Z(n_2368
		));
	notech_and3 i_501(.A(n_30706), .B(n_30685), .C(n_2305), .Z(n_1924));
	notech_and2 i_508(.A(n_2327), .B(n_4047), .Z(n_1923));
	notech_and4 i_515(.A(n_30712), .B(n_1958), .C(n_2377), .D(n_30693), .Z(n_960
		));
	notech_nao3 i_532(.A(n_30659), .B(n_2375), .C(n_2286), .Z(n_2113));
	notech_and2 i_792(.A(n_2411), .B(n_1603), .Z(n_2834));
	notech_or4 i_536(.A(n_58581), .B(n_2338), .C(n_58550), .D(n_30845), .Z(n_2234
		));
	notech_and2 i_545(.A(n_2216), .B(n_30792), .Z(n_1656));
	notech_and2 i_550(.A(n_2132), .B(n_2789), .Z(n_455));
	notech_and4 i_555(.A(n_4027), .B(n_4036), .C(n_4076), .D(n_2091), .Z(n_894
		));
	notech_and4 i_562(.A(n_2233), .B(n_1938), .C(n_4079), .D(n_4058), .Z(n_2047
		));
	notech_and3 i_567(.A(n_3838), .B(n_3973), .C(n_1798), .Z(n_3697));
	notech_and3 i_692(.A(n_4025), .B(n_30723), .C(n_2357), .Z(n_2831));
	notech_and2 i_606(.A(n_2380), .B(n_30856), .Z(n_1593));
	notech_and3 i_94(.A(n_3992), .B(n_1895), .C(n_1831), .Z(n_2829));
	notech_ao4 i_604(.A(n_2387), .B(n_30789), .C(n_2382), .D(n_30791), .Z(n_2827
		));
	notech_ao4 i_618(.A(n_30785), .B(n_2407), .C(n_2485), .D(n_30787), .Z(n_1306
		));
	notech_and2 i_625(.A(n_3982), .B(n_30692), .Z(n_1537));
	notech_and3 i_634(.A(n_3993), .B(n_4040), .C(n_2103), .Z(n_730));
	notech_and3 i_637(.A(n_3992), .B(n_2123), .C(n_30680), .Z(n_1712));
	notech_and4 i_780(.A(n_1949), .B(n_1796), .C(n_3880), .D(n_30665), .Z(n_2826
		));
	notech_or2 i_658(.A(n_3958), .B(n_2355), .Z(n_3672));
	notech_or4 i_659(.A(n_2316), .B(n_2276), .C(n_2373), .D(n_2333), .Z(n_2052
		));
	notech_or2 i_684(.A(n_2400), .B(n_2359), .Z(n_3665));
	notech_ao4 i_708(.A(n_2400), .B(n_3845), .C(n_30794), .D(n_2286), .Z(n_1543
		));
	notech_or4 i_729(.A(n_4010), .B(n_4018), .C(n_3950), .D(n_4015), .Z(n_1262
		));
	notech_and2 i_736(.A(n_3979), .B(n_4032), .Z(n_861));
	notech_and2 i_748(.A(n_2246), .B(n_1984), .Z(n_520));
	notech_and2 i_750(.A(n_2665), .B(n_2394), .Z(n_719));
	notech_and3 i_751(.A(n_2790), .B(n_1993), .C(n_3105), .Z(n_703));
	notech_ao4 i_753(.A(n_2291), .B(n_30800), .C(n_2118), .D(n_2363), .Z(n_673
		));
	notech_and2 i_755(.A(n_4002), .B(n_4048), .Z(n_2080));
	notech_ao4 i_757(.A(n_2422), .B(n_2384), .C(n_2499), .D(n_2382), .Z(n_574
		));
	notech_and2 i_768(.A(n_1936), .B(n_30685), .Z(n_215));
	notech_and3 i_769(.A(n_4041), .B(n_4036), .C(n_2056), .Z(n_1284));
	notech_and3 i_779(.A(n_3880), .B(n_3374), .C(n_2213), .Z(n_218));
	notech_and2 i_781(.A(n_2206), .B(n_733), .Z(n_709));
	notech_and3 i_782(.A(n_2625), .B(n_3779), .C(n_2073), .Z(n_533));
	notech_and3 i_791(.A(n_3979), .B(n_3980), .C(n_4082), .Z(n_1815));
	notech_or4 i_1318(.A(n_30813), .B(n_2817), .C(n_1998), .D(n_2000), .Z(n_2820
		));
	notech_and3 i_804(.A(n_4055), .B(n_2538), .C(n_3834), .Z(n_1340));
	notech_and3 i_810(.A(n_2166), .B(n_2108), .C(n_2380), .Z(n_466));
	notech_and3 i_812(.A(n_1886), .B(n_2686), .C(n_1887), .Z(n_2246));
	notech_and4 i_813(.A(n_3834), .B(n_2036), .C(n_1924), .D(n_3984), .Z(n_1920
		));
	notech_and3 i_818(.A(n_2025), .B(n_2103), .C(n_4027), .Z(n_1346));
	notech_and4 i_2932(.A(n_4047), .B(n_2091), .C(n_1999), .D(n_30714), .Z(n_1996
		));
	notech_or4 i_1315(.A(n_30754), .B(n_30771), .C(n_30808), .D(n_2814), .Z(n_2817
		));
	notech_nao3 i_1313(.A(n_1678), .B(n_2588), .C(n_2812), .Z(n_2814));
	notech_or4 i_1311(.A(n_1997), .B(n_30783), .C(n_2809), .D(n_2078), .Z(n_2812
		));
	notech_nao3 i_1308(.A(n_3777), .B(n_2808), .C(n_222394222), .Z(n_2809)
		);
	notech_and4 i_1307(.A(n_3665), .B(n_1923), .C(n_2804), .D(n_30719), .Z(n_2808
		));
	notech_and4 i_1304(.A(n_2627), .B(n_1995), .C(n_3965), .D(n_2801), .Z(n_2804
		));
	notech_ao3 i_1300(.A(n_2799), .B(n_2216), .C(n_1933), .Z(n_2801));
	notech_and4 i_1298(.A(n_2516), .B(n_2797), .C(n_3998), .D(n_2794), .Z(n_2799
		));
	notech_and4 i_1292(.A(n_30709), .B(n_30707), .C(n_1990), .D(n_1994), .Z(n_2797
		));
	notech_ao4 i_1290(.A(n_58482), .B(n_2734), .C(n_2140), .D(n_58470), .Z(n_2794
		));
	notech_and2 i_237(.A(n_2791), .B(n_2790), .Z(n_2792));
	notech_ao4 i_486(.A(n_2384), .B(n_30787), .C(n_2403), .D(n_30738), .Z(n_2791
		));
	notech_and2 i_43(.A(n_2789), .B(n_1982), .Z(n_2790));
	notech_and3 i_349(.A(n_1901), .B(n_4087), .C(n_3931), .Z(n_2789));
	notech_or4 i_1262(.A(n_222994228), .B(n_1975), .C(n_1976), .D(n_2782), .Z
		(n_2785));
	notech_nand3 i_1259(.A(n_2780), .B(n_2729), .C(n_222794226), .Z(n_2782)
		);
	notech_and4 i_1257(.A(n_2778), .B(n_2212), .C(n_30680), .D(n_2532), .Z(n_2780
		));
	notech_and4 i_1254(.A(n_2765), .B(n_1978), .C(n_2136), .D(n_2777), .Z(n_2778
		));
	notech_and4 i_1253(.A(n_2192), .B(n_2775), .C(n_2744), .D(n_2305), .Z(n_2777
		));
	notech_and4 i_1248(.A(n_1877), .B(n_2772), .C(n_3996), .D(n_30691), .Z(n_2775
		));
	notech_and4 i_1245(.A(n_2768), .B(n_3993), .C(n_2771), .D(n_30724), .Z(n_2772
		));
	notech_ao4 i_1244(.A(n_2458), .B(n_2299), .C(n_2383), .D(n_2621), .Z(n_2771
		));
	notech_ao4 i_1240(.A(n_2734), .B(n_30841), .C(n_2140), .D(n_30844), .Z(n_2768
		));
	notech_and3 i_173(.A(n_2216), .B(n_2733), .C(n_2730), .Z(n_2765));
	notech_and4 i_3740(.A(n_223492236), .B(n_1792), .C(n_2151), .D(n_30699),
		 .Z(n_2760));
	notech_and4 i_226(.A(n_30714), .B(n_30694), .C(n_2091), .D(n_3994), .Z(n_2759
		));
	notech_and2 i_478(.A(n_1993), .B(n_2665), .Z(n_2757));
	notech_and4 i_1213(.A(n_2751), .B(n_222794226), .C(n_2729), .D(n_1955), 
		.Z(n_2754));
	notech_and4 i_1210(.A(n_30797), .B(n_2749), .C(n_30724), .D(n_1954), .Z(n_2751
		));
	notech_and4 i_1208(.A(n_1930), .B(n_2741), .C(n_2747), .D(n_1737), .Z(n_2749
		));
	notech_and4 i_1206(.A(n_1949), .B(n_2744), .C(n_1952), .D(n_2743), .Z(n_2747
		));
	notech_and2 i_251(.A(n_1932), .B(n_30755), .Z(n_2744));
	notech_and2 i_138(.A(n_2192), .B(n_2305), .Z(n_2743));
	notech_and4 i_1203(.A(n_2730), .B(n_2731), .C(n_3965), .D(n_2739), .Z(n_2741
		));
	notech_and4 i_1200(.A(n_3993), .B(n_3992), .C(n_2736), .D(n_3980), .Z(n_2739
		));
	notech_and3 i_1194(.A(n_2733), .B(n_2234), .C(n_1947), .Z(n_2736));
	notech_ao4 i_218(.A(n_2403), .B(n_2389), .C(n_58498), .D(n_2646), .Z(n_2734
		));
	notech_ao4 i_543(.A(n_30729), .B(n_2446), .C(n_2325), .D(n_2282), .Z(n_2733
		));
	notech_ao4 i_1196(.A(n_2166), .B(n_30824), .C(n_2290), .D(n_2464), .Z(n_2731
		));
	notech_ao4 i_696(.A(n_2318), .B(n_2286), .C(n_30729), .D(n_2519), .Z(n_2730
		));
	notech_and4 i_157(.A(n_4084), .B(n_2377), .C(n_3751), .D(n_2727), .Z(n_2729
		));
	notech_ao4 i_1154(.A(n_2118), .B(n_2027), .C(n_2362), .D(n_2331), .Z(n_2727
		));
	notech_and4 i_1173(.A(n_30712), .B(n_1780), .C(n_2395), .D(n_2414), .Z(n_2726
		));
	notech_and2 i_485(.A(n_4002), .B(n_1797), .Z(n_2723));
	notech_and3 i_300(.A(n_3967), .B(n_2171), .C(n_2479), .Z(n_2722));
	notech_and4 i_1182(.A(n_2141), .B(n_4013), .C(n_2015), .D(n_1941), .Z(n_2719
		));
	notech_and4 i_348(.A(n_2195), .B(n_2714), .C(n_2611), .D(n_2713), .Z(n_2717
		));
	notech_ao4 i_1177(.A(n_2384), .B(n_1937), .C(n_2052), .D(n_2331), .Z(n_2714
		));
	notech_and2 i_701(.A(n_4016), .B(n_3972), .Z(n_2713));
	notech_and2 i_452(.A(n_1798), .B(n_2111), .Z(n_2709));
	notech_and4 i_387(.A(n_2190), .B(n_3973), .C(n_2463), .D(n_2675), .Z(n_2707
		));
	notech_and2 i_646(.A(n_2703), .B(n_2543), .Z(n_2704));
	notech_and4 i_473(.A(n_1873), .B(n_2555), .C(n_1874), .D(n_2702), .Z(n_2703
		));
	notech_and2 i_233(.A(n_1800), .B(n_2563), .Z(n_2702));
	notech_and4 i_1127(.A(n_2417), .B(n_2695), .C(n_2198), .D(n_2696), .Z(n_2699
		));
	notech_and4 i_1124(.A(n_2073), .B(n_4067), .C(n_2202), .D(n_30713), .Z(n_2696
		));
	notech_and2 i_399(.A(n_1796), .B(n_4029), .Z(n_2695));
	notech_and2 i_566(.A(n_2157), .B(n_1930), .Z(n_2694));
	notech_and3 i_3466(.A(n_3994), .B(n_30694), .C(n_30714), .Z(n_2690));
	notech_or4 i_101(.A(n_2386), .B(n_2037), .C(n_30844), .D(n_30851), .Z(n_2689
		));
	notech_and2 i_288(.A(n_2246), .B(n_2264), .Z(n_2688));
	notech_ao4 i_376(.A(n_2553), .B(n_2685), .C(n_2557), .D(n_2037), .Z(n_2686
		));
	notech_nand2 i_936(.A(n_1885), .B(modrm[1]), .Z(n_2685));
	notech_and4 i_711(.A(n_2681), .B(n_2675), .C(n_2665), .D(n_2664), .Z(n_2684
		));
	notech_and4 i_1021(.A(n_2179), .B(n_2678), .C(n_2457), .D(n_2022), .Z(n_2681
		));
	notech_and3 i_193(.A(n_2676), .B(n_2189), .C(n_2190), .Z(n_2678));
	notech_and2 i_54(.A(n_2188), .B(n_1907), .Z(n_2676));
	notech_and4 i_358(.A(n_4055), .B(n_1857), .C(n_3977), .D(n_2673), .Z(n_2675
		));
	notech_and4 i_877(.A(n_1855), .B(n_1854), .C(n_2668), .D(n_2238), .Z(n_2673
		));
	notech_ao4 i_137(.A(n_2667), .B(n_2300), .C(n_2666), .D(n_2292), .Z(n_2668
		));
	notech_nand2 i_868(.A(n_2530), .B(n_58532), .Z(n_2667));
	notech_nand2 i_867(.A(n_30841), .B(n_2536), .Z(n_2666));
	notech_and2 i_758(.A(n_2024), .B(n_1911), .Z(n_2665));
	notech_and2 i_614(.A(n_2663), .B(n_2352), .Z(n_2664));
	notech_ao4 i_52(.A(n_2291), .B(n_2052), .C(n_2278), .D(n_2337), .Z(n_2663
		));
	notech_and4 i_1111(.A(n_2484), .B(n_2549), .C(n_2483), .D(n_2661), .Z(n_2662
		));
	notech_and4 i_1108(.A(n_2658), .B(n_2619), .C(n_2607), .D(n_2567), .Z(n_2661
		));
	notech_and4 i_1100(.A(n_2654), .B(n_2157), .C(n_2650), .D(n_2656), .Z(n_2658
		));
	notech_and2 i_602(.A(n_2655), .B(n_4025), .Z(n_2656));
	notech_ao4 i_356(.A(n_2391), .B(n_2303), .C(n_2291), .D(n_30703), .Z(n_2655
		));
	notech_and2 i_293(.A(n_2030), .B(n_3991), .Z(n_2654));
	notech_and4 i_1093(.A(n_2648), .B(n_2643), .C(n_2304), .D(n_2620), .Z(n_2650
		));
	notech_and4 i_383(.A(n_4002), .B(n_4048), .C(n_2076), .D(n_30680), .Z(n_2648
		));
	notech_or4 i_997(.A(n_58581), .B(n_58568), .C(n_30844), .D(n_58591), .Z(n_2646
		));
	notech_and4 i_1087(.A(n_2625), .B(n_2634), .C(n_2332), .D(n_2641), .Z(n_2643
		));
	notech_and4 i_1084(.A(n_4058), .B(n_2049), .C(n_2639), .D(n_3981), .Z(n_2641
		));
	notech_and2 i_242(.A(n_2638), .B(n_2014), .Z(n_2639));
	notech_ao4 i_215(.A(n_2325), .B(n_2384), .C(n_2383), .D(n_2428), .Z(n_2638
		));
	notech_and2 i_616(.A(n_2233), .B(n_1938), .Z(n_2637));
	notech_and4 i_1081(.A(n_2631), .B(n_2628), .C(n_2357), .D(n_30723), .Z(n_2634
		));
	notech_and3 i_302(.A(n_2433), .B(n_2140), .C(n_4064), .Z(n_2631));
	notech_and2 i_569(.A(n_2433), .B(n_2140), .Z(n_2630));
	notech_nor2 i_426(.A(n_4010), .B(n_4018), .Z(n_2629));
	notech_and3 i_774(.A(n_3993), .B(n_4040), .C(n_3733), .Z(n_2628));
	notech_and2 i_410(.A(n_3993), .B(n_4040), .Z(n_2627));
	notech_and2 i_134(.A(n_1877), .B(n_1831), .Z(n_2625));
	notech_and2 i_45(.A(n_30706), .B(n_30685), .Z(n_2623));
	notech_or4 i_923(.A(n_2386), .B(n_30844), .C(n_58601), .D(n_58592), .Z(n_2621
		));
	notech_and2 i_509(.A(n_3987), .B(n_4029), .Z(n_2620));
	notech_and4 i_36692324(.A(n_2611), .B(n_2379), .C(n_2614), .D(n_2616), .Z
		(n_2619));
	notech_and4 i_978(.A(n_4027), .B(n_4036), .C(n_30689), .D(n_30688), .Z(n_2616
		));
	notech_and2 i_783(.A(n_4027), .B(n_4036), .Z(n_2615));
	notech_and3 i_430(.A(n_4041), .B(n_1896), .C(n_4026), .Z(n_2614));
	notech_and4 i_196(.A(n_4044), .B(n_2609), .C(n_2108), .D(n_30721), .Z(n_2611
		));
	notech_and4 i_802(.A(n_4044), .B(n_4051), .C(n_30721), .D(n_4085), .Z(n_2610
		));
	notech_and2 i_458(.A(n_4051), .B(n_4085), .Z(n_2609));
	notech_and4 i_1102(.A(n_2572), .B(n_1969), .C(n_2605), .D(n_2309), .Z(n_2607
		));
	notech_and4 i_63(.A(n_2591), .B(n_2602), .C(n_2588), .D(n_2587), .Z(n_2605
		));
	notech_and4 i_1076(.A(n_3931), .B(n_2598), .C(n_2171), .D(n_2601), .Z(n_2602
		));
	notech_and3 i_1075(.A(n_2192), .B(n_4017), .C(n_2195), .Z(n_2601));
	notech_and3 i_199(.A(n_2103), .B(n_2159), .C(n_1851), .Z(n_2598));
	notech_and2 i_830(.A(n_2103), .B(n_2159), .Z(n_2597));
	notech_or4 i_823(.A(n_58498), .B(n_2486), .C(n_58514), .D(n_30841), .Z(n_2596
		));
	notech_or4 i_863(.A(n_2302), .B(n_58550), .C(n_30806), .D(modrm[5]), .Z(n_2594
		));
	notech_and4 i_787(.A(n_2162), .B(n_30726), .C(n_30691), .D(n_30725), .Z(n_2591
		));
	notech_and3 i_598(.A(n_3970), .B(n_1806), .C(n_30696), .Z(n_2588));
	notech_and2 i_152(.A(n_1825), .B(n_2070), .Z(n_2587));
	notech_or4 i_1069(.A(n_58498), .B(n_2283), .C(n_30738), .D(n_30851), .Z(n_2586
		));
	notech_and3 i_223(.A(n_3979), .B(n_30722), .C(n_1978), .Z(n_2579));
	notech_or4 i_910(.A(n_58498), .B(n_30842), .C(n_30841), .D(adz), .Z(n_2577
		));
	notech_or4 i_663(.A(n_58581), .B(n_58550), .C(n_30845), .D(n_30779), .Z(n_2574
		));
	notech_and4 i_378(.A(n_1984), .B(n_1801), .C(n_4019), .D(n_30792), .Z(n_2572
		));
	notech_and2 i_517(.A(n_1984), .B(n_1801), .Z(n_2571));
	notech_and2 i_3478(.A(n_4019), .B(n_30792), .Z(n_2569));
	notech_and3 i_377(.A(n_2565), .B(n_2563), .C(n_2562), .Z(n_2567));
	notech_and3 i_759(.A(n_4067), .B(n_2166), .C(n_30713), .Z(n_2565));
	notech_or4 i_499(.A(n_58581), .B(n_2282), .C(n_58568), .D(n_30844), .Z(n_2564
		));
	notech_ao4 i_442(.A(n_2494), .B(n_2315), .C(n_2489), .D(n_2373), .Z(n_2563
		));
	notech_and4 i_723(.A(n_1873), .B(n_2555), .C(n_1874), .D(n_1800), .Z(n_2562
		));
	notech_or4 i_108(.A(n_2497), .B(n_2333), .C(modrm[1]), .D(modrm[0]), .Z(n_2560
		));
	notech_or4 i_109(.A(n_2497), .B(n_2333), .C(modrm[1]), .D(n_30847), .Z(n_2557
		));
	notech_and2 i_291(.A(n_1869), .B(n_1871), .Z(n_2555));
	notech_or2 i_496(.A(n_2497), .B(n_2333), .Z(n_2553));
	notech_and4 i_1101(.A(n_2510), .B(n_2500), .C(n_2547), .D(n_2498), .Z(n_2549
		));
	notech_and4 i_1095(.A(n_2534), .B(n_2522), .C(n_2526), .D(n_2545), .Z(n_2547
		));
	notech_and4 i_1088(.A(n_2538), .B(n_2111), .C(n_3982), .D(n_2543), .Z(n_2545
		));
	notech_and2 i_433(.A(n_3880), .B(n_30665), .Z(n_2543));
	notech_nor2 i_832(.A(n_2486), .B(n_2288), .Z(n_2542));
	notech_ao3 i_829(.A(modrm[2]), .B(n_2287), .C(n_2333), .Z(n_2541));
	notech_and3 i_608(.A(n_1798), .B(n_1796), .C(n_2111), .Z(n_2539));
	notech_and2 i_190(.A(n_1798), .B(n_1796), .Z(n_2538));
	notech_and4 i_84(.A(n_58482), .B(n_2431), .C(n_30842), .D(n_30851), .Z(n_2536
		));
	notech_and4 i_362(.A(n_2206), .B(n_4028), .C(n_2532), .D(n_3777), .Z(n_2534
		));
	notech_and4 i_638(.A(n_2206), .B(n_4028), .C(n_3992), .D(n_2123), .Z(n_2533
		));
	notech_and2 i_423(.A(n_3992), .B(n_2123), .Z(n_2532));
	notech_nand2 i_963(.A(n_30841), .B(n_30659), .Z(n_2531));
	notech_and4 i_83(.A(n_2431), .B(n_58482), .C(n_30842), .D(modrm[5]), .Z(n_2530
		));
	notech_and4 i_315(.A(n_3665), .B(n_2216), .C(n_3672), .D(n_2212), .Z(n_2526
		));
	notech_nand3 i_833(.A(n_2310), .B(n_30660), .C(n_58568), .Z(n_2523));
	notech_and4 i_298(.A(n_4004), .B(n_2398), .C(n_2513), .D(n_2518), .Z(n_2522
		));
	notech_or4 i_187(.A(n_58581), .B(n_2244), .C(n_58550), .D(n_30845), .Z(n_2519
		));
	notech_and2 i_713(.A(n_2516), .B(n_1890), .Z(n_2518));
	notech_or4 i_495(.A(n_58581), .B(n_2289), .C(n_58550), .D(n_30845), .Z(n_2517
		));
	notech_and2 i_903(.A(n_2515), .B(n_2032), .Z(n_2516));
	notech_or4 i_580(.A(n_2279), .B(n_58498), .C(n_30844), .D(n_58592), .Z(n_2515
		));
	notech_and2 i_703(.A(n_2234), .B(n_4005), .Z(n_2513));
	notech_and2 i_392(.A(n_2289), .B(n_30779), .Z(n_2512));
	notech_and4 i_380(.A(n_1901), .B(n_4087), .C(n_2198), .D(n_3972), .Z(n_2510
		));
	notech_or4 i_991(.A(n_2410), .B(modrm[3]), .C(modrm[4]), .D(modrm[5]), .Z
		(n_2505));
	notech_xor2 i_432(.A(n_30852), .B(modrm[7]), .Z(n_2504));
	notech_or4 i_90(.A(n_2410), .B(modrm[3]), .C(n_30850), .D(n_30851), .Z(n_2501
		));
	notech_and2 i_213(.A(n_3834), .B(n_3984), .Z(n_2500));
	notech_or4 i_87(.A(n_2386), .B(n_2315), .C(n_30844), .D(n_30851), .Z(n_2499
		));
	notech_and2 i_771(.A(n_1993), .B(n_1915), .Z(n_2498));
	notech_or4 i_48(.A(n_2329), .B(n_2292), .C(n_58601), .D(n_58592), .Z(n_2497
		));
	notech_and2 i_418(.A(n_2373), .B(n_2372), .Z(n_2495));
	notech_or4 i_578(.A(n_2486), .B(n_2485), .C(modrm[1]), .D(n_30847), .Z(n_2494
		));
	notech_and2 i_403(.A(n_30849), .B(n_30850), .Z(n_2492));
	notech_or4 i_885(.A(n_58550), .B(n_30806), .C(n_30851), .D(modrm[1]), .Z
		(n_2490));
	notech_or2 i_106(.A(n_2488), .B(modrm[0]), .Z(n_2489));
	notech_or4 i_836(.A(n_2325), .B(n_2485), .C(n_30851), .D(n_30848), .Z(n_2488
		));
	notech_or4 i_40(.A(n_58581), .B(n_58568), .C(n_58550), .D(n_30851), .Z(n_2486
		));
	notech_or4 i_49(.A(n_2329), .B(n_2300), .C(n_58601), .D(n_58592), .Z(n_2485
		));
	notech_and4 i_799(.A(n_1919), .B(n_3998), .C(n_30720), .D(n_30724), .Z(n_2484
		));
	notech_and4 i_319(.A(n_3967), .B(n_2480), .C(n_2479), .D(n_2415), .Z(n_2483
		));
	notech_ao4 i_129(.A(n_2027), .B(n_2393), .C(n_2346), .D(n_2387), .Z(n_2480
		));
	notech_and2 i_611(.A(n_3876), .B(n_4022), .Z(n_2479));
	notech_nand3 i_803(.A(n_2450), .B(n_2036), .C(n_2474), .Z(n_2475));
	notech_and3 i_795(.A(n_247292237), .B(n_2465), .C(n_1848), .Z(n_2474));
	notech_and3 i_800(.A(n_4025), .B(n_30709), .C(n_30707), .Z(n_247292237)
		);
	notech_and2 i_831(.A(cpl[1]), .B(cpl[0]), .Z(n_2469));
	notech_ao3 i_408(.A(n_58581), .B(n_2272), .C(n_2383), .Z(n_2466));
	notech_and4 i_504(.A(n_3965), .B(n_30726), .C(n_30691), .D(n_30725), .Z(n_2465
		));
	notech_or4 i_530(.A(n_58498), .B(n_30738), .C(n_58514), .D(n_30841), .Z(n_2464
		));
	notech_and4 i_119(.A(n_2189), .B(n_2206), .C(n_2179), .D(n_2457), .Z(n_2463
		));
	notech_or4 i_528(.A(n_58581), .B(n_58568), .C(n_58550), .D(n_30729), .Z(n_2458
		));
	notech_and3 i_316(.A(n_2255), .B(n_1805), .C(n_3975), .Z(n_2457));
	notech_or4 i_99(.A(n_58498), .B(n_58550), .C(n_30806), .D(n_58514), .Z(n_2455
		));
	notech_ao3 i_470(.A(n_3970), .B(n_1806), .C(n_1807), .Z(n_2450));
	notech_nand3 i_150(.A(n_2310), .B(n_58568), .C(n_30653), .Z(n_2448));
	notech_or4 i_849(.A(n_58497), .B(n_2311), .C(n_58514), .D(n_58519), .Z(n_2447
		));
	notech_nao3 i_457(.A(n_58601), .B(n_58592), .C(n_2311), .Z(n_2446));
	notech_or4 i_801(.A(n_30700), .B(n_30783), .C(n_2442), .D(n_3986), .Z(n_2445
		));
	notech_nao3 i_784(.A(n_2440), .B(n_2430), .C(n_1846), .Z(n_2442));
	notech_and4 i_775(.A(n_1843), .B(n_2437), .C(n_2140), .D(n_30724), .Z(n_2440
		));
	notech_and4 i_761(.A(n_2435), .B(n_1960), .C(n_3993), .D(n_2305), .Z(n_2437
		));
	notech_and2 i_44973062(.A(n_2234), .B(n_2398), .Z(n_2435));
	notech_and2 i_69073044(.A(n_3993), .B(n_2305), .Z(n_2434));
	notech_or2 i_250(.A(n_2403), .B(n_2389), .Z(n_2433));
	notech_nor2 i_579(.A(n_58581), .B(n_2403), .Z(n_2431));
	notech_ao4 i_773(.A(n_30842), .B(n_1842), .C(n_2383), .D(n_2428), .Z(n_2430
		));
	notech_or4 i_527(.A(n_58482), .B(n_58470), .C(n_30844), .D(n_30806), .Z(n_2428
		));
	notech_and3 i_674(.A(n_30844), .B(n_2324), .C(n_2369), .Z(n_2427));
	notech_and4 i_636(.A(n_4062), .B(n_4093), .C(n_30695), .D(n_30706), .Z(n_2426
		));
	notech_or4 i_352(.A(n_2386), .B(n_2372), .C(n_58537), .D(n_30851), .Z(n_2422
		));
	notech_and4 i_127(.A(n_58581), .B(n_30845), .C(n_58537), .D(n_2354), .Z(n_2418
		));
	notech_and2 i_594(.A(n_1938), .B(n_1835), .Z(n_2417));
	notech_and3 i_450(.A(n_2137), .B(n_2045), .C(n_2411), .Z(n_2415));
	notech_and2 i_307(.A(n_2137), .B(n_2045), .Z(n_2414));
	notech_and2 i_398(.A(n_2302), .B(n_30801), .Z(n_2413));
	notech_or4 i_194(.A(n_58492), .B(n_2325), .C(n_58532), .D(n_30842), .Z(n_2412
		));
	notech_and3 i_142(.A(n_2231), .B(n_1833), .C(n_2026), .Z(n_2411));
	notech_nao3 i_730(.A(n_30842), .B(n_58532), .C(n_2276), .Z(n_2408));
	notech_or4 i_77(.A(n_58581), .B(n_2290), .C(n_58550), .D(n_30845), .Z(n_2407
		));
	notech_and4 i_246(.A(n_2395), .B(n_2402), .C(n_2392), .D(n_2379), .Z(n_2406
		));
	notech_ao4 i_725(.A(n_2401), .B(n_3958), .C(n_3963), .D(n_2396), .Z(n_2402
		));
	notech_or4 i_67(.A(n_2329), .B(n_58592), .C(n_58482), .D(n_30659), .Z(n_2401
		));
	notech_and2 i_390(.A(n_30791), .B(n_2399), .Z(n_2400));
	notech_or4 i_96(.A(n_2410), .B(n_30849), .C(n_30850), .D(modrm[5]), .Z(n_2399
		));
	notech_or4 i_691(.A(n_58577), .B(n_2299), .C(n_58568), .D(n_58546), .Z(n_2396
		));
	notech_and3 i_434(.A(n_1829), .B(n_1828), .C(n_1958), .Z(n_2395));
	notech_ao4 i_132(.A(n_2297), .B(n_2393), .C(n_2346), .D(n_2299), .Z(n_2394
		));
	notech_or4 i_107(.A(n_2347), .B(n_2313), .C(n_2282), .D(n_30845), .Z(n_2393
		));
	notech_ao4 i_778(.A(n_2391), .B(n_2387), .C(n_30787), .D(n_4090), .Z(n_2392
		));
	notech_and2 i_429(.A(n_30703), .B(n_30789), .Z(n_2391));
	notech_and4 i_100(.A(n_58577), .B(n_30845), .C(n_58546), .D(n_2354), .Z(n_2390
		));
	notech_nand3 i_664(.A(n_58577), .B(n_30845), .C(n_58546), .Z(n_2389));
	notech_and2 i_185(.A(n_2278), .B(n_2299), .Z(n_2387));
	notech_nand2 i_369(.A(n_58577), .B(n_58568), .Z(n_2386));
	notech_nand2 i_419(.A(n_2372), .B(n_2315), .Z(n_2385));
	notech_nao3 i_95(.A(modrm[6]), .B(modrm[7]), .C(n_2381), .Z(n_2384));
	notech_or4 i_85(.A(n_2329), .B(n_58482), .C(n_58470), .D(n_2271), .Z(n_2382
		));
	notech_or4 i_661(.A(n_58492), .B(n_2283), .C(n_58482), .D(n_58470), .Z(n_2381
		));
	notech_and4 i_325(.A(n_4031), .B(n_4056), .C(n_4084), .D(n_2377), .Z(n_2379
		));
	notech_and2 i_339(.A(n_4066), .B(n_30687), .Z(n_2377));
	notech_or4 i_344(.A(n_2286), .B(n_30659), .C(n_2346), .D(n_30851), .Z(n_2376
		));
	notech_nor2 i_705(.A(n_2346), .B(n_58390), .Z(n_2375));
	notech_xor2 i_389(.A(n_30850), .B(modrm[3]), .Z(n_2374));
	notech_nand2 i_46(.A(n_30849), .B(modrm[4]), .Z(n_2373));
	notech_nand2 i_183(.A(n_30849), .B(n_30850), .Z(n_2372));
	notech_or4 i_693(.A(n_2279), .B(n_58532), .C(n_30842), .D(n_58537), .Z(n_2371
		));
	notech_and2 i_168(.A(n_1817), .B(n_2364), .Z(n_2365));
	notech_and2 i_756(.A(n_3991), .B(n_1813), .Z(n_2364));
	notech_and2 i_459(.A(n_2275), .B(n_2302), .Z(n_2363));
	notech_or4 i_86(.A(n_2347), .B(n_2360), .C(n_2282), .D(n_30845), .Z(n_2362
		));
	notech_nand2 i_535(.A(n_58519), .B(n_58514), .Z(n_2360));
	notech_or4 i_71(.A(n_2329), .B(n_58601), .C(n_58592), .D(n_2271), .Z(n_2359
		));
	notech_or4 i_66(.A(n_2329), .B(n_58592), .C(n_58482), .D(n_2271), .Z(n_2355
		));
	notech_and4 i_64(.A(n_223492236), .B(n_1792), .C(n_30699), .D(n_1797), .Z
		(n_2352));
	notech_or4 i_577(.A(n_2348), .B(n_2284), .C(n_30779), .D(n_30659), .Z(n_2350
		));
	notech_nor2 i_111(.A(n_2348), .B(n_2284), .Z(n_2349));
	notech_nao3 i_13(.A(n_58537), .B(n_58564), .C(n_58577), .Z(n_2348));
	notech_or2 i_600(.A(n_58577), .B(n_58546), .Z(n_2347));
	notech_or4 i_79(.A(n_2282), .B(n_2280), .C(n_58514), .D(n_58519), .Z(n_2346
		));
	notech_and4 i_351(.A(n_2141), .B(n_4013), .C(n_2058), .D(n_2343), .Z(n_2344
		));
	notech_and4 i_683(.A(n_2340), .B(n_2233), .C(n_2195), .D(n_2099), .Z(n_2343
		));
	notech_and2 i_513(.A(n_4044), .B(n_30721), .Z(n_2340));
	notech_nao3 i_671(.A(n_58573), .B(n_2272), .C(n_2338), .Z(n_2339));
	notech_nao3 i_151(.A(n_30842), .B(n_58519), .C(n_2282), .Z(n_2338));
	notech_or4 i_585(.A(n_2316), .B(n_2276), .C(n_2037), .D(n_2333), .Z(n_2337
		));
	notech_or4 i_32(.A(n_58573), .B(n_58564), .C(n_58546), .D(modrm[5]), .Z(n_2333
		));
	notech_nao3 i_574(.A(modrm[7]), .B(modrm[6]), .C(n_2290), .Z(n_2331));
	notech_or4 i_121(.A(n_58487), .B(n_2283), .C(n_58601), .D(n_58470), .Z(n_2330
		));
	notech_nao3 i_1(.A(n_58514), .B(n_58532), .C(n_58487), .Z(n_2329));
	notech_or4 i_0(.A(twobyte), .B(fpu), .C(ipg_fault), .D(n_30846), .Z(n_2328
		));
	notech_nao3 i_3(.A(n_58555), .B(n_58537), .C(n_58573), .Z(n_2325));
	notech_nor2 i_449(.A(n_58577), .B(n_58564), .Z(n_2324));
	notech_nor2 i_599(.A(opz[0]), .B(opz[2]), .Z(n_2322));
	notech_and2 i_73(.A(opz[2]), .B(n_2319), .Z(n_2321));
	notech_nor2 i_597(.A(opz[0]), .B(opz[1]), .Z(n_2319));
	notech_or4 i_92(.A(n_2403), .B(n_2311), .C(n_58514), .D(n_58532), .Z(n_2318
		));
	notech_nand2 i_584(.A(n_30842), .B(n_58519), .Z(n_2316));
	notech_nand2 i_446(.A(n_58456), .B(n_58532), .Z(n_2313));
	notech_nand3 i_41(.A(n_58573), .B(n_58537), .C(n_58564), .Z(n_2311));
	notech_and2 i_382(.A(n_58577), .B(n_58537), .Z(n_2310));
	notech_and4 i_436(.A(n_2141), .B(n_4013), .C(n_2308), .D(n_2294), .Z(n_2309
		));
	notech_and3 i_657(.A(n_4037), .B(n_1820), .C(n_1824), .Z(n_2308));
	notech_ao4 i_405(.A(n_2290), .B(n_2300), .C(n_2289), .D(n_30659), .Z(n_2303
		));
	notech_ao3 i_91(.A(n_58482), .B(n_58470), .C(n_2300), .Z(n_2301));
	notech_nao3 i_282(.A(modrm[7]), .B(modrm[6]), .C(modrm[2]), .Z(n_2300)
		);
	notech_nand3 i_68(.A(n_58465), .B(n_58601), .C(n_2271), .Z(n_2299));
	notech_nand3 i_59(.A(n_58601), .B(n_58592), .C(n_2271), .Z(n_2297));
	notech_and2 i_5(.A(n_58597), .B(n_58592), .Z(n_2296));
	notech_nao3 i_468(.A(modrm[2]), .B(n_2271), .C(n_2286), .Z(n_2295));
	notech_and2 i_790(.A(n_2258), .B(n_1821), .Z(n_2294));
	notech_nao3 i_88(.A(n_58482), .B(n_58465), .C(n_2292), .Z(n_2293));
	notech_nand3 i_276(.A(modrm[7]), .B(modrm[2]), .C(modrm[6]), .Z(n_2292)
		);
	notech_and2 i_393(.A(n_2278), .B(n_30702), .Z(n_2291));
	notech_nand2 i_2(.A(n_58481), .B(n_58465), .Z(n_2290));
	notech_nand2 i_6(.A(n_58465), .B(n_58597), .Z(n_2289));
	notech_or4 i_590(.A(modrm[2]), .B(n_58597), .C(n_58465), .D(n_30659), .Z
		(n_2288));
	notech_and4 i_120(.A(modrm[7]), .B(n_58476), .C(n_58592), .D(modrm[6]), 
		.Z(n_2287));
	notech_nand2 i_773161(.A(n_58476), .B(n_58592), .Z(n_2286));
	notech_or4 i_75(.A(n_58363), .B(n_2280), .C(n_58456), .D(n_58519), .Z(n_2285
		));
	notech_nao3 i_856(.A(n_58510), .B(n_58532), .C(n_58363), .Z(n_2284));
	notech_nand2 i_589(.A(n_58510), .B(n_58532), .Z(n_2283));
	notech_or4 i_9(.A(fpu), .B(ipg_fault), .C(n_30846), .D(n_30854), .Z(n_2282
		));
	notech_nao3 i_44(.A(n_58564), .B(n_58546), .C(n_58577), .Z(n_2280));
	notech_or2 i_593(.A(n_58577), .B(n_58555), .Z(n_2279));
	notech_or4 i_857(.A(fpu), .B(ipg_fault), .C(op[7]), .D(n_30854), .Z(n_2276
		));
	notech_and2 i_537(.A(n_58555), .B(n_58537), .Z(n_2272));
	notech_and2 i_230(.A(modrm[7]), .B(modrm[6]), .Z(n_2271));
	notech_and4 i_281(.A(n_3591), .B(n_3560), .C(n_717), .D(n_1593), .Z(n_2270
		));
	notech_or2 i_2397(.A(n_2398), .B(n_58476), .Z(n_2269));
	notech_nand3 i_308(.A(n_2757), .B(n_3548), .C(n_1951), .Z(\udeco[8] ));
	notech_nand2 i_2345(.A(modrm[3]), .B(n_3174), .Z(n_2267));
	notech_nao3 i_2349(.A(opz[1]), .B(n_2322), .C(n_2247), .Z(n_2266));
	notech_or4 i_2341(.A(n_2410), .B(n_2373), .C(n_3954), .D(n_58390), .Z(n_2265
		));
	notech_or2 i_335(.A(n_2485), .B(n_2333), .Z(n_2264));
	notech_or4 i_2350(.A(n_58492), .B(n_2248), .C(n_58510), .D(n_58532), .Z(n_2263
		));
	notech_nand2 i_2353(.A(n_58586), .B(n_2251), .Z(n_2262));
	notech_or4 i_144(.A(n_2286), .B(modrm[2]), .C(n_2285), .D(n_58399), .Z(n_2258
		));
	notech_or4 i_2344(.A(n_2412), .B(n_58476), .C(n_58465), .D(n_2271), .Z(n_2257
		));
	notech_or4 i_2342(.A(n_58492), .B(n_2316), .C(n_2389), .D(n_2278), .Z(n_2256
		));
	notech_or4 i_23111195(.A(n_2313), .B(n_58476), .C(n_2271), .D(n_30799), 
		.Z(n_2255));
	notech_or4 i_2351(.A(n_58492), .B(n_58528), .C(n_58456), .D(n_2249), .Z(n_2254
		));
	notech_or4 i_2346(.A(n_2347), .B(n_2338), .C(n_2512), .D(n_58555), .Z(n_2253
		));
	notech_or4 i_822(.A(n_2280), .B(n_58492), .C(n_58586), .D(n_58510), .Z(n_2252
		));
	notech_nand2 i_202(.A(n_2433), .B(n_2678), .Z(n_2251));
	notech_and3 i_203(.A(n_2141), .B(n_4013), .C(n_2140), .Z(n_2250));
	notech_and2 i_205(.A(n_2448), .B(n_2243), .Z(n_2249));
	notech_ao4 i_209(.A(n_2486), .B(n_2288), .C(n_2348), .D(n_2289), .Z(n_2248
		));
	notech_ao4 i_219(.A(n_2318), .B(n_2297), .C(n_2401), .D(n_2101), .Z(n_2247
		));
	notech_ao3 i_222(.A(n_2275), .B(n_2302), .C(n_2301), .Z(n_2245));
	notech_and2 i_404(.A(n_58372), .B(n_30779), .Z(n_2244));
	notech_nao3 i_2339(.A(n_2310), .B(n_58564), .C(n_2244), .Z(n_2243));
	notech_and4 i_320(.A(n_2484), .B(n_2703), .C(n_3500), .D(n_3465), .Z(n_2241
		));
	notech_nand2 i_2293(.A(n_3174), .B(modrm[4]), .Z(n_2240));
	notech_or4 i_2294(.A(n_2410), .B(n_2373), .C(n_2230), .D(n_58390), .Z(n_2239
		));
	notech_or4 i_287(.A(n_2383), .B(n_2486), .C(n_2290), .D(n_2300), .Z(n_2238
		));
	notech_nand2 i_2291(.A(n_58546), .B(n_30766), .Z(n_2237));
	notech_or4 i_23111324(.A(n_2348), .B(n_2320), .C(n_2275), .D(n_2284), .Z
		(n_223492236));
	notech_or4 i_23111438(.A(n_58399), .B(n_2337), .C(n_58597), .D(n_58586),
		 .Z(n_2233));
	notech_or4 i_2290(.A(n_2285), .B(n_58476), .C(n_58465), .D(n_2271), .Z(n_2232
		));
	notech_or4 i_23111390(.A(n_2347), .B(n_2290), .C(n_2408), .D(n_58555), .Z
		(n_2231));
	notech_and2 i_200(.A(n_2382), .B(n_2485), .Z(n_2230));
	notech_or4 i_2286(.A(n_58372), .B(n_2329), .C(n_2325), .D(n_58417), .Z(n_2229
		));
	notech_or4 i_2285(.A(n_2285), .B(n_58586), .C(n_58476), .D(n_58399), .Z(n_2228
		));
	notech_and4 i_334(.A(n_2694), .B(n_3458), .C(n_3429), .D(n_2704), .Z(n_2227
		));
	notech_nand2 i_2248(.A(n_3174), .B(modrm[5]), .Z(n_2226));
	notech_nao3 i_2249(.A(n_30658), .B(n_30790), .C(n_2499), .Z(n_2223));
	notech_or2 i_2243(.A(n_2065), .B(n_58456), .Z(n_2222));
	notech_or4 i_2247(.A(n_2360), .B(n_58487), .C(n_58381), .D(n_2297), .Z(n_2221
		));
	notech_or4 i_2250(.A(n_2316), .B(n_2276), .C(n_2289), .D(n_2280), .Z(n_2220
		));
	notech_and4 i_345(.A(n_2904), .B(n_2703), .C(n_2484), .D(n_3425), .Z(n_221992235
		));
	notech_or4 i_149(.A(n_2244), .B(n_2185), .C(n_58537), .D(n_2386), .Z(n_2218
		));
	notech_or2 i_2216(.A(n_2065), .B(n_58465), .Z(n_2217));
	notech_or4 i_23110652(.A(n_2329), .B(n_58586), .C(n_58476), .D(n_2389), 
		.Z(n_2216));
	notech_and4 i_431(.A(n_2689), .B(n_2501), .C(n_2499), .D(n_2422), .Z(n_2215
		));
	notech_or2 i_2215(.A(n_2215), .B(n_2359), .Z(n_2213));
	notech_and4 i_363(.A(n_2484), .B(n_3397), .C(n_2904), .D(n_2704), .Z(n_2208
		));
	notech_or2 i_2183(.A(n_2215), .B(n_2497), .Z(n_2207));
	notech_or4 i_23111192(.A(n_2316), .B(n_58476), .C(n_30799), .D(n_58417),
		 .Z(n_2206));
	notech_and2 i_353(.A(n_2295), .B(n_2293), .Z(n_2205));
	notech_or4 i_361(.A(n_58372), .B(n_2292), .C(n_2329), .D(n_30787), .Z(n_2202
		));
	notech_nand3 i_385(.A(n_3364), .B(n_3343), .C(n_1951), .Z(\udeco[16] )
		);
	notech_nao3 i_2126(.A(opz[1]), .B(n_2322), .C(n_2187), .Z(n_2200));
	notech_or2 i_2123(.A(n_2883), .B(n_30849), .Z(n_2199));
	notech_or2 i_297(.A(n_4090), .B(n_30787), .Z(n_2198));
	notech_or4 i_2125(.A(n_2373), .B(n_58390), .C(n_2410), .D(n_2115), .Z(n_2197
		));
	notech_or4 i_2120(.A(n_58354), .B(n_2037), .C(n_3954), .D(n_58390), .Z(n_2196
		));
	notech_or4 i_153(.A(n_58577), .B(n_2330), .C(n_58568), .D(n_58546), .Z(n_2195
		));
	notech_or4 i_2119(.A(n_2292), .B(n_2285), .C(n_58597), .D(n_58586), .Z(n_2193
		));
	notech_or4 i_677(.A(n_30738), .B(n_58586), .C(n_58476), .D(n_30785), .Z(n_2192
		));
	notech_or2 i_2982(.A(n_2300), .B(n_30777), .Z(n_2190));
	notech_or4 i_1241(.A(n_58476), .B(n_30799), .C(n_58510), .D(n_58399), .Z
		(n_2189));
	notech_or4 i_179(.A(n_58577), .B(n_2403), .C(n_2360), .D(n_58597), .Z(n_2188
		));
	notech_ao4 i_181(.A(n_4065), .B(n_2297), .C(n_2098), .D(n_2101), .Z(n_2187
		));
	notech_and2 i_524(.A(n_2668), .B(n_3154), .Z(n_2186));
	notech_and3 i_394(.A(n_2383), .B(n_30785), .C(n_30729), .Z(n_2185));
	notech_or4 i_2116(.A(n_2285), .B(n_58597), .C(n_58586), .D(n_58417), .Z(n_2183
		));
	notech_nao3 i_2115(.A(opz[1]), .B(n_2322), .C(n_2350), .Z(n_2181));
	notech_nand3 i_2110(.A(n_3895), .B(n_58568), .C(n_2310), .Z(n_2180));
	notech_or4 i_39(.A(n_2458), .B(n_58481), .C(n_58465), .D(n_58417), .Z(n_2179
		));
	notech_and4 i_400(.A(n_3309), .B(n_3302), .C(n_3273), .D(n_2562), .Z(n_2177
		));
	notech_or2 i_2061(.A(n_2883), .B(n_30850), .Z(n_2175));
	notech_or4 i_2060(.A(n_58354), .B(n_2373), .C(n_3836), .D(n_58390), .Z(n_2174
		));
	notech_nand2 i_2064(.A(n_58546), .B(n_30812), .Z(n_2173));
	notech_nao3 i_2062(.A(n_2321), .B(n_30793), .C(n_2101), .Z(n_2172));
	notech_or4 i_2063(.A(n_2403), .B(n_2161), .C(n_2313), .D(n_2311), .Z(n_2170
		));
	notech_or4 i_2058(.A(n_58354), .B(n_2037), .C(n_58390), .D(n_2355), .Z(n_2169
		));
	notech_nao3 i_2056(.A(n_2385), .B(n_30656), .C(n_2214), .Z(n_2168));
	notech_or4 i_227(.A(n_58381), .B(n_58417), .C(n_30779), .D(n_30785), .Z(n_2166
		));
	notech_or4 i_2059(.A(n_58597), .B(n_58586), .C(n_58417), .D(n_30703), .Z
		(n_2163));
	notech_ao4 i_518(.A(n_2297), .B(n_30807), .C(n_2275), .D(n_2149), .Z(n_2161
		));
	notech_or4 i_224(.A(n_58372), .B(n_2486), .C(n_58417), .D(n_30729), .Z(n_2159
		));
	notech_or4 i_2050(.A(n_58487), .B(n_2594), .C(n_58510), .D(n_58528), .Z(n_2155
		));
	notech_and2 i_290(.A(n_2285), .B(n_30703), .Z(n_2154));
	notech_and2 i_328(.A(n_2320), .B(n_30807), .Z(n_2149));
	notech_and4 i_414(.A(n_2757), .B(n_3257), .C(n_1504), .D(n_520), .Z(n_2146
		));
	notech_or2 i_2004(.A(n_2883), .B(n_58390), .Z(n_2145));
	notech_or4 i_2002(.A(n_58354), .B(n_2037), .C(n_3836), .D(n_58390), .Z(n_2144
		));
	notech_nand2 i_2005(.A(n_58568), .B(n_30812), .Z(n_2143));
	notech_and3 i_2003(.A(n_2287), .B(n_2375), .C(n_2385), .Z(n_2142));
	notech_nao3 i_1250(.A(n_2397), .B(n_58417), .C(n_2276), .Z(n_2141));
	notech_or4 i_180(.A(n_58577), .B(n_2403), .C(n_2283), .D(n_58564), .Z(n_2140
		));
	notech_and3 i_326(.A(n_2485), .B(n_2401), .C(n_2497), .Z(n_2139));
	notech_or4 i_675(.A(n_58408), .B(n_58487), .C(n_58381), .D(n_2027), .Z(n_2137
		));
	notech_or2 i_591(.A(n_2497), .B(n_30787), .Z(n_2136));
	notech_and4 i_438(.A(n_530), .B(n_2703), .C(n_3213), .D(n_537), .Z(n_2135
		));
	notech_or4 i_1968(.A(n_58354), .B(n_2373), .C(n_3954), .D(modrm[5]), .Z(n_2134
		));
	notech_or4 i_1967(.A(n_58597), .B(n_58586), .C(n_58417), .D(n_30800), .Z
		(n_2132));
	notech_nao3 i_1935(.A(n_30849), .B(n_30850), .C(n_2376), .Z(n_2131));
	notech_or4 i_1934(.A(n_58354), .B(n_2373), .C(n_2384), .D(n_58390), .Z(n_2130
		));
	notech_or4 i_1933(.A(n_58408), .B(n_58487), .C(n_58381), .D(n_2302), .Z(n_2129
		));
	notech_ao3 i_1931(.A(n_2299), .B(n_2297), .C(n_2301), .Z(n_2128));
	notech_and4 i_48310343(.A(n_719), .B(n_3171), .C(n_3143), .D(n_1950), .Z
		(n_2127));
	notech_nand3 i_1902(.A(opz[1]), .B(n_2322), .C(n_2117), .Z(n_2126));
	notech_or2 i_1898(.A(n_3728), .B(n_30849), .Z(n_2125));
	notech_or4 i_1901(.A(n_58354), .B(n_2037), .C(n_2115), .D(n_58390), .Z(n_2122
		));
	notech_or2 i_1899(.A(n_3697), .B(n_58465), .Z(n_2121));
	notech_or2 i_1897(.A(n_2151), .B(n_58481), .Z(n_2120));
	notech_or2 i_1900(.A(n_2052), .B(n_30702), .Z(n_2119));
	notech_nand2 i_169(.A(n_2988), .B(n_2350), .Z(n_2117));
	notech_and3 i_174(.A(n_2497), .B(n_2359), .C(n_2355), .Z(n_2115));
	notech_nand3 i_124(.A(n_58399), .B(n_58528), .C(n_2536), .Z(n_2111));
	notech_nao3 i_472(.A(n_1718), .B(n_3141), .C(n_4024), .Z(\udeco[25] ));
	notech_nand2 i_1860(.A(modrm[4]), .B(n_30715), .Z(n_2109));
	notech_or4 i_838(.A(n_58577), .B(n_58564), .C(n_58546), .D(n_2098), .Z(n_2108
		));
	notech_nand2 i_1861(.A(n_58546), .B(n_30716), .Z(n_2107));
	notech_nao3 i_1197(.A(opz[2]), .B(n_2319), .C(n_2350), .Z(n_2106));
	notech_or2 i_1858(.A(n_2151), .B(n_58519), .Z(n_2105));
	notech_nao3 i_827(.A(n_2287), .B(n_2375), .C(n_2374), .Z(n_2104));
	notech_or4 i_47(.A(n_2596), .B(n_58597), .C(n_58465), .D(n_58417), .Z(n_2103
		));
	notech_ao3 i_16373106(.A(opz[2]), .B(n_2319), .C(n_2083), .Z(n_2102));
	notech_and2 i_633(.A(n_2499), .B(n_2422), .Z(n_2101));
	notech_ao3 i_1824(.A(n_30658), .B(n_30662), .C(n_2499), .Z(n_2100));
	notech_and2 i_329(.A(n_2401), .B(n_2355), .Z(n_2098));
	notech_or4 i_1823(.A(n_58354), .B(n_2315), .C(n_3836), .D(n_58390), .Z(n_2097
		));
	notech_and4 i_1811(.A(n_2278), .B(n_2275), .C(n_30702), .D(n_2293), .Z(n_2095
		));
	notech_and4 i_546(.A(n_3091), .B(n_2903), .C(n_30838), .D(n_30798), .Z(n_2092
		));
	notech_or2 i_416(.A(n_3957), .B(n_2098), .Z(n_2091));
	notech_nao3 i_1775(.A(opz[1]), .B(n_2322), .C(n_2083), .Z(n_2090));
	notech_or4 i_1776(.A(n_2348), .B(n_58408), .C(n_58363), .D(n_2291), .Z(n_2089
		));
	notech_or4 i_1778(.A(n_2311), .B(n_3963), .C(n_58597), .D(n_58586), .Z(n_2087
		));
	notech_or4 i_1777(.A(n_58408), .B(n_2280), .C(n_58363), .D(n_30801), .Z(n_2086
		));
	notech_ao4 i_516(.A(n_2101), .B(n_2355), .C(n_4065), .D(n_2027), .Z(n_2083
		));
	notech_nand3 i_745(.A(n_3054), .B(n_2079), .C(n_30856), .Z(\udeco[108] )
		);
	notech_nand2 i_1646(.A(opz[0]), .B(n_2067), .Z(n_2079));
	notech_nor2 i_192(.A(n_2400), .B(n_3845), .Z(n_2078));
	notech_ao4 i_1647(.A(n_2418), .B(n_30803), .C(n_2301), .D(n_3908), .Z(n_2077
		));
	notech_or2 i_1648(.A(n_2359), .B(n_2069), .Z(n_2075));
	notech_or2 i_1645(.A(n_2523), .B(n_3961), .Z(n_2074));
	notech_or4 i_55(.A(modrm[2]), .B(n_2330), .C(n_58399), .D(n_30787), .Z(n_2073
		));
	notech_or4 i_1649(.A(n_2347), .B(n_58372), .C(n_3963), .D(n_58555), .Z(n_2072
		));
	notech_or4 i_23110742(.A(n_30738), .B(n_2329), .C(n_2331), .D(modrm[5]),
		 .Z(n_2071));
	notech_or4 i_23110745(.A(n_2586), .B(n_58601), .C(n_58586), .D(n_58399),
		 .Z(n_2070));
	notech_and3 i_163(.A(n_2400), .B(n_30738), .C(n_30787), .Z(n_2069));
	notech_nand3 i_165(.A(n_3018), .B(n_3013), .C(n_2955), .Z(n_2067));
	notech_or4 i_1629(.A(n_58487), .B(n_2574), .C(n_58510), .D(n_58519), .Z(n_2063
		));
	notech_nand2 i_1627(.A(n_2407), .B(n_2061), .Z(n_2062));
	notech_or4 i_254(.A(n_58577), .B(n_58372), .C(n_58546), .D(n_58555), .Z(n_2061
		));
	notech_and2 i_294(.A(n_2383), .B(n_2329), .Z(n_2059));
	notech_nao3 i_1622(.A(n_30660), .B(n_30855), .C(n_2407), .Z(n_2057));
	notech_or4 i_1620(.A(n_58487), .B(n_2407), .C(n_58510), .D(n_58528), .Z(n_2056
		));
	notech_and4 i_762(.A(n_3005), .B(n_2987), .C(n_2054), .D(n_30856), .Z(n_2055
		));
	notech_nand2 i_1590(.A(opz[1]), .B(n_30817), .Z(n_2054));
	notech_nao3 i_1586(.A(opz[1]), .B(n_2322), .C(n_2988), .Z(n_2053));
	notech_or2 i_1584(.A(adz), .B(n_2036), .Z(n_2051));
	notech_nao3 i_1585(.A(n_30847), .B(n_2037), .C(n_2488), .Z(n_2050));
	notech_or4 i_1228(.A(n_2485), .B(n_2490), .C(n_2492), .D(modrm[0]), .Z(n_2046
		));
	notech_or4 i_854(.A(n_58408), .B(n_58487), .C(n_58381), .D(n_2413), .Z(n_2045
		));
	notech_or4 i_1589(.A(n_58487), .B(n_2313), .C(n_2486), .D(n_2288), .Z(n_2042
		));
	notech_or4 i_1592(.A(n_58381), .B(n_3963), .C(n_58390), .D(n_2295), .Z(n_2041
		));
	notech_or4 i_1587(.A(n_58492), .B(n_2428), .C(n_58456), .D(n_58519), .Z(n_2040
		));
	notech_and4 i_158(.A(n_2309), .B(n_2958), .C(n_2975), .D(n_2955), .Z(n_2038
		));
	notech_nand2 i_564(.A(modrm[3]), .B(modrm[4]), .Z(n_2037));
	notech_and3 i_197(.A(n_2327), .B(n_4047), .C(n_3981), .Z(n_2036));
	notech_nand3 i_1566(.A(n_58577), .B(n_2272), .C(n_30662), .Z(n_2034));
	notech_or2 i_1567(.A(n_2523), .B(n_2512), .Z(n_2033));
	notech_or4 i_826(.A(n_2279), .B(n_58492), .C(n_58537), .D(n_58465), .Z(n_2032
		));
	notech_or4 i_1562(.A(n_2347), .B(n_2512), .C(n_58555), .D(n_2059), .Z(n_2031
		));
	notech_or4 i_1282(.A(n_2348), .B(n_58363), .C(n_1888), .D(n_58408), .Z(n_2030
		));
	notech_or4 i_1553(.A(n_3963), .B(n_2027), .C(n_58546), .D(n_30806), .Z(n_2028
		));
	notech_and2 i_301(.A(n_2275), .B(n_2297), .Z(n_2027));
	notech_or4 i_845(.A(n_2313), .B(n_58363), .C(n_2348), .D(n_2387), .Z(n_2026
		));
	notech_or4 i_1543(.A(n_2214), .B(n_2497), .C(modrm[3]), .D(n_30850), .Z(n_2025
		));
	notech_or4 i_1541(.A(n_2280), .B(n_58492), .C(n_58591), .D(n_58456), .Z(n_2021
		));
	notech_and4 i_796(.A(n_2939), .B(n_2936), .C(n_1718), .D(n_2890), .Z(n_2020
		));
	notech_or2 i_1174(.A(n_2400), .B(n_2401), .Z(n_2019));
	notech_or4 i_834(.A(n_58372), .B(n_58537), .C(n_30806), .D(n_30729), .Z(n_2014
		));
	notech_ao4 i_178(.A(n_2542), .B(n_2541), .C(n_2369), .D(n_2354), .Z(n_2013
		));
	notech_nand3 i_873(.A(n_2881), .B(n_1593), .C(n_2011), .Z(\udeco[117] )
		);
	notech_nand2 i_1366(.A(n_30768), .B(n_30819), .Z(n_2011));
	notech_nand2 i_1367(.A(modrm[4]), .B(n_3773), .Z(n_2010));
	notech_nand2 i_1368(.A(modrm[1]), .B(n_2007), .Z(n_2009));
	notech_or4 i_1365(.A(n_58363), .B(n_30738), .C(n_58470), .D(n_58519), .Z
		(n_2008));
	notech_nand3 i_140(.A(n_2099), .B(n_3736), .C(n_2654), .Z(n_2007));
	notech_mux2 i_396(.S(n_58528), .A(n_30850), .B(n_30848), .Z(n_2006));
	notech_or4 i_1361(.A(n_58408), .B(n_58492), .C(n_2519), .D(n_30855), .Z(n_2005
		));
	notech_or4 i_90810265(.A(n_2002), .B(n_2001), .C(n_2820), .D(n_1180), .Z
		(\udeco[120] ));
	notech_and2 i_1287(.A(n_3763), .B(n_1968), .Z(n_2002));
	notech_and2 i_1281(.A(n_30705), .B(n_30704), .Z(n_2001));
	notech_and2 i_1285(.A(modrm[0]), .B(n_30820), .Z(n_2000));
	notech_and2 i_1286(.A(modrm[3]), .B(n_1988), .Z(n_1998));
	notech_nor2 i_1288(.A(n_2362), .B(n_1989), .Z(n_1997));
	notech_or4 i_1141(.A(n_58408), .B(n_2280), .C(n_58363), .D(n_2413), .Z(n_1995
		));
	notech_or4 i_1280(.A(n_58497), .B(n_2517), .C(n_58514), .D(n_58528), .Z(n_1994
		));
	notech_or4 i_1284(.A(n_2347), .B(n_2338), .C(n_2244), .D(n_58555), .Z(n_1990
		));
	notech_and4 i_116(.A(n_2275), .B(n_2297), .C(n_2278), .D(n_2299), .Z(n_1989
		));
	notech_nand3 i_118(.A(n_2480), .B(n_1777), .C(n_2415), .Z(n_1988));
	notech_and4 i_655(.A(n_2309), .B(n_2760), .C(n_2717), .D(n_2759), .Z(n_1986
		));
	notech_or4 i_1275(.A(n_2315), .B(n_2214), .C(n_2330), .D(n_58399), .Z(n_1985
		));
	notech_or2 i_1273(.A(n_2382), .B(n_30787), .Z(n_1982));
	notech_or4 i_1272(.A(n_2372), .B(n_2214), .C(n_2330), .D(n_58399), .Z(n_1981
		));
	notech_or4 i_908(.A(n_1979), .B(n_1321), .C(n_1977), .D(n_2785), .Z(\udeco[121] 
		));
	notech_and2 i_1239(.A(n_1968), .B(n_30821), .Z(n_1979));
	notech_and2 i_1231(.A(n_30704), .B(n_30819), .Z(n_1977));
	notech_and2 i_1237(.A(modrm[1]), .B(n_30820), .Z(n_1976));
	notech_and2 i_1238(.A(modrm[4]), .B(n_1964), .Z(n_1975));
	notech_nand3 i_114(.A(n_2688), .B(n_2757), .C(n_2166), .Z(n_1968));
	notech_mux2 i_422(.S(n_58528), .A(n_30848), .B(n_30850), .Z(n_1965));
	notech_nand3 i_115(.A(n_2395), .B(n_1777), .C(n_2415), .Z(n_1964));
	notech_or4 i_483(.A(n_1326), .B(n_222994228), .C(n_1956), .D(n_30760), .Z
		(\udeco[122] ));
	notech_and2 i_1192(.A(modrm[2]), .B(n_1946), .Z(n_1956));
	notech_nand2 i_1191(.A(modrm[5]), .B(n_1945), .Z(n_1955));
	notech_nand2 i_1189(.A(n_1944), .B(n_30795), .Z(n_1954));
	notech_or4 i_1190(.A(n_2387), .B(n_58546), .C(n_30806), .D(n_30729), .Z(n_1952
		));
	notech_or4 i_1187(.A(n_58497), .B(n_58381), .C(n_58514), .D(n_3761), .Z(n_1949
		));
	notech_or2 i_1186(.A(n_2734), .B(n_58456), .Z(n_1947));
	notech_nand3 i_104(.A(n_2719), .B(n_2717), .C(n_2091), .Z(n_1946));
	notech_nand3 i_112(.A(n_2723), .B(n_4017), .C(n_2726), .Z(n_1945));
	notech_mux2 i_506(.S(n_58528), .A(n_58426), .B(modrm[2]), .Z(n_1944));
	notech_mux2 i_505(.S(n_58528), .A(modrm[2]), .B(n_58426), .Z(n_1943));
	notech_or2 i_1180(.A(n_1940), .B(n_2285), .Z(n_1941));
	notech_and4 i_113(.A(n_2027), .B(n_2387), .C(n_2302), .D(n_30702), .Z(n_1940
		));
	notech_or4 i_23111444(.A(n_58399), .B(n_2052), .C(n_58597), .D(n_58591),
		 .Z(n_1938));
	notech_and2 i_313(.A(n_2422), .B(n_2325), .Z(n_1937));
	notech_or4 i_1170(.A(n_2393), .B(n_58591), .C(n_58481), .D(n_30659), .Z(n_1936
		));
	notech_and4 i_1157(.A(n_58546), .B(n_2324), .C(n_2296), .D(n_30660), .Z(n_1933
		));
	notech_or2 i_1156(.A(n_2101), .B(n_2382), .Z(n_1932));
	notech_or2 i_1123(.A(n_3845), .B(n_30787), .Z(n_1930));
	notech_or4 i_1116(.A(n_58408), .B(n_58492), .C(n_30738), .D(n_2289), .Z(n_1921
		));
	notech_or4 i_1057(.A(n_2214), .B(n_2382), .C(n_30849), .D(n_30850), .Z(n_1919
		));
	notech_or4 i_1044(.A(n_2348), .B(n_30779), .C(adz), .D(n_2059), .Z(n_1918
		));
	notech_or4 i_284(.A(n_58492), .B(n_2286), .C(n_58528), .D(n_58456), .Z(n_1917
		));
	notech_and2 i_1042(.A(n_2330), .B(n_1917), .Z(n_1916));
	notech_or2 i_1030(.A(n_3836), .B(n_30787), .Z(n_1915));
	notech_or2 i_1028(.A(n_2494), .B(n_1913), .Z(n_1914));
	notech_and3 i_311(.A(n_2373), .B(n_2372), .C(n_2037), .Z(n_1913));
	notech_nao3 i_1027(.A(n_30847), .B(n_2385), .C(n_2488), .Z(n_1912));
	notech_or2 i_1018(.A(n_2497), .B(n_2486), .Z(n_1911));
	notech_or4 i_1011(.A(n_58528), .B(n_58456), .C(n_58481), .D(n_30799), .Z
		(n_1907));
	notech_ao4 i_1003(.A(n_2037), .B(n_2486), .C(n_58537), .D(n_2279), .Z(n_1902
		));
	notech_or4 i_992(.A(n_2330), .B(modrm[6]), .C(modrm[7]), .D(n_2505), .Z(n_1901
		));
	notech_and2 i_989(.A(modrm[6]), .B(modrm[7]), .Z(n_1900));
	notech_or4 i_975(.A(n_2412), .B(n_58591), .C(n_58481), .D(n_58417), .Z(n_1896
		));
	notech_or4 i_968(.A(n_2458), .B(n_58591), .C(n_58481), .D(n_58417), .Z(n_1895
		));
	notech_or4 i_956(.A(n_2313), .B(n_58363), .C(n_2280), .D(n_2387), .Z(n_1892
		));
	notech_or2 i_946(.A(n_3935), .B(n_3963), .Z(n_1890));
	notech_and4 i_940(.A(n_2027), .B(n_2387), .C(n_30702), .D(n_2413), .Z(n_1888
		));
	notech_or4 i_938(.A(modrm[1]), .B(n_2553), .C(n_30847), .D(n_2495), .Z(n_1887
		));
	notech_or4 i_937(.A(modrm[1]), .B(n_2553), .C(modrm[0]), .D(n_2492), .Z(n_1886
		));
	notech_mux2 i_321(.S(modrm[0]), .A(n_1882), .B(n_2037), .Z(n_1885));
	notech_nand3 i_322(.A(n_2372), .B(n_2315), .C(n_2037), .Z(n_1882));
	notech_nand2 i_932(.A(n_2037), .B(modrm[0]), .Z(n_1879));
	notech_or4 i_922(.A(n_2300), .B(n_2455), .C(n_58597), .D(n_58591), .Z(n_1877
		));
	notech_or4 i_913(.A(n_2360), .B(n_58492), .C(n_30738), .D(n_58372), .Z(n_1875
		));
	notech_or4 i_898(.A(modrm[1]), .B(n_2553), .C(modrm[0]), .D(n_2372), .Z(n_1874
		));
	notech_or4 i_897(.A(modrm[1]), .B(n_2553), .C(n_2315), .D(n_30847), .Z(n_1873
		));
	notech_mux2 i_312(.S(modrm[0]), .A(n_2373), .B(n_2037), .Z(n_1872));
	notech_or4 i_894(.A(n_2497), .B(n_2333), .C(n_1872), .D(n_30848), .Z(n_1871
		));
	notech_or4 i_893(.A(n_2485), .B(n_2372), .C(n_2490), .D(modrm[0]), .Z(n_1869
		));
	notech_ao4 i_881(.A(n_2333), .B(n_2288), .C(n_2486), .D(n_2295), .Z(n_1858
		));
	notech_or4 i_875(.A(n_2383), .B(n_2333), .C(n_2290), .D(n_2300), .Z(n_1857
		));
	notech_nao3 i_870(.A(n_58519), .B(n_2530), .C(n_2300), .Z(n_1855));
	notech_nao3 i_869(.A(n_58528), .B(n_2536), .C(n_2292), .Z(n_1854));
	notech_or4 i_825(.A(n_58381), .B(n_2302), .C(n_3963), .D(n_58426), .Z(n_1851
		));
	notech_or4 i_954(.A(n_2475), .B(n_2445), .C(n_1849), .D(n_1838), .Z(\udeco[126] 
		));
	notech_and2 i_752(.A(modrm[2]), .B(n_30826), .Z(n_1849));
	notech_nand2 i_741(.A(n_1943), .B(n_30795), .Z(n_1848));
	notech_and4 i_743(.A(n_58399), .B(n_1944), .C(n_2296), .D(n_2427), .Z(n_1846
		));
	notech_or2 i_740(.A(n_2433), .B(n_58591), .Z(n_1843));
	notech_and2 i_69(.A(n_2032), .B(n_3733), .Z(n_1842));
	notech_and4 i_81(.A(n_1837), .B(n_2417), .C(n_2415), .D(n_2406), .Z(n_1841
		));
	notech_and4 i_82(.A(n_2352), .B(n_2344), .C(n_1905), .D(n_1825), .Z(n_1840
		));
	notech_and2 i_749(.A(n_58426), .B(n_30827), .Z(n_1838));
	notech_or4 i_735(.A(n_58492), .B(n_2316), .C(n_30738), .D(n_2387), .Z(n_1837
		));
	notech_nand3 i_734(.A(n_58577), .B(n_2272), .C(n_30790), .Z(n_1835));
	notech_or4 i_731(.A(n_2276), .B(n_2407), .C(n_58514), .D(n_58528), .Z(n_1833
		));
	notech_or4 i_673(.A(n_2299), .B(n_3963), .C(n_58546), .D(n_30806), .Z(n_1831
		));
	notech_or4 i_718(.A(n_2393), .B(n_58481), .C(n_58465), .D(n_58399), .Z(n_1829
		));
	notech_or4 i_717(.A(n_2313), .B(n_58363), .C(n_2280), .D(n_2299), .Z(n_1828
		));
	notech_nao3 i_851(.A(n_58577), .B(n_2272), .C(n_4072), .Z(n_1825));
	notech_or2 i_656(.A(n_2303), .B(n_2285), .Z(n_1824));
	notech_and3 i_340(.A(n_2278), .B(n_2293), .C(n_30702), .Z(n_1822));
	notech_or2 i_652(.A(n_2285), .B(n_1822), .Z(n_1821));
	notech_or2 i_651(.A(n_2285), .B(n_2027), .Z(n_1820));
	notech_and2 i_647(.A(n_2295), .B(n_2302), .Z(n_1819));
	notech_and2 i_286(.A(n_2297), .B(n_30801), .Z(n_1818));
	notech_or4 i_621(.A(n_2348), .B(n_58408), .C(n_58363), .D(n_1818), .Z(n_1817
		));
	notech_or4 i_620(.A(n_2348), .B(n_58408), .C(n_58363), .D(n_2299), .Z(n_1813
		));
	notech_and4 i_615(.A(n_2278), .B(n_2275), .C(n_2302), .D(n_30702), .Z(n_1812
		));
	notech_ao3 i_531(.A(n_58546), .B(n_2324), .C(n_2330), .Z(n_1807));
	notech_or4 i_529(.A(n_58354), .B(n_2185), .C(n_58481), .D(n_58465), .Z(n_1806
		));
	notech_or4 i_502(.A(n_58492), .B(n_58381), .C(n_2297), .D(n_58514), .Z(n_1805
		));
	notech_and2 i_463(.A(n_2289), .B(n_2290), .Z(n_1802));
	notech_or2 i_23111435(.A(n_2337), .B(n_30702), .Z(n_1801));
	notech_or4 i_184(.A(n_2488), .B(n_30849), .C(n_30850), .D(n_30847), .Z(n_1800
		));
	notech_nand3 i_145(.A(n_58399), .B(n_2530), .C(n_58528), .Z(n_1798));
	notech_or4 i_839(.A(n_2313), .B(n_58363), .C(n_2280), .D(n_2290), .Z(n_1797
		));
	notech_or4 i_855(.A(n_2292), .B(n_2455), .C(n_58597), .D(n_58591), .Z(n_1796
		));
	notech_ao3 i_1104(.A(n_30790), .B(n_2321), .C(n_2101), .Z(n_1795));
	notech_or4 i_1225(.A(adz), .B(n_58555), .C(n_2347), .D(n_1916), .Z(n_1794
		));
	notech_or4 i_1291(.A(n_58492), .B(n_2448), .C(n_58510), .D(n_58528), .Z(n_1793
		));
	notech_or4 i_1233(.A(n_2347), .B(n_2284), .C(n_2018), .D(n_58555), .Z(n_1792
		));
	notech_nand3 i_520(.A(n_2278), .B(n_2299), .C(n_3761), .Z(n_1791));
	notech_and4 i_78572358(.A(n_1778), .B(n_3280), .C(n_3109), .D(n_1785), .Z
		(n_1789));
	notech_and4 i_78172362(.A(n_1950), .B(n_1638), .C(n_738), .D(n_3994), .Z
		(n_1785));
	notech_and4 i_78072363(.A(n_811), .B(n_3098), .C(n_2579), .D(n_3079), .Z
		(n_1778));
	notech_and4 i_11573087(.A(n_2571), .B(n_4013), .C(n_2394), .D(n_2365), .Z
		(n_1770));
	notech_and4 i_67372444(.A(n_1741), .B(n_1738), .C(n_176192234), .D(n_30728
		), .Z(n_1762));
	notech_and4 i_67072445(.A(n_1745), .B(n_1744), .C(n_1759), .D(n_1702), .Z
		(n_176192234));
	notech_and4 i_66872447(.A(n_3993), .B(n_1757), .C(n_2305), .D(n_1751), .Z
		(n_1759));
	notech_and4 i_66072454(.A(n_1793), .B(n_2894), .C(n_2136), .D(n_3152), .Z
		(n_1757));
	notech_and4 i_65972455(.A(n_2609), .B(n_2928), .C(n_1792), .D(n_2629), .Z
		(n_1751));
	notech_ao4 i_65872456(.A(n_30792), .B(n_58519), .C(n_30791), .D(n_4072),
		 .Z(n_1745));
	notech_ao4 i_65672457(.A(n_30794), .B(n_1802), .C(n_2124), .D(n_58537), 
		.Z(n_1744));
	notech_and4 i_66272452(.A(n_30836), .B(n_69848720), .C(n_30679), .D(n_2365
		), .Z(n_1741));
	notech_and4 i_66172453(.A(n_4056), .B(n_4036), .C(n_872), .D(n_30719), .Z
		(n_1738));
	notech_and3 i_31373069(.A(n_4014), .B(n_208149924), .C(n_30698), .Z(n_1734
		));
	notech_and4 i_46572613(.A(n_2894), .B(n_4055), .C(n_1725), .D(n_1699), .Z
		(n_1730));
	notech_and4 i_46072617(.A(n_4030), .B(n_2569), .C(n_1950), .D(n_30692), 
		.Z(n_1725));
	notech_nand3 i_25473074(.A(n_2076), .B(n_4055), .C(n_2620), .Z(n_1722)
		);
	notech_ao3 i_46472614(.A(n_1719), .B(n_1714), .C(n_1640), .Z(n_1721));
	notech_and4 i_45972618(.A(n_4031), .B(n_1014), .C(n_3993), .D(n_30720), 
		.Z(n_1719));
	notech_and4 i_45872619(.A(n_4026), .B(n_2760), .C(n_2479), .D(n_2690), .Z
		(n_1714));
	notech_and4 i_31273071(.A(n_4007), .B(n_4047), .C(n_2340), .D(n_2609), .Z
		(n_1709));
	notech_and4 i_11673086(.A(n_4086), .B(n_2538), .C(n_30722), .D(n_1704), 
		.Z(n_1708));
	notech_and3 i_8173089(.A(n_4002), .B(n_4076), .C(n_4027), .Z(n_1704));
	notech_and4 i_73573039(.A(n_30712), .B(n_1958), .C(n_2377), .D(n_30691),
		 .Z(n_1702));
	notech_and2 i_62273051(.A(n_2365), .B(n_30689), .Z(n_1699));
	notech_and4 i_13972901(.A(n_1801), .B(n_3402), .C(n_1694), .D(n_4093), .Z
		(n_1695));
	notech_and4 i_13772903(.A(n_2664), .B(n_2637), .C(n_2357), .D(n_3124), .Z
		(n_1694));
	notech_or4 i_13872902(.A(n_1795), .B(n_4024), .C(n_1626), .D(n_1625), .Z
		(n_1689));
	notech_and4 i_12572915(.A(n_2611), .B(n_2949), .C(n_2166), .D(n_2463), .Z
		(n_1684));
	notech_and4 i_12672914(.A(n_3013), .B(n_2480), .C(n_2729), .D(n_2959), .Z
		(n_1681));
	notech_ao3 i_8772946(.A(n_2743), .B(n_2623), .C(n_1675), .Z(n_1676));
	notech_nand3 i_32673067(.A(n_2019), .B(n_1616), .C(n_1618), .Z(n_1675)
		);
	notech_and4 i_8572948(.A(n_1671), .B(n_1668), .C(n_1664), .D(n_1661), .Z
		(n_1673));
	notech_and4 i_8072951(.A(n_247292237), .B(n_2045), .C(n_2591), .D(n_4030
		), .Z(n_1671));
	notech_and4 i_7972952(.A(n_2588), .B(n_3360), .C(n_2627), .D(n_30680), .Z
		(n_1668));
	notech_and4 i_7872953(.A(n_2744), .B(n_2140), .C(n_2516), .D(n_1942), .Z
		(n_1664));
	notech_ao3 i_7772954(.A(n_30664), .B(n_1619), .C(n_30813), .Z(n_1661));
	notech_and4 i_5972970(.A(n_4048), .B(n_164992233), .C(n_2036), .D(n_1653
		), .Z(n_1654));
	notech_and4 i_5772972(.A(n_30836), .B(n_2831), .C(n_2450), .D(n_2426), .Z
		(n_1653));
	notech_and2 i_5072978(.A(n_2398), .B(n_1834), .Z(n_164992233));
	notech_and4 i_5872971(.A(n_1644), .B(n_2305), .C(n_1612), .D(n_3984), .Z
		(n_1647));
	notech_ao4 i_5372975(.A(n_2166), .B(n_2006), .C(n_4071), .D(n_1965), .Z(n_1644
		));
	notech_nand3 i_52373060(.A(n_4025), .B(n_2629), .C(n_30723), .Z(n_1640)
		);
	notech_and4 i_50273113(.A(n_1770), .B(n_1789), .C(n_1709), .D(n_3197), .Z
		(n_1639));
	notech_or2 i_77372368(.A(n_2151), .B(n_58465), .Z(n_1638));
	notech_or2 i_71172419(.A(n_3958), .B(n_2359), .Z(n_1637));
	notech_nand3 i_55373118(.A(n_1762), .B(n_1734), .C(n_1629), .Z(\udeco[33] 
		));
	notech_nand2 i_64472465(.A(modrm[4]), .B(n_221894218), .Z(n_1629));
	notech_and4 i_60373126(.A(n_1730), .B(n_1709), .C(n_1708), .D(n_1721), .Z
		(n_1628));
	notech_or4 i_77673155(.A(n_1689), .B(n_1621), .C(n_30832), .D(n_2102), .Z
		(\udeco[110] ));
	notech_and2 i_12972911(.A(adz), .B(n_30823), .Z(n_1626));
	notech_and2 i_12872912(.A(adz), .B(n_30718), .Z(n_1625));
	notech_and4 i_373025(.A(n_2484), .B(n_1684), .C(n_1681), .D(n_1995), .Z(n_1622
		));
	notech_and2 i_13072910(.A(opz[2]), .B(n_30857), .Z(n_1621));
	notech_and4 i_91573158(.A(n_1676), .B(n_1673), .C(n_30681), .D(n_2435), 
		.Z(n_1620));
	notech_or4 i_6872962(.A(n_2289), .B(n_58381), .C(n_58399), .D(n_30785), 
		.Z(n_1619));
	notech_or4 i_6572965(.A(n_2311), .B(n_58481), .C(n_58465), .D(n_30785), 
		.Z(n_1618));
	notech_nao3 i_6672964(.A(n_58481), .B(n_58591), .C(n_3277), .Z(n_1616)
		);
	notech_and4 i_94373159(.A(n_1654), .B(n_1647), .C(n_1613), .D(n_1606), .Z
		(n_1614));
	notech_nand2 i_4772981(.A(modrm[1]), .B(n_30858), .Z(n_1613));
	notech_or2 i_4572983(.A(n_4070), .B(n_58519), .Z(n_1612));
	notech_and4 i_073028(.A(n_4034), .B(n_1865), .C(n_1604), .D(n_2883), .Z(n_1608
		));
	notech_nand3 i_63882(.A(n_2398), .B(n_2380), .C(n_30685), .Z(\udeco[4] )
		);
	notech_and4 i_64115(.A(n_2366), .B(n_1960), .C(n_30722), .D(n_122993389)
		, .Z(udeco_73100251));
	notech_and2 i_1073018(.A(modrm[4]), .B(n_30742), .Z(n_118493346));
	notech_or4 i_64146(.A(n_4024), .B(n_214994159), .C(n_3971), .D(n_118493346
		), .Z(\udeco[84] ));
	notech_and2 i_1373015(.A(n_58426), .B(n_30742), .Z(n_118593347));
	notech_or4 i_64151(.A(n_3971), .B(n_4045), .C(n_118593347), .D(n_123493393
		), .Z(\udeco[85] ));
	notech_nao3 i_10373100(.A(n_1960), .B(n_3998), .C(n_4057), .Z(\udeco[88] 
		));
	notech_or2 i_64163(.A(\udeco[88] ), .B(\udeco[5] ), .Z(\udeco[89] ));
	notech_or4 i_6973099(.A(n_30781), .B(\udeco[5] ), .C(n_30757), .D(n_3971
		), .Z(\udeco[91] ));
	notech_nao3 i_64166(.A(n_30696), .B(n_30724), .C(n_30788), .Z(\udeco[92] 
		));
	notech_nao3 i_11373098(.A(n_3998), .B(n_30696), .C(n_30788), .Z(\udeco[90] 
		));
	notech_or2 i_64168(.A(n_4057), .B(\udeco[90] ), .Z(\udeco[93] ));
	notech_or2 i_64169(.A(n_4057), .B(\udeco[91] ), .Z(\udeco[95] ));
	notech_nao3 i_64170(.A(n_3998), .B(n_1960), .C(n_4010), .Z(\udeco[96] )
		);
	notech_or2 i_64172(.A(n_4010), .B(\udeco[88] ), .Z(\udeco[98] ));
	notech_or4 i_64174(.A(n_4024), .B(n_4057), .C(n_3971), .D(n_3985), .Z(\udeco[100] 
		));
	notech_and4 i_64175(.A(n_30797), .B(n_2623), .C(n_1960), .D(n_30724), .Z
		(udeco_101100250));
	notech_or4 i_64176(.A(n_4018), .B(n_3950), .C(\udeco[88] ), .D(n_4010), 
		.Z(\udeco[102] ));
	notech_nao3 i_28673160(.A(n_30859), .B(n_124593404), .C(n_124093399), .Z
		(\udeco[127] ));
	notech_nand3 i_273026(.A(n_2099), .B(n_3736), .C(n_1905), .Z(n_118693348
		));
	notech_nor2 i_9072943(.A(n_1984), .B(n_30842), .Z(n_118793349));
	notech_nand2 i_9172942(.A(n_58426), .B(n_3956), .Z(n_118893350));
	notech_and2 i_9272941(.A(modrm[2]), .B(n_118693348), .Z(n_118993351));
	notech_or4 i_88073157(.A(n_124093399), .B(n_126193417), .C(n_125493411),
		 .D(n_125193408), .Z(\udeco[118] ));
	notech_or4 i_69873156(.A(n_4024), .B(n_4057), .C(n_1675), .D(n_30734), .Z
		(\udeco[115] ));
	notech_or4 i_56173154(.A(n_128793438), .B(n_30737), .C(n_127393426), .D(n_207949923
		), .Z(\udeco[107] ));
	notech_nao3 i_16272881(.A(n_58591), .B(n_2397), .C(n_2403), .Z(n_119093352
		));
	notech_or4 i_16472880(.A(n_58354), .B(n_4090), .C(n_2315), .D(modrm[5]),
		 .Z(n_119193353));
	notech_nand2 i_16872877(.A(opz[2]), .B(n_30708), .Z(n_119293354));
	notech_nand3 i_20273153(.A(n_119193353), .B(n_119093352), .C(n_129793447
		), .Z(\udeco[106] ));
	notech_or2 i_17872869(.A(n_2278), .B(n_2052), .Z(n_119493355));
	notech_nand2 i_17972868(.A(opz[1]), .B(n_30708), .Z(n_119593356));
	notech_nand3 i_72573152(.A(n_119193353), .B(n_130993454), .C(n_119093352
		), .Z(\udeco[105] ));
	notech_and4 i_20573151(.A(n_1969), .B(n_2623), .C(n_1960), .D(n_30797), 
		.Z(udeco_103100249));
	notech_and2 i_19272855(.A(modrm[7]), .B(n_30742), .Z(n_119693357));
	notech_or4 i_72173150(.A(n_30788), .B(n_214994159), .C(n_3971), .D(n_119693357
		), .Z(\udeco[87] ));
	notech_and2 i_19572852(.A(modrm[6]), .B(n_30742), .Z(n_119793358));
	notech_or4 i_72110268(.A(n_30788), .B(n_214994159), .C(n_3971), .D(n_119793358
		), .Z(\udeco[86] ));
	notech_or4 i_64173(.A(n_4024), .B(n_4057), .C(n_4010), .D(n_3971), .Z(\udeco[99] 
		));
	notech_nand2 i_19972848(.A(modrm[3]), .B(n_30742), .Z(n_119893359));
	notech_or4 i_71873149(.A(n_214994159), .B(n_4009), .C(\udeco[99] ), .D(n_131593460
		), .Z(\udeco[83] ));
	notech_nand2 i_21172841(.A(modrm[2]), .B(n_30742), .Z(n_120193362));
	notech_nand3 i_71573148(.A(n_131893463), .B(n_131793462), .C(n_132293465
		), .Z(\udeco[82] ));
	notech_or4 i_21772835(.A(n_2386), .B(n_58372), .C(n_58537), .D(n_30729),
		 .Z(n_120293363));
	notech_or4 i_22072833(.A(n_58492), .B(n_2182), .C(n_58528), .D(n_58456),
		 .Z(n_120493365));
	notech_and2 i_22172832(.A(modrm[1]), .B(n_30742), .Z(n_120593366));
	notech_or4 i_71273147(.A(n_30835), .B(n_120593366), .C(n_30788), .D(n_133193471
		), .Z(\udeco[81] ));
	notech_or4 i_22273146(.A(n_4011), .B(n_4018), .C(\udeco[91] ), .D(n_30739
		), .Z(\udeco[80] ));
	notech_nao3 i_10473093(.A(n_122993389), .B(n_1960), .C(n_133793475), .Z(\udeco[74] 
		));
	notech_or4 i_21610271(.A(n_30684), .B(n_30683), .C(\udeco[74] ), .D(n_3968
		), .Z(\udeco[78] ));
	notech_nao3 i_20510274(.A(n_30726), .B(n_30859), .C(n_133893476), .Z(\udeco[77] 
		));
	notech_or4 i_22873145(.A(n_133893476), .B(n_1326), .C(n_3971), .D(n_3978
		), .Z(\udeco[75] ));
	notech_nand3 i_22210283(.A(n_131793462), .B(n_135393486), .C(n_122993389
		), .Z(\udeco[72] ));
	notech_or4 i_70973144(.A(n_124093399), .B(n_136293494), .C(n_30683), .D(n_3969
		), .Z(\udeco[70] ));
	notech_nao3 i_11473092(.A(n_30709), .B(n_30691), .C(n_136293494), .Z(\udeco[71] 
		));
	notech_or4 i_70573143(.A(n_4009), .B(n_3969), .C(n_136293494), .D(n_3968
		), .Z(\udeco[68] ));
	notech_or4 i_20973142(.A(n_30683), .B(\udeco[71] ), .C(\udeco[5] ), .D(n_214994159
		), .Z(\udeco[67] ));
	notech_or4 i_20210290(.A(n_4045), .B(n_136293494), .C(n_136393495), .D(n_30684
		), .Z(\udeco[69] ));
	notech_or2 i_70273141(.A(n_4057), .B(\udeco[69] ), .Z(\udeco[66] ));
	notech_or4 i_69810294(.A(n_135693488), .B(n_30762), .C(n_136093492), .D(n_137393504
		), .Z(\udeco[65] ));
	notech_or4 i_69810298(.A(n_135693488), .B(n_30762), .C(n_136093492), .D(n_137793508
		), .Z(\udeco[64] ));
	notech_or4 i_69473140(.A(n_4054), .B(n_139393521), .C(n_4015), .D(n_138993517
		), .Z(\udeco[63] ));
	notech_or4 i_68373139(.A(n_121193371), .B(n_139393521), .C(n_124093399),
		 .D(n_138993517), .Z(\udeco[62] ));
	notech_nao3 i_68973138(.A(n_140093528), .B(n_30741), .C(n_124093399), .Z
		(\udeco[61] ));
	notech_or4 i_59273137(.A(n_140593532), .B(n_140293530), .C(n_4015), .D(n_4054
		), .Z(\udeco[60] ));
	notech_nand3 i_68310303(.A(n_138493512), .B(n_141293539), .C(n_30740), .Z
		(\udeco[59] ));
	notech_nand3 i_67873136(.A(n_2579), .B(n_138493512), .C(n_142393548), .Z
		(\udeco[58] ));
	notech_or4 i_67273135(.A(n_135893490), .B(n_135793489), .C(n_140293530),
		 .D(n_142693550), .Z(\udeco[57] ));
	notech_ao4 i_105873031(.A(n_2210), .B(n_3959), .C(n_30793), .D(n_30656),
		 .Z(n_121193371));
	notech_or4 i_66773134(.A(n_142993553), .B(n_121193371), .C(n_143293556),
		 .D(n_140293530), .Z(\udeco[56] ));
	notech_or4 i_66210308(.A(n_144193564), .B(n_4011), .C(n_1640), .D(n_30825
		), .Z(\udeco[55] ));
	notech_nao3 i_65773133(.A(n_143893561), .B(n_144893571), .C(n_124093399)
		, .Z(\udeco[54] ));
	notech_or4 i_65273132(.A(n_30746), .B(n_146193583), .C(n_221894218), .D(n_30762
		), .Z(\udeco[53] ));
	notech_or4 i_64573131(.A(n_146493586), .B(n_30825), .C(n_30745), .D(n_122893388
		), .Z(\udeco[52] ));
	notech_or4 i_64173130(.A(n_135893490), .B(n_135793489), .C(n_30825), .D(n_148393599
		), .Z(\udeco[51] ));
	notech_ao3 i_39472679(.A(n_30850), .B(modrm[3]), .C(n_2113), .Z(n_121293372
		));
	notech_or4 i_63573129(.A(n_30762), .B(n_30746), .C(n_124093399), .D(n_149993613
		), .Z(\udeco[50] ));
	notech_or4 i_41172662(.A(n_2118), .B(n_58597), .C(n_58465), .D(n_58417),
		 .Z(n_121393373));
	notech_nao3 i_61973128(.A(n_150993622), .B(n_143893561), .C(n_30825), .Z
		(\udeco[48] ));
	notech_or4 i_62373127(.A(n_152493637), .B(n_151293625), .C(n_139193519),
		 .D(n_30730), .Z(\udeco[47] ));
	notech_or4 i_61910312(.A(n_1640), .B(n_30751), .C(n_152793639), .D(n_153693647
		), .Z(\udeco[46] ));
	notech_or4 i_61573125(.A(n_155193657), .B(n_151793630), .C(n_154993655),
		 .D(n_30730), .Z(\udeco[44] ));
	notech_or4 i_35373124(.A(n_221894218), .B(n_30727), .C(n_30756), .D(n_157293675
		), .Z(\udeco[43] ));
	notech_or2 i_49872580(.A(n_5254), .B(n_58390), .Z(n_121493374));
	notech_or4 i_60973123(.A(n_30756), .B(n_157493677), .C(n_159193691), .D(n_30731
		), .Z(\udeco[42] ));
	notech_or4 i_60310319(.A(n_30825), .B(n_151793630), .C(n_161093706), .D(n_135993491
		), .Z(\udeco[41] ));
	notech_ao4 i_473024(.A(n_4065), .B(n_2320), .C(n_58363), .D(n_2371), .Z(n_121893378
		));
	notech_nor2 i_54372542(.A(n_5254), .B(n_30849), .Z(n_121993379));
	notech_nor2 i_54472541(.A(n_2275), .B(n_121893378), .Z(n_122093380));
	notech_or4 i_59673122(.A(n_161693711), .B(n_162593717), .C(n_152793639),
		 .D(n_151293625), .Z(\udeco[40] ));
	notech_nand3 i_59210324(.A(n_163993728), .B(n_163693725), .C(n_163293722
		), .Z(\udeco[39] ));
	notech_or4 i_58773121(.A(n_164893737), .B(n_164593734), .C(n_155193657),
		 .D(n_30761), .Z(\udeco[38] ));
	notech_nao3 i_57573120(.A(n_1734), .B(n_166593751), .C(n_221894218), .Z(\udeco[36] 
		));
	notech_nao3 i_61072488(.A(n_58399), .B(n_58591), .C(n_2564), .Z(n_122193381
		));
	notech_and4 i_56873119(.A(n_1193), .B(n_168393768), .C(n_167593761), .D(n_1734
		), .Z(udeco_35100248));
	notech_nand3 i_53973117(.A(n_170793789), .B(n_169193776), .C(n_1960), .Z
		(\udeco[31] ));
	notech_or4 i_53173116(.A(n_221894218), .B(n_30774), .C(n_204849898), .D(n_172793805
		), .Z(\udeco[30] ));
	notech_and4 i_52273115(.A(n_169093775), .B(n_1770), .C(n_174393818), .D(n_3109
		), .Z(udeco_29100247));
	notech_and4 i_51273114(.A(n_175093824), .B(n_176293834), .C(n_3510), .D(n_169193776
		), .Z(udeco_28100246));
	notech_or4 i_78872355(.A(n_2347), .B(n_2338), .C(n_3961), .D(n_58555), .Z
		(n_122293382));
	notech_nao3 i_46173112(.A(n_179193853), .B(n_1699), .C(n_30770), .Z(\udeco[22] 
		));
	notech_and4 i_45173111(.A(n_179493856), .B(n_182093879), .C(n_1925), .D(n_222294221
		), .Z(udeco_21100245));
	notech_or4 i_42473110(.A(n_30774), .B(n_30825), .C(n_30773), .D(n_184393897
		), .Z(\udeco[19] ));
	notech_and4 i_37273109(.A(n_185993912), .B(n_185593909), .C(n_185393907)
		, .D(n_3403), .Z(udeco_15100244));
	notech_and4 i_36973108(.A(n_187293922), .B(n_186793919), .C(n_151893631)
		, .D(n_3403), .Z(udeco_14100243));
	notech_nor2 i_88672262(.A(n_3954), .B(n_3958), .Z(n_122393383));
	notech_and4 i_35310362(.A(n_188093930), .B(n_187793927), .C(n_189293942)
		, .D(n_30698), .Z(udeco_12100242));
	notech_nand2 i_29510367(.A(n_68), .B(n_30782), .Z(\udeco[6] ));
	notech_or2 i_91272236(.A(n_2398), .B(n_58465), .Z(n_122493384));
	notech_nand3 i_29073107(.A(n_122493384), .B(n_30706), .C(n_30782), .Z(\udeco[3] 
		));
	notech_nor2 i_91672233(.A(n_2398), .B(n_58456), .Z(n_122593385));
	notech_or4 i_29010371(.A(n_1967), .B(n_30783), .C(n_122593385), .D(n_189793947
		), .Z(\udeco[2] ));
	notech_nor2 i_92072229(.A(n_2398), .B(n_58519), .Z(n_122693386));
	notech_or4 i_28610376(.A(n_190093949), .B(n_4006), .C(n_122693386), .D(n_30784
		), .Z(\udeco[1] ));
	notech_nand2 i_35473066(.A(n_1958), .B(n_4066), .Z(n_122893388));
	notech_and3 i_68673046(.A(n_3992), .B(n_3876), .C(n_30732), .Z(n_122993389
		));
	notech_nao3 i_1573013(.A(n_1950), .B(n_2380), .C(n_214994159), .Z(n_123493393
		));
	notech_nao3 i_6373090(.A(n_30709), .B(n_30707), .C(n_1640), .Z(n_124093399
		));
	notech_and4 i_3472994(.A(n_4017), .B(n_1920), .C(n_2450), .D(n_30725), .Z
		(n_124393402));
	notech_and4 i_3672992(.A(n_4048), .B(n_2195), .C(n_124393402), .D(n_2435
		), .Z(n_124593404));
	notech_or4 i_10072933(.A(n_30750), .B(n_4003), .C(n_1180), .D(n_3985), .Z
		(n_125193408));
	notech_or4 i_10172932(.A(n_222594224), .B(n_30818), .C(n_30822), .D(n_4080
		), .Z(n_125493411));
	notech_and4 i_9972934(.A(n_2516), .B(n_3733), .C(n_2332), .D(n_118893350
		), .Z(n_125893415));
	notech_or4 i_10672929(.A(n_118793349), .B(n_118993351), .C(n_3974), .D(n_30733
		), .Z(n_126193417));
	notech_and4 i_11272923(.A(n_1543), .B(n_1923), .C(n_4061), .D(n_1545), .Z
		(n_126993422));
	notech_or4 i_15272889(.A(n_222994228), .B(n_30735), .C(n_1262), .D(n_30736
		), .Z(n_127393426));
	notech_and4 i_15372888(.A(n_4084), .B(n_3991), .C(n_2162), .D(n_4004), .Z
		(n_127693429));
	notech_nand2 i_14472896(.A(n_4061), .B(n_2792), .Z(n_128193434));
	notech_or4 i_15472887(.A(n_4024), .B(n_30710), .C(n_30697), .D(n_128193434
		), .Z(n_128393436));
	notech_or4 i_16072883(.A(n_30828), .B(n_4009), .C(n_128393436), .D(n_30770
		), .Z(n_128793438));
	notech_and4 i_17572872(.A(n_1678), .B(n_208394100), .C(n_2623), .D(n_30724
		), .Z(n_129693446));
	notech_and4 i_17672871(.A(n_129693446), .B(n_30709), .C(n_4087), .D(n_119293354
		), .Z(n_129793447));
	notech_and4 i_18572862(.A(n_4043), .B(n_4087), .C(n_1678), .D(n_208394100
		), .Z(n_130193449));
	notech_and3 i_18472863(.A(n_2049), .B(n_3998), .C(n_119593356), .Z(n_130793452
		));
	notech_and4 i_18772860(.A(n_119493355), .B(n_130793452), .C(n_130193449)
		, .D(n_2380), .Z(n_130993454));
	notech_nao3 i_20472846(.A(n_4093), .B(n_119893359), .C(n_30684), .Z(n_131593460
		));
	notech_and2 i_69173043(.A(n_2366), .B(n_30856), .Z(n_131793462));
	notech_ao4 i_21372839(.A(n_2383), .B(n_2167), .C(n_3963), .D(n_2182), .Z
		(n_131893463));
	notech_and4 i_21472838(.A(n_30726), .B(n_30722), .C(n_2357), .D(n_120193362
		), .Z(n_132293465));
	notech_ao4 i_22572829(.A(n_2383), .B(n_2182), .C(n_2167), .D(n_30785), .Z
		(n_133093470));
	notech_nand3 i_22772827(.A(n_120293363), .B(n_133093470), .C(n_30722), .Z
		(n_133193471));
	notech_ao4 i_23372823(.A(n_1953), .B(n_30847), .C(n_2577), .D(n_3935), .Z
		(n_133493473));
	notech_nao3 i_80373033(.A(n_2629), .B(n_1953), .C(n_4011), .Z(n_133793475
		));
	notech_nao3 i_16973080(.A(n_5254), .B(n_30732), .C(n_133793475), .Z(n_133893476
		));
	notech_and3 i_25072806(.A(n_3970), .B(n_120493365), .C(n_30792), .Z(n_134993482
		));
	notech_ao4 i_24972807(.A(n_30729), .B(n_2167), .C(n_58354), .D(n_2368), 
		.Z(n_135193484));
	notech_and4 i_25272804(.A(n_135193484), .B(n_2151), .C(n_30829), .D(n_134993482
		), .Z(n_135393486));
	notech_nand2 i_55173058(.A(n_2123), .B(n_4034), .Z(n_135693488));
	notech_or2 i_80573032(.A(n_135693488), .B(n_30762), .Z(n_135793489));
	notech_or2 i_25772801(.A(n_30717), .B(n_4024), .Z(n_135893490));
	notech_or4 i_15673083(.A(n_4024), .B(n_30717), .C(n_135693488), .D(n_30762
		), .Z(n_135993491));
	notech_nand3 i_64273049(.A(n_4056), .B(n_4044), .C(n_3964), .Z(n_136093492
		));
	notech_or4 i_235573029(.A(n_4091), .B(n_136093492), .C(n_135893490), .D(n_135793489
		), .Z(n_136293494));
	notech_or4 i_25972799(.A(n_4011), .B(n_1640), .C(n_4009), .D(n_3969), .Z
		(n_136393495));
	notech_nand3 i_65173047(.A(n_5254), .B(n_2377), .C(n_1958), .Z(n_136893500
		));
	notech_or2 i_73073041(.A(n_30717), .B(n_30757), .Z(n_136993501));
	notech_or4 i_27272787(.A(n_30781), .B(n_3978), .C(n_136993501), .D(n_136893500
		), .Z(n_137393504));
	notech_or4 i_27772782(.A(n_30781), .B(n_4091), .C(n_136993501), .D(n_133793475
		), .Z(n_137793508));
	notech_and4 i_8273088(.A(n_2094), .B(n_210394118), .C(n_2569), .D(n_1905
		), .Z(n_138493512));
	notech_and4 i_28572775(.A(n_3979), .B(n_30725), .C(n_30691), .D(n_1978),
		 .Z(n_138793515));
	notech_nand3 i_11773085(.A(n_138493512), .B(n_138793515), .C(n_1193), .Z
		(n_138993517));
	notech_and2 i_62073053(.A(n_30693), .B(n_30688), .Z(n_139093518));
	notech_or2 i_59773056(.A(n_4006), .B(n_4024), .Z(n_139193519));
	notech_or4 i_28872773(.A(n_4024), .B(n_4006), .C(n_4091), .D(n_30752), .Z
		(n_139393521));
	notech_and4 i_29772765(.A(n_2327), .B(n_2623), .C(n_30692), .D(n_2305), 
		.Z(n_139793525));
	notech_and4 i_30072762(.A(n_139793525), .B(n_131793462), .C(n_139093518)
		, .D(n_30740), .Z(n_140093528));
	notech_nand2 i_62173052(.A(n_2579), .B(n_138493512), .Z(n_140293530));
	notech_or4 i_30472758(.A(n_4006), .B(n_4091), .C(n_222494223), .D(n_30752
		), .Z(n_140593532));
	notech_and4 i_31172751(.A(n_1978), .B(n_30836), .C(n_2304), .D(n_1816), 
		.Z(n_141193538));
	notech_and4 i_31472750(.A(n_141193538), .B(n_1953), .C(n_2623), .D(n_30693
		), .Z(n_141293539));
	notech_and3 i_81473030(.A(n_30695), .B(n_30688), .C(n_2380), .Z(n_141593542
		));
	notech_and4 i_32172743(.A(n_139793525), .B(n_30836), .C(n_2357), .D(n_30743
		), .Z(n_142193546));
	notech_and4 i_32572740(.A(n_30740), .B(n_1193), .C(n_141593542), .D(n_142193546
		), .Z(n_142393548));
	notech_nao3 i_32972737(.A(n_30692), .B(n_139093518), .C(n_4091), .Z(n_142693550
		));
	notech_nao3 i_33572731(.A(n_1953), .B(n_1950), .C(n_4009), .Z(n_142993553
		));
	notech_or4 i_33672730(.A(n_4091), .B(n_2307), .C(n_30717), .D(n_2165), .Z
		(n_143293556));
	notech_and4 i_32273068(.A(n_4031), .B(n_69848720), .C(n_2304), .D(n_30706
		), .Z(n_143893561));
	notech_or4 i_34472722(.A(n_3986), .B(n_210194116), .C(n_30769), .D(n_30744
		), .Z(n_144193564));
	notech_and4 i_35072716(.A(n_30712), .B(n_30721), .C(n_2365), .D(n_1972),
		 .Z(n_144693569));
	notech_and4 i_35272714(.A(n_30798), .B(n_144693569), .C(n_30732), .D(n_30720
		), .Z(n_144893571));
	notech_nand2 i_35872710(.A(n_222794226), .B(n_4016), .Z(n_145193573));
	notech_and4 i_36472704(.A(n_2365), .B(n_2099), .C(n_2327), .D(n_30721), 
		.Z(n_145593577));
	notech_nao3 i_36772702(.A(n_145593577), .B(n_2380), .C(n_145193573), .Z(n_145693578
		));
	notech_or4 i_36672703(.A(n_4045), .B(n_210194116), .C(n_4091), .D(n_30718
		), .Z(n_145993581));
	notech_or4 i_37072700(.A(n_145993581), .B(n_30828), .C(n_4009), .D(n_145693578
		), .Z(n_146193583));
	notech_or4 i_37872694(.A(n_30830), .B(n_30814), .C(n_30816), .D(n_4024),
		 .Z(n_146493586));
	notech_and4 i_37972693(.A(n_3360), .B(n_2099), .C(n_69848720), .D(n_30691
		), .Z(n_146993589));
	notech_and4 i_38872685(.A(n_222794226), .B(n_1737), .C(n_5254), .D(n_4031
		), .Z(n_147993596));
	notech_and4 i_38972684(.A(n_3982), .B(n_147993596), .C(n_2614), .D(n_30706
		), .Z(n_148193597));
	notech_nand3 i_39172682(.A(n_148193597), .B(n_141593542), .C(n_1702), .Z
		(n_148393599));
	notech_or4 i_39572678(.A(n_4023), .B(n_30815), .C(n_30828), .D(n_3990), 
		.Z(n_148693602));
	notech_or4 i_40472669(.A(n_121293372), .B(n_148693602), .C(n_1326), .D(n_4045
		), .Z(n_148893604));
	notech_or4 i_40372670(.A(n_4091), .B(n_3968), .C(n_4088), .D(n_30748), .Z
		(n_149593610));
	notech_or4 i_40572668(.A(n_209694112), .B(n_4052), .C(n_145193573), .D(n_149593610
		), .Z(n_149793611));
	notech_or4 i_40872665(.A(n_148893604), .B(n_30769), .C(n_149793611), .D(n_135693488
		), .Z(n_149993613));
	notech_and4 i_41772656(.A(n_3979), .B(n_2366), .C(n_30836), .D(n_210094115
		), .Z(n_150393617));
	notech_ao3 i_41672657(.A(n_210494119), .B(n_121393373), .C(n_222394222),
		 .Z(n_150793620));
	notech_and4 i_41972654(.A(n_150393617), .B(n_150793620), .C(n_2380), .D(n_30722
		), .Z(n_150993622));
	notech_nand3 i_25373075(.A(n_843), .B(n_4047), .C(n_4067), .Z(n_151293625
		));
	notech_and4 i_42872646(.A(n_4051), .B(n_4007), .C(n_4025), .D(n_4085), .Z
		(n_151693629));
	notech_nand3 i_17473079(.A(n_3993), .B(n_4055), .C(n_151693629), .Z(n_151793630
		));
	notech_and2 i_73773038(.A(n_30714), .B(n_30699), .Z(n_151893631));
	notech_and4 i_43272642(.A(n_4019), .B(n_1014), .C(n_2116), .D(n_30720), 
		.Z(n_152193634));
	notech_nao3 i_43372641(.A(n_30709), .B(n_152193634), .C(n_4088), .Z(n_152293635
		));
	notech_or4 i_43672638(.A(n_4035), .B(n_151793630), .C(n_4033), .D(n_152293635
		), .Z(n_152493637));
	notech_nand2 i_73873037(.A(n_4085), .B(n_1704), .Z(n_152793639));
	notech_and4 i_44372631(.A(n_3982), .B(n_1623), .C(n_30709), .D(n_30721),
		 .Z(n_153393644));
	notech_and4 i_44472630(.A(n_3064), .B(n_3360), .C(n_153393644), .D(n_30688
		), .Z(n_153493645));
	notech_or2 i_44672628(.A(n_139193519), .B(n_30767), .Z(n_153693647));
	notech_and4 i_47372605(.A(n_2017), .B(n_30699), .C(n_30714), .D(n_3980),
		 .Z(n_154293650));
	notech_and4 i_47472604(.A(n_5254), .B(n_4019), .C(n_3064), .D(n_2304), .Z
		(n_154793653));
	notech_nao3 i_47672602(.A(n_154793653), .B(n_154293650), .C(n_151293625)
		, .Z(n_154993655));
	notech_or4 i_36573065(.A(n_4050), .B(n_4054), .C(n_4059), .D(n_4024), .Z
		(n_155193657));
	notech_or4 i_48772591(.A(n_4023), .B(n_4059), .C(n_30831), .D(n_223094229
		), .Z(n_155893663));
	notech_or4 i_49272586(.A(n_1987), .B(n_30802), .C(n_1722), .D(n_155893663
		), .Z(n_156093665));
	notech_nand3 i_48372595(.A(n_1798), .B(n_1796), .C(n_4025), .Z(n_156393667
		));
	notech_or4 i_48972589(.A(n_2307), .B(n_222394222), .C(n_30815), .D(n_30839
		), .Z(n_156793671));
	notech_or4 i_49172587(.A(n_30830), .B(n_4050), .C(n_156393667), .D(n_156793671
		), .Z(n_156893672));
	notech_or4 i_49572583(.A(n_156093665), .B(n_156893672), .C(n_1086), .D(n_30767
		), .Z(n_157293675));
	notech_or4 i_51072569(.A(n_4035), .B(n_4033), .C(n_30717), .D(n_30757), 
		.Z(n_157493677));
	notech_and4 i_50672573(.A(n_210394118), .B(n_69848720), .C(n_2365), .D(n_3993
		), .Z(n_158393683));
	notech_and4 i_50872571(.A(n_3994), .B(n_3996), .C(n_158393683), .D(n_121493374
		), .Z(n_158493684));
	notech_and4 i_50772572(.A(n_2623), .B(n_30725), .C(n_30726), .D(n_4030),
		 .Z(n_158893688));
	notech_and4 i_51372567(.A(n_158893688), .B(n_141593542), .C(n_2116), .D(n_30709
		), .Z(n_159093690));
	notech_nand3 i_51572565(.A(n_222294221), .B(n_158493684), .C(n_159093690
		), .Z(n_159193691));
	notech_ao4 i_52872554(.A(n_5254), .B(n_30850), .C(n_4065), .D(n_2018), .Z
		(n_159493693));
	notech_and4 i_52972553(.A(n_1728), .B(n_4032), .C(n_4056), .D(n_4082), .Z
		(n_159793696));
	notech_and4 i_53072552(.A(n_2760), .B(n_3064), .C(n_214594156), .D(n_30689
		), .Z(n_160193700));
	notech_and4 i_53272551(.A(n_2569), .B(n_30692), .C(n_222794226), .D(n_4086
		), .Z(n_160693703));
	notech_and4 i_53572548(.A(n_160693703), .B(n_160193700), .C(n_159793696)
		, .D(n_159493693), .Z(n_160893705));
	notech_nand2 i_53672547(.A(n_160893705), .B(n_1704), .Z(n_161093706));
	notech_or4 i_55672531(.A(n_156393667), .B(n_4006), .C(n_30833), .D(n_122093380
		), .Z(n_161693711));
	notech_and4 i_55272534(.A(n_1014), .B(n_1951), .C(n_4007), .D(n_1815), .Z
		(n_162293716));
	notech_or4 i_55572532(.A(n_4001), .B(n_2164), .C(n_121993379), .D(n_30758
		), .Z(n_162593717));
	notech_and4 i_57172519(.A(n_2036), .B(n_2569), .C(n_30691), .D(n_30856),
		 .Z(n_163293722));
	notech_and4 i_56972521(.A(n_1332), .B(n_3967), .C(n_212094132), .D(n_211794130
		), .Z(n_163693725));
	notech_and4 i_57072520(.A(n_2176), .B(n_3979), .C(n_901), .D(n_3965), .Z
		(n_163993728));
	notech_and4 i_58072511(.A(n_2176), .B(n_901), .C(n_894), .D(n_212494135)
		, .Z(n_164493733));
	notech_nand3 i_58272509(.A(n_2036), .B(n_164493733), .C(n_30722), .Z(n_164593734
		));
	notech_or4 i_58172510(.A(n_30822), .B(n_1987), .C(n_30830), .D(n_4060), 
		.Z(n_164893737));
	notech_and4 i_60172495(.A(n_2569), .B(n_2015), .C(n_214594156), .D(n_30693
		), .Z(n_165393741));
	notech_and4 i_59872497(.A(n_1329), .B(n_3977), .C(n_861), .D(n_1537), .Z
		(n_165893744));
	notech_and4 i_59172501(.A(n_2663), .B(n_2327), .C(n_214094151), .D(n_853
		), .Z(n_165993745));
	notech_and4 i_60272494(.A(n_3967), .B(n_3965), .C(n_165993745), .D(n_165893744
		), .Z(n_166293748));
	notech_and4 i_60672491(.A(n_166293748), .B(n_165393741), .C(n_30753), .D
		(n_3107), .Z(n_166593751));
	notech_and4 i_63072475(.A(n_69848720), .B(n_1816), .C(n_30726), .D(n_30721
		), .Z(n_166993755));
	notech_and4 i_62772478(.A(n_222694225), .B(n_4051), .C(n_4029), .D(n_872
		), .Z(n_167393759));
	notech_and4 i_63372472(.A(n_167393759), .B(n_166993755), .C(n_2305), .D(n_122193381
		), .Z(n_167593761));
	notech_and4 i_61472484(.A(n_3062), .B(n_2500), .C(n_3736), .D(n_1905), .Z
		(n_167793763));
	notech_and4 i_62972476(.A(n_3994), .B(n_1593), .C(n_1329), .D(n_30719), 
		.Z(n_168293767));
	notech_and4 i_63272473(.A(n_2076), .B(n_4036), .C(n_167793763), .D(n_168293767
		), .Z(n_168393768));
	notech_and4 i_68172437(.A(n_3970), .B(n_1806), .C(n_730), .D(n_3079), .Z
		(n_168893773));
	notech_and4 i_68472435(.A(n_733), .B(n_738), .C(n_168893773), .D(n_3197)
		, .Z(n_169093775));
	notech_and2 i_26973073(.A(n_3109), .B(n_169093775), .Z(n_169193776));
	notech_and4 i_70172426(.A(n_2327), .B(n_4032), .C(n_853), .D(n_214094151
		), .Z(n_169493779));
	notech_and4 i_69972428(.A(n_717), .B(n_2246), .C(n_4014), .D(n_4013), .Z
		(n_169793782));
	notech_and3 i_69272432(.A(n_1984), .B(n_1801), .C(n_1993), .Z(n_169893783
		));
	notech_and4 i_70372425(.A(n_4034), .B(n_169793782), .C(n_4085), .D(n_169893783
		), .Z(n_170393786));
	notech_and4 i_70772422(.A(n_222294221), .B(n_169493779), .C(n_208149924)
		, .D(n_170393786), .Z(n_170793789));
	notech_and4 i_72372411(.A(n_214394154), .B(n_3992), .C(n_202794052), .D(n_692
		), .Z(n_171693795));
	notech_nand3 i_72772408(.A(n_171693795), .B(n_2627), .C(n_30695), .Z(n_171793796
		));
	notech_and4 i_72472410(.A(n_709), .B(n_719), .C(n_703), .D(n_4008), .Z(n_172193799
		));
	notech_and4 i_72672409(.A(n_2760), .B(n_4032), .C(n_3143), .D(n_3980), .Z
		(n_172493802));
	notech_or4 i_73372404(.A(n_30765), .B(n_171793796), .C(n_155193657), .D(n_30764
		), .Z(n_172793805));
	notech_and4 i_74772393(.A(n_4041), .B(n_4036), .C(n_720), .D(n_673), .Z(n_173393809
		));
	notech_and4 i_74872392(.A(n_214394154), .B(n_4028), .C(n_1718), .D(n_222894227
		), .Z(n_173893813));
	notech_and2 i_74572395(.A(n_1332), .B(n_212094132), .Z(n_174093815));
	notech_and4 i_75172389(.A(n_222694225), .B(n_4029), .C(n_174093815), .D(n_173893813
		), .Z(n_174293817));
	notech_and4 i_75272388(.A(n_173393809), .B(n_174293817), .C(n_1950), .D(n_30696
		), .Z(n_174393818));
	notech_and4 i_76372377(.A(n_2099), .B(n_4016), .C(n_4026), .D(n_2538), .Z
		(n_174793822));
	notech_and4 i_76872373(.A(n_4055), .B(n_2894), .C(n_174793822), .D(n_1770
		), .Z(n_175093824));
	notech_and4 i_76172379(.A(n_1290), .B(n_4014), .C(n_720), .D(n_1999), .Z
		(n_175693828));
	notech_and4 i_76272378(.A(n_1718), .B(n_3967), .C(n_30719), .D(n_2760), 
		.Z(n_175993831));
	notech_and4 i_77072371(.A(n_175993831), .B(n_175693828), .C(n_1960), .D(n_30698
		), .Z(n_176293834));
	notech_and2 i_77573035(.A(n_1434), .B(n_122293382), .Z(n_176693837));
	notech_and4 i_79872346(.A(n_4053), .B(n_200294031), .C(n_4027), .D(n_1615
		), .Z(n_177593843));
	notech_and4 i_80172343(.A(n_493), .B(n_4084), .C(n_177593843), .D(n_497)
		, .Z(n_177693844));
	notech_and2 i_79372350(.A(n_4038), .B(n_191193959), .Z(n_178193846));
	notech_and4 i_80072344(.A(n_1537), .B(n_2760), .C(n_2928), .D(n_2571), .Z
		(n_178793850));
	notech_and4 i_80272342(.A(n_178193846), .B(n_178793850), .C(n_2080), .D(n_1996
		), .Z(n_178993851));
	notech_and4 i_80872338(.A(n_177693844), .B(n_176693837), .C(n_3280), .D(n_178993851
		), .Z(n_179193853));
	notech_and4 i_82872319(.A(n_2928), .B(n_853), .C(n_730), .D(n_4047), .Z(n_179493856
		));
	notech_and4 i_82372324(.A(n_2678), .B(n_2791), .C(n_533), .D(n_2884), .Z
		(n_180093861));
	notech_and4 i_81272334(.A(n_2631), .B(n_1780), .C(n_2137), .D(n_2757), .Z
		(n_180393864));
	notech_and4 i_82572322(.A(n_2157), .B(n_2212), .C(n_4049), .D(n_2029), .Z
		(n_180793868));
	notech_and4 i_83072317(.A(n_574), .B(n_466), .C(n_180393864), .D(n_180793868
		), .Z(n_180893869));
	notech_and4 i_83372314(.A(n_4004), .B(n_2538), .C(n_180093861), .D(n_180893869
		), .Z(n_180993870));
	notech_and4 i_82672321(.A(n_3987), .B(n_537), .C(n_202094047), .D(n_1777
		), .Z(n_181293873));
	notech_and4 i_82772320(.A(n_3973), .B(n_4037), .C(n_1504), .D(n_4005), .Z
		(n_181793876));
	notech_and4 i_83672311(.A(n_181793876), .B(n_181293873), .C(n_2435), .D(n_180993870
		), .Z(n_182093879));
	notech_and4 i_85672291(.A(n_2398), .B(n_4004), .C(n_4084), .D(n_1923), .Z
		(n_182493882));
	notech_and4 i_85172296(.A(n_4002), .B(n_4076), .C(n_2377), .D(n_4064), .Z
		(n_183093887));
	notech_and4 i_85272295(.A(n_1970), .B(n_1526), .C(n_530), .D(n_2058), .Z
		(n_183593891));
	notech_ao3 i_84372304(.A(n_2216), .B(n_455), .C(n_1987), .Z(n_183893893)
		);
	notech_and4 i_85872289(.A(n_183593891), .B(n_1603), .C(n_3975), .D(n_183893893
		), .Z(n_184193895));
	notech_and4 i_86172286(.A(n_4017), .B(n_183093887), .C(n_184193895), .D(n_2380
		), .Z(n_184293896));
	notech_nand3 i_86372284(.A(n_182493882), .B(n_176693837), .C(n_184293896
		), .Z(n_184393897));
	notech_ao4 i_84572302(.A(n_3957), .B(n_3954), .C(n_3963), .D(n_2517), .Z
		(n_184593899));
	notech_and4 i_85572292(.A(n_3993), .B(n_493), .C(n_3973), .D(n_4085), .Z
		(n_184993903));
	notech_and4 i_85972288(.A(n_1306), .B(n_184593899), .C(n_184993903), .D(n_1340
		), .Z(n_185093904));
	notech_and3 i_76673036(.A(n_2141), .B(n_4013), .C(n_2484), .Z(n_185393907
		));
	notech_and4 i_86972278(.A(n_3374), .B(n_3880), .C(n_4079), .D(n_3981), .Z
		(n_185593909));
	notech_and4 i_87072277(.A(n_4046), .B(n_4053), .C(n_2171), .D(n_4058), .Z
		(n_185993912));
	notech_and4 i_87872269(.A(n_4084), .B(n_2394), .C(n_520), .D(n_3982), .Z
		(n_186493917));
	notech_and4 i_88372265(.A(n_444), .B(n_4046), .C(n_186493917), .D(n_185393907
		), .Z(n_186793919));
	notech_and4 i_87972268(.A(n_2024), .B(n_2047), .C(n_1780), .D(n_201494043
		), .Z(n_187293922));
	notech_and4 i_89672252(.A(n_1346), .B(n_204), .C(n_1284), .D(n_215), .Z(n_187793927
		));
	notech_and4 i_89772251(.A(n_2171), .B(n_530), .C(n_218), .D(n_254), .Z(n_188093930
		));
	notech_and4 i_89872250(.A(n_3975), .B(n_4085), .C(n_30721), .D(n_1615), 
		.Z(n_188593935));
	notech_ao3 i_89572253(.A(n_1130), .B(n_30699), .C(n_122393383), .Z(n_188993939
		));
	notech_and3 i_89972249(.A(n_69848720), .B(n_4004), .C(n_188993939), .Z(n_189093940
		));
	notech_and4 i_90472244(.A(n_189093940), .B(n_185393907), .C(n_2434), .D(n_188593935
		), .Z(n_189293942));
	notech_nao3 i_90672242(.A(n_1919), .B(n_30720), .C(n_2164), .Z(n_189493944
		));
	notech_or4 i_90972239(.A(n_30700), .B(n_189493944), .C(n_30718), .D(n_30780
		), .Z(n_189693946));
	notech_or4 i_14873084(.A(n_4011), .B(n_1640), .C(n_4009), .D(n_189693946
		), .Z(n_189793947));
	notech_or4 i_15873082(.A(n_124093399), .B(n_30781), .C(\udeco[5] ), .D(n_189693946
		), .Z(n_190093949));
	notech_nand3 i_10393453(.A(n_3779), .B(n_1865), .C(n_194993992), .Z(n_190893956
		));
	notech_and4 i_10293454(.A(n_2352), .B(n_2654), .C(n_1856), .D(n_2344), .Z
		(n_190993957));
	notech_or4 i_118393456(.A(n_58492), .B(n_3935), .C(n_58510), .D(n_58519)
		, .Z(n_191193959));
	notech_nand2 i_114093458(.A(modrm[3]), .B(n_30786), .Z(n_191393961));
	notech_and2 i_113793459(.A(n_3763), .B(n_30704), .Z(n_191493962));
	notech_and2 i_113993460(.A(modrm[0]), .B(n_190893956), .Z(n_191593963)
		);
	notech_or4 i_92993461(.A(n_1321), .B(n_191493962), .C(n_191593963), .D(n_30796
		), .Z(\udeco[124] ));
	notech_and3 i_33693463(.A(n_2302), .B(n_30801), .C(n_30702), .Z(n_191793965
		));
	notech_or4 i_116493464(.A(n_2348), .B(n_58408), .C(n_58363), .D(n_191793965
		), .Z(n_191893966));
	notech_nao3 i_116393465(.A(n_30658), .B(n_30655), .C(n_2318), .Z(n_191993967
		));
	notech_and4 i_89293466(.A(n_199894027), .B(n_199494024), .C(n_2694), .D(n_1942
		), .Z(udeco_119100241));
	notech_nand3 i_14893467(.A(n_3736), .B(n_2099), .C(n_1905), .Z(n_192193968
		));
	notech_or4 i_141093469(.A(n_58492), .B(n_2316), .C(n_2389), .D(n_3761), 
		.Z(n_192693970));
	notech_nand2 i_141293470(.A(modrm[0]), .B(n_192193968), .Z(n_192793971)
		);
	notech_and2 i_140993471(.A(modrm[3]), .B(n_3773), .Z(n_192993972));
	notech_and2 i_141193472(.A(n_30705), .B(n_30768), .Z(n_193093973));
	notech_or4 i_85093473(.A(n_1321), .B(n_192993972), .C(n_30804), .D(n_193093973
		), .Z(\udeco[116] ));
	notech_or4 i_144393474(.A(n_58354), .B(n_2373), .C(n_58390), .D(n_2401),
		 .Z(n_193193974));
	notech_and4 i_84293475(.A(n_204594069), .B(n_201794045), .C(n_2684), .D(n_2890
		), .Z(udeco_114100240));
	notech_and4 i_82093476(.A(n_2704), .B(n_2684), .C(n_207794095), .D(n_2890
		), .Z(udeco_113100239));
	notech_or4 i_168293477(.A(n_58354), .B(n_2373), .C(n_3845), .D(n_58426),
		 .Z(n_193293975));
	notech_or4 i_168693478(.A(n_58492), .B(n_2313), .C(n_58372), .D(n_2348),
		 .Z(n_193393976));
	notech_and2 i_168593479(.A(opz[0]), .B(n_30708), .Z(n_193493977));
	notech_or4 i_66293480(.A(n_193493977), .B(n_209294109), .C(n_30813), .D(n_30810
		), .Z(\udeco[104] ));
	notech_and2 i_12693481(.A(n_3992), .B(n_3876), .Z(n_5254));
	notech_nao3 i_62893485(.A(n_211494128), .B(n_5254), .C(n_210194116), .Z(\udeco[49] 
		));
	notech_or4 i_172393486(.A(n_58354), .B(n_2037), .C(n_4072), .D(n_58426),
		 .Z(n_193893981));
	notech_and4 i_58293487(.A(n_193893981), .B(n_213894149), .C(n_1593), .D(n_894
		), .Z(udeco_37100238));
	notech_nao3 i_175093490(.A(n_30658), .B(n_30793), .C(n_2499), .Z(n_194193984
		));
	notech_or2 i_174793491(.A(n_2124), .B(n_58555), .Z(n_194293985));
	notech_or4 i_174993492(.A(n_58354), .B(n_2315), .C(n_58390), .D(n_3836),
		 .Z(n_194393986));
	notech_nao3 i_56110332(.A(n_216894173), .B(n_214394154), .C(n_1326), .Z(\udeco[34] 
		));
	notech_or2 i_182693493(.A(n_2151), .B(n_58456), .Z(n_194493987));
	notech_or2 i_182893494(.A(n_3697), .B(n_58555), .Z(n_194593988));
	notech_or2 i_182793495(.A(n_3728), .B(n_58390), .Z(n_194693989));
	notech_nao3 i_49493496(.A(n_717), .B(n_219694198), .C(n_1326), .Z(\udeco[26] 
		));
	notech_and4 i_47210354(.A(n_520), .B(n_537), .C(n_2567), .D(n_221594215)
		, .Z(udeco_23100237));
	notech_nao3 i_34693497(.A(n_1951), .B(n_2380), .C(n_4057), .Z(n_1326));
	notech_or4 i_17293499(.A(n_1326), .B(n_30818), .C(n_30701), .D(n_3978), 
		.Z(n_1321));
	notech_ao3 i_113193501(.A(n_3777), .B(n_3987), .C(n_3846), .Z(n_194993992
		));
	notech_ao4 i_114293505(.A(n_58481), .B(n_4070), .C(n_2348), .D(n_2338), 
		.Z(n_195693996));
	notech_ao4 i_114393506(.A(n_2166), .B(n_3760), .C(n_30785), .D(n_3935), 
		.Z(n_195793997));
	notech_and4 i_114693509(.A(n_195793997), .B(n_195693996), .C(n_3834), .D
		(n_247292237), .Z(n_196294000));
	notech_and4 i_114993512(.A(n_2450), .B(n_196294000), .C(n_1834), .D(n_191393961
		), .Z(n_196594003));
	notech_and3 i_116693516(.A(n_2676), .B(n_191993967), .C(n_191893966), .Z
		(n_197394007));
	notech_nand2 i_14393518(.A(n_2629), .B(n_30723), .Z(n_1249));
	notech_nand2 i_22193520(.A(n_30836), .B(n_30726), .Z(n_1180));
	notech_and4 i_26693523(.A(n_2216), .B(n_2709), .C(n_2151), .D(n_30792), 
		.Z(n_1130));
	notech_and4 i_133193524(.A(n_2231), .B(n_1833), .C(n_2188), .D(n_1907), 
		.Z(n_197794011));
	notech_and4 i_133393527(.A(n_2630), .B(n_3733), .C(n_3993), .D(n_197794011
		), .Z(n_198194014));
	notech_and4 i_133693530(.A(n_198194014), .B(n_2638), .C(n_1130), .D(n_2065
		), .Z(n_198594017));
	notech_and3 i_133893532(.A(n_4002), .B(n_2166), .C(n_2829), .Z(n_198894019
		));
	notech_and4 i_134093534(.A(n_2827), .B(n_198594017), .C(n_198894019), .D
		(n_2414), .Z(n_199094021));
	notech_and4 i_134693537(.A(n_2826), .B(n_199094021), .C(n_2707), .D(n_1920
		), .Z(n_199494024));
	notech_and4 i_134593540(.A(n_2522), .B(n_2831), .C(n_2510), .D(n_2605), 
		.Z(n_199894027));
	notech_and2 i_61093543(.A(n_4029), .B(n_3967), .Z(n_200294031));
	notech_ao4 i_141393544(.A(n_1984), .B(n_58481), .C(n_2383), .D(n_2865), 
		.Z(n_200394032));
	notech_and4 i_141693547(.A(n_200394032), .B(n_2857), .C(n_192693970), .D
		(n_30706), .Z(n_200694035));
	notech_and4 i_141893549(.A(n_2479), .B(n_200694035), .C(n_30724), .D(n_30797
		), .Z(n_200894037));
	notech_and4 i_142193552(.A(n_200294031), .B(n_200894037), .C(n_2884), .D
		(n_192793971), .Z(n_201194040));
	notech_and2 i_61293555(.A(n_1993), .B(n_4040), .Z(n_201494043));
	notech_and4 i_146693557(.A(n_1993), .B(n_4040), .C(n_2309), .D(n_2483), 
		.Z(n_201794045));
	notech_and4 i_25793559(.A(n_1886), .B(n_2686), .C(n_2572), .D(n_2899), .Z
		(n_202094047));
	notech_and4 i_71093564(.A(n_4007), .B(n_3672), .C(n_1537), .D(n_193193974
		), .Z(n_202794052));
	notech_and4 i_144893567(.A(n_2629), .B(n_3964), .C(n_2709), .D(n_30709),
		 .Z(n_203194055));
	notech_and4 i_145193570(.A(n_2765), .B(n_3867), .C(n_203194055), .D(n_2124
		), .Z(n_203494058));
	notech_and3 i_145393572(.A(n_1949), .B(n_1796), .C(n_3880), .Z(n_203694060
		));
	notech_and4 i_145693574(.A(n_3777), .B(n_203494058), .C(n_1526), .D(n_203694060
		), .Z(n_203894062));
	notech_and4 i_145993577(.A(n_203894062), .B(n_198894019), .C(n_2655), .D
		(n_202794052), .Z(n_204194065));
	notech_and4 i_146593580(.A(n_2903), .B(n_2605), .C(n_204194065), .D(n_1504
		), .Z(n_204494068));
	notech_and4 i_146793581(.A(n_2898), .B(n_202094047), .C(n_2893), .D(n_204494068
		), .Z(n_204594069));
	notech_and4 i_148693587(.A(n_3994), .B(n_2839), .C(n_202794052), .D(n_2852
		), .Z(n_205494075));
	notech_ao3 i_147293590(.A(n_2516), .B(n_30707), .C(n_4010), .Z(n_205794078
		));
	notech_and4 i_147593593(.A(n_2765), .B(n_3931), .C(n_3751), .D(n_205794078
		), .Z(n_206194081));
	notech_and4 i_147893596(.A(n_2625), .B(n_2176), .C(n_206194081), .D(n_2591
		), .Z(n_206494084));
	notech_and4 i_148293599(.A(n_2332), .B(n_206494084), .C(n_2534), .D(n_2539
		), .Z(n_206894087));
	notech_and4 i_148793601(.A(n_2572), .B(n_1969), .C(n_206894087), .D(n_2656
		), .Z(n_207094089));
	notech_and4 i_149093604(.A(n_2722), .B(n_2898), .C(n_207094089), .D(n_2850
		), .Z(n_207394092));
	notech_and4 i_149293605(.A(n_4040), .B(n_205494075), .C(n_207394092), .D
		(n_1993), .Z(n_207494093));
	notech_and4 i_149493607(.A(n_2834), .B(n_2893), .C(n_207494093), .D(n_2688
		), .Z(n_207794095));
	notech_and2 i_72093610(.A(n_3973), .B(n_4029), .Z(n_843));
	notech_and4 i_26493613(.A(n_2327), .B(n_193293975), .C(n_3665), .D(n_30856
		), .Z(n_208394100));
	notech_and4 i_168993616(.A(n_3998), .B(n_193393976), .C(n_3890), .D(n_30709
		), .Z(n_208694103));
	notech_and4 i_169293619(.A(n_208694103), .B(n_1290), .C(n_2162), .D(n_2380
		), .Z(n_208994106));
	notech_or4 i_169593622(.A(n_3820), .B(n_30710), .C(n_1249), .D(n_30811),
		 .Z(n_209294109));
	notech_nand3 i_4353(.A(n_223492236), .B(n_1792), .C(n_1999), .Z(n_209694112
		));
	notech_and4 i_4356(.A(n_30712), .B(n_4019), .C(n_30713), .D(n_1972), .Z(n_210094115
		));
	notech_or4 i_37393627(.A(n_30830), .B(n_30814), .C(n_30816), .D(n_1180),
		 .Z(n_210194116));
	notech_and2 i_4347(.A(n_4026), .B(n_3982), .Z(n_69848720));
	notech_and2 i_4298(.A(n_3838), .B(n_3987), .Z(n_210394118));
	notech_ao4 i_65093629(.A(n_2113), .B(n_2373), .C(n_2278), .D(n_2346), .Z
		(n_210494119));
	notech_ao4 i_170693630(.A(n_2275), .B(n_2118), .C(n_2564), .D(n_58417), 
		.Z(n_210594120));
	notech_and4 i_170993633(.A(n_210594120), .B(n_210494119), .C(n_4031), .D
		(n_1816), .Z(n_210894123));
	notech_and4 i_171393636(.A(n_2340), .B(n_210894123), .C(n_2099), .D(n_210394118
		), .Z(n_211194126));
	notech_and4 i_171593638(.A(n_4032), .B(n_4030), .C(n_211194126), .D(n_69848720
		), .Z(n_211494128));
	notech_and4 i_80793640(.A(n_4076), .B(n_193893981), .C(n_2615), .D(n_2091
		), .Z(n_211794130));
	notech_ao3 i_4572(.A(n_4014), .B(n_1329), .C(n_30661), .Z(n_212094132)
		);
	notech_and4 i_173893643(.A(n_872), .B(n_2500), .C(n_212094132), .D(n_200294031
		), .Z(n_212294134));
	notech_and2 i_74293644(.A(n_3994), .B(n_4085), .Z(n_692));
	notech_and3 i_4510(.A(n_2629), .B(n_4086), .C(n_30723), .Z(n_212494135)
		);
	notech_and4 i_172693648(.A(n_3973), .B(n_3736), .C(n_4031), .D(n_1114), 
		.Z(n_212894139));
	notech_and4 i_172993651(.A(n_212894139), .B(n_2743), .C(n_3061), .D(n_30714
		), .Z(n_213194142));
	notech_and4 i_173393654(.A(n_4034), .B(n_213194142), .C(n_2465), .D(n_861
		), .Z(n_213494145));
	notech_and4 i_173793656(.A(n_2036), .B(n_1014), .C(n_213494145), .D(n_30838
		), .Z(n_213694147));
	notech_and4 i_174093658(.A(n_3994), .B(n_213694147), .C(n_212294134), .D
		(n_4085), .Z(n_213894149));
	notech_and4 i_4614(.A(n_2192), .B(n_4017), .C(n_2500), .D(n_3981), .Z(n_214094151
		));
	notech_and4 i_4656(.A(n_2663), .B(n_2327), .C(n_214094151), .D(n_30797),
		 .Z(n_214394154));
	notech_ao3 i_4531(.A(n_4041), .B(n_1896), .C(n_222394222), .Z(n_214594156
		));
	notech_nand2 i_351093665(.A(n_30726), .B(n_30722), .Z(n_214994159));
	notech_ao4 i_175193666(.A(n_58456), .B(n_30792), .C(n_58390), .D(n_30834
		), .Z(n_215094160));
	notech_and4 i_175493669(.A(n_215094160), .B(n_3992), .C(n_194193984), .D
		(n_30829), .Z(n_215494163));
	notech_and4 i_175993672(.A(n_215494163), .B(n_194293985), .C(n_2017), .D
		(n_194393986), .Z(n_215894166));
	notech_and4 i_176093673(.A(n_811), .B(n_2340), .C(n_214594156), .D(n_215894166
		), .Z(n_215994167));
	notech_and4 i_176393675(.A(n_4055), .B(n_2538), .C(n_843), .D(n_215994167
		), .Z(n_216194169));
	notech_and4 i_176493676(.A(n_2099), .B(n_216194169), .C(n_3736), .D(n_2116
		), .Z(n_216294170));
	notech_and4 i_176793679(.A(n_960), .B(n_894), .C(n_2903), .D(n_216294170
		), .Z(n_216894173));
	notech_and3 i_184493682(.A(n_3102), .B(n_738), .C(n_2588), .Z(n_217294176
		));
	notech_and4 i_184893684(.A(n_30797), .B(n_217294176), .C(n_3098), .D(n_30693
		), .Z(n_217494178));
	notech_and4 i_183193688(.A(n_4026), .B(n_4041), .C(n_4013), .D(n_3980), 
		.Z(n_217994182));
	notech_and3 i_183493690(.A(n_217994182), .B(n_2305), .C(n_30719), .Z(n_218194184
		));
	notech_and4 i_183893692(.A(n_1290), .B(n_194493987), .C(n_218194184), .D
		(n_194593988), .Z(n_218494186));
	notech_and4 i_183993696(.A(n_3103), .B(n_853), .C(n_2099), .D(n_2533), .Z
		(n_218894190));
	notech_and4 i_184393698(.A(n_218894190), .B(n_2465), .C(n_218494186), .D
		(n_2015), .Z(n_219094192));
	notech_and4 i_184993701(.A(n_219094192), .B(n_222894227), .C(n_30720), .D
		(n_194693989), .Z(n_219394195));
	notech_and4 i_185293704(.A(n_703), .B(n_2246), .C(n_219394195), .D(n_217494178
		), .Z(n_219694198));
	notech_and4 i_195593708(.A(n_3049), .B(n_2723), .C(n_2928), .D(n_2024), 
		.Z(n_220094202));
	notech_and3 i_194793711(.A(n_4048), .B(n_4047), .C(n_4019), .Z(n_220394205
		));
	notech_and4 i_195093714(.A(n_2365), .B(n_3739), .C(n_4049), .D(n_220394205
		), .Z(n_220694208));
	notech_and4 i_195693717(.A(n_2212), .B(n_2522), .C(n_200294031), .D(n_220694208
		), .Z(n_220994211));
	notech_and4 i_195993719(.A(n_2157), .B(n_220994211), .C(n_3177), .D(n_220094202
		), .Z(n_221194213));
	notech_and4 i_196193721(.A(n_1993), .B(n_4040), .C(n_221194213), .D(n_530
		), .Z(n_221594215));
	notech_nand3 i_20073105(.A(n_2123), .B(n_4034), .C(n_4022), .Z(n_221894218
		));
	notech_and2 i_413973095(.A(n_30695), .B(n_4062), .Z(n_2219));
	notech_and3 i_4288(.A(n_3992), .B(n_3876), .C(n_2377), .Z(n_222194220)
		);
	notech_and3 i_61773054(.A(n_4067), .B(n_4022), .C(n_30713), .Z(n_222294221
		));
	notech_and4 i_173027(.A(n_2344), .B(n_3279), .C(n_3545), .D(n_1856), .Z(n_1607
		));
	notech_ao3 i_16193724(.A(n_30855), .B(n_3895), .C(n_2348), .Z(n_222394222
		));
	notech_or2 i_3625(.A(n_4089), .B(n_4024), .Z(n_222494223));
	notech_nand3 i_3834(.A(n_2073), .B(n_2202), .C(n_4082), .Z(n_222594224)
		);
	notech_ao4 i_4638(.A(n_2303), .B(n_30800), .C(n_30789), .D(n_2291), .Z(n_222694225
		));
	notech_nand2 i_4672982(.A(modrm[4]), .B(n_30875), .Z(n_1606));
	notech_ao4 i_41793725(.A(n_4072), .B(n_30787), .C(n_30791), .D(n_4090), 
		.Z(n_222794226));
	notech_ao4 i_55993726(.A(n_3954), .B(n_3957), .C(n_2339), .D(n_2299), .Z
		(n_222894227));
	notech_nand3 i_69593727(.A(n_2587), .B(n_197394007), .C(n_2722), .Z(n_222994228
		));
	notech_nand3 i_79793728(.A(n_4086), .B(n_4044), .C(n_30797), .Z(n_223094229
		));
	notech_nand2 i_4172987(.A(n_2390), .B(n_1791), .Z(n_1604));
	notech_inv i_36373(.A(n_1614), .Z(\udeco[125] ));
	notech_inv i_36374(.A(n_1620), .Z(\udeco[123] ));
	notech_inv i_36375(.A(n_1628), .Z(\udeco[45] ));
	notech_inv i_36376(.A(n_1802), .Z(n_30653));
	notech_inv i_36377(.A(n_1639), .Z(\udeco[27] ));
	notech_inv i_36378(.A(n_2027), .Z(n_30655));
	notech_inv i_36379(.A(n_2359), .Z(n_30656));
	notech_inv i_36380(.A(n_2469), .Z(n_30657));
	notech_inv i_36381(.A(n_2149), .Z(n_30658));
	notech_inv i_36382(.A(n_58417), .Z(n_30659));
	notech_inv i_36383(.A(n_2059), .Z(n_30660));
	notech_inv i_36384(.A(n_2005), .Z(n_30661));
	notech_inv i_36385(.A(n_2098), .Z(n_30662));
	notech_inv i_36386(.A(n_2202), .Z(n_30663));
	notech_inv i_36387(.A(n_2078), .Z(n_30664));
	notech_inv i_36388(.A(n_2013), .Z(n_30665));
	notech_inv i_36389(.A(n_2020), .Z(\udeco[112] ));
	notech_inv i_36390(.A(n_2055), .Z(\udeco[109] ));
	notech_inv i_36391(.A(n_2092), .Z(\udeco[32] ));
	notech_inv i_36392(.A(n_2127), .Z(\udeco[24] ));
	notech_inv i_36393(.A(n_2135), .Z(\udeco[20] ));
	notech_inv i_36394(.A(n_2146), .Z(\udeco[18] ));
	notech_inv i_36395(.A(n_2177), .Z(\udeco[17] ));
	notech_inv i_36396(.A(n_2208), .Z(\udeco[13] ));
	notech_inv i_36397(.A(n_221992235), .Z(\udeco[11] ));
	notech_inv i_36398(.A(n_2227), .Z(\udeco[10] ));
	notech_inv i_36399(.A(n_2241), .Z(\udeco[9] ));
	notech_inv i_36400(.A(n_2270), .Z(\udeco[0] ));
	notech_inv i_36401(.A(n_4003), .Z(n_30678));
	notech_inv i_36402(.A(n_4080), .Z(n_30679));
	notech_inv i_36403(.A(n_3974), .Z(n_30680));
	notech_inv i_36404(.A(n_207949923), .Z(n_30681));
	notech_inv i_36405(.A(n_4018), .Z(n_30682));
	notech_inv i_36406(.A(n_4093), .Z(n_30683));
	notech_inv i_36407(.A(n_4062), .Z(n_30684));
	notech_inv i_36408(.A(n_4057), .Z(n_30685));
	notech_inv i_36409(.A(n_4052), .Z(n_30686));
	notech_inv i_36410(.A(n_4091), .Z(n_30687));
	notech_inv i_36411(.A(n_4054), .Z(n_30688));
	notech_inv i_36412(.A(n_4050), .Z(n_30689));
	notech_inv i_36413(.A(n_4065), .Z(n_30690));
	notech_inv i_36414(.A(n_3969), .Z(n_30691));
	notech_inv i_36415(.A(n_4060), .Z(n_30692));
	notech_inv i_36416(.A(n_4015), .Z(n_30693));
	notech_inv i_36417(.A(n_4059), .Z(n_30694));
	notech_inv i_36418(.A(n_4045), .Z(n_30695));
	notech_inv i_36419(.A(n_3971), .Z(n_30696));
	notech_inv i_36420(.A(n_3981), .Z(n_30697));
	notech_inv i_36421(.A(n_204849898), .Z(n_30698));
	notech_inv i_36422(.A(n_4033), .Z(n_30699));
	notech_inv i_36423(.A(n_3984), .Z(n_30700));
	notech_inv i_36424(.A(n_4082), .Z(n_30701));
	notech_inv i_36425(.A(n_3908), .Z(n_30702));
	notech_inv i_36426(.A(n_3846), .Z(n_30703));
	notech_inv i_36427(.A(n_4071), .Z(n_30704));
	notech_inv i_36428(.A(n_3760), .Z(n_30705));
	notech_inv i_36429(.A(n_4006), .Z(n_30706));
	notech_inv i_36430(.A(n_4011), .Z(n_30707));
	notech_inv i_36431(.A(n_3955), .Z(n_30708));
	notech_inv i_36432(.A(n_4009), .Z(n_30709));
	notech_inv i_36433(.A(n_3972), .Z(n_30710));
	notech_inv i_36434(.A(n_3820), .Z(n_30711));
	notech_inv i_36435(.A(n_3990), .Z(n_30712));
	notech_inv i_36436(.A(n_4023), .Z(n_30713));
	notech_inv i_36437(.A(n_4035), .Z(n_30714));
	notech_inv i_36438(.A(n_3728), .Z(n_30715));
	notech_inv i_36439(.A(n_3697), .Z(n_30716));
	notech_inv i_36440(.A(n_3980), .Z(n_30717));
	notech_inv i_36441(.A(n_2305), .Z(n_30718));
	notech_inv i_36442(.A(n_4001), .Z(n_30719));
	notech_inv i_36443(.A(n_3986), .Z(n_30720));
	notech_inv i_36444(.A(n_4088), .Z(n_30721));
	notech_inv i_36445(.A(n_3978), .Z(n_30722));
	notech_inv i_36446(.A(n_3950), .Z(n_30723));
	notech_inv i_36447(.A(n_3985), .Z(n_30724));
	notech_inv i_36448(.A(n_4089), .Z(n_30725));
	notech_inv i_36449(.A(n_3968), .Z(n_30726));
	notech_inv i_36450(.A(n_4085), .Z(n_30727));
	notech_inv i_36451(.A(n_2102), .Z(n_30728));
	notech_inv i_36452(.A(n_2354), .Z(n_30729));
	notech_inv i_36453(.A(n_1708), .Z(n_30730));
	notech_inv i_36454(.A(n_1709), .Z(n_30731));
	notech_inv i_36455(.A(n_122893388), .Z(n_30732));
	notech_inv i_36456(.A(n_125893415), .Z(n_30733));
	notech_inv i_36457(.A(n_126993422), .Z(n_30734));
	notech_inv i_36458(.A(n_1712), .Z(n_30735));
	notech_inv i_36459(.A(n_1870), .Z(n_30736));
	notech_inv i_36460(.A(n_127693429), .Z(n_30737));
	notech_inv i_36461(.A(n_2397), .Z(n_30738));
	notech_inv i_36462(.A(n_133493473), .Z(n_30739));
	notech_inv i_36463(.A(n_136893500), .Z(n_30740));
	notech_inv i_36464(.A(n_138993517), .Z(n_30741));
	notech_inv i_36465(.A(n_1953), .Z(n_30742));
	notech_inv i_36466(.A(n_121193371), .Z(n_30743));
	notech_inv i_36467(.A(n_143893561), .Z(n_30744));
	notech_inv i_36468(.A(n_146993589), .Z(n_30745));
	notech_inv i_36469(.A(n_2614), .Z(n_30746));
	notech_inv i_36470(.A(n_2878), .Z(n_30747));
	notech_inv i_36471(.A(n_1978), .Z(n_30748));
	notech_inv i_36472(.A(n_2854), .Z(n_30749));
	notech_inv i_36473(.A(n_1623), .Z(n_30750));
	notech_inv i_36474(.A(n_153493645), .Z(n_30751));
	notech_inv i_36475(.A(n_2304), .Z(n_30752));
	notech_inv i_36476(.A(n_155193657), .Z(n_30753));
	notech_inv i_36477(.A(n_1981), .Z(n_30754));
	notech_inv i_36478(.A(n_1933), .Z(n_30755));
	notech_inv i_36479(.A(n_1704), .Z(n_30756));
	notech_inv i_36480(.A(n_1951), .Z(n_30757));
	notech_inv i_36481(.A(n_162293716), .Z(n_30758));
	notech_inv i_36482(.A(n_2759), .Z(n_30759));
	notech_inv i_36483(.A(n_2754), .Z(n_30760));
	notech_inv i_36484(.A(n_1702), .Z(n_30761));
	notech_inv i_36485(.A(n_3107), .Z(n_30762));
	notech_inv i_36486(.A(n_2713), .Z(n_30763));
	notech_inv i_36487(.A(n_172193799), .Z(n_30764));
	notech_inv i_36488(.A(n_172493802), .Z(n_30765));
	notech_inv i_36489(.A(n_2678), .Z(n_30766));
	notech_inv i_36490(.A(n_3510), .Z(n_30767));
	notech_inv i_36491(.A(n_1718), .Z(n_30768));
	notech_inv i_36492(.A(n_1699), .Z(n_30769));
	notech_inv i_36493(.A(n_1263), .Z(n_30770));
	notech_inv i_36494(.A(n_2620), .Z(n_30771));
	notech_inv i_36495(.A(n_2615), .Z(n_30772));
	notech_inv i_36496(.A(n_185093904), .Z(n_30773));
	notech_inv i_36497(.A(n_696), .Z(n_30774));
	notech_inv i_36498(.A(n_2543), .Z(n_30775));
	notech_inv i_36499(.A(n_2541), .Z(n_30776));
	notech_inv i_36500(.A(n_2536), .Z(n_30777));
	notech_inv i_36501(.A(n_1615), .Z(n_30778));
	notech_inv i_36502(.A(n_2296), .Z(n_30779));
	notech_inv i_36503(.A(n_1923), .Z(n_30780));
	notech_inv i_36504(.A(n_2022), .Z(n_30781));
	notech_inv i_36505(.A(n_190093949), .Z(n_30782));
	notech_inv i_36506(.A(n_2426), .Z(n_30783));
	notech_inv i_36507(.A(n_1969), .Z(n_30784));
	notech_inv i_36508(.A(n_2369), .Z(n_30785));
	notech_inv i_36509(.A(n_190993957), .Z(n_30786));
	notech_inv i_36510(.A(n_3959), .Z(n_30787));
	notech_inv i_36511(.A(n_1942), .Z(n_30788));
	notech_inv i_36512(.A(n_2390), .Z(n_30789));
	notech_inv i_36513(.A(n_2401), .Z(n_30790));
	notech_inv i_36514(.A(n_2210), .Z(n_30791));
	notech_inv i_36515(.A(n_1987), .Z(n_30792));
	notech_inv i_36516(.A(n_2355), .Z(n_30793));
	notech_inv i_36517(.A(n_2466), .Z(n_30794));
	notech_inv i_36518(.A(n_2463), .Z(n_30795));
	notech_inv i_36519(.A(n_196594003), .Z(n_30796));
	notech_inv i_36520(.A(n_1249), .Z(n_30797));
	notech_inv i_36521(.A(n_1180), .Z(n_30798));
	notech_inv i_36522(.A(n_2431), .Z(n_30799));
	notech_inv i_36523(.A(n_2418), .Z(n_30800));
	notech_inv i_36524(.A(n_2287), .Z(n_30801));
	notech_inv i_36525(.A(n_1905), .Z(n_30802));
	notech_inv i_36526(.A(n_2391), .Z(n_30803));
	notech_inv i_36527(.A(n_201194040), .Z(n_30804));
	notech_inv i_36528(.A(n_2852), .Z(n_30805));
	notech_inv i_36529(.A(n_2324), .Z(n_30806));
	notech_inv i_36530(.A(n_2321), .Z(n_30807));
	notech_inv i_36531(.A(n_2656), .Z(n_30808));
	notech_inv i_36532(.A(n_2850), .Z(n_30809));
	notech_inv i_36533(.A(n_208394100), .Z(n_30810));
	notech_inv i_36534(.A(n_208994106), .Z(n_30811));
	notech_inv i_36535(.A(n_2186), .Z(n_30812));
	notech_inv i_36536(.A(n_2792), .Z(n_30813));
	notech_inv i_36537(.A(n_1999), .Z(n_30814));
	notech_inv i_36538(.A(n_1972), .Z(n_30815));
	notech_inv i_36539(.A(n_210094115), .Z(n_30816));
	notech_inv i_36540(.A(n_2038), .Z(n_30817));
	notech_inv i_36541(.A(n_1816), .Z(n_30818));
	notech_inv i_36542(.A(n_2006), .Z(n_30819));
	notech_inv i_36543(.A(n_1986), .Z(n_30820));
	notech_inv i_36544(.A(n_1965), .Z(n_30821));
	notech_inv i_36545(.A(n_1624), .Z(n_30822));
	notech_inv i_36546(.A(n_2036), .Z(n_30823));
	notech_inv i_36547(.A(n_1943), .Z(n_30824));
	notech_inv i_36548(.A(n_1114), .Z(n_30825));
	notech_inv i_36549(.A(n_1841), .Z(n_30826));
	notech_inv i_36550(.A(n_1840), .Z(n_30827));
	notech_inv i_36551(.A(n_2116), .Z(n_30828));
	notech_inv i_36552(.A(n_214994159), .Z(n_30829));
	notech_inv i_36553(.A(n_2017), .Z(n_30830));
	notech_inv i_36554(.A(n_960), .Z(n_30831));
	notech_inv i_36555(.A(n_1695), .Z(n_30832));
	notech_inv i_36556(.A(n_2365), .Z(n_30833));
	notech_inv i_36557(.A(n_221894218), .Z(n_30834));
	notech_inv i_36558(.A(n_2357), .Z(n_30835));
	notech_inv i_36559(.A(n_222494223), .Z(n_30836));
	notech_inv i_36560(.A(n_2380), .Z(\udeco[5] ));
	notech_inv i_36561(.A(n_223094229), .Z(n_30838));
	notech_inv i_36562(.A(n_1950), .Z(n_30839));
	notech_inv i_36564(.A(n_58528), .Z(n_30841));
	notech_inv i_36565(.A(n_58514), .Z(n_30842));
	notech_inv i_36567(.A(n_58546), .Z(n_30844));
	notech_inv i_36568(.A(n_58568), .Z(n_30845));
	notech_inv i_36569(.A(op[7]), .Z(n_30846));
	notech_inv i_36570(.A(modrm[0]), .Z(n_30847));
	notech_inv i_36571(.A(modrm[1]), .Z(n_30848));
	notech_inv i_36572(.A(modrm[3]), .Z(n_30849));
	notech_inv i_36573(.A(modrm[4]), .Z(n_30850));
	notech_inv i_36574(.A(n_58426), .Z(n_30851));
	notech_inv i_36575(.A(modrm[6]), .Z(n_30852));
	notech_inv i_36576(.A(ipg_fault), .Z(n_30853));
	notech_inv i_36577(.A(twobyte), .Z(n_30854));
	notech_inv i_36578(.A(adz), .Z(n_30855));
	notech_inv i_36579(.A(n_4024), .Z(n_30856));
	notech_inv i_36580(.A(n_1622), .Z(n_30857));
	notech_inv i_36581(.A(n_1608), .Z(n_30858));
	notech_inv i_36582(.A(\udeco[91] ), .Z(n_30859));
	notech_inv i_36583(.A(udeco_73100251), .Z(\udeco[73] ));
	notech_inv i_36584(.A(udeco_101100250), .Z(\udeco[101] ));
	notech_inv i_36585(.A(udeco_103100249), .Z(\udeco[103] ));
	notech_inv i_36586(.A(udeco_35100248), .Z(\udeco[35] ));
	notech_inv i_36587(.A(udeco_29100247), .Z(\udeco[29] ));
	notech_inv i_36588(.A(udeco_28100246), .Z(\udeco[28] ));
	notech_inv i_36589(.A(udeco_21100245), .Z(\udeco[21] ));
	notech_inv i_36590(.A(udeco_15100244), .Z(\udeco[15] ));
	notech_inv i_36591(.A(udeco_14100243), .Z(\udeco[14] ));
	notech_inv i_36592(.A(udeco_12100242), .Z(\udeco[12] ));
	notech_inv i_36593(.A(udeco_119100241), .Z(\udeco[119] ));
	notech_inv i_36594(.A(udeco_114100240), .Z(\udeco[114] ));
	notech_inv i_36595(.A(udeco_113100239), .Z(\udeco[113] ));
	notech_inv i_36596(.A(udeco_37100238), .Z(\udeco[37] ));
	notech_inv i_36597(.A(udeco_23100237), .Z(\udeco[23] ));
	notech_inv i_36598(.A(n_1607), .Z(n_30875));
endmodule
module deco(clk, rstn, useq_ptr, in128, adz, pc_req, ivect, int_main, iack, ie, pg_fault
		, ipg_fault, cpl, cr0, valid_len, to_vliw, lenpc_out, immediate,
		 to_acu, operand_size, reps, over_seg, valid_op, term, start, ready_vliw
		);

	input clk;
	input rstn;
	output [3:0] useq_ptr;
	input [127:0] in128;
	input adz;
	input pc_req;
	input [7:0] ivect;
	input int_main;
	output iack;
	input ie;
	input pg_fault;
	input ipg_fault;
	input [1:0] cpl;
	input [31:0] cr0;
	input [5:0] valid_len;
	output [127:0] to_vliw;
	output [31:0] lenpc_out;
	output [63:0] immediate;
	output [210:0] to_acu;
	output [2:0] operand_size;
	output [2:0] reps;
	output [5:0] over_seg;
	output valid_op;
	input term;
	output start;
	input ready_vliw;

	wire [210:0] to_acu2;
	wire [31:0] lenpc2;
	wire [2:0] opz2;
	wire [2:0] reps1;
	wire [127:0] inst_deco1;
	wire [2:0] opz1;
	wire [127:0] inst_deco2;
	wire [210:0] to_acu1;
	wire [3:0] i_ptr;
	wire [5:0] int_excl;
	wire [1:0] idx_deco;
	wire [2:0] reps2;
	wire [7:0] ififo_rvect1;
	wire [4:0] fsm;
	wire [31:0] lenpc1;
	wire [210:0] to_acu0;
	wire [127:0] inst_deco;
	wire [2:0] opz0;
	wire [2:0] reps0;
	wire [31:0] lenpc;
	wire [7:0] ififo_rvect2;
	wire [7:0] ififo_rvect3;
	wire [7:0] ififo_rvect4;
	wire [127:0] udeco;
	wire [2:0] displc;
	wire [2:0] opz;
	wire [2:0] imm_sz;
	wire [4:0] pfx_sz;



	notech_inv i_15589(.A(n_62280), .Z(n_62343));
	notech_inv i_15587(.A(n_62280), .Z(n_62341));
	notech_inv i_15584(.A(n_62280), .Z(n_62338));
	notech_inv i_15582(.A(n_62280), .Z(n_62336));
	notech_inv i_15579(.A(n_62280), .Z(n_62333));
	notech_inv i_15577(.A(n_62280), .Z(n_62331));
	notech_inv i_15573(.A(n_62280), .Z(n_62327));
	notech_inv i_15571(.A(n_62280), .Z(n_62325));
	notech_inv i_15568(.A(n_62280), .Z(n_62322));
	notech_inv i_15566(.A(n_62280), .Z(n_62320));
	notech_inv i_15563(.A(n_62280), .Z(n_62317));
	notech_inv i_15561(.A(n_62280), .Z(n_62315));
	notech_inv i_15557(.A(n_62280), .Z(n_62311));
	notech_inv i_15555(.A(n_62280), .Z(n_62309));
	notech_inv i_15552(.A(n_62280), .Z(n_62306));
	notech_inv i_15550(.A(n_62280), .Z(n_62304));
	notech_inv i_15547(.A(n_62280), .Z(n_62301));
	notech_inv i_15545(.A(n_62280), .Z(n_62299));
	notech_inv i_15541(.A(n_62282), .Z(n_62295));
	notech_inv i_15539(.A(n_62282), .Z(n_62293));
	notech_inv i_15536(.A(n_62282), .Z(n_62290));
	notech_inv i_15534(.A(n_62282), .Z(n_62288));
	notech_inv i_15531(.A(n_62282), .Z(n_62285));
	notech_inv i_15529(.A(n_62282), .Z(n_62283));
	notech_inv i_15528(.A(n_62281), .Z(n_62282));
	notech_inv i_15527(.A(n_62280), .Z(n_62281));
	notech_inv i_15526(.A(clk), .Z(n_62280));
	notech_inv i_15524(.A(n_62215), .Z(n_62278));
	notech_inv i_15522(.A(n_62215), .Z(n_62276));
	notech_inv i_15519(.A(n_62215), .Z(n_62273));
	notech_inv i_15517(.A(n_62215), .Z(n_62271));
	notech_inv i_15514(.A(n_62215), .Z(n_62268));
	notech_inv i_15512(.A(n_62215), .Z(n_62266));
	notech_inv i_15508(.A(n_62215), .Z(n_62262));
	notech_inv i_15506(.A(n_62215), .Z(n_62260));
	notech_inv i_15503(.A(n_62215), .Z(n_62257));
	notech_inv i_15501(.A(n_62215), .Z(n_62255));
	notech_inv i_15498(.A(n_62215), .Z(n_62252));
	notech_inv i_15496(.A(n_62215), .Z(n_62250));
	notech_inv i_15492(.A(n_62215), .Z(n_62246));
	notech_inv i_15490(.A(n_62215), .Z(n_62244));
	notech_inv i_15487(.A(n_62215), .Z(n_62241));
	notech_inv i_15485(.A(n_62215), .Z(n_62239));
	notech_inv i_15482(.A(n_62215), .Z(n_62236));
	notech_inv i_15480(.A(n_62215), .Z(n_62234));
	notech_inv i_15476(.A(n_62217), .Z(n_62230));
	notech_inv i_15474(.A(n_62217), .Z(n_62228));
	notech_inv i_15471(.A(n_62217), .Z(n_62225));
	notech_inv i_15469(.A(n_62217), .Z(n_62223));
	notech_inv i_15466(.A(n_62217), .Z(n_62220));
	notech_inv i_15464(.A(n_62217), .Z(n_62218));
	notech_inv i_15463(.A(n_62239), .Z(n_62217));
	notech_inv i_15461(.A(clk), .Z(n_62215));
	notech_inv i_15459(.A(n_62150), .Z(n_62213));
	notech_inv i_15457(.A(n_62150), .Z(n_62211));
	notech_inv i_15454(.A(n_62150), .Z(n_62208));
	notech_inv i_15452(.A(n_62150), .Z(n_62206));
	notech_inv i_15449(.A(n_62150), .Z(n_62203));
	notech_inv i_15447(.A(n_62150), .Z(n_62201));
	notech_inv i_15443(.A(n_62150), .Z(n_62197));
	notech_inv i_15441(.A(n_62150), .Z(n_62195));
	notech_inv i_15438(.A(n_62150), .Z(n_62192));
	notech_inv i_15436(.A(n_62150), .Z(n_62190));
	notech_inv i_15433(.A(n_62150), .Z(n_62187));
	notech_inv i_15431(.A(n_62150), .Z(n_62185));
	notech_inv i_15427(.A(n_62150), .Z(n_62181));
	notech_inv i_15425(.A(n_62150), .Z(n_62179));
	notech_inv i_15422(.A(n_62150), .Z(n_62176));
	notech_inv i_15420(.A(n_62150), .Z(n_62174));
	notech_inv i_15417(.A(n_62150), .Z(n_62171));
	notech_inv i_15415(.A(n_62150), .Z(n_62169));
	notech_inv i_15411(.A(n_62152), .Z(n_62165));
	notech_inv i_15409(.A(n_62152), .Z(n_62163));
	notech_inv i_15406(.A(n_62152), .Z(n_62160));
	notech_inv i_15404(.A(n_62152), .Z(n_62158));
	notech_inv i_15401(.A(n_62152), .Z(n_62155));
	notech_inv i_15399(.A(n_62152), .Z(n_62153));
	notech_inv i_15398(.A(n_62174), .Z(n_62152));
	notech_inv i_15396(.A(clk), .Z(n_62150));
	notech_inv i_14743(.A(n_61732), .Z(n_61796));
	notech_inv i_14741(.A(n_61732), .Z(n_61794));
	notech_inv i_14740(.A(n_61732), .Z(n_61793));
	notech_inv i_14736(.A(n_61732), .Z(n_61789));
	notech_inv i_14735(.A(n_61732), .Z(n_61788));
	notech_inv i_14731(.A(n_61732), .Z(n_61784));
	notech_inv i_14730(.A(n_61732), .Z(n_61783));
	notech_inv i_14726(.A(n_61732), .Z(n_61779));
	notech_inv i_14724(.A(n_61732), .Z(n_61777));
	notech_inv i_14721(.A(n_61732), .Z(n_61774));
	notech_inv i_14719(.A(n_61732), .Z(n_61772));
	notech_inv i_14716(.A(n_61732), .Z(n_61769));
	notech_inv i_14714(.A(n_61732), .Z(n_61767));
	notech_inv i_14710(.A(n_61732), .Z(n_61763));
	notech_inv i_14708(.A(n_61732), .Z(n_61761));
	notech_inv i_14705(.A(n_61732), .Z(n_61758));
	notech_inv i_14703(.A(n_61732), .Z(n_61756));
	notech_inv i_14700(.A(n_61732), .Z(n_61753));
	notech_inv i_14698(.A(n_61732), .Z(n_61751));
	notech_inv i_14694(.A(n_61734), .Z(n_61747));
	notech_inv i_14692(.A(n_61734), .Z(n_61745));
	notech_inv i_14689(.A(n_61734), .Z(n_61742));
	notech_inv i_14687(.A(n_61734), .Z(n_61740));
	notech_inv i_14684(.A(n_61734), .Z(n_61737));
	notech_inv i_14682(.A(n_61734), .Z(n_61735));
	notech_inv i_14681(.A(n_61751), .Z(n_61734));
	notech_inv i_14679(.A(rstn), .Z(n_61732));
	notech_inv i_14677(.A(n_61667), .Z(n_61730));
	notech_inv i_14675(.A(n_61667), .Z(n_61728));
	notech_inv i_14672(.A(n_61667), .Z(n_61725));
	notech_inv i_14670(.A(n_61667), .Z(n_61723));
	notech_inv i_14667(.A(n_61667), .Z(n_61720));
	notech_inv i_14665(.A(n_61667), .Z(n_61718));
	notech_inv i_14661(.A(n_61667), .Z(n_61714));
	notech_inv i_14659(.A(n_61667), .Z(n_61712));
	notech_inv i_14656(.A(n_61667), .Z(n_61709));
	notech_inv i_14654(.A(n_61667), .Z(n_61707));
	notech_inv i_14651(.A(n_61667), .Z(n_61704));
	notech_inv i_14649(.A(n_61667), .Z(n_61702));
	notech_inv i_14645(.A(n_61667), .Z(n_61698));
	notech_inv i_14643(.A(n_61667), .Z(n_61696));
	notech_inv i_14640(.A(n_61667), .Z(n_61693));
	notech_inv i_14638(.A(n_61667), .Z(n_61691));
	notech_inv i_14635(.A(n_61667), .Z(n_61688));
	notech_inv i_14633(.A(n_61667), .Z(n_61686));
	notech_inv i_14629(.A(n_61669), .Z(n_61682));
	notech_inv i_14627(.A(n_61669), .Z(n_61680));
	notech_inv i_14624(.A(n_61669), .Z(n_61677));
	notech_inv i_14622(.A(n_61669), .Z(n_61675));
	notech_inv i_14619(.A(n_61669), .Z(n_61672));
	notech_inv i_14617(.A(n_61669), .Z(n_61670));
	notech_inv i_14616(.A(n_61691), .Z(n_61669));
	notech_inv i_14614(.A(rstn), .Z(n_61667));
	notech_inv i_14612(.A(n_61602), .Z(n_61665));
	notech_inv i_14610(.A(n_61602), .Z(n_61663));
	notech_inv i_14607(.A(n_61602), .Z(n_61660));
	notech_inv i_14605(.A(n_61602), .Z(n_61658));
	notech_inv i_14602(.A(n_61602), .Z(n_61655));
	notech_inv i_14600(.A(n_61602), .Z(n_61653));
	notech_inv i_14596(.A(n_61602), .Z(n_61649));
	notech_inv i_14594(.A(n_61602), .Z(n_61647));
	notech_inv i_14591(.A(n_61602), .Z(n_61644));
	notech_inv i_14589(.A(n_61602), .Z(n_61642));
	notech_inv i_14586(.A(n_61602), .Z(n_61639));
	notech_inv i_14584(.A(n_61602), .Z(n_61637));
	notech_inv i_14580(.A(n_61602), .Z(n_61633));
	notech_inv i_14578(.A(n_61602), .Z(n_61631));
	notech_inv i_14575(.A(n_61602), .Z(n_61628));
	notech_inv i_14573(.A(n_61602), .Z(n_61626));
	notech_inv i_14570(.A(n_61602), .Z(n_61623));
	notech_inv i_14568(.A(n_61602), .Z(n_61621));
	notech_inv i_14564(.A(n_61604), .Z(n_61617));
	notech_inv i_14562(.A(n_61604), .Z(n_61615));
	notech_inv i_14559(.A(n_61604), .Z(n_61612));
	notech_inv i_14557(.A(n_61604), .Z(n_61610));
	notech_inv i_14554(.A(n_61604), .Z(n_61607));
	notech_inv i_14552(.A(n_61604), .Z(n_61605));
	notech_inv i_14551(.A(n_61626), .Z(n_61604));
	notech_inv i_14549(.A(rstn), .Z(n_61602));
	notech_inv i_14055(.A(n_61033), .Z(n_61098));
	notech_inv i_14054(.A(n_61033), .Z(n_61097));
	notech_inv i_14049(.A(n_61033), .Z(n_61092));
	notech_inv i_14044(.A(n_61033), .Z(n_61087));
	notech_inv i_14043(.A(n_61033), .Z(n_61086));
	notech_inv i_14038(.A(n_61033), .Z(n_61081));
	notech_inv i_14033(.A(n_61033), .Z(n_61076));
	notech_inv i_14032(.A(n_61033), .Z(n_61075));
	notech_inv i_14027(.A(n_61033), .Z(n_61070));
	notech_inv i_14021(.A(n_61033), .Z(n_61064));
	notech_inv i_14020(.A(n_61033), .Z(n_61063));
	notech_inv i_14015(.A(n_61033), .Z(n_61058));
	notech_inv i_14010(.A(n_61033), .Z(n_61053));
	notech_inv i_14009(.A(n_61033), .Z(n_61052));
	notech_inv i_14004(.A(n_61033), .Z(n_61047));
	notech_inv i_13999(.A(n_61033), .Z(n_61042));
	notech_inv i_13998(.A(n_61033), .Z(n_61041));
	notech_inv i_13993(.A(n_61033), .Z(n_61036));
	notech_inv i_13990(.A(term), .Z(n_61033));
	notech_inv i_13987(.A(n_60999), .Z(n_61030));
	notech_inv i_13986(.A(n_60999), .Z(n_61029));
	notech_inv i_13981(.A(n_60999), .Z(n_61024));
	notech_inv i_13976(.A(n_60999), .Z(n_61019));
	notech_inv i_13975(.A(n_60999), .Z(n_61018));
	notech_inv i_13970(.A(n_60999), .Z(n_61013));
	notech_inv i_13965(.A(n_60999), .Z(n_61008));
	notech_inv i_13964(.A(n_60999), .Z(n_61007));
	notech_inv i_13959(.A(n_60999), .Z(n_61002));
	notech_inv i_13956(.A(term), .Z(n_60999));
	notech_inv i_13105(.A(n_60052), .Z(n_60068));
	notech_inv i_13103(.A(n_60052), .Z(n_60066));
	notech_inv i_13102(.A(n_60052), .Z(n_60065));
	notech_inv i_13098(.A(n_60052), .Z(n_60061));
	notech_inv i_13096(.A(n_60052), .Z(n_60059));
	notech_inv i_13093(.A(n_60052), .Z(n_60056));
	notech_inv i_13091(.A(n_60052), .Z(n_60054));
	notech_inv i_13090(.A(n_60052), .Z(n_60053));
	notech_inv i_13089(.A(n_274294699), .Z(n_60052));
	notech_inv i_13080(.A(n_60041), .Z(n_60042));
	notech_inv i_13079(.A(n_2226), .Z(n_60041));
	notech_inv i_13076(.A(n_59972), .Z(n_60037));
	notech_inv i_13075(.A(n_59972), .Z(n_60036));
	notech_inv i_13070(.A(n_59972), .Z(n_60031));
	notech_inv i_13065(.A(n_59972), .Z(n_60026));
	notech_inv i_13064(.A(n_59972), .Z(n_60025));
	notech_inv i_13059(.A(n_59972), .Z(n_60020));
	notech_inv i_13054(.A(n_59972), .Z(n_60015));
	notech_inv i_13053(.A(n_59972), .Z(n_60014));
	notech_inv i_13048(.A(n_59972), .Z(n_60009));
	notech_inv i_13042(.A(n_59972), .Z(n_60003));
	notech_inv i_13041(.A(n_59972), .Z(n_60002));
	notech_inv i_13036(.A(n_59972), .Z(n_59997));
	notech_inv i_13031(.A(n_59972), .Z(n_59992));
	notech_inv i_13030(.A(n_59972), .Z(n_59991));
	notech_inv i_13025(.A(n_59972), .Z(n_59986));
	notech_inv i_13020(.A(n_59972), .Z(n_59981));
	notech_inv i_13019(.A(n_59972), .Z(n_59980));
	notech_inv i_13014(.A(n_59972), .Z(n_59975));
	notech_inv i_13011(.A(n_40926), .Z(n_59972));
	notech_inv i_13008(.A(n_59938), .Z(n_59969));
	notech_inv i_13007(.A(n_59938), .Z(n_59968));
	notech_inv i_13002(.A(n_59938), .Z(n_59963));
	notech_inv i_12996(.A(n_59938), .Z(n_59957));
	notech_inv i_12991(.A(n_59938), .Z(n_59952));
	notech_inv i_12985(.A(n_59938), .Z(n_59946));
	notech_inv i_12980(.A(n_59938), .Z(n_59941));
	notech_inv i_12977(.A(n_40926), .Z(n_59938));
	notech_inv i_12755(.A(n_59650), .Z(n_59704));
	notech_inv i_12754(.A(n_59650), .Z(n_59703));
	notech_inv i_12750(.A(n_59650), .Z(n_59699));
	notech_inv i_12746(.A(n_59650), .Z(n_59695));
	notech_inv i_12745(.A(n_59650), .Z(n_59694));
	notech_inv i_12741(.A(n_59650), .Z(n_59690));
	notech_inv i_12737(.A(n_59650), .Z(n_59686));
	notech_inv i_12736(.A(n_59650), .Z(n_59685));
	notech_inv i_12732(.A(n_59650), .Z(n_59681));
	notech_inv i_12727(.A(n_59650), .Z(n_59676));
	notech_inv i_12726(.A(n_59650), .Z(n_59675));
	notech_inv i_12722(.A(n_59650), .Z(n_59671));
	notech_inv i_12718(.A(n_59650), .Z(n_59667));
	notech_inv i_12717(.A(n_59650), .Z(n_59666));
	notech_inv i_12713(.A(n_59650), .Z(n_59662));
	notech_inv i_12709(.A(n_59650), .Z(n_59658));
	notech_inv i_12708(.A(n_59650), .Z(n_59657));
	notech_inv i_12704(.A(n_59650), .Z(n_59653));
	notech_inv i_12701(.A(n_5770), .Z(n_59650));
	notech_inv i_12699(.A(n_59622), .Z(n_59648));
	notech_inv i_12698(.A(n_59622), .Z(n_59647));
	notech_inv i_12694(.A(n_59622), .Z(n_59643));
	notech_inv i_12685(.A(n_59633), .Z(n_59634));
	notech_inv i_12684(.A(n_59632), .Z(n_59633));
	notech_inv i_12683(.A(n_59622), .Z(n_59632));
	notech_inv i_12676(.A(n_59624), .Z(n_59625));
	notech_inv i_12675(.A(n_59623), .Z(n_59624));
	notech_inv i_12674(.A(n_59622), .Z(n_59623));
	notech_inv i_12673(.A(n_5770), .Z(n_59622));
	notech_inv i_12671(.A(n_59531), .Z(n_59619));
	notech_inv i_12669(.A(n_59531), .Z(n_59617));
	notech_inv i_12666(.A(n_59531), .Z(n_59614));
	notech_inv i_12664(.A(n_59531), .Z(n_59612));
	notech_inv i_12660(.A(n_59531), .Z(n_59608));
	notech_inv i_12658(.A(n_59531), .Z(n_59606));
	notech_inv i_12655(.A(n_59531), .Z(n_59603));
	notech_inv i_12653(.A(n_59531), .Z(n_59601));
	notech_inv i_12649(.A(n_59531), .Z(n_59597));
	notech_inv i_12647(.A(n_59531), .Z(n_59595));
	notech_inv i_12644(.A(n_59531), .Z(n_59592));
	notech_inv i_12642(.A(n_59531), .Z(n_59590));
	notech_inv i_12638(.A(n_59531), .Z(n_59586));
	notech_inv i_12636(.A(n_59531), .Z(n_59584));
	notech_inv i_12633(.A(n_59531), .Z(n_59581));
	notech_inv i_12631(.A(n_59531), .Z(n_59579));
	notech_inv i_12626(.A(n_59566), .Z(n_59574));
	notech_inv i_12624(.A(n_59566), .Z(n_59572));
	notech_inv i_12621(.A(n_59566), .Z(n_59569));
	notech_inv i_12619(.A(n_59566), .Z(n_59567));
	notech_inv i_12618(.A(n_59612), .Z(n_59566));
	notech_inv i_12615(.A(n_59566), .Z(n_59563));
	notech_inv i_12613(.A(n_59566), .Z(n_59561));
	notech_inv i_12610(.A(n_59566), .Z(n_59558));
	notech_inv i_12608(.A(n_59566), .Z(n_59556));
	notech_inv i_12604(.A(n_59566), .Z(n_59552));
	notech_inv i_12602(.A(n_59566), .Z(n_59550));
	notech_inv i_12599(.A(n_59566), .Z(n_59547));
	notech_inv i_12597(.A(n_59566), .Z(n_59545));
	notech_inv i_12593(.A(n_59531), .Z(n_59541));
	notech_inv i_12591(.A(n_59531), .Z(n_59539));
	notech_inv i_12588(.A(n_59531), .Z(n_59536));
	notech_inv i_12586(.A(n_59531), .Z(n_59534));
	notech_inv i_12583(.A(n_5769), .Z(n_59531));
	notech_inv i_12581(.A(n_59486), .Z(n_59529));
	notech_inv i_12579(.A(n_59486), .Z(n_59527));
	notech_inv i_12576(.A(n_59486), .Z(n_59524));
	notech_inv i_12574(.A(n_59486), .Z(n_59522));
	notech_inv i_12570(.A(n_59486), .Z(n_59518));
	notech_inv i_12568(.A(n_59486), .Z(n_59516));
	notech_inv i_12565(.A(n_59486), .Z(n_59513));
	notech_inv i_12563(.A(n_59486), .Z(n_59511));
	notech_inv i_12559(.A(n_59486), .Z(n_59507));
	notech_inv i_12557(.A(n_59486), .Z(n_59505));
	notech_inv i_12554(.A(n_59486), .Z(n_59502));
	notech_inv i_12552(.A(n_59486), .Z(n_59500));
	notech_inv i_12548(.A(n_59486), .Z(n_59496));
	notech_inv i_12546(.A(n_59486), .Z(n_59494));
	notech_inv i_12542(.A(n_59486), .Z(n_59490));
	notech_inv i_12538(.A(n_5769), .Z(n_59486));
	notech_inv i_12134(.A(n_59075), .Z(n_59091));
	notech_inv i_12132(.A(n_59075), .Z(n_59089));
	notech_inv i_12131(.A(n_59075), .Z(n_59088));
	notech_inv i_12127(.A(n_59075), .Z(n_59084));
	notech_inv i_12125(.A(n_59075), .Z(n_59082));
	notech_inv i_12122(.A(n_59075), .Z(n_59079));
	notech_inv i_12120(.A(n_59075), .Z(n_59077));
	notech_inv i_12119(.A(n_59075), .Z(n_59076));
	notech_inv i_12118(.A(n_5768), .Z(n_59075));
	notech_inv i_12111(.A(n_59066), .Z(n_59067));
	notech_inv i_12110(.A(n_3185), .Z(n_59066));
	notech_inv i_12108(.A(n_59045), .Z(n_59063));
	notech_inv i_12106(.A(n_59045), .Z(n_59061));
	notech_inv i_12103(.A(n_59045), .Z(n_59058));
	notech_inv i_12101(.A(n_59045), .Z(n_59056));
	notech_inv i_12098(.A(n_59045), .Z(n_59053));
	notech_inv i_12096(.A(n_59045), .Z(n_59051));
	notech_inv i_12093(.A(n_59045), .Z(n_59048));
	notech_inv i_12091(.A(n_59045), .Z(n_59046));
	notech_inv i_12090(.A(n_3184), .Z(n_59045));
	notech_inv i_12083(.A(n_59036), .Z(n_59037));
	notech_inv i_12082(.A(n_3273), .Z(n_59036));
	notech_inv i_12075(.A(n_59027), .Z(n_59028));
	notech_inv i_12074(.A(n_1448), .Z(n_59027));
	notech_inv i_12070(.A(n_1953), .Z(n_59022));
	notech_inv i_12065(.A(n_1953), .Z(n_59017));
	notech_inv i_12062(.A(n_58997), .Z(n_59013));
	notech_inv i_12060(.A(n_58997), .Z(n_59011));
	notech_inv i_12059(.A(n_58997), .Z(n_59010));
	notech_inv i_12055(.A(n_58997), .Z(n_59006));
	notech_inv i_12053(.A(n_58997), .Z(n_59004));
	notech_inv i_12050(.A(n_58997), .Z(n_59001));
	notech_inv i_12048(.A(n_58997), .Z(n_58999));
	notech_inv i_12047(.A(n_58997), .Z(n_58998));
	notech_inv i_12046(.A(n_5276), .Z(n_58997));
	notech_inv i_12041(.A(n_58990), .Z(n_58991));
	notech_inv i_12040(.A(fpu), .Z(n_58990));
	notech_inv i_11540(.A(n_58450), .Z(n_58452));
	notech_inv i_11539(.A(n_58450), .Z(n_58451));
	notech_inv i_11538(.A(in128[10]), .Z(n_58450));
	notech_inv i_11448(.A(n_58284), .Z(n_58349));
	notech_inv i_11447(.A(n_58284), .Z(n_58348));
	notech_inv i_11442(.A(n_58284), .Z(n_58343));
	notech_inv i_11437(.A(n_58284), .Z(n_58338));
	notech_inv i_11436(.A(n_58284), .Z(n_58337));
	notech_inv i_11431(.A(n_58284), .Z(n_58332));
	notech_inv i_11426(.A(n_58284), .Z(n_58327));
	notech_inv i_11425(.A(n_58284), .Z(n_58326));
	notech_inv i_11420(.A(n_58284), .Z(n_58321));
	notech_inv i_11414(.A(n_58284), .Z(n_58315));
	notech_inv i_11413(.A(n_58284), .Z(n_58314));
	notech_inv i_11408(.A(n_58284), .Z(n_58309));
	notech_inv i_11403(.A(n_58284), .Z(n_58304));
	notech_inv i_11402(.A(n_58284), .Z(n_58303));
	notech_inv i_11397(.A(n_58284), .Z(n_58298));
	notech_inv i_11392(.A(n_58284), .Z(n_58293));
	notech_inv i_11391(.A(n_58284), .Z(n_58292));
	notech_inv i_11386(.A(n_58284), .Z(n_58287));
	notech_inv i_11383(.A(\nbus_13540[0] ), .Z(n_58284));
	notech_inv i_11380(.A(n_58250), .Z(n_58281));
	notech_inv i_11379(.A(n_58250), .Z(n_58280));
	notech_inv i_11369(.A(n_58250), .Z(n_58270));
	notech_inv i_11368(.A(n_58250), .Z(n_58269));
	notech_inv i_11363(.A(n_58250), .Z(n_58264));
	notech_inv i_11358(.A(n_58250), .Z(n_58259));
	notech_inv i_11357(.A(n_58250), .Z(n_58258));
	notech_inv i_11352(.A(n_58250), .Z(n_58253));
	notech_inv i_11349(.A(\nbus_13540[0] ), .Z(n_58250));
	notech_inv i_11347(.A(n_58159), .Z(n_58247));
	notech_inv i_11345(.A(n_58159), .Z(n_58245));
	notech_inv i_11342(.A(n_58159), .Z(n_58242));
	notech_inv i_11340(.A(n_58159), .Z(n_58240));
	notech_inv i_11336(.A(n_58159), .Z(n_58236));
	notech_inv i_11334(.A(n_58159), .Z(n_58234));
	notech_inv i_11331(.A(n_58159), .Z(n_58231));
	notech_inv i_11329(.A(n_58159), .Z(n_58229));
	notech_inv i_11325(.A(n_58159), .Z(n_58225));
	notech_inv i_11323(.A(n_58159), .Z(n_58223));
	notech_inv i_11320(.A(n_58159), .Z(n_58220));
	notech_inv i_11318(.A(n_58159), .Z(n_58218));
	notech_inv i_11314(.A(n_58159), .Z(n_58214));
	notech_inv i_11312(.A(n_58159), .Z(n_58212));
	notech_inv i_11309(.A(n_58159), .Z(n_58209));
	notech_inv i_11307(.A(n_58159), .Z(n_58207));
	notech_inv i_11302(.A(n_58194), .Z(n_58202));
	notech_inv i_11300(.A(n_58194), .Z(n_58200));
	notech_inv i_11297(.A(n_58194), .Z(n_58197));
	notech_inv i_11295(.A(n_58194), .Z(n_58195));
	notech_inv i_11294(.A(n_58240), .Z(n_58194));
	notech_inv i_11291(.A(n_58194), .Z(n_58191));
	notech_inv i_11289(.A(n_58194), .Z(n_58189));
	notech_inv i_11286(.A(n_58194), .Z(n_58186));
	notech_inv i_11284(.A(n_58194), .Z(n_58184));
	notech_inv i_11280(.A(n_58194), .Z(n_58180));
	notech_inv i_11278(.A(n_58194), .Z(n_58178));
	notech_inv i_11275(.A(n_58194), .Z(n_58175));
	notech_inv i_11273(.A(n_58194), .Z(n_58173));
	notech_inv i_11269(.A(n_58159), .Z(n_58169));
	notech_inv i_11267(.A(n_58159), .Z(n_58167));
	notech_inv i_11264(.A(n_58159), .Z(n_58164));
	notech_inv i_11262(.A(n_58159), .Z(n_58162));
	notech_inv i_11259(.A(n_5630), .Z(n_58159));
	notech_inv i_11257(.A(n_58114), .Z(n_58157));
	notech_inv i_11255(.A(n_58114), .Z(n_58155));
	notech_inv i_11252(.A(n_58114), .Z(n_58152));
	notech_inv i_11250(.A(n_58114), .Z(n_58150));
	notech_inv i_11246(.A(n_58114), .Z(n_58146));
	notech_inv i_11244(.A(n_58114), .Z(n_58144));
	notech_inv i_11241(.A(n_58114), .Z(n_58141));
	notech_inv i_11239(.A(n_58114), .Z(n_58139));
	notech_inv i_11235(.A(n_58114), .Z(n_58135));
	notech_inv i_11233(.A(n_58114), .Z(n_58133));
	notech_inv i_11229(.A(n_58114), .Z(n_58129));
	notech_inv i_11223(.A(n_58114), .Z(n_58123));
	notech_inv i_11222(.A(n_58114), .Z(n_58122));
	notech_inv i_11217(.A(n_58114), .Z(n_58117));
	notech_inv i_11214(.A(n_5630), .Z(n_58114));
	notech_inv i_10449(.A(n_57100), .Z(n_57101));
	notech_inv i_10448(.A(n_2884), .Z(n_57100));
	notech_inv i_9082(.A(n_55754), .Z(n_55755));
	notech_inv i_9081(.A(n_162496319), .Z(n_55754));
	notech_inv i_9072(.A(n_55743), .Z(n_55744));
	notech_inv i_9071(.A(\nbus_13535[0] ), .Z(n_55743));
	notech_inv i_9045(.A(n_55716), .Z(n_55717));
	notech_inv i_9044(.A(\nbus_13534[0] ), .Z(n_55716));
	notech_inv i_9040(.A(n_55716), .Z(n_55712));
	notech_inv i_9036(.A(n_55716), .Z(n_55708));
	notech_inv i_9031(.A(n_55716), .Z(n_55703));
	notech_inv i_9027(.A(n_55716), .Z(n_55699));
	notech_inv i_9017(.A(n_55688), .Z(n_55689));
	notech_inv i_9016(.A(n_55669), .Z(n_55688));
	notech_inv i_9012(.A(n_55688), .Z(n_55684));
	notech_inv i_9008(.A(n_55688), .Z(n_55680));
	notech_inv i_9003(.A(n_55688), .Z(n_55675));
	notech_inv i_8999(.A(n_55688), .Z(n_55671));
	notech_inv i_8997(.A(n_55716), .Z(n_55669));
	notech_inv i_8989(.A(n_55660), .Z(n_55661));
	notech_inv i_8988(.A(n_55641), .Z(n_55660));
	notech_inv i_8984(.A(n_55660), .Z(n_55656));
	notech_inv i_8980(.A(n_55660), .Z(n_55652));
	notech_inv i_8975(.A(n_55660), .Z(n_55647));
	notech_inv i_8971(.A(n_55660), .Z(n_55643));
	notech_inv i_8969(.A(n_55716), .Z(n_55641));
	notech_inv i_8466(.A(n_55058), .Z(n_55123));
	notech_inv i_8465(.A(n_55058), .Z(n_55122));
	notech_inv i_8460(.A(n_55058), .Z(n_55117));
	notech_inv i_8455(.A(n_55058), .Z(n_55112));
	notech_inv i_8454(.A(n_55058), .Z(n_55111));
	notech_inv i_8449(.A(n_55058), .Z(n_55106));
	notech_inv i_8444(.A(n_55058), .Z(n_55101));
	notech_inv i_8443(.A(n_55058), .Z(n_55100));
	notech_inv i_8438(.A(n_55058), .Z(n_55095));
	notech_inv i_8432(.A(n_55058), .Z(n_55089));
	notech_inv i_8431(.A(n_55058), .Z(n_55088));
	notech_inv i_8426(.A(n_55058), .Z(n_55083));
	notech_inv i_8421(.A(n_55058), .Z(n_55078));
	notech_inv i_8420(.A(n_55058), .Z(n_55077));
	notech_inv i_8415(.A(n_55058), .Z(n_55072));
	notech_inv i_8410(.A(n_55058), .Z(n_55067));
	notech_inv i_8409(.A(n_55058), .Z(n_55066));
	notech_inv i_8404(.A(n_55058), .Z(n_55061));
	notech_inv i_8401(.A(\nbus_13541[0] ), .Z(n_55058));
	notech_inv i_8398(.A(n_55024), .Z(n_55055));
	notech_inv i_8397(.A(n_55024), .Z(n_55054));
	notech_inv i_8387(.A(n_55024), .Z(n_55044));
	notech_inv i_8386(.A(n_55024), .Z(n_55043));
	notech_inv i_8381(.A(n_55024), .Z(n_55038));
	notech_inv i_8376(.A(n_55024), .Z(n_55033));
	notech_inv i_8375(.A(n_55024), .Z(n_55032));
	notech_inv i_8370(.A(n_55024), .Z(n_55027));
	notech_inv i_8367(.A(\nbus_13541[0] ), .Z(n_55024));
	notech_inv i_7962(.A(n_54628), .Z(n_54629));
	notech_inv i_7961(.A(n_40487), .Z(n_54628));
	notech_inv i_7943(.A(n_54556), .Z(n_54557));
	notech_inv i_7942(.A(n_3123), .Z(n_54556));
	notech_ao4 i_2627697(.A(n_2122), .B(n_59579), .C(n_58207), .D(n_39285), 
		.Z(n_3282));
	notech_ao4 i_1727688(.A(n_2125), .B(n_59574), .C(n_58207), .D(n_39272), 
		.Z(n_3283));
	notech_ao4 i_1527686(.A(n_2126), .B(n_59579), .C(n_58207), .D(n_39269), 
		.Z(n_3284));
	notech_ao4 i_12725521(.A(n_59579), .B(n_40721), .C(n_58207), .D(n_39612)
		, .Z(n_3285));
	notech_ao4 i_12625520(.A(n_59579), .B(n_40720), .C(n_58207), .D(n_39610)
		, .Z(n_3286));
	notech_ao4 i_12525519(.A(n_59574), .B(n_40719), .C(n_58202), .D(n_39609)
		, .Z(n_3287));
	notech_ao4 i_12425518(.A(n_59574), .B(n_40718), .C(n_58202), .D(n_39607)
		, .Z(n_3288));
	notech_ao4 i_12325517(.A(n_59574), .B(n_40717), .C(n_58202), .D(n_39606)
		, .Z(n_3289));
	notech_ao4 i_12225516(.A(n_59574), .B(n_40716), .C(n_58207), .D(n_39604)
		, .Z(n_3290));
	notech_ao4 i_12125515(.A(n_59574), .B(n_40715), .C(n_58207), .D(n_39603)
		, .Z(n_3291));
	notech_ao4 i_12025514(.A(n_59579), .B(n_40714), .C(n_58207), .D(n_39601)
		, .Z(n_3292));
	notech_ao4 i_11925513(.A(n_59579), .B(n_40713), .C(n_58207), .D(n_39600)
		, .Z(n_3293));
	notech_ao4 i_11825512(.A(n_59579), .B(n_40712), .C(n_58209), .D(n_39598)
		, .Z(n_3294));
	notech_ao4 i_11725511(.A(n_59579), .B(n_40711), .C(n_58209), .D(n_39597)
		, .Z(n_3295));
	notech_ao4 i_11625510(.A(n_59579), .B(n_40710), .C(n_58209), .D(n_39595)
		, .Z(n_3296));
	notech_ao4 i_11525509(.A(n_59579), .B(n_40709), .C(n_58207), .D(n_39594)
		, .Z(n_3297));
	notech_ao4 i_11425508(.A(n_59579), .B(n_40708), .C(n_58207), .D(n_39592)
		, .Z(n_3298));
	notech_ao4 i_11325507(.A(n_59579), .B(n_40707), .C(n_58207), .D(n_39591)
		, .Z(n_3299));
	notech_ao4 i_11225506(.A(n_59579), .B(n_40706), .C(n_58207), .D(n_39589)
		, .Z(n_3300));
	notech_ao4 i_11125505(.A(n_59579), .B(n_40705), .C(n_58207), .D(n_39588)
		, .Z(n_3301));
	notech_ao3 i_3403(.A(n_60009), .B(udeco[110]), .C(n_59681), .Z(n_3302)
		);
	notech_ao4 i_11025504(.A(n_59574), .B(n_40704), .C(n_58202), .D(n_39586)
		, .Z(n_3303));
	notech_ao4 i_10925503(.A(n_59572), .B(n_40703), .C(n_58200), .D(n_39585)
		, .Z(n_3304));
	notech_ao4 i_10825502(.A(n_59572), .B(n_40702), .C(n_58200), .D(n_39583)
		, .Z(n_3305));
	notech_ao3 i_3400(.A(n_60009), .B(udeco[107]), .C(n_59681), .Z(n_3306)
		);
	notech_ao4 i_10725501(.A(n_59572), .B(n_40701), .C(n_58200), .D(n_39582)
		, .Z(n_3307));
	notech_ao4 i_10625500(.A(n_59572), .B(n_40700), .C(n_58200), .D(n_39580)
		, .Z(n_3308));
	notech_ao4 i_10525499(.A(n_59572), .B(n_40699), .C(n_58200), .D(n_39579)
		, .Z(n_3309));
	notech_ao4 i_10425498(.A(n_59572), .B(n_40698), .C(n_58200), .D(n_39577)
		, .Z(n_3310));
	notech_ao4 i_10325497(.A(n_59572), .B(n_40697), .C(n_58200), .D(n_39575)
		, .Z(n_3311));
	notech_ao4 i_10225496(.A(n_59572), .B(n_40696), .C(n_58200), .D(n_39573)
		, .Z(n_3312));
	notech_ao4 i_10125495(.A(n_59572), .B(n_40695), .C(n_58200), .D(n_39572)
		, .Z(n_3313));
	notech_ao4 i_10025494(.A(n_59572), .B(n_40694), .C(n_58200), .D(n_39570)
		, .Z(n_3314));
	notech_ao4 i_9925493(.A(n_59574), .B(n_40693), .C(n_58202), .D(n_39569),
		 .Z(n_3315));
	notech_ao4 i_9825492(.A(n_59574), .B(n_40692), .C(n_58202), .D(n_39567),
		 .Z(n_3316));
	notech_ao4 i_9725491(.A(n_59574), .B(n_40691), .C(n_58202), .D(n_39566),
		 .Z(n_3317));
	notech_ao4 i_9625490(.A(n_59574), .B(n_40690), .C(n_58202), .D(n_39564),
		 .Z(n_3318));
	notech_ao4 i_9525489(.A(n_59574), .B(n_40689), .C(n_58202), .D(n_39563),
		 .Z(n_3319));
	notech_ao4 i_9425488(.A(n_59572), .B(n_40688), .C(n_58202), .D(n_39561),
		 .Z(n_3320));
	notech_ao4 i_9325487(.A(n_59572), .B(n_40687), .C(n_58202), .D(n_39560),
		 .Z(n_3321));
	notech_ao4 i_9225486(.A(n_59572), .B(n_40686), .C(n_58202), .D(n_39558),
		 .Z(n_3322));
	notech_ao4 i_9125485(.A(n_59574), .B(n_40685), .C(n_58202), .D(n_39557),
		 .Z(n_3323));
	notech_ao4 i_9025484(.A(n_59574), .B(n_40684), .C(n_58202), .D(n_39555),
		 .Z(n_3324));
	notech_ao4 i_8925483(.A(n_59581), .B(n_40683), .C(n_58214), .D(n_39554),
		 .Z(n_3325));
	notech_ao3 i_3382(.A(n_60009), .B(udeco[88]), .C(n_59681), .Z(n_3326));
	notech_ao4 i_8825482(.A(n_59586), .B(n_40682), .C(n_58214), .D(n_39552),
		 .Z(n_3327));
	notech_ao4 i_8725481(.A(n_59584), .B(n_40681), .C(n_58214), .D(n_39551),
		 .Z(n_3328));
	notech_ao3 i_3380(.A(n_60009), .B(udeco[86]), .C(n_59681), .Z(n_3329));
	notech_ao4 i_8625480(.A(n_59586), .B(n_40680), .C(n_58214), .D(n_39549),
		 .Z(n_3330));
	notech_ao4 i_8525479(.A(n_59586), .B(n_40679), .C(n_58214), .D(n_39548),
		 .Z(n_3331));
	notech_ao3 i_3378(.A(n_60009), .B(udeco[84]), .C(n_59681), .Z(n_3332));
	notech_ao4 i_8425478(.A(n_59586), .B(n_40678), .C(n_58212), .D(n_39546),
		 .Z(n_3333));
	notech_ao4 i_8325477(.A(n_59584), .B(n_40677), .C(n_58212), .D(n_39545),
		 .Z(n_3334));
	notech_ao4 i_8225476(.A(n_59584), .B(n_40676), .C(n_58212), .D(n_39543),
		 .Z(n_3335));
	notech_ao4 i_8125475(.A(n_59584), .B(n_40675), .C(n_58214), .D(n_39542),
		 .Z(n_3336));
	notech_ao4 i_8025474(.A(n_59584), .B(n_40674), .C(n_58212), .D(n_39540),
		 .Z(n_3337));
	notech_ao4 i_7925473(.A(n_59584), .B(n_40673), .C(n_58214), .D(n_39539),
		 .Z(n_3338));
	notech_ao4 i_7825472(.A(n_59586), .B(n_40672), .C(n_58214), .D(n_39537),
		 .Z(n_3339));
	notech_ao4 i_7725471(.A(n_59586), .B(n_40671), .C(n_58214), .D(n_39536),
		 .Z(n_3340));
	notech_ao4 i_7625470(.A(n_59586), .B(n_40670), .C(n_58218), .D(n_39534),
		 .Z(n_3341));
	notech_ao4 i_7525469(.A(n_59586), .B(n_40669), .C(n_58218), .D(n_39533),
		 .Z(n_3342));
	notech_ao4 i_7425468(.A(n_59586), .B(n_40668), .C(n_58214), .D(n_39531),
		 .Z(n_3343));
	notech_ao4 i_7325467(.A(n_59586), .B(n_40667), .C(n_58214), .D(n_39530),
		 .Z(n_3344));
	notech_ao4 i_7225466(.A(n_59586), .B(n_40666), .C(n_58214), .D(n_39528),
		 .Z(n_3345));
	notech_ao4 i_7125465(.A(n_59586), .B(n_40665), .C(n_58214), .D(n_39527),
		 .Z(n_3346));
	notech_ao4 i_7025464(.A(n_59586), .B(n_40664), .C(n_58214), .D(n_39525),
		 .Z(n_3347));
	notech_ao4 i_6925463(.A(n_59586), .B(n_40663), .C(n_58212), .D(n_39524),
		 .Z(n_3348));
	notech_ao4 i_6825462(.A(n_59584), .B(n_40662), .C(n_58209), .D(n_39522),
		 .Z(n_3349));
	notech_ao3 i_3361(.A(n_60009), .B(udeco[67]), .C(n_59681), .Z(n_3350));
	notech_ao4 i_6725461(.A(n_59581), .B(n_40661), .C(n_58209), .D(n_39521),
		 .Z(n_3351));
	notech_ao3 i_3360(.A(n_60009), .B(udeco[66]), .C(n_59681), .Z(n_3352));
	notech_ao4 i_6625460(.A(n_59581), .B(n_40660), .C(n_58209), .D(n_39519),
		 .Z(n_3353));
	notech_ao3 i_3359(.A(n_60014), .B(udeco[65]), .C(n_59681), .Z(n_3354));
	notech_ao4 i_6525459(.A(n_59581), .B(n_40659), .C(n_58209), .D(n_39518),
		 .Z(n_3355));
	notech_ao3 i_3358(.A(n_60014), .B(udeco[64]), .C(n_59681), .Z(n_3356));
	notech_ao4 i_6425458(.A(n_59581), .B(n_40658), .C(n_58209), .D(n_39516),
		 .Z(n_3357));
	notech_ao3 i_3357(.A(n_60009), .B(udeco[63]), .C(n_59681), .Z(n_3358));
	notech_ao4 i_6325457(.A(n_59581), .B(n_40657), .C(n_58209), .D(n_39515),
		 .Z(n_3359));
	notech_ao3 i_3356(.A(n_60009), .B(udeco[62]), .C(n_59681), .Z(n_3360));
	notech_ao4 i_6225456(.A(n_59581), .B(n_40656), .C(n_58209), .D(n_39513),
		 .Z(n_3361));
	notech_ao3 i_3355(.A(n_60009), .B(udeco[61]), .C(n_59676), .Z(n_3362));
	notech_ao4 i_6125455(.A(n_59581), .B(n_40655), .C(n_58209), .D(n_39512),
		 .Z(n_3363));
	notech_ao3 i_3354(.A(n_60009), .B(udeco[60]), .C(n_59676), .Z(n_3364));
	notech_ao4 i_6025454(.A(n_59581), .B(n_40654), .C(n_58209), .D(n_39510),
		 .Z(n_3365));
	notech_ao3 i_3353(.A(n_60003), .B(udeco[59]), .C(n_59676), .Z(n_3366));
	notech_ao4 i_5925453(.A(n_59581), .B(n_40653), .C(n_58209), .D(n_39509),
		 .Z(n_3367));
	notech_ao3 i_3352(.A(n_60003), .B(udeco[58]), .C(n_59676), .Z(n_3368));
	notech_ao4 i_5825452(.A(n_59581), .B(n_40652), .C(n_58212), .D(n_39507),
		 .Z(n_3369));
	notech_ao3 i_3351(.A(n_60003), .B(udeco[57]), .C(n_59676), .Z(n_3370));
	notech_ao4 i_5725451(.A(n_59584), .B(n_40651), .C(n_58212), .D(n_39506),
		 .Z(n_3371));
	notech_ao3 i_3350(.A(n_60003), .B(udeco[56]), .C(n_59676), .Z(n_3372));
	notech_ao4 i_5625450(.A(n_59584), .B(n_40650), .C(n_58212), .D(n_39504),
		 .Z(n_3373));
	notech_ao3 i_3349(.A(n_60003), .B(udeco[55]), .C(n_59676), .Z(n_3374));
	notech_ao4 i_5525449(.A(n_59584), .B(n_40649), .C(n_58212), .D(n_39503),
		 .Z(n_3375));
	notech_ao3 i_3348(.A(n_60003), .B(udeco[54]), .C(n_59681), .Z(n_3376));
	notech_ao4 i_5425448(.A(n_59584), .B(n_40648), .C(n_58212), .D(n_39501),
		 .Z(n_3377));
	notech_ao3 i_3347(.A(n_60003), .B(udeco[53]), .C(n_59676), .Z(n_3378));
	notech_ao4 i_5325447(.A(n_59584), .B(n_40647), .C(n_58212), .D(n_39500),
		 .Z(n_3379));
	notech_ao3 i_3346(.A(n_60003), .B(udeco[52]), .C(n_59676), .Z(n_3380));
	notech_ao4 i_5225446(.A(n_59581), .B(n_40646), .C(n_58209), .D(n_39498),
		 .Z(n_3381));
	notech_ao3 i_3345(.A(n_60009), .B(udeco[51]), .C(n_59676), .Z(n_3382));
	notech_ao4 i_5125445(.A(n_59581), .B(n_40645), .C(n_58212), .D(n_39497),
		 .Z(n_3383));
	notech_ao3 i_3344(.A(n_60003), .B(udeco[50]), .C(n_59681), .Z(n_3384));
	notech_ao4 i_5025444(.A(n_59581), .B(n_40644), .C(n_58212), .D(n_39495),
		 .Z(n_3385));
	notech_ao3 i_3343(.A(n_60003), .B(udeco[49]), .C(n_59685), .Z(n_3386));
	notech_ao4 i_4925443(.A(n_59584), .B(n_40643), .C(n_58212), .D(n_39494),
		 .Z(n_3387));
	notech_ao3 i_3342(.A(n_60003), .B(udeco[48]), .C(n_59686), .Z(n_3388));
	notech_ao4 i_4825442(.A(n_59584), .B(n_40642), .C(n_58200), .D(n_39492),
		 .Z(n_3389));
	notech_ao3 i_3341(.A(n_60014), .B(udeco[47]), .C(n_59685), .Z(n_3390));
	notech_ao4 i_4725441(.A(n_59572), .B(n_40641), .C(n_58189), .D(n_39491),
		 .Z(n_3391));
	notech_ao3 i_3340(.A(n_60015), .B(udeco[46]), .C(n_59685), .Z(n_3392));
	notech_ao4 i_4625440(.A(n_59561), .B(n_40640), .C(n_58189), .D(n_39489),
		 .Z(n_3393));
	notech_ao3 i_3339(.A(n_60015), .B(udeco[45]), .C(n_59685), .Z(n_3394));
	notech_ao4 i_4525439(.A(n_59558), .B(n_40639), .C(n_58189), .D(n_39488),
		 .Z(n_3395));
	notech_ao3 i_3338(.A(n_60015), .B(udeco[44]), .C(n_59686), .Z(n_3396));
	notech_ao4 i_4425438(.A(n_59561), .B(n_40638), .C(n_58189), .D(n_39486),
		 .Z(n_3397));
	notech_ao3 i_3337(.A(n_60014), .B(udeco[43]), .C(n_59686), .Z(n_3398));
	notech_ao4 i_4325437(.A(n_59561), .B(n_40637), .C(n_58189), .D(n_39485),
		 .Z(n_3399));
	notech_ao3 i_3336(.A(n_60014), .B(udeco[42]), .C(n_59686), .Z(n_3400));
	notech_ao4 i_4225436(.A(n_59561), .B(n_40636), .C(n_58186), .D(n_39483),
		 .Z(n_3401));
	notech_ao3 i_3335(.A(n_60015), .B(udeco[41]), .C(n_59686), .Z(n_3402));
	notech_ao4 i_4125435(.A(n_59558), .B(n_40635), .C(n_58186), .D(n_39482),
		 .Z(n_3403));
	notech_ao3 i_3334(.A(n_60015), .B(udeco[40]), .C(n_59686), .Z(n_3404));
	notech_ao4 i_4025434(.A(n_59558), .B(n_40634), .C(n_58189), .D(n_39480),
		 .Z(n_3405));
	notech_ao3 i_3333(.A(n_60015), .B(udeco[39]), .C(n_59686), .Z(n_3406));
	notech_ao4 i_3925433(.A(n_59558), .B(n_40633), .C(n_58189), .D(n_39479),
		 .Z(n_3407));
	notech_ao3 i_3332(.A(n_60015), .B(udeco[38]), .C(n_59685), .Z(n_3408));
	notech_ao4 i_3725431(.A(n_59558), .B(n_40631), .C(n_58189), .D(n_39476),
		 .Z(n_3409));
	notech_ao3 i_3330(.A(n_60015), .B(udeco[36]), .C(n_59685), .Z(n_3410));
	notech_ao4 i_3625430(.A(n_59558), .B(n_40630), .C(n_58191), .D(n_39474),
		 .Z(n_3411));
	notech_ao3 i_3329(.A(n_60015), .B(udeco[35]), .C(n_59685), .Z(n_3412));
	notech_ao4 i_3525429(.A(n_59561), .B(n_40629), .C(n_58189), .D(n_39473),
		 .Z(n_3413));
	notech_ao3 i_3328(.A(n_60015), .B(udeco[34]), .C(n_59681), .Z(n_3414));
	notech_ao4 i_3425428(.A(n_59561), .B(n_40628), .C(n_58191), .D(n_39471),
		 .Z(n_3415));
	notech_ao3 i_3327(.A(n_60014), .B(udeco[33]), .C(n_59685), .Z(n_3416));
	notech_ao4 i_3225426(.A(n_59561), .B(n_40626), .C(n_58191), .D(n_39468),
		 .Z(n_3417));
	notech_ao3 i_3325(.A(n_60014), .B(udeco[31]), .C(n_59685), .Z(n_3418));
	notech_ao4 i_3125425(.A(n_59561), .B(n_40625), .C(n_58191), .D(n_39467),
		 .Z(n_3419));
	notech_ao3 i_3324(.A(n_60014), .B(udeco[30]), .C(n_59685), .Z(n_3420));
	notech_ao4 i_3025424(.A(n_59561), .B(n_40624), .C(n_58189), .D(n_39465),
		 .Z(n_3421));
	notech_ao3 i_3323(.A(n_60014), .B(udeco[29]), .C(n_59685), .Z(n_3422));
	notech_ao4 i_2925423(.A(n_59561), .B(n_40623), .C(n_58189), .D(n_39464),
		 .Z(n_3423));
	notech_ao3 i_3322(.A(n_60014), .B(udeco[28]), .C(n_59685), .Z(n_3424));
	notech_ao4 i_2825422(.A(n_59561), .B(n_40622), .C(n_58189), .D(n_39462),
		 .Z(n_3425));
	notech_ao3 i_3321(.A(n_60014), .B(udeco[27]), .C(n_59685), .Z(n_3426));
	notech_ao4 i_2725421(.A(n_59561), .B(n_40621), .C(n_58189), .D(n_39461),
		 .Z(n_3427));
	notech_ao3 i_3320(.A(n_60014), .B(udeco[26]), .C(n_59685), .Z(n_3428));
	notech_ao4 i_2225416(.A(n_59561), .B(n_40616), .C(n_58189), .D(n_39453),
		 .Z(n_3429));
	notech_ao4 i_2125415(.A(n_59561), .B(n_40615), .C(n_58186), .D(n_39452),
		 .Z(n_3430));
	notech_ao3 i_3314(.A(n_60014), .B(udeco[20]), .C(n_59676), .Z(n_3431));
	notech_ao4 i_2025414(.A(n_59558), .B(n_40614), .C(n_58184), .D(n_39450),
		 .Z(n_3432));
	notech_ao4 i_1825412(.A(n_59556), .B(n_40612), .C(n_58184), .D(n_39447),
		 .Z(n_3433));
	notech_ao4 i_1725411(.A(n_59556), .B(n_40611), .C(n_58184), .D(n_39446),
		 .Z(n_3434));
	notech_ao3 i_3310(.A(n_60014), .B(udeco[16]), .C(n_59671), .Z(n_3435));
	notech_ao4 i_1625410(.A(n_59556), .B(n_40610), .C(n_58186), .D(n_39444),
		 .Z(n_3436));
	notech_ao4 i_1525409(.A(n_59556), .B(n_40609), .C(n_58184), .D(n_39443),
		 .Z(n_3437));
	notech_ao4 i_1425408(.A(n_59556), .B(n_40608), .C(n_58184), .D(n_39441),
		 .Z(n_3438));
	notech_ao4 i_1325407(.A(n_59556), .B(n_40607), .C(n_58184), .D(n_39440),
		 .Z(n_3439));
	notech_ao3 i_3306(.A(n_60014), .B(udeco[12]), .C(n_59671), .Z(n_3440));
	notech_ao4 i_1225406(.A(n_59556), .B(n_40606), .C(n_58184), .D(n_39438),
		 .Z(n_3441));
	notech_ao4 i_1125405(.A(n_59556), .B(n_40605), .C(n_58184), .D(n_39437),
		 .Z(n_3442));
	notech_ao4 i_1025404(.A(n_59556), .B(n_40604), .C(n_58184), .D(n_39435),
		 .Z(n_3443));
	notech_ao4 i_925403(.A(n_59556), .B(n_40603), .C(n_58186), .D(n_39434), 
		.Z(n_3444));
	notech_ao4 i_825402(.A(n_59558), .B(n_40602), .C(n_58186), .D(n_39432), 
		.Z(n_3445));
	notech_ao4 i_725401(.A(n_59558), .B(n_40601), .C(n_58186), .D(n_39431), 
		.Z(n_3446));
	notech_ao4 i_625400(.A(n_59558), .B(n_40600), .C(n_58186), .D(n_39429), 
		.Z(n_3447));
	notech_ao4 i_525399(.A(n_59558), .B(n_40599), .C(n_58186), .D(n_39428), 
		.Z(n_3448));
	notech_ao4 i_425398(.A(n_59558), .B(n_40598), .C(n_58186), .D(n_39426), 
		.Z(n_3449));
	notech_ao4 i_325397(.A(n_59556), .B(n_40597), .C(n_58186), .D(n_39425), 
		.Z(n_3450));
	notech_ao4 i_225396(.A(n_59556), .B(n_40596), .C(n_58186), .D(n_39423), 
		.Z(n_3451));
	notech_ao4 i_125395(.A(n_59556), .B(n_40595), .C(n_58186), .D(n_39422), 
		.Z(n_3452));
	notech_ao4 i_21126328(.A(n_59558), .B(n_40838), .C(n_58186), .D(n_40171)
		, .Z(n_3453));
	notech_ao4 i_3627707(.A(n_3123), .B(n_40312), .C(n_58197), .D(n_39300), 
		.Z(n_3281));
	notech_ao4 i_21026327(.A(n_59558), .B(n_40837), .C(n_58197), .D(n_40170)
		, .Z(n_3454));
	notech_ao3 i_11574039(.A(n_60014), .B(in128[126]), .C(n_59667), .Z(n_48392
		));
	notech_ao4 i_20926326(.A(n_59563), .B(n_40836), .C(n_58197), .D(n_40168)
		, .Z(n_3455));
	notech_ao3 i_11674038(.A(n_60014), .B(in128[125]), .C(n_59667), .Z(n_48386
		));
	notech_ao4 i_20826325(.A(n_59569), .B(n_40835), .C(n_58197), .D(n_40167)
		, .Z(n_3456));
	notech_ao4 i_20726324(.A(n_59567), .B(n_40834), .C(n_58197), .D(n_40165)
		, .Z(n_3457));
	notech_ao3 i_11874036(.A(n_60014), .B(in128[123]), .C(n_59667), .Z(n_48374
		));
	notech_ao4 i_20626323(.A(n_59569), .B(n_40833), .C(n_58195), .D(n_40164)
		, .Z(n_3458));
	notech_ao4 i_20526322(.A(n_59569), .B(n_40832), .C(n_58195), .D(n_40162)
		, .Z(n_3459));
	notech_ao3 i_12074034(.A(n_60003), .B(in128[121]), .C(n_59671), .Z(n_48362
		));
	notech_ao4 i_20426321(.A(n_59569), .B(n_40831), .C(n_58195), .D(n_40161)
		, .Z(n_3460));
	notech_ao3 i_12174033(.A(n_59997), .B(in128[120]), .C(n_59671), .Z(n_3461
		));
	notech_ao4 i_20326320(.A(n_59567), .B(n_40830), .C(n_58197), .D(n_40159)
		, .Z(n_3462));
	notech_ao3 i_12274032(.A(n_59997), .B(in128[119]), .C(n_59671), .Z(n_3463
		));
	notech_ao4 i_20226319(.A(n_59567), .B(n_40829), .C(n_58197), .D(n_40158)
		, .Z(n_3464));
	notech_ao3 i_12374031(.A(n_59997), .B(in128[118]), .C(n_59671), .Z(n_3465
		));
	notech_ao4 i_20126318(.A(n_59567), .B(n_40828), .C(n_58197), .D(n_40156)
		, .Z(n_3466));
	notech_ao3 i_12474030(.A(n_59992), .B(in128[117]), .C(n_59671), .Z(n_3467
		));
	notech_ao4 i_20026317(.A(n_59567), .B(n_40827), .C(n_58197), .D(n_40155)
		, .Z(n_3468));
	notech_ao3 i_12574029(.A(n_59992), .B(in128[116]), .C(n_59671), .Z(n_3469
		));
	notech_ao4 i_19926316(.A(n_59567), .B(n_40826), .C(n_58200), .D(n_40153)
		, .Z(n_3470));
	notech_ao3 i_12674028(.A(n_59997), .B(in128[115]), .C(n_59667), .Z(n_3471
		));
	notech_ao4 i_19826315(.A(n_59569), .B(n_40825), .C(n_58200), .D(n_40152)
		, .Z(n_3472));
	notech_ao3 i_12774027(.A(n_59997), .B(in128[114]), .C(n_59667), .Z(n_3473
		));
	notech_ao4 i_19726314(.A(n_59569), .B(n_40824), .C(n_58200), .D(n_40150)
		, .Z(n_3474));
	notech_ao3 i_12874026(.A(n_59997), .B(in128[113]), .C(n_59667), .Z(n_3475
		));
	notech_ao4 i_19526312(.A(n_59569), .B(n_40822), .C(n_58197), .D(n_40147)
		, .Z(n_3476));
	notech_ao3 i_12974025(.A(n_59997), .B(in128[111]), .C(n_59667), .Z(n_3477
		));
	notech_ao4 i_19426311(.A(n_59569), .B(n_40821), .C(n_58197), .D(n_40146)
		, .Z(n_3478));
	notech_ao3 i_13074024(.A(n_59997), .B(in128[110]), .C(n_59667), .Z(n_3479
		));
	notech_ao4 i_19326310(.A(n_59569), .B(n_40820), .C(n_58197), .D(n_40144)
		, .Z(n_3480));
	notech_ao3 i_13174023(.A(n_59997), .B(in128[109]), .C(n_59667), .Z(n_3481
		));
	notech_ao4 i_19226309(.A(n_59569), .B(n_40819), .C(n_58197), .D(n_40143)
		, .Z(n_3482));
	notech_ao3 i_13274022(.A(n_59997), .B(in128[108]), .C(n_59667), .Z(n_3483
		));
	notech_ao4 i_19126308(.A(n_59569), .B(n_40818), .C(n_58197), .D(n_40141)
		, .Z(n_3484));
	notech_ao3 i_13374021(.A(n_59992), .B(in128[107]), .C(n_59667), .Z(n_3485
		));
	notech_ao4 i_19026307(.A(n_59569), .B(n_40817), .C(n_58195), .D(n_40140)
		, .Z(n_3486));
	notech_ao3 i_13474020(.A(n_59992), .B(in128[106]), .C(n_59667), .Z(n_3487
		));
	notech_ao4 i_18926306(.A(n_59569), .B(n_40816), .C(n_58191), .D(n_40138)
		, .Z(n_3488));
	notech_ao3 i_13574019(.A(n_59992), .B(in128[105]), .C(n_59667), .Z(n_3489
		));
	notech_ao4 i_18826305(.A(n_59569), .B(n_40815), .C(n_58191), .D(n_40137)
		, .Z(n_3490));
	notech_ao3 i_13674018(.A(n_59992), .B(in128[104]), .C(n_59667), .Z(n_3491
		));
	notech_ao4 i_18726304(.A(n_59567), .B(n_40814), .C(n_58191), .D(n_40135)
		, .Z(n_3492));
	notech_ao3 i_13774017(.A(n_59992), .B(in128[103]), .C(n_59671), .Z(n_3493
		));
	notech_ao4 i_18626303(.A(n_59563), .B(n_40813), .C(n_58191), .D(n_40134)
		, .Z(n_3494));
	notech_ao3 i_13874016(.A(n_59992), .B(in128[102]), .C(n_59675), .Z(n_3495
		));
	notech_ao4 i_18526302(.A(n_59563), .B(n_40812), .C(n_58191), .D(n_40132)
		, .Z(n_3496));
	notech_ao3 i_13974015(.A(n_59992), .B(in128[101]), .C(n_59675), .Z(n_3497
		));
	notech_ao4 i_18426301(.A(n_59563), .B(n_40811), .C(n_58191), .D(n_40131)
		, .Z(n_3498));
	notech_ao3 i_14074014(.A(n_59992), .B(in128[100]), .C(n_59675), .Z(n_3499
		));
	notech_ao4 i_18326300(.A(n_59563), .B(n_40810), .C(n_58191), .D(n_40129)
		, .Z(n_3500));
	notech_ao3 i_14174013(.A(n_59992), .B(in128[99]), .C(n_59675), .Z(n_3501
		));
	notech_ao4 i_18226299(.A(n_59563), .B(n_40809), .C(n_58191), .D(n_40128)
		, .Z(n_3502));
	notech_ao3 i_14274012(.A(n_59992), .B(in128[98]), .C(n_59675), .Z(n_3503
		));
	notech_ao4 i_18026297(.A(n_59563), .B(n_40807), .C(n_58191), .D(n_40125)
		, .Z(n_3504));
	notech_ao3 i_14374011(.A(n_59992), .B(in128[96]), .C(n_59675), .Z(n_3505
		));
	notech_ao4 i_17926296(.A(n_59563), .B(n_40806), .C(n_58191), .D(n_40123)
		, .Z(n_3506));
	notech_ao3 i_14474010(.A(n_59992), .B(in128[95]), .C(n_59676), .Z(n_3507
		));
	notech_ao4 i_17826295(.A(n_59563), .B(n_40805), .C(n_58195), .D(n_40122)
		, .Z(n_3508));
	notech_ao3 i_14574009(.A(n_59992), .B(in128[94]), .C(n_59676), .Z(n_3509
		));
	notech_ao4 i_17726294(.A(n_59563), .B(n_40804), .C(n_58195), .D(n_40120)
		, .Z(n_3510));
	notech_ao4 i_17626293(.A(n_59563), .B(n_40803), .C(n_58195), .D(n_40119)
		, .Z(n_3511));
	notech_ao3 i_14674008(.A(n_59997), .B(in128[92]), .C(n_59676), .Z(n_3512
		));
	notech_ao4 i_17526292(.A(n_59567), .B(n_40802), .C(n_58195), .D(n_40117)
		, .Z(n_3513));
	notech_ao3 i_14774007(.A(n_60002), .B(in128[91]), .C(n_59675), .Z(n_3514
		));
	notech_ao4 i_17426291(.A(n_59567), .B(n_40801), .C(n_58195), .D(n_40116)
		, .Z(n_3515));
	notech_ao3 i_14874006(.A(n_60002), .B(in128[90]), .C(n_59675), .Z(n_3516
		));
	notech_ao4 i_17326290(.A(n_59567), .B(n_40800), .C(n_58195), .D(n_40114)
		, .Z(n_3517));
	notech_ao4 i_17226289(.A(n_59567), .B(n_40799), .C(n_58195), .D(n_40113)
		, .Z(n_3518));
	notech_ao3 i_14974005(.A(n_60002), .B(in128[88]), .C(n_59671), .Z(n_3519
		));
	notech_ao4 i_17126288(.A(n_59567), .B(n_40798), .C(n_58195), .D(n_40111)
		, .Z(n_3520));
	notech_ao3 i_5674098(.A(n_60002), .B(in128[87]), .C(n_59671), .Z(n_3521)
		);
	notech_ao4 i_17026287(.A(n_59563), .B(n_40797), .C(n_58195), .D(n_40110)
		, .Z(n_3522));
	notech_ao3 i_4574109(.A(n_60002), .B(in128[86]), .C(n_59671), .Z(n_3523)
		);
	notech_ao4 i_16926286(.A(n_59563), .B(n_40796), .C(n_58195), .D(n_40109)
		, .Z(n_3524));
	notech_ao4 i_16826285(.A(n_59563), .B(n_40795), .C(n_58218), .D(n_40108)
		, .Z(n_3525));
	notech_ao3 i_4674108(.A(n_60002), .B(in128[84]), .C(n_59671), .Z(n_3526)
		);
	notech_ao4 i_16726284(.A(n_58240), .B(n_40107), .C(n_59567), .D(n_40794)
		, .Z(n_3527));
	notech_ao4 i_16626283(.A(n_58240), .B(n_40106), .C(n_59567), .D(n_40793)
		, .Z(n_3528));
	notech_ao4 i_16326280(.A(n_59590), .B(n_40790), .C(n_58240), .D(n_40103)
		, .Z(n_3529));
	notech_ao4 i_16226279(.A(n_59612), .B(n_40789), .C(n_58240), .D(n_40102)
		, .Z(n_3530));
	notech_ao4 i_16126278(.A(n_59608), .B(n_40788), .C(n_58240), .D(n_40101)
		, .Z(n_3531));
	notech_ao4 i_16026277(.A(n_59612), .B(n_40787), .C(n_58236), .D(n_40100)
		, .Z(n_3532));
	notech_ao4 i_15926276(.A(n_59612), .B(n_40786), .C(n_58236), .D(n_40099)
		, .Z(n_3533));
	notech_ao3 i_4874106(.A(n_60003), .B(in128[75]), .C(n_59671), .Z(n_3534)
		);
	notech_ao4 i_15826275(.A(n_59612), .B(n_40785), .C(n_58236), .D(n_40098)
		, .Z(n_3535));
	notech_ao4 i_15626273(.A(n_59608), .B(n_40783), .C(n_58236), .D(n_40096)
		, .Z(n_3536));
	notech_ao4 i_15526272(.A(n_59608), .B(n_40782), .C(n_58236), .D(n_40095)
		, .Z(n_3537));
	notech_ao4 i_15426271(.A(n_59608), .B(n_40781), .C(n_58240), .D(n_40094)
		, .Z(n_3538));
	notech_ao4 i_15026267(.A(n_59608), .B(n_40777), .C(n_58240), .D(n_40090)
		, .Z(n_3539));
	notech_ao4 i_14926266(.A(n_59608), .B(n_40776), .C(n_58240), .D(n_40089)
		, .Z(n_3540));
	notech_ao4 i_14826265(.A(n_59612), .B(n_40775), .C(n_58242), .D(n_40088)
		, .Z(n_3541));
	notech_ao4 i_14726264(.A(n_59612), .B(n_40774), .C(n_58240), .D(n_40087)
		, .Z(n_3542));
	notech_ao4 i_14626263(.A(n_59612), .B(n_40773), .C(n_58240), .D(n_40086)
		, .Z(n_3543));
	notech_ao4 i_14526262(.A(n_59612), .B(n_40772), .C(n_58240), .D(n_40084)
		, .Z(n_3544));
	notech_ao4 i_14426261(.A(n_59612), .B(n_40771), .C(n_58240), .D(n_40083)
		, .Z(n_3545));
	notech_ao4 i_14326260(.A(n_59612), .B(n_40770), .C(n_58240), .D(n_40081)
		, .Z(n_3546));
	notech_ao4 i_14226259(.A(n_59612), .B(n_40769), .C(n_58240), .D(n_40080)
		, .Z(n_3547));
	notech_ao4 i_14126258(.A(n_59612), .B(n_40768), .C(n_58236), .D(n_40079)
		, .Z(n_3548));
	notech_ao4 i_14026257(.A(n_59612), .B(n_40767), .C(n_58234), .D(n_40078)
		, .Z(n_3549));
	notech_ao4 i_13926256(.A(n_59612), .B(n_40766), .C(n_58234), .D(n_40077)
		, .Z(n_3550));
	notech_ao4 i_13826255(.A(n_59608), .B(n_40765), .C(n_58234), .D(n_40076)
		, .Z(n_3551));
	notech_ao4 i_13726254(.A(n_59606), .B(n_40764), .C(n_58234), .D(n_40075)
		, .Z(n_3552));
	notech_ao4 i_13626253(.A(n_59606), .B(n_40763), .C(n_58234), .D(n_40074)
		, .Z(n_3553));
	notech_ao4 i_13526252(.A(n_59606), .B(n_40762), .C(n_58234), .D(n_40072)
		, .Z(n_3554));
	notech_ao4 i_13426251(.A(n_59606), .B(n_40761), .C(n_58234), .D(n_40071)
		, .Z(n_3555));
	notech_ao4 i_13326250(.A(n_59606), .B(n_40760), .C(n_58234), .D(n_40069)
		, .Z(n_3556));
	notech_ao4 i_13226249(.A(n_59606), .B(n_40759), .C(n_58234), .D(n_40068)
		, .Z(n_3557));
	notech_ao4 i_13126248(.A(n_59606), .B(n_40758), .C(n_58234), .D(n_40066)
		, .Z(n_3558));
	notech_ao4 i_13026247(.A(n_59606), .B(n_40757), .C(n_58236), .D(n_40065)
		, .Z(n_3559));
	notech_ao4 i_12926246(.A(n_59606), .B(n_40756), .C(n_58236), .D(n_40063)
		, .Z(n_3560));
	notech_ao4 i_12826245(.A(n_59606), .B(n_40755), .C(n_58236), .D(n_40062)
		, .Z(n_3561));
	notech_ao4 i_12726244(.A(n_59608), .B(n_40754), .C(n_58236), .D(n_40060)
		, .Z(n_3562));
	notech_ao4 i_12626243(.A(n_59608), .B(n_40753), .C(n_58236), .D(n_40059)
		, .Z(n_3563));
	notech_ao4 i_12426241(.A(n_59608), .B(n_40751), .C(n_58234), .D(n_40056)
		, .Z(n_3564));
	notech_ao4 i_12326240(.A(n_59608), .B(n_40750), .C(n_58234), .D(n_40054)
		, .Z(n_3565));
	notech_ao4 i_12226239(.A(n_59608), .B(n_40749), .C(n_58236), .D(n_40053)
		, .Z(n_3566));
	notech_ao4 i_12026237(.A(n_59606), .B(n_40747), .C(n_58236), .D(n_40050)
		, .Z(n_3567));
	notech_ao4 i_11426231(.A(n_59606), .B(n_40741), .C(n_58236), .D(n_40041)
		, .Z(n_3568));
	notech_ao4 i_11326230(.A(n_59606), .B(n_40740), .C(n_58247), .D(n_40039)
		, .Z(n_3569));
	notech_ao4 i_11226229(.A(n_59608), .B(n_40739), .C(n_58245), .D(n_40038)
		, .Z(n_3570));
	notech_ao4 i_11126228(.A(n_59608), .B(n_40738), .C(n_58247), .D(n_40036)
		, .Z(n_3571));
	notech_ao4 i_11026227(.A(n_59614), .B(n_40737), .C(n_58247), .D(n_40035)
		, .Z(n_3572));
	notech_ao4 i_10826225(.A(n_59619), .B(n_40735), .C(n_58247), .D(n_40031)
		, .Z(n_3573));
	notech_ao4 i_9026207(.A(n_59617), .B(n_40856), .C(n_58245), .D(n_39996),
		 .Z(n_3574));
	notech_ao3 i_15174003(.A(n_60003), .B(in128[6]), .C(n_59675), .Z(n_3575)
		);
	notech_ao4 i_8926206(.A(n_59619), .B(n_40857), .C(n_58245), .D(n_39994),
		 .Z(n_3576));
	notech_ao3 i_15274002(.A(n_60003), .B(in128[5]), .C(n_59675), .Z(n_3577)
		);
	notech_ao4 i_8826205(.A(n_59619), .B(n_40858), .C(n_58245), .D(n_39993),
		 .Z(n_3578));
	notech_ao3 i_15374001(.A(n_60003), .B(in128[4]), .C(n_59675), .Z(n_3579)
		);
	notech_ao4 i_8726204(.A(n_59619), .B(n_40859), .C(n_58245), .D(n_39991),
		 .Z(n_3580));
	notech_ao3 i_15474000(.A(n_60003), .B(in128[3]), .C(n_59675), .Z(n_3581)
		);
	notech_ao4 i_8626203(.A(n_59617), .B(n_40918), .C(n_58245), .D(n_39990),
		 .Z(n_3582));
	notech_ao3 i_6374091(.A(n_60003), .B(in128[2]), .C(n_59675), .Z(n_3583)
		);
	notech_ao4 i_8426201(.A(n_59617), .B(n_40839), .C(n_58247), .D(n_39986),
		 .Z(n_3584));
	notech_ao3 i_5774097(.A(n_60002), .B(in128[0]), .C(n_59675), .Z(n_3585)
		);
	notech_ao4 i_8326200(.A(n_59617), .B(n_40920), .C(n_58247), .D(n_39984),
		 .Z(n_3586));
	notech_ao3 i_11374041(.A(n_60002), .B(mod_dec), .C(n_59699), .Z(n_3587)
		);
	notech_ao4 i_8226199(.A(n_59617), .B(n_40919), .C(n_58247), .D(n_39983),
		 .Z(n_3588));
	notech_ao3 i_11474040(.A(n_60002), .B(sib_dec), .C(n_59699), .Z(n_3589)
		);
	notech_ao4 i_8126198(.A(n_59617), .B(n_40873), .C(n_58247), .D(n_39981),
		 .Z(n_3590));
	notech_ao3 i_9574059(.A(n_60002), .B(\to_acu2_0[80] ), .C(n_59699), .Z(n_3591
		));
	notech_ao4 i_8026197(.A(n_59619), .B(n_40889), .C(n_58247), .D(n_39980),
		 .Z(n_3592));
	notech_ao3 i_9174063(.A(n_59997), .B(\to_acu2_0[79] ), .C(n_59699), .Z(n_3593
		));
	notech_ao4 i_7926196(.A(n_59619), .B(n_40891), .C(n_58247), .D(n_39978),
		 .Z(n_3594));
	notech_ao3 i_9074064(.A(n_60002), .B(\to_acu2_0[78] ), .C(n_59699), .Z(n_3595
		));
	notech_ao4 i_7826195(.A(n_59619), .B(n_40840), .C(n_58247), .D(n_39977),
		 .Z(n_3596));
	notech_ao3 i_15573999(.A(n_60002), .B(\to_acu2_0[77] ), .C(n_59699), .Z(n_3597
		));
	notech_ao4 i_7726194(.A(n_59619), .B(n_40862), .C(n_58247), .D(n_39975),
		 .Z(n_3598));
	notech_ao3 i_8974065(.A(n_60002), .B(\to_acu2_0[76] ), .C(n_59703), .Z(n_3599
		));
	notech_ao4 i_7626193(.A(n_59619), .B(n_40855), .C(n_58247), .D(n_39974),
		 .Z(n_3600));
	notech_ao3 i_9374061(.A(n_60002), .B(\to_acu2_0[75] ), .C(n_59703), .Z(n_3601
		));
	notech_ao4 i_7526192(.A(n_59619), .B(n_40865), .C(n_58247), .D(n_39972),
		 .Z(n_3602));
	notech_ao3 i_7074084(.A(n_60002), .B(\to_acu2_0[74] ), .C(n_59703), .Z(n_3603
		));
	notech_ao4 i_7426191(.A(n_59619), .B(n_40864), .C(n_58245), .D(n_39971),
		 .Z(n_3604));
	notech_ao3 i_6774087(.A(n_60002), .B(\to_acu2_0[73] ), .C(n_59703), .Z(n_3605
		));
	notech_ao4 i_7326190(.A(n_59619), .B(n_40863), .C(n_58242), .D(n_39969),
		 .Z(n_3606));
	notech_ao3 i_8874066(.A(n_60002), .B(\to_acu2_0[72] ), .C(n_59703), .Z(n_3607
		));
	notech_ao4 i_7226189(.A(n_59619), .B(n_40853), .C(n_58242), .D(n_39968),
		 .Z(n_3608));
	notech_ao3 i_5274102(.A(n_60002), .B(\to_acu2_0[71] ), .C(n_59699), .Z(n_3609
		));
	notech_ao4 i_7126188(.A(n_59619), .B(n_40854), .C(n_58242), .D(n_39966),
		 .Z(n_3610));
	notech_ao3 i_9274062(.A(n_60015), .B(\to_acu2_0[70] ), .C(n_59699), .Z(n_3611
		));
	notech_ao4 i_7026187(.A(n_59617), .B(n_40914), .C(n_58242), .D(n_39965),
		 .Z(n_3612));
	notech_ao3 i_10474050(.A(n_60036), .B(\to_acu2_0[69] ), .C(n_59695), .Z(n_3613
		));
	notech_ao4 i_6926186(.A(n_59614), .B(n_40906), .C(n_58242), .D(n_39963),
		 .Z(n_3614));
	notech_ao3 i_8774067(.A(n_60036), .B(\to_acu2_0[68] ), .C(n_59695), .Z(n_3615
		));
	notech_ao4 i_6826185(.A(n_59614), .B(n_40841), .C(n_58242), .D(n_39962),
		 .Z(n_3616));
	notech_ao3 i_15673998(.A(n_60036), .B(\to_acu2_0[67] ), .C(n_59695), .Z(n_3617
		));
	notech_ao4 i_6726184(.A(n_59614), .B(n_40842), .C(n_58242), .D(n_39960),
		 .Z(n_3618));
	notech_ao3 i_15773997(.A(n_60031), .B(\to_acu2_0[66] ), .C(n_59699), .Z(n_3619
		));
	notech_ao4 i_6626183(.A(n_59614), .B(n_40843), .C(n_58242), .D(n_39959),
		 .Z(n_3620));
	notech_ao3 i_15873996(.A(n_60031), .B(\to_acu2_0[65] ), .C(n_59699), .Z(n_3621
		));
	notech_ao4 i_6526182(.A(n_59614), .B(n_40844), .C(n_58242), .D(n_39957),
		 .Z(n_3622));
	notech_ao3 i_15973995(.A(n_60036), .B(\to_acu2_0[64] ), .C(n_59699), .Z(n_3623
		));
	notech_ao4 i_6426181(.A(n_59614), .B(n_40845), .C(n_58242), .D(n_39956),
		 .Z(n_3624));
	notech_ao3 i_16073994(.A(n_60036), .B(\to_acu2_0[63] ), .C(n_59699), .Z(n_3625
		));
	notech_ao4 i_6326180(.A(n_59614), .B(n_40913), .C(n_58245), .D(n_39954),
		 .Z(n_3626));
	notech_ao3 i_10574049(.A(n_60036), .B(\to_acu2_0[62] ), .C(n_59699), .Z(n_3627
		));
	notech_ao4 i_6226179(.A(n_59614), .B(n_40890), .C(n_58245), .D(n_39953),
		 .Z(n_3628));
	notech_ao3 i_8674068(.A(n_60036), .B(\to_acu2_0[61] ), .C(n_59699), .Z(n_3629
		));
	notech_ao4 i_6126178(.A(n_59614), .B(n_40846), .C(n_58245), .D(n_39951),
		 .Z(n_3630));
	notech_ao3 i_16173993(.A(n_60036), .B(\to_acu2_0[60] ), .C(n_59703), .Z(n_3631
		));
	notech_ao4 i_6026177(.A(n_59614), .B(n_40872), .C(n_58245), .D(n_39950),
		 .Z(n_3632));
	notech_ao3 i_8574069(.A(n_60036), .B(\to_acu2_0[59] ), .C(n_59704), .Z(n_3633
		));
	notech_ao4 i_5926176(.A(n_59617), .B(n_40921), .C(n_58245), .D(n_39948),
		 .Z(n_3634));
	notech_ao4 i_5826175(.A(n_59617), .B(n_40866), .C(n_58242), .D(n_39947),
		 .Z(n_3635));
	notech_ao3 i_7174083(.A(n_60036), .B(\to_acu2_0[57] ), .C(n_59704), .Z(n_3636
		));
	notech_ao4 i_5726174(.A(n_59617), .B(n_40860), .C(n_58242), .D(n_39945),
		 .Z(n_3637));
	notech_ao3 i_9474060(.A(n_60031), .B(\to_acu2_0[56] ), .C(n_59704), .Z(n_3638
		));
	notech_ao4 i_5626173(.A(n_59617), .B(n_40870), .C(n_58242), .D(n_39944),
		 .Z(n_3639));
	notech_ao3 i_4074114(.A(n_60031), .B(\to_acu2_0[55] ), .C(n_59704), .Z(n_3640
		));
	notech_ao4 i_5526172(.A(n_59617), .B(n_40871), .C(n_58245), .D(n_39942),
		 .Z(n_3641));
	notech_ao3 i_3574119(.A(n_60031), .B(\to_acu2_0[54] ), .C(n_59704), .Z(n_3642
		));
	notech_ao4 i_5426171(.A(n_59614), .B(n_40869), .C(n_58245), .D(n_39941),
		 .Z(n_3643));
	notech_ao3 i_6074094(.A(n_60031), .B(\to_acu2_0[53] ), .C(n_59704), .Z(n_3644
		));
	notech_ao4 i_5326170(.A(n_59614), .B(n_40867), .C(n_58234), .D(n_39939),
		 .Z(n_3645));
	notech_ao3 i_4974105(.A(n_60026), .B(\to_acu2_0[52] ), .C(n_59704), .Z(n_3646
		));
	notech_ao4 i_5226169(.A(n_59614), .B(n_40868), .C(n_58223), .D(n_39938),
		 .Z(n_3647));
	notech_ao3 i_6174093(.A(n_60026), .B(\to_acu2_0[51] ), .C(n_59704), .Z(n_3648
		));
	notech_ao4 i_5126168(.A(n_59617), .B(n_40861), .C(n_58223), .D(n_39936),
		 .Z(n_3649));
	notech_ao3 i_5974095(.A(n_60026), .B(\to_acu2_0[50] ), .C(n_59704), .Z(n_3650
		));
	notech_ao4 i_5026167(.A(n_59617), .B(n_40847), .C(n_58223), .D(n_39935),
		 .Z(n_3651));
	notech_ao3 i_16273992(.A(n_60031), .B(\to_acu2_0[49] ), .C(n_59704), .Z(n_3652
		));
	notech_ao4 i_4926166(.A(n_59606), .B(n_40874), .C(n_58223), .D(n_39933),
		 .Z(n_3653));
	notech_ao3 i_8474070(.A(n_60031), .B(\to_acu2_0[48] ), .C(n_59704), .Z(n_3654
		));
	notech_ao4 i_4826165(.A(n_59595), .B(n_40888), .C(n_58223), .D(n_39932),
		 .Z(n_3655));
	notech_ao3 i_6274092(.A(n_60031), .B(\to_acu2_0[47] ), .C(n_59703), .Z(n_3656
		));
	notech_ao4 i_4726164(.A(n_59592), .B(n_40886), .C(n_58220), .D(n_39930),
		 .Z(n_3657));
	notech_ao3 i_5074104(.A(n_60031), .B(\to_acu2_0[46] ), .C(n_59703), .Z(n_3658
		));
	notech_ao4 i_4626163(.A(n_59595), .B(n_40887), .C(n_58220), .D(n_39929),
		 .Z(n_3659));
	notech_ao3 i_4174113(.A(n_60031), .B(\to_acu2_0[45] ), .C(n_59703), .Z(n_3660
		));
	notech_ao4 i_4526162(.A(n_59595), .B(n_40885), .C(n_58220), .D(n_39927),
		 .Z(n_3661));
	notech_ao3 i_3674118(.A(n_60031), .B(\to_acu2_0[44] ), .C(n_59703), .Z(n_3662
		));
	notech_ao4 i_4426161(.A(n_59595), .B(n_40883), .C(n_58223), .D(n_39926),
		 .Z(n_3663));
	notech_ao3 i_3374121(.A(n_60036), .B(\to_acu2_0[43] ), .C(n_59703), .Z(n_3664
		));
	notech_ao4 i_4326160(.A(n_59592), .B(n_40884), .C(n_58220), .D(n_39924),
		 .Z(n_3665));
	notech_ao3 i_11274042(.A(n_60037), .B(\to_acu2_0[42] ), .C(n_59703), .Z(n_3666
		));
	notech_ao4 i_4226159(.A(n_59592), .B(n_40882), .C(n_58223), .D(n_39923),
		 .Z(n_3667));
	notech_ao3 i_2974125(.A(n_60037), .B(\to_acu2_0[41] ), .C(n_59704), .Z(n_3668
		));
	notech_ao4 i_4126158(.A(n_59592), .B(n_40880), .C(n_58223), .D(n_39921),
		 .Z(n_3669));
	notech_ao3 i_11174043(.A(n_60037), .B(\to_acu2_0[40] ), .C(n_59704), .Z(n_3670
		));
	notech_ao4 i_3926156(.A(n_59592), .B(n_40881), .C(n_58223), .D(n_39919),
		 .Z(n_3671));
	notech_ao3 i_11074044(.A(n_60037), .B(\to_acu2_0[38] ), .C(n_59704), .Z(n_3672
		));
	notech_ao4 i_3826155(.A(n_59592), .B(n_40878), .C(n_58225), .D(n_39918),
		 .Z(n_3673));
	notech_ao3 i_10974045(.A(n_60037), .B(\to_acu2_0[37] ), .C(n_59703), .Z(n_3674
		));
	notech_ao4 i_3726154(.A(n_59595), .B(n_40879), .C(n_58225), .D(n_39916),
		 .Z(n_3675));
	notech_ao3 i_10874046(.A(n_60037), .B(\to_acu2_0[36] ), .C(n_59703), .Z(n_3676
		));
	notech_ao4 i_3626153(.A(n_59595), .B(n_40876), .C(n_58223), .D(n_39915),
		 .Z(n_3677));
	notech_ao3 i_10774047(.A(n_60037), .B(\to_acu2_0[35] ), .C(n_59695), .Z(n_3678
		));
	notech_ao4 i_3526152(.A(n_59595), .B(n_40877), .C(n_58223), .D(n_39913),
		 .Z(n_3679));
	notech_ao3 i_10674048(.A(n_60037), .B(\to_acu2_0[34] ), .C(n_59690), .Z(n_3680
		));
	notech_ao4 i_3426151(.A(n_59595), .B(n_40848), .C(n_58223), .D(n_39912),
		 .Z(n_3681));
	notech_ao3 i_16373991(.A(n_60037), .B(\to_acu2_0[33] ), .C(n_59690), .Z(n_3682
		));
	notech_ao4 i_3326150(.A(n_59595), .B(n_40849), .C(n_58223), .D(n_39910),
		 .Z(n_3683));
	notech_ao3 i_16473990(.A(n_60037), .B(\to_acu2_0[32] ), .C(n_59690), .Z(n_3684
		));
	notech_ao4 i_3226149(.A(n_59595), .B(n_40850), .C(n_58223), .D(n_39909),
		 .Z(n_3685));
	notech_ao3 i_16573989(.A(n_60037), .B(\to_acu2_0[31] ), .C(n_59690), .Z(n_3686
		));
	notech_ao4 i_3126148(.A(n_59595), .B(n_40851), .C(n_58220), .D(n_39907),
		 .Z(n_3687));
	notech_ao3 i_16673988(.A(n_60037), .B(\to_acu2_0[30] ), .C(n_59690), .Z(n_3688
		));
	notech_ao4 i_3026147(.A(n_59595), .B(n_40852), .C(n_58218), .D(n_39906),
		 .Z(n_3689));
	notech_ao3 i_16773987(.A(n_60037), .B(\to_acu2_0[29] ), .C(n_59690), .Z(n_3690
		));
	notech_ao4 i_2926146(.A(n_59595), .B(n_40911), .C(n_58218), .D(n_39904),
		 .Z(n_3691));
	notech_ao3 i_8374071(.A(n_60036), .B(\to_acu2_0[28] ), .C(n_59690), .Z(n_3692
		));
	notech_ao4 i_2826145(.A(n_59595), .B(n_40907), .C(n_58218), .D(n_39903),
		 .Z(n_3693));
	notech_ao3 i_8274072(.A(n_60036), .B(\to_acu2_0[27] ), .C(n_59694), .Z(n_3694
		));
	notech_ao4 i_2726144(.A(n_59592), .B(n_40908), .C(n_58218), .D(n_39901),
		 .Z(n_3695));
	notech_ao3 i_4274112(.A(n_60036), .B(\to_acu2_0[26] ), .C(n_59690), .Z(n_3696
		));
	notech_ao4 i_2626143(.A(n_59590), .B(n_40910), .C(n_58218), .D(n_39900),
		 .Z(n_3697));
	notech_ao3 i_8174073(.A(n_60036), .B(\to_acu2_0[25] ), .C(n_59690), .Z(n_3698
		));
	notech_ao4 i_2526142(.A(n_59590), .B(n_40909), .C(n_58218), .D(n_39898),
		 .Z(n_3699));
	notech_ao3 i_8074074(.A(n_60036), .B(\to_acu2_0[24] ), .C(n_59690), .Z(n_3700
		));
	notech_ao4 i_2426141(.A(n_59590), .B(n_40904), .C(n_58218), .D(n_39897),
		 .Z(n_3701));
	notech_ao3 i_10374051(.A(n_60036), .B(\to_acu2_0[23] ), .C(n_59686), .Z(n_3702
		));
	notech_ao4 i_2326140(.A(n_59590), .B(n_40905), .C(n_58218), .D(n_39895),
		 .Z(n_3703));
	notech_ao3 i_10274052(.A(n_60037), .B(\to_acu2_0[22] ), .C(n_59686), .Z(n_3704
		));
	notech_ao4 i_2226139(.A(n_59590), .B(n_40903), .C(n_58218), .D(n_39894),
		 .Z(n_3705));
	notech_ao3 i_10174053(.A(n_60037), .B(\to_acu2_0[21] ), .C(n_59686), .Z(n_3706
		));
	notech_ao4 i_2126138(.A(n_59590), .B(n_40902), .C(n_58218), .D(n_39892),
		 .Z(n_3707));
	notech_ao3 i_7974075(.A(n_60037), .B(\to_acu2_0[20] ), .C(n_59686), .Z(n_3708
		));
	notech_ao4 i_2026137(.A(n_59590), .B(n_40901), .C(n_58220), .D(n_39891),
		 .Z(n_3709));
	notech_ao3 i_7874076(.A(n_60036), .B(\to_acu2_0[19] ), .C(n_59686), .Z(n_3710
		));
	notech_ao4 i_1926136(.A(n_59590), .B(n_40899), .C(n_58220), .D(n_39889),
		 .Z(n_3711));
	notech_ao3 i_10074054(.A(n_60037), .B(\to_acu2_0[18] ), .C(n_59686), .Z(n_3712
		));
	notech_ao4 i_1826135(.A(n_59590), .B(n_40898), .C(n_58220), .D(n_39888),
		 .Z(n_3713));
	notech_ao3 i_9974055(.A(n_60037), .B(\to_acu2_0[17] ), .C(n_59690), .Z(n_3714
		));
	notech_ao4 i_1726134(.A(n_59590), .B(n_40912), .C(n_58220), .D(n_39886),
		 .Z(n_3715));
	notech_ao3 i_6574089(.A(n_60026), .B(\to_acu2_0[16] ), .C(n_59690), .Z(n_3716
		));
	notech_ao4 i_1626133(.A(n_59592), .B(n_40895), .C(n_58220), .D(n_39885),
		 .Z(n_3717));
	notech_ao3 i_9874056(.A(n_60020), .B(\to_acu2_0[15] ), .C(n_59690), .Z(n_3718
		));
	notech_ao4 i_1526132(.A(n_59592), .B(n_40896), .C(n_58220), .D(n_39883),
		 .Z(n_3719));
	notech_ao3 i_9774057(.A(n_60020), .B(\to_acu2_0[14] ), .C(n_59686), .Z(n_3720
		));
	notech_ao4 i_1426131(.A(n_59592), .B(n_40897), .C(n_58218), .D(n_39882),
		 .Z(n_3721));
	notech_ao3 i_3774117(.A(n_60020), .B(\to_acu2_0[13] ), .C(n_59690), .Z(n_3722
		));
	notech_ao4 i_1326130(.A(n_59592), .B(n_40900), .C(n_58220), .D(n_39880),
		 .Z(n_3723));
	notech_ao3 i_7774077(.A(n_60020), .B(\to_acu2_0[12] ), .C(n_59694), .Z(n_3724
		));
	notech_ao4 i_1226129(.A(n_59592), .B(n_40915), .C(n_58220), .D(n_39879),
		 .Z(n_3725));
	notech_ao3 i_9674058(.A(n_60020), .B(\to_acu2_0[11] ), .C(n_59695), .Z(n_3726
		));
	notech_ao4 i_1126128(.A(n_59590), .B(n_40922), .C(n_58220), .D(n_39877),
		 .Z(n_3727));
	notech_ao4 i_1026127(.A(n_59590), .B(n_40916), .C(n_58231), .D(n_39876),
		 .Z(n_3728));
	notech_ao4 i_4627845(.A(n_2116), .B(n_59590), .C(n_58231), .D(n_39242), 
		.Z(n_3729));
	notech_ao4 i_4227841(.A(n_2119), .B(n_59592), .C(n_58231), .D(n_39234), 
		.Z(n_3730));
	notech_ao4 i_2627825(.A(n_2122), .B(n_59592), .C(n_58231), .D(n_39202), 
		.Z(n_3731));
	notech_ao4 i_2027819(.A(n_59597), .B(n_242894385), .C(n_58231), .D(n_39192
		), .Z(n_3732));
	notech_ao4 i_1727816(.A(n_2125), .B(n_59603), .C(n_58229), .D(n_39189), 
		.Z(n_3733));
	notech_ao4 i_1527814(.A(n_2126), .B(n_59601), .C(n_58229), .D(n_39187), 
		.Z(n_3734));
	notech_ao4 i_20826536(.A(n_59603), .B(n_40835), .C(n_58229), .D(n_40464)
		, .Z(n_3735));
	notech_ao4 i_20626534(.A(n_59603), .B(n_40833), .C(n_58229), .D(n_40462)
		, .Z(n_3736));
	notech_ao4 i_20126529(.A(n_59603), .B(n_40828), .C(n_58229), .D(n_40457)
		, .Z(n_3737));
	notech_ao4 i_19926527(.A(n_59601), .B(n_40826), .C(n_58231), .D(n_40455)
		, .Z(n_3738));
	notech_ao4 i_19826526(.A(n_59601), .B(n_40825), .C(n_58231), .D(n_40454)
		, .Z(n_3739));
	notech_ao4 i_19726525(.A(n_59601), .B(n_40824), .C(n_58231), .D(n_40453)
		, .Z(n_3740));
	notech_ao4 i_19526523(.A(n_59601), .B(n_40822), .C(n_58234), .D(n_40450)
		, .Z(n_3741));
	notech_ao4 i_19426522(.A(n_59601), .B(n_40821), .C(n_58231), .D(n_40449)
		, .Z(n_3742));
	notech_ao4 i_19326521(.A(n_59603), .B(n_40820), .C(n_58231), .D(n_40448)
		, .Z(n_3743));
	notech_ao4 i_19226520(.A(n_59603), .B(n_40819), .C(n_58231), .D(n_40447)
		, .Z(n_3744));
	notech_ao4 i_19126519(.A(n_59603), .B(n_40818), .C(n_58231), .D(n_40446)
		, .Z(n_3745));
	notech_ao4 i_19026518(.A(n_59603), .B(n_40817), .C(n_58231), .D(n_40445)
		, .Z(n_3746));
	notech_ao4 i_18926517(.A(n_59603), .B(n_40816), .C(n_58231), .D(n_40444)
		, .Z(n_3747));
	notech_ao4 i_18826516(.A(n_59603), .B(n_40815), .C(n_58229), .D(n_40443)
		, .Z(n_3748));
	notech_ao4 i_18726515(.A(n_59603), .B(n_40814), .C(n_58225), .D(n_40442)
		, .Z(n_3749));
	notech_ao4 i_18626514(.A(n_59603), .B(n_40813), .C(n_58225), .D(n_40441)
		, .Z(n_3750));
	notech_ao4 i_18526513(.A(n_59603), .B(n_40812), .C(n_58225), .D(n_40440)
		, .Z(n_3751));
	notech_ao4 i_18426512(.A(n_59603), .B(n_40811), .C(n_58225), .D(n_40439)
		, .Z(n_3752));
	notech_ao4 i_18326511(.A(n_59601), .B(n_40810), .C(n_58225), .D(n_40438)
		, .Z(n_3753));
	notech_ao4 i_18226510(.A(n_59597), .B(n_40809), .C(n_58225), .D(n_40437)
		, .Z(n_3754));
	notech_ao4 i_18126509(.A(n_59597), .B(n_40808), .C(n_58225), .D(n_40436)
		, .Z(n_3755));
	notech_ao4 i_18026508(.A(n_59597), .B(n_40807), .C(n_58225), .D(n_40435)
		, .Z(n_3756));
	notech_ao4 i_17926507(.A(n_59597), .B(n_40806), .C(n_58225), .D(n_40434)
		, .Z(n_3757));
	notech_ao4 i_17826506(.A(n_59597), .B(n_40805), .C(n_58225), .D(n_40433)
		, .Z(n_3758));
	notech_ao4 i_17626504(.A(n_59597), .B(n_40803), .C(n_58229), .D(n_40431)
		, .Z(n_3759));
	notech_ao4 i_17526503(.A(n_59597), .B(n_40802), .C(n_58229), .D(n_40430)
		, .Z(n_3760));
	notech_ao4 i_17426502(.A(n_59597), .B(n_40801), .C(n_58229), .D(n_40429)
		, .Z(n_3761));
	notech_ao4 i_17226500(.A(n_59597), .B(n_40799), .C(n_58229), .D(n_40427)
		, .Z(n_3762));
	notech_ao4 i_17126499(.A(n_59597), .B(n_40798), .C(n_58229), .D(n_40426)
		, .Z(n_3763));
	notech_ao4 i_17026498(.A(n_59601), .B(n_40797), .C(n_58225), .D(n_40425)
		, .Z(n_3764));
	notech_ao4 i_16826496(.A(n_59601), .B(n_40795), .C(n_58225), .D(n_40423)
		, .Z(n_3765));
	notech_ao4 i_16726495(.A(n_58229), .B(n_40422), .C(n_59601), .D(n_40794)
		, .Z(n_3766));
	notech_ao4 i_16626494(.A(n_58229), .B(n_40421), .C(n_59601), .D(n_40793)
		, .Z(n_3767));
	notech_ao4 i_16526493(.A(n_58229), .B(n_40420), .C(n_59601), .D(n_40792)
		, .Z(n_3768));
	notech_ao4 i_16426492(.A(n_58139), .B(n_40418), .C(n_59597), .D(n_40791)
		, .Z(n_3769));
	notech_ao4 i_15926487(.A(n_59597), .B(n_40786), .C(n_58139), .D(n_40412)
		, .Z(n_3770));
	notech_ao4 i_15726485(.A(n_59597), .B(n_40784), .C(n_58139), .D(n_40410)
		, .Z(n_3771));
	notech_ao3 i_3174123(.A(n_60020), .B(in128[73]), .C(n_59695), .Z(n_48074
		));
	notech_ao4 i_15226480(.A(n_58139), .B(n_40403), .C(n_59601), .D(n_40779)
		, .Z(n_3772));
	notech_ao4 i_10926437(.A(n_58139), .B(n_40351), .C(n_59601), .D(n_40736)
		, .Z(n_3773));
	notech_ao4 i_10726435(.A(n_58139), .B(n_40348), .C(n_59511), .D(n_40734)
		, .Z(n_3774));
	notech_ao4 i_10626434(.A(n_58139), .B(n_40346), .C(n_59511), .D(n_40733)
		, .Z(n_3775));
	notech_ao4 i_10526433(.A(n_58139), .B(n_40344), .C(n_59511), .D(n_40732)
		, .Z(n_3776));
	notech_ao4 i_10426432(.A(n_58139), .B(n_40342), .C(n_59511), .D(n_40731)
		, .Z(n_3777));
	notech_ao4 i_10326431(.A(n_58139), .B(n_40340), .C(n_59511), .D(n_40730)
		, .Z(n_3778));
	notech_ao4 i_10226430(.A(n_58141), .B(n_40338), .C(n_59507), .D(n_40729)
		, .Z(n_3779));
	notech_ao4 i_10126429(.A(n_58141), .B(n_40336), .C(n_59507), .D(n_40728)
		, .Z(n_3780));
	notech_ao4 i_10026428(.A(n_58141), .B(n_40334), .C(n_59507), .D(n_40727)
		, .Z(n_3781));
	notech_ao4 i_9926427(.A(n_58141), .B(n_40332), .C(n_59507), .D(n_40892),
		 .Z(n_3782));
	notech_ao4 i_9826426(.A(n_58141), .B(n_40330), .C(n_59507), .D(n_40893),
		 .Z(n_3783));
	notech_ao4 i_9726425(.A(n_58139), .B(n_40328), .C(n_59511), .D(n_40936),
		 .Z(n_3784));
	notech_ao4 i_9626424(.A(n_58139), .B(n_40325), .C(n_59511), .D(n_40935),
		 .Z(n_3785));
	notech_ao4 i_9526423(.A(n_58141), .B(n_40323), .C(n_59511), .D(n_40934),
		 .Z(n_3786));
	notech_ao4 i_9326421(.A(n_58141), .B(n_40318), .C(n_59513), .D(n_40928),
		 .Z(n_3787));
	notech_ao4 i_9126419(.A(n_58141), .B(n_40314), .C(n_59511), .D(n_40947),
		 .Z(n_3788));
	notech_ao4 i_6326391(.A(n_59511), .B(n_40913), .C(n_58139), .D(n_40273),
		 .Z(n_3789));
	notech_ao4 i_5526383(.A(n_59511), .B(n_40871), .C(n_58135), .D(n_40264),
		 .Z(n_3790));
	notech_ao4 i_5426382(.A(n_59511), .B(n_40869), .C(n_58135), .D(n_40263),
		 .Z(n_3791));
	notech_ao4 i_5226380(.A(n_59511), .B(n_40868), .C(n_58135), .D(n_40261),
		 .Z(n_3792));
	notech_ao4 i_5126379(.A(n_59511), .B(n_40861), .C(n_58135), .D(n_40260),
		 .Z(n_3793));
	notech_ao4 i_4826376(.A(n_59507), .B(n_40888), .C(n_58135), .D(n_40257),
		 .Z(n_3794));
	notech_ao4 i_4726375(.A(n_59505), .B(n_40886), .C(n_58133), .D(n_40256),
		 .Z(n_3795));
	notech_ao4 i_4626374(.A(n_59505), .B(n_40887), .C(n_58133), .D(n_40255),
		 .Z(n_3796));
	notech_ao4 i_4326371(.A(n_59505), .B(n_40884), .C(n_58133), .D(n_40252),
		 .Z(n_3797));
	notech_ao4 i_4226370(.A(n_59505), .B(n_40882), .C(n_58133), .D(n_40251),
		 .Z(n_3798));
	notech_ao4 i_4126369(.A(n_59505), .B(n_40880), .C(n_58133), .D(n_40250),
		 .Z(n_3799));
	notech_ao4 i_3926367(.A(n_59505), .B(n_40881), .C(n_58135), .D(n_40249),
		 .Z(n_3800));
	notech_ao4 i_3826366(.A(n_59505), .B(n_40878), .C(n_58135), .D(n_40248),
		 .Z(n_3801));
	notech_ao4 i_3726365(.A(n_59505), .B(n_40879), .C(n_58135), .D(n_40247),
		 .Z(n_3802));
	notech_ao4 i_3626364(.A(n_59505), .B(n_40876), .C(n_58139), .D(n_40245),
		 .Z(n_3803));
	notech_ao4 i_3526363(.A(n_59505), .B(n_40877), .C(n_58135), .D(n_40243),
		 .Z(n_3804));
	notech_ao4 i_3426362(.A(n_59507), .B(n_40848), .C(n_58135), .D(n_40241),
		 .Z(n_3805));
	notech_ao4 i_3326361(.A(n_59507), .B(n_40849), .C(n_58135), .D(n_40239),
		 .Z(n_3806));
	notech_ao4 i_3226360(.A(n_59507), .B(n_40850), .C(n_58135), .D(n_40237),
		 .Z(n_3807));
	notech_ao4 i_3126359(.A(n_59507), .B(n_40851), .C(n_58135), .D(n_40235),
		 .Z(n_3808));
	notech_ao4 i_3026358(.A(n_59507), .B(n_40852), .C(n_58135), .D(n_40233),
		 .Z(n_3809));
	notech_ao4 i_2926357(.A(n_59505), .B(n_40911), .C(n_58146), .D(n_40231),
		 .Z(n_3810));
	notech_ao4 i_2826356(.A(n_59505), .B(n_40907), .C(n_58146), .D(n_40229),
		 .Z(n_3811));
	notech_ao4 i_2726355(.A(n_59507), .B(n_40908), .C(n_58146), .D(n_40227),
		 .Z(n_3812));
	notech_ao4 i_2626354(.A(n_59507), .B(n_40910), .C(n_58146), .D(n_40225),
		 .Z(n_3813));
	notech_ao4 i_2526353(.A(n_59507), .B(n_40909), .C(n_58146), .D(n_40223),
		 .Z(n_3814));
	notech_ao4 i_2426352(.A(n_59513), .B(n_40904), .C(n_58146), .D(n_40221),
		 .Z(n_3815));
	notech_ao4 i_2126349(.A(n_59518), .B(n_40902), .C(n_58146), .D(n_40215),
		 .Z(n_3816));
	notech_ao4 i_2026348(.A(n_59518), .B(n_40901), .C(n_58146), .D(n_40213),
		 .Z(n_3817));
	notech_ao4 i_1826346(.A(n_59518), .B(n_40898), .C(n_58146), .D(n_40209),
		 .Z(n_3818));
	notech_ao4 i_1726345(.A(n_59518), .B(n_40912), .C(n_58146), .D(n_40207),
		 .Z(n_3819));
	notech_ao3 i_3312(.A(n_60025), .B(udeco[18]), .C(n_59695), .Z(n_43300)
		);
	notech_ao3 i_3316(.A(n_60025), .B(udeco[22]), .C(n_59694), .Z(n_43324)
		);
	notech_ao3 i_3317(.A(n_60025), .B(udeco[23]), .C(n_59695), .Z(n_43330)
		);
	notech_ao3 i_3318(.A(n_60025), .B(udeco[24]), .C(n_59695), .Z(n_43336)
		);
	notech_ao3 i_3319(.A(n_60025), .B(udeco[25]), .C(n_59695), .Z(n_43342)
		);
	notech_ao3 i_3326(.A(n_60025), .B(udeco[32]), .C(n_59695), .Z(n_43384)
		);
	notech_ao3 i_3331(.A(n_60020), .B(udeco[37]), .C(n_59695), .Z(n_43414)
		);
	notech_ao4 i_4227713(.A(n_2119), .B(n_59518), .C(n_58150), .D(n_39309), 
		.Z(n_3280));
	notech_ao4 i_65991(.A(n_224196468), .B(n_2917), .C(n_2915), .D(n_40501),
		 .Z(n_2027));
	notech_ao3 i_228(.A(n_60015), .B(\to_acu2_0[6] ), .C(n_59695), .Z(n_2022
		));
	notech_ao3 i_248(.A(n_60015), .B(in128[89]), .C(n_59695), .Z(n_2021));
	notech_ao3 i_252(.A(n_60015), .B(in128[93]), .C(n_59694), .Z(n_2020));
	notech_nor2 i_333(.A(n_2948), .B(n_40488), .Z(n_2019));
	notech_ao3 i_355(.A(n_60015), .B(\to_acu2_0[10] ), .C(n_59694), .Z(n_2018
		));
	notech_ao3 i_356(.A(n_60015), .B(\to_acu2_0[8] ), .C(n_59694), .Z(n_2017
		));
	notech_ao3 i_378(.A(n_60015), .B(in128[27]), .C(n_59694), .Z(n_2016));
	notech_ao3 i_379(.A(n_60020), .B(in128[49]), .C(n_59694), .Z(n_2015));
	notech_ao3 i_380(.A(n_60020), .B(in128[28]), .C(n_59694), .Z(n_2014));
	notech_ao3 i_383(.A(n_60020), .B(in128[53]), .C(n_59694), .Z(n_2013));
	notech_ao3 i_384(.A(n_60015), .B(in128[40]), .C(n_59694), .Z(n_2012));
	notech_ao3 i_385(.A(n_60020), .B(\to_acu2_0[3] ), .C(n_59694), .Z(n_2011
		));
	notech_ao4 i_4627717(.A(n_2116), .B(n_59516), .C(n_58150), .D(n_39315), 
		.Z(n_3279));
	notech_ao3 i_386(.A(n_60020), .B(in128[48]), .C(n_59694), .Z(n_2010));
	notech_ao3 i_387(.A(n_60025), .B(in128[54]), .C(n_59694), .Z(n_2009));
	notech_ao3 i_391(.A(n_60026), .B(in128[34]), .C(n_59666), .Z(n_2008));
	notech_ao3 i_392(.A(n_60026), .B(in128[33]), .C(n_59632), .Z(n_2007));
	notech_ao3 i_393(.A(n_60026), .B(in128[32]), .C(n_59632), .Z(n_2006));
	notech_ao3 i_395(.A(n_60026), .B(\to_acu2_0[4] ), .C(n_59632), .Z(n_2005
		));
	notech_nor2 i_33574156(.A(n_2116), .B(n_59516), .Z(n_3278));
	notech_ao3 i_396(.A(n_60026), .B(in128[74]), .C(n_59632), .Z(n_2004));
	notech_ao3 i_397(.A(n_60026), .B(in128[37]), .C(n_59632), .Z(n_2003));
	notech_ao3 i_398(.A(n_60026), .B(in128[43]), .C(n_59632), .Z(n_2002));
	notech_ao3 i_399(.A(n_60026), .B(in128[36]), .C(n_59632), .Z(n_2001));
	notech_ao3 i_400(.A(n_60026), .B(in128[38]), .C(n_59632), .Z(n_2000));
	notech_ao3 i_401(.A(n_60026), .B(in128[50]), .C(n_59632), .Z(n_1999));
	notech_ao3 i_402(.A(n_60026), .B(in128[76]), .C(n_59632), .Z(n_1998));
	notech_ao3 i_403(.A(n_60026), .B(in128[42]), .C(n_59632), .Z(n_1997));
	notech_ao3 i_404(.A(n_60026), .B(in128[51]), .C(n_59634), .Z(n_1996));
	notech_ao3 i_406(.A(n_60025), .B(in128[35]), .C(n_59634), .Z(n_1995));
	notech_ao3 i_407(.A(n_60025), .B(in128[63]), .C(n_59634), .Z(n_1994));
	notech_ao3 i_408(.A(n_60025), .B(in128[62]), .C(n_59634), .Z(n_1993));
	notech_ao3 i_409(.A(n_60025), .B(in128[60]), .C(n_59634), .Z(n_1992));
	notech_ao3 i_410(.A(n_60025), .B(in128[59]), .C(n_59634), .Z(n_1991));
	notech_ao3 i_411(.A(n_60025), .B(in128[57]), .C(n_59632), .Z(n_1990));
	notech_ao3 i_412(.A(n_60025), .B(in128[56]), .C(n_59632), .Z(n_1989));
	notech_ao3 i_413(.A(n_60025), .B(in128[31]), .C(n_59632), .Z(n_1988));
	notech_ao3 i_414(.A(n_60026), .B(in128[44]), .C(n_59634), .Z(n_1987));
	notech_ao3 i_415(.A(n_60025), .B(in128[39]), .C(n_59634), .Z(n_1986));
	notech_ao3 i_418(.A(n_60025), .B(in128[78]), .C(n_59632), .Z(n_1985));
	notech_ao3 i_419(.A(n_60025), .B(\to_acu2_0[0] ), .C(n_59643), .Z(n_1984
		));
	notech_nor2 i_30674159(.A(n_2125), .B(n_59516), .Z(n_3277));
	notech_ao3 i_426(.A(n_59992), .B(in128[55]), .C(n_59643), .Z(n_1983));
	notech_ao3 i_427(.A(n_59957), .B(in128[64]), .C(n_59643), .Z(n_1982));
	notech_ao3 i_428(.A(n_59957), .B(in128[47]), .C(n_59643), .Z(n_1981));
	notech_ao3 i_430(.A(n_59957), .B(\to_acu2_0[2] ), .C(n_59643), .Z(n_1980
		));
	notech_ao3 i_27174161(.A(n_59957), .B(in128[112]), .C(n_59647), .Z(n_3276
		));
	notech_ao3 i_432(.A(n_59957), .B(in128[26]), .C(n_59647), .Z(n_1979));
	notech_ao3 i_433(.A(n_59957), .B(in128[45]), .C(n_59647), .Z(n_1978));
	notech_ao3 i_436(.A(n_59957), .B(in128[69]), .C(n_59647), .Z(n_1977));
	notech_ao3 i_437(.A(n_59957), .B(\to_acu2_0[1] ), .C(n_59647), .Z(n_1976
		));
	notech_ao3 i_438(.A(n_59957), .B(\to_acu2_0[9] ), .C(n_59647), .Z(n_1975
		));
	notech_ao3 i_439(.A(n_59957), .B(in128[30]), .C(n_59643), .Z(n_1974));
	notech_ao3 i_442(.A(n_59957), .B(in128[29]), .C(n_59643), .Z(n_1973));
	notech_ao3 i_443(.A(n_59957), .B(in128[71]), .C(n_59632), .Z(n_1972));
	notech_ao3 i_444(.A(n_59957), .B(in128[46]), .C(n_59632), .Z(n_1971));
	notech_ao3 i_448(.A(n_59952), .B(in128[72]), .C(n_59632), .Z(n_1970));
	notech_ao3 i_451(.A(n_59952), .B(in128[52]), .C(n_59643), .Z(n_1969));
	notech_ao3 i_452(.A(n_59952), .B(in128[41]), .C(n_59643), .Z(n_1968));
	notech_ao3 i_453(.A(n_59952), .B(in128[70]), .C(n_59643), .Z(n_1967));
	notech_ao3 i_454(.A(n_59952), .B(in128[61]), .C(n_59643), .Z(n_1966));
	notech_ao3 i_456(.A(n_59952), .B(in128[58]), .C(n_59643), .Z(n_1965));
	notech_ao3 i_460(.A(n_59957), .B(in128[77]), .C(n_59643), .Z(n_1964));
	notech_ao3 i_461(.A(n_59957), .B(in128[85]), .C(n_59634), .Z(n_1963));
	notech_ao3 i_466(.A(n_59957), .B(in128[24]), .C(n_59625), .Z(n_1962));
	notech_ao3 i_467(.A(n_59952), .B(in128[67]), .C(n_59625), .Z(n_1961));
	notech_ao3 i_468(.A(n_59952), .B(\to_acu2_0[5] ), .C(n_59625), .Z(n_1960
		));
	notech_ao3 i_469(.A(n_59957), .B(in128[66]), .C(n_59625), .Z(n_1959));
	notech_ao3 i_473(.A(n_59957), .B(\to_acu2_0[58] ), .C(n_59625), .Z(n_1958
		));
	notech_ao3 i_476(.A(n_59968), .B(\to_acu2_0[7] ), .C(n_59625), .Z(n_1957
		));
	notech_ao3 i_25674162(.A(n_59968), .B(in128[97]), .C(n_59623), .Z(n_3275
		));
	notech_ao3 i_477(.A(n_59968), .B(in128[79]), .C(n_59623), .Z(n_1956));
	notech_ao3 i_485(.A(n_59968), .B(in128[65]), .C(n_59623), .Z(n_1955));
	notech_nor2 i_3729806(.A(int_excl[2]), .B(n_5423), .Z(n_1954));
	notech_nor2 i_66875(.A(idx_deco[1]), .B(n_39370), .Z(n_5414));
	notech_ao4 i_1(.A(n_2870), .B(n_39133), .C(n_2871), .D(n_2865), .Z(n_1953
		));
	notech_nand2 i_6351(.A(idx_deco[1]), .B(n_39370), .Z(n_5408));
	notech_ao3 i_286(.A(n_59968), .B(in128[127]), .C(n_59625), .Z(n_48398)
		);
	notech_ao3 i_69(.A(n_59968), .B(udeco[68]), .C(n_59623), .Z(n_43600));
	notech_ao3 i_70(.A(n_59968), .B(udeco[69]), .C(n_59625), .Z(n_43606));
	notech_ao3 i_71(.A(n_59968), .B(udeco[70]), .C(n_59625), .Z(n_43612));
	notech_ao3 i_72(.A(n_59968), .B(udeco[71]), .C(n_59625), .Z(n_43618));
	notech_ao3 i_73(.A(n_59968), .B(udeco[72]), .C(n_59625), .Z(n_43624));
	notech_ao3 i_74(.A(n_59968), .B(udeco[73]), .C(n_59625), .Z(n_43630));
	notech_ao3 i_75(.A(n_59968), .B(udeco[74]), .C(n_59625), .Z(n_43636));
	notech_ao3 i_76(.A(n_59963), .B(udeco[75]), .C(n_59625), .Z(n_43642));
	notech_ao3 i_77(.A(n_59963), .B(udeco[76]), .C(n_59625), .Z(n_43648));
	notech_ao3 i_78(.A(n_59963), .B(udeco[77]), .C(n_59625), .Z(n_43654));
	notech_ao3 i_79(.A(n_59963), .B(udeco[78]), .C(n_59625), .Z(n_43660));
	notech_ao3 i_80(.A(n_59957), .B(udeco[79]), .C(n_59625), .Z(n_43666));
	notech_ao3 i_81(.A(n_59957), .B(udeco[80]), .C(n_59623), .Z(n_43672));
	notech_ao3 i_82(.A(n_59963), .B(udeco[81]), .C(n_59634), .Z(n_43678));
	notech_ao3 i_83(.A(n_59963), .B(udeco[82]), .C(n_59634), .Z(n_43684));
	notech_ao3 i_84(.A(n_59963), .B(udeco[83]), .C(n_59634), .Z(n_43690));
	notech_ao3 i_86(.A(n_59963), .B(udeco[85]), .C(n_59623), .Z(n_43702));
	notech_ao3 i_88(.A(n_59963), .B(udeco[87]), .C(n_59623), .Z(n_43714));
	notech_ao3 i_90(.A(n_59963), .B(udeco[89]), .C(n_59634), .Z(n_43726));
	notech_ao3 i_91(.A(n_59963), .B(udeco[90]), .C(n_59634), .Z(n_43732));
	notech_ao3 i_92(.A(n_59952), .B(udeco[91]), .C(n_59634), .Z(n_43738));
	notech_ao3 i_93(.A(n_59941), .B(udeco[92]), .C(n_59634), .Z(n_43744));
	notech_ao3 i_94(.A(n_59941), .B(udeco[93]), .C(n_59634), .Z(n_43750));
	notech_ao3 i_95(.A(n_59941), .B(udeco[94]), .C(n_59634), .Z(n_43756));
	notech_ao3 i_96(.A(n_59941), .B(udeco[95]), .C(n_59623), .Z(n_43762));
	notech_ao3 i_97(.A(n_59941), .B(udeco[96]), .C(n_59623), .Z(n_43768));
	notech_ao3 i_98(.A(n_59941), .B(udeco[97]), .C(n_59623), .Z(n_43774));
	notech_ao3 i_99(.A(n_59946), .B(udeco[98]), .C(n_59623), .Z(n_43780));
	notech_ao3 i_100(.A(n_59946), .B(udeco[99]), .C(n_59623), .Z(n_43786));
	notech_ao3 i_101(.A(n_59946), .B(udeco[100]), .C(n_59623), .Z(n_43792)
		);
	notech_ao3 i_102(.A(n_59941), .B(udeco[101]), .C(n_59623), .Z(n_43798)
		);
	notech_ao3 i_103(.A(n_59946), .B(udeco[102]), .C(n_59623), .Z(n_43804)
		);
	notech_ao3 i_105(.A(n_59946), .B(udeco[104]), .C(n_59623), .Z(n_43816)
		);
	notech_ao3 i_106(.A(n_59941), .B(udeco[105]), .C(n_59623), .Z(n_43822)
		);
	notech_ao3 i_107(.A(n_59941), .B(udeco[106]), .C(n_59623), .Z(n_43828)
		);
	notech_ao3 i_109(.A(n_59941), .B(udeco[108]), .C(n_59658), .Z(n_43840)
		);
	notech_ao3 i_110(.A(n_59941), .B(udeco[109]), .C(n_59658), .Z(n_43846)
		);
	notech_ao3 i_112(.A(n_59941), .B(udeco[111]), .C(n_59658), .Z(n_43858)
		);
	notech_ao3 i_113(.A(n_59941), .B(udeco[112]), .C(n_59658), .Z(n_43864)
		);
	notech_ao3 i_114(.A(n_59941), .B(udeco[113]), .C(n_59658), .Z(n_43870)
		);
	notech_ao3 i_115(.A(n_59941), .B(udeco[114]), .C(n_59658), .Z(n_43876)
		);
	notech_ao3 i_116(.A(n_59941), .B(udeco[115]), .C(n_59662), .Z(n_43882)
		);
	notech_ao3 i_117(.A(n_59941), .B(udeco[116]), .C(n_59662), .Z(n_43888)
		);
	notech_ao3 i_118(.A(n_59941), .B(udeco[117]), .C(n_59662), .Z(n_43894)
		);
	notech_ao3 i_119(.A(n_59941), .B(udeco[118]), .C(n_59658), .Z(n_43900)
		);
	notech_ao3 i_120(.A(n_59941), .B(udeco[119]), .C(n_59662), .Z(n_43906)
		);
	notech_ao3 i_121(.A(n_59946), .B(udeco[120]), .C(n_59657), .Z(n_43912)
		);
	notech_ao3 i_122(.A(n_59952), .B(udeco[121]), .C(n_59658), .Z(n_43918)
		);
	notech_ao3 i_123(.A(n_59952), .B(udeco[122]), .C(n_59657), .Z(n_43924)
		);
	notech_ao3 i_124(.A(n_59952), .B(udeco[123]), .C(n_59657), .Z(n_43930)
		);
	notech_ao3 i_125(.A(n_59946), .B(udeco[124]), .C(n_59657), .Z(n_43936)
		);
	notech_ao3 i_126(.A(n_59952), .B(udeco[125]), .C(n_59658), .Z(n_43942)
		);
	notech_ao3 i_127(.A(n_59952), .B(udeco[126]), .C(n_59658), .Z(n_43948)
		);
	notech_ao3 i_416(.A(in128[1]), .B(in128[2]), .C(n_59516), .Z(n_49787));
	notech_ao3 i_200(.A(n_59952), .B(in128[1]), .C(n_59658), .Z(n_47642));
	notech_ao3 i_227(.A(n_59952), .B(repz), .C(n_59658), .Z(n_49793));
	notech_ao3 i_207(.A(n_59952), .B(udeco[103]), .C(n_59658), .Z(n_43810)
		);
	notech_ao3 i_127194(.A(n_59952), .B(\nbus_12182[0] ), .C(n_59658), .Z(n_44841
		));
	notech_ao3 i_227195(.A(n_59952), .B(\nbus_12182[1] ), .C(n_59662), .Z(n_44847
		));
	notech_ao3 i_327196(.A(n_59952), .B(\nbus_12182[2] ), .C(n_59666), .Z(n_44853
		));
	notech_ao3 i_427197(.A(n_59946), .B(\nbus_12182[3] ), .C(n_59666), .Z(n_44859
		));
	notech_ao3 i_527198(.A(n_59946), .B(\nbus_12182[4] ), .C(n_59666), .Z(n_44865
		));
	notech_ao3 i_627199(.A(n_59946), .B(\nbus_12182[5] ), .C(n_59666), .Z(n_44871
		));
	notech_nand3 i_2515(.A(n_2226), .B(n_59946), .C(n_40937), .Z(n_1949));
	notech_or2 i_6369(.A(idx_deco[1]), .B(idx_deco[0]), .Z(n_5396));
	notech_nor2 i_290(.A(n_227894235), .B(n_59516), .Z(n_44449));
	notech_nor2 i_291(.A(n_228694243), .B(n_59518), .Z(n_44455));
	notech_nor2 i_292(.A(n_229494251), .B(n_59518), .Z(n_44461));
	notech_nor2 i_293(.A(n_230294259), .B(n_59518), .Z(n_44467));
	notech_nor2 i_294(.A(n_231094267), .B(n_59522), .Z(n_44473));
	notech_nor2 i_295(.A(n_231894275), .B(n_59518), .Z(n_44479));
	notech_nor2 i_296(.A(n_232694283), .B(n_59518), .Z(n_44485));
	notech_nor2 i_297(.A(n_233494291), .B(n_59518), .Z(n_44491));
	notech_nor2 i_298(.A(n_234294299), .B(n_59518), .Z(n_44497));
	notech_nor2 i_299(.A(n_235094307), .B(n_59518), .Z(n_44503));
	notech_nor2 i_300(.A(n_235894315), .B(n_59518), .Z(n_44509));
	notech_nor2 i_301(.A(n_236694323), .B(n_59516), .Z(n_44515));
	notech_nor2 i_302(.A(n_237494331), .B(n_59513), .Z(n_44521));
	notech_nor2 i_303(.A(n_238294339), .B(n_59513), .Z(n_44527));
	notech_nor2 i_305(.A(n_239494351), .B(n_59513), .Z(n_44539));
	notech_nor2 i_307(.A(n_240894365), .B(n_59513), .Z(n_44551));
	notech_nor2 i_308(.A(n_241894375), .B(n_59513), .Z(n_44557));
	notech_nor2 i_309(.A(n_242894385), .B(n_59513), .Z(n_44563));
	notech_nor2 i_310(.A(n_243894395), .B(n_59513), .Z(n_44569));
	notech_nor2 i_311(.A(n_244894405), .B(n_59513), .Z(n_44575));
	notech_nor2 i_312(.A(n_245894415), .B(n_59513), .Z(n_44581));
	notech_nor2 i_313(.A(n_246894425), .B(n_59513), .Z(n_44587));
	notech_nor2 i_314(.A(n_247894435), .B(n_59516), .Z(n_44593));
	notech_nor2 i_316(.A(n_248894445), .B(n_59516), .Z(n_44605));
	notech_nor2 i_317(.A(n_249894455), .B(n_59516), .Z(n_44611));
	notech_nor2 i_318(.A(n_250894465), .B(n_59516), .Z(n_44617));
	notech_nor2 i_319(.A(n_251894475), .B(n_59516), .Z(n_44623));
	notech_nor2 i_320(.A(n_252894485), .B(n_59513), .Z(n_44629));
	notech_nor2 i_321(.A(n_254094497), .B(n_59513), .Z(n_44635));
	notech_nor2 i_322(.A(n_3123), .B(n_40326), .Z(n_44641));
	notech_nor2 i_323(.A(n_3123), .B(n_40319), .Z(n_44647));
	notech_nor2 i_325(.A(n_3123), .B(n_40312), .Z(n_44659));
	notech_nor2 i_326(.A(n_3123), .B(n_40309), .Z(n_44665));
	notech_nor2 i_327(.A(n_3123), .B(n_40307), .Z(n_44671));
	notech_nor2 i_328(.A(n_3123), .B(n_40304), .Z(n_44677));
	notech_nor2 i_329(.A(n_3123), .B(n_40300), .Z(n_44683));
	notech_nor2 i_330(.A(n_2948), .B(n_40298), .Z(n_44689));
	notech_nor2 i_332(.A(n_2948), .B(n_40295), .Z(n_44701));
	notech_nor2 i_336(.A(n_2948), .B(n_40293), .Z(n_44725));
	notech_nor2 i_337(.A(n_2948), .B(n_40290), .Z(n_44731));
	notech_or4 i_151(.A(n_2870), .B(pg_fault), .C(pc_req), .D(n_227296437), 
		.Z(n_2025));
	notech_or2 i_2461(.A(int_excl[5]), .B(n_224496465), .Z(n_1940));
	notech_nand3 i_11(.A(n_40937), .B(n_59946), .C(n_59022), .Z(n_5276));
	notech_nand2 i_210237(.A(n_1940), .B(start), .Z(n_5392));
	notech_nand2 i_65723(.A(n_2858), .B(n_2855), .Z(n_1932));
	notech_nand2 i_65730(.A(n_40863), .B(n_40862), .Z(n_1931));
	notech_and2 i_95610218(.A(\to_acu2_0[0] ), .B(\to_acu2_0[1] ), .Z(n_1925
		));
	notech_nor2 i_334(.A(n_2948), .B(n_40281), .Z(n_44713));
	notech_nor2 i_324(.A(n_3123), .B(n_40279), .Z(n_44653));
	notech_and2 i_202(.A(n_5408), .B(n_5396), .Z(n_1952));
	notech_ao3 i_225(.A(udeco[103]), .B(rep), .C(n_59516), .Z(n_49799));
	notech_ao3 i_3420(.A(n_59946), .B(udeco[127]), .C(n_59666), .Z(n_43954)
		);
	notech_nor2 i_226(.A(n_59516), .B(n_40469), .Z(n_45938));
	notech_nand2 i_393732(.A(n_2226), .B(n_59946), .Z(n_5630));
	notech_nao3 i_8(.A(n_59946), .B(n_40937), .C(n_59666), .Z(n_5768));
	notech_nor2 i_13(.A(n_2884), .B(pc_req), .Z(n_41563));
	notech_nao3 i_21175785(.A(n_59946), .B(n_40937), .C(n_1512), .Z(n_3274)
		);
	notech_and2 i_31(.A(n_2184), .B(n_40864), .Z(n_1773));
	notech_and3 i_134(.A(n_40943), .B(n_40941), .C(n_258294539), .Z(n_1772)
		);
	notech_or2 i_155(.A(int_excl[1]), .B(int_excl[0]), .Z(n_5423));
	notech_ao3 i_166(.A(n_258194538), .B(n_39148), .C(\fpu_indrm[2] ), .Z(n_1768
		));
	notech_nand2 i_189(.A(n_2181), .B(n_2180), .Z(n_1763));
	notech_and2 i_208(.A(n_40943), .B(n_40941), .Z(n_1757));
	notech_nand3 i_223(.A(n_59666), .B(n_2870), .C(n_59946), .Z(n_1753));
	notech_and3 i_3080(.A(n_2226), .B(lenpc2[31]), .C(n_59946), .Z(n_44289)
		);
	notech_nor2 i_3514(.A(n_2171), .B(n_40468), .Z(n_42972));
	notech_or4 i_6337(.A(fsm[2]), .B(n_2864), .C(fsm[0]), .D(n_39374), .Z(n_5770
		));
	notech_and2 i_775787(.A(n_2025), .B(n_40937), .Z(n_3273));
	notech_ao4 i_123151(.A(n_40918), .B(n_39987), .C(n_58150), .D(n_39415), 
		.Z(n_3272));
	notech_ao4 i_223152(.A(n_59516), .B(n_39380), .C(n_58150), .D(n_39418), 
		.Z(n_3271));
	notech_nand2 i_1125661(.A(n_60065), .B(n_1642), .Z(n_3270));
	notech_nand2 i_1425664(.A(n_60065), .B(n_1641), .Z(n_3269));
	notech_nand3 i_3125681(.A(n_60065), .B(n_1448), .C(n_1640), .Z(n_3268)
		);
	notech_nand2 i_5225702(.A(n_60065), .B(n_1639), .Z(n_3267));
	notech_nand3 i_5925709(.A(n_60065), .B(n_3273), .C(n_1638), .Z(n_3266)
		);
	notech_nand2 i_6025710(.A(n_60065), .B(n_1637), .Z(n_3265));
	notech_nand2 i_6125711(.A(n_60065), .B(n_1636), .Z(n_3264));
	notech_nand2 i_6625716(.A(n_60065), .B(n_1635), .Z(n_3263));
	notech_nand2 i_7425724(.A(n_60066), .B(n_1634), .Z(n_3262));
	notech_nand3 i_8125731(.A(n_60065), .B(n_1632), .C(n_1540), .Z(n_3261)
		);
	notech_nand3 i_8225732(.A(n_16151033), .B(n_1630), .C(n_1543), .Z(n_3260
		));
	notech_nand3 i_8325733(.A(n_16151033), .B(n_1628), .C(n_1546), .Z(n_3259
		));
	notech_nand3 i_8425734(.A(n_16151033), .B(n_1626), .C(n_1549), .Z(n_3258
		));
	notech_nand3 i_8525735(.A(n_60066), .B(n_1624), .C(n_1552), .Z(n_3257)
		);
	notech_nand3 i_8625736(.A(n_60066), .B(n_1622), .C(n_1555), .Z(n_3256)
		);
	notech_nand3 i_8725737(.A(n_60065), .B(n_1620), .C(n_1558), .Z(n_3255)
		);
	notech_nand3 i_8825738(.A(n_60065), .B(n_1618), .C(n_1561), .Z(n_3254)
		);
	notech_nand2 i_8925739(.A(n_60065), .B(n_1617), .Z(n_3253));
	notech_nand2 i_9025740(.A(n_60065), .B(n_1616), .Z(n_3252));
	notech_nand2 i_9125741(.A(n_60065), .B(n_1615), .Z(n_3251));
	notech_nand2 i_9325743(.A(n_60061), .B(n_1614), .Z(n_3250));
	notech_nand2 i_9425744(.A(n_60061), .B(n_1613), .Z(n_3249));
	notech_nand2 i_9525745(.A(n_60061), .B(n_1612), .Z(n_3248));
	notech_nand2 i_9625746(.A(n_60061), .B(n_1611), .Z(n_3247));
	notech_nand2 i_9725747(.A(n_60061), .B(n_1610), .Z(n_3246));
	notech_nand2 i_9825748(.A(n_60061), .B(n_1609), .Z(n_3245));
	notech_nand2 i_9925749(.A(n_137396068), .B(n_1608), .Z(n_3244));
	notech_nand2 i_10025750(.A(n_137396068), .B(n_1607), .Z(n_3243));
	notech_ao4 i_123148(.A(n_59505), .B(n_40725), .C(n_58150), .D(n_40496), 
		.Z(n_3242));
	notech_ao4 i_223149(.A(n_59494), .B(n_40726), .C(n_58146), .D(n_40497), 
		.Z(n_3241));
	notech_ao4 i_123145(.A(n_59494), .B(n_40725), .C(n_58146), .D(n_40494), 
		.Z(n_3240));
	notech_ao3 i_38875788(.A(n_59946), .B(opz[0]), .C(n_59666), .Z(n_3239)
		);
	notech_ao4 i_223146(.A(n_59494), .B(n_40726), .C(n_58146), .D(n_40495), 
		.Z(n_3238));
	notech_or2 i_075797(.A(n_59666), .B(pc_req), .Z(n_5769));
	notech_ao3 i_43175789(.A(n_59946), .B(opz[1]), .C(n_59666), .Z(n_3237)
		);
	notech_ao4 i_122118(.A(n_59494), .B(n_40933), .C(n_58150), .D(n_39388), 
		.Z(n_3236));
	notech_ao4 i_222119(.A(n_59494), .B(n_40932), .C(n_58150), .D(n_39390), 
		.Z(n_3235));
	notech_ao4 i_322120(.A(n_59490), .B(n_40931), .C(n_58146), .D(n_39391), 
		.Z(n_3234));
	notech_ao4 i_422121(.A(n_59490), .B(n_40946), .C(n_58144), .D(n_39393), 
		.Z(n_3233));
	notech_ao4 i_522122(.A(n_59490), .B(n_40930), .C(n_58141), .D(n_39394), 
		.Z(n_3232));
	notech_ao4 i_622123(.A(n_59490), .B(n_40929), .C(n_58144), .D(n_39396), 
		.Z(n_3231));
	notech_ao4 i_127800(.A(n_59490), .B(n_227894235), .C(n_58144), .D(n_39172
		), .Z(n_3230));
	notech_ao4 i_227801(.A(n_59494), .B(n_228694243), .C(n_58144), .D(n_39174
		), .Z(n_3229));
	notech_ao4 i_327802(.A(n_59494), .B(n_229494251), .C(n_58141), .D(n_39175
		), .Z(n_3228));
	notech_ao4 i_427803(.A(n_59494), .B(n_230294259), .C(n_58141), .D(n_39176
		), .Z(n_3227));
	notech_ao4 i_527804(.A(n_59496), .B(n_231094267), .C(n_58141), .D(n_39177
		), .Z(n_3226));
	notech_ao4 i_627805(.A(n_59494), .B(n_231894275), .C(n_58141), .D(n_39178
		), .Z(n_3225));
	notech_ao4 i_727806(.A(n_59494), .B(n_232694283), .C(n_58141), .D(n_39179
		), .Z(n_3224));
	notech_ao4 i_827807(.A(n_59494), .B(n_233494291), .C(n_58144), .D(n_39180
		), .Z(n_3223));
	notech_ao4 i_927808(.A(n_234294299), .B(n_59494), .C(n_58144), .D(n_39181
		), .Z(n_3222));
	notech_ao4 i_1027809(.A(n_235094307), .B(n_59494), .C(n_58144), .D(n_39182
		), .Z(n_3221));
	notech_ao4 i_1127810(.A(n_235894315), .B(n_59494), .C(n_58144), .D(n_39183
		), .Z(n_3220));
	notech_ao4 i_1227811(.A(n_236694323), .B(n_59490), .C(n_58144), .D(n_39184
		), .Z(n_3219));
	notech_ao4 i_1327812(.A(n_237494331), .B(n_59490), .C(n_58144), .D(n_39185
		), .Z(n_3218));
	notech_ao4 i_1427813(.A(n_238294339), .B(n_59496), .C(n_58144), .D(n_39186
		), .Z(n_3217));
	notech_ao4 i_1627815(.A(n_239494351), .B(n_59490), .C(n_58144), .D(n_39188
		), .Z(n_3216));
	notech_ao4 i_1827817(.A(n_59490), .B(n_240894365), .C(n_58144), .D(n_39190
		), .Z(n_3215));
	notech_ao4 i_1927818(.A(n_59490), .B(n_241894375), .C(n_58144), .D(n_39191
		), .Z(n_3214));
	notech_ao4 i_2127820(.A(n_59496), .B(n_243894395), .C(n_58133), .D(n_39193
		), .Z(n_3213));
	notech_ao4 i_2227821(.A(n_59496), .B(n_244894405), .C(n_58122), .D(n_39194
		), .Z(n_3212));
	notech_ao4 i_2327822(.A(n_59496), .B(n_245894415), .C(n_58122), .D(n_39196
		), .Z(n_3211));
	notech_ao4 i_2427823(.A(n_59496), .B(n_246894425), .C(n_58122), .D(n_39198
		), .Z(n_3210));
	notech_ao4 i_2527824(.A(n_59496), .B(n_247894435), .C(n_58123), .D(n_39200
		), .Z(n_3209));
	notech_ao4 i_2727826(.A(n_59490), .B(n_248894445), .C(n_58122), .D(n_39204
		), .Z(n_3208));
	notech_ao4 i_2827827(.A(n_59490), .B(n_249894455), .C(n_58122), .D(n_39206
		), .Z(n_3207));
	notech_ao4 i_2927828(.A(n_59490), .B(n_250894465), .C(n_58122), .D(n_39208
		), .Z(n_3206));
	notech_ao4 i_3027829(.A(n_59490), .B(n_251894475), .C(n_58122), .D(n_39210
		), .Z(n_3205));
	notech_ao4 i_3127830(.A(n_59490), .B(n_252894485), .C(n_58122), .D(n_39212
		), .Z(n_3204));
	notech_ao4 i_3227831(.A(n_59490), .B(n_254094497), .C(n_58122), .D(n_39214
		), .Z(n_3203));
	notech_ao4 i_3327832(.A(n_3123), .B(n_40326), .C(n_58123), .D(n_39216), 
		.Z(n_3202));
	notech_ao4 i_3427833(.A(n_3123), .B(n_40319), .C(n_58123), .D(n_39218), 
		.Z(n_3201));
	notech_ao4 i_3627835(.A(n_3123), .B(n_40312), .C(n_58123), .D(n_39222), 
		.Z(n_3200));
	notech_ao4 i_3727836(.A(n_54557), .B(n_40309), .C(n_58123), .D(n_39224),
		 .Z(n_3199));
	notech_ao4 i_3827837(.A(n_54557), .B(n_40307), .C(n_58123), .D(n_39226),
		 .Z(n_3198));
	notech_ao4 i_3927838(.A(n_54557), .B(n_40304), .C(n_58123), .D(n_39228),
		 .Z(n_3197));
	notech_ao4 i_4027839(.A(n_54557), .B(n_40300), .C(n_58123), .D(n_39230),
		 .Z(n_3196));
	notech_ao4 i_4127840(.A(n_2948), .B(n_40298), .C(n_58123), .D(n_39232), 
		.Z(n_3195));
	notech_ao4 i_4327842(.A(n_2948), .B(n_40295), .C(n_58123), .D(n_39236), 
		.Z(n_3194));
	notech_ao4 i_4427843(.A(n_2948), .B(n_40488), .C(n_58123), .D(n_39238), 
		.Z(n_3193));
	notech_ao4 i_4727846(.A(n_2948), .B(n_40293), .C(n_58122), .D(n_39244), 
		.Z(n_3192));
	notech_ao4 i_4827847(.A(n_2948), .B(n_40290), .C(n_58117), .D(n_39246), 
		.Z(n_3191));
	notech_ao4 i_126118(.A(n_59490), .B(n_40942), .C(n_58117), .D(n_39862), 
		.Z(n_3190));
	notech_ao4 i_226119(.A(n_59490), .B(n_40925), .C(n_58117), .D(n_39864), 
		.Z(n_3189));
	notech_ao4 i_626123(.A(n_59490), .B(n_40875), .C(n_58117), .D(n_39870), 
		.Z(n_3188));
	notech_ao4 i_726124(.A(n_59490), .B(n_40924), .C(n_58117), .D(n_39871), 
		.Z(n_3187));
	notech_ao4 i_926126(.A(n_59496), .B(n_40923), .C(n_58117), .D(n_39874), 
		.Z(n_3186));
	notech_and2 i_429882(.A(cpl[0]), .B(cpl[1]), .Z(n_14051012));
	notech_or4 i_19875790(.A(twobyte), .B(fpu), .C(n_40559), .D(n_2176), .Z(n_17551047
		));
	notech_and2 i_22275791(.A(n_1597), .B(n_1505), .Z(n_3185));
	notech_and3 i_72603(.A(n_3185), .B(n_40937), .C(n_59968), .Z(n_3184));
	notech_and4 i_74326(.A(n_60061), .B(n_224396466), .C(n_18051052), .D(n_1506
		), .Z(n_3183));
	notech_and3 i_75543(.A(n_59088), .B(n_1600), .C(n_40559), .Z(n_3182));
	notech_and3 i_71458(.A(n_16151033), .B(n_1595), .C(n_1588), .Z(n_3181)
		);
	notech_and4 i_72241(.A(n_60061), .B(n_224396466), .C(n_18051052), .D(n_1514
		), .Z(n_3180));
	notech_and4 i_71477(.A(n_60065), .B(n_224396466), .C(n_18051052), .D(n_1515
		), .Z(n_3179));
	notech_and4 i_70763(.A(n_18051052), .B(n_1520), .C(n_1591), .D(n_2225), 
		.Z(n_3178));
	notech_and4 i_70741(.A(n_60065), .B(n_18051052), .C(n_224396466), .D(n_1516
		), .Z(n_3177));
	notech_and4 i_72065(.A(n_18051052), .B(n_1591), .C(n_1520), .D(n_2230), 
		.Z(n_3176));
	notech_nand2 i_1340(.A(n_2910), .B(n_1507), .Z(n_3173));
	notech_ao4 i_1335(.A(ipg_fault), .B(n_40468), .C(pc_req), .D(n_2908), .Z
		(n_3172));
	notech_or2 i_1311(.A(\fpu_indrm[4] ), .B(n_39065), .Z(n_3170));
	notech_ao4 i_1317(.A(n_40468), .B(n_269994656), .C(n_1772), .D(n_3153), 
		.Z(n_3168));
	notech_ao4 i_1304(.A(n_3157), .B(n_3139), .C(n_269294649), .D(n_40938), 
		.Z(n_3165));
	notech_ao4 i_194(.A(n_3153), .B(\to_acu2_0[4] ), .C(n_3161), .D(n_3135),
		 .Z(n_3162));
	notech_or4 i_1299(.A(n_268594642), .B(fpu), .C(n_40499), .D(n_40940), .Z
		(n_3161));
	notech_ao4 i_1294(.A(n_3153), .B(n_40940), .C(n_1757), .D(n_3158), .Z(n_3159
		));
	notech_nao3 i_29(.A(db67), .B(n_41563), .C(n_3157), .Z(n_3158));
	notech_or4 i_1287(.A(n_268594642), .B(fpu), .C(n_40499), .D(n_1925), .Z(n_3157
		));
	notech_ao4 i_205(.A(n_3139), .B(n_3154), .C(n_3153), .D(n_1772), .Z(n_3155
		));
	notech_nand2 i_1285(.A(n_39065), .B(fpu), .Z(n_3154));
	notech_or4 i_36(.A(n_2960), .B(n_3139), .C(fpu), .D(n_40499), .Z(n_3153)
		);
	notech_xor2 i_1241(.A(int_excl[2]), .B(n_5423), .Z(n_3150));
	notech_ao4 i_1165(.A(n_261494571), .B(in128[50]), .C(n_3122), .D(in128[
		42]), .Z(n_3149));
	notech_ao4 i_1146(.A(n_259594552), .B(in128[52]), .C(n_2941), .D(in128[
		60]), .Z(n_3148));
	notech_nand2 i_1138(.A(n_40938), .B(\to_acu2_0[4] ), .Z(n_3147));
	notech_nand2 i_1133(.A(\fpu_indrm[4] ), .B(n_1768), .Z(n_3146));
	notech_and3 i_1104(.A(\fpu_indrm[7] ), .B(\fpu_modrm[2] ), .C(\fpu_indrm[0] 
		), .Z(n_3142));
	notech_nao3 i_27(.A(db67), .B(n_59981), .C(n_2884), .Z(n_3139));
	notech_or4 i_3925(.A(db67), .B(n_40468), .C(\to_acu2_0[4] ), .D(\to_acu2_0[3] 
		), .Z(n_3137));
	notech_or4 i_175(.A(n_2884), .B(db67), .C(pc_req), .D(\to_acu2_0[4] ), .Z
		(n_3136));
	notech_or2 i_143(.A(db67), .B(n_40468), .Z(n_3135));
	notech_ao4 i_1094(.A(n_257594532), .B(in128[55]), .C(n_2941), .D(in128[
		63]), .Z(n_3134));
	notech_ao4 i_1090(.A(n_257294529), .B(in128[54]), .C(n_2941), .D(in128[
		62]), .Z(n_3133));
	notech_ao4 i_1086(.A(n_256994526), .B(in128[50]), .C(n_2941), .D(in128[
		58]), .Z(n_3132));
	notech_ao4 i_1082(.A(n_256694523), .B(in128[48]), .C(n_2941), .D(in128[
		56]), .Z(n_3131));
	notech_ao4 i_1078(.A(n_256394520), .B(in128[55]), .C(n_3122), .D(in128[
		47]), .Z(n_3130));
	notech_ao4 i_1074(.A(n_256094517), .B(in128[54]), .C(n_3122), .D(in128[
		46]), .Z(n_3129));
	notech_ao4 i_1070(.A(n_255794514), .B(in128[45]), .C(n_2941), .D(in128[
		53]), .Z(n_3128));
	notech_ao4 i_1066(.A(n_255494511), .B(in128[52]), .C(n_3122), .D(in128[
		44]), .Z(n_3127));
	notech_ao4 i_1062(.A(n_255194508), .B(in128[51]), .C(n_3122), .D(in128[
		43]), .Z(n_3126));
	notech_ao4 i_1058(.A(n_254894505), .B(in128[41]), .C(n_2941), .D(in128[
		49]), .Z(n_3125));
	notech_ao4 i_1054(.A(n_254594502), .B(in128[48]), .C(n_3122), .D(in128[
		40]), .Z(n_3124));
	notech_nao3 i_4(.A(n_59981), .B(n_254494501), .C(n_59666), .Z(n_3123));
	notech_and4 i_184(.A(n_239994356), .B(n_2945), .C(n_40520), .D(n_2943), 
		.Z(n_3122));
	notech_and2 i_1043(.A(n_3117), .B(n_253594492), .Z(n_3118));
	notech_ao4 i_1042(.A(n_3047), .B(n_40790), .C(n_253194488), .D(n_40758),
		 .Z(n_3117));
	notech_and2 i_1031(.A(n_3112), .B(n_252494481), .Z(n_3113));
	notech_ao4 i_1030(.A(n_3047), .B(n_40789), .C(n_253194488), .D(n_40757),
		 .Z(n_3112));
	notech_and2 i_1019(.A(n_3107), .B(n_251494471), .Z(n_3108));
	notech_ao4 i_1018(.A(n_3047), .B(n_40788), .C(n_253194488), .D(n_40756),
		 .Z(n_3107));
	notech_and2 i_1007(.A(n_3102), .B(n_250494461), .Z(n_3103));
	notech_ao4 i_1006(.A(n_3047), .B(n_40787), .C(n_253194488), .D(n_40755),
		 .Z(n_3102));
	notech_and2 i_995(.A(n_3097), .B(n_249494451), .Z(n_3098));
	notech_ao4 i_994(.A(n_3047), .B(n_40786), .C(n_253194488), .D(n_40754), 
		.Z(n_3097));
	notech_and2 i_983(.A(n_3092), .B(n_248494441), .Z(n_3093));
	notech_ao4 i_982(.A(n_3047), .B(n_40785), .C(n_253194488), .D(n_40753), 
		.Z(n_3092));
	notech_and2 i_971(.A(n_3087), .B(n_247494431), .Z(n_3088));
	notech_ao4 i_970(.A(n_3047), .B(n_40783), .C(n_253194488), .D(n_40751), 
		.Z(n_3087));
	notech_and2 i_954(.A(n_3082), .B(n_246494421), .Z(n_3083));
	notech_ao4 i_953(.A(n_3048), .B(n_40750), .C(n_3047), .D(n_40782), .Z(n_3082
		));
	notech_and2 i_942(.A(n_3077), .B(n_245494411), .Z(n_3078));
	notech_ao4 i_941(.A(n_3048), .B(n_40749), .C(n_3047), .D(n_40781), .Z(n_3077
		));
	notech_and2 i_930(.A(n_3072), .B(n_244494401), .Z(n_3073));
	notech_ao4 i_929(.A(n_3048), .B(n_40748), .C(n_3047), .D(n_40780), .Z(n_3072
		));
	notech_and2 i_918(.A(n_3067), .B(n_243494391), .Z(n_3068));
	notech_ao4 i_917(.A(n_3048), .B(n_40747), .C(n_3047), .D(n_40779), .Z(n_3067
		));
	notech_and2 i_906(.A(n_3062), .B(n_242494381), .Z(n_3063));
	notech_ao4 i_905(.A(n_3048), .B(n_40746), .C(n_3047), .D(n_40778), .Z(n_3062
		));
	notech_and2 i_894(.A(n_3057), .B(n_241494371), .Z(n_3058));
	notech_ao4 i_893(.A(n_3048), .B(n_40745), .C(n_3047), .D(n_40777), .Z(n_3057
		));
	notech_or2 i_146(.A(n_239994356), .B(n_2968), .Z(n_3055));
	notech_or2 i_145(.A(n_40492), .B(n_2168), .Z(n_3053));
	notech_or2 i_147(.A(n_239994356), .B(n_2972), .Z(n_3052));
	notech_and2 i_882(.A(n_3049), .B(n_240494361), .Z(n_3050));
	notech_ao4 i_881(.A(n_3048), .B(n_40744), .C(n_3047), .D(n_40776), .Z(n_3049
		));
	notech_or4 i_186(.A(n_225196458), .B(n_225096459), .C(n_40490), .D(n_239894355
		), .Z(n_3048));
	notech_or2 i_150(.A(n_239994356), .B(n_2965), .Z(n_3047));
	notech_nao3 i_148(.A(n_40487), .B(n_2962), .C(n_239994356), .Z(n_3046)
		);
	notech_or4 i_154(.A(n_40479), .B(n_2961), .C(n_40487), .D(n_239994356), 
		.Z(n_3045));
	notech_ao4 i_871(.A(n_40766), .B(n_238994346), .C(n_40758), .D(n_238894345
		), .Z(n_3042));
	notech_ao4 i_870(.A(n_238794344), .B(n_40782), .C(n_238694343), .D(n_40734
		), .Z(n_3041));
	notech_ao4 i_873(.A(n_40750), .B(n_2173), .C(n_40742), .D(n_2174), .Z(n_3040
		));
	notech_ao4 i_861(.A(n_238894345), .B(n_40756), .C(n_238994346), .D(n_40764
		), .Z(n_3037));
	notech_ao4 i_860(.A(n_238794344), .B(n_40780), .C(n_238694343), .D(n_40732
		), .Z(n_3036));
	notech_ao4 i_863(.A(n_2172), .B(n_40772), .C(n_2174), .D(n_40740), .Z(n_3035
		));
	notech_ao4 i_851(.A(n_238994346), .B(n_40763), .C(n_238894345), .D(n_40755
		), .Z(n_3032));
	notech_ao4 i_850(.A(n_238794344), .B(n_40779), .C(n_238694343), .D(n_40731
		), .Z(n_3031));
	notech_ao4 i_853(.A(n_2173), .B(n_40747), .C(n_2174), .D(n_40739), .Z(n_3030
		));
	notech_ao4 i_841(.A(n_238994346), .B(n_40762), .C(n_238894345), .D(n_40754
		), .Z(n_3027));
	notech_ao4 i_840(.A(n_238794344), .B(n_40778), .C(n_238694343), .D(n_40730
		), .Z(n_3026));
	notech_ao4 i_843(.A(n_2173), .B(n_40746), .C(n_2174), .D(n_40738), .Z(n_3025
		));
	notech_ao4 i_831(.A(n_238694343), .B(n_40729), .C(n_238994346), .D(n_40761
		), .Z(n_3022));
	notech_ao4 i_830(.A(n_238894345), .B(n_40753), .C(n_238794344), .D(n_40777
		), .Z(n_3021));
	notech_ao4 i_833(.A(n_2173), .B(n_40745), .C(n_2174), .D(n_40737), .Z(n_3020
		));
	notech_ao4 i_821(.A(n_238694343), .B(n_40728), .C(n_238894345), .D(n_40752
		), .Z(n_3017));
	notech_ao4 i_820(.A(n_238994346), .B(n_40760), .C(n_238794344), .D(n_40776
		), .Z(n_3016));
	notech_ao4 i_823(.A(n_40768), .B(n_2172), .C(n_2173), .D(n_40744), .Z(n_3015
		));
	notech_ao4 i_811(.A(n_238694343), .B(n_40727), .C(n_238994346), .D(n_40759
		), .Z(n_3012));
	notech_ao4 i_810(.A(n_238894345), .B(n_40751), .C(n_40775), .D(n_238794344
		), .Z(n_3011));
	notech_ao4 i_813(.A(n_2173), .B(n_40743), .C(n_2174), .D(n_40735), .Z(n_3010
		));
	notech_ao4 i_803(.A(n_40758), .B(n_2972), .C(n_40492), .D(n_40892), .Z(n_3008
		));
	notech_and2 i_801(.A(n_3005), .B(n_233394290), .Z(n_3006));
	notech_ao4 i_800(.A(n_2968), .B(n_40774), .C(n_40766), .D(n_2965), .Z(n_3005
		));
	notech_ao4 i_793(.A(n_2972), .B(n_40757), .C(n_40492), .D(n_40893), .Z(n_3003
		));
	notech_and2 i_791(.A(n_3000), .B(n_232594282), .Z(n_3001));
	notech_ao4 i_790(.A(n_2968), .B(n_40773), .C(n_40765), .D(n_2965), .Z(n_3000
		));
	notech_ao4 i_783(.A(n_2972), .B(n_40756), .C(n_40492), .D(n_40936), .Z(n_2998
		));
	notech_and2 i_781(.A(n_2995), .B(n_231794274), .Z(n_2996));
	notech_ao4 i_780(.A(n_2968), .B(n_40772), .C(n_40764), .D(n_2965), .Z(n_2995
		));
	notech_ao4 i_773(.A(n_2972), .B(n_40755), .C(n_40492), .D(n_40935), .Z(n_2993
		));
	notech_and2 i_771(.A(n_2990), .B(n_230994266), .Z(n_2991));
	notech_ao4 i_770(.A(n_2968), .B(n_40771), .C(n_40763), .D(n_2965), .Z(n_2990
		));
	notech_ao4 i_763(.A(n_2972), .B(n_40754), .C(n_40492), .D(n_40934), .Z(n_2988
		));
	notech_and2 i_761(.A(n_2985), .B(n_230194258), .Z(n_2986));
	notech_ao4 i_760(.A(n_2968), .B(n_40770), .C(n_40762), .D(n_2965), .Z(n_2985
		));
	notech_ao4 i_753(.A(n_40753), .B(n_2972), .C(n_40492), .D(n_40927), .Z(n_2983
		));
	notech_and2 i_751(.A(n_2980), .B(n_229394250), .Z(n_2981));
	notech_ao4 i_750(.A(n_2968), .B(n_40769), .C(n_40761), .D(n_2965), .Z(n_2980
		));
	notech_ao4 i_743(.A(n_40752), .B(n_2972), .C(n_40492), .D(n_40928), .Z(n_2978
		));
	notech_and2 i_741(.A(n_2975), .B(n_228594242), .Z(n_2976));
	notech_ao4 i_740(.A(n_2968), .B(n_40768), .C(n_40760), .D(n_2965), .Z(n_2975
		));
	notech_ao4 i_733(.A(n_40751), .B(n_2972), .C(n_40492), .D(n_40894), .Z(n_2973
		));
	notech_nao3 i_32(.A(n_40479), .B(n_2938), .C(n_40487), .Z(n_2972));
	notech_and2 i_730(.A(n_2969), .B(n_227794234), .Z(n_2970));
	notech_ao4 i_729(.A(n_2968), .B(n_40767), .C(n_40759), .D(n_2965), .Z(n_2969
		));
	notech_or4 i_131(.A(n_2937), .B(n_227396436), .C(n_40487), .D(n_2933), .Z
		(n_2968));
	notech_nand2 i_130(.A(n_40479), .B(n_2942), .Z(n_2965));
	notech_nor2 i_19(.A(n_2961), .B(n_40479), .Z(n_2962));
	notech_or2 i_721(.A(n_2937), .B(n_227396436), .Z(n_2961));
	notech_nao3 i_539(.A(\to_acu2_0[0] ), .B(\to_acu2_0[1] ), .C(n_268594642
		), .Z(n_2960));
	notech_nand3 i_65818(.A(n_226796442), .B(n_2957), .C(n_2178), .Z(n_2959)
		);
	notech_and4 i_649(.A(n_40912), .B(n_40911), .C(n_40910), .D(n_40909), .Z
		(n_2957));
	notech_and4 i_643(.A(n_40912), .B(n_40902), .C(n_40901), .D(n_40900), .Z
		(n_2952));
	notech_ao4 i_574(.A(n_226196448), .B(in128[51]), .C(n_2941), .D(in128[59
		]), .Z(n_2949));
	notech_nao3 i_7(.A(n_59981), .B(n_226096449), .C(n_59662), .Z(n_2948));
	notech_and4 i_182(.A(imm_sz[1]), .B(n_2943), .C(n_224696463), .D(n_240094357
		), .Z(n_2947));
	notech_ao4 i_567(.A(n_40591), .B(n_2936), .C(n_2944), .D(n_40592), .Z(n_2945
		));
	notech_nand2 i_563(.A(n_40591), .B(n_40593), .Z(n_2944));
	notech_nor2 i_18(.A(n_40479), .B(n_40490), .Z(n_2943));
	notech_ao3 i_569(.A(n_2937), .B(n_40487), .C(n_227396436), .Z(n_2942));
	notech_and4 i_153(.A(imm_sz[1]), .B(imm_sz[2]), .C(n_40591), .D(n_2940),
		 .Z(n_2941));
	notech_ao3 i_21(.A(n_2938), .B(n_2935), .C(n_40479), .Z(n_2940));
	notech_and2 i_6(.A(n_2937), .B(n_40486), .Z(n_2938));
	notech_xor2 i_2229756(.A(displc[1]), .B(n_2931), .Z(n_2937));
	notech_nand2 i_559(.A(n_40593), .B(n_40592), .Z(n_2936));
	notech_xor2 i_2129755(.A(displc[0]), .B(n_2934), .Z(n_2935));
	notech_xor2 i_216(.A(n_40920), .B(sib_dec), .Z(n_2934));
	notech_nor2 i_2329757(.A(n_225196458), .B(n_225096459), .Z(n_2933));
	notech_nand2 i_276(.A(displc[1]), .B(n_40493), .Z(n_2932));
	notech_nao3 i_26675528(.A(cpl[0]), .B(cpl[1]), .C(n_2025), .Z(n_22894934
		));
	notech_or2 i_29275502(.A(n_3273), .B(n_14051012), .Z(n_22994935));
	notech_or2 i_36575429(.A(n_17551047), .B(n_40853), .Z(n_24494950));
	notech_or4 i_36675428(.A(n_59088), .B(idx_deco[1]), .C(n_223996470), .D(idx_deco
		[0]), .Z(n_24594951));
	notech_nao3 i_36775427(.A(idx_deco[1]), .B(n_39370), .C(n_18051052), .Z(n_24694952
		));
	notech_or4 i_36875426(.A(idx_deco[1]), .B(n_59088), .C(n_39370), .D(n_223996470
		), .Z(n_24794953));
	notech_or2 i_123474562(.A(n_17551047), .B(n_40854), .Z(n_111195806));
	notech_or2 i_124274554(.A(n_17551047), .B(n_40855), .Z(n_111295807));
	notech_and3 i_288793973(.A(n_2226), .B(to_acu1[39]), .C(n_59981), .Z(n_111395808
		));
	notech_nand3 i_24775547(.A(n_2885), .B(inst_deco1[106]), .C(n_59022), .Z
		(n_126695961));
	notech_nand3 i_26275532(.A(n_2885), .B(inst_deco1[113]), .C(n_59022), .Z
		(n_128195976));
	notech_and2 i_302993974(.A(lenpc1[6]), .B(n_59022), .Z(n_131296007));
	notech_and2 i_303093975(.A(lenpc1[7]), .B(n_59022), .Z(n_131396008));
	notech_and2 i_303193976(.A(lenpc1[8]), .B(n_59022), .Z(n_131496009));
	notech_and2 i_303293977(.A(lenpc1[9]), .B(n_59022), .Z(n_131596010));
	notech_and2 i_303393978(.A(lenpc1[10]), .B(n_59022), .Z(n_131696011));
	notech_and2 i_303493979(.A(lenpc1[11]), .B(n_59022), .Z(n_131796012));
	notech_and2 i_303593980(.A(lenpc1[12]), .B(n_59022), .Z(n_131896013));
	notech_and2 i_303693981(.A(lenpc1[13]), .B(n_59022), .Z(n_131996014));
	notech_and2 i_303793982(.A(lenpc1[14]), .B(n_59022), .Z(n_132096015));
	notech_and2 i_303893983(.A(lenpc1[15]), .B(n_59022), .Z(n_132196016));
	notech_and2 i_303993984(.A(lenpc1[16]), .B(n_59022), .Z(n_132296017));
	notech_and2 i_304093985(.A(lenpc1[17]), .B(n_59022), .Z(n_132396018));
	notech_and2 i_304193986(.A(lenpc1[18]), .B(n_59022), .Z(n_132496019));
	notech_and2 i_304293987(.A(lenpc1[19]), .B(n_59022), .Z(n_132596020));
	notech_and2 i_304393988(.A(lenpc1[20]), .B(n_59022), .Z(n_132696021));
	notech_and2 i_304493989(.A(lenpc1[21]), .B(n_59022), .Z(n_132796022));
	notech_and2 i_304593990(.A(lenpc1[22]), .B(n_59022), .Z(n_132896023));
	notech_and2 i_304693991(.A(lenpc1[23]), .B(n_59017), .Z(n_132996024));
	notech_and2 i_304793992(.A(lenpc1[24]), .B(n_59017), .Z(n_133096025));
	notech_and2 i_304893993(.A(lenpc1[25]), .B(n_59017), .Z(n_133196026));
	notech_and2 i_304993994(.A(lenpc1[26]), .B(n_59017), .Z(n_133296027));
	notech_and2 i_305093995(.A(lenpc1[27]), .B(n_59017), .Z(n_133396028));
	notech_and2 i_305193996(.A(lenpc1[28]), .B(n_59017), .Z(n_133496029));
	notech_and2 i_305293997(.A(lenpc1[29]), .B(n_59017), .Z(n_133596030));
	notech_and2 i_305393998(.A(lenpc1[30]), .B(n_59017), .Z(n_133696031));
	notech_and2 i_305493999(.A(lenpc1[31]), .B(n_59017), .Z(n_133796032));
	notech_and3 i_305594000(.A(lenpc2[6]), .B(n_2226), .C(n_59981), .Z(n_133896033
		));
	notech_and3 i_305794001(.A(n_2226), .B(lenpc2[8]), .C(n_59981), .Z(n_133996034
		));
	notech_and3 i_306294002(.A(n_2226), .B(lenpc2[13]), .C(n_59986), .Z(n_134096035
		));
	notech_and3 i_306394003(.A(n_2226), .B(lenpc2[14]), .C(n_59986), .Z(n_134196036
		));
	notech_and3 i_306494004(.A(n_2226), .B(lenpc2[15]), .C(n_59986), .Z(n_134296037
		));
	notech_and3 i_306594005(.A(n_2226), .B(lenpc2[16]), .C(n_59986), .Z(n_134396038
		));
	notech_and3 i_306694006(.A(n_2226), .B(lenpc2[17]), .C(n_59986), .Z(n_134496039
		));
	notech_and3 i_306794007(.A(n_2226), .B(lenpc2[18]), .C(n_59986), .Z(n_134596040
		));
	notech_and3 i_306994008(.A(n_2226), .B(lenpc2[20]), .C(n_59981), .Z(n_134696041
		));
	notech_and3 i_307094009(.A(n_2226), .B(lenpc2[21]), .C(n_59981), .Z(n_134796042
		));
	notech_and3 i_307194010(.A(n_2226), .B(lenpc2[22]), .C(n_59981), .Z(n_134896043
		));
	notech_and3 i_307294011(.A(n_2226), .B(lenpc2[23]), .C(n_59981), .Z(n_134996044
		));
	notech_and3 i_307494012(.A(n_60042), .B(lenpc2[25]), .C(n_59980), .Z(n_135096045
		));
	notech_and3 i_307694013(.A(n_60042), .B(lenpc2[27]), .C(n_59981), .Z(n_135196046
		));
	notech_and3 i_307794014(.A(n_60042), .B(lenpc2[28]), .C(n_59981), .Z(n_135296047
		));
	notech_and3 i_307894015(.A(n_60042), .B(lenpc2[29]), .C(n_59981), .Z(n_135396048
		));
	notech_and3 i_307994016(.A(n_60042), .B(lenpc2[30]), .C(n_59981), .Z(n_135496049
		));
	notech_ao4 i_138074416(.A(n_59010), .B(n_39861), .C(n_59088), .D(n_40722
		), .Z(n_135696051));
	notech_ao4 i_137974417(.A(n_59010), .B(n_39859), .C(n_59088), .D(n_40721
		), .Z(n_135896053));
	notech_ao4 i_137874418(.A(n_59010), .B(n_39857), .C(n_59088), .D(n_40720
		), .Z(n_135996054));
	notech_ao4 i_137774419(.A(n_59010), .B(n_39855), .C(n_59088), .D(n_40719
		), .Z(n_136096055));
	notech_ao4 i_137674420(.A(n_59010), .B(n_39853), .C(n_59088), .D(n_40718
		), .Z(n_136196056));
	notech_ao4 i_137574421(.A(n_59010), .B(n_39851), .C(n_59089), .D(n_40717
		), .Z(n_136296057));
	notech_ao4 i_137474422(.A(n_59010), .B(n_39849), .C(n_59088), .D(n_40716
		), .Z(n_136396058));
	notech_ao4 i_137374423(.A(n_59010), .B(n_39847), .C(n_59089), .D(n_40715
		), .Z(n_136496059));
	notech_ao4 i_137274424(.A(n_59011), .B(n_39845), .C(n_59089), .D(n_40714
		), .Z(n_136596060));
	notech_ao4 i_137174425(.A(n_59011), .B(n_39843), .C(n_59088), .D(n_40713
		), .Z(n_136696061));
	notech_ao4 i_137074426(.A(n_59010), .B(n_39841), .C(n_59088), .D(n_40712
		), .Z(n_136796062));
	notech_ao4 i_136974427(.A(n_59010), .B(n_39839), .C(n_59088), .D(n_40711
		), .Z(n_136896063));
	notech_ao4 i_136874428(.A(n_59010), .B(n_39837), .C(n_59088), .D(n_40710
		), .Z(n_136996064));
	notech_ao4 i_136774429(.A(n_59010), .B(n_39835), .C(n_59084), .D(n_40709
		), .Z(n_137196066));
	notech_ao4 i_136674430(.A(n_59084), .B(n_40708), .C(n_2025), .D(n_14051012
		), .Z(n_137296067));
	notech_mux2 i_20475778(.S(pg_fault), .A(n_59981), .B(n_39063), .Z(n_137396068
		));
	notech_ao4 i_136474432(.A(n_59010), .B(n_39832), .C(n_59084), .D(n_40707
		), .Z(n_137596070));
	notech_ao4 i_136274434(.A(n_59006), .B(n_39830), .C(n_59084), .D(n_40706
		), .Z(n_137796072));
	notech_ao4 i_136174435(.A(n_59006), .B(n_39828), .C(n_59084), .D(n_40705
		), .Z(n_137896073));
	notech_ao4 i_136074436(.A(n_59006), .B(n_39826), .C(n_59084), .D(n_40704
		), .Z(n_137996074));
	notech_ao4 i_135974437(.A(n_59006), .B(n_39824), .C(n_59084), .D(n_40703
		), .Z(n_138096075));
	notech_ao4 i_135874438(.A(n_59006), .B(n_39822), .C(n_59084), .D(n_40702
		), .Z(n_138196076));
	notech_ao4 i_135774439(.A(n_59088), .B(n_40701), .C(n_14051012), .D(n_40937
		), .Z(n_138296077));
	notech_ao4 i_135574441(.A(n_59006), .B(n_39819), .C(n_59088), .D(n_40700
		), .Z(n_138496079));
	notech_ao4 i_135474442(.A(n_59006), .B(n_39817), .C(n_59088), .D(n_40699
		), .Z(n_138596080));
	notech_ao4 i_135374443(.A(n_59010), .B(n_39815), .C(n_59088), .D(n_40698
		), .Z(n_138696081));
	notech_ao4 i_135274444(.A(n_59010), .B(n_39813), .C(n_59084), .D(n_40697
		), .Z(n_138796082));
	notech_ao4 i_135174445(.A(n_59010), .B(n_39811), .C(n_59084), .D(n_40696
		), .Z(n_138896083));
	notech_ao4 i_135074446(.A(n_59006), .B(n_39809), .C(n_59088), .D(n_40695
		), .Z(n_138996084));
	notech_ao4 i_132274474(.A(n_59006), .B(n_39776), .C(n_59084), .D(n_40674
		), .Z(n_139096085));
	notech_ao4 i_132174475(.A(n_59006), .B(n_39774), .C(n_59089), .D(n_40673
		), .Z(n_139196086));
	notech_ao4 i_132074476(.A(n_59006), .B(n_39772), .C(n_59091), .D(n_40672
		), .Z(n_139296087));
	notech_ao4 i_131974477(.A(n_59011), .B(n_39770), .C(n_59091), .D(n_40671
		), .Z(n_139396088));
	notech_ao4 i_131874478(.A(n_59013), .B(n_39768), .C(n_59091), .D(n_40670
		), .Z(n_139496089));
	notech_ao4 i_131774479(.A(n_59013), .B(n_39766), .C(n_59091), .D(n_40669
		), .Z(n_139596090));
	notech_ao4 i_131574481(.A(n_59013), .B(n_39761), .C(n_59091), .D(n_40666
		), .Z(n_139696091));
	notech_ao4 i_131474482(.A(n_59013), .B(n_39759), .C(n_59091), .D(n_40665
		), .Z(n_139796092));
	notech_ao4 i_131374483(.A(n_59013), .B(n_39757), .C(n_59091), .D(n_40664
		), .Z(n_139896093));
	notech_ao4 i_131274484(.A(n_59013), .B(n_39755), .C(n_59091), .D(n_40663
		), .Z(n_139996094));
	notech_ao4 i_131174485(.A(n_59013), .B(n_39753), .C(n_59091), .D(n_40662
		), .Z(n_140096095));
	notech_ao4 i_131074486(.A(n_59013), .B(n_39751), .C(n_59091), .D(n_40661
		), .Z(n_140196096));
	notech_ao4 i_130874488(.A(n_59013), .B(n_39747), .C(n_59091), .D(n_40659
		), .Z(n_140296097));
	notech_ao4 i_130774489(.A(n_59013), .B(n_39745), .C(n_59091), .D(n_40658
		), .Z(n_140396098));
	notech_ao4 i_130674490(.A(n_59013), .B(n_39743), .C(n_59091), .D(n_40657
		), .Z(n_140496099));
	notech_ao4 i_130574491(.A(n_59013), .B(n_39741), .C(n_59091), .D(n_40656
		), .Z(n_140596100));
	notech_ao4 i_130174495(.A(n_59013), .B(n_39733), .C(n_59091), .D(n_40652
		), .Z(n_140696101));
	notech_ao4 i_130074496(.A(n_59013), .B(n_39731), .C(n_59091), .D(n_40651
		), .Z(n_140796102));
	notech_ao4 i_129974497(.A(n_59013), .B(n_39729), .C(n_59089), .D(n_40650
		), .Z(n_140896103));
	notech_ao4 i_129874498(.A(n_59011), .B(n_39727), .C(n_59089), .D(n_40649
		), .Z(n_140996104));
	notech_ao4 i_129774499(.A(n_59011), .B(n_39725), .C(n_59089), .D(n_40648
		), .Z(n_141096105));
	notech_ao4 i_129674500(.A(n_59011), .B(n_39723), .C(n_59089), .D(n_40647
		), .Z(n_141196106));
	notech_ao4 i_129474502(.A(n_59011), .B(n_39719), .C(n_59089), .D(n_40645
		), .Z(n_141296107));
	notech_ao4 i_129374503(.A(n_59011), .B(n_39717), .C(n_59089), .D(n_40644
		), .Z(n_141396108));
	notech_ao4 i_129274504(.A(n_59011), .B(n_39715), .C(n_59089), .D(n_40643
		), .Z(n_141496109));
	notech_ao4 i_129174505(.A(n_59011), .B(n_39713), .C(n_59089), .D(n_40642
		), .Z(n_141596110));
	notech_ao4 i_129074506(.A(n_59011), .B(n_39711), .C(n_59089), .D(n_40641
		), .Z(n_141696111));
	notech_ao4 i_128974507(.A(n_59011), .B(n_39709), .C(n_59089), .D(n_40640
		), .Z(n_141796112));
	notech_ao4 i_128874508(.A(n_59013), .B(n_39707), .C(n_59091), .D(n_40639
		), .Z(n_141896113));
	notech_ao4 i_128774509(.A(n_59011), .B(n_39705), .C(n_59091), .D(n_40638
		), .Z(n_141996114));
	notech_ao4 i_128674510(.A(n_59011), .B(n_39703), .C(n_59089), .D(n_40637
		), .Z(n_142096115));
	notech_ao4 i_128574511(.A(n_59011), .B(n_39701), .C(n_59089), .D(n_40636
		), .Z(n_142196116));
	notech_ao4 i_128474512(.A(n_59011), .B(n_39699), .C(n_59089), .D(n_40635
		), .Z(n_142296117));
	notech_ao4 i_128374513(.A(n_58999), .B(n_39697), .C(n_59089), .D(n_40634
		), .Z(n_142396118));
	notech_ao4 i_128274514(.A(n_58999), .B(n_39695), .C(n_59084), .D(n_40633
		), .Z(n_142496119));
	notech_ao4 i_128174515(.A(n_58999), .B(n_39693), .C(n_59077), .D(n_40632
		), .Z(n_142596120));
	notech_ao4 i_128074516(.A(n_58999), .B(n_39690), .C(n_59077), .D(n_40631
		), .Z(n_142696121));
	notech_ao4 i_127974517(.A(n_58999), .B(n_39688), .C(n_59077), .D(n_40630
		), .Z(n_142796122));
	notech_ao4 i_127874518(.A(n_58999), .B(n_39686), .C(n_59077), .D(n_40629
		), .Z(n_142896123));
	notech_ao4 i_127774519(.A(n_58999), .B(n_39684), .C(n_59077), .D(n_40628
		), .Z(n_142996124));
	notech_ao4 i_127674520(.A(n_59001), .B(n_39682), .C(n_59077), .D(n_40627
		), .Z(n_143096125));
	notech_ao4 i_127574521(.A(n_59001), .B(n_39680), .C(n_59077), .D(n_40626
		), .Z(n_143196126));
	notech_ao4 i_127374523(.A(n_59001), .B(n_39676), .C(n_59077), .D(n_40624
		), .Z(n_143296127));
	notech_ao4 i_127274524(.A(n_59001), .B(n_39674), .C(n_59079), .D(n_40623
		), .Z(n_143396128));
	notech_ao4 i_127174525(.A(n_59001), .B(n_39672), .C(n_59079), .D(n_40622
		), .Z(n_143496129));
	notech_ao4 i_127074526(.A(n_59001), .B(n_39670), .C(n_59079), .D(n_40621
		), .Z(n_143596130));
	notech_ao4 i_126974527(.A(n_59001), .B(n_39668), .C(n_59079), .D(n_40620
		), .Z(n_143696131));
	notech_ao4 i_126874528(.A(n_58999), .B(n_39665), .C(n_59079), .D(n_40619
		), .Z(n_143796132));
	notech_ao4 i_126774529(.A(n_58998), .B(n_39663), .C(n_59079), .D(n_40618
		), .Z(n_143896133));
	notech_ao4 i_126674530(.A(n_58998), .B(n_39660), .C(n_59079), .D(n_40617
		), .Z(n_143996134));
	notech_ao4 i_126574531(.A(n_58998), .B(n_39658), .C(n_59079), .D(n_40616
		), .Z(n_144096135));
	notech_ao4 i_126474532(.A(n_58998), .B(n_39656), .C(n_59076), .D(n_40615
		), .Z(n_144196136));
	notech_ao4 i_126374533(.A(n_58998), .B(n_39654), .C(n_59076), .D(n_40614
		), .Z(n_144296137));
	notech_ao4 i_126274534(.A(n_58998), .B(n_39652), .C(n_59076), .D(n_40613
		), .Z(n_144396138));
	notech_ao4 i_126174535(.A(n_58998), .B(n_39649), .C(n_59076), .D(n_40612
		), .Z(n_144496139));
	notech_ao4 i_126074536(.A(n_58999), .B(n_39647), .C(n_59076), .D(n_40611
		), .Z(n_144596140));
	notech_ao4 i_125974537(.A(n_58999), .B(n_39645), .C(n_59076), .D(n_40610
		), .Z(n_144696141));
	notech_ao4 i_125874538(.A(n_58999), .B(n_39643), .C(n_59076), .D(n_40609
		), .Z(n_144796142));
	notech_ao4 i_125674540(.A(n_58999), .B(n_39639), .C(n_59076), .D(n_40607
		), .Z(n_144896143));
	notech_ao4 i_125574541(.A(n_58999), .B(n_39637), .C(n_59077), .D(n_40606
		), .Z(n_144996144));
	notech_ao4 i_125374543(.A(n_58999), .B(n_39633), .C(n_59077), .D(n_40604
		), .Z(n_145096145));
	notech_ao4 i_125274544(.A(n_58999), .B(n_39631), .C(n_59077), .D(n_40603
		), .Z(n_145196146));
	notech_ao4 i_125174545(.A(n_59001), .B(n_39629), .C(n_59077), .D(n_40602
		), .Z(n_145296147));
	notech_ao4 i_125074546(.A(n_59004), .B(n_39627), .C(n_59077), .D(n_40601
		), .Z(n_145396148));
	notech_ao4 i_124974547(.A(n_59004), .B(n_39625), .C(n_59077), .D(n_40600
		), .Z(n_145496149));
	notech_ao4 i_124874548(.A(n_59004), .B(n_39623), .C(n_59077), .D(n_40599
		), .Z(n_145596150));
	notech_ao4 i_124774549(.A(n_59004), .B(n_39621), .C(n_59077), .D(n_40598
		), .Z(n_145696151));
	notech_ao4 i_124674550(.A(n_59004), .B(n_39619), .C(n_59079), .D(n_40597
		), .Z(n_145796152));
	notech_ao4 i_124574551(.A(n_59004), .B(n_39617), .C(n_59082), .D(n_40596
		), .Z(n_145896153));
	notech_ao4 i_124474552(.A(n_59004), .B(n_39615), .C(n_59082), .D(n_40595
		), .Z(n_145996154));
	notech_or4 i_66774(.A(trig_it), .B(intff), .C(n_39322), .D(n_40945), .Z(n_146096155
		));
	notech_xor2 i_17273982(.A(int_excl[3]), .B(n_1954), .Z(n_146196156));
	notech_and3 i_308494017(.A(n_60042), .B(to_acu2[39]), .C(n_59981), .Z(n_160996304
		));
	notech_ao3 i_5474100(.A(n_59981), .B(in128[8]), .C(n_59662), .Z(n_161096305
		));
	notech_ao3 i_7274082(.A(n_59981), .B(n_58452), .C(n_59662), .Z(n_161196306
		));
	notech_ao3 i_3517(.A(n_1940), .B(n_146196156), .C(n_2027), .Z(n_161296307
		));
	notech_ao3 i_3518(.A(int_excl[5]), .B(n_224496465), .C(n_2027), .Z(n_161596310
		));
	notech_and2 i_3524(.A(ififo_rvect3[0]), .B(n_162496319), .Z(n_161696311)
		);
	notech_and2 i_3529(.A(ififo_rvect3[1]), .B(n_162496319), .Z(n_161796312)
		);
	notech_and2 i_3530(.A(ififo_rvect3[2]), .B(n_162496319), .Z(n_161896313)
		);
	notech_and2 i_3531(.A(ififo_rvect3[3]), .B(n_162496319), .Z(n_161996314)
		);
	notech_and2 i_3532(.A(ififo_rvect3[4]), .B(n_162496319), .Z(n_162096315)
		);
	notech_and2 i_3533(.A(ififo_rvect3[5]), .B(n_162496319), .Z(n_162196316)
		);
	notech_and2 i_3534(.A(ififo_rvect3[6]), .B(n_162496319), .Z(n_162296317)
		);
	notech_and2 i_3535(.A(ififo_rvect3[7]), .B(n_162496319), .Z(n_162396318)
		);
	notech_nand2 i_210222(.A(trig_it), .B(n_39321), .Z(n_162496319));
	notech_or4 i_2874126(.A(int_excl[1]), .B(int_excl[0]), .C(int_excl[3]), 
		.D(int_excl[2]), .Z(n_162796322));
	notech_xor2 i_94073224(.A(int_excl[4]), .B(n_162796322), .Z(n_162896323)
		);
	notech_xor2 i_27994018(.A(pfx_sz[2]), .B(n_171996413), .Z(n_163096325)
		);
	notech_xor2 i_28094019(.A(pfx_sz[3]), .B(n_172096414), .Z(n_163196326)
		);
	notech_xor2 i_28194020(.A(pfx_sz[4]), .B(n_172196415), .Z(n_163296327)
		);
	notech_xor2 i_28394021(.A(int_excl[1]), .B(int_excl[0]), .Z(n_163396328)
		);
	notech_mux2 i_28494022(.S(fpu), .A(n_39059), .B(n_39065), .Z(n_163496329
		));
	notech_mux2 i_28594027(.S(n_1925), .A(n_1757), .B(n_1772), .Z(n_163996334
		));
	notech_and4 i_222715(.A(n_59662), .B(n_2870), .C(n_59986), .D(n_40726), 
		.Z(n_44339));
	notech_and4 i_125694031(.A(n_39060), .B(adz), .C(n_40864), .D(n_39061), 
		.Z(n_164396338));
	notech_xor2 i_26594032(.A(opz[1]), .B(opz[2]), .Z(n_164496339));
	notech_and3 i_125494033(.A(twobyte), .B(\to_acu2_0[16] ), .C(n_41563), .Z
		(n_164596340));
	notech_and4 i_125794034(.A(n_41563), .B(n_169796392), .C(n_1931), .D(n_164496339
		), .Z(n_164696341));
	notech_ao3 i_125594035(.A(opz[2]), .B(n_39060), .C(n_1773), .Z(n_164796342
		));
	notech_or4 i_323174(.A(n_164696341), .B(n_164596340), .C(n_164796342), .D
		(n_164396338), .Z(n_49859));
	notech_or4 i_126894036(.A(adz), .B(\to_acu2_0[73] ), .C(n_169996394), .D
		(n_170196396), .Z(n_164896343));
	notech_or4 i_126594037(.A(twobyte), .B(n_2851), .C(n_40861), .D(n_40468)
		, .Z(n_164996344));
	notech_nao3 i_126694038(.A(n_1931), .B(n_40726), .C(n_169896393), .Z(n_165096345
		));
	notech_or4 i_126794039(.A(n_1931), .B(n_169896393), .C(n_40726), .D(n_1773
		), .Z(n_165196346));
	notech_and4 i_223173(.A(n_164996344), .B(n_165196346), .C(n_164896343), 
		.D(n_165096345), .Z(n_49853));
	notech_or4 i_127794040(.A(n_1931), .B(n_169896393), .C(\to_acu2_0[73] ),
		 .D(n_40865), .Z(n_165296347));
	notech_nand3 i_26694041(.A(n_1773), .B(n_40863), .C(n_40862), .Z(n_165396348
		));
	notech_nao3 i_127694042(.A(n_59991), .B(n_1763), .C(n_2884), .Z(n_165496349
		));
	notech_nao3 i_127894043(.A(opz[0]), .B(n_165396348), .C(n_169896393), .Z
		(n_165596350));
	notech_nand3 i_123172(.A(n_165596350), .B(n_165496349), .C(n_165296347),
		 .Z(n_49847));
	notech_or4 i_132294044(.A(n_59662), .B(pc_req), .C(pg_fault), .D(n_165796352
		), .Z(n_165696351));
	notech_xor2 i_27194045(.A(n_39370), .B(idx_deco[1]), .Z(n_165796352));
	notech_nao3 i_132194046(.A(idx_deco[1]), .B(idx_deco[0]), .C(n_59006), .Z
		(n_165896353));
	notech_nand3 i_222701(.A(n_2025), .B(n_165896353), .C(n_165696351), .Z(n_42953
		));
	notech_or4 i_132594047(.A(n_59662), .B(pc_req), .C(pg_fault), .D(n_1952)
		, .Z(n_165996354));
	notech_nao3 i_132694048(.A(idx_deco[1]), .B(n_39370), .C(n_59006), .Z(n_166096355
		));
	notech_nand3 i_122700(.A(n_2025), .B(n_166096355), .C(n_165996354), .Z(n_42947
		));
	notech_ao4 i_226976(.A(n_40468), .B(n_172296416), .C(n_172396417), .D(n_40724
		), .Z(n_43076));
	notech_ao4 i_323144(.A(n_58117), .B(n_39413), .C(n_39381), .D(n_39576), 
		.Z(n_50758));
	notech_ao4 i_223143(.A(n_58117), .B(n_39412), .C(n_59502), .D(n_39380), 
		.Z(n_50752));
	notech_ao4 i_627217(.A(n_58117), .B(n_40470), .C(n_59502), .D(n_40469), 
		.Z(n_43160));
	notech_ao4 i_69118(.A(n_59666), .B(n_40946), .C(n_1953), .D(n_40476), .Z
		(n_46424));
	notech_ao4 i_16926497(.A(n_58117), .B(n_40424), .C(n_59502), .D(n_40796)
		, .Z(n_42611));
	notech_ao4 i_16226490(.A(n_58122), .B(n_40415), .C(n_59502), .D(n_40789)
		, .Z(n_42569));
	notech_ao4 i_16126489(.A(n_58122), .B(n_40414), .C(n_59502), .D(n_40788)
		, .Z(n_42563));
	notech_ao4 i_16026488(.A(n_58122), .B(n_40413), .C(n_59500), .D(n_40787)
		, .Z(n_42557));
	notech_ao4 i_15826486(.A(n_58122), .B(n_40411), .C(n_59500), .D(n_40785)
		, .Z(n_42545));
	notech_ao4 i_15626484(.A(n_58122), .B(n_40408), .C(n_59500), .D(n_40783)
		, .Z(n_42533));
	notech_ao4 i_15526483(.A(n_58117), .B(n_40407), .C(n_59500), .D(n_40782)
		, .Z(n_42527));
	notech_ao4 i_15026478(.A(n_58117), .B(n_40399), .C(n_59500), .D(n_40777)
		, .Z(n_42497));
	notech_ao4 i_14926477(.A(n_58122), .B(n_40398), .C(n_59502), .D(n_40776)
		, .Z(n_42491));
	notech_ao4 i_14526473(.A(n_58122), .B(n_40394), .C(n_59502), .D(n_40772)
		, .Z(n_42467));
	notech_ao4 i_14426472(.A(n_58122), .B(n_40393), .C(n_59502), .D(n_40771)
		, .Z(n_42461));
	notech_ao4 i_14326471(.A(n_58129), .B(n_40392), .C(n_59505), .D(n_40770)
		, .Z(n_42455));
	notech_ao4 i_14126469(.A(n_58129), .B(n_40390), .C(n_59502), .D(n_40768)
		, .Z(n_42443));
	notech_ao4 i_13026458(.A(n_58129), .B(n_40379), .C(n_59502), .D(n_40757)
		, .Z(n_42377));
	notech_ao4 i_12926457(.A(n_58129), .B(n_40378), .C(n_59502), .D(n_40756)
		, .Z(n_42371));
	notech_ao4 i_12826456(.A(n_58129), .B(n_40377), .C(n_59502), .D(n_40755)
		, .Z(n_42365));
	notech_ao4 i_12726455(.A(n_58129), .B(n_40376), .C(n_59502), .D(n_40754)
		, .Z(n_42359));
	notech_ao4 i_12626454(.A(n_58129), .B(n_40375), .C(n_59502), .D(n_40753)
		, .Z(n_42353));
	notech_ao4 i_12426452(.A(n_58129), .B(n_40372), .C(n_59500), .D(n_40751)
		, .Z(n_42341));
	notech_ao4 i_12326451(.A(n_58129), .B(n_40371), .C(n_59496), .D(n_40750)
		, .Z(n_42335));
	notech_ao4 i_1026338(.A(n_58129), .B(n_40193), .C(n_59496), .D(n_40916),
		 .Z(n_41657));
	notech_ao4 i_626334(.A(n_58133), .B(n_40185), .C(n_59496), .D(n_40875), 
		.Z(n_41633));
	notech_ao4 i_126329(.A(n_58133), .B(n_40173), .C(n_59496), .D(n_40942), 
		.Z(n_41603));
	notech_ao3 i_125194085(.A(n_40861), .B(n_40939), .C(n_2851), .Z(n_169796392
		));
	notech_nao3 i_16994086(.A(n_169796392), .B(n_59991), .C(n_2884), .Z(n_169896393
		));
	notech_nao3 i_20694087(.A(n_40863), .B(n_40862), .C(n_169896393), .Z(n_169996394
		));
	notech_nand3 i_28994089(.A(n_2858), .B(n_2855), .C(n_40865), .Z(n_170196396
		));
	notech_and2 i_3436(.A(pfx_sz[0]), .B(pfx_sz[1]), .Z(n_171996413));
	notech_and3 i_1794106(.A(pfx_sz[0]), .B(pfx_sz[2]), .C(pfx_sz[1]), .Z(n_172096414
		));
	notech_and4 i_28294107(.A(pfx_sz[1]), .B(pfx_sz[0]), .C(pfx_sz[2]), .D(pfx_sz
		[3]), .Z(n_172196415));
	notech_nand2 i_135094108(.A(pfx_sz[0]), .B(n_40724), .Z(n_172296416));
	notech_nand3 i_73299(.A(n_18051052), .B(n_1591), .C(n_111295807), .Z(n_46391
		));
	notech_nand2 i_72093(.A(n_60065), .B(n_1949), .Z(n_44084));
	notech_nand3 i_72219(.A(n_18051052), .B(n_1591), .C(n_111195806), .Z(\nbus_13545[1] 
		));
	notech_nand3 i_71547(.A(n_18051052), .B(n_1591), .C(n_17551047), .Z(\nbus_13539[0] 
		));
	notech_mux2 i_122086(.S(n_61070), .A(lenpc[0]), .B(lenpc1[0]), .Z(lenpc_out
		[0]));
	notech_mux2 i_222087(.S(n_61070), .A(lenpc[1]), .B(lenpc1[1]), .Z(lenpc_out
		[1]));
	notech_mux2 i_322088(.S(n_61070), .A(lenpc[2]), .B(lenpc1[2]), .Z(lenpc_out
		[2]));
	notech_mux2 i_422089(.S(n_61064), .A(lenpc[3]), .B(lenpc1[3]), .Z(lenpc_out
		[3]));
	notech_mux2 i_522090(.S(n_61064), .A(lenpc[4]), .B(lenpc1[4]), .Z(lenpc_out
		[4]));
	notech_mux2 i_622091(.S(n_61064), .A(lenpc[5]), .B(lenpc1[5]), .Z(lenpc_out
		[5]));
	notech_mux2 i_722092(.S(n_61070), .A(lenpc[6]), .B(lenpc1[6]), .Z(lenpc_out
		[6]));
	notech_mux2 i_822093(.S(n_61070), .A(lenpc[7]), .B(lenpc1[7]), .Z(lenpc_out
		[7]));
	notech_mux2 i_922094(.S(n_61070), .A(lenpc[8]), .B(lenpc1[8]), .Z(lenpc_out
		[8]));
	notech_mux2 i_1022095(.S(n_61070), .A(lenpc[9]), .B(lenpc1[9]), .Z(lenpc_out
		[9]));
	notech_mux2 i_1122096(.S(n_61070), .A(lenpc[10]), .B(lenpc1[10]), .Z(lenpc_out
		[10]));
	notech_mux2 i_1222097(.S(n_61070), .A(lenpc[11]), .B(lenpc1[11]), .Z(lenpc_out
		[11]));
	notech_mux2 i_1322098(.S(n_61070), .A(lenpc[12]), .B(lenpc1[12]), .Z(lenpc_out
		[12]));
	notech_mux2 i_1422099(.S(n_61064), .A(lenpc[13]), .B(lenpc1[13]), .Z(lenpc_out
		[13]));
	notech_mux2 i_1522100(.S(n_61064), .A(lenpc[14]), .B(lenpc1[14]), .Z(lenpc_out
		[14]));
	notech_mux2 i_1622101(.S(n_61064), .A(lenpc[15]), .B(lenpc1[15]), .Z(lenpc_out
		[15]));
	notech_mux2 i_1722102(.S(n_61064), .A(lenpc[16]), .B(lenpc1[16]), .Z(lenpc_out
		[16]));
	notech_mux2 i_1822103(.S(n_61064), .A(lenpc[17]), .B(lenpc1[17]), .Z(lenpc_out
		[17]));
	notech_mux2 i_1922104(.S(n_61064), .A(lenpc[18]), .B(lenpc1[18]), .Z(lenpc_out
		[18]));
	notech_mux2 i_2022105(.S(n_61064), .A(lenpc[19]), .B(lenpc1[19]), .Z(lenpc_out
		[19]));
	notech_mux2 i_2122106(.S(n_61064), .A(lenpc[20]), .B(lenpc1[20]), .Z(lenpc_out
		[20]));
	notech_mux2 i_2222107(.S(n_61064), .A(lenpc[21]), .B(lenpc1[21]), .Z(lenpc_out
		[21]));
	notech_mux2 i_2322108(.S(n_61064), .A(lenpc[22]), .B(lenpc1[22]), .Z(lenpc_out
		[22]));
	notech_mux2 i_2422109(.S(n_61064), .A(lenpc[23]), .B(lenpc1[23]), .Z(lenpc_out
		[23]));
	notech_mux2 i_2522110(.S(n_61064), .A(lenpc[24]), .B(lenpc1[24]), .Z(lenpc_out
		[24]));
	notech_mux2 i_2622111(.S(n_61064), .A(lenpc[25]), .B(lenpc1[25]), .Z(lenpc_out
		[25]));
	notech_mux2 i_2722112(.S(n_61070), .A(lenpc[26]), .B(lenpc1[26]), .Z(lenpc_out
		[26]));
	notech_mux2 i_2822113(.S(n_61075), .A(lenpc[27]), .B(lenpc1[27]), .Z(lenpc_out
		[27]));
	notech_mux2 i_2922114(.S(n_61075), .A(lenpc[28]), .B(lenpc1[28]), .Z(lenpc_out
		[28]));
	notech_mux2 i_3022115(.S(n_61075), .A(lenpc[29]), .B(lenpc1[29]), .Z(lenpc_out
		[29]));
	notech_mux2 i_3122116(.S(n_61075), .A(lenpc[30]), .B(lenpc1[30]), .Z(lenpc_out
		[30]));
	notech_mux2 i_3222117(.S(n_61075), .A(lenpc[31]), .B(lenpc1[31]), .Z(lenpc_out
		[31]));
	notech_mux2 i_123118(.S(n_61075), .A(reps0[0]), .B(reps1[0]), .Z(reps[0]
		));
	notech_mux2 i_223119(.S(n_61076), .A(reps0[1]), .B(reps1[1]), .Z(reps[1]
		));
	notech_mux2 i_323120(.S(n_61076), .A(reps0[2]), .B(reps1[2]), .Z(reps[2]
		));
	notech_mux2 i_123121(.S(n_61076), .A(opz0[0]), .B(opz1[0]), .Z(operand_size
		[0]));
	notech_mux2 i_223122(.S(n_61076), .A(opz0[1]), .B(opz1[1]), .Z(operand_size
		[1]));
	notech_mux2 i_323123(.S(n_61076), .A(opz0[2]), .B(opz1[2]), .Z(operand_size
		[2]));
	notech_mux2 i_125267(.S(n_61076), .A(inst_deco[0]), .B(inst_deco1[0]), .Z
		(to_vliw[0]));
	notech_mux2 i_225268(.S(n_61076), .A(inst_deco[1]), .B(inst_deco1[1]), .Z
		(to_vliw[1]));
	notech_mux2 i_325269(.S(n_61075), .A(inst_deco[2]), .B(inst_deco1[2]), .Z
		(to_vliw[2]));
	notech_mux2 i_425270(.S(n_61075), .A(inst_deco[3]), .B(inst_deco1[3]), .Z
		(to_vliw[3]));
	notech_mux2 i_525271(.S(n_61075), .A(inst_deco[4]), .B(inst_deco1[4]), .Z
		(to_vliw[4]));
	notech_mux2 i_625272(.S(n_61070), .A(inst_deco[5]), .B(inst_deco1[5]), .Z
		(to_vliw[5]));
	notech_mux2 i_725273(.S(n_61075), .A(inst_deco[6]), .B(inst_deco1[6]), .Z
		(to_vliw[6]));
	notech_mux2 i_825274(.S(n_61075), .A(inst_deco[7]), .B(inst_deco1[7]), .Z
		(to_vliw[7]));
	notech_mux2 i_925275(.S(n_61075), .A(inst_deco[8]), .B(inst_deco1[8]), .Z
		(to_vliw[8]));
	notech_mux2 i_1025276(.S(n_61075), .A(inst_deco[9]), .B(inst_deco1[9]), 
		.Z(to_vliw[9]));
	notech_mux2 i_1125277(.S(n_61075), .A(inst_deco[10]), .B(inst_deco1[10])
		, .Z(to_vliw[10]));
	notech_mux2 i_1225278(.S(n_61075), .A(inst_deco[11]), .B(inst_deco1[11])
		, .Z(to_vliw[11]));
	notech_mux2 i_1325279(.S(n_61075), .A(inst_deco[12]), .B(inst_deco1[12])
		, .Z(to_vliw[12]));
	notech_mux2 i_1425280(.S(n_61075), .A(inst_deco[13]), .B(inst_deco1[13])
		, .Z(to_vliw[13]));
	notech_mux2 i_1525281(.S(n_61075), .A(inst_deco[14]), .B(inst_deco1[14])
		, .Z(to_vliw[14]));
	notech_mux2 i_1625282(.S(n_61064), .A(inst_deco[15]), .B(inst_deco1[15])
		, .Z(to_vliw[15]));
	notech_mux2 i_1725283(.S(n_61053), .A(inst_deco[16]), .B(inst_deco1[16])
		, .Z(to_vliw[16]));
	notech_mux2 i_1825284(.S(n_61053), .A(inst_deco[17]), .B(inst_deco1[17])
		, .Z(to_vliw[17]));
	notech_mux2 i_1925285(.S(n_61053), .A(inst_deco[18]), .B(inst_deco1[18])
		, .Z(to_vliw[18]));
	notech_mux2 i_2025286(.S(n_61053), .A(inst_deco[19]), .B(inst_deco1[19])
		, .Z(to_vliw[19]));
	notech_mux2 i_2125287(.S(n_61053), .A(inst_deco[20]), .B(inst_deco1[20])
		, .Z(to_vliw[20]));
	notech_mux2 i_2225288(.S(n_61053), .A(inst_deco[21]), .B(inst_deco1[21])
		, .Z(to_vliw[21]));
	notech_mux2 i_2325289(.S(n_61053), .A(inst_deco[22]), .B(inst_deco1[22])
		, .Z(to_vliw[22]));
	notech_mux2 i_2425290(.S(n_61058), .A(inst_deco[23]), .B(inst_deco1[23])
		, .Z(to_vliw[23]));
	notech_mux2 i_2525291(.S(n_61058), .A(inst_deco[24]), .B(inst_deco1[24])
		, .Z(to_vliw[24]));
	notech_mux2 i_2625292(.S(n_61058), .A(inst_deco[25]), .B(inst_deco1[25])
		, .Z(to_vliw[25]));
	notech_mux2 i_2725293(.S(n_61053), .A(inst_deco[26]), .B(inst_deco1[26])
		, .Z(to_vliw[26]));
	notech_mux2 i_2825294(.S(n_61053), .A(inst_deco[27]), .B(inst_deco1[27])
		, .Z(to_vliw[27]));
	notech_mux2 i_2925295(.S(n_61058), .A(inst_deco[28]), .B(inst_deco1[28])
		, .Z(to_vliw[28]));
	notech_mux2 i_3025296(.S(n_61052), .A(inst_deco[29]), .B(inst_deco1[29])
		, .Z(to_vliw[29]));
	notech_mux2 i_3125297(.S(n_61053), .A(inst_deco[30]), .B(inst_deco1[30])
		, .Z(to_vliw[30]));
	notech_mux2 i_3225298(.S(n_61053), .A(inst_deco[31]), .B(inst_deco1[31])
		, .Z(to_vliw[31]));
	notech_mux2 i_3325299(.S(n_61052), .A(inst_deco[32]), .B(inst_deco1[32])
		, .Z(to_vliw[32]));
	notech_mux2 i_3425300(.S(n_61052), .A(inst_deco[33]), .B(inst_deco1[33])
		, .Z(to_vliw[33]));
	notech_mux2 i_3525301(.S(n_61052), .A(inst_deco[34]), .B(inst_deco1[34])
		, .Z(to_vliw[34]));
	notech_mux2 i_3625302(.S(n_61053), .A(inst_deco[35]), .B(inst_deco1[35])
		, .Z(to_vliw[35]));
	notech_mux2 i_3725303(.S(n_61053), .A(inst_deco[36]), .B(inst_deco1[36])
		, .Z(to_vliw[36]));
	notech_mux2 i_3825304(.S(n_61053), .A(inst_deco[37]), .B(inst_deco1[37])
		, .Z(to_vliw[37]));
	notech_mux2 i_3925305(.S(n_61053), .A(inst_deco[38]), .B(inst_deco1[38])
		, .Z(to_vliw[38]));
	notech_mux2 i_4025306(.S(n_61053), .A(inst_deco[39]), .B(inst_deco1[39])
		, .Z(to_vliw[39]));
	notech_mux2 i_4125307(.S(n_61053), .A(inst_deco[40]), .B(inst_deco1[40])
		, .Z(to_vliw[40]));
	notech_mux2 i_4225308(.S(n_61053), .A(inst_deco[41]), .B(inst_deco1[41])
		, .Z(to_vliw[41]));
	notech_mux2 i_4325309(.S(n_61058), .A(inst_deco[42]), .B(inst_deco1[42])
		, .Z(to_vliw[42]));
	notech_mux2 i_4425310(.S(n_61063), .A(inst_deco[43]), .B(inst_deco1[43])
		, .Z(to_vliw[43]));
	notech_mux2 i_4525311(.S(n_61063), .A(inst_deco[44]), .B(inst_deco1[44])
		, .Z(to_vliw[44]));
	notech_mux2 i_4625312(.S(n_61063), .A(inst_deco[45]), .B(inst_deco1[45])
		, .Z(to_vliw[45]));
	notech_mux2 i_4725313(.S(n_61063), .A(inst_deco[46]), .B(inst_deco1[46])
		, .Z(to_vliw[46]));
	notech_mux2 i_4825314(.S(n_61063), .A(inst_deco[47]), .B(inst_deco1[47])
		, .Z(to_vliw[47]));
	notech_mux2 i_4925315(.S(n_61063), .A(inst_deco[48]), .B(inst_deco1[48])
		, .Z(to_vliw[48]));
	notech_mux2 i_5025316(.S(n_61063), .A(inst_deco[49]), .B(inst_deco1[49])
		, .Z(to_vliw[49]));
	notech_mux2 i_5125317(.S(n_61063), .A(inst_deco[50]), .B(inst_deco1[50])
		, .Z(to_vliw[50]));
	notech_mux2 i_5225318(.S(n_61063), .A(inst_deco[51]), .B(inst_deco1[51])
		, .Z(to_vliw[51]));
	notech_mux2 i_5325319(.S(n_61064), .A(inst_deco[52]), .B(inst_deco1[52])
		, .Z(to_vliw[52]));
	notech_mux2 i_5425320(.S(n_61063), .A(inst_deco[53]), .B(inst_deco1[53])
		, .Z(to_vliw[53]));
	notech_mux2 i_5525321(.S(n_61063), .A(inst_deco[54]), .B(inst_deco1[54])
		, .Z(to_vliw[54]));
	notech_mux2 i_5625322(.S(n_61063), .A(inst_deco[55]), .B(inst_deco1[55])
		, .Z(to_vliw[55]));
	notech_mux2 i_5725323(.S(n_61058), .A(inst_deco[56]), .B(inst_deco1[56])
		, .Z(to_vliw[56]));
	notech_mux2 i_5825324(.S(n_61058), .A(inst_deco[57]), .B(inst_deco1[57])
		, .Z(to_vliw[57]));
	notech_mux2 i_5925325(.S(n_61058), .A(inst_deco[58]), .B(inst_deco1[58])
		, .Z(to_vliw[58]));
	notech_mux2 i_6025326(.S(n_61058), .A(inst_deco[59]), .B(inst_deco1[59])
		, .Z(to_vliw[59]));
	notech_mux2 i_6125327(.S(n_61058), .A(inst_deco[60]), .B(inst_deco1[60])
		, .Z(to_vliw[60]));
	notech_mux2 i_6225328(.S(n_61058), .A(inst_deco[61]), .B(inst_deco1[61])
		, .Z(to_vliw[61]));
	notech_mux2 i_6325329(.S(n_61058), .A(inst_deco[62]), .B(inst_deco1[62])
		, .Z(to_vliw[62]));
	notech_mux2 i_6425330(.S(n_61063), .A(inst_deco[63]), .B(inst_deco1[63])
		, .Z(to_vliw[63]));
	notech_mux2 i_6525331(.S(n_61063), .A(inst_deco[64]), .B(inst_deco1[64])
		, .Z(to_vliw[64]));
	notech_mux2 i_6625332(.S(n_61063), .A(inst_deco[65]), .B(inst_deco1[65])
		, .Z(to_vliw[65]));
	notech_mux2 i_6725333(.S(n_61063), .A(inst_deco[66]), .B(inst_deco1[66])
		, .Z(to_vliw[66]));
	notech_mux2 i_6825334(.S(n_61063), .A(inst_deco[67]), .B(inst_deco1[67])
		, .Z(to_vliw[67]));
	notech_mux2 i_6925335(.S(n_61063), .A(inst_deco[68]), .B(inst_deco1[68])
		, .Z(to_vliw[68]));
	notech_mux2 i_7025336(.S(n_61092), .A(inst_deco[69]), .B(inst_deco1[69])
		, .Z(to_vliw[69]));
	notech_mux2 i_7125337(.S(n_61097), .A(inst_deco[70]), .B(inst_deco1[70])
		, .Z(to_vliw[70]));
	notech_mux2 i_7225338(.S(n_61097), .A(inst_deco[71]), .B(inst_deco1[71])
		, .Z(to_vliw[71]));
	notech_mux2 i_7325339(.S(n_61092), .A(inst_deco[72]), .B(inst_deco1[72])
		, .Z(to_vliw[72]));
	notech_mux2 i_7425340(.S(n_61092), .A(inst_deco[73]), .B(inst_deco1[73])
		, .Z(to_vliw[73]));
	notech_mux2 i_7525341(.S(n_61092), .A(inst_deco[74]), .B(inst_deco1[74])
		, .Z(to_vliw[74]));
	notech_mux2 i_7625342(.S(n_61097), .A(inst_deco[75]), .B(inst_deco1[75])
		, .Z(to_vliw[75]));
	notech_mux2 i_7725343(.S(n_61097), .A(inst_deco[76]), .B(inst_deco1[76])
		, .Z(to_vliw[76]));
	notech_mux2 i_7825344(.S(n_61097), .A(inst_deco[77]), .B(inst_deco1[77])
		, .Z(to_vliw[77]));
	notech_mux2 i_7925345(.S(n_61097), .A(inst_deco[78]), .B(inst_deco1[78])
		, .Z(to_vliw[78]));
	notech_mux2 i_8025346(.S(n_61097), .A(inst_deco[79]), .B(inst_deco1[79])
		, .Z(to_vliw[79]));
	notech_mux2 i_8125347(.S(n_61097), .A(inst_deco[80]), .B(inst_deco1[80])
		, .Z(to_vliw[80]));
	notech_mux2 i_8225348(.S(n_61097), .A(inst_deco[81]), .B(inst_deco1[81])
		, .Z(to_vliw[81]));
	notech_mux2 i_8325349(.S(n_61087), .A(inst_deco[82]), .B(inst_deco1[82])
		, .Z(to_vliw[82]));
	notech_mux2 i_8425350(.S(n_61087), .A(inst_deco[83]), .B(inst_deco1[83])
		, .Z(to_vliw[83]));
	notech_mux2 i_8525351(.S(n_61092), .A(inst_deco[84]), .B(inst_deco1[84])
		, .Z(to_vliw[84]));
	notech_mux2 i_8625352(.S(n_61087), .A(inst_deco[85]), .B(inst_deco1[85])
		, .Z(to_vliw[85]));
	notech_mux2 i_8725353(.S(n_61087), .A(inst_deco[86]), .B(inst_deco1[86])
		, .Z(to_vliw[86]));
	notech_mux2 i_8825354(.S(n_61087), .A(inst_deco[87]), .B(inst_deco1[87])
		, .Z(to_vliw[87]));
	notech_mux2 i_8925355(.S(n_61092), .A(inst_deco[88]), .B(inst_deco1[88])
		, .Z(to_vliw[88]));
	notech_mux2 i_9025356(.S(n_61092), .A(inst_deco[89]), .B(inst_deco1[89])
		, .Z(to_vliw[89]));
	notech_mux2 i_9125357(.S(n_61092), .A(inst_deco[90]), .B(inst_deco1[90])
		, .Z(to_vliw[90]));
	notech_mux2 i_9225358(.S(n_61092), .A(inst_deco[91]), .B(inst_deco1[91])
		, .Z(to_vliw[91]));
	notech_mux2 i_9325359(.S(n_61092), .A(inst_deco[92]), .B(inst_deco1[92])
		, .Z(to_vliw[92]));
	notech_mux2 i_9425360(.S(n_61092), .A(inst_deco[93]), .B(inst_deco1[93])
		, .Z(to_vliw[93]));
	notech_mux2 i_9525361(.S(n_61092), .A(inst_deco[94]), .B(inst_deco1[94])
		, .Z(to_vliw[94]));
	notech_mux2 i_9625362(.S(n_61097), .A(inst_deco[95]), .B(inst_deco1[95])
		, .Z(to_vliw[95]));
	notech_mux2 i_9725363(.S(n_61098), .A(inst_deco[96]), .B(inst_deco1[96])
		, .Z(to_vliw[96]));
	notech_mux2 i_9825364(.S(n_61098), .A(inst_deco[97]), .B(inst_deco1[97])
		, .Z(to_vliw[97]));
	notech_mux2 i_9925365(.S(n_61098), .A(inst_deco[98]), .B(inst_deco1[98])
		, .Z(to_vliw[98]));
	notech_mux2 i_10025366(.S(n_61098), .A(inst_deco[99]), .B(inst_deco1[99]
		), .Z(to_vliw[99]));
	notech_mux2 i_10125367(.S(n_61098), .A(inst_deco[100]), .B(inst_deco1[
		100]), .Z(to_vliw[100]));
	notech_mux2 i_10225368(.S(n_61098), .A(inst_deco[101]), .B(inst_deco1[
		101]), .Z(to_vliw[101]));
	notech_mux2 i_10325369(.S(n_61098), .A(inst_deco[102]), .B(inst_deco1[
		102]), .Z(to_vliw[102]));
	notech_mux2 i_10425370(.S(n_61098), .A(inst_deco[103]), .B(inst_deco1[
		103]), .Z(to_vliw[103]));
	notech_mux2 i_10525371(.S(n_61098), .A(inst_deco[104]), .B(inst_deco1[
		104]), .Z(to_vliw[104]));
	notech_mux2 i_10625372(.S(n_61098), .A(inst_deco[105]), .B(inst_deco1[
		105]), .Z(to_vliw[105]));
	notech_mux2 i_10725373(.S(n_61098), .A(inst_deco[106]), .B(inst_deco1[
		106]), .Z(to_vliw[106]));
	notech_mux2 i_10825374(.S(n_61098), .A(inst_deco[107]), .B(inst_deco1[
		107]), .Z(to_vliw[107]));
	notech_mux2 i_10925375(.S(n_61098), .A(inst_deco[108]), .B(inst_deco1[
		108]), .Z(to_vliw[108]));
	notech_mux2 i_11025376(.S(n_61097), .A(inst_deco[109]), .B(inst_deco1[
		109]), .Z(to_vliw[109]));
	notech_mux2 i_11125377(.S(n_61097), .A(inst_deco[110]), .B(inst_deco1[
		110]), .Z(to_vliw[110]));
	notech_mux2 i_11225378(.S(n_61097), .A(inst_deco[111]), .B(inst_deco1[
		111]), .Z(to_vliw[111]));
	notech_mux2 i_11325379(.S(n_61097), .A(inst_deco[112]), .B(inst_deco1[
		112]), .Z(to_vliw[112]));
	notech_mux2 i_11425380(.S(n_61097), .A(inst_deco[113]), .B(inst_deco1[
		113]), .Z(to_vliw[113]));
	notech_mux2 i_11525381(.S(n_61097), .A(inst_deco[114]), .B(inst_deco1[
		114]), .Z(to_vliw[114]));
	notech_mux2 i_11625382(.S(n_61097), .A(inst_deco[115]), .B(inst_deco1[
		115]), .Z(to_vliw[115]));
	notech_mux2 i_11725383(.S(n_61098), .A(inst_deco[116]), .B(inst_deco1[
		116]), .Z(to_vliw[116]));
	notech_mux2 i_11825384(.S(n_61098), .A(inst_deco[117]), .B(inst_deco1[
		117]), .Z(to_vliw[117]));
	notech_mux2 i_11925385(.S(n_61098), .A(inst_deco[118]), .B(inst_deco1[
		118]), .Z(to_vliw[118]));
	notech_mux2 i_12025386(.S(n_61097), .A(inst_deco[119]), .B(inst_deco1[
		119]), .Z(to_vliw[119]));
	notech_mux2 i_12125387(.S(n_61098), .A(inst_deco[120]), .B(inst_deco1[
		120]), .Z(to_vliw[120]));
	notech_mux2 i_12225388(.S(n_61098), .A(inst_deco[121]), .B(inst_deco1[
		121]), .Z(to_vliw[121]));
	notech_mux2 i_12325389(.S(n_61087), .A(inst_deco[122]), .B(inst_deco1[
		122]), .Z(to_vliw[122]));
	notech_mux2 i_12425390(.S(n_61081), .A(inst_deco[123]), .B(inst_deco1[
		123]), .Z(to_vliw[123]));
	notech_mux2 i_12525391(.S(n_61081), .A(inst_deco[124]), .B(inst_deco1[
		124]), .Z(to_vliw[124]));
	notech_mux2 i_12625392(.S(n_61081), .A(inst_deco[125]), .B(inst_deco1[
		125]), .Z(to_vliw[125]));
	notech_mux2 i_12725393(.S(n_61081), .A(inst_deco[126]), .B(inst_deco1[
		126]), .Z(to_vliw[126]));
	notech_mux2 i_12825394(.S(n_61081), .A(inst_deco[127]), .B(inst_deco1[
		127]), .Z(to_vliw[127]));
	notech_mux2 i_125907(.S(n_61081), .A(to_acu0[0]), .B(to_acu1[0]), .Z(to_acu
		[0]));
	notech_mux2 i_225908(.S(n_61081), .A(to_acu0[1]), .B(to_acu1[1]), .Z(to_acu
		[1]));
	notech_mux2 i_325909(.S(n_61086), .A(to_acu0[2]), .B(to_acu1[2]), .Z(to_acu
		[2]));
	notech_mux2 i_425910(.S(n_61086), .A(to_acu0[3]), .B(to_acu1[3]), .Z(to_acu
		[3]));
	notech_mux2 i_525911(.S(n_61086), .A(to_acu0[4]), .B(to_acu1[4]), .Z(to_acu
		[4]));
	notech_mux2 i_625912(.S(n_61081), .A(to_acu0[5]), .B(to_acu1[5]), .Z(to_acu
		[5]));
	notech_mux2 i_725913(.S(n_61081), .A(to_acu0[6]), .B(to_acu1[6]), .Z(to_acu
		[6]));
	notech_mux2 i_825914(.S(n_61081), .A(to_acu0[7]), .B(to_acu1[7]), .Z(to_acu
		[7]));
	notech_mux2 i_925915(.S(n_61076), .A(to_acu0[8]), .B(to_acu1[8]), .Z(to_acu
		[8]));
	notech_mux2 i_1025916(.S(n_61076), .A(to_acu0[9]), .B(to_acu1[9]), .Z(to_acu
		[9]));
	notech_mux2 i_1125917(.S(n_61076), .A(to_acu0[10]), .B(to_acu1[10]), .Z(to_acu
		[10]));
	notech_mux2 i_1225918(.S(n_61076), .A(to_acu0[11]), .B(to_acu1[11]), .Z(to_acu
		[11]));
	notech_mux2 i_1325919(.S(n_61076), .A(to_acu0[12]), .B(to_acu1[12]), .Z(to_acu
		[12]));
	notech_mux2 i_1425920(.S(n_61076), .A(to_acu0[13]), .B(to_acu1[13]), .Z(to_acu
		[13]));
	notech_mux2 i_1525921(.S(n_61076), .A(to_acu0[14]), .B(to_acu1[14]), .Z(to_acu
		[14]));
	notech_mux2 i_1625922(.S(n_61076), .A(to_acu0[15]), .B(to_acu1[15]), .Z(to_acu
		[15]));
	notech_mux2 i_1725923(.S(n_61081), .A(to_acu0[16]), .B(to_acu1[16]), .Z(to_acu
		[16]));
	notech_mux2 i_1825924(.S(n_61081), .A(to_acu0[17]), .B(to_acu1[17]), .Z(to_acu
		[17]));
	notech_mux2 i_1925925(.S(n_61076), .A(to_acu0[18]), .B(to_acu1[18]), .Z(to_acu
		[18]));
	notech_mux2 i_2025926(.S(n_61076), .A(to_acu0[19]), .B(to_acu1[19]), .Z(to_acu
		[19]));
	notech_mux2 i_2125927(.S(n_61076), .A(to_acu0[20]), .B(to_acu1[20]), .Z(to_acu
		[20]));
	notech_mux2 i_2225928(.S(n_61086), .A(to_acu0[21]), .B(to_acu1[21]), .Z(to_acu
		[21]));
	notech_mux2 i_2325929(.S(n_61087), .A(to_acu0[22]), .B(to_acu1[22]), .Z(to_acu
		[22]));
	notech_mux2 i_2425930(.S(n_61087), .A(to_acu0[23]), .B(to_acu1[23]), .Z(to_acu
		[23]));
	notech_mux2 i_2525931(.S(n_61087), .A(to_acu0[24]), .B(to_acu1[24]), .Z(to_acu
		[24]));
	notech_mux2 i_2625932(.S(n_61086), .A(to_acu0[25]), .B(to_acu1[25]), .Z(to_acu
		[25]));
	notech_mux2 i_2725933(.S(n_61087), .A(to_acu0[26]), .B(to_acu1[26]), .Z(to_acu
		[26]));
	notech_mux2 i_2825934(.S(n_61087), .A(to_acu0[27]), .B(to_acu1[27]), .Z(to_acu
		[27]));
	notech_mux2 i_2925935(.S(n_61087), .A(to_acu0[28]), .B(to_acu1[28]), .Z(to_acu
		[28]));
	notech_mux2 i_3025936(.S(n_61087), .A(to_acu0[29]), .B(to_acu1[29]), .Z(to_acu
		[29]));
	notech_mux2 i_3125937(.S(n_61087), .A(to_acu0[30]), .B(to_acu1[30]), .Z(to_acu
		[30]));
	notech_mux2 i_3225938(.S(n_61087), .A(to_acu0[31]), .B(to_acu1[31]), .Z(to_acu
		[31]));
	notech_mux2 i_3325939(.S(n_61087), .A(to_acu0[32]), .B(to_acu1[32]), .Z(to_acu
		[32]));
	notech_mux2 i_3425940(.S(n_61087), .A(to_acu0[33]), .B(to_acu1[33]), .Z(to_acu
		[33]));
	notech_mux2 i_3525941(.S(n_61087), .A(to_acu0[34]), .B(to_acu1[34]), .Z(to_acu
		[34]));
	notech_mux2 i_3625942(.S(n_61086), .A(to_acu0[35]), .B(to_acu1[35]), .Z(to_acu
		[35]));
	notech_mux2 i_3725943(.S(n_61086), .A(to_acu0[36]), .B(to_acu1[36]), .Z(to_acu
		[36]));
	notech_mux2 i_3825944(.S(n_61086), .A(to_acu0[37]), .B(to_acu1[37]), .Z(to_acu
		[37]));
	notech_mux2 i_3925945(.S(n_61086), .A(to_acu0[38]), .B(to_acu1[38]), .Z(to_acu
		[38]));
	notech_mux2 i_4025946(.S(n_61086), .A(to_acu0[39]), .B(to_acu1[39]), .Z(to_acu
		[39]));
	notech_mux2 i_4125947(.S(n_61086), .A(to_acu0[40]), .B(to_acu1[40]), .Z(to_acu
		[40]));
	notech_mux2 i_4225948(.S(n_61086), .A(to_acu0[41]), .B(to_acu1[41]), .Z(to_acu
		[41]));
	notech_mux2 i_4325949(.S(n_61086), .A(to_acu0[42]), .B(to_acu1[42]), .Z(to_acu
		[42]));
	notech_mux2 i_4425950(.S(n_61086), .A(to_acu0[43]), .B(to_acu1[43]), .Z(to_acu
		[43]));
	notech_mux2 i_4525951(.S(n_61086), .A(to_acu0[44]), .B(to_acu1[44]), .Z(to_acu
		[44]));
	notech_mux2 i_4625952(.S(n_61086), .A(to_acu0[45]), .B(to_acu1[45]), .Z(to_acu
		[45]));
	notech_mux2 i_4725953(.S(n_61086), .A(to_acu0[46]), .B(to_acu1[46]), .Z(to_acu
		[46]));
	notech_mux2 i_4825954(.S(n_61086), .A(to_acu0[47]), .B(to_acu1[47]), .Z(to_acu
		[47]));
	notech_mux2 i_4925955(.S(n_61052), .A(to_acu0[48]), .B(to_acu1[48]), .Z(to_acu
		[48]));
	notech_mux2 i_5025956(.S(n_61018), .A(to_acu0[49]), .B(to_acu1[49]), .Z(to_acu
		[49]));
	notech_mux2 i_5125957(.S(n_61018), .A(to_acu0[50]), .B(to_acu1[50]), .Z(to_acu
		[50]));
	notech_mux2 i_5225958(.S(n_61018), .A(to_acu0[51]), .B(to_acu1[51]), .Z(to_acu
		[51]));
	notech_mux2 i_5325959(.S(n_61018), .A(to_acu0[52]), .B(to_acu1[52]), .Z(to_acu
		[52]));
	notech_mux2 i_5425960(.S(n_61018), .A(to_acu0[53]), .B(to_acu1[53]), .Z(to_acu
		[53]));
	notech_mux2 i_5525961(.S(n_61018), .A(to_acu0[54]), .B(to_acu1[54]), .Z(to_acu
		[54]));
	notech_mux2 i_5625962(.S(n_61018), .A(to_acu0[55]), .B(to_acu1[55]), .Z(to_acu
		[55]));
	notech_mux2 i_5725963(.S(n_61019), .A(to_acu0[56]), .B(to_acu1[56]), .Z(to_acu
		[56]));
	notech_mux2 i_5825964(.S(n_61019), .A(to_acu0[57]), .B(to_acu1[57]), .Z(to_acu
		[57]));
	notech_mux2 i_5925965(.S(n_61019), .A(to_acu0[58]), .B(to_acu1[58]), .Z(to_acu
		[58]));
	notech_mux2 i_6025966(.S(n_61018), .A(to_acu0[59]), .B(to_acu1[59]), .Z(to_acu
		[59]));
	notech_mux2 i_6125967(.S(n_61019), .A(to_acu0[60]), .B(to_acu1[60]), .Z(to_acu
		[60]));
	notech_mux2 i_6225968(.S(n_61019), .A(to_acu0[61]), .B(to_acu1[61]), .Z(to_acu
		[61]));
	notech_mux2 i_6325969(.S(n_61018), .A(to_acu0[62]), .B(to_acu1[62]), .Z(to_acu
		[62]));
	notech_mux2 i_6425970(.S(n_61018), .A(to_acu0[63]), .B(to_acu1[63]), .Z(to_acu
		[63]));
	notech_mux2 i_6525971(.S(n_61018), .A(to_acu0[64]), .B(to_acu1[64]), .Z(to_acu
		[64]));
	notech_mux2 i_6625972(.S(n_61013), .A(to_acu0[65]), .B(to_acu1[65]), .Z(to_acu
		[65]));
	notech_mux2 i_6725973(.S(n_61013), .A(to_acu0[66]), .B(to_acu1[66]), .Z(to_acu
		[66]));
	notech_mux2 i_6825974(.S(n_61013), .A(to_acu0[67]), .B(to_acu1[67]), .Z(to_acu
		[67]));
	notech_mux2 i_6925975(.S(n_61018), .A(to_acu0[68]), .B(to_acu1[68]), .Z(to_acu
		[68]));
	notech_mux2 i_7025976(.S(n_61018), .A(to_acu0[69]), .B(to_acu1[69]), .Z(to_acu
		[69]));
	notech_mux2 i_7125977(.S(n_61018), .A(to_acu0[70]), .B(to_acu1[70]), .Z(to_acu
		[70]));
	notech_mux2 i_7225978(.S(n_61018), .A(to_acu0[71]), .B(to_acu1[71]), .Z(to_acu
		[71]));
	notech_mux2 i_7325979(.S(n_61018), .A(to_acu0[72]), .B(to_acu1[72]), .Z(to_acu
		[72]));
	notech_mux2 i_7425980(.S(n_61018), .A(to_acu0[73]), .B(to_acu1[73]), .Z(to_acu
		[73]));
	notech_mux2 i_7525981(.S(n_61018), .A(to_acu0[74]), .B(to_acu1[74]), .Z(to_acu
		[74]));
	notech_mux2 i_7625982(.S(n_61019), .A(to_acu0[75]), .B(to_acu1[75]), .Z(to_acu
		[75]));
	notech_mux2 i_7725983(.S(n_61024), .A(to_acu0[76]), .B(to_acu1[76]), .Z(to_acu
		[76]));
	notech_mux2 i_7825984(.S(n_61024), .A(to_acu0[77]), .B(to_acu1[77]), .Z(to_acu
		[77]));
	notech_mux2 i_7925985(.S(n_61024), .A(to_acu0[78]), .B(to_acu1[78]), .Z(to_acu
		[78]));
	notech_mux2 i_8025986(.S(n_61024), .A(to_acu0[79]), .B(to_acu1[79]), .Z(to_acu
		[79]));
	notech_mux2 i_8125987(.S(n_61024), .A(to_acu0[80]), .B(to_acu1[80]), .Z(to_acu
		[80]));
	notech_mux2 i_8225988(.S(n_61024), .A(to_acu0[81]), .B(to_acu1[81]), .Z(to_acu
		[81]));
	notech_mux2 i_8325989(.S(n_61024), .A(to_acu0[82]), .B(to_acu1[82]), .Z(to_acu
		[82]));
	notech_mux2 i_8425990(.S(n_61024), .A(to_acu0[83]), .B(to_acu1[83]), .Z(to_acu
		[83]));
	notech_mux2 i_8525991(.S(n_61029), .A(to_acu0[84]), .B(to_acu1[84]), .Z(to_acu
		[84]));
	notech_mux2 i_8625992(.S(n_61029), .A(to_acu0[85]), .B(to_acu1[85]), .Z(to_acu
		[85]));
	notech_mux2 i_8725993(.S(n_61024), .A(to_acu0[86]), .B(to_acu1[86]), .Z(to_acu
		[86]));
	notech_mux2 i_8825994(.S(n_61024), .A(to_acu0[87]), .B(to_acu1[87]), .Z(to_acu
		[87]));
	notech_mux2 i_8925995(.S(n_61024), .A(to_acu0[88]), .B(to_acu1[88]), .Z(to_acu
		[88]));
	notech_mux2 i_9025996(.S(n_61019), .A(to_acu0[89]), .B(to_acu1[89]), .Z(to_acu
		[89]));
	notech_mux2 i_9125997(.S(n_61019), .A(to_acu0[90]), .B(to_acu1[90]), .Z(to_acu
		[90]));
	notech_mux2 i_9225998(.S(n_61019), .A(to_acu0[91]), .B(to_acu1[91]), .Z(to_acu
		[91]));
	notech_mux2 i_9325999(.S(n_61019), .A(to_acu0[92]), .B(to_acu1[92]), .Z(to_acu
		[92]));
	notech_mux2 i_9426000(.S(n_61019), .A(to_acu0[93]), .B(to_acu1[93]), .Z(to_acu
		[93]));
	notech_mux2 i_9526001(.S(n_61019), .A(to_acu0[94]), .B(to_acu1[94]), .Z(to_acu
		[94]));
	notech_mux2 i_9626002(.S(n_61019), .A(to_acu0[95]), .B(to_acu1[95]), .Z(to_acu
		[95]));
	notech_mux2 i_9726003(.S(n_61019), .A(to_acu0[96]), .B(to_acu1[96]), .Z(to_acu
		[96]));
	notech_mux2 i_9826004(.S(n_61019), .A(to_acu0[97]), .B(to_acu1[97]), .Z(to_acu
		[97]));
	notech_mux2 i_9926005(.S(n_61024), .A(to_acu0[98]), .B(to_acu1[98]), .Z(to_acu
		[98]));
	notech_mux2 i_10026006(.S(n_61019), .A(to_acu0[99]), .B(to_acu1[99]), .Z
		(to_acu[99]));
	notech_mux2 i_10126007(.S(n_61019), .A(to_acu0[100]), .B(to_acu1[100]), 
		.Z(to_acu[100]));
	notech_mux2 i_10226008(.S(n_61019), .A(to_acu0[101]), .B(to_acu1[101]), 
		.Z(to_acu[101]));
	notech_mux2 i_10326009(.S(n_61013), .A(to_acu0[102]), .B(to_acu1[102]), 
		.Z(to_acu[102]));
	notech_mux2 i_10426010(.S(n_61007), .A(to_acu0[103]), .B(to_acu1[103]), 
		.Z(to_acu[103]));
	notech_mux2 i_10526011(.S(n_61007), .A(to_acu0[104]), .B(to_acu1[104]), 
		.Z(to_acu[104]));
	notech_mux2 i_10626012(.S(n_61007), .A(to_acu0[105]), .B(to_acu1[105]), 
		.Z(to_acu[105]));
	notech_mux2 i_10726013(.S(n_61007), .A(to_acu0[106]), .B(to_acu1[106]), 
		.Z(to_acu[106]));
	notech_mux2 i_10826014(.S(n_61007), .A(to_acu0[107]), .B(to_acu1[107]), 
		.Z(to_acu[107]));
	notech_mux2 i_10926015(.S(n_61007), .A(to_acu0[108]), .B(to_acu1[108]), 
		.Z(to_acu[108]));
	notech_mux2 i_11026016(.S(n_61007), .A(to_acu0[109]), .B(to_acu1[109]), 
		.Z(to_acu[109]));
	notech_mux2 i_11126017(.S(n_61007), .A(to_acu0[110]), .B(to_acu1[110]), 
		.Z(to_acu[110]));
	notech_mux2 i_11226018(.S(n_61007), .A(to_acu0[111]), .B(to_acu1[111]), 
		.Z(to_acu[111]));
	notech_mux2 i_11326019(.S(n_61007), .A(to_acu0[112]), .B(to_acu1[112]), 
		.Z(to_acu[112]));
	notech_mux2 i_11426020(.S(n_61007), .A(to_acu0[113]), .B(to_acu1[113]), 
		.Z(to_acu[113]));
	notech_mux2 i_11526021(.S(n_61007), .A(to_acu0[114]), .B(to_acu1[114]), 
		.Z(to_acu[114]));
	notech_mux2 i_11626022(.S(n_61007), .A(to_acu0[115]), .B(to_acu1[115]), 
		.Z(to_acu[115]));
	notech_mux2 i_11726023(.S(n_61002), .A(to_acu0[116]), .B(to_acu1[116]), 
		.Z(to_acu[116]));
	notech_mux2 i_11826024(.S(n_61002), .A(to_acu0[117]), .B(to_acu1[117]), 
		.Z(to_acu[117]));
	notech_mux2 i_11926025(.S(n_61002), .A(to_acu0[118]), .B(to_acu1[118]), 
		.Z(to_acu[118]));
	notech_mux2 i_12026026(.S(n_61002), .A(to_acu0[119]), .B(to_acu1[119]), 
		.Z(to_acu[119]));
	notech_mux2 i_12126027(.S(n_61002), .A(to_acu0[120]), .B(to_acu1[120]), 
		.Z(to_acu[120]));
	notech_mux2 i_12226028(.S(n_61002), .A(to_acu0[121]), .B(to_acu1[121]), 
		.Z(to_acu[121]));
	notech_mux2 i_12326029(.S(n_61002), .A(to_acu0[122]), .B(to_acu1[122]), 
		.Z(to_acu[122]));
	notech_mux2 i_12426030(.S(n_61007), .A(to_acu0[123]), .B(to_acu1[123]), 
		.Z(to_acu[123]));
	notech_mux2 i_12526031(.S(n_61007), .A(to_acu0[124]), .B(to_acu1[124]), 
		.Z(to_acu[124]));
	notech_mux2 i_12626032(.S(n_61007), .A(to_acu0[125]), .B(to_acu1[125]), 
		.Z(to_acu[125]));
	notech_mux2 i_12726033(.S(n_61002), .A(to_acu0[126]), .B(to_acu1[126]), 
		.Z(to_acu[126]));
	notech_mux2 i_12826034(.S(n_61002), .A(to_acu0[127]), .B(to_acu1[127]), 
		.Z(to_acu[127]));
	notech_mux2 i_12926035(.S(n_61002), .A(to_acu0[128]), .B(to_acu1[128]), 
		.Z(to_acu[128]));
	notech_mux2 i_13026036(.S(n_61007), .A(to_acu0[129]), .B(to_acu1[129]), 
		.Z(to_acu[129]));
	notech_mux2 i_13126037(.S(n_61008), .A(to_acu0[130]), .B(to_acu1[130]), 
		.Z(to_acu[130]));
	notech_mux2 i_13226038(.S(n_61008), .A(to_acu0[131]), .B(to_acu1[131]), 
		.Z(to_acu[131]));
	notech_mux2 i_13326039(.S(n_61013), .A(to_acu0[132]), .B(to_acu1[132]), 
		.Z(to_acu[132]));
	notech_mux2 i_13426040(.S(n_61008), .A(to_acu0[133]), .B(to_acu1[133]), 
		.Z(to_acu[133]));
	notech_mux2 i_13526041(.S(n_61008), .A(to_acu0[134]), .B(to_acu1[134]), 
		.Z(to_acu[134]));
	notech_mux2 i_13626042(.S(n_61008), .A(to_acu0[135]), .B(to_acu1[135]), 
		.Z(to_acu[135]));
	notech_mux2 i_13726043(.S(n_61013), .A(to_acu0[136]), .B(to_acu1[136]), 
		.Z(to_acu[136]));
	notech_mux2 i_13826044(.S(n_61013), .A(to_acu0[137]), .B(to_acu1[137]), 
		.Z(to_acu[137]));
	notech_mux2 i_13926045(.S(n_61013), .A(to_acu0[138]), .B(to_acu1[138]), 
		.Z(to_acu[138]));
	notech_mux2 i_14026046(.S(n_61013), .A(to_acu0[139]), .B(to_acu1[139]), 
		.Z(to_acu[139]));
	notech_mux2 i_14126047(.S(n_61013), .A(to_acu0[140]), .B(to_acu1[140]), 
		.Z(to_acu[140]));
	notech_mux2 i_14226048(.S(n_61013), .A(to_acu0[141]), .B(to_acu1[141]), 
		.Z(to_acu[141]));
	notech_mux2 i_14326049(.S(n_61013), .A(to_acu0[142]), .B(to_acu1[142]), 
		.Z(to_acu[142]));
	notech_mux2 i_14426050(.S(n_61008), .A(to_acu0[143]), .B(to_acu1[143]), 
		.Z(to_acu[143]));
	notech_mux2 i_14526051(.S(n_61008), .A(to_acu0[144]), .B(to_acu1[144]), 
		.Z(to_acu[144]));
	notech_mux2 i_14626052(.S(n_61008), .A(to_acu0[145]), .B(to_acu1[145]), 
		.Z(to_acu[145]));
	notech_mux2 i_14726053(.S(n_61008), .A(to_acu0[146]), .B(to_acu1[146]), 
		.Z(to_acu[146]));
	notech_mux2 i_14826054(.S(n_61008), .A(to_acu0[147]), .B(to_acu1[147]), 
		.Z(to_acu[147]));
	notech_mux2 i_14926055(.S(n_61008), .A(to_acu0[148]), .B(to_acu1[148]), 
		.Z(to_acu[148]));
	notech_mux2 i_15026056(.S(n_61008), .A(to_acu0[149]), .B(to_acu1[149]), 
		.Z(to_acu[149]));
	notech_mux2 i_15126057(.S(n_61008), .A(to_acu0[150]), .B(to_acu1[150]), 
		.Z(to_acu[150]));
	notech_mux2 i_15226058(.S(n_61008), .A(to_acu0[151]), .B(to_acu1[151]), 
		.Z(to_acu[151]));
	notech_mux2 i_15326059(.S(n_61008), .A(to_acu0[152]), .B(to_acu1[152]), 
		.Z(to_acu[152]));
	notech_mux2 i_15426060(.S(n_61008), .A(to_acu0[153]), .B(to_acu1[153]), 
		.Z(to_acu[153]));
	notech_mux2 i_15526061(.S(n_61008), .A(to_acu0[154]), .B(to_acu1[154]), 
		.Z(to_acu[154]));
	notech_mux2 i_15626062(.S(n_61008), .A(to_acu0[155]), .B(to_acu1[155]), 
		.Z(to_acu[155]));
	notech_mux2 i_15726063(.S(n_61042), .A(to_acu0[156]), .B(to_acu1[156]), 
		.Z(to_acu[156]));
	notech_mux2 i_15826064(.S(n_61042), .A(to_acu0[157]), .B(to_acu1[157]), 
		.Z(to_acu[157]));
	notech_mux2 i_15926065(.S(n_61042), .A(to_acu0[158]), .B(to_acu1[158]), 
		.Z(to_acu[158]));
	notech_mux2 i_16026066(.S(n_61042), .A(to_acu0[159]), .B(to_acu1[159]), 
		.Z(to_acu[159]));
	notech_mux2 i_16126067(.S(n_61042), .A(to_acu0[160]), .B(to_acu1[160]), 
		.Z(to_acu[160]));
	notech_mux2 i_16226068(.S(n_61042), .A(to_acu0[161]), .B(to_acu1[161]), 
		.Z(to_acu[161]));
	notech_mux2 i_16326069(.S(n_61042), .A(to_acu0[162]), .B(to_acu1[162]), 
		.Z(to_acu[162]));
	notech_mux2 i_16426070(.S(n_61042), .A(to_acu0[163]), .B(to_acu1[163]), 
		.Z(to_acu[163]));
	notech_mux2 i_16526071(.S(n_61042), .A(to_acu0[164]), .B(to_acu1[164]), 
		.Z(to_acu[164]));
	notech_mux2 i_16626072(.S(n_61042), .A(to_acu0[165]), .B(to_acu1[165]), 
		.Z(to_acu[165]));
	notech_mux2 i_16726073(.S(n_61042), .A(to_acu0[166]), .B(to_acu1[166]), 
		.Z(to_acu[166]));
	notech_mux2 i_16826074(.S(n_61042), .A(to_acu0[167]), .B(to_acu1[167]), 
		.Z(to_acu[167]));
	notech_mux2 i_16926075(.S(n_61042), .A(to_acu0[168]), .B(to_acu1[168]), 
		.Z(to_acu[168]));
	notech_mux2 i_17026076(.S(n_61041), .A(to_acu0[169]), .B(to_acu1[169]), 
		.Z(to_acu[169]));
	notech_mux2 i_17126077(.S(n_61041), .A(to_acu0[170]), .B(to_acu1[170]), 
		.Z(to_acu[170]));
	notech_mux2 i_17226078(.S(n_61041), .A(to_acu0[171]), .B(to_acu1[171]), 
		.Z(to_acu[171]));
	notech_mux2 i_17326079(.S(n_61041), .A(to_acu0[172]), .B(to_acu1[172]), 
		.Z(to_acu[172]));
	notech_mux2 i_17426080(.S(n_61041), .A(to_acu0[173]), .B(to_acu1[173]), 
		.Z(to_acu[173]));
	notech_mux2 i_17526081(.S(n_61041), .A(to_acu0[174]), .B(to_acu1[174]), 
		.Z(to_acu[174]));
	notech_mux2 i_17626082(.S(n_61041), .A(to_acu0[175]), .B(to_acu1[175]), 
		.Z(to_acu[175]));
	notech_mux2 i_17726083(.S(n_61042), .A(to_acu0[176]), .B(to_acu1[176]), 
		.Z(to_acu[176]));
	notech_mux2 i_17826084(.S(n_61042), .A(to_acu0[177]), .B(to_acu1[177]), 
		.Z(to_acu[177]));
	notech_mux2 i_17926085(.S(n_61042), .A(to_acu0[178]), .B(to_acu1[178]), 
		.Z(to_acu[178]));
	notech_mux2 i_18026086(.S(n_61041), .A(to_acu0[179]), .B(to_acu1[179]), 
		.Z(to_acu[179]));
	notech_mux2 i_18126087(.S(n_61041), .A(to_acu0[180]), .B(to_acu1[180]), 
		.Z(to_acu[180]));
	notech_mux2 i_18226088(.S(n_61041), .A(to_acu0[181]), .B(to_acu1[181]), 
		.Z(to_acu[181]));
	notech_mux2 i_18326089(.S(n_61042), .A(to_acu0[182]), .B(to_acu1[182]), 
		.Z(to_acu[182]));
	notech_mux2 i_18426090(.S(n_61052), .A(to_acu0[183]), .B(to_acu1[183]), 
		.Z(to_acu[183]));
	notech_mux2 i_18526091(.S(n_61052), .A(to_acu0[184]), .B(to_acu1[184]), 
		.Z(to_acu[184]));
	notech_mux2 i_18626092(.S(n_61052), .A(to_acu0[185]), .B(to_acu1[185]), 
		.Z(to_acu[185]));
	notech_mux2 i_18726093(.S(n_61052), .A(to_acu0[186]), .B(to_acu1[186]), 
		.Z(to_acu[186]));
	notech_mux2 i_18826094(.S(n_61052), .A(to_acu0[187]), .B(to_acu1[187]), 
		.Z(to_acu[187]));
	notech_mux2 i_18926095(.S(n_61052), .A(to_acu0[188]), .B(to_acu1[188]), 
		.Z(to_acu[188]));
	notech_mux2 i_19026096(.S(n_61052), .A(to_acu0[189]), .B(to_acu1[189]), 
		.Z(to_acu[189]));
	notech_mux2 i_19126097(.S(n_61052), .A(to_acu0[190]), .B(to_acu1[190]), 
		.Z(to_acu[190]));
	notech_mux2 i_19226098(.S(n_61052), .A(to_acu0[191]), .B(to_acu1[191]), 
		.Z(to_acu[191]));
	notech_mux2 i_19326099(.S(n_61052), .A(to_acu0[192]), .B(to_acu1[192]), 
		.Z(to_acu[192]));
	notech_mux2 i_19426100(.S(n_61052), .A(to_acu0[193]), .B(to_acu1[193]), 
		.Z(to_acu[193]));
	notech_mux2 i_19526101(.S(n_61052), .A(to_acu0[194]), .B(to_acu1[194]), 
		.Z(to_acu[194]));
	notech_mux2 i_19626102(.S(n_61052), .A(to_acu0[195]), .B(to_acu1[195]), 
		.Z(to_acu[195]));
	notech_mux2 i_19726103(.S(n_61047), .A(to_acu0[196]), .B(to_acu1[196]), 
		.Z(to_acu[196]));
	notech_mux2 i_19826104(.S(n_61047), .A(to_acu0[197]), .B(to_acu1[197]), 
		.Z(to_acu[197]));
	notech_mux2 i_19926105(.S(n_61047), .A(to_acu0[198]), .B(to_acu1[198]), 
		.Z(to_acu[198]));
	notech_mux2 i_20026106(.S(n_61042), .A(to_acu0[199]), .B(to_acu1[199]), 
		.Z(to_acu[199]));
	notech_mux2 i_20126107(.S(n_61047), .A(to_acu0[200]), .B(to_acu1[200]), 
		.Z(to_acu[200]));
	notech_mux2 i_20226108(.S(n_61047), .A(to_acu0[201]), .B(to_acu1[201]), 
		.Z(to_acu[201]));
	notech_mux2 i_20326109(.S(n_61047), .A(to_acu0[202]), .B(to_acu1[202]), 
		.Z(to_acu[202]));
	notech_mux2 i_20426110(.S(n_61047), .A(to_acu0[203]), .B(to_acu1[203]), 
		.Z(to_acu[203]));
	notech_mux2 i_20526111(.S(n_61047), .A(to_acu0[204]), .B(to_acu1[204]), 
		.Z(to_acu[204]));
	notech_mux2 i_20626112(.S(n_61047), .A(to_acu0[205]), .B(to_acu1[205]), 
		.Z(to_acu[205]));
	notech_mux2 i_20726113(.S(n_61047), .A(to_acu0[206]), .B(to_acu1[206]), 
		.Z(to_acu[206]));
	notech_mux2 i_20826114(.S(n_61047), .A(to_acu0[207]), .B(to_acu1[207]), 
		.Z(to_acu[207]));
	notech_mux2 i_20926115(.S(n_61047), .A(to_acu0[208]), .B(to_acu1[208]), 
		.Z(to_acu[208]));
	notech_mux2 i_21026116(.S(n_61041), .A(to_acu0[209]), .B(to_acu1[209]), 
		.Z(to_acu[209]));
	notech_mux2 i_21126117(.S(n_61030), .A(to_acu0[210]), .B(to_acu1[210]), 
		.Z(to_acu[210]));
	notech_mux2 i_627211(.S(n_61030), .A(\over_seg0[5] ), .B(\over_seg1[5] )
		, .Z(over_seg[5]));
	notech_mux2 i_127608(.S(n_61030), .A(\imm0[0] ), .B(\imm1[0] ), .Z(immediate
		[0]));
	notech_mux2 i_227609(.S(n_61029), .A(\imm0[1] ), .B(\imm1[1] ), .Z(immediate
		[1]));
	notech_mux2 i_327610(.S(n_61029), .A(\imm0[2] ), .B(\imm1[2] ), .Z(immediate
		[2]));
	notech_mux2 i_427611(.S(n_61029), .A(\imm0[3] ), .B(\imm1[3] ), .Z(immediate
		[3]));
	notech_mux2 i_527612(.S(n_61030), .A(\imm0[4] ), .B(\imm1[4] ), .Z(immediate
		[4]));
	notech_mux2 i_627613(.S(n_61030), .A(\imm0[5] ), .B(\imm1[5] ), .Z(immediate
		[5]));
	notech_mux2 i_727614(.S(n_61030), .A(\imm0[6] ), .B(\imm1[6] ), .Z(immediate
		[6]));
	notech_mux2 i_827615(.S(n_61030), .A(\imm0[7] ), .B(\imm1[7] ), .Z(immediate
		[7]));
	notech_mux2 i_927616(.S(n_61030), .A(\imm0[8] ), .B(\imm1[8] ), .Z(immediate
		[8]));
	notech_mux2 i_1027617(.S(n_61030), .A(\imm0[9] ), .B(\imm1[9] ), .Z(immediate
		[9]));
	notech_mux2 i_1127618(.S(n_61030), .A(\imm0[10] ), .B(\imm1[10] ), .Z(immediate
		[10]));
	notech_mux2 i_1227619(.S(n_61029), .A(\imm0[11] ), .B(\imm1[11] ), .Z(immediate
		[11]));
	notech_mux2 i_1327620(.S(n_61029), .A(\imm0[12] ), .B(\imm1[12] ), .Z(immediate
		[12]));
	notech_mux2 i_1427621(.S(n_61029), .A(\imm0[13] ), .B(\imm1[13] ), .Z(immediate
		[13]));
	notech_mux2 i_1527622(.S(n_61029), .A(\imm0[14] ), .B(\imm1[14] ), .Z(immediate
		[14]));
	notech_mux2 i_1627623(.S(n_61029), .A(\imm0[15] ), .B(\imm1[15] ), .Z(immediate
		[15]));
	notech_mux2 i_1727624(.S(n_61029), .A(\imm0[16] ), .B(\imm1[16] ), .Z(immediate
		[16]));
	notech_mux2 i_1827625(.S(n_61029), .A(\imm0[17] ), .B(\imm1[17] ), .Z(immediate
		[17]));
	notech_mux2 i_1927626(.S(n_61029), .A(\imm0[18] ), .B(\imm1[18] ), .Z(immediate
		[18]));
	notech_mux2 i_2027627(.S(n_61029), .A(\imm0[19] ), .B(\imm1[19] ), .Z(immediate
		[19]));
	notech_mux2 i_2127628(.S(n_61029), .A(\imm0[20] ), .B(\imm1[20] ), .Z(immediate
		[20]));
	notech_mux2 i_2227629(.S(n_61029), .A(\imm0[21] ), .B(\imm1[21] ), .Z(immediate
		[21]));
	notech_mux2 i_2327630(.S(n_61029), .A(\imm0[22] ), .B(\imm1[22] ), .Z(immediate
		[22]));
	notech_mux2 i_2427631(.S(n_61029), .A(\imm0[23] ), .B(\imm1[23] ), .Z(immediate
		[23]));
	notech_mux2 i_2527632(.S(n_61030), .A(\imm0[24] ), .B(\imm1[24] ), .Z(immediate
		[24]));
	notech_mux2 i_2627633(.S(n_61036), .A(\imm0[25] ), .B(\imm1[25] ), .Z(immediate
		[25]));
	notech_mux2 i_2727634(.S(n_61036), .A(\imm0[26] ), .B(\imm1[26] ), .Z(immediate
		[26]));
	notech_mux2 i_2827635(.S(n_61036), .A(\imm0[27] ), .B(\imm1[27] ), .Z(immediate
		[27]));
	notech_mux2 i_2927636(.S(n_61036), .A(\imm0[28] ), .B(\imm1[28] ), .Z(immediate
		[28]));
	notech_mux2 i_3027637(.S(n_61036), .A(\imm0[29] ), .B(\imm1[29] ), .Z(immediate
		[29]));
	notech_mux2 i_3127638(.S(n_61036), .A(\imm0[30] ), .B(\imm1[30] ), .Z(immediate
		[30]));
	notech_mux2 i_3227639(.S(n_61041), .A(\imm0[31] ), .B(\imm1[31] ), .Z(immediate
		[31]));
	notech_mux2 i_3327640(.S(n_61041), .A(\imm0[32] ), .B(\imm1[32] ), .Z(immediate
		[32]));
	notech_mux2 i_3427641(.S(n_61041), .A(\imm0[33] ), .B(\imm1[33] ), .Z(immediate
		[33]));
	notech_mux2 i_3527642(.S(n_61041), .A(\imm0[34] ), .B(\imm1[34] ), .Z(immediate
		[34]));
	notech_mux2 i_3627643(.S(n_61041), .A(\imm0[35] ), .B(\imm1[35] ), .Z(immediate
		[35]));
	notech_mux2 i_3727644(.S(n_61041), .A(\imm0[36] ), .B(\imm1[36] ), .Z(immediate
		[36]));
	notech_mux2 i_3827645(.S(n_61041), .A(\imm0[37] ), .B(\imm1[37] ), .Z(immediate
		[37]));
	notech_mux2 i_3927646(.S(n_61030), .A(\imm0[38] ), .B(\imm1[38] ), .Z(immediate
		[38]));
	notech_mux2 i_4027647(.S(n_61030), .A(\imm0[39] ), .B(\imm1[39] ), .Z(immediate
		[39]));
	notech_mux2 i_4127648(.S(n_61030), .A(\imm0[40] ), .B(\imm1[40] ), .Z(immediate
		[40]));
	notech_mux2 i_4227649(.S(n_61030), .A(\imm0[41] ), .B(\imm1[41] ), .Z(immediate
		[41]));
	notech_mux2 i_4327650(.S(n_61030), .A(\imm0[42] ), .B(\imm1[42] ), .Z(immediate
		[42]));
	notech_mux2 i_4427651(.S(n_61030), .A(\imm0[43] ), .B(\imm1[43] ), .Z(immediate
		[43]));
	notech_mux2 i_4527652(.S(n_61030), .A(\imm0[44] ), .B(\imm1[44] ), .Z(immediate
		[44]));
	notech_mux2 i_4627653(.S(n_61036), .A(\imm0[45] ), .B(\imm1[45] ), .Z(immediate
		[45]));
	notech_mux2 i_4727654(.S(n_61036), .A(\imm0[46] ), .B(\imm1[46] ), .Z(immediate
		[46]));
	notech_mux2 i_4827655(.S(n_61036), .A(\imm0[47] ), .B(\imm1[47] ), .Z(immediate
		[47]));
	notech_ao4 i_2830(.A(n_224996460), .B(n_40920), .C(n_40919), .D(n_40594)
		, .Z(n_2931));
	notech_nand3 i_15975796(.A(n_3274), .B(n_60065), .C(n_24794953), .Z(\nbus_13540[0] 
		));
	notech_nand3 i_16075795(.A(n_3274), .B(n_60061), .C(n_24694952), .Z(\nbus_13541[0] 
		));
	notech_nand3 i_17075794(.A(n_60061), .B(n_24594951), .C(n_3274), .Z(\nbus_13534[0] 
		));
	notech_nand3 i_22075793(.A(n_18051052), .B(n_1591), .C(n_24494950), .Z(n_44067
		));
	notech_ao4 i_69106(.A(n_1953), .B(n_40473), .C(n_59666), .D(n_40933), .Z
		(n_46406));
	notech_ao4 i_69110(.A(n_1953), .B(n_40474), .C(n_59662), .D(n_40932), .Z
		(n_46412));
	notech_ao4 i_69114(.A(n_1953), .B(n_40475), .C(n_59662), .D(n_40931), .Z
		(n_46418));
	notech_ao4 i_69122(.A(n_1953), .B(n_40477), .C(n_59662), .D(n_40930), .Z
		(n_46430));
	notech_ao4 i_69126(.A(n_1953), .B(n_40478), .C(n_59657), .D(n_40929), .Z
		(n_46436));
	notech_ao4 i_826125(.A(n_58133), .B(n_39873), .C(n_59496), .D(n_40944), 
		.Z(n_48483));
	notech_ao4 i_526122(.A(n_58133), .B(n_39868), .C(n_59496), .D(n_40940), 
		.Z(n_48465));
	notech_ao4 i_426121(.A(n_58133), .B(n_39867), .C(n_59496), .D(n_40941), 
		.Z(n_48459));
	notech_ao4 i_326120(.A(n_58129), .B(n_39865), .C(n_59496), .D(n_40943), 
		.Z(n_48453));
	notech_nand3 i_12825778(.A(n_60061), .B(n_3273), .C(n_135696051), .Z(n_45834
		));
	notech_nand3 i_12725777(.A(n_60061), .B(n_22994935), .C(n_135896053), .Z
		(n_45828));
	notech_nand3 i_12625776(.A(n_60068), .B(n_3273), .C(n_135996054), .Z(n_45822
		));
	notech_nand3 i_12525775(.A(n_60068), .B(n_22994935), .C(n_136096055), .Z
		(n_45816));
	notech_nand3 i_12425774(.A(n_60068), .B(n_22994935), .C(n_136196056), .Z
		(n_45810));
	notech_nand3 i_12325773(.A(n_60068), .B(n_1448), .C(n_136296057), .Z(n_45804
		));
	notech_nand2 i_12225772(.A(n_60068), .B(n_136396058), .Z(n_45798));
	notech_nand3 i_12125771(.A(n_60068), .B(n_22994935), .C(n_136496059), .Z
		(n_45792));
	notech_nand3 i_12025770(.A(n_60068), .B(n_3273), .C(n_136596060), .Z(n_45786
		));
	notech_nand3 i_11925769(.A(n_60068), .B(n_3273), .C(n_136696061), .Z(n_45780
		));
	notech_nand3 i_11825768(.A(n_60068), .B(n_3273), .C(n_136796062), .Z(n_45774
		));
	notech_nand3 i_11725767(.A(n_60068), .B(n_1448), .C(n_136896063), .Z(n_45768
		));
	notech_nand2 i_11625766(.A(n_60068), .B(n_136996064), .Z(n_45762));
	notech_nand3 i_11525765(.A(n_16151033), .B(n_22894934), .C(n_137196066),
		 .Z(n_45756));
	notech_nand3 i_11425764(.A(n_137296067), .B(n_137396068), .C(n_128195976
		), .Z(n_45750));
	notech_nand3 i_11325763(.A(n_60068), .B(n_2025), .C(n_137596070), .Z(n_45744
		));
	notech_nand2 i_11225762(.A(n_60068), .B(n_137796072), .Z(n_45738));
	notech_nand3 i_11125761(.A(n_60068), .B(n_3273), .C(n_137896073), .Z(n_45732
		));
	notech_nand2 i_11025760(.A(n_60068), .B(n_137996074), .Z(n_45726));
	notech_nand2 i_10925759(.A(n_60068), .B(n_138096075), .Z(n_45720));
	notech_nand3 i_10825758(.A(n_138196076), .B(n_16151033), .C(n_22894934),
		 .Z(n_45714));
	notech_nand3 i_10725757(.A(n_60068), .B(n_138296077), .C(n_126695961), .Z
		(n_45708));
	notech_nand2 i_10625756(.A(n_60066), .B(n_138496079), .Z(n_45702));
	notech_nand3 i_10525755(.A(n_60066), .B(n_1448), .C(n_138596080), .Z(n_45696
		));
	notech_nand3 i_10425754(.A(n_60066), .B(n_1448), .C(n_138696081), .Z(n_45690
		));
	notech_nand3 i_10325753(.A(n_60066), .B(n_1448), .C(n_138796082), .Z(n_45684
		));
	notech_nand3 i_10225752(.A(n_60066), .B(n_1448), .C(n_138896083), .Z(n_45678
		));
	notech_nand2 i_10125751(.A(n_60066), .B(n_138996084), .Z(n_45672));
	notech_nand3 i_8025730(.A(n_60066), .B(n_1448), .C(n_139096085), .Z(n_45546
		));
	notech_nand3 i_7925729(.A(n_60066), .B(n_1448), .C(n_139196086), .Z(n_45540
		));
	notech_nand3 i_7825728(.A(n_60066), .B(n_1448), .C(n_139296087), .Z(n_45534
		));
	notech_nand3 i_7725727(.A(n_60066), .B(n_1448), .C(n_139396088), .Z(n_45528
		));
	notech_nand3 i_7625726(.A(n_60068), .B(n_1448), .C(n_139496089), .Z(n_45522
		));
	notech_nand3 i_7525725(.A(n_60066), .B(n_1448), .C(n_139596090), .Z(n_45516
		));
	notech_nand3 i_7225722(.A(n_60066), .B(n_22994935), .C(n_139696091), .Z(n_45498
		));
	notech_nand3 i_7125721(.A(n_60066), .B(n_3273), .C(n_139796092), .Z(n_45492
		));
	notech_nand3 i_7025720(.A(n_60066), .B(n_3273), .C(n_139896093), .Z(n_45486
		));
	notech_nand3 i_6925719(.A(n_60066), .B(n_22994935), .C(n_139996094), .Z(n_45480
		));
	notech_nand3 i_6825718(.A(n_60054), .B(n_22994935), .C(n_140096095), .Z(n_45474
		));
	notech_nand3 i_6725717(.A(n_60054), .B(n_3273), .C(n_140196096), .Z(n_45468
		));
	notech_nand3 i_6525715(.A(n_60056), .B(n_59028), .C(n_140296097), .Z(n_45456
		));
	notech_nand2 i_6425714(.A(n_60054), .B(n_140396098), .Z(n_45450));
	notech_nand3 i_6325713(.A(n_60054), .B(n_59037), .C(n_140496099), .Z(n_45444
		));
	notech_nand3 i_6225712(.A(n_60054), .B(n_59037), .C(n_140596100), .Z(n_45438
		));
	notech_nand2 i_5825708(.A(n_60054), .B(n_140696101), .Z(n_45414));
	notech_nand3 i_5725707(.A(n_60054), .B(n_22994935), .C(n_140796102), .Z(n_45408
		));
	notech_nand3 i_5625706(.A(n_60056), .B(n_59028), .C(n_140896103), .Z(n_45402
		));
	notech_nand3 i_5525705(.A(n_60056), .B(n_59037), .C(n_140996104), .Z(n_45396
		));
	notech_nand3 i_5425704(.A(n_60056), .B(n_22994935), .C(n_141096105), .Z(n_45390
		));
	notech_nand2 i_5325703(.A(n_60056), .B(n_141196106), .Z(n_45384));
	notech_nand3 i_5125701(.A(n_60056), .B(n_59037), .C(n_141296107), .Z(n_45372
		));
	notech_nand2 i_5025700(.A(n_60056), .B(n_141396108), .Z(n_45366));
	notech_nand2 i_4925699(.A(n_60056), .B(n_141496109), .Z(n_45360));
	notech_nand3 i_4825698(.A(n_60056), .B(n_22994935), .C(n_141596110), .Z(n_45354
		));
	notech_nand3 i_4725697(.A(n_60054), .B(n_59037), .C(n_141696111), .Z(n_45348
		));
	notech_nand3 i_4625696(.A(n_60053), .B(n_59028), .C(n_141796112), .Z(n_45342
		));
	notech_nand2 i_4525695(.A(n_60053), .B(n_141896113), .Z(n_45336));
	notech_nand3 i_4425694(.A(n_60053), .B(n_59028), .C(n_141996114), .Z(n_45330
		));
	notech_nand3 i_4325693(.A(n_60053), .B(n_142096115), .C(n_22994935), .Z(n_45324
		));
	notech_nand2 i_4225692(.A(n_60053), .B(n_142196116), .Z(n_45318));
	notech_nand2 i_4125691(.A(n_60053), .B(n_142296117), .Z(n_45312));
	notech_nand2 i_4025690(.A(n_60053), .B(n_142396118), .Z(n_45306));
	notech_nand3 i_3925689(.A(n_60053), .B(n_59028), .C(n_142496119), .Z(n_45300
		));
	notech_nand3 i_3825688(.A(n_60054), .B(n_59028), .C(n_142596120), .Z(n_45294
		));
	notech_nand2 i_3725687(.A(n_60054), .B(n_142696121), .Z(n_45288));
	notech_nand2 i_3625686(.A(n_60054), .B(n_142796122), .Z(n_45282));
	notech_nand3 i_3525685(.A(n_60054), .B(n_59028), .C(n_142896123), .Z(n_45276
		));
	notech_nand3 i_3425684(.A(n_60054), .B(n_59028), .C(n_142996124), .Z(n_45270
		));
	notech_nand3 i_3325683(.A(n_60054), .B(n_59028), .C(n_143096125), .Z(n_45264
		));
	notech_nand2 i_3225682(.A(n_60054), .B(n_143196126), .Z(n_45258));
	notech_nand3 i_3025680(.A(n_60054), .B(n_59028), .C(n_143296127), .Z(n_45246
		));
	notech_nand2 i_2925679(.A(n_60059), .B(n_143396128), .Z(n_45240));
	notech_nand2 i_2825678(.A(n_60059), .B(n_143496129), .Z(n_45234));
	notech_nand3 i_2725677(.A(n_60059), .B(n_59028), .C(n_143596130), .Z(n_45228
		));
	notech_nand3 i_2625676(.A(n_60059), .B(n_143696131), .C(n_59028), .Z(n_45222
		));
	notech_nand2 i_2525675(.A(n_60059), .B(n_143796132), .Z(n_45216));
	notech_nand2 i_2425674(.A(n_60059), .B(n_143896133), .Z(n_45210));
	notech_nand2 i_2325673(.A(n_60059), .B(n_143996134), .Z(n_45204));
	notech_nand2 i_2225672(.A(n_60059), .B(n_144096135), .Z(n_45198));
	notech_nand2 i_2125671(.A(n_60061), .B(n_144196136), .Z(n_45192));
	notech_nand2 i_2025670(.A(n_60061), .B(n_144296137), .Z(n_45186));
	notech_nand2 i_1925669(.A(n_60061), .B(n_144396138), .Z(n_45180));
	notech_nand2 i_1825668(.A(n_60061), .B(n_144496139), .Z(n_45174));
	notech_nand2 i_1725667(.A(n_60059), .B(n_144596140), .Z(n_45168));
	notech_nand2 i_1625666(.A(n_60059), .B(n_144696141), .Z(n_45162));
	notech_nand2 i_1525665(.A(n_60061), .B(n_144796142), .Z(n_45156));
	notech_nand2 i_1325663(.A(n_60061), .B(n_144896143), .Z(n_45144));
	notech_nand2 i_1225662(.A(n_60059), .B(n_144996144), .Z(n_45138));
	notech_nand2 i_1025660(.A(n_60056), .B(n_145096145), .Z(n_45126));
	notech_nand2 i_925659(.A(n_60056), .B(n_145196146), .Z(n_45120));
	notech_nand3 i_825658(.A(n_60056), .B(n_59037), .C(n_145296147), .Z(n_45114
		));
	notech_nand3 i_725657(.A(n_60056), .B(n_59037), .C(n_145396148), .Z(n_45108
		));
	notech_nand2 i_625656(.A(n_60056), .B(n_145496149), .Z(n_45102));
	notech_nand2 i_525655(.A(n_60056), .B(n_145596150), .Z(n_45096));
	notech_nand3 i_425654(.A(n_60056), .B(n_3273), .C(n_145696151), .Z(n_45090
		));
	notech_nand3 i_325653(.A(n_60056), .B(n_59037), .C(n_145796152), .Z(n_45084
		));
	notech_nand3 i_225652(.A(n_60059), .B(n_145896153), .C(n_59037), .Z(n_45078
		));
	notech_nand2 i_125651(.A(n_145996154), .B(n_60059), .Z(n_45072));
	notech_ao4 i_21126539(.A(n_59496), .B(n_40838), .C(n_58129), .D(n_40467)
		, .Z(n_42863));
	notech_ao4 i_8526413(.A(n_58133), .B(n_40303), .C(n_59496), .D(n_40917),
		 .Z(n_42107));
	notech_and2 i_538(.A(n_39344), .B(n_39342), .Z(n_2926));
	notech_and4 i_541(.A(n_39347), .B(n_39345), .C(n_39350), .D(n_39348), .Z
		(n_2925));
	notech_nao3 i_9(.A(ie), .B(n_40937), .C(ipg_fault), .Z(n_2922));
	notech_nand2 i_525(.A(n_40591), .B(n_40592), .Z(n_2918));
	notech_nand2 i_522(.A(n_61036), .B(term_f), .Z(n_2917));
	notech_nao3 i_520(.A(n_39370), .B(n_40498), .C(idx_deco[1]), .Z(n_2916)
		);
	notech_or2 i_422(.A(n_2870), .B(pc_req), .Z(n_2915));
	notech_and4 i_511(.A(n_60059), .B(n_2837), .C(n_2228), .D(n_2229), .Z(n_2912
		));
	notech_nao3 i_171(.A(n_2224), .B(n_40500), .C(n_2171), .Z(n_2910));
	notech_nao3 i_65873(.A(fsm[0]), .B(n_39374), .C(n_2865), .Z(n_2908));
	notech_nand2 i_22(.A(n_40938), .B(n_2905), .Z(n_2906));
	notech_ao3 i_39(.A(n_2224), .B(n_40500), .C(n_2171), .Z(n_2905));
	notech_or2 i_162(.A(twobyte), .B(fpu), .Z(n_2901));
	notech_and4 i_1129737(.A(n_40894), .B(n_40893), .C(in128[9]), .D(n_2895)
		, .Z(n_2898));
	notech_and2 i_488(.A(n_40892), .B(n_58452), .Z(n_2895));
	notech_or2 i_472(.A(valid_len[3]), .B(valid_len[4]), .Z(n_2890));
	notech_or2 i_24(.A(ipg_fault), .B(n_2887), .Z(n_2888));
	notech_and2 i_6323(.A(n_61036), .B(n_39139), .Z(n_2887));
	notech_ao3 i_3884(.A(n_40937), .B(n_59991), .C(n_2884), .Z(n_2886));
	notech_nand2 i_75073(.A(n_162496319), .B(n_5392), .Z(\nbus_13565[0] ));
	notech_nand2 i_18874163(.A(n_162496319), .B(n_146096155), .Z(\nbus_13535[0] 
		));
	notech_mux2 i_828079(.S(n_162496319), .A(ififo_rvect4[7]), .B(ififo_rvect2
		[7]), .Z(n_44005));
	notech_mux2 i_728078(.S(n_162496319), .A(ififo_rvect4[6]), .B(ififo_rvect2
		[6]), .Z(n_43999));
	notech_mux2 i_628077(.S(n_162496319), .A(ififo_rvect4[5]), .B(ififo_rvect2
		[5]), .Z(n_43993));
	notech_mux2 i_528076(.S(n_162496319), .A(ififo_rvect4[4]), .B(ififo_rvect2
		[4]), .Z(n_43987));
	notech_mux2 i_428075(.S(n_162496319), .A(ififo_rvect4[3]), .B(ififo_rvect2
		[3]), .Z(n_43981));
	notech_mux2 i_328074(.S(n_162496319), .A(ififo_rvect4[2]), .B(ififo_rvect2
		[2]), .Z(n_43975));
	notech_mux2 i_228073(.S(n_162496319), .A(ififo_rvect4[1]), .B(ififo_rvect2
		[1]), .Z(n_43969));
	notech_mux2 i_128072(.S(n_55755), .A(ififo_rvect4[0]), .B(ififo_rvect2[0
		]), .Z(n_43963));
	notech_mux2 i_828039(.S(n_55755), .A(ififo_rvect3[7]), .B(ififo_rvect1[7
		]), .Z(n_42913));
	notech_mux2 i_728038(.S(n_55755), .A(ififo_rvect3[6]), .B(ififo_rvect1[6
		]), .Z(n_42907));
	notech_mux2 i_628037(.S(n_55755), .A(ififo_rvect3[5]), .B(ififo_rvect1[5
		]), .Z(n_42901));
	notech_mux2 i_528036(.S(n_55755), .A(ififo_rvect3[4]), .B(ififo_rvect1[4
		]), .Z(n_42895));
	notech_mux2 i_428035(.S(n_55755), .A(ififo_rvect3[3]), .B(ififo_rvect1[3
		]), .Z(n_42889));
	notech_mux2 i_328034(.S(n_55755), .A(ififo_rvect3[2]), .B(ififo_rvect1[2
		]), .Z(n_42883));
	notech_mux2 i_228033(.S(n_55755), .A(ififo_rvect3[1]), .B(ififo_rvect1[1
		]), .Z(n_42877));
	notech_mux2 i_128032(.S(n_55755), .A(ififo_rvect3[0]), .B(ififo_rvect1[0
		]), .Z(n_42871));
	notech_mux2 i_828047(.S(n_55755), .A(ififo_rvect2[7]), .B(ivect[7]), .Z(n_44409
		));
	notech_mux2 i_728046(.S(n_55755), .A(ififo_rvect2[6]), .B(ivect[6]), .Z(n_44403
		));
	notech_mux2 i_628045(.S(n_162496319), .A(ififo_rvect2[5]), .B(ivect[5]),
		 .Z(n_44397));
	notech_mux2 i_528044(.S(n_55755), .A(ififo_rvect2[4]), .B(ivect[4]), .Z(n_44391
		));
	notech_mux2 i_428043(.S(n_55755), .A(ififo_rvect2[3]), .B(ivect[3]), .Z(n_44385
		));
	notech_mux2 i_328042(.S(n_55755), .A(ififo_rvect2[2]), .B(ivect[2]), .Z(n_44379
		));
	notech_mux2 i_228041(.S(n_55755), .A(ififo_rvect2[1]), .B(ivect[1]), .Z(n_44373
		));
	notech_mux2 i_128040(.S(n_55755), .A(ififo_rvect2[0]), .B(ivect[0]), .Z(n_44367
		));
	notech_nao3 i_527192(.A(n_162896323), .B(n_1940), .C(n_2027), .Z(n_49899
		));
	notech_ao4 i_3825432(.A(n_59500), .B(n_40632), .C(n_58133), .D(n_39477),
		 .Z(n_50143));
	notech_ao4 i_3325427(.A(n_59500), .B(n_40627), .C(n_58133), .D(n_39470),
		 .Z(n_50113));
	notech_ao4 i_2625420(.A(n_59500), .B(n_40620), .C(n_58129), .D(n_39459),
		 .Z(n_50071));
	notech_ao4 i_2525419(.A(n_59500), .B(n_40619), .C(n_58123), .D(n_39458),
		 .Z(n_50065));
	notech_ao4 i_2425418(.A(n_59500), .B(n_40618), .C(n_58123), .D(n_39456),
		 .Z(n_50059));
	notech_ao4 i_2325417(.A(n_59496), .B(n_40617), .C(n_58135), .D(n_39455),
		 .Z(n_50053));
	notech_ao4 i_1925413(.A(n_59496), .B(n_40613), .C(n_58135), .D(n_39449),
		 .Z(n_50029));
	notech_ao4 i_19626313(.A(n_59500), .B(n_40823), .C(n_58135), .D(n_40149)
		, .Z(n_49611));
	notech_ao4 i_16526282(.A(n_59500), .B(n_40792), .C(n_58123), .D(n_40105)
		, .Z(n_49425));
	notech_ao4 i_16426281(.A(n_59500), .B(n_40791), .C(n_58123), .D(n_40104)
		, .Z(n_49419));
	notech_ao4 i_15726274(.A(n_59522), .B(n_40784), .C(n_58123), .D(n_40097)
		, .Z(n_49377));
	notech_ao4 i_15326270(.A(n_58123), .B(n_40093), .C(n_59545), .D(n_40780)
		, .Z(n_49353));
	notech_ao4 i_15226269(.A(n_59545), .B(n_40779), .C(n_58123), .D(n_40092)
		, .Z(n_49347));
	notech_ao4 i_15126268(.A(n_58129), .B(n_40091), .C(n_59545), .D(n_40778)
		, .Z(n_49341));
	notech_ao4 i_12526242(.A(n_58129), .B(n_40057), .C(n_59545), .D(n_40752)
		, .Z(n_49185));
	notech_ao4 i_12126238(.A(n_58129), .B(n_40051), .C(n_59545), .D(n_40748)
		, .Z(n_49161));
	notech_ao4 i_11926236(.A(n_58129), .B(n_40048), .C(n_59541), .D(n_40746)
		, .Z(n_49149));
	notech_ao4 i_11826235(.A(n_58129), .B(n_40047), .C(n_59541), .D(n_40745)
		, .Z(n_49143));
	notech_ao4 i_11726234(.A(n_58135), .B(n_40045), .C(n_59541), .D(n_40744)
		, .Z(n_49137));
	notech_ao4 i_11626233(.A(n_58135), .B(n_40044), .C(n_59541), .D(n_40743)
		, .Z(n_49131));
	notech_ao4 i_11526232(.A(n_58135), .B(n_40042), .C(n_59541), .D(n_40742)
		, .Z(n_49125));
	notech_ao4 i_10926226(.A(n_59545), .B(n_40736), .C(n_58129), .D(n_40033)
		, .Z(n_49089));
	notech_ao4 i_10726224(.A(n_59545), .B(n_40734), .C(n_58129), .D(n_40030)
		, .Z(n_49077));
	notech_ao4 i_10626223(.A(n_59545), .B(n_40733), .C(n_58150), .D(n_40028)
		, .Z(n_49071));
	notech_ao4 i_10526222(.A(n_59547), .B(n_40732), .C(n_58173), .D(n_40026)
		, .Z(n_49065));
	notech_ao4 i_10426221(.A(n_59545), .B(n_40731), .C(n_58173), .D(n_40024)
		, .Z(n_49059));
	notech_ao4 i_10326220(.A(n_59545), .B(n_40730), .C(n_58173), .D(n_40022)
		, .Z(n_49053));
	notech_ao4 i_10226219(.A(n_59545), .B(n_40729), .C(n_58173), .D(n_40020)
		, .Z(n_49047));
	notech_ao4 i_10126218(.A(n_59545), .B(n_40728), .C(n_58173), .D(n_40018)
		, .Z(n_49041));
	notech_ao4 i_10026217(.A(n_59545), .B(n_40727), .C(n_58173), .D(n_40016)
		, .Z(n_49035));
	notech_ao4 i_9926216(.A(n_59545), .B(n_40892), .C(n_58173), .D(n_40014),
		 .Z(n_49029));
	notech_ao4 i_9826215(.A(n_59541), .B(n_40893), .C(n_58173), .D(n_40012),
		 .Z(n_49023));
	notech_ao4 i_9726214(.A(n_59539), .B(n_40936), .C(n_58173), .D(n_40010),
		 .Z(n_49017));
	notech_ao4 i_9626213(.A(n_59539), .B(n_40935), .C(n_58173), .D(n_40008),
		 .Z(n_49011));
	notech_ao4 i_9526212(.A(n_59539), .B(n_40934), .C(n_58175), .D(n_40006),
		 .Z(n_49005));
	notech_ao4 i_9426211(.A(n_59539), .B(n_40927), .C(n_58175), .D(n_40004),
		 .Z(n_48999));
	notech_ao4 i_9326210(.A(n_59539), .B(n_40928), .C(n_58175), .D(n_40002),
		 .Z(n_48993));
	notech_ao4 i_9226209(.A(n_59539), .B(n_40894), .C(n_58175), .D(n_40000),
		 .Z(n_48987));
	notech_ao4 i_9126208(.A(n_59539), .B(n_40947), .C(n_58175), .D(n_39998),
		 .Z(n_48981));
	notech_ao4 i_8526202(.A(n_58173), .B(n_39988), .C(n_59539), .D(n_40917),
		 .Z(n_48945));
	notech_ao4 i_21026538(.A(n_59539), .B(n_40837), .C(n_58173), .D(n_40466)
		, .Z(n_42857));
	notech_ao4 i_20926537(.A(n_59539), .B(n_40836), .C(n_58173), .D(n_40465)
		, .Z(n_42851));
	notech_ao4 i_20726535(.A(n_59541), .B(n_40834), .C(n_58175), .D(n_40463)
		, .Z(n_42839));
	notech_ao4 i_20526533(.A(n_59541), .B(n_40832), .C(n_58173), .D(n_40461)
		, .Z(n_42827));
	notech_ao4 i_20426532(.A(n_59541), .B(n_40831), .C(n_58169), .D(n_40460)
		, .Z(n_42821));
	notech_ao4 i_20326531(.A(n_59541), .B(n_40830), .C(n_58167), .D(n_40459)
		, .Z(n_42815));
	notech_ao4 i_20226530(.A(n_59541), .B(n_40829), .C(n_58167), .D(n_40458)
		, .Z(n_42809));
	notech_ao4 i_20026528(.A(n_59539), .B(n_40827), .C(n_58169), .D(n_40456)
		, .Z(n_42797));
	notech_ao4 i_9426422(.A(n_59539), .B(n_40927), .C(n_58169), .D(n_40321),
		 .Z(n_42161));
	notech_ao4 i_9226420(.A(n_59541), .B(n_40894), .C(n_58169), .D(n_40316),
		 .Z(n_42149));
	notech_ao4 i_9026418(.A(n_59541), .B(n_40856), .C(n_58167), .D(n_40311),
		 .Z(n_42137));
	notech_ao4 i_8926417(.A(n_59541), .B(n_40857), .C(n_58167), .D(n_40310),
		 .Z(n_42131));
	notech_ao4 i_8826416(.A(n_59547), .B(n_40858), .C(n_58167), .D(n_40308),
		 .Z(n_42125));
	notech_ao4 i_8726415(.A(n_59552), .B(n_40859), .C(n_58167), .D(n_40306),
		 .Z(n_42119));
	notech_ao4 i_8626414(.A(n_59552), .B(n_40918), .C(n_58167), .D(n_40305),
		 .Z(n_42113));
	notech_ao4 i_8426412(.A(n_59552), .B(n_40839), .C(n_58169), .D(n_40301),
		 .Z(n_42101));
	notech_ao4 i_8326411(.A(n_59552), .B(n_40920), .C(n_58169), .D(n_40299),
		 .Z(n_42095));
	notech_ao4 i_8226410(.A(n_59552), .B(n_40919), .C(n_58169), .D(n_40297),
		 .Z(n_42089));
	notech_ao4 i_8126409(.A(n_59550), .B(n_40873), .C(n_58169), .D(n_40296),
		 .Z(n_42083));
	notech_ao4 i_8026408(.A(n_59550), .B(n_40889), .C(n_58169), .D(n_40294),
		 .Z(n_42077));
	notech_ao4 i_7926407(.A(n_59550), .B(n_40891), .C(n_58169), .D(n_40292),
		 .Z(n_42071));
	notech_ao4 i_7826406(.A(n_59550), .B(n_40840), .C(n_58169), .D(n_40291),
		 .Z(n_42065));
	notech_ao4 i_7726405(.A(n_59550), .B(n_40862), .C(n_58169), .D(n_40289),
		 .Z(n_42059));
	notech_ao4 i_7626404(.A(n_59552), .B(n_40855), .C(n_58169), .D(n_40288),
		 .Z(n_42053));
	notech_ao4 i_7526403(.A(n_59552), .B(n_40865), .C(n_58169), .D(n_40287),
		 .Z(n_42047));
	notech_ao4 i_7426402(.A(n_59552), .B(n_40864), .C(n_58180), .D(n_40286),
		 .Z(n_42041));
	notech_ao4 i_7326401(.A(n_59556), .B(n_40863), .C(n_58180), .D(n_40285),
		 .Z(n_42035));
	notech_ao4 i_7226400(.A(n_59552), .B(n_40853), .C(n_58180), .D(n_40284),
		 .Z(n_42029));
	notech_ao4 i_7126399(.A(n_59552), .B(n_40854), .C(n_58180), .D(n_40283),
		 .Z(n_42023));
	notech_ao4 i_7026398(.A(n_59552), .B(n_40914), .C(n_58180), .D(n_40282),
		 .Z(n_42017));
	notech_ao4 i_6926397(.A(n_59552), .B(n_40906), .C(n_58180), .D(n_40280),
		 .Z(n_42011));
	notech_ao4 i_6826396(.A(n_59552), .B(n_40841), .C(n_58178), .D(n_40278),
		 .Z(n_42005));
	notech_ao4 i_6726395(.A(n_59552), .B(n_40842), .C(n_58180), .D(n_40277),
		 .Z(n_41999));
	notech_ao4 i_6626394(.A(n_59550), .B(n_40843), .C(n_58180), .D(n_40276),
		 .Z(n_41993));
	notech_ao4 i_6526393(.A(n_59547), .B(n_40844), .C(n_58180), .D(n_40275),
		 .Z(n_41987));
	notech_ao4 i_6426392(.A(n_59547), .B(n_40845), .C(n_58184), .D(n_40274),
		 .Z(n_41981));
	notech_ao4 i_6226390(.A(n_59547), .B(n_40890), .C(n_58184), .D(n_40272),
		 .Z(n_41969));
	notech_ao4 i_6126389(.A(n_59547), .B(n_40846), .C(n_58184), .D(n_40271),
		 .Z(n_41963));
	notech_ao4 i_6026388(.A(n_59547), .B(n_40872), .C(n_58184), .D(n_40270),
		 .Z(n_41957));
	notech_ao4 i_5826386(.A(n_59547), .B(n_40866), .C(n_58184), .D(n_40268),
		 .Z(n_41945));
	notech_ao4 i_5726385(.A(n_59547), .B(n_40860), .C(n_58180), .D(n_40266),
		 .Z(n_41939));
	notech_ao4 i_5626384(.A(n_59547), .B(n_40870), .C(n_58180), .D(n_40265),
		 .Z(n_41933));
	notech_ao4 i_5326381(.A(n_59547), .B(n_40867), .C(n_58180), .D(n_40262),
		 .Z(n_41915));
	notech_ao4 i_5026378(.A(n_59547), .B(n_40847), .C(n_58180), .D(n_40259),
		 .Z(n_41897));
	notech_ao4 i_4926377(.A(n_59550), .B(n_40874), .C(n_58180), .D(n_40258),
		 .Z(n_41891));
	notech_ao4 i_4526373(.A(n_59550), .B(n_40885), .C(n_58178), .D(n_40254),
		 .Z(n_41867));
	notech_ao4 i_4426372(.A(n_59550), .B(n_40883), .C(n_58175), .D(n_40253),
		 .Z(n_41861));
	notech_ao4 i_2326351(.A(n_59550), .B(n_40905), .C(n_58175), .D(n_40219),
		 .Z(n_41735));
	notech_ao4 i_2226350(.A(n_59550), .B(n_40903), .C(n_58175), .D(n_40217),
		 .Z(n_41729));
	notech_ao4 i_1926347(.A(n_59547), .B(n_40899), .C(n_58178), .D(n_40211),
		 .Z(n_41711));
	notech_ao4 i_1626344(.A(n_59547), .B(n_40895), .C(n_58178), .D(n_40205),
		 .Z(n_41693));
	notech_ao4 i_1526343(.A(n_59550), .B(n_40896), .C(n_58175), .D(n_40203),
		 .Z(n_41687));
	notech_ao4 i_1426342(.A(n_59550), .B(n_40897), .C(n_58175), .D(n_40201),
		 .Z(n_41681));
	notech_ao4 i_1326341(.A(n_59550), .B(n_40900), .C(n_58175), .D(n_40199),
		 .Z(n_41675));
	notech_ao4 i_1226340(.A(n_59539), .B(n_40915), .C(n_58175), .D(n_40197),
		 .Z(n_41669));
	notech_and2 i_5(.A(n_40937), .B(n_59991), .Z(n_2885));
	notech_ao3 i_3074124(.A(n_59991), .B(in128[81]), .C(n_59648), .Z(n_73850748
		));
	notech_ao3 i_3274122(.A(n_59991), .B(in128[22]), .C(n_59648), .Z(n_73650746
		));
	notech_ao3 i_3474120(.A(n_59991), .B(in128[82]), .C(n_59648), .Z(n_73450744
		));
	notech_ao3 i_3874116(.A(n_59992), .B(in128[12]), .C(n_59648), .Z(n_73050740
		));
	notech_ao3 i_3974115(.A(n_59992), .B(in128[83]), .C(n_59648), .Z(n_72950739
		));
	notech_ao3 i_4374111(.A(n_59991), .B(in128[23]), .C(n_59648), .Z(n_72550735
		));
	notech_ao3 i_4474110(.A(n_59991), .B(in128[13]), .C(n_59648), .Z(n_72450734
		));
	notech_ao3 i_4774107(.A(n_59991), .B(in128[80]), .C(n_59648), .Z(n_72150731
		));
	notech_ao3 i_5174103(.A(n_59991), .B(in128[19]), .C(n_59648), .Z(n_71750727
		));
	notech_ao3 i_5374101(.A(n_59986), .B(in128[15]), .C(n_59648), .Z(n_71550725
		));
	notech_ao3 i_5574099(.A(n_59986), .B(in128[11]), .C(n_59648), .Z(n_71350723
		));
	notech_ao3 i_5874096(.A(n_59991), .B(in128[17]), .C(n_59647), .Z(n_71050720
		));
	notech_ao3 i_6474090(.A(n_59986), .B(in128[18]), .C(n_59647), .Z(n_70450714
		));
	notech_ao3 i_6674088(.A(n_59986), .B(in128[14]), .C(n_59647), .Z(n_70250712
		));
	notech_ao3 i_6874086(.A(n_59986), .B(in128[25]), .C(n_59647), .Z(n_70050710
		));
	notech_ao3 i_6974085(.A(n_59991), .B(in128[20]), .C(n_59647), .Z(n_69950709
		));
	notech_ao3 i_7374081(.A(n_59991), .B(in128[9]), .C(n_59647), .Z(n_69550705
		));
	notech_ao3 i_7474080(.A(n_59991), .B(in128[68]), .C(n_59648), .Z(n_69450704
		));
	notech_ao3 i_7574079(.A(n_59991), .B(in128[16]), .C(n_59648), .Z(n_69350703
		));
	notech_ao3 i_7674078(.A(n_59991), .B(in128[21]), .C(n_59648), .Z(n_69250702
		));
	notech_ao3 i_15074004(.A(n_59991), .B(in128[7]), .C(n_59647), .Z(n_61750629
		));
	notech_or4 i_65879(.A(fsm[2]), .B(fsm[1]), .C(fsm[0]), .D(n_2864), .Z(n_2884
		));
	notech_xor2 i_6334(.A(n_2872), .B(n_2879), .Z(n_2880));
	notech_xor2 i_214(.A(imm_sz[1]), .B(i_ptr[1]), .Z(n_2879));
	notech_xor2 i_6333(.A(n_2873), .B(n_2877), .Z(n_2878));
	notech_xor2 i_20(.A(imm_sz[2]), .B(i_ptr[2]), .Z(n_2877));
	notech_xor2 i_6332(.A(i_ptr[3]), .B(n_2874), .Z(n_2876));
	notech_nand2 i_6330(.A(i_ptr[3]), .B(n_40505), .Z(n_2875));
	notech_ao4 i_6331(.A(n_2197), .B(n_40506), .C(n_40593), .D(n_39368), .Z(n_2874
		));
	notech_ao4 i_2129836(.A(n_2872), .B(n_2194), .C(i_ptr[1]), .D(imm_sz[1])
		, .Z(n_2873));
	notech_and2 i_6329(.A(i_ptr[0]), .B(imm_sz[0]), .Z(n_2872));
	notech_nand2 i_496(.A(fsm[0]), .B(fsm[1]), .Z(n_2871));
	notech_or4 i_6339(.A(fsm[3]), .B(fsm[0]), .C(fsm[1]), .D(n_2867), .Z(n_2870
		));
	notech_nand2 i_494(.A(fsm[2]), .B(n_39377), .Z(n_2867));
	notech_or2 i_167(.A(fsm[2]), .B(n_2864), .Z(n_2865));
	notech_or2 i_464(.A(fsm[4]), .B(fsm[3]), .Z(n_2864));
	notech_and3 i_376(.A(n_40865), .B(n_40860), .C(n_40861), .Z(n_2860));
	notech_and4 i_373(.A(n_2183), .B(n_40871), .C(n_40870), .D(n_40869), .Z(n_2858
		));
	notech_and4 i_372(.A(n_40868), .B(n_40867), .C(n_40866), .D(n_40921), .Z
		(n_2855));
	notech_or4 i_65731(.A(n_2849), .B(n_2846), .C(n_2842), .D(n_2839), .Z(n_2851
		));
	notech_or2 i_3432(.A(n_40468), .B(pfx_sz[0]), .Z(n_172396417));
	notech_ao3 i_3434(.A(n_59980), .B(n_163096325), .C(n_2884), .Z(n_172496418
		));
	notech_ao3 i_3435(.A(n_59969), .B(n_163196326), .C(n_2884), .Z(n_172596419
		));
	notech_ao3 i_3437(.A(n_163296327), .B(n_59969), .C(n_2884), .Z(n_172696420
		));
	notech_ao3 i_3439(.A(n_59969), .B(in128[0]), .C(n_2884), .Z(n_172796421)
		);
	notech_ao3 i_3512(.A(opz[2]), .B(n_59969), .C(n_2884), .Z(n_172896422)
		);
	notech_nor2 i_3515(.A(n_5392), .B(int_excl[0]), .Z(n_172996423));
	notech_nor2 i_3516(.A(n_5392), .B(n_163396328), .Z(n_173096424));
	notech_ao3 i_3536(.A(n_39133), .B(n_2887), .C(n_2915), .Z(n_173196425)
		);
	notech_ao3 i_3763(.A(n_59969), .B(n_40938), .C(n_57101), .Z(n_173296426)
		);
	notech_and3 i_3783(.A(db67), .B(n_41563), .C(n_163496329), .Z(n_173396427
		));
	notech_ao3 i_3791(.A(n_59969), .B(in128[16]), .C(n_57101), .Z(n_173496428
		));
	notech_ao3 i_3792(.A(n_59969), .B(in128[17]), .C(n_57101), .Z(n_173596429
		));
	notech_ao3 i_3793(.A(n_59975), .B(in128[18]), .C(n_57101), .Z(n_173696430
		));
	notech_ao3 i_3794(.A(n_59975), .B(\to_acu2_0[0] ), .C(n_57101), .Z(n_173796431
		));
	notech_ao3 i_3797(.A(n_59969), .B(\to_acu2_0[2] ), .C(n_57101), .Z(n_173896432
		));
	notech_ao3 i_3798(.A(n_59969), .B(\to_acu2_0[3] ), .C(n_2884), .Z(n_173996433
		));
	notech_ao3 i_3799(.A(n_59969), .B(\to_acu2_0[4] ), .C(n_57101), .Z(n_174096434
		));
	notech_ao3 i_3800(.A(n_59969), .B(\to_acu2_0[7] ), .C(n_57101), .Z(n_174196435
		));
	notech_or4 i_361(.A(\to_acu2_0[79] ), .B(\to_acu2_0[47] ), .C(\to_acu2_0[45] 
		), .D(\to_acu2_0[46] ), .Z(n_2849));
	notech_or4 i_360(.A(\to_acu2_0[44] ), .B(\to_acu2_0[42] ), .C(\to_acu2_0[43] 
		), .D(\to_acu2_0[41] ), .Z(n_2846));
	notech_reg term_f_reg(.CP(n_62285), .D(n_61036), .CD(n_61737), .Q(term_f
		));
	notech_reg db67_reg(.CP(n_62285), .D(n_30898), .CD(n_61737), .Q(db67));
	notech_mux2 i_36606(.S(n_46391), .A(db67), .B(n_258094537), .Z(n_30898)
		);
	notech_reg_set fpu_indrm_reg_0(.CP(n_62285), .D(n_30904), .SD(1'b1), .Q(\fpu_indrm[0] 
		));
	notech_mux2 i_36614(.S(\nbus_13559[0] ), .A(\fpu_indrm[0] ), .B(n_173796431
		), .Z(n_30904));
	notech_reg_set fpu_indrm_reg_2(.CP(n_62285), .D(n_30910), .SD(1'b1), .Q(\fpu_indrm[2] 
		));
	notech_mux2 i_36622(.S(\nbus_13559[0] ), .A(\fpu_indrm[2] ), .B(n_173896432
		), .Z(n_30910));
	notech_reg_set fpu_indrm_reg_3(.CP(n_62285), .D(n_30916), .SD(1'b1), .Q(\fpu_indrm[3] 
		));
	notech_mux2 i_36630(.S(\nbus_13559[0] ), .A(\fpu_indrm[3] ), .B(n_173996433
		), .Z(n_30916));
	notech_or4 i_359(.A(\to_acu2_0[38] ), .B(\to_acu2_0[40] ), .C(\to_acu2_0[36] 
		), .D(\to_acu2_0[37] ), .Z(n_2842));
	notech_reg_set fpu_indrm_reg_4(.CP(n_62285), .D(n_30922), .SD(1'b1), .Q(\fpu_indrm[4] 
		));
	notech_mux2 i_36638(.S(\nbus_13559[0] ), .A(\fpu_indrm[4] ), .B(n_174096434
		), .Z(n_30922));
	notech_reg_set fpu_indrm_reg_7(.CP(n_62285), .D(n_30928), .SD(1'b1), .Q(\fpu_indrm[7] 
		));
	notech_mux2 i_36646(.S(\nbus_13559[0] ), .A(\fpu_indrm[7] ), .B(n_174196435
		), .Z(n_30928));
	notech_reg_set fpu_modrm_reg_0(.CP(n_62285), .D(n_30934), .SD(1'b1), .Q(\fpu_modrm[0] 
		));
	notech_mux2 i_36654(.S(\nbus_13559[0] ), .A(\fpu_modrm[0] ), .B(n_173496428
		), .Z(n_30934));
	notech_nand3 i_358(.A(n_40877), .B(n_40876), .C(n_2179), .Z(n_2839));
	notech_reg_set fpu_modrm_reg_1(.CP(n_62285), .D(n_30940), .SD(1'b1), .Q(\fpu_modrm[1] 
		));
	notech_mux2 i_36662(.S(\nbus_13559[0] ), .A(\fpu_modrm[1] ), .B(n_173596429
		), .Z(n_30940));
	notech_reg_set fpu_modrm_reg_2(.CP(n_62285), .D(n_30946), .SD(1'b1), .Q(\fpu_modrm[2] 
		));
	notech_mux2 i_36670(.S(\nbus_13559[0] ), .A(\fpu_modrm[2] ), .B(n_173696430
		), .Z(n_30946));
	notech_nao3 i_156(.A(n_2905), .B(n_2222), .C(fpu), .Z(n_2837));
	notech_reg displc_reg_0(.CP(n_62285), .D(n_30952), .CD(n_61737), .Q(displc
		[0]));
	notech_mux2 i_36678(.S(n_3176), .A(n_39173), .B(displc[0]), .Z(n_30952)
		);
	notech_ao4 i_226330(.A(n_58175), .B(n_40175), .C(n_59527), .D(n_40925), 
		.Z(n_2836));
	notech_reg displc_reg_1(.CP(n_62283), .D(n_30958), .CD(n_61737), .Q(displc
		[1]));
	notech_mux2 i_36686(.S(n_3176), .A(n_44046), .B(displc[1]), .Z(n_30958)
		);
	notech_reg displc_reg_2(.CP(n_62283), .D(n_30964), .CD(n_61737), .Q(displc
		[2]));
	notech_mux2 i_36694(.S(n_3176), .A(n_173396427), .B(displc[2]), .Z(n_30964
		));
	notech_ao4 i_326331(.A(n_58178), .B(n_40178), .C(n_59527), .D(n_40943), 
		.Z(n_2834));
	notech_reg sib_dec_reg(.CP(n_62283), .D(n_30970), .CD(n_61737), .Q(sib_dec
		));
	notech_mux2 i_36702(.S(n_3177), .A(n_41563), .B(sib_dec), .Z(n_30970));
	notech_reg mod_dec_reg(.CP(n_62283), .D(n_30976), .CD(n_61737), .Q(mod_dec
		));
	notech_mux2 i_36710(.S(n_3178), .A(n_173296426), .B(mod_dec), .Z(n_30976
		));
	notech_ao4 i_426332(.A(n_58178), .B(n_40180), .C(n_59527), .D(n_40941), 
		.Z(n_2832));
	notech_reg imm1_reg_0(.CP(n_62283), .D(n_30982), .CD(n_61737), .Q(\imm1[0] 
		));
	notech_mux2 i_36718(.S(n_58321), .A(\imm1[0] ), .B(n_39123), .Z(n_30982)
		);
	notech_reg imm1_reg_1(.CP(n_62285), .D(n_30988), .CD(n_61737), .Q(\imm1[1] 
		));
	notech_mux2 i_36726(.S(n_58321), .A(\imm1[1] ), .B(n_39124), .Z(n_30988)
		);
	notech_ao4 i_526333(.A(n_58178), .B(n_40183), .C(n_59527), .D(n_40940), 
		.Z(n_2830));
	notech_reg imm1_reg_2(.CP(n_62285), .D(n_30994), .CD(n_61737), .Q(\imm1[2] 
		));
	notech_mux2 i_36734(.S(n_58321), .A(\imm1[2] ), .B(n_39125), .Z(n_30994)
		);
	notech_reg imm1_reg_3(.CP(n_62283), .D(n_31000), .CD(n_61737), .Q(\imm1[3] 
		));
	notech_mux2 i_36742(.S(n_58315), .A(\imm1[3] ), .B(n_39126), .Z(n_31000)
		);
	notech_ao4 i_726335(.A(n_58178), .B(n_40187), .C(n_59527), .D(n_40924), 
		.Z(n_2828));
	notech_reg imm1_reg_4(.CP(n_62283), .D(n_31006), .CD(n_61735), .Q(\imm1[4] 
		));
	notech_mux2 i_36750(.S(n_58315), .A(\imm1[4] ), .B(n_39127), .Z(n_31006)
		);
	notech_reg imm1_reg_5(.CP(n_62283), .D(n_31012), .CD(n_61735), .Q(\imm1[5] 
		));
	notech_mux2 i_36758(.S(n_58315), .A(\imm1[5] ), .B(n_39129), .Z(n_31012)
		);
	notech_ao4 i_826336(.A(n_58178), .B(n_40189), .C(n_59524), .D(n_40944), 
		.Z(n_2826));
	notech_reg imm1_reg_6(.CP(n_62288), .D(n_31018), .CD(n_61735), .Q(\imm1[6] 
		));
	notech_mux2 i_36766(.S(n_58321), .A(\imm1[6] ), .B(n_39130), .Z(n_31018)
		);
	notech_reg imm1_reg_7(.CP(n_62288), .D(n_31024), .CD(n_61735), .Q(\imm1[7] 
		));
	notech_mux2 i_36774(.S(n_58321), .A(\imm1[7] ), .B(n_39132), .Z(n_31024)
		);
	notech_ao4 i_926337(.A(n_58178), .B(n_40191), .C(n_59524), .D(n_40923), 
		.Z(n_2824));
	notech_reg imm1_reg_8(.CP(n_62288), .D(n_31030), .CD(n_61735), .Q(\imm1[8] 
		));
	notech_mux2 i_36782(.S(n_58321), .A(\imm1[8] ), .B(n_39134), .Z(n_31030)
		);
	notech_reg imm1_reg_9(.CP(n_62288), .D(n_31036), .CD(n_61737), .Q(\imm1[9] 
		));
	notech_mux2 i_36790(.S(n_58321), .A(\imm1[9] ), .B(n_39136), .Z(n_31036)
		);
	notech_ao4 i_1126339(.A(n_58178), .B(n_40195), .C(n_59524), .D(n_40922),
		 .Z(n_2822));
	notech_reg imm1_reg_10(.CP(n_62288), .D(n_31042), .CD(n_61737), .Q(\imm1[10] 
		));
	notech_mux2 i_36798(.S(n_58321), .A(\imm1[10] ), .B(n_39137), .Z(n_31042
		));
	notech_reg imm1_reg_11(.CP(n_62288), .D(n_31048), .CD(n_61737), .Q(\imm1[11] 
		));
	notech_mux2 i_36806(.S(n_58321), .A(\imm1[11] ), .B(n_39138), .Z(n_31048
		));
	notech_ao4 i_5926387(.A(n_58178), .B(n_40269), .C(n_59524), .D(n_40921),
		 .Z(n_2820));
	notech_reg imm1_reg_12(.CP(n_62288), .D(n_31054), .CD(n_61735), .Q(\imm1[12] 
		));
	notech_mux2 i_36814(.S(n_58321), .A(\imm1[12] ), .B(n_39140), .Z(n_31054
		));
	notech_reg imm1_reg_13(.CP(n_62288), .D(n_31060), .CD(n_61737), .Q(\imm1[13] 
		));
	notech_mux2 i_36822(.S(n_58315), .A(\imm1[13] ), .B(n_39141), .Z(n_31060
		));
	notech_ao4 i_10826436(.A(n_58178), .B(n_40349), .C(n_59524), .D(n_40735)
		, .Z(n_2818));
	notech_reg imm1_reg_14(.CP(n_62288), .D(n_31066), .CD(n_61740), .Q(\imm1[14] 
		));
	notech_mux2 i_36830(.S(n_58315), .A(\imm1[14] ), .B(n_40058), .Z(n_31066
		));
	notech_reg imm1_reg_15(.CP(n_62288), .D(n_31072), .CD(n_61740), .Q(\imm1[15] 
		));
	notech_mux2 i_36838(.S(n_58315), .A(\imm1[15] ), .B(n_39142), .Z(n_31072
		));
	notech_ao4 i_11026438(.A(n_58178), .B(n_40352), .C(n_59527), .D(n_40737)
		, .Z(n_2816));
	notech_reg imm1_reg_16(.CP(n_62288), .D(n_31078), .CD(n_61740), .Q(\imm1[16] 
		));
	notech_mux2 i_36846(.S(n_58315), .A(\imm1[16] ), .B(n_40061), .Z(n_31078
		));
	notech_reg imm1_reg_17(.CP(n_62285), .D(n_31084), .CD(n_61740), .Q(\imm1[17] 
		));
	notech_mux2 i_36854(.S(n_58315), .A(\imm1[17] ), .B(n_39144), .Z(n_31084
		));
	notech_ao4 i_11126439(.A(n_58167), .B(n_40353), .C(n_59527), .D(n_40738)
		, .Z(n_2814));
	notech_reg imm1_reg_18(.CP(n_62285), .D(n_31090), .CD(n_61740), .Q(\imm1[18] 
		));
	notech_mux2 i_36862(.S(n_58315), .A(\imm1[18] ), .B(n_39145), .Z(n_31090
		));
	notech_reg imm1_reg_19(.CP(n_62285), .D(n_31096), .CD(n_61740), .Q(\imm1[19] 
		));
	notech_mux2 i_36870(.S(n_58315), .A(\imm1[19] ), .B(n_39146), .Z(n_31096
		));
	notech_ao4 i_11226440(.A(n_58155), .B(n_40354), .C(n_59527), .D(n_40739)
		, .Z(n_2812));
	notech_reg imm1_reg_20(.CP(n_62285), .D(n_31102), .CD(n_61740), .Q(\imm1[20] 
		));
	notech_mux2 i_36878(.S(n_58315), .A(\imm1[20] ), .B(n_39147), .Z(n_31102
		));
	notech_reg imm1_reg_21(.CP(n_62285), .D(n_31108), .CD(n_61740), .Q(\imm1[21] 
		));
	notech_mux2 i_36886(.S(n_58315), .A(\imm1[21] ), .B(n_39149), .Z(n_31108
		));
	notech_ao4 i_11326441(.A(n_58155), .B(n_40355), .C(n_59529), .D(n_40740)
		, .Z(n_2810));
	notech_reg imm1_reg_22(.CP(n_62288), .D(n_31114), .CD(n_61740), .Q(\imm1[22] 
		));
	notech_mux2 i_36894(.S(n_58315), .A(\imm1[22] ), .B(n_39150), .Z(n_31114
		));
	notech_reg imm1_reg_23(.CP(n_62288), .D(n_31120), .CD(n_61740), .Q(\imm1[23] 
		));
	notech_mux2 i_36902(.S(n_58315), .A(\imm1[23] ), .B(n_39151), .Z(n_31120
		));
	notech_ao4 i_11426442(.A(n_58155), .B(n_40356), .C(n_59527), .D(n_40741)
		, .Z(n_2808));
	notech_reg imm1_reg_24(.CP(n_62288), .D(n_31126), .CD(n_61740), .Q(\imm1[24] 
		));
	notech_mux2 i_36910(.S(n_58315), .A(\imm1[24] ), .B(n_39152), .Z(n_31126
		));
	notech_reg imm1_reg_25(.CP(n_62285), .D(n_31132), .CD(n_61737), .Q(\imm1[25] 
		));
	notech_mux2 i_36918(.S(n_58315), .A(\imm1[25] ), .B(n_40064), .Z(n_31132
		));
	notech_ao4 i_11526443(.A(n_58155), .B(n_40358), .C(n_59527), .D(n_40742)
		, .Z(n_2806));
	notech_reg imm1_reg_26(.CP(n_62285), .D(n_31138), .CD(n_61737), .Q(\imm1[26] 
		));
	notech_mux2 i_36926(.S(n_58321), .A(\imm1[26] ), .B(n_39153), .Z(n_31138
		));
	notech_reg imm1_reg_27(.CP(n_62283), .D(n_31144), .CD(n_61737), .Q(\imm1[27] 
		));
	notech_mux2 i_36934(.S(n_58326), .A(\imm1[27] ), .B(n_39154), .Z(n_31144
		));
	notech_ao4 i_11626444(.A(n_58155), .B(n_40360), .C(n_59527), .D(n_40743)
		, .Z(n_2804));
	notech_reg imm1_reg_28(.CP(n_62278), .D(n_31150), .CD(n_61737), .Q(\imm1[28] 
		));
	notech_mux2 i_36942(.S(n_58326), .A(\imm1[28] ), .B(n_39155), .Z(n_31150
		));
	notech_reg imm1_reg_29(.CP(n_62278), .D(n_31156), .CD(n_61737), .Q(\imm1[29] 
		));
	notech_mux2 i_36950(.S(n_58326), .A(\imm1[29] ), .B(n_39156), .Z(n_31156
		));
	notech_ao4 i_11726445(.A(n_58155), .B(n_40362), .C(n_59527), .D(n_40744)
		, .Z(n_2802));
	notech_reg imm1_reg_30(.CP(n_62278), .D(n_31162), .CD(n_61740), .Q(\imm1[30] 
		));
	notech_mux2 i_36958(.S(n_58326), .A(\imm1[30] ), .B(n_39157), .Z(n_31162
		));
	notech_reg imm1_reg_31(.CP(n_62278), .D(n_31168), .CD(n_61740), .Q(\imm1[31] 
		));
	notech_mux2 i_36966(.S(n_58326), .A(\imm1[31] ), .B(n_39158), .Z(n_31168
		));
	notech_ao4 i_11826446(.A(n_58155), .B(n_40364), .C(n_59527), .D(n_40745)
		, .Z(n_2800));
	notech_reg imm1_reg_32(.CP(n_62278), .D(n_31174), .CD(n_61740), .Q(\imm1[32] 
		));
	notech_mux2 i_36974(.S(n_58326), .A(\imm1[32] ), .B(n_39159), .Z(n_31174
		));
	notech_reg imm1_reg_33(.CP(n_62278), .D(n_31180), .CD(n_61740), .Q(\imm1[33] 
		));
	notech_mux2 i_36982(.S(n_58327), .A(\imm1[33] ), .B(n_39160), .Z(n_31180
		));
	notech_ao4 i_11926447(.A(n_58155), .B(n_40366), .C(n_59527), .D(n_40746)
		, .Z(n_2798));
	notech_reg imm1_reg_34(.CP(n_62278), .D(n_31186), .CD(n_61740), .Q(\imm1[34] 
		));
	notech_mux2 i_36990(.S(n_58327), .A(\imm1[34] ), .B(n_39161), .Z(n_31186
		));
	notech_reg imm1_reg_35(.CP(n_62278), .D(n_31192), .CD(n_61730), .Q(\imm1[35] 
		));
	notech_mux2 i_36998(.S(n_58327), .A(\imm1[35] ), .B(n_40067), .Z(n_31192
		));
	notech_ao4 i_12026448(.A(n_58155), .B(n_40367), .C(n_59524), .D(n_40747)
		, .Z(n_2796));
	notech_reg imm1_reg_36(.CP(n_62278), .D(n_31198), .CD(n_61730), .Q(\imm1[36] 
		));
	notech_mux2 i_37006(.S(n_58327), .A(\imm1[36] ), .B(n_39162), .Z(n_31198
		));
	notech_reg imm1_reg_37(.CP(n_62278), .D(n_31204), .CD(n_61730), .Q(\imm1[37] 
		));
	notech_mux2 i_37014(.S(n_58327), .A(\imm1[37] ), .B(n_39163), .Z(n_31204
		));
	notech_ao4 i_12126449(.A(n_58155), .B(n_40369), .C(n_59522), .D(n_40748)
		, .Z(n_2794));
	notech_reg imm1_reg_38(.CP(n_62276), .D(n_31210), .CD(n_61730), .Q(\imm1[38] 
		));
	notech_mux2 i_37022(.S(n_58327), .A(\imm1[38] ), .B(n_39164), .Z(n_31210
		));
	notech_reg imm1_reg_39(.CP(n_62276), .D(n_31216), .CD(n_61730), .Q(\imm1[39] 
		));
	notech_mux2 i_37030(.S(n_58327), .A(\imm1[39] ), .B(n_39165), .Z(n_31216
		));
	notech_ao4 i_12226450(.A(n_58157), .B(n_40370), .C(n_59522), .D(n_40749)
		, .Z(n_2792));
	notech_reg imm1_reg_40(.CP(n_62276), .D(n_31222), .CD(n_61730), .Q(\imm1[40] 
		));
	notech_mux2 i_37038(.S(n_58326), .A(\imm1[40] ), .B(n_39166), .Z(n_31222
		));
	notech_reg imm1_reg_41(.CP(n_62276), .D(n_31228), .CD(n_61730), .Q(\imm1[41] 
		));
	notech_mux2 i_37046(.S(n_58326), .A(\imm1[41] ), .B(n_40070), .Z(n_31228
		));
	notech_ao4 i_12526453(.A(n_58157), .B(n_40374), .C(n_59522), .D(n_40752)
		, .Z(n_2790));
	notech_reg imm1_reg_42(.CP(n_62276), .D(n_31234), .CD(n_61730), .Q(\imm1[42] 
		));
	notech_mux2 i_37054(.S(n_58326), .A(\imm1[42] ), .B(n_39167), .Z(n_31234
		));
	notech_reg imm1_reg_43(.CP(n_62276), .D(n_31240), .CD(n_61730), .Q(\imm1[43] 
		));
	notech_mux2 i_37062(.S(n_58321), .A(\imm1[43] ), .B(n_39168), .Z(n_31240
		));
	notech_ao4 i_13126459(.A(n_58157), .B(n_40380), .C(n_59522), .D(n_40758)
		, .Z(n_2788));
	notech_reg imm1_reg_44(.CP(n_62276), .D(n_31246), .CD(n_61730), .Q(\imm1[44] 
		));
	notech_mux2 i_37070(.S(n_58326), .A(\imm1[44] ), .B(n_39169), .Z(n_31246
		));
	notech_reg imm1_reg_45(.CP(n_62276), .D(n_31252), .CD(n_61730), .Q(\imm1[45] 
		));
	notech_mux2 i_37078(.S(n_58326), .A(\imm1[45] ), .B(n_40073), .Z(n_31252
		));
	notech_ao4 i_13226460(.A(n_58157), .B(n_40381), .C(n_59522), .D(n_40759)
		, .Z(n_2786));
	notech_reg imm1_reg_46(.CP(n_62276), .D(n_31258), .CD(n_61728), .Q(\imm1[46] 
		));
	notech_mux2 i_37086(.S(n_58326), .A(\imm1[46] ), .B(n_39170), .Z(n_31258
		));
	notech_reg imm1_reg_47(.CP(n_62276), .D(n_31264), .CD(n_61728), .Q(\imm1[47] 
		));
	notech_mux2 i_37094(.S(n_58326), .A(\imm1[47] ), .B(n_39171), .Z(n_31264
		));
	notech_ao4 i_13326461(.A(n_58157), .B(n_40382), .C(n_59522), .D(n_40760)
		, .Z(n_2784));
	notech_reg imm2_reg_0(.CP(n_62276), .D(n_31270), .CD(n_61728), .Q(\imm2[0] 
		));
	notech_mux2 i_37102(.S(n_55095), .A(\imm2[0] ), .B(n_44449), .Z(n_31270)
		);
	notech_reg imm2_reg_1(.CP(n_62283), .D(n_31276), .CD(n_61728), .Q(\imm2[1] 
		));
	notech_mux2 i_37110(.S(n_55095), .A(\imm2[1] ), .B(n_44455), .Z(n_31276)
		);
	notech_ao4 i_13426462(.A(n_58155), .B(n_40383), .C(n_59522), .D(n_40761)
		, .Z(n_2782));
	notech_reg imm2_reg_2(.CP(n_62283), .D(n_31282), .CD(n_61728), .Q(\imm2[2] 
		));
	notech_mux2 i_37118(.S(n_55095), .A(\imm2[2] ), .B(n_44461), .Z(n_31282)
		);
	notech_reg imm2_reg_3(.CP(n_62283), .D(n_31288), .CD(n_61730), .Q(\imm2[3] 
		));
	notech_mux2 i_37126(.S(n_55089), .A(\imm2[3] ), .B(n_44467), .Z(n_31288)
		);
	notech_ao4 i_13526463(.A(n_58155), .B(n_40384), .C(n_59522), .D(n_40762)
		, .Z(n_2780));
	notech_reg imm2_reg_4(.CP(n_62283), .D(n_31294), .CD(n_61730), .Q(\imm2[4] 
		));
	notech_mux2 i_37134(.S(n_55089), .A(\imm2[4] ), .B(n_44473), .Z(n_31294)
		);
	notech_reg imm2_reg_5(.CP(n_62283), .D(n_31300), .CD(n_61728), .Q(\imm2[5] 
		));
	notech_mux2 i_37142(.S(n_55089), .A(\imm2[5] ), .B(n_44479), .Z(n_31300)
		);
	notech_ao4 i_13626464(.A(n_58155), .B(n_40385), .C(n_59522), .D(n_40763)
		, .Z(n_2778));
	notech_reg imm2_reg_6(.CP(n_62283), .D(n_31306), .CD(n_61728), .Q(\imm2[6] 
		));
	notech_mux2 i_37150(.S(n_55095), .A(\imm2[6] ), .B(n_44485), .Z(n_31306)
		);
	notech_reg imm2_reg_7(.CP(n_62283), .D(n_31312), .CD(n_61728), .Q(\imm2[7] 
		));
	notech_mux2 i_37158(.S(n_55095), .A(\imm2[7] ), .B(n_44491), .Z(n_31312)
		);
	notech_ao4 i_13726465(.A(n_58157), .B(n_40386), .C(n_59522), .D(n_40764)
		, .Z(n_2776));
	notech_reg imm2_reg_8(.CP(n_62283), .D(n_31318), .CD(n_61735), .Q(\imm2[8] 
		));
	notech_mux2 i_37166(.S(n_55095), .A(\imm2[8] ), .B(n_44497), .Z(n_31318)
		);
	notech_reg imm2_reg_9(.CP(n_62283), .D(n_31324), .CD(n_61735), .Q(\imm2[9] 
		));
	notech_mux2 i_37174(.S(n_55095), .A(\imm2[9] ), .B(n_44503), .Z(n_31324)
		);
	notech_ao4 i_13826466(.A(n_58157), .B(n_40387), .C(n_59524), .D(n_40765)
		, .Z(n_2774));
	notech_reg imm2_reg_10(.CP(n_62283), .D(n_31330), .CD(n_61735), .Q(\imm2[10] 
		));
	notech_mux2 i_37182(.S(n_55095), .A(\imm2[10] ), .B(n_44509), .Z(n_31330
		));
	notech_reg imm2_reg_11(.CP(n_62283), .D(n_31336), .CD(n_61735), .Q(\imm2[11] 
		));
	notech_mux2 i_37190(.S(n_55095), .A(\imm2[11] ), .B(n_44515), .Z(n_31336
		));
	notech_ao4 i_13926467(.A(n_58155), .B(n_40388), .C(n_59524), .D(n_40766)
		, .Z(n_2772));
	notech_reg imm2_reg_12(.CP(n_62278), .D(n_31342), .CD(n_61735), .Q(\imm2[12] 
		));
	notech_mux2 i_37198(.S(n_55095), .A(\imm2[12] ), .B(n_44521), .Z(n_31342
		));
	notech_reg imm2_reg_13(.CP(n_62278), .D(n_31348), .CD(n_61735), .Q(\imm2[13] 
		));
	notech_mux2 i_37206(.S(n_55089), .A(\imm2[13] ), .B(n_44527), .Z(n_31348
		));
	notech_ao4 i_14026468(.A(n_58152), .B(n_40389), .C(n_59524), .D(n_40767)
		, .Z(n_2770));
	notech_reg imm2_reg_14(.CP(n_62278), .D(n_31354), .CD(n_61735), .Q(\imm2[14] 
		));
	notech_mux2 i_37214(.S(n_55089), .A(\imm2[14] ), .B(n_44533), .Z(n_31354
		));
	notech_reg imm2_reg_15(.CP(n_62278), .D(n_31360), .CD(n_61735), .Q(\imm2[15] 
		));
	notech_mux2 i_37222(.S(n_55089), .A(\imm2[15] ), .B(n_44539), .Z(n_31360
		));
	notech_ao4 i_14226470(.A(n_58150), .B(n_40391), .C(n_59524), .D(n_40769)
		, .Z(n_2768));
	notech_reg imm2_reg_16(.CP(n_62278), .D(n_31366), .CD(n_61735), .Q(\imm2[16] 
		));
	notech_mux2 i_37230(.S(n_55089), .A(\imm2[16] ), .B(n_3277), .Z(n_31366)
		);
	notech_reg imm2_reg_17(.CP(n_62278), .D(n_31372), .CD(n_61735), .Q(\imm2[17] 
		));
	notech_mux2 i_37238(.S(n_55089), .A(\imm2[17] ), .B(n_44551), .Z(n_31372
		));
	notech_ao4 i_14626474(.A(n_58152), .B(n_40395), .C(n_59524), .D(n_40773)
		, .Z(n_2766));
	notech_reg imm2_reg_18(.CP(n_62278), .D(n_31378), .CD(n_61735), .Q(\imm2[18] 
		));
	notech_mux2 i_37246(.S(n_55089), .A(\imm2[18] ), .B(n_44557), .Z(n_31378
		));
	notech_reg imm2_reg_19(.CP(n_62278), .D(n_31384), .CD(n_61730), .Q(\imm2[19] 
		));
	notech_mux2 i_37254(.S(n_55089), .A(\imm2[19] ), .B(n_44563), .Z(n_31384
		));
	notech_ao4 i_14726475(.A(n_58152), .B(n_40396), .C(n_59522), .D(n_40774)
		, .Z(n_2764));
	notech_reg imm2_reg_20(.CP(n_62278), .D(n_31390), .CD(n_61730), .Q(\imm2[20] 
		));
	notech_mux2 i_37262(.S(n_55089), .A(\imm2[20] ), .B(n_44569), .Z(n_31390
		));
	notech_reg imm2_reg_21(.CP(n_62278), .D(n_31396), .CD(n_61730), .Q(\imm2[21] 
		));
	notech_mux2 i_37270(.S(n_55089), .A(\imm2[21] ), .B(n_44575), .Z(n_31396
		));
	notech_ao4 i_14826476(.A(n_58152), .B(n_40397), .C(n_59522), .D(n_40775)
		, .Z(n_2762));
	notech_reg imm2_reg_22(.CP(n_62295), .D(n_31402), .CD(n_61730), .Q(\imm2[22] 
		));
	notech_mux2 i_37278(.S(n_55089), .A(\imm2[22] ), .B(n_44581), .Z(n_31402
		));
	notech_reg imm2_reg_23(.CP(n_62295), .D(n_31408), .CD(n_61730), .Q(\imm2[23] 
		));
	notech_mux2 i_37286(.S(n_55089), .A(\imm2[23] ), .B(n_44587), .Z(n_31408
		));
	notech_ao4 i_15126479(.A(n_58150), .B(n_40401), .C(n_59524), .D(n_40778)
		, .Z(n_2760));
	notech_reg imm2_reg_24(.CP(n_62295), .D(n_31414), .CD(n_61735), .Q(\imm2[24] 
		));
	notech_mux2 i_37294(.S(n_55089), .A(\imm2[24] ), .B(n_44593), .Z(n_31414
		));
	notech_reg imm2_reg_25(.CP(n_62295), .D(n_31420), .CD(n_61735), .Q(\imm2[25] 
		));
	notech_mux2 i_37302(.S(n_55089), .A(\imm2[25] ), .B(n_44599), .Z(n_31420
		));
	notech_ao4 i_15326481(.A(n_58150), .B(n_40405), .C(n_59524), .D(n_40780)
		, .Z(n_2758));
	notech_reg imm2_reg_26(.CP(n_62295), .D(n_31426), .CD(n_61735), .Q(\imm2[26] 
		));
	notech_mux2 i_37310(.S(n_55095), .A(\imm2[26] ), .B(n_44605), .Z(n_31426
		));
	notech_reg imm2_reg_27(.CP(n_62295), .D(n_31432), .CD(n_61730), .Q(\imm2[27] 
		));
	notech_mux2 i_37318(.S(n_55100), .A(\imm2[27] ), .B(n_44611), .Z(n_31432
		));
	notech_ao4 i_15426482(.A(n_58150), .B(n_40406), .C(n_59524), .D(n_40781)
		, .Z(n_2756));
	notech_reg imm2_reg_28(.CP(n_62295), .D(n_31438), .CD(n_61730), .Q(\imm2[28] 
		));
	notech_mux2 i_37326(.S(n_55100), .A(\imm2[28] ), .B(n_44617), .Z(n_31438
		));
	notech_reg imm2_reg_29(.CP(n_62295), .D(n_31444), .CD(n_61740), .Q(\imm2[29] 
		));
	notech_mux2 i_37334(.S(n_55100), .A(\imm2[29] ), .B(n_44623), .Z(n_31444
		));
	notech_ao4 i_16326491(.A(n_58150), .B(n_40416), .C(n_59529), .D(n_40790)
		, .Z(n_2754));
	notech_reg imm2_reg_30(.CP(n_62295), .D(n_31450), .CD(n_61747), .Q(\imm2[30] 
		));
	notech_mux2 i_37342(.S(n_55100), .A(\imm2[30] ), .B(n_44629), .Z(n_31450
		));
	notech_reg imm2_reg_31(.CP(n_62295), .D(n_31456), .CD(n_61747), .Q(\imm2[31] 
		));
	notech_mux2 i_37350(.S(n_55100), .A(\imm2[31] ), .B(n_44635), .Z(n_31456
		));
	notech_ao4 i_17326501(.A(n_58150), .B(n_40428), .C(n_59536), .D(n_40800)
		, .Z(n_2752));
	notech_reg imm2_reg_32(.CP(n_62295), .D(n_31462), .CD(n_61747), .Q(\imm2[32] 
		));
	notech_mux2 i_37358(.S(n_55100), .A(\imm2[32] ), .B(n_44641), .Z(n_31462
		));
	notech_reg imm2_reg_33(.CP(n_62295), .D(n_31468), .CD(n_61747), .Q(\imm2[33] 
		));
	notech_mux2 i_37366(.S(n_55101), .A(\imm2[33] ), .B(n_44647), .Z(n_31468
		));
	notech_ao4 i_17726505(.A(n_58152), .B(n_40432), .C(n_59536), .D(n_40804)
		, .Z(n_275094707));
	notech_reg imm2_reg_34(.CP(n_62295), .D(n_31474), .CD(n_61747), .Q(\imm2[34] 
		));
	notech_mux2 i_37374(.S(n_55101), .A(\imm2[34] ), .B(n_44653), .Z(n_31474
		));
	notech_reg imm2_reg_35(.CP(n_62293), .D(n_31480), .CD(n_61747), .Q(\imm2[35] 
		));
	notech_mux2 i_37382(.S(n_55101), .A(\imm2[35] ), .B(n_44659), .Z(n_31480
		));
	notech_ao4 i_19626524(.A(n_59536), .B(n_40823), .C(n_58152), .D(n_40452)
		, .Z(n_274894705));
	notech_reg imm2_reg_36(.CP(n_62293), .D(n_31486), .CD(n_61747), .Q(\imm2[36] 
		));
	notech_mux2 i_37390(.S(n_55101), .A(\imm2[36] ), .B(n_44665), .Z(n_31486
		));
	notech_reg imm2_reg_37(.CP(n_62293), .D(n_31492), .CD(n_61747), .Q(\imm2[37] 
		));
	notech_mux2 i_37398(.S(n_55101), .A(\imm2[37] ), .B(n_44671), .Z(n_31492
		));
	notech_ao4 i_323153(.A(n_58152), .B(n_39420), .C(n_39381), .D(n_39576), 
		.Z(n_274694703));
	notech_reg imm2_reg_38(.CP(n_62295), .D(n_31498), .CD(n_61747), .Q(\imm2[38] 
		));
	notech_mux2 i_37406(.S(n_55101), .A(\imm2[38] ), .B(n_44677), .Z(n_31498
		));
	notech_reg imm2_reg_39(.CP(n_62295), .D(n_31504), .CD(n_61747), .Q(\imm2[39] 
		));
	notech_mux2 i_37414(.S(n_55101), .A(\imm2[39] ), .B(n_44683), .Z(n_31504
		));
	notech_nand3 i_7325723(.A(n_60059), .B(n_274394700), .C(n_274194698), .Z
		(n_274494701));
	notech_reg imm2_reg_40(.CP(n_62295), .D(n_31510), .CD(n_61747), .Q(\imm2[40] 
		));
	notech_mux2 i_37422(.S(n_55100), .A(\imm2[40] ), .B(n_44689), .Z(n_31510
		));
	notech_nand3 i_1391(.A(inst_deco1[72]), .B(n_59017), .C(n_2885), .Z(n_274394700
		));
	notech_reg imm2_reg_41(.CP(n_62295), .D(n_31516), .CD(n_61747), .Q(\imm2[41] 
		));
	notech_mux2 i_37430(.S(n_55100), .A(\imm2[41] ), .B(n_44695), .Z(n_31516
		));
	notech_nand2 i_10(.A(n_40937), .B(pc_req), .Z(n_274294699));
	notech_reg imm2_reg_42(.CP(n_62295), .D(n_31522), .CD(n_61747), .Q(\imm2[42] 
		));
	notech_mux2 i_37438(.S(n_55100), .A(\imm2[42] ), .B(n_44701), .Z(n_31522
		));
	notech_or4 i_1390(.A(n_59647), .B(pc_req), .C(pg_fault), .D(n_40667), .Z
		(n_274194698));
	notech_reg imm2_reg_43(.CP(n_62299), .D(n_31528), .CD(n_61747), .Q(\imm2[43] 
		));
	notech_mux2 i_37446(.S(n_55095), .A(\imm2[43] ), .B(n_2019), .Z(n_31528)
		);
	notech_nand3 i_9225742(.A(n_60059), .B(n_273994696), .C(n_273894695), .Z
		(n_274094697));
	notech_reg imm2_reg_44(.CP(n_62299), .D(n_31534), .CD(n_61745), .Q(\imm2[44] 
		));
	notech_mux2 i_37454(.S(n_55100), .A(\imm2[44] ), .B(n_44713), .Z(n_31534
		));
	notech_nand3 i_1385(.A(n_2885), .B(inst_deco1[91]), .C(n_59017), .Z(n_273994696
		));
	notech_reg imm2_reg_45(.CP(n_62299), .D(n_31540), .CD(n_61747), .Q(\imm2[45] 
		));
	notech_mux2 i_37462(.S(n_55100), .A(\imm2[45] ), .B(n_3278), .Z(n_31540)
		);
	notech_or4 i_1384(.A(n_59653), .B(pc_req), .C(pg_fault), .D(n_40686), .Z
		(n_273894695));
	notech_reg imm2_reg_46(.CP(n_62299), .D(n_31546), .CD(n_61747), .Q(\imm2[46] 
		));
	notech_mux2 i_37470(.S(n_55100), .A(\imm2[46] ), .B(n_44725), .Z(n_31546
		));
	notech_nand3 i_323150(.A(n_273294689), .B(n_59968), .C(n_273694693), .Z(n_273794694
		));
	notech_reg imm2_reg_47(.CP(n_62299), .D(n_31552), .CD(n_61747), .Q(\imm2[47] 
		));
	notech_mux2 i_37478(.S(n_55100), .A(\imm2[47] ), .B(n_44731), .Z(n_31552
		));
	notech_nand3 i_1382(.A(n_60042), .B(opz1[2]), .C(n_59968), .Z(n_273694693
		));
	notech_reg trig_it_reg(.CP(n_62299), .D(n_31558), .CD(n_61747), .Q(trig_it
		));
	notech_mux2 i_37486(.S(n_44084), .A(trig_it), .B(n_173196425), .Z(n_31558
		));
	notech_nand3 i_323147(.A(n_273294689), .B(n_59969), .C(n_273494691), .Z(n_273594692
		));
	notech_reg trig_itf_reg(.CP(n_62299), .D(trig_it), .CD(n_61747), .Q(trig_itf
		));
	notech_reg intf_reg(.CP(n_62299), .D(int_main), .CD(n_61747), .Q(intf)
		);
	notech_reg_set intff_reg(.CP(n_62299), .D(n_31568), .SD(1'b1), .Q(intff)
		);
	notech_mux2 i_37502(.S(n_61751), .A(intff), .B(intf), .Z(n_31568));
	notech_nand3 i_1380(.A(n_60042), .B(opz2[2]), .C(n_59968), .Z(n_273494691
		));
	notech_reg ififo_rvect4_reg_0(.CP(n_62299), .D(n_31574), .CD(n_61751), .Q
		(ififo_rvect4[0]));
	notech_mux2 i_37510(.S(\nbus_13535[0] ), .A(ififo_rvect4[0]), .B(n_161696311
		), .Z(n_31574));
	notech_nand2 i_203(.A(n_273294689), .B(n_59968), .Z(n_273394690));
	notech_reg ififo_rvect4_reg_1(.CP(n_62299), .D(n_31580), .CD(n_61751), .Q
		(ififo_rvect4[1]));
	notech_mux2 i_37518(.S(\nbus_13535[0] ), .A(ififo_rvect4[1]), .B(n_161796312
		), .Z(n_31580));
	notech_nao3 i_1378(.A(opz[2]), .B(n_59968), .C(n_59657), .Z(n_273294689)
		);
	notech_reg ififo_rvect4_reg_2(.CP(n_62299), .D(n_31586), .CD(n_61751), .Q
		(ififo_rvect4[2]));
	notech_mux2 i_37526(.S(\nbus_13535[0] ), .A(ififo_rvect4[2]), .B(n_161896313
		), .Z(n_31586));
	notech_ao4 i_3527834(.A(n_58152), .B(n_39220), .C(n_54557), .D(n_40279),
		 .Z(n_273194688));
	notech_reg ififo_rvect4_reg_3(.CP(n_62299), .D(n_31592), .CD(n_61751), .Q
		(ififo_rvect4[3]));
	notech_mux2 i_37534(.S(\nbus_13535[0] ), .A(ififo_rvect4[3]), .B(n_161996314
		), .Z(n_31592));
	notech_reg ififo_rvect4_reg_4(.CP(n_62299), .D(n_31598), .CD(n_61753), .Q
		(ififo_rvect4[4]));
	notech_mux2 i_37542(.S(\nbus_13535[0] ), .A(ififo_rvect4[4]), .B(n_162096315
		), .Z(n_31598));
	notech_ao4 i_4527844(.A(n_58152), .B(n_39240), .C(n_2948), .D(n_40281), 
		.Z(n_272994686));
	notech_reg ififo_rvect4_reg_5(.CP(n_62295), .D(n_31604), .CD(n_61753), .Q
		(ififo_rvect4[5]));
	notech_mux2 i_37550(.S(\nbus_13535[0] ), .A(ififo_rvect4[5]), .B(n_162196316
		), .Z(n_31604));
	notech_reg ififo_rvect4_reg_6(.CP(n_62295), .D(n_31610), .CD(n_61751), .Q
		(ififo_rvect4[6]));
	notech_mux2 i_37558(.S(\nbus_13535[0] ), .A(ififo_rvect4[6]), .B(n_162296317
		), .Z(n_31610));
	notech_ao4 i_627223(.A(n_58152), .B(n_40472), .C(n_59536), .D(n_40469), 
		.Z(n_272794684));
	notech_reg ififo_rvect4_reg_7(.CP(n_62299), .D(n_31616), .CD(n_61751), .Q
		(ififo_rvect4[7]));
	notech_mux2 i_37566(.S(\nbus_13535[0] ), .A(ififo_rvect4[7]), .B(n_162396318
		), .Z(n_31616));
	notech_reg ififo_rvect3_reg_0(.CP(n_62299), .D(n_31622), .CD(n_61751), .Q
		(ififo_rvect3[0]));
	notech_mux2 i_37574(.S(\nbus_13535[0] ), .A(ififo_rvect3[0]), .B(n_43963
		), .Z(n_31622));
	notech_ao4 i_18126298(.A(n_59536), .B(n_40808), .C(n_58152), .D(n_40126)
		, .Z(n_272594682));
	notech_reg ififo_rvect3_reg_1(.CP(n_62299), .D(n_31628), .CD(n_61751), .Q
		(ififo_rvect3[1]));
	notech_mux2 i_37582(.S(\nbus_13535[0] ), .A(ififo_rvect3[1]), .B(n_43969
		), .Z(n_31628));
	notech_reg ififo_rvect3_reg_2(.CP(n_62299), .D(n_31634), .CD(n_61751), .Q
		(ififo_rvect3[2]));
	notech_mux2 i_37590(.S(\nbus_13535[0] ), .A(ififo_rvect3[2]), .B(n_43975
		), .Z(n_31634));
	notech_ao4 i_12825522(.A(n_58152), .B(n_39613), .C(n_59534), .D(n_40722)
		, .Z(n_272394680));
	notech_reg ififo_rvect3_reg_3(.CP(n_62299), .D(n_31640), .CD(n_61751), .Q
		(ififo_rvect3[3]));
	notech_mux2 i_37598(.S(\nbus_13535[0] ), .A(ififo_rvect3[3]), .B(n_43981
		), .Z(n_31640));
	notech_reg ififo_rvect3_reg_4(.CP(n_62293), .D(n_31646), .CD(n_61751), .Q
		(ififo_rvect3[4]));
	notech_mux2 i_37606(.S(\nbus_13535[0] ), .A(ififo_rvect3[4]), .B(n_43987
		), .Z(n_31646));
	notech_ao4 i_123142(.A(n_58152), .B(n_39410), .C(n_40918), .D(n_39987), 
		.Z(n_272194678));
	notech_reg ififo_rvect3_reg_5(.CP(n_62290), .D(n_31652), .CD(n_61751), .Q
		(ififo_rvect3[5]));
	notech_mux2 i_37614(.S(\nbus_13535[0] ), .A(ififo_rvect3[5]), .B(n_43993
		), .Z(n_31652));
	notech_reg ififo_rvect3_reg_6(.CP(n_62290), .D(n_31658), .CD(n_61751), .Q
		(ififo_rvect3[6]));
	notech_mux2 i_37622(.S(\nbus_13535[0] ), .A(ififo_rvect3[6]), .B(n_43999
		), .Z(n_31658));
	notech_ao4 i_123109(.A(n_40468), .B(n_3173), .C(n_271194668), .D(n_40501
		), .Z(n_271994676));
	notech_reg ififo_rvect3_reg_7(.CP(n_62290), .D(n_31664), .CD(n_61751), .Q
		(ififo_rvect3[7]));
	notech_mux2 i_37630(.S(\nbus_13535[0] ), .A(ififo_rvect3[7]), .B(n_44005
		), .Z(n_31664));
	notech_reg ififo_rvect2_reg_0(.CP(n_62290), .D(n_31670), .CD(n_61751), .Q
		(ififo_rvect2[0]));
	notech_mux2 i_37638(.S(n_55744), .A(ififo_rvect2[0]), .B(n_42871), .Z(n_31670
		));
	notech_ao4 i_223110(.A(n_40468), .B(n_271694673), .C(n_271194668), .D(n_40501
		), .Z(n_271794674));
	notech_reg ififo_rvect2_reg_1(.CP(n_62290), .D(n_31676), .CD(n_61751), .Q
		(ififo_rvect2[1]));
	notech_mux2 i_37646(.S(n_55744), .A(ififo_rvect2[1]), .B(n_42877), .Z(n_31676
		));
	notech_nor2 i_275(.A(ipg_fault), .B(n_271494671), .Z(n_271694673));
	notech_reg ififo_rvect2_reg_2(.CP(n_62290), .D(n_31682), .CD(n_61751), .Q
		(ififo_rvect2[2]));
	notech_mux2 i_37654(.S(n_55744), .A(ififo_rvect2[2]), .B(n_42883), .Z(n_31682
		));
	notech_reg ififo_rvect2_reg_3(.CP(n_62290), .D(n_31688), .CD(n_61751), .Q
		(ififo_rvect2[3]));
	notech_mux2 i_37662(.S(n_55744), .A(ififo_rvect2[3]), .B(n_42889), .Z(n_31688
		));
	notech_and2 i_1336(.A(n_1507), .B(n_2905), .Z(n_271494671));
	notech_reg ififo_rvect2_reg_4(.CP(n_62290), .D(n_31694), .CD(n_61742), .Q
		(ififo_rvect2[4]));
	notech_mux2 i_37670(.S(n_55744), .A(ififo_rvect2[4]), .B(n_42895), .Z(n_31694
		));
	notech_reg ififo_rvect2_reg_5(.CP(n_62290), .D(n_31700), .CD(n_61742), .Q
		(ififo_rvect2[5]));
	notech_mux2 i_37678(.S(n_55744), .A(ififo_rvect2[5]), .B(n_42901), .Z(n_31700
		));
	notech_reg ififo_rvect2_reg_6(.CP(n_62290), .D(n_31706), .CD(n_61742), .Q
		(ififo_rvect2[6]));
	notech_mux2 i_37686(.S(n_55744), .A(ififo_rvect2[6]), .B(n_42907), .Z(n_31706
		));
	notech_and2 i_1334(.A(n_59534), .B(n_3172), .Z(n_271194668));
	notech_reg ififo_rvect2_reg_7(.CP(n_62290), .D(n_31712), .CD(n_61742), .Q
		(ififo_rvect2[7]));
	notech_mux2 i_37694(.S(n_55744), .A(ififo_rvect2[7]), .B(n_42913), .Z(n_31712
		));
	notech_ao4 i_323111(.A(n_270994666), .B(n_2219), .C(n_227296437), .D(n_2915
		), .Z(n_271094667));
	notech_reg ififo_rvect1_reg_0(.CP(n_62288), .D(n_31718), .CD(n_61742), .Q
		(ififo_rvect1[0]));
	notech_mux2 i_37702(.S(n_55744), .A(ififo_rvect1[0]), .B(n_44367), .Z(n_31718
		));
	notech_ao4 i_272(.A(n_59534), .B(n_2887), .C(n_40468), .D(n_2888), .Z(n_270994666
		));
	notech_reg ififo_rvect1_reg_1(.CP(n_62288), .D(n_31724), .CD(n_61742), .Q
		(ififo_rvect1[1]));
	notech_mux2 i_37710(.S(n_55744), .A(ififo_rvect1[1]), .B(n_44373), .Z(n_31724
		));
	notech_reg ififo_rvect1_reg_2(.CP(n_62288), .D(n_31730), .CD(n_61742), .Q
		(ififo_rvect1[2]));
	notech_mux2 i_37718(.S(n_55744), .A(ififo_rvect1[2]), .B(n_44379), .Z(n_31730
		));
	notech_reg ififo_rvect1_reg_3(.CP(n_62288), .D(n_31736), .CD(n_61742), .Q
		(ififo_rvect1[3]));
	notech_mux2 i_37726(.S(n_55744), .A(ififo_rvect1[3]), .B(n_44385), .Z(n_31736
		));
	notech_reg ififo_rvect1_reg_4(.CP(n_62288), .D(n_31742), .CD(n_61742), .Q
		(ififo_rvect1[4]));
	notech_mux2 i_37734(.S(n_55744), .A(ififo_rvect1[4]), .B(n_44391), .Z(n_31742
		));
	notech_reg ififo_rvect1_reg_5(.CP(n_62290), .D(n_31748), .CD(n_61742), .Q
		(ififo_rvect1[5]));
	notech_mux2 i_37742(.S(n_55744), .A(ififo_rvect1[5]), .B(n_44397), .Z(n_31748
		));
	notech_and4 i_123226(.A(n_3162), .B(n_270294659), .C(n_3168), .D(n_270394660
		), .Z(n_270494661));
	notech_reg ififo_rvect1_reg_6(.CP(n_62290), .D(n_31754), .CD(n_61742), .Q
		(ififo_rvect1[6]));
	notech_mux2 i_37750(.S(n_55744), .A(ififo_rvect1[6]), .B(n_44403), .Z(n_31754
		));
	notech_or2 i_1314(.A(n_270094657), .B(n_40938), .Z(n_270394660));
	notech_reg ififo_rvect1_reg_7(.CP(n_62290), .D(n_31760), .CD(n_61742), .Q
		(ififo_rvect1[7]));
	notech_mux2 i_37758(.S(n_55744), .A(ififo_rvect1[7]), .B(n_44409), .Z(n_31760
		));
	notech_or4 i_1315(.A(n_3158), .B(\to_acu2_0[2] ), .C(\to_acu2_0[3] ), .D
		(n_40940), .Z(n_270294659));
	notech_reg int_excl_reg_0(.CP(n_62288), .D(n_31766), .CD(n_61742), .Q(int_excl
		[0]));
	notech_mux2 i_37766(.S(\nbus_13565[0] ), .A(int_excl[0]), .B(n_172996423
		), .Z(n_31766));
	notech_reg int_excl_reg_1(.CP(n_62290), .D(n_31772), .CD(n_61740), .Q(int_excl
		[1]));
	notech_mux2 i_37774(.S(\nbus_13565[0] ), .A(int_excl[1]), .B(n_173096424
		), .Z(n_31772));
	notech_ao4 i_268(.A(n_3139), .B(n_3170), .C(n_269794654), .D(n_3135), .Z
		(n_270094657));
	notech_reg int_excl_reg_2(.CP(n_62293), .D(n_31778), .CD(n_61740), .Q(int_excl
		[2]));
	notech_mux2 i_37782(.S(\nbus_13565[0] ), .A(int_excl[2]), .B(n_268294639
		), .Z(n_31778));
	notech_nor2 i_269(.A(n_2910), .B(n_269594652), .Z(n_269994656));
	notech_reg int_excl_reg_3(.CP(n_62293), .D(n_31784), .CD(n_61740), .Q(int_excl
		[3]));
	notech_mux2 i_37790(.S(\nbus_13565[0] ), .A(int_excl[3]), .B(n_161296307
		), .Z(n_31784));
	notech_reg int_excl_reg_4(.CP(n_62293), .D(n_31790), .CD(n_61742), .Q(int_excl
		[4]));
	notech_mux2 i_37798(.S(\nbus_13565[0] ), .A(int_excl[4]), .B(n_49899), .Z
		(n_31790));
	notech_and2 i_270(.A(n_40941), .B(n_40267), .Z(n_269794654));
	notech_reg int_excl_reg_5(.CP(n_62293), .D(n_31796), .CD(n_61742), .Q(int_excl
		[5]));
	notech_mux2 i_37806(.S(\nbus_13565[0] ), .A(int_excl[5]), .B(n_161596310
		), .Z(n_31796));
	notech_reg fpu_reg(.CP(n_62293), .D(n_31802), .CD(n_61742), .Q(fpu));
	notech_mux2 i_37814(.S(n_3179), .A(n_42972), .B(n_58991), .Z(n_31802));
	notech_and3 i_1308(.A(n_268594642), .B(n_40938), .C(n_2905), .Z(n_269594652
		));
	notech_reg twobyte_reg(.CP(n_62293), .D(n_31808), .CD(n_61742), .Q(twobyte
		));
	notech_mux2 i_37822(.S(n_3180), .A(n_41563), .B(twobyte), .Z(n_31808));
	notech_and4 i_223227(.A(n_269394650), .B(n_3165), .C(n_3162), .D(n_3155)
		, .Z(n_269494651));
	notech_reg opz_reg_0(.CP(n_62293), .D(n_31817), .CD(n_61742), .Q(opz[0])
		);
	notech_and4 i_37832(.A(n_60056), .B(n_224396466), .C(n_18051052), .D(opz
		[0]), .Z(n_31817));
	notech_or4 i_1302(.A(n_268594642), .B(n_3137), .C(n_2906), .D(n_2898), .Z
		(n_269394650));
	notech_reg opz_reg_1(.CP(n_62293), .D(n_31820), .CD(n_61745), .Q(opz[1])
		);
	notech_mux2 i_37838(.S(\nbus_13545[1] ), .A(opz[1]), .B(n_172896422), .Z
		(n_31820));
	notech_ao4 i_191(.A(n_3139), .B(n_3146), .C(db67), .D(n_40468), .Z(n_269294649
		));
	notech_reg_set opz_reg_2(.CP(n_62293), .D(n_31826), .SD(n_61745), .Q(opz
		[2]));
	notech_mux2 i_37846(.S(\nbus_13545[1] ), .A(opz[2]), .B(n_39361), .Z(n_31826
		));
	notech_reg imm_sz_reg_0(.CP(n_62293), .D(n_31832), .CD(n_61745), .Q(imm_sz
		[0]));
	notech_mux2 i_37854(.S(n_2191), .A(n_49847), .B(imm_sz[0]), .Z(n_31832)
		);
	notech_reg imm_sz_reg_1(.CP(n_62293), .D(n_31838), .CD(n_61745), .Q(imm_sz
		[1]));
	notech_mux2 i_37862(.S(n_2191), .A(n_39363), .B(imm_sz[1]), .Z(n_31838)
		);
	notech_nand3 i_323228(.A(n_3155), .B(n_3159), .C(n_268694643), .Z(n_268994646
		));
	notech_reg imm_sz_reg_2(.CP(n_62290), .D(n_31844), .CD(n_61745), .Q(imm_sz
		[2]));
	notech_mux2 i_37870(.S(n_2191), .A(n_49859), .B(imm_sz[2]), .Z(n_31844)
		);
	notech_reg i_ptr_reg_0(.CP(n_62290), .D(n_31850), .CD(n_61745), .Q(i_ptr
		[0]));
	notech_mux2 i_37878(.S(n_223196478), .A(n_39121), .B(i_ptr[0]), .Z(n_31850
		));
	notech_reg i_ptr_reg_1(.CP(n_62290), .D(n_31856), .CD(n_61745), .Q(i_ptr
		[1]));
	notech_mux2 i_37886(.S(n_223196478), .A(n_39122), .B(i_ptr[1]), .Z(n_31856
		));
	notech_or4 i_1291(.A(n_268594642), .B(n_1644), .C(n_58991), .D(n_40499),
		 .Z(n_268694643));
	notech_reg i_ptr_reg_2(.CP(n_62290), .D(n_31862), .CD(n_61745), .Q(i_ptr
		[2]));
	notech_mux2 i_37894(.S(n_223196478), .A(n_268994646), .B(i_ptr[2]), .Z(n_31862
		));
	notech_mux2 i_523(.S(twobyte), .A(n_226996440), .B(n_2959), .Z(n_268594642
		));
	notech_reg i_ptr_reg_3(.CP(n_62290), .D(n_31871), .CD(n_61745), .Q(i_ptr
		[3]));
	notech_and2 i_37904(.A(n_223196478), .B(i_ptr[3]), .Z(n_31871));
	notech_reg idx_deco_reg_0(.CP(n_62293), .D(n_31874), .CD(n_61745), .Q(idx_deco
		[0]));
	notech_mux2 i_37910(.S(n_3181), .A(n_42947), .B(idx_deco[0]), .Z(n_31874
		));
	notech_reg idx_deco_reg_1(.CP(n_62293), .D(n_31880), .CD(n_61745), .Q(idx_deco
		[1]));
	notech_mux2 i_37918(.S(n_3181), .A(n_42953), .B(idx_deco[1]), .Z(n_31880
		));
	notech_nao3 i_327190(.A(n_1940), .B(n_3150), .C(n_2027), .Z(n_268294639)
		);
	notech_reg fsm_reg_0(.CP(n_62293), .D(n_31886), .CD(n_61745), .Q(fsm[0])
		);
	notech_mux2 i_37926(.S(n_3182), .A(n_39118), .B(fsm[0]), .Z(n_31886));
	notech_reg fsm_reg_1(.CP(n_62293), .D(n_31892), .CD(n_61745), .Q(fsm[1])
		);
	notech_mux2 i_37934(.S(n_3182), .A(n_39119), .B(fsm[1]), .Z(n_31892));
	notech_ao4 i_127672(.A(n_58152), .B(n_39248), .C(n_227894235), .D(n_59534
		), .Z(n_268094637));
	notech_reg fsm_reg_2(.CP(n_62293), .D(n_31898), .CD(n_61745), .Q(fsm[2])
		);
	notech_mux2 i_37942(.S(n_3182), .A(n_39120), .B(fsm[2]), .Z(n_31898));
	notech_reg fsm_reg_3(.CP(n_62260), .D(n_31907), .CD(n_61742), .Q(fsm[3])
		);
	notech_and2 i_37952(.A(n_3182), .B(fsm[3]), .Z(n_31907));
	notech_ao4 i_227673(.A(n_58164), .B(n_39249), .C(n_228694243), .D(n_59534
		), .Z(n_267894635));
	notech_reg fsm_reg_4(.CP(n_62260), .D(n_31913), .CD(n_61742), .Q(fsm[4])
		);
	notech_and2 i_37960(.A(n_3182), .B(fsm[4]), .Z(n_31913));
	notech_reg repz_reg(.CP(n_62260), .D(n_31916), .CD(n_61745), .Q(repz));
	notech_mux2 i_37966(.S(n_44067), .A(repz), .B(n_172796421), .Z(n_31916)
		);
	notech_ao4 i_327674(.A(n_58164), .B(n_39251), .C(n_229494251), .D(n_59536
		), .Z(n_267694633));
	notech_reg rep_reg(.CP(n_62260), .D(n_31922), .CD(n_61745), .Q(rep));
	notech_mux2 i_37974(.S(n_44067), .A(rep), .B(n_41563), .Z(n_31922));
	notech_reg pfx_sz_reg_0(.CP(n_62260), .D(n_31928), .CD(n_61745), .Q(pfx_sz
		[0]));
	notech_mux2 i_37982(.S(\nbus_13539[0] ), .A(pfx_sz[0]), .B(n_39131), .Z(n_31928
		));
	notech_ao4 i_427675(.A(n_58164), .B(n_39252), .C(n_230294259), .D(n_59536
		), .Z(n_267494631));
	notech_reg pfx_sz_reg_1(.CP(n_62262), .D(n_31934), .CD(n_61745), .Q(pfx_sz
		[1]));
	notech_mux2 i_37990(.S(\nbus_13539[0] ), .A(pfx_sz[1]), .B(n_39384), .Z(n_31934
		));
	notech_reg pfx_sz_reg_2(.CP(n_62262), .D(n_31940), .CD(n_61745), .Q(pfx_sz
		[2]));
	notech_mux2 i_37998(.S(\nbus_13539[0] ), .A(pfx_sz[2]), .B(n_172496418),
		 .Z(n_31940));
	notech_ao4 i_527676(.A(n_58164), .B(n_39254), .C(n_231094267), .D(n_59536
		), .Z(n_267294629));
	notech_reg pfx_sz_reg_3(.CP(n_62262), .D(n_31946), .CD(n_61728), .Q(pfx_sz
		[3]));
	notech_mux2 i_38006(.S(\nbus_13539[0] ), .A(pfx_sz[3]), .B(n_172596419),
		 .Z(n_31946));
	notech_reg pfx_sz_reg_4(.CP(n_62260), .D(n_31952), .CD(n_61712), .Q(pfx_sz
		[4]));
	notech_mux2 i_38014(.S(\nbus_13539[0] ), .A(pfx_sz[4]), .B(n_172696420),
		 .Z(n_31952));
	notech_ao4 i_627677(.A(n_58164), .B(n_39255), .C(n_231894275), .D(n_59539
		), .Z(n_267094627));
	notech_reg lenpc2_reg_0(.CP(n_62260), .D(n_31958), .CD(n_61712), .Q(lenpc2
		[0]));
	notech_mux2 i_38022(.S(n_55100), .A(lenpc2[0]), .B(n_44841), .Z(n_31958)
		);
	notech_reg lenpc2_reg_1(.CP(n_62260), .D(n_31964), .CD(n_61712), .Q(lenpc2
		[1]));
	notech_mux2 i_38030(.S(n_55100), .A(lenpc2[1]), .B(n_44847), .Z(n_31964)
		);
	notech_ao4 i_727678(.A(n_58164), .B(n_39257), .C(n_232694283), .D(n_59536
		), .Z(n_266894625));
	notech_reg lenpc2_reg_2(.CP(n_62260), .D(n_31970), .CD(n_61712), .Q(lenpc2
		[2]));
	notech_mux2 i_38038(.S(n_55100), .A(lenpc2[2]), .B(n_44853), .Z(n_31970)
		);
	notech_reg lenpc2_reg_3(.CP(n_62260), .D(n_31976), .CD(n_61712), .Q(lenpc2
		[3]));
	notech_mux2 i_38046(.S(n_55100), .A(lenpc2[3]), .B(n_44859), .Z(n_31976)
		);
	notech_ao4 i_827679(.A(n_58164), .B(n_39258), .C(n_233494291), .D(n_59536
		), .Z(n_266694623));
	notech_reg lenpc2_reg_4(.CP(n_62260), .D(n_31982), .CD(n_61714), .Q(lenpc2
		[4]));
	notech_mux2 i_38054(.S(n_55100), .A(lenpc2[4]), .B(n_44865), .Z(n_31982)
		);
	notech_reg lenpc2_reg_5(.CP(n_62260), .D(n_31988), .CD(n_61714), .Q(lenpc2
		[5]));
	notech_mux2 i_38062(.S(n_55078), .A(lenpc2[5]), .B(n_44871), .Z(n_31988)
		);
	notech_ao4 i_927680(.A(n_58164), .B(n_39260), .C(n_234294299), .D(n_59536
		), .Z(n_266494621));
	notech_reg lenpc2_reg_6(.CP(n_62260), .D(n_31998), .CD(n_61714), .Q(lenpc2
		[6]));
	notech_ao3 i_38074(.A(lenpc2[6]), .B(1'b1), .C(n_55078), .Z(n_31998));
	notech_reg lenpc2_reg_7(.CP(n_62260), .D(n_32004), .CD(n_61712), .Q(lenpc2
		[7]));
	notech_ao4 i_1027681(.A(n_58164), .B(n_39261), .C(n_235094307), .D(n_59536
		), .Z(n_266294619));
	notech_ao3 i_38082(.A(lenpc2[7]), .B(1'b1), .C(n_55078), .Z(n_32004));
	notech_reg lenpc2_reg_8(.CP(n_62260), .D(n_32010), .CD(n_61714), .Q(lenpc2
		[8]));
	notech_ao3 i_38090(.A(lenpc2[8]), .B(1'b1), .C(n_55078), .Z(n_32010));
	notech_reg lenpc2_reg_9(.CP(n_62260), .D(n_32016), .CD(n_61712), .Q(lenpc2
		[9]));
	notech_ao4 i_1127682(.A(n_58164), .B(n_39263), .C(n_235894315), .D(n_59536
		), .Z(n_266094617));
	notech_ao3 i_38098(.A(lenpc2[9]), .B(1'b1), .C(n_55078), .Z(n_32016));
	notech_reg lenpc2_reg_10(.CP(n_62260), .D(n_32022), .CD(n_61712), .Q(lenpc2
		[10]));
	notech_ao3 i_38106(.A(lenpc2[10]), .B(1'b1), .C(n_55078), .Z(n_32022));
	notech_reg lenpc2_reg_11(.CP(n_62260), .D(n_32028), .CD(n_61712), .Q(lenpc2
		[11]));
	notech_ao4 i_1227683(.A(n_58167), .B(n_39264), .C(n_236694323), .D(n_59536
		), .Z(n_265894615));
	notech_ao3 i_38114(.A(lenpc2[11]), .B(1'b1), .C(n_55078), .Z(n_32028));
	notech_reg lenpc2_reg_12(.CP(n_62262), .D(n_32034), .CD(n_61712), .Q(lenpc2
		[12]));
	notech_ao3 i_38122(.A(lenpc2[12]), .B(1'b1), .C(n_55083), .Z(n_32034));
	notech_reg lenpc2_reg_13(.CP(n_62262), .D(n_32040), .CD(n_61712), .Q(lenpc2
		[13]));
	notech_ao4 i_1327684(.A(n_58167), .B(n_39266), .C(n_237494331), .D(n_59534
		), .Z(n_265694613));
	notech_ao3 i_38130(.A(lenpc2[13]), .B(1'b1), .C(n_55083), .Z(n_32040));
	notech_reg lenpc2_reg_14(.CP(n_62262), .D(n_32046), .CD(n_61712), .Q(lenpc2
		[14]));
	notech_ao3 i_38138(.A(lenpc2[14]), .B(1'b1), .C(n_55083), .Z(n_32046));
	notech_reg lenpc2_reg_15(.CP(n_62262), .D(n_32052), .CD(n_61712), .Q(lenpc2
		[15]));
	notech_ao4 i_1427685(.A(n_58167), .B(n_39267), .C(n_238294339), .D(n_59529
		), .Z(n_265494611));
	notech_ao3 i_38146(.A(lenpc2[15]), .B(1'b1), .C(n_55078), .Z(n_32052));
	notech_reg lenpc2_reg_16(.CP(n_62262), .D(n_32058), .CD(n_61712), .Q(lenpc2
		[16]));
	notech_ao3 i_38154(.A(lenpc2[16]), .B(1'b1), .C(n_55083), .Z(n_32058));
	notech_reg lenpc2_reg_17(.CP(n_62266), .D(n_32064), .CD(n_61712), .Q(lenpc2
		[17]));
	notech_ao4 i_1627687(.A(n_58167), .B(n_39270), .C(n_239494351), .D(n_59529
		), .Z(n_265294609));
	notech_ao3 i_38162(.A(lenpc2[17]), .B(1'b1), .C(n_55083), .Z(n_32064));
	notech_reg lenpc2_reg_18(.CP(n_62266), .D(n_32070), .CD(n_61712), .Q(lenpc2
		[18]));
	notech_ao3 i_38170(.A(lenpc2[18]), .B(1'b1), .C(n_55078), .Z(n_32070));
	notech_reg lenpc2_reg_19(.CP(n_62266), .D(n_32076), .CD(n_61712), .Q(lenpc2
		[19]));
	notech_ao4 i_1827689(.A(n_58167), .B(n_39273), .C(n_240894365), .D(n_59529
		), .Z(n_265094607));
	notech_ao3 i_38178(.A(lenpc2[19]), .B(1'b1), .C(n_55078), .Z(n_32076));
	notech_reg lenpc2_reg_20(.CP(n_62262), .D(n_32082), .CD(n_61714), .Q(lenpc2
		[20]));
	notech_ao3 i_38186(.A(lenpc2[20]), .B(1'b1), .C(n_55078), .Z(n_32082));
	notech_reg lenpc2_reg_21(.CP(n_62266), .D(n_32088), .CD(n_61718), .Q(lenpc2
		[21]));
	notech_ao4 i_1927690(.A(n_58164), .B(n_39275), .C(n_241894375), .D(n_59529
		), .Z(n_264894605));
	notech_ao3 i_38194(.A(lenpc2[21]), .B(1'b1), .C(n_55077), .Z(n_32088));
	notech_reg lenpc2_reg_22(.CP(n_62262), .D(n_32094), .CD(n_61714), .Q(lenpc2
		[22]));
	notech_ao3 i_38202(.A(lenpc2[22]), .B(1'b1), .C(n_55077), .Z(n_32094));
	notech_reg lenpc2_reg_23(.CP(n_62262), .D(n_32100), .CD(n_61714), .Q(lenpc2
		[23]));
	notech_ao4 i_2027691(.A(n_58164), .B(n_39276), .C(n_242894385), .D(n_59529
		), .Z(n_264694603));
	notech_ao3 i_38210(.A(lenpc2[23]), .B(1'b1), .C(n_55077), .Z(n_32100));
	notech_reg lenpc2_reg_24(.CP(n_62262), .D(n_32106), .CD(n_61714), .Q(lenpc2
		[24]));
	notech_ao3 i_38218(.A(lenpc2[24]), .B(1'b1), .C(n_55078), .Z(n_32106));
	notech_reg lenpc2_reg_25(.CP(n_62262), .D(n_32112), .CD(n_61718), .Q(lenpc2
		[25]));
	notech_ao4 i_2127692(.A(n_58164), .B(n_39278), .C(n_243894395), .D(n_59529
		), .Z(n_264494601));
	notech_ao3 i_38226(.A(lenpc2[25]), .B(1'b1), .C(n_55078), .Z(n_32112));
	notech_reg lenpc2_reg_26(.CP(n_62262), .D(n_32118), .CD(n_61718), .Q(lenpc2
		[26]));
	notech_ao3 i_38234(.A(lenpc2[26]), .B(1'b1), .C(n_55078), .Z(n_32118));
	notech_reg lenpc2_reg_27(.CP(n_62262), .D(n_32124), .CD(n_61718), .Q(lenpc2
		[27]));
	notech_ao4 i_2227693(.A(n_58167), .B(n_39279), .C(n_244894405), .D(n_59529
		), .Z(n_264294599));
	notech_ao3 i_38242(.A(lenpc2[27]), .B(1'b1), .C(n_55078), .Z(n_32124));
	notech_reg lenpc2_reg_28(.CP(n_62262), .D(n_32130), .CD(n_61718), .Q(lenpc2
		[28]));
	notech_ao3 i_38250(.A(lenpc2[28]), .B(1'b1), .C(n_55078), .Z(n_32130));
	notech_reg lenpc2_reg_29(.CP(n_62262), .D(n_32136), .CD(n_61718), .Q(lenpc2
		[29]));
	notech_ao4 i_2327694(.A(n_58164), .B(n_39281), .C(n_245894415), .D(n_59529
		), .Z(n_264094597));
	notech_ao3 i_38258(.A(lenpc2[29]), .B(1'b1), .C(n_55078), .Z(n_32136));
	notech_reg lenpc2_reg_30(.CP(n_62262), .D(n_32142), .CD(n_61714), .Q(lenpc2
		[30]));
	notech_ao3 i_38266(.A(lenpc2[30]), .B(1'b1), .C(n_55078), .Z(n_32142));
	notech_reg lenpc2_reg_31(.CP(n_62262), .D(n_32148), .CD(n_61714), .Q(lenpc2
		[31]));
	notech_ao4 i_2427695(.A(n_58162), .B(n_39282), .C(n_246894425), .D(n_59529
		), .Z(n_263894595));
	notech_ao3 i_38274(.A(lenpc2[31]), .B(1'b1), .C(n_55083), .Z(n_32148));
	notech_reg reps2_reg_0(.CP(n_62262), .D(n_32150), .CD(n_61714), .Q(reps2
		[0]));
	notech_mux2 i_38278(.S(n_55088), .A(reps2[0]), .B(n_49787), .Z(n_32150)
		);
	notech_reg reps2_reg_1(.CP(n_62260), .D(n_32156), .CD(n_61714), .Q(reps2
		[1]));
	notech_mux2 i_38286(.S(n_55088), .A(reps2[1]), .B(n_49793), .Z(n_32156)
		);
	notech_ao4 i_2527696(.A(n_58157), .B(n_39284), .C(n_247894435), .D(n_59529
		), .Z(n_263694593));
	notech_reg reps2_reg_2(.CP(n_62255), .D(n_32162), .CD(n_61714), .Q(reps2
		[2]));
	notech_mux2 i_38294(.S(n_55088), .A(reps2[2]), .B(n_49799), .Z(n_32162)
		);
	notech_reg reps1_reg_0(.CP(n_62255), .D(n_32168), .CD(n_61714), .Q(reps1
		[0]));
	notech_mux2 i_38302(.S(n_58326), .A(reps1[0]), .B(n_39117), .Z(n_32168)
		);
	notech_ao4 i_2727698(.A(n_58157), .B(n_39287), .C(n_248894445), .D(n_59534
		), .Z(n_263494591));
	notech_reg reps1_reg_1(.CP(n_62255), .D(n_32174), .CD(n_61714), .Q(reps1
		[1]));
	notech_mux2 i_38310(.S(n_58326), .A(reps1[1]), .B(n_39417), .Z(n_32174)
		);
	notech_reg reps1_reg_2(.CP(n_62255), .D(n_32180), .CD(n_61714), .Q(reps1
		[2]));
	notech_mux2 i_38318(.S(n_58326), .A(reps1[2]), .B(n_39419), .Z(n_32180)
		);
	notech_ao4 i_2827699(.A(n_58162), .B(n_39288), .C(n_249894455), .D(n_59534
		), .Z(n_263294589));
	notech_reg inst_deco2_reg_0(.CP(n_62255), .D(n_32186), .CD(n_61714), .Q(inst_deco2
		[0]));
	notech_mux2 i_38326(.S(n_55088), .A(inst_deco2[0]), .B(n_43192), .Z(n_32186
		));
	notech_reg inst_deco2_reg_1(.CP(n_62255), .D(n_32192), .CD(n_61714), .Q(inst_deco2
		[1]));
	notech_mux2 i_38334(.S(n_55088), .A(inst_deco2[1]), .B(n_43198), .Z(n_32192
		));
	notech_ao4 i_2927700(.A(n_58162), .B(n_39290), .C(n_250894465), .D(n_59534
		), .Z(n_263094587));
	notech_reg inst_deco2_reg_2(.CP(n_62255), .D(n_32198), .CD(n_61714), .Q(inst_deco2
		[2]));
	notech_mux2 i_38342(.S(n_55088), .A(inst_deco2[2]), .B(n_43204), .Z(n_32198
		));
	notech_reg inst_deco2_reg_3(.CP(n_62255), .D(n_32204), .CD(n_61707), .Q(inst_deco2
		[3]));
	notech_mux2 i_38350(.S(n_55088), .A(inst_deco2[3]), .B(n_43210), .Z(n_32204
		));
	notech_ao4 i_3027701(.A(n_58162), .B(n_39291), .C(n_251894475), .D(n_59534
		), .Z(n_262894585));
	notech_reg inst_deco2_reg_4(.CP(n_62255), .D(n_32210), .CD(n_61707), .Q(inst_deco2
		[4]));
	notech_mux2 i_38358(.S(n_55088), .A(inst_deco2[4]), .B(n_43216), .Z(n_32210
		));
	notech_reg inst_deco2_reg_5(.CP(n_62255), .D(n_32216), .CD(n_61707), .Q(inst_deco2
		[5]));
	notech_mux2 i_38366(.S(n_55089), .A(inst_deco2[5]), .B(n_43222), .Z(n_32216
		));
	notech_ao4 i_3127702(.A(n_58157), .B(n_39293), .C(n_252894485), .D(n_59534
		), .Z(n_262694583));
	notech_reg inst_deco2_reg_6(.CP(n_62255), .D(n_32222), .CD(n_61707), .Q(inst_deco2
		[6]));
	notech_mux2 i_38374(.S(n_55089), .A(inst_deco2[6]), .B(n_43228), .Z(n_32222
		));
	notech_reg inst_deco2_reg_7(.CP(n_62255), .D(n_32228), .CD(n_61707), .Q(inst_deco2
		[7]));
	notech_mux2 i_38382(.S(n_55088), .A(inst_deco2[7]), .B(n_43234), .Z(n_32228
		));
	notech_ao4 i_3227703(.A(n_58157), .B(n_39294), .C(n_254094497), .D(n_59529
		), .Z(n_262494581));
	notech_reg inst_deco2_reg_8(.CP(n_62255), .D(n_32234), .CD(n_61707), .Q(inst_deco2
		[8]));
	notech_mux2 i_38390(.S(n_55088), .A(inst_deco2[8]), .B(n_43240), .Z(n_32234
		));
	notech_reg inst_deco2_reg_9(.CP(n_62255), .D(n_32240), .CD(n_61707), .Q(inst_deco2
		[9]));
	notech_mux2 i_38398(.S(n_55088), .A(inst_deco2[9]), .B(n_43246), .Z(n_32240
		));
	notech_ao4 i_3327704(.A(n_58157), .B(n_39296), .C(n_54557), .D(n_40326),
		 .Z(n_262294579));
	notech_reg inst_deco2_reg_10(.CP(n_62252), .D(n_32246), .CD(n_61707), .Q
		(inst_deco2[10]));
	notech_mux2 i_38406(.S(n_55083), .A(inst_deco2[10]), .B(n_43252), .Z(n_32246
		));
	notech_reg inst_deco2_reg_11(.CP(n_62252), .D(n_32252), .CD(n_61707), .Q
		(inst_deco2[11]));
	notech_mux2 i_38414(.S(n_55083), .A(inst_deco2[11]), .B(n_43258), .Z(n_32252
		));
	notech_ao4 i_3427705(.A(n_58157), .B(n_39297), .C(n_54557), .D(n_40319),
		 .Z(n_262094577));
	notech_reg inst_deco2_reg_12(.CP(n_62255), .D(n_32258), .CD(n_61707), .Q
		(inst_deco2[12]));
	notech_mux2 i_38422(.S(n_55083), .A(inst_deco2[12]), .B(n_3440), .Z(n_32258
		));
	notech_reg inst_deco2_reg_13(.CP(n_62255), .D(n_32264), .CD(n_61707), .Q
		(inst_deco2[13]));
	notech_mux2 i_38430(.S(n_55083), .A(inst_deco2[13]), .B(n_43270), .Z(n_32264
		));
	notech_ao4 i_3527706(.A(n_58157), .B(n_39299), .C(n_54557), .D(n_40279),
		 .Z(n_261894575));
	notech_reg inst_deco2_reg_14(.CP(n_62255), .D(n_32270), .CD(n_61704), .Q
		(inst_deco2[14]));
	notech_mux2 i_38438(.S(n_55083), .A(inst_deco2[14]), .B(n_43276), .Z(n_32270
		));
	notech_reg inst_deco2_reg_15(.CP(n_62255), .D(n_32276), .CD(n_61704), .Q
		(inst_deco2[15]));
	notech_mux2 i_38446(.S(n_55083), .A(inst_deco2[15]), .B(n_43282), .Z(n_32276
		));
	notech_reg inst_deco2_reg_16(.CP(n_62255), .D(n_32282), .CD(n_61704), .Q
		(inst_deco2[16]));
	notech_mux2 i_38454(.S(n_55088), .A(inst_deco2[16]), .B(n_3435), .Z(n_32282
		));
	notech_reg inst_deco2_reg_17(.CP(n_62257), .D(n_32288), .CD(n_61704), .Q
		(inst_deco2[17]));
	notech_mux2 i_38462(.S(n_55088), .A(inst_deco2[17]), .B(n_43294), .Z(n_32288
		));
	notech_and2 i_264(.A(in128[42]), .B(n_2941), .Z(n_261494571));
	notech_reg inst_deco2_reg_18(.CP(n_62257), .D(n_32294), .CD(n_61704), .Q
		(inst_deco2[18]));
	notech_mux2 i_38470(.S(n_55088), .A(inst_deco2[18]), .B(n_43300), .Z(n_32294
		));
	notech_ao4 i_3727708(.A(n_58162), .B(n_39302), .C(n_54557), .D(n_40309),
		 .Z(n_261394570));
	notech_reg inst_deco2_reg_19(.CP(n_62257), .D(n_32300), .CD(n_61707), .Q
		(inst_deco2[19]));
	notech_mux2 i_38478(.S(n_55088), .A(inst_deco2[19]), .B(n_43306), .Z(n_32300
		));
	notech_reg inst_deco2_reg_20(.CP(n_62257), .D(n_32306), .CD(n_61707), .Q
		(inst_deco2[20]));
	notech_mux2 i_38486(.S(n_55088), .A(inst_deco2[20]), .B(n_3431), .Z(n_32306
		));
	notech_ao4 i_3827709(.A(n_58162), .B(n_39303), .C(n_54557), .D(n_40307),
		 .Z(n_261194568));
	notech_reg inst_deco2_reg_21(.CP(n_62257), .D(n_32312), .CD(n_61707), .Q
		(inst_deco2[21]));
	notech_mux2 i_38494(.S(n_55088), .A(inst_deco2[21]), .B(n_43318), .Z(n_32312
		));
	notech_reg inst_deco2_reg_22(.CP(n_62257), .D(n_32318), .CD(n_61707), .Q
		(inst_deco2[22]));
	notech_mux2 i_38502(.S(n_55088), .A(inst_deco2[22]), .B(n_43324), .Z(n_32318
		));
	notech_ao4 i_3927710(.A(n_58162), .B(n_39305), .C(n_54557), .D(n_40304),
		 .Z(n_260994566));
	notech_reg inst_deco2_reg_23(.CP(n_62260), .D(n_32324), .CD(n_61707), .Q
		(inst_deco2[23]));
	notech_mux2 i_38510(.S(n_55101), .A(inst_deco2[23]), .B(n_43330), .Z(n_32324
		));
	notech_reg inst_deco2_reg_24(.CP(n_62257), .D(n_32330), .CD(n_61709), .Q
		(inst_deco2[24]));
	notech_mux2 i_38518(.S(n_55117), .A(inst_deco2[24]), .B(n_43336), .Z(n_32330
		));
	notech_ao4 i_4027711(.A(n_58162), .B(n_39306), .C(n_54557), .D(n_40300),
		 .Z(n_260794564));
	notech_reg inst_deco2_reg_25(.CP(n_62257), .D(n_32336), .CD(n_61709), .Q
		(inst_deco2[25]));
	notech_mux2 i_38526(.S(n_55122), .A(inst_deco2[25]), .B(n_43342), .Z(n_32336
		));
	notech_reg inst_deco2_reg_26(.CP(n_62257), .D(n_32342), .CD(n_61709), .Q
		(inst_deco2[26]));
	notech_mux2 i_38534(.S(n_55122), .A(inst_deco2[26]), .B(n_3428), .Z(n_32342
		));
	notech_ao4 i_4127712(.A(n_58162), .B(n_39308), .C(n_2948), .D(n_40298), 
		.Z(n_260594562));
	notech_reg inst_deco2_reg_27(.CP(n_62257), .D(n_32348), .CD(n_61709), .Q
		(inst_deco2[27]));
	notech_mux2 i_38542(.S(n_55117), .A(inst_deco2[27]), .B(n_3426), .Z(n_32348
		));
	notech_reg inst_deco2_reg_28(.CP(n_62257), .D(n_32354), .CD(n_61709), .Q
		(inst_deco2[28]));
	notech_mux2 i_38550(.S(n_55117), .A(inst_deco2[28]), .B(n_3424), .Z(n_32354
		));
	notech_ao4 i_4327714(.A(n_58162), .B(n_39311), .C(n_2948), .D(n_40295), 
		.Z(n_260394560));
	notech_reg inst_deco2_reg_29(.CP(n_62257), .D(n_32360), .CD(n_61709), .Q
		(inst_deco2[29]));
	notech_mux2 i_38558(.S(n_55117), .A(inst_deco2[29]), .B(n_3422), .Z(n_32360
		));
	notech_reg inst_deco2_reg_30(.CP(n_62257), .D(n_32366), .CD(n_61712), .Q
		(inst_deco2[30]));
	notech_mux2 i_38566(.S(n_55122), .A(inst_deco2[30]), .B(n_3420), .Z(n_32366
		));
	notech_ao4 i_4427715(.A(n_58162), .B(n_39312), .C(n_2948), .D(n_40488), 
		.Z(n_260194558));
	notech_reg inst_deco2_reg_31(.CP(n_62257), .D(n_32372), .CD(n_61709), .Q
		(inst_deco2[31]));
	notech_mux2 i_38574(.S(n_55122), .A(inst_deco2[31]), .B(n_3418), .Z(n_32372
		));
	notech_reg inst_deco2_reg_32(.CP(n_62257), .D(n_32378), .CD(n_61709), .Q
		(inst_deco2[32]));
	notech_mux2 i_38582(.S(n_55122), .A(inst_deco2[32]), .B(n_43384), .Z(n_32378
		));
	notech_ao4 i_4527716(.A(n_58162), .B(n_39314), .C(n_2948), .D(n_40281), 
		.Z(n_259994556));
	notech_reg inst_deco2_reg_33(.CP(n_62257), .D(n_32384), .CD(n_61709), .Q
		(inst_deco2[33]));
	notech_mux2 i_38590(.S(n_55122), .A(inst_deco2[33]), .B(n_3416), .Z(n_32384
		));
	notech_reg inst_deco2_reg_34(.CP(n_62257), .D(n_32390), .CD(n_61709), .Q
		(inst_deco2[34]));
	notech_mux2 i_38598(.S(n_55122), .A(inst_deco2[34]), .B(n_3414), .Z(n_32390
		));
	notech_reg inst_deco2_reg_35(.CP(n_62257), .D(n_32396), .CD(n_61709), .Q
		(inst_deco2[35]));
	notech_mux2 i_38606(.S(n_55122), .A(inst_deco2[35]), .B(n_3412), .Z(n_32396
		));
	notech_reg inst_deco2_reg_36(.CP(n_62257), .D(n_32402), .CD(n_61709), .Q
		(inst_deco2[36]));
	notech_mux2 i_38614(.S(n_55122), .A(inst_deco2[36]), .B(n_3410), .Z(n_32402
		));
	notech_and2 i_263(.A(in128[60]), .B(n_2947), .Z(n_259594552));
	notech_reg inst_deco2_reg_37(.CP(n_62257), .D(n_32408), .CD(n_61709), .Q
		(inst_deco2[37]));
	notech_mux2 i_38622(.S(n_55112), .A(inst_deco2[37]), .B(n_43414), .Z(n_32408
		));
	notech_ao4 i_4727718(.A(n_58162), .B(n_39317), .C(n_2948), .D(n_40293), 
		.Z(n_259494551));
	notech_reg inst_deco2_reg_38(.CP(n_62273), .D(n_32414), .CD(n_61707), .Q
		(inst_deco2[38]));
	notech_mux2 i_38630(.S(n_55112), .A(inst_deco2[38]), .B(n_3408), .Z(n_32414
		));
	notech_reg inst_deco2_reg_39(.CP(n_62273), .D(n_32420), .CD(n_61707), .Q
		(inst_deco2[39]));
	notech_mux2 i_38638(.S(n_55117), .A(inst_deco2[39]), .B(n_3406), .Z(n_32420
		));
	notech_ao4 i_4827719(.A(n_58162), .B(n_39318), .C(n_2948), .D(n_40290), 
		.Z(n_259294549));
	notech_reg inst_deco2_reg_40(.CP(n_62273), .D(n_32426), .CD(n_61709), .Q
		(inst_deco2[40]));
	notech_mux2 i_38646(.S(n_55112), .A(inst_deco2[40]), .B(n_3404), .Z(n_32426
		));
	notech_reg inst_deco2_reg_41(.CP(n_62271), .D(n_32432), .CD(n_61709), .Q
		(inst_deco2[41]));
	notech_mux2 i_38654(.S(n_55112), .A(inst_deco2[41]), .B(n_3402), .Z(n_32432
		));
	notech_ao4 i_123166(.A(n_258994546), .B(n_3147), .C(n_269294649), .D(n_40938
		), .Z(n_259094547));
	notech_reg inst_deco2_reg_42(.CP(n_62271), .D(n_32438), .CD(n_61709), .Q
		(inst_deco2[42]));
	notech_mux2 i_38662(.S(n_55112), .A(inst_deco2[42]), .B(n_3400), .Z(n_32438
		));
	notech_ao4 i_261(.A(n_3139), .B(n_258694543), .C(db67), .D(n_40468), .Z(n_258994546
		));
	notech_reg inst_deco2_reg_43(.CP(n_62273), .D(n_32444), .CD(n_61709), .Q
		(inst_deco2[43]));
	notech_mux2 i_38670(.S(n_55117), .A(inst_deco2[43]), .B(n_3398), .Z(n_32444
		));
	notech_reg inst_deco2_reg_44(.CP(n_62273), .D(n_32450), .CD(n_61709), .Q
		(inst_deco2[44]));
	notech_mux2 i_38678(.S(n_55117), .A(inst_deco2[44]), .B(n_3396), .Z(n_32450
		));
	notech_reg inst_deco2_reg_45(.CP(n_62273), .D(n_32456), .CD(n_61718), .Q
		(inst_deco2[45]));
	notech_mux2 i_38686(.S(n_55117), .A(inst_deco2[45]), .B(n_3394), .Z(n_32456
		));
	notech_nor2 i_262(.A(n_1772), .B(n_258494541), .Z(n_258694543));
	notech_reg inst_deco2_reg_46(.CP(n_62273), .D(n_32462), .CD(n_61725), .Q
		(inst_deco2[46]));
	notech_mux2 i_38694(.S(n_55117), .A(inst_deco2[46]), .B(n_3392), .Z(n_32462
		));
	notech_reg inst_deco2_reg_47(.CP(n_62273), .D(n_32468), .CD(n_61725), .Q
		(inst_deco2[47]));
	notech_mux2 i_38702(.S(n_55117), .A(inst_deco2[47]), .B(n_3390), .Z(n_32468
		));
	notech_ao3 i_1134(.A(n_40943), .B(n_40941), .C(n_1925), .Z(n_258494541)
		);
	notech_reg inst_deco2_reg_48(.CP(n_62271), .D(n_32474), .CD(n_61725), .Q
		(inst_deco2[48]));
	notech_mux2 i_38710(.S(n_55117), .A(inst_deco2[48]), .B(n_3388), .Z(n_32474
		));
	notech_reg inst_deco2_reg_49(.CP(n_62271), .D(n_32480), .CD(n_61725), .Q
		(inst_deco2[49]));
	notech_mux2 i_38718(.S(n_55117), .A(inst_deco2[49]), .B(n_3386), .Z(n_32480
		));
	notech_or4 i_1106(.A(in128[17]), .B(n_40944), .C(n_40729), .D(n_40727), 
		.Z(n_258294539));
	notech_reg inst_deco2_reg_50(.CP(n_62271), .D(n_32486), .CD(n_61725), .Q
		(inst_deco2[50]));
	notech_mux2 i_38726(.S(n_55122), .A(inst_deco2[50]), .B(n_3384), .Z(n_32486
		));
	notech_nao3 i_1101(.A(\fpu_modrm[0] ), .B(n_3142), .C(\fpu_modrm[1] ), .Z
		(n_258194538));
	notech_reg inst_deco2_reg_51(.CP(n_62271), .D(n_32492), .CD(n_61725), .Q
		(inst_deco2[51]));
	notech_mux2 i_38734(.S(n_55123), .A(inst_deco2[51]), .B(n_3382), .Z(n_32492
		));
	notech_mux2 i_70614(.S(adz), .A(n_41563), .B(n_1753), .Z(n_258094537));
	notech_reg inst_deco2_reg_52(.CP(n_62271), .D(n_32498), .CD(n_61725), .Q
		(inst_deco2[52]));
	notech_mux2 i_38742(.S(n_55123), .A(inst_deco2[52]), .B(n_3380), .Z(n_32498
		));
	notech_reg inst_deco2_reg_53(.CP(n_62271), .D(n_32504), .CD(n_61725), .Q
		(inst_deco2[53]));
	notech_mux2 i_38750(.S(n_55123), .A(inst_deco2[53]), .B(n_3378), .Z(n_32504
		));
	notech_reg inst_deco2_reg_54(.CP(n_62271), .D(n_32510), .CD(n_61725), .Q
		(inst_deco2[54]));
	notech_mux2 i_38758(.S(n_55123), .A(inst_deco2[54]), .B(n_3376), .Z(n_32510
		));
	notech_reg inst_deco2_reg_55(.CP(n_62271), .D(n_32516), .CD(n_61725), .Q
		(inst_deco2[55]));
	notech_mux2 i_38766(.S(n_55123), .A(inst_deco2[55]), .B(n_3374), .Z(n_32516
		));
	notech_reg inst_deco2_reg_56(.CP(n_62271), .D(n_32522), .CD(n_61723), .Q
		(inst_deco2[56]));
	notech_mux2 i_38774(.S(n_55123), .A(inst_deco2[56]), .B(n_3372), .Z(n_32522
		));
	notech_and2 i_247(.A(in128[63]), .B(n_2947), .Z(n_257594532));
	notech_reg inst_deco2_reg_57(.CP(n_62271), .D(n_32528), .CD(n_61723), .Q
		(inst_deco2[57]));
	notech_mux2 i_38782(.S(n_55123), .A(inst_deco2[57]), .B(n_3370), .Z(n_32528
		));
	notech_reg inst_deco2_reg_58(.CP(n_62271), .D(n_32534), .CD(n_61723), .Q
		(inst_deco2[58]));
	notech_mux2 i_38790(.S(n_55123), .A(inst_deco2[58]), .B(n_3368), .Z(n_32534
		));
	notech_reg inst_deco2_reg_59(.CP(n_62276), .D(n_32540), .CD(n_61723), .Q
		(inst_deco2[59]));
	notech_mux2 i_38798(.S(n_55123), .A(inst_deco2[59]), .B(n_3366), .Z(n_32540
		));
	notech_and2 i_246(.A(in128[62]), .B(n_2947), .Z(n_257294529));
	notech_reg inst_deco2_reg_60(.CP(n_62276), .D(n_32546), .CD(n_61723), .Q
		(inst_deco2[60]));
	notech_mux2 i_38806(.S(n_55123), .A(inst_deco2[60]), .B(n_3364), .Z(n_32546
		));
	notech_reg inst_deco2_reg_61(.CP(n_62276), .D(n_32552), .CD(n_61723), .Q
		(inst_deco2[61]));
	notech_mux2 i_38814(.S(n_55123), .A(inst_deco2[61]), .B(n_3362), .Z(n_32552
		));
	notech_reg inst_deco2_reg_62(.CP(n_62273), .D(n_32558), .CD(n_61723), .Q
		(inst_deco2[62]));
	notech_mux2 i_38822(.S(n_55123), .A(inst_deco2[62]), .B(n_3360), .Z(n_32558
		));
	notech_and2 i_245(.A(in128[58]), .B(n_2947), .Z(n_256994526));
	notech_reg inst_deco2_reg_63(.CP(n_62276), .D(n_32564), .CD(n_61723), .Q
		(inst_deco2[63]));
	notech_mux2 i_38830(.S(n_55123), .A(inst_deco2[63]), .B(n_3358), .Z(n_32564
		));
	notech_reg inst_deco2_reg_64(.CP(n_62276), .D(n_32570), .CD(n_61723), .Q
		(inst_deco2[64]));
	notech_mux2 i_38838(.S(n_55122), .A(inst_deco2[64]), .B(n_3356), .Z(n_32570
		));
	notech_reg inst_deco2_reg_65(.CP(n_62276), .D(n_32576), .CD(n_61723), .Q
		(inst_deco2[65]));
	notech_mux2 i_38846(.S(n_55122), .A(inst_deco2[65]), .B(n_3354), .Z(n_32576
		));
	notech_and2 i_244(.A(in128[56]), .B(n_2947), .Z(n_256694523));
	notech_reg inst_deco2_reg_66(.CP(n_62276), .D(n_32582), .CD(n_61723), .Q
		(inst_deco2[66]));
	notech_mux2 i_38854(.S(n_55122), .A(inst_deco2[66]), .B(n_3352), .Z(n_32582
		));
	notech_reg inst_deco2_reg_67(.CP(n_62276), .D(n_32588), .CD(n_61728), .Q
		(inst_deco2[67]));
	notech_mux2 i_38862(.S(n_55122), .A(inst_deco2[67]), .B(n_3350), .Z(n_32588
		));
	notech_reg inst_deco2_reg_68(.CP(n_62276), .D(n_32594), .CD(n_61728), .Q
		(inst_deco2[68]));
	notech_mux2 i_38870(.S(n_55122), .A(inst_deco2[68]), .B(n_43600), .Z(n_32594
		));
	notech_and2 i_243(.A(in128[47]), .B(n_2941), .Z(n_256394520));
	notech_reg inst_deco2_reg_69(.CP(n_62273), .D(n_32600), .CD(n_61728), .Q
		(inst_deco2[69]));
	notech_mux2 i_38878(.S(n_55122), .A(inst_deco2[69]), .B(n_43606), .Z(n_32600
		));
	notech_reg inst_deco2_reg_70(.CP(n_62273), .D(n_32606), .CD(n_61728), .Q
		(inst_deco2[70]));
	notech_mux2 i_38886(.S(n_55122), .A(inst_deco2[70]), .B(n_43612), .Z(n_32606
		));
	notech_reg inst_deco2_reg_71(.CP(n_62273), .D(n_32612), .CD(n_61728), .Q
		(inst_deco2[71]));
	notech_mux2 i_38894(.S(n_55123), .A(inst_deco2[71]), .B(n_43618), .Z(n_32612
		));
	notech_and2 i_242(.A(n_2941), .B(in128[46]), .Z(n_256094517));
	notech_reg inst_deco2_reg_72(.CP(n_62273), .D(n_32618), .CD(n_61728), .Q
		(inst_deco2[72]));
	notech_mux2 i_38902(.S(n_55123), .A(inst_deco2[72]), .B(n_43624), .Z(n_32618
		));
	notech_reg inst_deco2_reg_73(.CP(n_62273), .D(n_32624), .CD(n_61728), .Q
		(inst_deco2[73]));
	notech_mux2 i_38910(.S(n_55123), .A(inst_deco2[73]), .B(n_43630), .Z(n_32624
		));
	notech_reg inst_deco2_reg_74(.CP(n_62273), .D(n_32630), .CD(n_61728), .Q
		(inst_deco2[74]));
	notech_mux2 i_38918(.S(n_55122), .A(inst_deco2[74]), .B(n_43636), .Z(n_32630
		));
	notech_and2 i_241(.A(n_3122), .B(in128[53]), .Z(n_255794514));
	notech_reg inst_deco2_reg_75(.CP(n_62273), .D(n_32636), .CD(n_61728), .Q
		(inst_deco2[75]));
	notech_mux2 i_38926(.S(n_55123), .A(inst_deco2[75]), .B(n_43642), .Z(n_32636
		));
	notech_reg inst_deco2_reg_76(.CP(n_62273), .D(n_32642), .CD(n_61728), .Q
		(inst_deco2[76]));
	notech_mux2 i_38934(.S(n_55123), .A(inst_deco2[76]), .B(n_43648), .Z(n_32642
		));
	notech_reg inst_deco2_reg_77(.CP(n_62273), .D(n_32648), .CD(n_61728), .Q
		(inst_deco2[77]));
	notech_mux2 i_38942(.S(n_55106), .A(inst_deco2[77]), .B(n_43654), .Z(n_32648
		));
	notech_and2 i_240(.A(n_2941), .B(in128[44]), .Z(n_255494511));
	notech_reg inst_deco2_reg_78(.CP(n_62273), .D(n_32654), .CD(n_61725), .Q
		(inst_deco2[78]));
	notech_mux2 i_38950(.S(n_55106), .A(inst_deco2[78]), .B(n_43660), .Z(n_32654
		));
	notech_reg inst_deco2_reg_79(.CP(n_62273), .D(n_32660), .CD(n_61725), .Q
		(inst_deco2[79]));
	notech_mux2 i_38958(.S(n_55106), .A(inst_deco2[79]), .B(n_43666), .Z(n_32660
		));
	notech_reg inst_deco2_reg_80(.CP(n_62271), .D(n_32666), .CD(n_61725), .Q
		(inst_deco2[80]));
	notech_mux2 i_38966(.S(n_55106), .A(inst_deco2[80]), .B(n_43672), .Z(n_32666
		));
	notech_and2 i_239(.A(n_2941), .B(in128[43]), .Z(n_255194508));
	notech_reg inst_deco2_reg_81(.CP(n_62266), .D(n_32672), .CD(n_61725), .Q
		(inst_deco2[81]));
	notech_mux2 i_38974(.S(n_55106), .A(inst_deco2[81]), .B(n_43678), .Z(n_32672
		));
	notech_reg inst_deco2_reg_82(.CP(n_62266), .D(n_32678), .CD(n_61725), .Q
		(inst_deco2[82]));
	notech_mux2 i_38982(.S(n_55106), .A(inst_deco2[82]), .B(n_43684), .Z(n_32678
		));
	notech_reg inst_deco2_reg_83(.CP(n_62266), .D(n_32684), .CD(n_61725), .Q
		(inst_deco2[83]));
	notech_mux2 i_38990(.S(n_55106), .A(inst_deco2[83]), .B(n_43690), .Z(n_32684
		));
	notech_and2 i_238(.A(n_3122), .B(in128[49]), .Z(n_254894505));
	notech_reg inst_deco2_reg_84(.CP(n_62266), .D(n_32690), .CD(n_61725), .Q
		(inst_deco2[84]));
	notech_mux2 i_38998(.S(n_55111), .A(inst_deco2[84]), .B(n_3332), .Z(n_32690
		));
	notech_reg inst_deco2_reg_85(.CP(n_62266), .D(n_32696), .CD(n_61725), .Q
		(inst_deco2[85]));
	notech_mux2 i_39006(.S(n_55111), .A(inst_deco2[85]), .B(n_43702), .Z(n_32696
		));
	notech_reg inst_deco2_reg_86(.CP(n_62268), .D(n_32702), .CD(n_61725), .Q
		(inst_deco2[86]));
	notech_mux2 i_39014(.S(n_55111), .A(inst_deco2[86]), .B(n_3329), .Z(n_32702
		));
	notech_and2 i_237(.A(n_2941), .B(in128[40]), .Z(n_254594502));
	notech_reg inst_deco2_reg_87(.CP(n_62268), .D(n_32708), .CD(n_61725), .Q
		(inst_deco2[87]));
	notech_mux2 i_39022(.S(n_55106), .A(inst_deco2[87]), .B(n_43714), .Z(n_32708
		));
	notech_or2 i_1051(.A(n_3122), .B(n_2941), .Z(n_254494501));
	notech_reg inst_deco2_reg_88(.CP(n_62268), .D(n_32714), .CD(n_61720), .Q
		(inst_deco2[88]));
	notech_mux2 i_39030(.S(n_55106), .A(inst_deco2[88]), .B(n_3326), .Z(n_32714
		));
	notech_and3 i_12(.A(n_40593), .B(imm_sz[0]), .C(imm_sz[1]), .Z(n_254394500
		));
	notech_reg inst_deco2_reg_89(.CP(n_62268), .D(n_32720), .CD(n_61720), .Q
		(inst_deco2[89]));
	notech_mux2 i_39038(.S(n_55111), .A(inst_deco2[89]), .B(n_43726), .Z(n_32720
		));
	notech_or2 i_234(.A(n_3055), .B(n_40798), .Z(n_254294499));
	notech_reg inst_deco2_reg_90(.CP(n_62268), .D(n_32726), .CD(n_61720), .Q
		(inst_deco2[90]));
	notech_mux2 i_39046(.S(n_55101), .A(inst_deco2[90]), .B(n_43732), .Z(n_32726
		));
	notech_ao4 i_235(.A(n_40782), .B(n_3052), .C(n_40750), .D(n_3053), .Z(n_254194498
		));
	notech_reg inst_deco2_reg_91(.CP(n_62266), .D(n_32732), .CD(n_61718), .Q
		(inst_deco2[91]));
	notech_mux2 i_39054(.S(n_55101), .A(inst_deco2[91]), .B(n_43738), .Z(n_32732
		));
	notech_and4 i_1047(.A(n_254194498), .B(n_254294499), .C(n_253294489), .D
		(n_3118), .Z(n_254094497));
	notech_reg inst_deco2_reg_92(.CP(n_62266), .D(n_32738), .CD(n_61718), .Q
		(inst_deco2[92]));
	notech_mux2 i_39062(.S(n_55101), .A(inst_deco2[92]), .B(n_43744), .Z(n_32738
		));
	notech_reg inst_deco2_reg_93(.CP(n_62266), .D(n_32744), .CD(n_61720), .Q
		(inst_deco2[93]));
	notech_mux2 i_39070(.S(n_55101), .A(inst_deco2[93]), .B(n_43750), .Z(n_32744
		));
	notech_reg inst_deco2_reg_94(.CP(n_62266), .D(n_32750), .CD(n_61720), .Q
		(inst_deco2[94]));
	notech_mux2 i_39078(.S(n_55101), .A(inst_deco2[94]), .B(n_43756), .Z(n_32750
		));
	notech_reg inst_deco2_reg_95(.CP(n_62266), .D(n_32756), .CD(n_61720), .Q
		(inst_deco2[95]));
	notech_mux2 i_39086(.S(n_55101), .A(inst_deco2[95]), .B(n_43762), .Z(n_32756
		));
	notech_reg inst_deco2_reg_96(.CP(n_62266), .D(n_32762), .CD(n_61720), .Q
		(inst_deco2[96]));
	notech_mux2 i_39094(.S(n_55101), .A(inst_deco2[96]), .B(n_43768), .Z(n_32762
		));
	notech_or2 i_1039(.A(n_3046), .B(n_40774), .Z(n_253594492));
	notech_reg inst_deco2_reg_97(.CP(n_62266), .D(n_32768), .CD(n_61720), .Q
		(inst_deco2[97]));
	notech_mux2 i_39102(.S(n_55106), .A(inst_deco2[97]), .B(n_43774), .Z(n_32768
		));
	notech_reg inst_deco2_reg_98(.CP(n_62266), .D(n_32774), .CD(n_61718), .Q
		(inst_deco2[98]));
	notech_mux2 i_39110(.S(n_55106), .A(inst_deco2[98]), .B(n_43780), .Z(n_32774
		));
	notech_reg inst_deco2_reg_99(.CP(n_62266), .D(n_32780), .CD(n_61718), .Q
		(inst_deco2[99]));
	notech_mux2 i_39118(.S(n_55106), .A(inst_deco2[99]), .B(n_43786), .Z(n_32780
		));
	notech_or2 i_1041(.A(n_3045), .B(n_40766), .Z(n_253294489));
	notech_reg inst_deco2_reg_100(.CP(n_62266), .D(n_32786), .CD(n_61718), .Q
		(inst_deco2[100]));
	notech_mux2 i_39126(.S(n_55101), .A(inst_deco2[100]), .B(n_43792), .Z(n_32786
		));
	notech_or4 i_18374153(.A(n_225196458), .B(n_225096459), .C(n_40490), .D(n_2123
		), .Z(n_253194488));
	notech_reg inst_deco2_reg_101(.CP(n_62266), .D(n_32792), .CD(n_61718), .Q
		(inst_deco2[101]));
	notech_mux2 i_39134(.S(n_55101), .A(inst_deco2[101]), .B(n_43798), .Z(n_32792
		));
	notech_or2 i_231(.A(n_3055), .B(n_40797), .Z(n_253094487));
	notech_reg inst_deco2_reg_102(.CP(n_62268), .D(n_32798), .CD(n_61718), .Q
		(inst_deco2[102]));
	notech_mux2 i_39142(.S(n_55101), .A(inst_deco2[102]), .B(n_43804), .Z(n_32798
		));
	notech_ao4 i_232(.A(n_3052), .B(n_40781), .C(n_3053), .D(n_40749), .Z(n_252994486
		));
	notech_reg inst_deco2_reg_103(.CP(n_62271), .D(n_32804), .CD(n_61718), .Q
		(inst_deco2[103]));
	notech_mux2 i_39150(.S(n_55111), .A(inst_deco2[103]), .B(n_43810), .Z(n_32804
		));
	notech_and4 i_1035(.A(n_252994486), .B(n_253094487), .C(n_252194478), .D
		(n_3113), .Z(n_252894485));
	notech_reg inst_deco2_reg_104(.CP(n_62268), .D(n_32810), .CD(n_61718), .Q
		(inst_deco2[104]));
	notech_mux2 i_39158(.S(n_55112), .A(inst_deco2[104]), .B(n_43816), .Z(n_32810
		));
	notech_reg inst_deco2_reg_105(.CP(n_62268), .D(n_32816), .CD(n_61718), .Q
		(inst_deco2[105]));
	notech_mux2 i_39166(.S(n_55112), .A(inst_deco2[105]), .B(n_43822), .Z(n_32816
		));
	notech_reg inst_deco2_reg_106(.CP(n_62268), .D(n_32822), .CD(n_61718), .Q
		(inst_deco2[106]));
	notech_mux2 i_39174(.S(n_55112), .A(inst_deco2[106]), .B(n_43828), .Z(n_32822
		));
	notech_reg inst_deco2_reg_107(.CP(n_62271), .D(n_32828), .CD(n_61718), .Q
		(inst_deco2[107]));
	notech_mux2 i_39182(.S(n_55112), .A(inst_deco2[107]), .B(n_3306), .Z(n_32828
		));
	notech_or2 i_1027(.A(n_3046), .B(n_40773), .Z(n_252494481));
	notech_reg inst_deco2_reg_108(.CP(n_62271), .D(n_32834), .CD(n_61718), .Q
		(inst_deco2[108]));
	notech_mux2 i_39190(.S(n_55112), .A(inst_deco2[108]), .B(n_43840), .Z(n_32834
		));
	notech_reg inst_deco2_reg_109(.CP(n_62271), .D(n_32840), .CD(n_61723), .Q
		(inst_deco2[109]));
	notech_mux2 i_39198(.S(n_55112), .A(inst_deco2[109]), .B(n_43846), .Z(n_32840
		));
	notech_reg inst_deco2_reg_110(.CP(n_62271), .D(n_32846), .CD(n_61723), .Q
		(inst_deco2[110]));
	notech_mux2 i_39206(.S(n_55112), .A(inst_deco2[110]), .B(n_3302), .Z(n_32846
		));
	notech_or2 i_1029(.A(n_3045), .B(n_40765), .Z(n_252194478));
	notech_reg inst_deco2_reg_111(.CP(n_62271), .D(n_32852), .CD(n_61723), .Q
		(inst_deco2[111]));
	notech_mux2 i_39214(.S(n_55112), .A(inst_deco2[111]), .B(n_43858), .Z(n_32852
		));
	notech_or2 i_224(.A(n_3055), .B(n_40796), .Z(n_252094477));
	notech_reg inst_deco2_reg_112(.CP(n_62268), .D(n_32858), .CD(n_61720), .Q
		(inst_deco2[112]));
	notech_mux2 i_39222(.S(n_55112), .A(inst_deco2[112]), .B(n_43864), .Z(n_32858
		));
	notech_ao4 i_229(.A(n_3052), .B(n_40780), .C(n_3053), .D(n_40748), .Z(n_251994476
		));
	notech_reg inst_deco2_reg_113(.CP(n_62268), .D(n_32864), .CD(n_61723), .Q
		(inst_deco2[113]));
	notech_mux2 i_39230(.S(n_55112), .A(inst_deco2[113]), .B(n_43870), .Z(n_32864
		));
	notech_and4 i_1023(.A(n_251994476), .B(n_252094477), .C(n_251194468), .D
		(n_3108), .Z(n_251894475));
	notech_reg inst_deco2_reg_114(.CP(n_62268), .D(n_32870), .CD(n_61723), .Q
		(inst_deco2[114]));
	notech_mux2 i_39238(.S(n_55112), .A(inst_deco2[114]), .B(n_43876), .Z(n_32870
		));
	notech_reg inst_deco2_reg_115(.CP(n_62268), .D(n_32876), .CD(n_61723), .Q
		(inst_deco2[115]));
	notech_mux2 i_39246(.S(n_55112), .A(inst_deco2[115]), .B(n_43882), .Z(n_32876
		));
	notech_reg inst_deco2_reg_116(.CP(n_62268), .D(n_32882), .CD(n_61723), .Q
		(inst_deco2[116]));
	notech_mux2 i_39254(.S(n_55112), .A(inst_deco2[116]), .B(n_43888), .Z(n_32882
		));
	notech_reg inst_deco2_reg_117(.CP(n_62268), .D(n_32888), .CD(n_61723), .Q
		(inst_deco2[117]));
	notech_mux2 i_39262(.S(n_55111), .A(inst_deco2[117]), .B(n_43894), .Z(n_32888
		));
	notech_or2 i_1015(.A(n_3046), .B(n_40772), .Z(n_251494471));
	notech_reg inst_deco2_reg_118(.CP(n_62268), .D(n_32894), .CD(n_61723), .Q
		(inst_deco2[118]));
	notech_mux2 i_39270(.S(n_55111), .A(inst_deco2[118]), .B(n_43900), .Z(n_32894
		));
	notech_reg inst_deco2_reg_119(.CP(n_62268), .D(n_32900), .CD(n_61720), .Q
		(inst_deco2[119]));
	notech_mux2 i_39278(.S(n_55111), .A(inst_deco2[119]), .B(n_43906), .Z(n_32900
		));
	notech_reg inst_deco2_reg_120(.CP(n_62268), .D(n_32906), .CD(n_61720), .Q
		(inst_deco2[120]));
	notech_mux2 i_39286(.S(n_55111), .A(inst_deco2[120]), .B(n_43912), .Z(n_32906
		));
	notech_or2 i_1017(.A(n_3045), .B(n_40764), .Z(n_251194468));
	notech_reg inst_deco2_reg_121(.CP(n_62268), .D(n_32912), .CD(n_61720), .Q
		(inst_deco2[121]));
	notech_mux2 i_39294(.S(n_55111), .A(inst_deco2[121]), .B(n_43918), .Z(n_32912
		));
	notech_or2 i_220(.A(n_3055), .B(n_40795), .Z(n_251094467));
	notech_reg inst_deco2_reg_122(.CP(n_62268), .D(n_32918), .CD(n_61720), .Q
		(inst_deco2[122]));
	notech_mux2 i_39302(.S(n_55111), .A(inst_deco2[122]), .B(n_43924), .Z(n_32918
		));
	notech_ao4 i_221(.A(n_3052), .B(n_40779), .C(n_3053), .D(n_40747), .Z(n_250994466
		));
	notech_reg inst_deco2_reg_123(.CP(n_62299), .D(n_32924), .CD(n_61720), .Q
		(inst_deco2[123]));
	notech_mux2 i_39310(.S(n_55111), .A(inst_deco2[123]), .B(n_43930), .Z(n_32924
		));
	notech_and4 i_1011(.A(n_250994466), .B(n_251094467), .C(n_250194458), .D
		(n_3103), .Z(n_250894465));
	notech_reg inst_deco2_reg_124(.CP(n_62331), .D(n_32930), .CD(n_61720), .Q
		(inst_deco2[124]));
	notech_mux2 i_39318(.S(n_55111), .A(inst_deco2[124]), .B(n_43936), .Z(n_32930
		));
	notech_reg inst_deco2_reg_125(.CP(n_62331), .D(n_32936), .CD(n_61720), .Q
		(inst_deco2[125]));
	notech_mux2 i_39326(.S(n_55111), .A(inst_deco2[125]), .B(n_43942), .Z(n_32936
		));
	notech_reg inst_deco2_reg_126(.CP(n_62331), .D(n_32942), .CD(n_61720), .Q
		(inst_deco2[126]));
	notech_mux2 i_39334(.S(n_55111), .A(inst_deco2[126]), .B(n_43948), .Z(n_32942
		));
	notech_reg inst_deco2_reg_127(.CP(n_62331), .D(n_32948), .CD(n_61720), .Q
		(inst_deco2[127]));
	notech_mux2 i_39342(.S(n_55111), .A(inst_deco2[127]), .B(n_43954), .Z(n_32948
		));
	notech_or2 i_1003(.A(n_3046), .B(n_40771), .Z(n_250494461));
	notech_reg inst_deco1_reg_0(.CP(n_62331), .D(n_32954), .CD(n_61720), .Q(inst_deco1
		[0]));
	notech_mux2 i_39350(.S(n_58326), .A(inst_deco1[0]), .B(n_39775), .Z(n_32954
		));
	notech_reg inst_deco1_reg_1(.CP(n_62331), .D(n_32960), .CD(n_61720), .Q(inst_deco1
		[1]));
	notech_mux2 i_39358(.S(n_58326), .A(inst_deco1[1]), .B(n_39777), .Z(n_32960
		));
	notech_reg inst_deco1_reg_2(.CP(n_62331), .D(n_32966), .CD(n_61783), .Q(inst_deco1
		[2]));
	notech_mux2 i_39366(.S(n_58304), .A(inst_deco1[2]), .B(n_39778), .Z(n_32966
		));
	notech_or2 i_1005(.A(n_3045), .B(n_40763), .Z(n_250194458));
	notech_reg inst_deco1_reg_3(.CP(n_62331), .D(n_32972), .CD(n_61783), .Q(inst_deco1
		[3]));
	notech_mux2 i_39374(.S(n_58304), .A(inst_deco1[3]), .B(n_39779), .Z(n_32972
		));
	notech_or2 i_215(.A(n_3055), .B(n_40794), .Z(n_250094457));
	notech_reg inst_deco1_reg_4(.CP(n_62331), .D(n_32978), .CD(n_61783), .Q(inst_deco1
		[4]));
	notech_mux2 i_39382(.S(n_58304), .A(inst_deco1[4]), .B(n_39780), .Z(n_32978
		));
	notech_ao4 i_217(.A(n_3052), .B(n_40778), .C(n_3053), .D(n_40746), .Z(n_249994456
		));
	notech_reg inst_deco1_reg_5(.CP(n_62331), .D(n_32984), .CD(n_61783), .Q(inst_deco1
		[5]));
	notech_mux2 i_39390(.S(n_58304), .A(inst_deco1[5]), .B(n_39781), .Z(n_32984
		));
	notech_and4 i_999(.A(n_249994456), .B(n_250094457), .C(n_249194448), .D(n_3098
		), .Z(n_249894455));
	notech_reg inst_deco1_reg_6(.CP(n_62331), .D(n_32990), .CD(n_61783), .Q(inst_deco1
		[6]));
	notech_mux2 i_39398(.S(n_58304), .A(inst_deco1[6]), .B(n_39782), .Z(n_32990
		));
	notech_reg inst_deco1_reg_7(.CP(n_62327), .D(n_32996), .CD(n_61784), .Q(inst_deco1
		[7]));
	notech_mux2 i_39406(.S(n_58304), .A(inst_deco1[7]), .B(n_39783), .Z(n_32996
		));
	notech_reg inst_deco1_reg_8(.CP(n_62327), .D(n_33002), .CD(n_61784), .Q(inst_deco1
		[8]));
	notech_mux2 i_39414(.S(n_58304), .A(inst_deco1[8]), .B(n_39784), .Z(n_33002
		));
	notech_reg inst_deco1_reg_9(.CP(n_62327), .D(n_33008), .CD(n_61784), .Q(inst_deco1
		[9]));
	notech_mux2 i_39422(.S(n_58309), .A(inst_deco1[9]), .B(n_39785), .Z(n_33008
		));
	notech_or2 i_991(.A(n_3046), .B(n_40770), .Z(n_249494451));
	notech_reg inst_deco1_reg_10(.CP(n_62327), .D(n_33014), .CD(n_61784), .Q
		(inst_deco1[10]));
	notech_mux2 i_39430(.S(n_58309), .A(inst_deco1[10]), .B(n_39787), .Z(n_33014
		));
	notech_reg inst_deco1_reg_11(.CP(n_62327), .D(n_33020), .CD(n_61784), .Q
		(inst_deco1[11]));
	notech_mux2 i_39438(.S(n_58309), .A(inst_deco1[11]), .B(n_39789), .Z(n_33020
		));
	notech_reg inst_deco1_reg_12(.CP(n_62331), .D(n_33026), .CD(n_61783), .Q
		(inst_deco1[12]));
	notech_mux2 i_39446(.S(n_58304), .A(inst_deco1[12]), .B(n_39791), .Z(n_33026
		));
	notech_or2 i_993(.A(n_3045), .B(n_40762), .Z(n_249194448));
	notech_reg inst_deco1_reg_13(.CP(n_62331), .D(n_33032), .CD(n_61779), .Q
		(inst_deco1[13]));
	notech_mux2 i_39454(.S(n_58309), .A(inst_deco1[13]), .B(n_39792), .Z(n_33032
		));
	notech_or2 i_210(.A(n_3055), .B(n_40793), .Z(n_249094447));
	notech_reg inst_deco1_reg_14(.CP(n_62331), .D(n_33038), .CD(n_61779), .Q
		(inst_deco1[14]));
	notech_mux2 i_39462(.S(n_58309), .A(inst_deco1[14]), .B(n_39794), .Z(n_33038
		));
	notech_ao4 i_211(.A(n_3052), .B(n_40777), .C(n_3053), .D(n_40745), .Z(n_248994446
		));
	notech_reg inst_deco1_reg_15(.CP(n_62327), .D(n_33044), .CD(n_61779), .Q
		(inst_deco1[15]));
	notech_mux2 i_39470(.S(n_58304), .A(inst_deco1[15]), .B(n_39796), .Z(n_33044
		));
	notech_and4 i_987(.A(n_248994446), .B(n_249094447), .C(n_248194438), .D(n_3093
		), .Z(n_248894445));
	notech_reg inst_deco1_reg_16(.CP(n_62327), .D(n_33050), .CD(n_61779), .Q
		(inst_deco1[16]));
	notech_mux2 i_39478(.S(n_58304), .A(inst_deco1[16]), .B(n_39798), .Z(n_33050
		));
	notech_reg inst_deco1_reg_17(.CP(n_62333), .D(n_33056), .CD(n_61779), .Q
		(inst_deco1[17]));
	notech_mux2 i_39486(.S(n_58304), .A(inst_deco1[17]), .B(n_39800), .Z(n_33056
		));
	notech_reg inst_deco1_reg_18(.CP(n_62333), .D(n_33062), .CD(n_61783), .Q
		(inst_deco1[18]));
	notech_mux2 i_39494(.S(n_58303), .A(inst_deco1[18]), .B(n_39651), .Z(n_33062
		));
	notech_reg inst_deco1_reg_19(.CP(n_62333), .D(n_33068), .CD(n_61783), .Q
		(inst_deco1[19]));
	notech_mux2 i_39502(.S(n_58303), .A(inst_deco1[19]), .B(n_39802), .Z(n_33068
		));
	notech_or2 i_979(.A(n_3046), .B(n_40769), .Z(n_248494441));
	notech_reg inst_deco1_reg_20(.CP(n_62333), .D(n_33074), .CD(n_61783), .Q
		(inst_deco1[20]));
	notech_mux2 i_39510(.S(n_58303), .A(inst_deco1[20]), .B(n_39804), .Z(n_33074
		));
	notech_reg inst_deco1_reg_21(.CP(n_62333), .D(n_33080), .CD(n_61779), .Q
		(inst_deco1[21]));
	notech_mux2 i_39518(.S(n_58304), .A(inst_deco1[21]), .B(n_39806), .Z(n_33080
		));
	notech_reg inst_deco1_reg_22(.CP(n_62333), .D(n_33086), .CD(n_61783), .Q
		(inst_deco1[22]));
	notech_mux2 i_39526(.S(n_58304), .A(inst_deco1[22]), .B(n_39659), .Z(n_33086
		));
	notech_or2 i_981(.A(n_3045), .B(n_40761), .Z(n_248194438));
	notech_reg inst_deco1_reg_23(.CP(n_62333), .D(n_33092), .CD(n_61784), .Q
		(inst_deco1[23]));
	notech_mux2 i_39534(.S(n_58304), .A(inst_deco1[23]), .B(n_39662), .Z(n_33092
		));
	notech_or2 i_201(.A(n_3055), .B(n_40791), .Z(n_248094437));
	notech_reg inst_deco1_reg_24(.CP(n_62333), .D(n_33098), .CD(n_61788), .Q
		(inst_deco1[24]));
	notech_mux2 i_39542(.S(n_58304), .A(inst_deco1[24]), .B(n_39664), .Z(n_33098
		));
	notech_ao4 i_204(.A(n_3052), .B(n_40775), .C(n_3053), .D(n_40743), .Z(n_247994436
		));
	notech_reg inst_deco1_reg_25(.CP(n_62333), .D(n_33104), .CD(n_61784), .Q
		(inst_deco1[25]));
	notech_mux2 i_39550(.S(n_58304), .A(inst_deco1[25]), .B(n_39667), .Z(n_33104
		));
	notech_and4 i_975(.A(n_247994436), .B(n_248094437), .C(n_247194428), .D(n_3088
		), .Z(n_247894435));
	notech_reg inst_deco1_reg_26(.CP(n_62333), .D(n_33110), .CD(n_61784), .Q
		(inst_deco1[26]));
	notech_mux2 i_39558(.S(n_58304), .A(inst_deco1[26]), .B(n_39808), .Z(n_33110
		));
	notech_reg inst_deco1_reg_27(.CP(n_62333), .D(n_33116), .CD(n_61784), .Q
		(inst_deco1[27]));
	notech_mux2 i_39566(.S(n_58304), .A(inst_deco1[27]), .B(n_39810), .Z(n_33116
		));
	notech_reg inst_deco1_reg_28(.CP(n_62331), .D(n_33122), .CD(n_61788), .Q
		(inst_deco1[28]));
	notech_mux2 i_39574(.S(n_58309), .A(inst_deco1[28]), .B(n_39812), .Z(n_33122
		));
	notech_reg inst_deco1_reg_29(.CP(n_62331), .D(n_33128), .CD(n_61788), .Q
		(inst_deco1[29]));
	notech_mux2 i_39582(.S(n_58314), .A(inst_deco1[29]), .B(n_39814), .Z(n_33128
		));
	notech_or2 i_967(.A(n_3046), .B(n_40767), .Z(n_247494431));
	notech_reg inst_deco1_reg_30(.CP(n_62331), .D(n_33134), .CD(n_61788), .Q
		(inst_deco1[30]));
	notech_mux2 i_39590(.S(n_58314), .A(inst_deco1[30]), .B(n_39816), .Z(n_33134
		));
	notech_reg inst_deco1_reg_31(.CP(n_62331), .D(n_33140), .CD(n_61788), .Q
		(inst_deco1[31]));
	notech_mux2 i_39598(.S(n_58314), .A(inst_deco1[31]), .B(n_39818), .Z(n_33140
		));
	notech_reg inst_deco1_reg_32(.CP(n_62331), .D(n_33146), .CD(n_61788), .Q
		(inst_deco1[32]));
	notech_mux2 i_39606(.S(n_58314), .A(inst_deco1[32]), .B(n_39681), .Z(n_33146
		));
	notech_or2 i_969(.A(n_3045), .B(n_40759), .Z(n_247194428));
	notech_reg inst_deco1_reg_33(.CP(n_62333), .D(n_33152), .CD(n_61784), .Q
		(inst_deco1[33]));
	notech_mux2 i_39614(.S(n_58314), .A(inst_deco1[33]), .B(n_39820), .Z(n_33152
		));
	notech_or2 i_197(.A(n_3055), .B(n_40790), .Z(n_247094427));
	notech_reg inst_deco1_reg_34(.CP(n_62333), .D(n_33158), .CD(n_61784), .Q
		(inst_deco1[34]));
	notech_mux2 i_39622(.S(n_58314), .A(inst_deco1[34]), .B(n_39821), .Z(n_33158
		));
	notech_ao4 i_198(.A(n_3053), .B(n_40742), .C(n_3052), .D(n_40774), .Z(n_246994426
		));
	notech_reg inst_deco1_reg_35(.CP(n_62333), .D(n_33164), .CD(n_61784), .Q
		(inst_deco1[35]));
	notech_mux2 i_39630(.S(n_58314), .A(inst_deco1[35]), .B(n_39823), .Z(n_33164
		));
	notech_and4 i_963(.A(n_246994426), .B(n_247094427), .C(n_246194418), .D(n_3083
		), .Z(n_246894425));
	notech_reg inst_deco1_reg_36(.CP(n_62331), .D(n_33170), .CD(n_61784), .Q
		(inst_deco1[36]));
	notech_mux2 i_39638(.S(n_58314), .A(inst_deco1[36]), .B(n_39825), .Z(n_33170
		));
	notech_reg inst_deco1_reg_37(.CP(n_62333), .D(n_33176), .CD(n_61784), .Q
		(inst_deco1[37]));
	notech_mux2 i_39646(.S(n_58315), .A(inst_deco1[37]), .B(n_39692), .Z(n_33176
		));
	notech_reg inst_deco1_reg_38(.CP(n_62327), .D(n_33182), .CD(n_61784), .Q
		(inst_deco1[38]));
	notech_mux2 i_39654(.S(n_58315), .A(inst_deco1[38]), .B(n_39827), .Z(n_33182
		));
	notech_reg inst_deco1_reg_39(.CP(n_62325), .D(n_33188), .CD(n_61784), .Q
		(inst_deco1[39]));
	notech_mux2 i_39662(.S(n_58314), .A(inst_deco1[39]), .B(n_39829), .Z(n_33188
		));
	notech_or2 i_949(.A(n_3046), .B(n_40766), .Z(n_246494421));
	notech_reg inst_deco1_reg_40(.CP(n_62325), .D(n_33194), .CD(n_61784), .Q
		(inst_deco1[40]));
	notech_mux2 i_39670(.S(n_58314), .A(inst_deco1[40]), .B(n_39831), .Z(n_33194
		));
	notech_reg inst_deco1_reg_41(.CP(n_62325), .D(n_33200), .CD(n_61784), .Q
		(inst_deco1[41]));
	notech_mux2 i_39678(.S(n_58314), .A(inst_deco1[41]), .B(n_39833), .Z(n_33200
		));
	notech_reg inst_deco1_reg_42(.CP(n_62325), .D(n_33206), .CD(n_61784), .Q
		(inst_deco1[42]));
	notech_mux2 i_39686(.S(n_58309), .A(inst_deco1[42]), .B(n_39834), .Z(n_33206
		));
	notech_or2 i_951(.A(n_3045), .B(n_40758), .Z(n_246194418));
	notech_reg inst_deco1_reg_43(.CP(n_62325), .D(n_33212), .CD(n_61784), .Q
		(inst_deco1[43]));
	notech_mux2 i_39694(.S(n_58309), .A(inst_deco1[43]), .B(n_39836), .Z(n_33212
		));
	notech_or2 i_192(.A(n_3055), .B(n_40789), .Z(n_246094417));
	notech_reg inst_deco1_reg_44(.CP(n_62325), .D(n_33218), .CD(n_61777), .Q
		(inst_deco1[44]));
	notech_mux2 i_39702(.S(n_58309), .A(inst_deco1[44]), .B(n_39838), .Z(n_33218
		));
	notech_ao4 i_193(.A(n_3053), .B(n_40741), .C(n_3052), .D(n_40773), .Z(n_245994416
		));
	notech_reg inst_deco1_reg_45(.CP(n_62325), .D(n_33224), .CD(n_61777), .Q
		(inst_deco1[45]));
	notech_mux2 i_39710(.S(n_58309), .A(inst_deco1[45]), .B(n_39840), .Z(n_33224
		));
	notech_and4 i_946(.A(n_245994416), .B(n_246094417), .C(n_245194408), .D(n_3078
		), .Z(n_245894415));
	notech_reg inst_deco1_reg_46(.CP(n_62325), .D(n_33230), .CD(n_61777), .Q
		(inst_deco1[46]));
	notech_mux2 i_39718(.S(n_58309), .A(inst_deco1[46]), .B(n_39842), .Z(n_33230
		));
	notech_reg inst_deco1_reg_47(.CP(n_62325), .D(n_33236), .CD(n_61777), .Q
		(inst_deco1[47]));
	notech_mux2 i_39726(.S(n_58309), .A(inst_deco1[47]), .B(n_39844), .Z(n_33236
		));
	notech_reg inst_deco1_reg_48(.CP(n_62325), .D(n_33242), .CD(n_61777), .Q
		(inst_deco1[48]));
	notech_mux2 i_39734(.S(n_58314), .A(inst_deco1[48]), .B(n_39846), .Z(n_33242
		));
	notech_reg inst_deco1_reg_49(.CP(n_62325), .D(n_33248), .CD(n_61777), .Q
		(inst_deco1[49]));
	notech_mux2 i_39742(.S(n_58314), .A(inst_deco1[49]), .B(n_39848), .Z(n_33248
		));
	notech_or2 i_937(.A(n_3046), .B(n_40765), .Z(n_245494411));
	notech_reg inst_deco1_reg_50(.CP(n_62322), .D(n_33254), .CD(n_61777), .Q
		(inst_deco1[50]));
	notech_mux2 i_39750(.S(n_58314), .A(inst_deco1[50]), .B(n_39850), .Z(n_33254
		));
	notech_reg inst_deco1_reg_51(.CP(n_62322), .D(n_33260), .CD(n_61777), .Q
		(inst_deco1[51]));
	notech_mux2 i_39758(.S(n_58314), .A(inst_deco1[51]), .B(n_39852), .Z(n_33260
		));
	notech_reg inst_deco1_reg_52(.CP(n_62322), .D(n_33266), .CD(n_61777), .Q
		(inst_deco1[52]));
	notech_mux2 i_39766(.S(n_58314), .A(inst_deco1[52]), .B(n_39854), .Z(n_33266
		));
	notech_or2 i_939(.A(n_3045), .B(n_40757), .Z(n_245194408));
	notech_reg inst_deco1_reg_53(.CP(n_62322), .D(n_33272), .CD(n_61777), .Q
		(inst_deco1[53]));
	notech_mux2 i_39774(.S(n_58314), .A(inst_deco1[53]), .B(n_39856), .Z(n_33272
		));
	notech_or2 i_187(.A(n_3055), .B(n_40788), .Z(n_245094407));
	notech_reg inst_deco1_reg_54(.CP(n_62322), .D(n_33278), .CD(n_61777), .Q
		(inst_deco1[54]));
	notech_mux2 i_39782(.S(n_58314), .A(inst_deco1[54]), .B(n_39858), .Z(n_33278
		));
	notech_ao4 i_188(.A(n_3053), .B(n_40740), .C(n_3052), .D(n_40772), .Z(n_244994406
		));
	notech_reg inst_deco1_reg_55(.CP(n_62322), .D(n_33284), .CD(n_61774), .Q
		(inst_deco1[55]));
	notech_mux2 i_39790(.S(n_58327), .A(inst_deco1[55]), .B(n_39860), .Z(n_33284
		));
	notech_and4 i_934(.A(n_244994406), .B(n_245094407), .C(n_244194398), .D(n_3073
		), .Z(n_244894405));
	notech_reg inst_deco1_reg_56(.CP(n_62322), .D(n_33290), .CD(n_61774), .Q
		(inst_deco1[56]));
	notech_mux2 i_39798(.S(n_58343), .A(inst_deco1[56]), .B(n_39863), .Z(n_33290
		));
	notech_reg inst_deco1_reg_57(.CP(n_62322), .D(n_33296), .CD(n_61774), .Q
		(inst_deco1[57]));
	notech_mux2 i_39806(.S(n_58348), .A(inst_deco1[57]), .B(n_39866), .Z(n_33296
		));
	notech_reg inst_deco1_reg_58(.CP(n_62322), .D(n_33302), .CD(n_61774), .Q
		(inst_deco1[58]));
	notech_mux2 i_39814(.S(n_58348), .A(inst_deco1[58]), .B(n_39869), .Z(n_33302
		));
	notech_reg inst_deco1_reg_59(.CP(n_62322), .D(n_33308), .CD(n_61774), .Q
		(inst_deco1[59]));
	notech_mux2 i_39822(.S(n_58343), .A(inst_deco1[59]), .B(n_39872), .Z(n_33308
		));
	notech_or2 i_925(.A(n_3046), .B(n_40764), .Z(n_244494401));
	notech_reg inst_deco1_reg_60(.CP(n_62327), .D(n_33314), .CD(n_61777), .Q
		(inst_deco1[60]));
	notech_mux2 i_39830(.S(n_58343), .A(inst_deco1[60]), .B(n_39875), .Z(n_33314
		));
	notech_reg inst_deco1_reg_61(.CP(n_62327), .D(n_33320), .CD(n_61777), .Q
		(inst_deco1[61]));
	notech_mux2 i_39838(.S(n_58343), .A(inst_deco1[61]), .B(n_39878), .Z(n_33320
		));
	notech_reg inst_deco1_reg_62(.CP(n_62327), .D(n_33326), .CD(n_61774), .Q
		(inst_deco1[62]));
	notech_mux2 i_39846(.S(n_58348), .A(inst_deco1[62]), .B(n_39881), .Z(n_33326
		));
	notech_or2 i_927(.A(n_3045), .B(n_40756), .Z(n_244194398));
	notech_reg inst_deco1_reg_63(.CP(n_62327), .D(n_33332), .CD(n_61774), .Q
		(inst_deco1[63]));
	notech_mux2 i_39854(.S(n_58348), .A(inst_deco1[63]), .B(n_39884), .Z(n_33332
		));
	notech_or2 i_181(.A(n_3055), .B(n_40787), .Z(n_244094397));
	notech_reg inst_deco1_reg_64(.CP(n_62327), .D(n_33338), .CD(n_61774), .Q
		(inst_deco1[64]));
	notech_mux2 i_39862(.S(n_58348), .A(inst_deco1[64]), .B(n_39887), .Z(n_33338
		));
	notech_ao4 i_183(.A(n_3053), .B(n_40739), .C(n_3052), .D(n_40771), .Z(n_243994396
		));
	notech_reg inst_deco1_reg_65(.CP(n_62327), .D(n_33344), .CD(n_61779), .Q
		(inst_deco1[65]));
	notech_mux2 i_39870(.S(n_58348), .A(inst_deco1[65]), .B(n_39890), .Z(n_33344
		));
	notech_and4 i_922(.A(n_243994396), .B(n_244094397), .C(n_243194388), .D(n_3068
		), .Z(n_243894395));
	notech_reg inst_deco1_reg_66(.CP(n_62327), .D(n_33350), .CD(n_61779), .Q
		(inst_deco1[66]));
	notech_mux2 i_39878(.S(n_58348), .A(inst_deco1[66]), .B(n_39893), .Z(n_33350
		));
	notech_reg inst_deco1_reg_67(.CP(n_62327), .D(n_33356), .CD(n_61779), .Q
		(inst_deco1[67]));
	notech_mux2 i_39886(.S(n_58348), .A(inst_deco1[67]), .B(n_39896), .Z(n_33356
		));
	notech_reg inst_deco1_reg_68(.CP(n_62327), .D(n_33362), .CD(n_61779), .Q
		(inst_deco1[68]));
	notech_mux2 i_39894(.S(n_58348), .A(inst_deco1[68]), .B(n_39899), .Z(n_33362
		));
	notech_reg inst_deco1_reg_69(.CP(n_62327), .D(n_33368), .CD(n_61779), .Q
		(inst_deco1[69]));
	notech_mux2 i_39902(.S(n_58338), .A(inst_deco1[69]), .B(n_39902), .Z(n_33368
		));
	notech_or2 i_913(.A(n_3046), .B(n_40763), .Z(n_243494391));
	notech_reg inst_deco1_reg_70(.CP(n_62327), .D(n_33374), .CD(n_61779), .Q
		(inst_deco1[70]));
	notech_mux2 i_39910(.S(n_58338), .A(inst_deco1[70]), .B(n_39905), .Z(n_33374
		));
	notech_reg inst_deco1_reg_71(.CP(n_62325), .D(n_33380), .CD(n_61779), .Q
		(inst_deco1[71]));
	notech_mux2 i_39918(.S(n_58343), .A(inst_deco1[71]), .B(n_39908), .Z(n_33380
		));
	notech_reg inst_deco1_reg_72(.CP(n_62325), .D(n_33386), .CD(n_61779), .Q
		(inst_deco1[72]));
	notech_mux2 i_39926(.S(n_58338), .A(inst_deco1[72]), .B(n_39911), .Z(n_33386
		));
	notech_or2 i_915(.A(n_3045), .B(n_40755), .Z(n_243194388));
	notech_reg inst_deco1_reg_73(.CP(n_62325), .D(n_33392), .CD(n_61779), .Q
		(inst_deco1[73]));
	notech_mux2 i_39934(.S(n_58338), .A(inst_deco1[73]), .B(n_39914), .Z(n_33392
		));
	notech_or2 i_178(.A(n_3055), .B(n_40786), .Z(n_243094387));
	notech_reg inst_deco1_reg_74(.CP(n_62325), .D(n_33398), .CD(n_61779), .Q
		(inst_deco1[74]));
	notech_mux2 i_39942(.S(n_58338), .A(inst_deco1[74]), .B(n_39917), .Z(n_33398
		));
	notech_ao4 i_179(.A(n_3053), .B(n_40738), .C(n_3052), .D(n_40770), .Z(n_242994386
		));
	notech_reg inst_deco1_reg_75(.CP(n_62325), .D(n_33404), .CD(n_61779), .Q
		(inst_deco1[75]));
	notech_mux2 i_39950(.S(n_58343), .A(inst_deco1[75]), .B(n_39920), .Z(n_33404
		));
	notech_and4 i_910(.A(n_242994386), .B(n_243094387), .C(n_242194378), .D(n_3063
		), .Z(n_242894385));
	notech_reg inst_deco1_reg_76(.CP(n_62325), .D(n_33410), .CD(n_61777), .Q
		(inst_deco1[76]));
	notech_mux2 i_39958(.S(n_58343), .A(inst_deco1[76]), .B(n_39922), .Z(n_33410
		));
	notech_reg inst_deco1_reg_77(.CP(n_62327), .D(n_33416), .CD(n_61777), .Q
		(inst_deco1[77]));
	notech_mux2 i_39966(.S(n_58343), .A(inst_deco1[77]), .B(n_39925), .Z(n_33416
		));
	notech_reg inst_deco1_reg_78(.CP(n_62325), .D(n_33422), .CD(n_61777), .Q
		(inst_deco1[78]));
	notech_mux2 i_39974(.S(n_58343), .A(inst_deco1[78]), .B(n_39928), .Z(n_33422
		));
	notech_reg inst_deco1_reg_79(.CP(n_62325), .D(n_33428), .CD(n_61777), .Q
		(inst_deco1[79]));
	notech_mux2 i_39982(.S(n_58343), .A(inst_deco1[79]), .B(n_39931), .Z(n_33428
		));
	notech_or2 i_901(.A(n_3046), .B(n_40762), .Z(n_242494381));
	notech_reg inst_deco1_reg_80(.CP(n_62325), .D(n_33434), .CD(n_61777), .Q
		(inst_deco1[80]));
	notech_mux2 i_39990(.S(n_58343), .A(inst_deco1[80]), .B(n_39934), .Z(n_33434
		));
	notech_reg inst_deco1_reg_81(.CP(n_62341), .D(n_33440), .CD(n_61779), .Q
		(inst_deco1[81]));
	notech_mux2 i_39998(.S(n_58343), .A(inst_deco1[81]), .B(n_39937), .Z(n_33440
		));
	notech_reg inst_deco1_reg_82(.CP(n_62341), .D(n_33446), .CD(n_61779), .Q
		(inst_deco1[82]));
	notech_mux2 i_40006(.S(n_58348), .A(inst_deco1[82]), .B(n_39940), .Z(n_33446
		));
	notech_or2 i_903(.A(n_3045), .B(n_40754), .Z(n_242194378));
	notech_reg inst_deco1_reg_83(.CP(n_62341), .D(n_33452), .CD(n_61779), .Q
		(inst_deco1[83]));
	notech_mux2 i_40014(.S(n_58349), .A(inst_deco1[83]), .B(n_39943), .Z(n_33452
		));
	notech_or2 i_173(.A(n_3055), .B(n_40785), .Z(n_242094377));
	notech_reg inst_deco1_reg_84(.CP(n_62341), .D(n_33458), .CD(n_61777), .Q
		(inst_deco1[84]));
	notech_mux2 i_40022(.S(n_58349), .A(inst_deco1[84]), .B(n_39946), .Z(n_33458
		));
	notech_ao4 i_174(.A(n_3053), .B(n_40737), .C(n_3052), .D(n_40769), .Z(n_241994376
		));
	notech_reg inst_deco1_reg_85(.CP(n_62341), .D(n_33464), .CD(n_61777), .Q
		(inst_deco1[85]));
	notech_mux2 i_40030(.S(n_58349), .A(inst_deco1[85]), .B(n_39949), .Z(n_33464
		));
	notech_and4 i_898(.A(n_241994376), .B(n_242094377), .C(n_241194368), .D(n_3058
		), .Z(n_241894375));
	notech_reg inst_deco1_reg_86(.CP(n_62341), .D(n_33470), .CD(n_61788), .Q
		(inst_deco1[86]));
	notech_mux2 i_40038(.S(n_58349), .A(inst_deco1[86]), .B(n_39952), .Z(n_33470
		));
	notech_reg inst_deco1_reg_87(.CP(n_62341), .D(n_33476), .CD(n_61794), .Q
		(inst_deco1[87]));
	notech_mux2 i_40046(.S(n_58349), .A(inst_deco1[87]), .B(n_39955), .Z(n_33476
		));
	notech_reg inst_deco1_reg_88(.CP(n_62341), .D(n_33482), .CD(n_61794), .Q
		(inst_deco1[88]));
	notech_mux2 i_40054(.S(n_58349), .A(inst_deco1[88]), .B(n_39958), .Z(n_33482
		));
	notech_reg inst_deco1_reg_89(.CP(n_62341), .D(n_33488), .CD(n_61794), .Q
		(inst_deco1[89]));
	notech_mux2 i_40062(.S(n_58349), .A(inst_deco1[89]), .B(n_39961), .Z(n_33488
		));
	notech_or2 i_889(.A(n_3046), .B(n_40761), .Z(n_241494371));
	notech_reg inst_deco1_reg_90(.CP(n_62341), .D(n_33494), .CD(n_61794), .Q
		(inst_deco1[90]));
	notech_mux2 i_40070(.S(n_58349), .A(inst_deco1[90]), .B(n_39964), .Z(n_33494
		));
	notech_reg inst_deco1_reg_91(.CP(n_62341), .D(n_33500), .CD(n_61794), .Q
		(inst_deco1[91]));
	notech_mux2 i_40078(.S(n_58349), .A(inst_deco1[91]), .B(n_39967), .Z(n_33500
		));
	notech_reg inst_deco1_reg_92(.CP(n_62341), .D(n_33506), .CD(n_61794), .Q
		(inst_deco1[92]));
	notech_mux2 i_40086(.S(n_58349), .A(inst_deco1[92]), .B(n_39970), .Z(n_33506
		));
	notech_or2 i_891(.A(n_3045), .B(n_40753), .Z(n_241194368));
	notech_reg inst_deco1_reg_93(.CP(n_62341), .D(n_33512), .CD(n_61794), .Q
		(inst_deco1[93]));
	notech_mux2 i_40094(.S(n_58349), .A(inst_deco1[93]), .B(n_39973), .Z(n_33512
		));
	notech_or2 i_165(.A(n_3055), .B(n_40784), .Z(n_241094367));
	notech_reg inst_deco1_reg_94(.CP(n_62341), .D(n_33518), .CD(n_61794), .Q
		(inst_deco1[94]));
	notech_mux2 i_40102(.S(n_58349), .A(inst_deco1[94]), .B(n_39976), .Z(n_33518
		));
	notech_ao4 i_170(.A(n_3052), .B(n_40768), .C(n_3053), .D(n_40736), .Z(n_240994366
		));
	notech_reg inst_deco1_reg_95(.CP(n_62338), .D(n_33524), .CD(n_61794), .Q
		(inst_deco1[95]));
	notech_mux2 i_40110(.S(n_58349), .A(inst_deco1[95]), .B(n_39979), .Z(n_33524
		));
	notech_and4 i_886(.A(n_240994366), .B(n_241094367), .C(n_240194358), .D(n_3050
		), .Z(n_240894365));
	notech_reg inst_deco1_reg_96(.CP(n_62338), .D(n_33530), .CD(n_61794), .Q
		(inst_deco1[96]));
	notech_mux2 i_40118(.S(n_58348), .A(inst_deco1[96]), .B(n_39982), .Z(n_33530
		));
	notech_reg inst_deco1_reg_97(.CP(n_62341), .D(n_33536), .CD(n_61793), .Q
		(inst_deco1[97]));
	notech_mux2 i_40126(.S(n_58348), .A(inst_deco1[97]), .B(n_39985), .Z(n_33536
		));
	notech_reg inst_deco1_reg_98(.CP(n_62341), .D(n_33542), .CD(n_61793), .Q
		(inst_deco1[98]));
	notech_mux2 i_40134(.S(n_58348), .A(inst_deco1[98]), .B(n_39989), .Z(n_33542
		));
	notech_reg inst_deco1_reg_99(.CP(n_62341), .D(n_33548), .CD(n_61793), .Q
		(inst_deco1[99]));
	notech_mux2 i_40142(.S(n_58348), .A(inst_deco1[99]), .B(n_39992), .Z(n_33548
		));
	notech_or2 i_877(.A(n_3046), .B(n_40760), .Z(n_240494361));
	notech_reg inst_deco1_reg_100(.CP(n_62341), .D(n_33554), .CD(n_61793), .Q
		(inst_deco1[100]));
	notech_mux2 i_40150(.S(n_58348), .A(inst_deco1[100]), .B(n_39995), .Z(n_33554
		));
	notech_reg inst_deco1_reg_101(.CP(n_62341), .D(n_33560), .CD(n_61793), .Q
		(inst_deco1[101]));
	notech_mux2 i_40158(.S(n_58348), .A(inst_deco1[101]), .B(n_39997), .Z(n_33560
		));
	notech_reg inst_deco1_reg_102(.CP(n_62343), .D(n_33566), .CD(n_61793), .Q
		(inst_deco1[102]));
	notech_mux2 i_40166(.S(n_58348), .A(inst_deco1[102]), .B(n_39999), .Z(n_33566
		));
	notech_or2 i_879(.A(n_3045), .B(n_40752), .Z(n_240194358));
	notech_reg inst_deco1_reg_103(.CP(n_62343), .D(n_33572), .CD(n_61793), .Q
		(inst_deco1[103]));
	notech_mux2 i_40174(.S(n_58349), .A(inst_deco1[103]), .B(n_40001), .Z(n_33572
		));
	notech_and2 i_141(.A(n_239994356), .B(n_2945), .Z(n_240094357));
	notech_reg inst_deco1_reg_104(.CP(n_62343), .D(n_33578), .CD(n_61793), .Q
		(inst_deco1[104]));
	notech_mux2 i_40182(.S(n_58349), .A(inst_deco1[104]), .B(n_40003), .Z(n_33578
		));
	notech_nand3 i_629759(.A(n_40591), .B(n_40592), .C(imm_sz[2]), .Z(n_239994356
		));
	notech_reg inst_deco1_reg_105(.CP(n_62343), .D(n_33584), .CD(n_61793), .Q
		(inst_deco1[105]));
	notech_mux2 i_40190(.S(n_58349), .A(inst_deco1[105]), .B(n_40005), .Z(n_33584
		));
	notech_and2 i_876(.A(n_239994356), .B(n_40534), .Z(n_239894355));
	notech_reg inst_deco1_reg_106(.CP(n_62343), .D(n_33590), .CD(n_61793), .Q
		(inst_deco1[106]));
	notech_mux2 i_40198(.S(n_58348), .A(inst_deco1[106]), .B(n_40007), .Z(n_33590
		));
	notech_or2 i_160(.A(n_2172), .B(n_40774), .Z(n_239794354));
	notech_reg inst_deco1_reg_107(.CP(n_62343), .D(n_33596), .CD(n_61793), .Q
		(inst_deco1[107]));
	notech_mux2 i_40206(.S(n_58349), .A(inst_deco1[107]), .B(n_40009), .Z(n_33596
		));
	notech_reg inst_deco1_reg_108(.CP(n_62343), .D(n_33602), .CD(n_61796), .Q
		(inst_deco1[108]));
	notech_mux2 i_40214(.S(n_58349), .A(inst_deco1[108]), .B(n_40011), .Z(n_33602
		));
	notech_reg inst_deco1_reg_109(.CP(n_62343), .D(n_33608), .CD(n_61796), .Q
		(inst_deco1[109]));
	notech_mux2 i_40222(.S(n_58332), .A(inst_deco1[109]), .B(n_40013), .Z(n_33608
		));
	notech_and4 i_872(.A(n_3042), .B(n_3041), .C(n_3040), .D(n_239794354), .Z
		(n_239494351));
	notech_reg inst_deco1_reg_110(.CP(n_62343), .D(n_33614), .CD(n_61796), .Q
		(inst_deco1[110]));
	notech_mux2 i_40230(.S(n_58332), .A(inst_deco1[110]), .B(n_40015), .Z(n_33614
		));
	notech_reg inst_deco1_reg_111(.CP(n_62343), .D(n_33620), .CD(n_61796), .Q
		(inst_deco1[111]));
	notech_mux2 i_40238(.S(n_58332), .A(inst_deco1[111]), .B(n_40017), .Z(n_33620
		));
	notech_reg inst_deco1_reg_112(.CP(n_62343), .D(n_33626), .CD(n_61796), .Q
		(inst_deco1[112]));
	notech_mux2 i_40246(.S(n_58332), .A(inst_deco1[112]), .B(n_40019), .Z(n_33626
		));
	notech_reg inst_deco1_reg_113(.CP(n_62343), .D(n_33632), .CD(n_61796), .Q
		(inst_deco1[113]));
	notech_mux2 i_40254(.S(n_58332), .A(inst_deco1[113]), .B(n_40021), .Z(n_33632
		));
	notech_reg inst_deco1_reg_114(.CP(n_62343), .D(n_33638), .CD(n_61796), .Q
		(inst_deco1[114]));
	notech_mux2 i_40262(.S(n_58332), .A(inst_deco1[114]), .B(n_40023), .Z(n_33638
		));
	notech_or2 i_4100(.A(n_2149), .B(n_2972), .Z(n_238994346));
	notech_reg inst_deco1_reg_115(.CP(n_62343), .D(n_33644), .CD(n_61796), .Q
		(inst_deco1[115]));
	notech_mux2 i_40270(.S(n_58332), .A(inst_deco1[115]), .B(n_40025), .Z(n_33644
		));
	notech_nao3 i_4102(.A(n_40487), .B(n_2962), .C(n_2149), .Z(n_238894345)
		);
	notech_reg inst_deco1_reg_116(.CP(n_62341), .D(n_33650), .CD(n_61796), .Q
		(inst_deco1[116]));
	notech_mux2 i_40278(.S(n_58337), .A(inst_deco1[116]), .B(n_40027), .Z(n_33650
		));
	notech_or2 i_4103(.A(n_2149), .B(n_2968), .Z(n_238794344));
	notech_reg inst_deco1_reg_117(.CP(n_62343), .D(n_33656), .CD(n_61796), .Q
		(inst_deco1[117]));
	notech_mux2 i_40286(.S(n_58337), .A(inst_deco1[117]), .B(n_40029), .Z(n_33656
		));
	notech_or2 i_18774152(.A(n_40492), .B(n_2127), .Z(n_238694343));
	notech_reg inst_deco1_reg_118(.CP(n_62343), .D(n_33662), .CD(n_61796), .Q
		(inst_deco1[118]));
	notech_mux2 i_40294(.S(n_58337), .A(inst_deco1[118]), .B(n_40032), .Z(n_33662
		));
	notech_or2 i_157(.A(n_2173), .B(n_40748), .Z(n_238594342));
	notech_reg inst_deco1_reg_119(.CP(n_62343), .D(n_33668), .CD(n_61794), .Q
		(inst_deco1[119]));
	notech_mux2 i_40302(.S(n_58332), .A(inst_deco1[119]), .B(n_40034), .Z(n_33668
		));
	notech_reg inst_deco1_reg_120(.CP(n_62343), .D(n_33674), .CD(n_61794), .Q
		(inst_deco1[120]));
	notech_mux2 i_40310(.S(n_58332), .A(inst_deco1[120]), .B(n_40037), .Z(n_33674
		));
	notech_reg inst_deco1_reg_121(.CP(n_62343), .D(n_33680), .CD(n_61794), .Q
		(inst_deco1[121]));
	notech_mux2 i_40318(.S(n_58337), .A(inst_deco1[121]), .B(n_40040), .Z(n_33680
		));
	notech_and4 i_862(.A(n_3037), .B(n_3036), .C(n_3035), .D(n_238594342), .Z
		(n_238294339));
	notech_reg inst_deco1_reg_122(.CP(n_62343), .D(n_33686), .CD(n_61794), .Q
		(inst_deco1[122]));
	notech_mux2 i_40326(.S(n_58327), .A(inst_deco1[122]), .B(n_40043), .Z(n_33686
		));
	notech_reg inst_deco1_reg_123(.CP(n_62338), .D(n_33692), .CD(n_61794), .Q
		(inst_deco1[123]));
	notech_mux2 i_40334(.S(n_58327), .A(inst_deco1[123]), .B(n_40046), .Z(n_33692
		));
	notech_reg inst_deco1_reg_124(.CP(n_62336), .D(n_33698), .CD(n_61794), .Q
		(inst_deco1[124]));
	notech_mux2 i_40342(.S(n_58327), .A(inst_deco1[124]), .B(n_40049), .Z(n_33698
		));
	notech_reg inst_deco1_reg_125(.CP(n_62336), .D(n_33704), .CD(n_61794), .Q
		(inst_deco1[125]));
	notech_mux2 i_40350(.S(n_58327), .A(inst_deco1[125]), .B(n_40052), .Z(n_33704
		));
	notech_reg inst_deco1_reg_126(.CP(n_62336), .D(n_33710), .CD(n_61794), .Q
		(inst_deco1[126]));
	notech_mux2 i_40358(.S(n_58327), .A(inst_deco1[126]), .B(n_40055), .Z(n_33710
		));
	notech_or2 i_142(.A(n_2172), .B(n_40771), .Z(n_237794334));
	notech_reg inst_deco1_reg_127(.CP(n_62336), .D(n_33716), .CD(n_61794), .Q
		(inst_deco1[127]));
	notech_mux2 i_40366(.S(n_58327), .A(inst_deco1[127]), .B(n_39116), .Z(n_33716
		));
	notech_reg to_acu2_reg_0(.CP(n_62336), .D(n_33722), .CD(n_61794), .Q(to_acu2
		[0]));
	notech_mux2 i_40374(.S(n_55111), .A(to_acu2[0]), .B(n_1984), .Z(n_33722)
		);
	notech_reg to_acu2_reg_1(.CP(n_62336), .D(n_33728), .CD(n_61789), .Q(to_acu2
		[1]));
	notech_mux2 i_40382(.S(n_55111), .A(to_acu2[1]), .B(n_1976), .Z(n_33728)
		);
	notech_and4 i_852(.A(n_3032), .B(n_3031), .C(n_3030), .D(n_237794334), .Z
		(n_237494331));
	notech_reg to_acu2_reg_2(.CP(n_62336), .D(n_33734), .CD(n_61789), .Q(to_acu2
		[2]));
	notech_mux2 i_40390(.S(n_55043), .A(to_acu2[2]), .B(n_1980), .Z(n_33734)
		);
	notech_reg to_acu2_reg_3(.CP(n_62336), .D(n_33740), .CD(n_61789), .Q(to_acu2
		[3]));
	notech_mux2 i_40398(.S(n_55043), .A(to_acu2[3]), .B(n_2011), .Z(n_33740)
		);
	notech_reg to_acu2_reg_4(.CP(n_62336), .D(n_33746), .CD(n_61788), .Q(to_acu2
		[4]));
	notech_mux2 i_40406(.S(n_55043), .A(to_acu2[4]), .B(n_2005), .Z(n_33746)
		);
	notech_reg to_acu2_reg_5(.CP(n_62336), .D(n_33752), .CD(n_61788), .Q(to_acu2
		[5]));
	notech_mux2 i_40414(.S(n_55043), .A(to_acu2[5]), .B(n_1960), .Z(n_33752)
		);
	notech_reg to_acu2_reg_6(.CP(n_62336), .D(n_33758), .CD(n_61789), .Q(to_acu2
		[6]));
	notech_mux2 i_40422(.S(n_55043), .A(to_acu2[6]), .B(n_2022), .Z(n_33758)
		);
	notech_or2 i_137(.A(n_2172), .B(n_40770), .Z(n_236994326));
	notech_reg to_acu2_reg_7(.CP(n_62333), .D(n_33764), .CD(n_61789), .Q(to_acu2
		[7]));
	notech_mux2 i_40430(.S(n_55043), .A(to_acu2[7]), .B(n_1957), .Z(n_33764)
		);
	notech_reg to_acu2_reg_8(.CP(n_62333), .D(n_33770), .CD(n_61789), .Q(to_acu2
		[8]));
	notech_mux2 i_40438(.S(n_55044), .A(to_acu2[8]), .B(n_2017), .Z(n_33770)
		);
	notech_reg to_acu2_reg_9(.CP(n_62333), .D(n_33776), .CD(n_61789), .Q(to_acu2
		[9]));
	notech_mux2 i_40446(.S(n_55044), .A(to_acu2[9]), .B(n_1975), .Z(n_33776)
		);
	notech_and4 i_842(.A(n_3027), .B(n_3026), .C(n_3025), .D(n_236994326), .Z
		(n_236694323));
	notech_reg to_acu2_reg_10(.CP(n_62333), .D(n_33782), .CD(n_61789), .Q(to_acu2
		[10]));
	notech_mux2 i_40454(.S(n_55044), .A(to_acu2[10]), .B(n_2018), .Z(n_33782
		));
	notech_reg to_acu2_reg_11(.CP(n_62333), .D(n_33788), .CD(n_61788), .Q(to_acu2
		[11]));
	notech_mux2 i_40462(.S(n_55044), .A(to_acu2[11]), .B(n_3726), .Z(n_33788
		));
	notech_reg to_acu2_reg_12(.CP(n_62336), .D(n_33794), .CD(n_61788), .Q(to_acu2
		[12]));
	notech_mux2 i_40470(.S(n_55044), .A(to_acu2[12]), .B(n_3724), .Z(n_33794
		));
	notech_reg to_acu2_reg_13(.CP(n_62336), .D(n_33800), .CD(n_61788), .Q(to_acu2
		[13]));
	notech_mux2 i_40478(.S(n_55044), .A(to_acu2[13]), .B(n_3722), .Z(n_33800
		));
	notech_reg to_acu2_reg_14(.CP(n_62336), .D(n_33806), .CD(n_61788), .Q(to_acu2
		[14]));
	notech_mux2 i_40486(.S(n_55044), .A(to_acu2[14]), .B(n_3720), .Z(n_33806
		));
	notech_or2 i_133(.A(n_2172), .B(n_40769), .Z(n_236194318));
	notech_reg to_acu2_reg_15(.CP(n_62336), .D(n_33812), .CD(n_61788), .Q(to_acu2
		[15]));
	notech_mux2 i_40494(.S(n_55043), .A(to_acu2[15]), .B(n_3718), .Z(n_33812
		));
	notech_reg to_acu2_reg_16(.CP(n_62336), .D(n_33818), .CD(n_61788), .Q(to_acu2
		[16]));
	notech_mux2 i_40502(.S(n_55043), .A(to_acu2[16]), .B(n_3716), .Z(n_33818
		));
	notech_reg to_acu2_reg_17(.CP(n_62338), .D(n_33824), .CD(n_61788), .Q(to_acu2
		[17]));
	notech_mux2 i_40510(.S(n_55043), .A(to_acu2[17]), .B(n_3714), .Z(n_33824
		));
	notech_and4 i_832(.A(n_3022), .B(n_3021), .C(n_3020), .D(n_236194318), .Z
		(n_235894315));
	notech_reg to_acu2_reg_18(.CP(n_62338), .D(n_33830), .CD(n_61788), .Q(to_acu2
		[18]));
	notech_mux2 i_40518(.S(n_55038), .A(to_acu2[18]), .B(n_3712), .Z(n_33830
		));
	notech_reg to_acu2_reg_19(.CP(n_62338), .D(n_33836), .CD(n_61788), .Q(to_acu2
		[19]));
	notech_mux2 i_40526(.S(n_55043), .A(to_acu2[19]), .B(n_3710), .Z(n_33836
		));
	notech_reg to_acu2_reg_20(.CP(n_62338), .D(n_33842), .CD(n_61788), .Q(to_acu2
		[20]));
	notech_mux2 i_40534(.S(n_55043), .A(to_acu2[20]), .B(n_3708), .Z(n_33842
		));
	notech_reg to_acu2_reg_21(.CP(n_62338), .D(n_33848), .CD(n_61788), .Q(to_acu2
		[21]));
	notech_mux2 i_40542(.S(n_55043), .A(to_acu2[21]), .B(n_3706), .Z(n_33848
		));
	notech_reg to_acu2_reg_22(.CP(n_62338), .D(n_33854), .CD(n_61793), .Q(to_acu2
		[22]));
	notech_mux2 i_40550(.S(n_55043), .A(to_acu2[22]), .B(n_3704), .Z(n_33854
		));
	notech_or4 i_111(.A(n_40479), .B(n_40490), .C(n_1643), .D(n_40736), .Z(n_235394310
		));
	notech_reg to_acu2_reg_23(.CP(n_62338), .D(n_33860), .CD(n_61793), .Q(to_acu2
		[23]));
	notech_mux2 i_40558(.S(n_55043), .A(to_acu2[23]), .B(n_3702), .Z(n_33860
		));
	notech_reg to_acu2_reg_24(.CP(n_62338), .D(n_33866), .CD(n_61793), .Q(to_acu2
		[24]));
	notech_mux2 i_40566(.S(n_55043), .A(to_acu2[24]), .B(n_3700), .Z(n_33866
		));
	notech_reg to_acu2_reg_25(.CP(n_62338), .D(n_33872), .CD(n_61789), .Q(to_acu2
		[25]));
	notech_mux2 i_40574(.S(n_55043), .A(to_acu2[25]), .B(n_3698), .Z(n_33872
		));
	notech_and4 i_822(.A(n_3017), .B(n_3016), .C(n_3015), .D(n_235394310), .Z
		(n_235094307));
	notech_reg to_acu2_reg_26(.CP(n_62338), .D(n_33878), .CD(n_61793), .Q(to_acu2
		[26]));
	notech_mux2 i_40582(.S(n_55043), .A(to_acu2[26]), .B(n_3696), .Z(n_33878
		));
	notech_reg to_acu2_reg_27(.CP(n_62338), .D(n_33884), .CD(n_61793), .Q(to_acu2
		[27]));
	notech_mux2 i_40590(.S(n_55043), .A(to_acu2[27]), .B(n_3694), .Z(n_33884
		));
	notech_reg to_acu2_reg_28(.CP(n_62336), .D(n_33890), .CD(n_61793), .Q(to_acu2
		[28]));
	notech_mux2 i_40598(.S(n_55044), .A(to_acu2[28]), .B(n_3692), .Z(n_33890
		));
	notech_reg to_acu2_reg_29(.CP(n_62338), .D(n_33896), .CD(n_61793), .Q(to_acu2
		[29]));
	notech_mux2 i_40606(.S(n_55027), .A(to_acu2[29]), .B(n_3690), .Z(n_33896
		));
	notech_reg to_acu2_reg_30(.CP(n_62336), .D(n_33902), .CD(n_61793), .Q(to_acu2
		[30]));
	notech_mux2 i_40614(.S(n_55027), .A(to_acu2[30]), .B(n_3688), .Z(n_33902
		));
	notech_or2 i_87(.A(n_2172), .B(n_40767), .Z(n_234594302));
	notech_reg to_acu2_reg_31(.CP(n_62336), .D(n_33908), .CD(n_61793), .Q(to_acu2
		[31]));
	notech_mux2 i_40622(.S(n_55027), .A(to_acu2[31]), .B(n_3686), .Z(n_33908
		));
	notech_reg to_acu2_reg_32(.CP(n_62336), .D(n_33914), .CD(n_61789), .Q(to_acu2
		[32]));
	notech_mux2 i_40630(.S(n_55027), .A(to_acu2[32]), .B(n_3684), .Z(n_33914
		));
	notech_reg to_acu2_reg_33(.CP(n_62338), .D(n_33920), .CD(n_61789), .Q(to_acu2
		[33]));
	notech_mux2 i_40638(.S(n_55027), .A(to_acu2[33]), .B(n_3682), .Z(n_33920
		));
	notech_and4 i_812(.A(n_3012), .B(n_3011), .C(n_3010), .D(n_234594302), .Z
		(n_234294299));
	notech_reg to_acu2_reg_34(.CP(n_62338), .D(n_33926), .CD(n_61789), .Q(to_acu2
		[34]));
	notech_mux2 i_40646(.S(n_55027), .A(to_acu2[34]), .B(n_3680), .Z(n_33926
		));
	notech_reg to_acu2_reg_35(.CP(n_62338), .D(n_33932), .CD(n_61789), .Q(to_acu2
		[35]));
	notech_mux2 i_40654(.S(n_55027), .A(to_acu2[35]), .B(n_3678), .Z(n_33932
		));
	notech_reg to_acu2_reg_36(.CP(n_62338), .D(n_33938), .CD(n_61789), .Q(to_acu2
		[36]));
	notech_mux2 i_40662(.S(n_55054), .A(to_acu2[36]), .B(n_3676), .Z(n_33938
		));
	notech_reg to_acu2_reg_37(.CP(n_62338), .D(n_33944), .CD(n_61789), .Q(to_acu2
		[37]));
	notech_mux2 i_40670(.S(n_55054), .A(to_acu2[37]), .B(n_3674), .Z(n_33944
		));
	notech_reg to_acu2_reg_38(.CP(n_62306), .D(n_33950), .CD(n_61789), .Q(to_acu2
		[38]));
	notech_mux2 i_40678(.S(n_55054), .A(to_acu2[38]), .B(n_3672), .Z(n_33950
		));
	notech_or4 i_85(.A(n_225196458), .B(n_225096459), .C(n_40490), .D(n_40734
		), .Z(n_233794294));
	notech_reg to_acu2_reg_39(.CP(n_62306), .D(n_33960), .CD(n_61789), .Q(to_acu2
		[39]));
	notech_ao3 i_40690(.A(to_acu2[39]), .B(1'b1), .C(n_55027), .Z(n_33960)
		);
	notech_reg to_acu2_reg_40(.CP(n_62306), .D(n_33962), .CD(n_61789), .Q(to_acu2
		[40]));
	notech_mux2 i_40694(.S(n_55027), .A(to_acu2[40]), .B(n_3670), .Z(n_33962
		));
	notech_reg to_acu2_reg_41(.CP(n_62306), .D(n_33968), .CD(n_61789), .Q(to_acu2
		[41]));
	notech_mux2 i_40702(.S(n_55054), .A(to_acu2[41]), .B(n_3668), .Z(n_33968
		));
	notech_and4 i_802(.A(n_3008), .B(n_233794294), .C(n_233094287), .D(n_3006
		), .Z(n_233494291));
	notech_reg to_acu2_reg_42(.CP(n_62306), .D(n_33974), .CD(n_61789), .Q(to_acu2
		[42]));
	notech_mux2 i_40710(.S(n_55044), .A(to_acu2[42]), .B(n_3666), .Z(n_33974
		));
	notech_or4 i_796(.A(n_40479), .B(n_2961), .C(n_40487), .D(n_40742), .Z(n_233394290
		));
	notech_reg to_acu2_reg_43(.CP(n_62309), .D(n_33980), .CD(n_61774), .Q(to_acu2
		[43]));
	notech_mux2 i_40718(.S(n_55044), .A(to_acu2[43]), .B(n_3664), .Z(n_33980
		));
	notech_reg to_acu2_reg_44(.CP(n_62309), .D(n_33986), .CD(n_61758), .Q(to_acu2
		[44]));
	notech_mux2 i_40726(.S(n_55044), .A(to_acu2[44]), .B(n_3662), .Z(n_33986
		));
	notech_reg to_acu2_reg_45(.CP(n_62309), .D(n_33992), .CD(n_61758), .Q(to_acu2
		[45]));
	notech_mux2 i_40734(.S(n_55044), .A(to_acu2[45]), .B(n_3660), .Z(n_33992
		));
	notech_nand3 i_797(.A(n_40487), .B(n_2962), .C(in128[39]), .Z(n_233094287
		));
	notech_reg to_acu2_reg_46(.CP(n_62306), .D(n_33998), .CD(n_61758), .Q(to_acu2
		[46]));
	notech_mux2 i_40742(.S(n_55044), .A(to_acu2[46]), .B(n_3658), .Z(n_33998
		));
	notech_or4 i_66(.A(n_225196458), .B(n_225096459), .C(n_40490), .D(n_40733
		), .Z(n_232994286));
	notech_reg to_acu2_reg_47(.CP(n_62309), .D(n_34004), .CD(n_61758), .Q(to_acu2
		[47]));
	notech_mux2 i_40750(.S(n_55044), .A(to_acu2[47]), .B(n_3656), .Z(n_34004
		));
	notech_reg to_acu2_reg_48(.CP(n_62306), .D(n_34010), .CD(n_61758), .Q(to_acu2
		[48]));
	notech_mux2 i_40758(.S(n_55044), .A(to_acu2[48]), .B(n_3654), .Z(n_34010
		));
	notech_reg to_acu2_reg_49(.CP(n_62306), .D(n_34016), .CD(n_61761), .Q(to_acu2
		[49]));
	notech_mux2 i_40766(.S(n_55027), .A(to_acu2[49]), .B(n_3652), .Z(n_34016
		));
	notech_and4 i_792(.A(n_3003), .B(n_232994286), .C(n_232294279), .D(n_3001
		), .Z(n_232694283));
	notech_reg to_acu2_reg_50(.CP(n_62306), .D(n_34022), .CD(n_61761), .Q(to_acu2
		[50]));
	notech_mux2 i_40774(.S(n_55027), .A(to_acu2[50]), .B(n_3650), .Z(n_34022
		));
	notech_or4 i_786(.A(n_40479), .B(n_2961), .C(n_40487), .D(n_40741), .Z(n_232594282
		));
	notech_reg to_acu2_reg_51(.CP(n_62306), .D(n_34028), .CD(n_61761), .Q(to_acu2
		[51]));
	notech_mux2 i_40782(.S(n_55027), .A(to_acu2[51]), .B(n_3648), .Z(n_34028
		));
	notech_reg to_acu2_reg_52(.CP(n_62306), .D(n_34034), .CD(n_61761), .Q(to_acu2
		[52]));
	notech_mux2 i_40790(.S(n_55044), .A(to_acu2[52]), .B(n_3646), .Z(n_34034
		));
	notech_reg to_acu2_reg_53(.CP(n_62306), .D(n_34040), .CD(n_61761), .Q(to_acu2
		[53]));
	notech_mux2 i_40798(.S(n_55044), .A(to_acu2[53]), .B(n_3644), .Z(n_34040
		));
	notech_nand3 i_787(.A(n_40487), .B(n_2962), .C(in128[38]), .Z(n_232294279
		));
	notech_reg to_acu2_reg_54(.CP(n_62306), .D(n_34046), .CD(n_61758), .Q(to_acu2
		[54]));
	notech_mux2 i_40806(.S(n_55044), .A(to_acu2[54]), .B(n_3642), .Z(n_34046
		));
	notech_or4 i_63(.A(n_225196458), .B(n_225096459), .C(n_40490), .D(n_40732
		), .Z(n_232194278));
	notech_reg to_acu2_reg_55(.CP(n_62306), .D(n_34052), .CD(n_61758), .Q(to_acu2
		[55]));
	notech_mux2 i_40814(.S(n_55032), .A(to_acu2[55]), .B(n_3640), .Z(n_34052
		));
	notech_reg to_acu2_reg_56(.CP(n_62306), .D(n_34058), .CD(n_61758), .Q(to_acu2
		[56]));
	notech_mux2 i_40822(.S(n_55032), .A(to_acu2[56]), .B(n_3638), .Z(n_34058
		));
	notech_reg to_acu2_reg_57(.CP(n_62306), .D(n_34064), .CD(n_61758), .Q(to_acu2
		[57]));
	notech_mux2 i_40830(.S(n_55032), .A(to_acu2[57]), .B(n_3636), .Z(n_34064
		));
	notech_and4 i_782(.A(n_2998), .B(n_232194278), .C(n_231494271), .D(n_2996
		), .Z(n_231894275));
	notech_reg to_acu2_reg_58(.CP(n_62306), .D(n_34070), .CD(n_61758), .Q(to_acu2
		[58]));
	notech_mux2 i_40838(.S(n_55032), .A(to_acu2[58]), .B(n_1958), .Z(n_34070
		));
	notech_or4 i_776(.A(n_40479), .B(n_2961), .C(n_40487), .D(n_40740), .Z(n_231794274
		));
	notech_reg to_acu2_reg_59(.CP(n_62309), .D(n_34076), .CD(n_61758), .Q(to_acu2
		[59]));
	notech_mux2 i_40846(.S(n_55032), .A(to_acu2[59]), .B(n_3633), .Z(n_34076
		));
	notech_reg to_acu2_reg_60(.CP(n_62309), .D(n_34082), .CD(n_61758), .Q(to_acu2
		[60]));
	notech_mux2 i_40854(.S(n_55032), .A(to_acu2[60]), .B(n_3631), .Z(n_34082
		));
	notech_reg to_acu2_reg_61(.CP(n_62309), .D(n_34088), .CD(n_61758), .Q(to_acu2
		[61]));
	notech_mux2 i_40862(.S(n_55032), .A(to_acu2[61]), .B(n_3629), .Z(n_34088
		));
	notech_nand3 i_777(.A(n_40487), .B(n_2962), .C(in128[37]), .Z(n_231494271
		));
	notech_reg to_acu2_reg_62(.CP(n_62309), .D(n_34094), .CD(n_61758), .Q(to_acu2
		[62]));
	notech_mux2 i_40870(.S(n_55032), .A(to_acu2[62]), .B(n_3627), .Z(n_34094
		));
	notech_or4 i_60(.A(n_225196458), .B(n_225096459), .C(n_40490), .D(n_40731
		), .Z(n_231394270));
	notech_reg to_acu2_reg_63(.CP(n_62309), .D(n_34100), .CD(n_61758), .Q(to_acu2
		[63]));
	notech_mux2 i_40878(.S(n_55032), .A(to_acu2[63]), .B(n_3625), .Z(n_34100
		));
	notech_reg to_acu2_reg_64(.CP(n_62311), .D(n_34106), .CD(n_61758), .Q(to_acu2
		[64]));
	notech_mux2 i_40886(.S(n_55033), .A(to_acu2[64]), .B(n_3623), .Z(n_34106
		));
	notech_reg to_acu2_reg_65(.CP(n_62311), .D(n_34112), .CD(n_61761), .Q(to_acu2
		[65]));
	notech_mux2 i_40894(.S(n_55032), .A(to_acu2[65]), .B(n_3621), .Z(n_34112
		));
	notech_and4 i_772(.A(n_2993), .B(n_231394270), .C(n_230694263), .D(n_2991
		), .Z(n_231094267));
	notech_reg to_acu2_reg_66(.CP(n_62311), .D(n_34118), .CD(n_61763), .Q(to_acu2
		[66]));
	notech_mux2 i_40902(.S(n_55032), .A(to_acu2[66]), .B(n_3619), .Z(n_34118
		));
	notech_or4 i_766(.A(n_40479), .B(n_2961), .C(n_54629), .D(n_40739), .Z(n_230994266
		));
	notech_reg to_acu2_reg_67(.CP(n_62311), .D(n_34124), .CD(n_61761), .Q(to_acu2
		[67]));
	notech_mux2 i_40910(.S(n_55032), .A(to_acu2[67]), .B(n_3617), .Z(n_34124
		));
	notech_reg to_acu2_reg_68(.CP(n_62311), .D(n_34130), .CD(n_61761), .Q(to_acu2
		[68]));
	notech_mux2 i_40918(.S(n_55027), .A(to_acu2[68]), .B(n_3615), .Z(n_34130
		));
	notech_reg to_acu2_reg_69(.CP(n_62309), .D(n_34136), .CD(n_61761), .Q(to_acu2
		[69]));
	notech_mux2 i_40926(.S(n_55027), .A(to_acu2[69]), .B(n_3613), .Z(n_34136
		));
	notech_nand3 i_767(.A(n_54629), .B(n_2962), .C(in128[36]), .Z(n_230694263
		));
	notech_reg to_acu2_reg_70(.CP(n_62309), .D(n_34142), .CD(n_61763), .Q(to_acu2
		[70]));
	notech_mux2 i_40934(.S(n_55032), .A(to_acu2[70]), .B(n_3611), .Z(n_34142
		));
	notech_or4 i_57(.A(n_225196458), .B(n_225096459), .C(n_40490), .D(n_40730
		), .Z(n_230594262));
	notech_reg to_acu2_reg_71(.CP(n_62309), .D(n_34148), .CD(n_61763), .Q(to_acu2
		[71]));
	notech_mux2 i_40942(.S(n_55027), .A(to_acu2[71]), .B(n_3609), .Z(n_34148
		));
	notech_reg to_acu2_reg_72(.CP(n_62309), .D(n_34154), .CD(n_61763), .Q(to_acu2
		[72]));
	notech_mux2 i_40950(.S(n_55027), .A(to_acu2[72]), .B(n_3607), .Z(n_34154
		));
	notech_reg to_acu2_reg_73(.CP(n_62309), .D(n_34160), .CD(n_61763), .Q(to_acu2
		[73]));
	notech_mux2 i_40958(.S(n_55027), .A(to_acu2[73]), .B(n_3605), .Z(n_34160
		));
	notech_and4 i_762(.A(n_2988), .B(n_230594262), .C(n_229894255), .D(n_2986
		), .Z(n_230294259));
	notech_reg to_acu2_reg_74(.CP(n_62309), .D(n_34166), .CD(n_61763), .Q(to_acu2
		[74]));
	notech_mux2 i_40966(.S(n_55032), .A(to_acu2[74]), .B(n_3603), .Z(n_34166
		));
	notech_or4 i_756(.A(n_40479), .B(n_2961), .C(n_54629), .D(n_40738), .Z(n_230194258
		));
	notech_reg to_acu2_reg_75(.CP(n_62309), .D(n_34172), .CD(n_61761), .Q(to_acu2
		[75]));
	notech_mux2 i_40974(.S(n_55032), .A(to_acu2[75]), .B(n_3601), .Z(n_34172
		));
	notech_reg to_acu2_reg_76(.CP(n_62309), .D(n_34178), .CD(n_61761), .Q(to_acu2
		[76]));
	notech_mux2 i_40982(.S(n_55032), .A(to_acu2[76]), .B(n_3599), .Z(n_34178
		));
	notech_reg to_acu2_reg_77(.CP(n_62309), .D(n_34184), .CD(n_61761), .Q(to_acu2
		[77]));
	notech_mux2 i_40990(.S(n_55032), .A(to_acu2[77]), .B(n_3597), .Z(n_34184
		));
	notech_nand3 i_757(.A(n_54629), .B(n_2962), .C(in128[35]), .Z(n_229894255
		));
	notech_reg to_acu2_reg_78(.CP(n_62309), .D(n_34190), .CD(n_61761), .Q(to_acu2
		[78]));
	notech_mux2 i_40998(.S(n_55032), .A(to_acu2[78]), .B(n_3595), .Z(n_34190
		));
	notech_or4 i_54(.A(n_225196458), .B(n_225096459), .C(n_40490), .D(n_40729
		), .Z(n_229794254));
	notech_reg to_acu2_reg_79(.CP(n_62309), .D(n_34196), .CD(n_61761), .Q(to_acu2
		[79]));
	notech_mux2 i_41006(.S(n_55032), .A(to_acu2[79]), .B(n_3593), .Z(n_34196
		));
	notech_reg to_acu2_reg_80(.CP(n_62306), .D(n_34202), .CD(n_61761), .Q(to_acu2
		[80]));
	notech_mux2 i_41014(.S(n_55032), .A(to_acu2[80]), .B(n_3591), .Z(n_34202
		));
	notech_reg to_acu2_reg_81(.CP(n_62301), .D(n_34208), .CD(n_61761), .Q(to_acu2
		[81]));
	notech_mux2 i_41022(.S(n_55033), .A(to_acu2[81]), .B(n_3589), .Z(n_34208
		));
	notech_and4 i_752(.A(n_2983), .B(n_229794254), .C(n_229094247), .D(n_2981
		), .Z(n_229494251));
	notech_reg to_acu2_reg_82(.CP(n_62301), .D(n_34214), .CD(n_61761), .Q(to_acu2
		[82]));
	notech_mux2 i_41030(.S(n_55038), .A(to_acu2[82]), .B(n_3587), .Z(n_34214
		));
	notech_or4 i_746(.A(n_40479), .B(n_2961), .C(n_54629), .D(n_40737), .Z(n_229394250
		));
	notech_reg to_acu2_reg_83(.CP(n_62301), .D(n_34220), .CD(n_61761), .Q(to_acu2
		[83]));
	notech_mux2 i_41038(.S(n_55038), .A(to_acu2[83]), .B(n_3585), .Z(n_34220
		));
	notech_reg to_acu2_reg_84(.CP(n_62301), .D(n_34226), .CD(n_61761), .Q(to_acu2
		[84]));
	notech_mux2 i_41046(.S(n_55038), .A(to_acu2[84]), .B(n_47642), .Z(n_34226
		));
	notech_reg to_acu2_reg_85(.CP(n_62301), .D(n_34232), .CD(n_61761), .Q(to_acu2
		[85]));
	notech_mux2 i_41054(.S(n_55033), .A(to_acu2[85]), .B(n_3583), .Z(n_34232
		));
	notech_nand3 i_747(.A(n_54629), .B(n_2962), .C(in128[34]), .Z(n_229094247
		));
	notech_reg to_acu2_reg_86(.CP(n_62301), .D(n_34238), .CD(n_61753), .Q(to_acu2
		[86]));
	notech_mux2 i_41062(.S(n_55033), .A(to_acu2[86]), .B(n_3581), .Z(n_34238
		));
	notech_or4 i_51(.A(n_225196458), .B(n_225096459), .C(n_40490), .D(n_40728
		), .Z(n_228994246));
	notech_reg to_acu2_reg_87(.CP(n_62304), .D(n_34244), .CD(n_61753), .Q(to_acu2
		[87]));
	notech_mux2 i_41070(.S(n_55038), .A(to_acu2[87]), .B(n_3579), .Z(n_34244
		));
	notech_reg to_acu2_reg_88(.CP(n_62301), .D(n_34250), .CD(n_61753), .Q(to_acu2
		[88]));
	notech_mux2 i_41078(.S(n_55038), .A(to_acu2[88]), .B(n_3577), .Z(n_34250
		));
	notech_reg to_acu2_reg_89(.CP(n_62301), .D(n_34256), .CD(n_61753), .Q(to_acu2
		[89]));
	notech_mux2 i_41086(.S(n_55038), .A(to_acu2[89]), .B(n_3575), .Z(n_34256
		));
	notech_and4 i_742(.A(n_2978), .B(n_228994246), .C(n_228294239), .D(n_2976
		), .Z(n_228694243));
	notech_reg to_acu2_reg_90(.CP(n_62301), .D(n_34262), .CD(n_61753), .Q(to_acu2
		[90]));
	notech_mux2 i_41094(.S(n_55038), .A(to_acu2[90]), .B(n_61750629), .Z(n_34262
		));
	notech_or4 i_736(.A(n_40479), .B(n_2961), .C(n_54629), .D(n_40736), .Z(n_228594242
		));
	notech_reg to_acu2_reg_91(.CP(n_62301), .D(n_34268), .CD(n_61756), .Q(to_acu2
		[91]));
	notech_mux2 i_41102(.S(n_55038), .A(to_acu2[91]), .B(n_161096305), .Z(n_34268
		));
	notech_reg to_acu2_reg_92(.CP(n_62301), .D(n_34274), .CD(n_61756), .Q(to_acu2
		[92]));
	notech_mux2 i_41110(.S(n_55038), .A(to_acu2[92]), .B(n_69550705), .Z(n_34274
		));
	notech_reg to_acu2_reg_93(.CP(n_62301), .D(n_34280), .CD(n_61756), .Q(to_acu2
		[93]));
	notech_mux2 i_41118(.S(n_55038), .A(to_acu2[93]), .B(n_161196306), .Z(n_34280
		));
	notech_nand3 i_737(.A(n_54629), .B(n_2962), .C(in128[33]), .Z(n_228294239
		));
	notech_reg to_acu2_reg_94(.CP(n_62301), .D(n_34286), .CD(n_61753), .Q(to_acu2
		[94]));
	notech_mux2 i_41126(.S(n_55038), .A(to_acu2[94]), .B(n_71350723), .Z(n_34286
		));
	notech_or4 i_48(.A(n_225196458), .B(n_225096459), .C(n_40490), .D(n_40727
		), .Z(n_228194238));
	notech_reg to_acu2_reg_95(.CP(n_62301), .D(n_34292), .CD(n_61753), .Q(to_acu2
		[95]));
	notech_mux2 i_41134(.S(n_55033), .A(to_acu2[95]), .B(n_73050740), .Z(n_34292
		));
	notech_reg to_acu2_reg_96(.CP(n_62301), .D(n_34298), .CD(n_61753), .Q(to_acu2
		[96]));
	notech_mux2 i_41142(.S(n_55033), .A(to_acu2[96]), .B(n_72450734), .Z(n_34298
		));
	notech_reg to_acu2_reg_97(.CP(n_62301), .D(n_34304), .CD(n_61753), .Q(to_acu2
		[97]));
	notech_mux2 i_41150(.S(n_55033), .A(to_acu2[97]), .B(n_70250712), .Z(n_34304
		));
	notech_and4 i_732(.A(n_2973), .B(n_228194238), .C(n_227494231), .D(n_2970
		), .Z(n_227894235));
	notech_reg to_acu2_reg_98(.CP(n_62301), .D(n_34310), .CD(n_61753), .Q(to_acu2
		[98]));
	notech_mux2 i_41158(.S(n_55033), .A(to_acu2[98]), .B(n_71550725), .Z(n_34310
		));
	notech_or4 i_725(.A(n_40479), .B(n_2961), .C(n_54629), .D(n_40735), .Z(n_227794234
		));
	notech_reg to_acu2_reg_99(.CP(n_62301), .D(n_34316), .CD(n_61753), .Q(to_acu2
		[99]));
	notech_mux2 i_41166(.S(n_55033), .A(to_acu2[99]), .B(n_69350703), .Z(n_34316
		));
	notech_reg to_acu2_reg_100(.CP(n_62301), .D(n_34322), .CD(n_61753), .Q(to_acu2
		[100]));
	notech_mux2 i_41174(.S(n_55033), .A(to_acu2[100]), .B(n_71050720), .Z(n_34322
		));
	notech_reg to_acu2_reg_101(.CP(n_62301), .D(n_34328), .CD(n_61753), .Q(to_acu2
		[101]));
	notech_mux2 i_41182(.S(n_55033), .A(to_acu2[101]), .B(n_70450714), .Z(n_34328
		));
	notech_nand3 i_726(.A(n_54629), .B(n_2962), .C(in128[32]), .Z(n_227494231
		));
	notech_reg to_acu2_reg_102(.CP(n_62304), .D(n_34334), .CD(n_61753), .Q(to_acu2
		[102]));
	notech_mux2 i_41190(.S(n_55033), .A(to_acu2[102]), .B(n_71750727), .Z(n_34334
		));
	notech_and3 i_629731(.A(n_40593), .B(n_40592), .C(n_40591), .Z(n_227396436
		));
	notech_reg to_acu2_reg_103(.CP(n_62304), .D(n_34340), .CD(n_61753), .Q(to_acu2
		[103]));
	notech_mux2 i_41198(.S(n_55033), .A(to_acu2[103]), .B(n_69950709), .Z(n_34340
		));
	notech_or4 i_210241(.A(int_excl[5]), .B(n_224496465), .C(n_224596464), .D
		(n_2922), .Z(n_227296437));
	notech_reg to_acu2_reg_104(.CP(n_62304), .D(n_34346), .CD(n_61753), .Q(to_acu2
		[104]));
	notech_mux2 i_41206(.S(n_55033), .A(to_acu2[104]), .B(n_69250702), .Z(n_34346
		));
	notech_reg to_acu2_reg_105(.CP(n_62304), .D(n_34352), .CD(n_61753), .Q(to_acu2
		[105]));
	notech_mux2 i_41214(.S(n_55033), .A(to_acu2[105]), .B(n_73650746), .Z(n_34352
		));
	notech_reg to_acu2_reg_106(.CP(n_62304), .D(n_34358), .CD(n_61753), .Q(to_acu2
		[106]));
	notech_mux2 i_41222(.S(n_55033), .A(to_acu2[106]), .B(n_72550735), .Z(n_34358
		));
	notech_and3 i_65832(.A(n_226596444), .B(n_2952), .C(n_2177), .Z(n_226996440
		));
	notech_reg to_acu2_reg_107(.CP(n_62306), .D(n_34364), .CD(n_61756), .Q(to_acu2
		[107]));
	notech_mux2 i_41230(.S(n_55033), .A(to_acu2[107]), .B(n_1962), .Z(n_34364
		));
	notech_reg to_acu2_reg_108(.CP(n_62306), .D(n_34370), .CD(n_61756), .Q(to_acu2
		[108]));
	notech_mux2 i_41238(.S(n_55054), .A(to_acu2[108]), .B(n_70050710), .Z(n_34370
		));
	notech_nand2 i_343(.A(n_226696443), .B(\to_acu2_0[26] ), .Z(n_226796442)
		);
	notech_reg to_acu2_reg_109(.CP(n_62304), .D(n_34376), .CD(n_61756), .Q(to_acu2
		[109]));
	notech_mux2 i_41246(.S(n_55067), .A(to_acu2[109]), .B(n_1979), .Z(n_34376
		));
	notech_nand2 i_646(.A(n_40907), .B(n_40906), .Z(n_226696443));
	notech_reg to_acu2_reg_110(.CP(n_62304), .D(n_34382), .CD(n_61756), .Q(to_acu2
		[110]));
	notech_mux2 i_41254(.S(n_55067), .A(to_acu2[110]), .B(n_2016), .Z(n_34382
		));
	notech_nand2 i_342(.A(\to_acu2_0[18] ), .B(\to_acu2_0[17] ), .Z(n_226596444
		));
	notech_reg to_acu2_reg_111(.CP(n_62304), .D(n_34388), .CD(n_61756), .Q(to_acu2
		[111]));
	notech_mux2 i_41262(.S(n_55067), .A(to_acu2[111]), .B(n_2014), .Z(n_34388
		));
	notech_nand2 i_640(.A(n_40896), .B(n_40895), .Z(n_226496445));
	notech_reg to_acu2_reg_112(.CP(n_62304), .D(n_34394), .CD(n_61758), .Q(to_acu2
		[112]));
	notech_mux2 i_41270(.S(n_55067), .A(to_acu2[112]), .B(n_1973), .Z(n_34394
		));
	notech_reg to_acu2_reg_113(.CP(n_62304), .D(n_34400), .CD(n_61758), .Q(to_acu2
		[113]));
	notech_mux2 i_41278(.S(n_55067), .A(to_acu2[113]), .B(n_1974), .Z(n_34400
		));
	notech_reg to_acu2_reg_114(.CP(n_62304), .D(n_34406), .CD(n_61758), .Q(to_acu2
		[114]));
	notech_mux2 i_41286(.S(n_55067), .A(to_acu2[114]), .B(n_1988), .Z(n_34406
		));
	notech_and2 i_45(.A(n_2947), .B(in128[59]), .Z(n_226196448));
	notech_reg to_acu2_reg_115(.CP(n_62304), .D(n_34412), .CD(n_61756), .Q(to_acu2
		[115]));
	notech_mux2 i_41294(.S(n_55067), .A(to_acu2[115]), .B(n_2006), .Z(n_34412
		));
	notech_nand2 i_571(.A(n_40489), .B(n_40491), .Z(n_226096449));
	notech_reg to_acu2_reg_116(.CP(n_62304), .D(n_34418), .CD(n_61758), .Q(to_acu2
		[116]));
	notech_mux2 i_41302(.S(n_55067), .A(to_acu2[116]), .B(n_2007), .Z(n_34418
		));
	notech_reg to_acu2_reg_117(.CP(n_62304), .D(n_34424), .CD(n_61756), .Q(to_acu2
		[117]));
	notech_mux2 i_41310(.S(n_55067), .A(to_acu2[117]), .B(n_2008), .Z(n_34424
		));
	notech_nand3 i_629764(.A(n_40591), .B(n_40593), .C(imm_sz[1]), .Z(n_225896451
		));
	notech_reg to_acu2_reg_118(.CP(n_62304), .D(n_34430), .CD(n_61756), .Q(to_acu2
		[118]));
	notech_mux2 i_41318(.S(n_55067), .A(to_acu2[118]), .B(n_1995), .Z(n_34430
		));
	notech_reg to_acu2_reg_119(.CP(n_62304), .D(n_34436), .CD(n_61756), .Q(to_acu2
		[119]));
	notech_mux2 i_41326(.S(n_55067), .A(to_acu2[119]), .B(n_2001), .Z(n_34436
		));
	notech_reg to_acu2_reg_120(.CP(n_62304), .D(n_34442), .CD(n_61756), .Q(to_acu2
		[120]));
	notech_mux2 i_41334(.S(n_55067), .A(to_acu2[120]), .B(n_2003), .Z(n_34442
		));
	notech_reg to_acu2_reg_121(.CP(n_62304), .D(n_34448), .CD(n_61756), .Q(to_acu2
		[121]));
	notech_mux2 i_41342(.S(n_55067), .A(to_acu2[121]), .B(n_2000), .Z(n_34448
		));
	notech_reg to_acu2_reg_122(.CP(n_62304), .D(n_34454), .CD(n_61756), .Q(to_acu2
		[122]));
	notech_mux2 i_41350(.S(n_55066), .A(to_acu2[122]), .B(n_1986), .Z(n_34454
		));
	notech_reg to_acu2_reg_123(.CP(n_62320), .D(n_34460), .CD(n_61756), .Q(to_acu2
		[123]));
	notech_mux2 i_41358(.S(n_55066), .A(to_acu2[123]), .B(n_2012), .Z(n_34460
		));
	notech_reg to_acu2_reg_124(.CP(n_62320), .D(n_34466), .CD(n_61756), .Q(to_acu2
		[124]));
	notech_mux2 i_41366(.S(n_55066), .A(to_acu2[124]), .B(n_1968), .Z(n_34466
		));
	notech_nor2 i_554(.A(displc[2]), .B(n_2932), .Z(n_225196458));
	notech_reg to_acu2_reg_125(.CP(n_62320), .D(n_34472), .CD(n_61756), .Q(to_acu2
		[125]));
	notech_mux2 i_41374(.S(n_55066), .A(to_acu2[125]), .B(n_1997), .Z(n_34472
		));
	notech_and2 i_553(.A(displc[2]), .B(n_2932), .Z(n_225096459));
	notech_reg to_acu2_reg_126(.CP(n_62317), .D(n_34478), .CD(n_61756), .Q(to_acu2
		[126]));
	notech_mux2 i_41382(.S(n_55066), .A(to_acu2[126]), .B(n_2002), .Z(n_34478
		));
	notech_and2 i_277(.A(n_40919), .B(n_40594), .Z(n_224996460));
	notech_reg to_acu2_reg_127(.CP(n_62320), .D(n_34484), .CD(n_61756), .Q(to_acu2
		[127]));
	notech_mux2 i_41390(.S(n_55066), .A(to_acu2[127]), .B(n_1987), .Z(n_34484
		));
	notech_reg to_acu2_reg_128(.CP(n_62320), .D(n_34490), .CD(n_61763), .Q(to_acu2
		[128]));
	notech_mux2 i_41398(.S(n_55066), .A(to_acu2[128]), .B(n_1978), .Z(n_34490
		));
	notech_reg to_acu2_reg_129(.CP(n_62320), .D(n_34496), .CD(n_61772), .Q(to_acu2
		[129]));
	notech_mux2 i_41406(.S(n_55067), .A(to_acu2[129]), .B(n_1971), .Z(n_34496
		));
	notech_nand2 i_546(.A(n_40593), .B(imm_sz[0]), .Z(n_224696463));
	notech_reg to_acu2_reg_130(.CP(n_62320), .D(n_34502), .CD(n_61772), .Q(to_acu2
		[130]));
	notech_mux2 i_41414(.S(n_55067), .A(to_acu2[130]), .B(n_1981), .Z(n_34502
		));
	notech_and4 i_23(.A(n_39341), .B(n_39339), .C(n_2926), .D(n_2925), .Z(n_224596464
		));
	notech_reg to_acu2_reg_131(.CP(n_62320), .D(n_34508), .CD(n_61772), .Q(to_acu2
		[131]));
	notech_mux2 i_41422(.S(n_55067), .A(to_acu2[131]), .B(n_2010), .Z(n_34508
		));
	notech_or4 i_168(.A(int_excl[2]), .B(int_excl[3]), .C(int_excl[4]), .D(n_5423
		), .Z(n_224496465));
	notech_reg to_acu2_reg_132(.CP(n_62320), .D(n_34514), .CD(n_61772), .Q(to_acu2
		[132]));
	notech_mux2 i_41430(.S(n_55066), .A(to_acu2[132]), .B(n_2015), .Z(n_34514
		));
	notech_nao3 i_139(.A(n_40937), .B(n_59969), .C(n_2870), .Z(n_224396466)
		);
	notech_reg to_acu2_reg_133(.CP(n_62317), .D(n_34520), .CD(n_61772), .Q(to_acu2
		[133]));
	notech_mux2 i_41438(.S(n_55067), .A(to_acu2[133]), .B(n_1999), .Z(n_34520
		));
	notech_nand3 i_829762(.A(n_40591), .B(imm_sz[1]), .C(imm_sz[2]), .Z(n_224296467
		));
	notech_reg to_acu2_reg_134(.CP(n_62317), .D(n_34526), .CD(n_61772), .Q(to_acu2
		[134]));
	notech_mux2 i_41446(.S(n_55067), .A(to_acu2[134]), .B(n_1996), .Z(n_34526
		));
	notech_ao4 i_43(.A(n_59529), .B(n_2916), .C(n_223796472), .D(pc_req), .Z
		(n_224196468));
	notech_reg to_acu2_reg_135(.CP(n_62317), .D(n_34532), .CD(n_61772), .Q(to_acu2
		[135]));
	notech_mux2 i_41454(.S(n_55072), .A(to_acu2[135]), .B(n_1969), .Z(n_34532
		));
	notech_reg to_acu2_reg_136(.CP(n_62317), .D(n_34538), .CD(n_61772), .Q(to_acu2
		[136]));
	notech_mux2 i_41462(.S(n_55077), .A(to_acu2[136]), .B(n_2013), .Z(n_34538
		));
	notech_ao3 i_3229868(.A(n_2218), .B(n_40723), .C(n_2215), .Z(n_223996470
		));
	notech_reg to_acu2_reg_137(.CP(n_62317), .D(n_34544), .CD(n_61772), .Q(to_acu2
		[137]));
	notech_mux2 i_41470(.S(n_55077), .A(to_acu2[137]), .B(n_2009), .Z(n_34544
		));
	notech_reg to_acu2_reg_138(.CP(n_62317), .D(n_34550), .CD(n_61772), .Q(to_acu2
		[138]));
	notech_mux2 i_41478(.S(n_55077), .A(to_acu2[138]), .B(n_1983), .Z(n_34550
		));
	notech_mux2 i_44(.S(n_5414), .A(n_223396476), .B(n_223596474), .Z(n_223796472
		));
	notech_reg to_acu2_reg_139(.CP(n_62317), .D(n_34556), .CD(n_61769), .Q(to_acu2
		[139]));
	notech_mux2 i_41486(.S(n_55077), .A(to_acu2[139]), .B(n_1989), .Z(n_34556
		));
	notech_reg to_acu2_reg_140(.CP(n_62317), .D(n_34562), .CD(n_61769), .Q(to_acu2
		[140]));
	notech_mux2 i_41494(.S(n_55077), .A(to_acu2[140]), .B(n_1990), .Z(n_34562
		));
	notech_ao3 i_65888(.A(fsm[0]), .B(fsm[1]), .C(n_2865), .Z(n_223596474)
		);
	notech_reg to_acu2_reg_141(.CP(n_62317), .D(n_34568), .CD(n_61769), .Q(to_acu2
		[141]));
	notech_mux2 i_41502(.S(n_55077), .A(to_acu2[141]), .B(n_1965), .Z(n_34568
		));
	notech_reg to_acu2_reg_142(.CP(n_62317), .D(n_34574), .CD(n_61769), .Q(to_acu2
		[142]));
	notech_mux2 i_41510(.S(n_55077), .A(to_acu2[142]), .B(n_1991), .Z(n_34574
		));
	notech_and2 i_4230(.A(n_5408), .B(n_2219), .Z(n_223396476));
	notech_reg to_acu2_reg_143(.CP(n_62317), .D(n_34580), .CD(n_61769), .Q(to_acu2
		[143]));
	notech_mux2 i_41518(.S(n_55077), .A(to_acu2[143]), .B(n_1992), .Z(n_34580
		));
	notech_reg to_acu2_reg_144(.CP(n_62322), .D(n_34586), .CD(n_61769), .Q(to_acu2
		[144]));
	notech_mux2 i_41526(.S(n_55077), .A(to_acu2[144]), .B(n_1966), .Z(n_34586
		));
	notech_and4 i_71506(.A(n_2912), .B(n_59082), .C(n_1949), .D(n_2230), .Z(n_223196478
		));
	notech_reg to_acu2_reg_145(.CP(n_62322), .D(n_34592), .CD(n_61769), .Q(to_acu2
		[145]));
	notech_mux2 i_41534(.S(n_55077), .A(to_acu2[145]), .B(n_1993), .Z(n_34592
		));
	notech_nao3 i_2842(.A(n_58991), .B(n_2170), .C(n_40559), .Z(n_2230));
	notech_reg to_acu2_reg_146(.CP(n_62322), .D(n_34598), .CD(n_61769), .Q(to_acu2
		[146]));
	notech_mux2 i_41542(.S(n_55077), .A(to_acu2[146]), .B(n_1994), .Z(n_34598
		));
	notech_nand2 i_509(.A(n_2910), .B(n_2222), .Z(n_2229));
	notech_reg to_acu2_reg_147(.CP(n_62322), .D(n_34604), .CD(n_61769), .Q(to_acu2
		[147]));
	notech_mux2 i_41550(.S(n_55077), .A(to_acu2[147]), .B(n_1982), .Z(n_34604
		));
	notech_nao3 i_508(.A(n_40937), .B(n_59969), .C(n_2908), .Z(n_2228));
	notech_reg to_acu2_reg_148(.CP(n_62322), .D(n_34610), .CD(n_61769), .Q(to_acu2
		[148]));
	notech_mux2 i_41558(.S(n_55077), .A(to_acu2[148]), .B(n_1955), .Z(n_34610
		));
	notech_nor2 i_163(.A(n_2171), .B(n_2223), .Z(n_2227));
	notech_reg to_acu2_reg_149(.CP(n_62322), .D(n_34616), .CD(n_61769), .Q(to_acu2
		[149]));
	notech_mux2 i_41566(.S(n_55072), .A(to_acu2[149]), .B(n_1959), .Z(n_34616
		));
	notech_nand2 i_497(.A(n_39195), .B(n_2870), .Z(n_2226));
	notech_reg to_acu2_reg_150(.CP(n_62322), .D(n_34622), .CD(n_61774), .Q(to_acu2
		[150]));
	notech_mux2 i_41574(.S(n_55072), .A(to_acu2[150]), .B(n_1961), .Z(n_34622
		));
	notech_nand2 i_212(.A(fpu), .B(n_2222), .Z(n_2225));
	notech_reg to_acu2_reg_151(.CP(n_62322), .D(n_34628), .CD(n_61774), .Q(to_acu2
		[151]));
	notech_mux2 i_41582(.S(n_55072), .A(to_acu2[151]), .B(n_69450704), .Z(n_34628
		));
	notech_nao3 i_483(.A(n_40938), .B(\to_acu2_0[62] ), .C(twobyte), .Z(n_2224
		));
	notech_reg to_acu2_reg_152(.CP(n_62322), .D(n_34634), .CD(n_61774), .Q(to_acu2
		[152]));
	notech_mux2 i_41590(.S(n_55072), .A(to_acu2[152]), .B(n_1977), .Z(n_34634
		));
	notech_ao3 i_482(.A(n_40938), .B(\to_acu2_0[69] ), .C(twobyte), .Z(n_2223
		));
	notech_reg to_acu2_reg_153(.CP(n_62322), .D(n_34640), .CD(n_61774), .Q(to_acu2
		[153]));
	notech_mux2 i_41598(.S(n_55072), .A(to_acu2[153]), .B(n_1967), .Z(n_34640
		));
	notech_and4 i_28(.A(n_2220), .B(n_1507), .C(n_2886), .D(n_40498), .Z(n_2222
		));
	notech_reg to_acu2_reg_154(.CP(n_62320), .D(n_34646), .CD(n_61774), .Q(to_acu2
		[154]));
	notech_mux2 i_41606(.S(n_55072), .A(to_acu2[154]), .B(n_1972), .Z(n_34646
		));
	notech_and2 i_347(.A(valid_len[0]), .B(valid_len[1]), .Z(n_2221));
	notech_reg to_acu2_reg_155(.CP(n_62320), .D(n_34652), .CD(n_61774), .Q(to_acu2
		[155]));
	notech_mux2 i_41614(.S(n_55072), .A(to_acu2[155]), .B(n_1970), .Z(n_34652
		));
	notech_or4 i_471(.A(valid_len[2]), .B(valid_len[5]), .C(n_2890), .D(n_2221
		), .Z(n_2220));
	notech_reg to_acu2_reg_156(.CP(n_62320), .D(n_34658), .CD(n_61774), .Q(to_acu2
		[156]));
	notech_mux2 i_41622(.S(n_55072), .A(to_acu2[156]), .B(n_48074), .Z(n_34658
		));
	notech_nand2 i_429870(.A(idx_deco[1]), .B(idx_deco[0]), .Z(n_2219));
	notech_reg to_acu2_reg_157(.CP(n_62320), .D(n_34664), .CD(n_61774), .Q(to_acu2
		[157]));
	notech_mux2 i_41630(.S(n_55077), .A(to_acu2[157]), .B(n_2004), .Z(n_34664
		));
	notech_nand2 i_458(.A(n_2875), .B(valid_len[4]), .Z(n_2218));
	notech_reg to_acu2_reg_158(.CP(n_62320), .D(n_34670), .CD(n_61774), .Q(to_acu2
		[158]));
	notech_mux2 i_41638(.S(n_55077), .A(to_acu2[158]), .B(n_3534), .Z(n_34670
		));
	notech_reg to_acu2_reg_159(.CP(n_62320), .D(n_34676), .CD(n_61774), .Q(to_acu2
		[159]));
	notech_mux2 i_41646(.S(n_55072), .A(to_acu2[159]), .B(n_1998), .Z(n_34676
		));
	notech_reg to_acu2_reg_160(.CP(n_62320), .D(n_34682), .CD(n_61774), .Q(to_acu2
		[160]));
	notech_mux2 i_41654(.S(n_55072), .A(to_acu2[160]), .B(n_1964), .Z(n_34682
		));
	notech_ao4 i_459(.A(n_2212), .B(n_2211), .C(valid_len[4]), .D(n_2875), .Z
		(n_2215));
	notech_reg to_acu2_reg_161(.CP(n_62320), .D(n_34688), .CD(n_61772), .Q(to_acu2
		[161]));
	notech_mux2 i_41662(.S(n_55072), .A(to_acu2[161]), .B(n_1985), .Z(n_34688
		));
	notech_reg to_acu2_reg_162(.CP(n_62320), .D(n_34694), .CD(n_61772), .Q(to_acu2
		[162]));
	notech_mux2 i_41670(.S(n_55055), .A(to_acu2[162]), .B(n_1956), .Z(n_34694
		));
	notech_reg to_acu2_reg_163(.CP(n_62320), .D(n_34700), .CD(n_61772), .Q(to_acu2
		[163]));
	notech_mux2 i_41678(.S(n_55055), .A(to_acu2[163]), .B(n_72150731), .Z(n_34700
		));
	notech_ao4 i_455(.A(n_2208), .B(n_2207), .C(valid_len[3]), .D(n_2876), .Z
		(n_2212));
	notech_reg to_acu2_reg_164(.CP(n_62320), .D(n_34706), .CD(n_61772), .Q(to_acu2
		[164]));
	notech_mux2 i_41686(.S(n_55055), .A(to_acu2[164]), .B(n_73850748), .Z(n_34706
		));
	notech_and2 i_450(.A(n_2876), .B(valid_len[3]), .Z(n_2211));
	notech_reg to_acu2_reg_165(.CP(n_62317), .D(n_34712), .CD(n_61772), .Q(to_acu2
		[165]));
	notech_mux2 i_41694(.S(n_55055), .A(to_acu2[165]), .B(n_73450744), .Z(n_34712
		));
	notech_reg to_acu2_reg_166(.CP(n_62311), .D(n_34718), .CD(n_61772), .Q(to_acu2
		[166]));
	notech_mux2 i_41702(.S(n_55055), .A(to_acu2[166]), .B(n_72950739), .Z(n_34718
		));
	notech_reg to_acu2_reg_167(.CP(n_62315), .D(n_34724), .CD(n_61772), .Q(to_acu2
		[167]));
	notech_mux2 i_41710(.S(n_55055), .A(to_acu2[167]), .B(n_3526), .Z(n_34724
		));
	notech_ao4 i_449(.A(valid_len[2]), .B(n_40504), .C(n_2204), .D(n_2203), 
		.Z(n_2208));
	notech_reg to_acu2_reg_168(.CP(n_62311), .D(n_34730), .CD(n_61772), .Q(to_acu2
		[168]));
	notech_mux2 i_41718(.S(n_55055), .A(to_acu2[168]), .B(n_1963), .Z(n_34730
		));
	notech_and2 i_447(.A(valid_len[2]), .B(n_40504), .Z(n_2207));
	notech_reg to_acu2_reg_169(.CP(n_62311), .D(n_34736), .CD(n_61772), .Q(to_acu2
		[169]));
	notech_mux2 i_41726(.S(n_55055), .A(to_acu2[169]), .B(n_3523), .Z(n_34736
		));
	notech_xor2 i_6335(.A(imm_sz[0]), .B(i_ptr[0]), .Z(n_2206));
	notech_reg to_acu2_reg_170(.CP(n_62311), .D(n_34742), .CD(n_61772), .Q(to_acu2
		[170]));
	notech_mux2 i_41734(.S(n_55055), .A(to_acu2[170]), .B(n_3521), .Z(n_34742
		));
	notech_or2 i_346(.A(valid_len[1]), .B(n_40503), .Z(n_2205));
	notech_reg to_acu2_reg_171(.CP(n_62315), .D(n_34748), .CD(n_61767), .Q(to_acu2
		[171]));
	notech_mux2 i_41742(.S(n_55055), .A(to_acu2[171]), .B(n_3519), .Z(n_34748
		));
	notech_ao3 i_445(.A(valid_len[0]), .B(n_2205), .C(n_2206), .Z(n_2204));
	notech_reg to_acu2_reg_172(.CP(n_62315), .D(n_34754), .CD(n_61767), .Q(to_acu2
		[172]));
	notech_mux2 i_41750(.S(n_55055), .A(to_acu2[172]), .B(n_2021), .Z(n_34754
		));
	notech_and2 i_441(.A(valid_len[1]), .B(n_40503), .Z(n_2203));
	notech_reg to_acu2_reg_173(.CP(n_62315), .D(n_34760), .CD(n_61767), .Q(to_acu2
		[173]));
	notech_mux2 i_41758(.S(n_55055), .A(to_acu2[173]), .B(n_3516), .Z(n_34760
		));
	notech_reg to_acu2_reg_174(.CP(n_62315), .D(n_34766), .CD(n_61763), .Q(to_acu2
		[174]));
	notech_mux2 i_41766(.S(n_55055), .A(to_acu2[174]), .B(n_3514), .Z(n_34766
		));
	notech_reg to_acu2_reg_175(.CP(n_62315), .D(n_34772), .CD(n_61763), .Q(to_acu2
		[175]));
	notech_mux2 i_41774(.S(n_55054), .A(to_acu2[175]), .B(n_3512), .Z(n_34772
		));
	notech_reg to_acu2_reg_176(.CP(n_62311), .D(n_34778), .CD(n_61767), .Q(to_acu2
		[176]));
	notech_mux2 i_41782(.S(n_55054), .A(to_acu2[176]), .B(n_2020), .Z(n_34778
		));
	notech_reg to_acu2_reg_177(.CP(n_62311), .D(n_34784), .CD(n_61767), .Q(to_acu2
		[177]));
	notech_mux2 i_41790(.S(n_55054), .A(to_acu2[177]), .B(n_3509), .Z(n_34784
		));
	notech_reg to_acu2_reg_178(.CP(n_62311), .D(n_34790), .CD(n_61767), .Q(to_acu2
		[178]));
	notech_mux2 i_41798(.S(n_55054), .A(to_acu2[178]), .B(n_3507), .Z(n_34790
		));
	notech_and2 i_288(.A(n_40593), .B(n_39368), .Z(n_2197));
	notech_reg to_acu2_reg_179(.CP(n_62311), .D(n_34796), .CD(n_61767), .Q(to_acu2
		[179]));
	notech_mux2 i_41806(.S(n_55054), .A(to_acu2[179]), .B(n_3505), .Z(n_34796
		));
	notech_reg to_acu2_reg_180(.CP(n_62311), .D(n_34802), .CD(n_61767), .Q(to_acu2
		[180]));
	notech_mux2 i_41814(.S(n_55054), .A(to_acu2[180]), .B(n_3275), .Z(n_34802
		));
	notech_reg to_acu2_reg_181(.CP(n_62311), .D(n_34808), .CD(n_61763), .Q(to_acu2
		[181]));
	notech_mux2 i_41822(.S(n_55054), .A(to_acu2[181]), .B(n_3503), .Z(n_34808
		));
	notech_and2 i_287(.A(i_ptr[1]), .B(imm_sz[1]), .Z(n_2194));
	notech_reg to_acu2_reg_182(.CP(n_62311), .D(n_34814), .CD(n_61763), .Q(to_acu2
		[182]));
	notech_mux2 i_41830(.S(n_55054), .A(to_acu2[182]), .B(n_3501), .Z(n_34814
		));
	notech_reg to_acu2_reg_183(.CP(n_62311), .D(n_34820), .CD(n_61763), .Q(to_acu2
		[183]));
	notech_mux2 i_41838(.S(n_55054), .A(to_acu2[183]), .B(n_3499), .Z(n_34820
		));
	notech_reg to_acu2_reg_184(.CP(n_62311), .D(n_34826), .CD(n_61763), .Q(to_acu2
		[184]));
	notech_mux2 i_41846(.S(n_55054), .A(to_acu2[184]), .B(n_3497), .Z(n_34826
		));
	notech_and4 i_75059(.A(n_60059), .B(n_224396466), .C(n_18051052), .D(n_2189
		), .Z(n_2191));
	notech_reg to_acu2_reg_185(.CP(n_62311), .D(n_34832), .CD(n_61763), .Q(to_acu2
		[185]));
	notech_mux2 i_41854(.S(n_55054), .A(to_acu2[185]), .B(n_3495), .Z(n_34832
		));
	notech_and4 i_40(.A(n_2181), .B(n_2180), .C(n_2188), .D(n_2185), .Z(n_2190
		));
	notech_reg to_acu2_reg_186(.CP(n_62311), .D(n_34838), .CD(n_61763), .Q(to_acu2
		[186]));
	notech_mux2 i_41862(.S(n_55054), .A(to_acu2[186]), .B(n_3493), .Z(n_34838
		));
	notech_or2 i_389(.A(n_2837), .B(n_2190), .Z(n_2189));
	notech_reg to_acu2_reg_187(.CP(n_62317), .D(n_34844), .CD(n_61763), .Q(to_acu2
		[187]));
	notech_mux2 i_41870(.S(n_55054), .A(to_acu2[187]), .B(n_3491), .Z(n_34844
		));
	notech_nand2 i_382(.A(twobyte), .B(n_2187), .Z(n_2188));
	notech_reg to_acu2_reg_188(.CP(n_62317), .D(n_34850), .CD(n_61763), .Q(to_acu2
		[188]));
	notech_mux2 i_41878(.S(n_55055), .A(to_acu2[188]), .B(n_3489), .Z(n_34850
		));
	notech_nand2 i_41(.A(n_40912), .B(n_40873), .Z(n_2187));
	notech_reg to_acu2_reg_189(.CP(n_62315), .D(n_34856), .CD(n_61763), .Q(to_acu2
		[189]));
	notech_mux2 i_41886(.S(n_55066), .A(to_acu2[189]), .B(n_3487), .Z(n_34856
		));
	notech_nao3 i_42(.A(n_1773), .B(n_2860), .C(n_1931), .Z(n_2186));
	notech_reg to_acu2_reg_190(.CP(n_62315), .D(n_34862), .CD(n_61763), .Q(to_acu2
		[190]));
	notech_mux2 i_41894(.S(n_55066), .A(to_acu2[190]), .B(n_3485), .Z(n_34862
		));
	notech_nao3 i_381(.A(n_40939), .B(n_2186), .C(n_2851), .Z(n_2185));
	notech_reg to_acu2_reg_191(.CP(n_62315), .D(n_34868), .CD(n_61763), .Q(to_acu2
		[191]));
	notech_mux2 i_41902(.S(n_55066), .A(to_acu2[191]), .B(n_3483), .Z(n_34868
		));
	notech_nand2 i_374(.A(n_1932), .B(n_40865), .Z(n_2184));
	notech_reg to_acu2_reg_192(.CP(n_62317), .D(n_34874), .CD(n_61769), .Q(to_acu2
		[192]));
	notech_mux2 i_41910(.S(n_55061), .A(to_acu2[192]), .B(n_3481), .Z(n_34874
		));
	notech_nand2 i_367(.A(\to_acu2_0[5] ), .B(\to_acu2_0[59] ), .Z(n_2183)
		);
	notech_reg to_acu2_reg_193(.CP(n_62317), .D(n_34880), .CD(n_61769), .Q(to_acu2
		[193]));
	notech_mux2 i_41918(.S(n_55061), .A(to_acu2[193]), .B(n_3479), .Z(n_34880
		));
	notech_nand2 i_278(.A(n_40891), .B(n_40890), .Z(n_2182));
	notech_reg to_acu2_reg_194(.CP(n_62317), .D(n_34886), .CD(n_61769), .Q(to_acu2
		[194]));
	notech_mux2 i_41926(.S(n_55061), .A(to_acu2[194]), .B(n_3477), .Z(n_34886
		));
	notech_nand3 i_365(.A(twobyte), .B(n_40912), .C(n_2182), .Z(n_2181));
	notech_reg to_acu2_reg_195(.CP(n_62317), .D(n_34892), .CD(n_61767), .Q(to_acu2
		[195]));
	notech_mux2 i_41934(.S(n_55066), .A(to_acu2[195]), .B(n_3276), .Z(n_34892
		));
	notech_nand2 i_364(.A(n_2851), .B(n_40939), .Z(n_2180));
	notech_reg to_acu2_reg_196(.CP(n_62317), .D(n_34898), .CD(n_61769), .Q(to_acu2
		[196]));
	notech_mux2 i_41942(.S(n_55066), .A(to_acu2[196]), .B(n_3475), .Z(n_34898
		));
	notech_nand2 i_348(.A(\to_acu2_0[5] ), .B(\to_acu2_0[48] ), .Z(n_2179)
		);
	notech_reg to_acu2_reg_197(.CP(n_62315), .D(n_34904), .CD(n_61769), .Q(to_acu2
		[197]));
	notech_mux2 i_41950(.S(n_55066), .A(to_acu2[197]), .B(n_3473), .Z(n_34904
		));
	notech_nand3 i_344(.A(\to_acu2_0[23] ), .B(\to_acu2_0[21] ), .C(\to_acu2_0[22] 
		), .Z(n_2178));
	notech_reg to_acu2_reg_198(.CP(n_62315), .D(n_34910), .CD(n_61769), .Q(to_acu2
		[198]));
	notech_mux2 i_41958(.S(n_55066), .A(to_acu2[198]), .B(n_3471), .Z(n_34910
		));
	notech_nand2 i_341(.A(n_226496445), .B(\to_acu2_0[13] ), .Z(n_2177));
	notech_reg to_acu2_reg_199(.CP(n_62315), .D(n_34916), .CD(n_61769), .Q(to_acu2
		[199]));
	notech_mux2 i_41966(.S(n_55066), .A(to_acu2[199]), .B(n_3469), .Z(n_34916
		));
	notech_and4 i_306(.A(n_40916), .B(n_40922), .C(n_40915), .D(n_40923), .Z
		(n_2176));
	notech_reg to_acu2_reg_200(.CP(n_62315), .D(n_34922), .CD(n_61769), .Q(to_acu2
		[200]));
	notech_mux2 i_41974(.S(n_55066), .A(to_acu2[200]), .B(n_3467), .Z(n_34922
		));
	notech_reg to_acu2_reg_201(.CP(n_62315), .D(n_34928), .CD(n_61769), .Q(to_acu2
		[201]));
	notech_mux2 i_41982(.S(n_55066), .A(to_acu2[201]), .B(n_3465), .Z(n_34928
		));
	notech_or4 i_4106(.A(n_40490), .B(n_1643), .C(n_225196458), .D(n_225096459
		), .Z(n_2174));
	notech_reg to_acu2_reg_202(.CP(n_62315), .D(n_34934), .CD(n_61767), .Q(to_acu2
		[202]));
	notech_mux2 i_41990(.S(n_55055), .A(to_acu2[202]), .B(n_3463), .Z(n_34934
		));
	notech_or4 i_4108(.A(n_40479), .B(n_2961), .C(n_54629), .D(n_2149), .Z(n_2173
		));
	notech_reg to_acu2_reg_203(.CP(n_62315), .D(n_34940), .CD(n_61767), .Q(to_acu2
		[203]));
	notech_mux2 i_41998(.S(n_55061), .A(to_acu2[203]), .B(n_3461), .Z(n_34940
		));
	notech_or2 i_4107(.A(n_2149), .B(n_2965), .Z(n_2172));
	notech_reg to_acu2_reg_204(.CP(n_62315), .D(n_34946), .CD(n_61767), .Q(to_acu2
		[204]));
	notech_mux2 i_42006(.S(n_55061), .A(to_acu2[204]), .B(n_48362), .Z(n_34946
		));
	notech_nor2 i_6336(.A(n_2176), .B(n_2901), .Z(n_2171));
	notech_reg to_acu2_reg_205(.CP(n_62315), .D(n_34952), .CD(n_61767), .Q(to_acu2
		[205]));
	notech_mux2 i_42014(.S(n_55055), .A(to_acu2[205]), .B(n_48368), .Z(n_34952
		));
	notech_or4 i_72045(.A(db67), .B(\to_acu2_0[4] ), .C(\to_acu2_0[3] ), .D(n_2898
		), .Z(n_2170));
	notech_reg to_acu2_reg_206(.CP(n_62315), .D(n_34958), .CD(n_61767), .Q(to_acu2
		[206]));
	notech_mux2 i_42022(.S(n_55055), .A(to_acu2[206]), .B(n_48374), .Z(n_34958
		));
	notech_nor2 i_33174157(.A(n_2119), .B(n_59534), .Z(n_44695));
	notech_reg to_acu2_reg_207(.CP(n_62315), .D(n_34964), .CD(n_61767), .Q(to_acu2
		[207]));
	notech_mux2 i_42030(.S(n_55055), .A(to_acu2[207]), .B(n_48380), .Z(n_34964
		));
	notech_nor2 i_31574158(.A(n_2122), .B(n_59534), .Z(n_44599));
	notech_reg to_acu2_reg_208(.CP(n_62252), .D(n_34970), .CD(n_61767), .Q(to_acu2
		[208]));
	notech_mux2 i_42038(.S(n_55061), .A(to_acu2[208]), .B(n_48386), .Z(n_34970
		));
	notech_nor2 i_30474160(.A(n_2126), .B(n_59534), .Z(n_44533));
	notech_reg to_acu2_reg_209(.CP(n_62185), .D(n_34976), .CD(n_61767), .Q(to_acu2
		[209]));
	notech_mux2 i_42046(.S(n_55061), .A(to_acu2[209]), .B(n_48392), .Z(n_34976
		));
	notech_reg to_acu2_reg_210(.CP(n_62185), .D(n_34982), .CD(n_61767), .Q(to_acu2
		[210]));
	notech_mux2 i_42054(.S(n_55061), .A(to_acu2[210]), .B(n_48398), .Z(n_34982
		));
	notech_and2 i_14(.A(n_239994356), .B(n_224296467), .Z(n_2168));
	notech_reg to_acu1_reg_0(.CP(n_62185), .D(n_34988), .CD(n_61767), .Q(to_acu1
		[0]));
	notech_mux2 i_42062(.S(n_58327), .A(to_acu1[0]), .B(n_40238), .Z(n_34988
		));
	notech_reg to_acu1_reg_1(.CP(n_62185), .D(n_34994), .CD(n_61767), .Q(to_acu1
		[1]));
	notech_mux2 i_42070(.S(n_58332), .A(to_acu1[1]), .B(n_40240), .Z(n_34994
		));
	notech_reg to_acu1_reg_2(.CP(n_62185), .D(n_35000), .CD(n_61637), .Q(to_acu1
		[2]));
	notech_mux2 i_42078(.S(n_58332), .A(to_acu1[2]), .B(n_40177), .Z(n_35000
		));
	notech_reg to_acu1_reg_3(.CP(n_62185), .D(n_35006), .CD(n_61637), .Q(to_acu1
		[3]));
	notech_mux2 i_42086(.S(n_58332), .A(to_acu1[3]), .B(n_40179), .Z(n_35006
		));
	notech_ao4 i_95273212(.A(n_40760), .B(n_3045), .C(n_40768), .D(n_3046), 
		.Z(n_2164));
	notech_reg to_acu1_reg_4(.CP(n_62185), .D(n_35012), .CD(n_61637), .Q(to_acu1
		[4]));
	notech_mux2 i_42094(.S(n_58327), .A(to_acu1[4]), .B(n_40182), .Z(n_35012
		));
	notech_reg to_acu1_reg_5(.CP(n_62185), .D(n_35018), .CD(n_61637), .Q(to_acu1
		[5]));
	notech_mux2 i_42102(.S(n_58327), .A(to_acu1[5]), .B(n_40242), .Z(n_35018
		));
	notech_ao4 i_95473210(.A(n_3053), .B(n_40744), .C(n_3055), .D(n_40792), 
		.Z(n_2162));
	notech_reg to_acu1_reg_6(.CP(n_62185), .D(n_35024), .CD(n_61637), .Q(to_acu1
		[6]));
	notech_mux2 i_42110(.S(n_58327), .A(to_acu1[6]), .B(n_40244), .Z(n_35024
		));
	notech_ao4 i_95573209(.A(n_3052), .B(n_40776), .C(n_3047), .D(n_40784), 
		.Z(n_2161));
	notech_reg to_acu1_reg_7(.CP(n_62185), .D(n_35030), .CD(n_61637), .Q(to_acu1
		[7]));
	notech_mux2 i_42118(.S(n_58337), .A(to_acu1[7]), .B(n_40188), .Z(n_35030
		));
	notech_reg to_acu1_reg_8(.CP(n_62185), .D(n_35036), .CD(n_61637), .Q(to_acu1
		[8]));
	notech_mux2 i_42126(.S(n_58338), .A(to_acu1[8]), .B(n_40246), .Z(n_35036
		));
	notech_ao4 i_957(.A(n_3055), .B(n_40783), .C(n_3052), .D(n_40767), .Z(n_2159
		));
	notech_reg to_acu1_reg_9(.CP(n_62185), .D(n_35042), .CD(n_61637), .Q(to_acu1
		[9]));
	notech_mux2 i_42134(.S(n_58338), .A(to_acu1[9]), .B(n_39376), .Z(n_35042
		));
	notech_reg to_acu1_reg_10(.CP(n_62185), .D(n_35048), .CD(n_61637), .Q(to_acu1
		[10]));
	notech_mux2 i_42142(.S(n_58338), .A(to_acu1[10]), .B(n_39378), .Z(n_35048
		));
	notech_ao4 i_959(.A(n_3046), .B(n_40759), .C(n_40775), .D(n_3047), .Z(n_2157
		));
	notech_reg to_acu1_reg_11(.CP(n_62181), .D(n_35054), .CD(n_61637), .Q(to_acu1
		[11]));
	notech_mux2 i_42150(.S(n_58338), .A(to_acu1[11]), .B(n_39379), .Z(n_35054
		));
	notech_ao4 i_960(.A(n_3045), .B(n_40751), .C(n_40743), .D(n_3048), .Z(n_2156
		));
	notech_reg to_acu1_reg_12(.CP(n_62181), .D(n_35060), .CD(n_61637), .Q(to_acu1
		[12]));
	notech_mux2 i_42158(.S(n_58338), .A(to_acu1[12]), .B(n_39382), .Z(n_35060
		));
	notech_reg to_acu1_reg_13(.CP(n_62181), .D(n_35066), .CD(n_61633), .Q(to_acu1
		[13]));
	notech_mux2 i_42166(.S(n_58338), .A(to_acu1[13]), .B(n_39383), .Z(n_35066
		));
	notech_ao4 i_96273207(.A(n_40733), .B(n_238694343), .C(n_2173), .D(n_40749
		), .Z(n_2154));
	notech_reg to_acu1_reg_14(.CP(n_62185), .D(n_35072), .CD(n_61637), .Q(to_acu1
		[14]));
	notech_mux2 i_42174(.S(n_58338), .A(to_acu1[14]), .B(n_39385), .Z(n_35072
		));
	notech_reg to_acu1_reg_15(.CP(n_62185), .D(n_35078), .CD(n_61633), .Q(to_acu1
		[15]));
	notech_mux2 i_42182(.S(n_58338), .A(to_acu1[15]), .B(n_39386), .Z(n_35078
		));
	notech_reg to_acu1_reg_16(.CP(n_62185), .D(n_35084), .CD(n_61633), .Q(to_acu1
		[16]));
	notech_mux2 i_42190(.S(n_58338), .A(to_acu1[16]), .B(n_39387), .Z(n_35084
		));
	notech_ao4 i_96473205(.A(n_2172), .B(n_40773), .C(n_238794344), .D(n_40781
		), .Z(n_2151));
	notech_reg to_acu1_reg_17(.CP(n_62185), .D(n_35090), .CD(n_61633), .Q(to_acu1
		[17]));
	notech_mux2 i_42198(.S(n_58338), .A(to_acu1[17]), .B(n_39389), .Z(n_35090
		));
	notech_ao4 i_96573204(.A(n_238894345), .B(n_40757), .C(n_238994346), .D(n_40765
		), .Z(n_2150));
	notech_reg to_acu1_reg_18(.CP(n_62185), .D(n_35096), .CD(n_61637), .Q(to_acu1
		[18]));
	notech_mux2 i_42206(.S(n_58338), .A(to_acu1[18]), .B(n_39392), .Z(n_35096
		));
	notech_ao4 i_474154(.A(n_2918), .B(n_40593), .C(n_2944), .D(n_40592), .Z
		(n_2149));
	notech_reg to_acu1_reg_19(.CP(n_62187), .D(n_35102), .CD(n_61637), .Q(to_acu1
		[19]));
	notech_mux2 i_42214(.S(n_58338), .A(to_acu1[19]), .B(n_39395), .Z(n_35102
		));
	notech_reg to_acu1_reg_20(.CP(n_62187), .D(n_35108), .CD(n_61637), .Q(to_acu1
		[20]));
	notech_mux2 i_42222(.S(n_58338), .A(to_acu1[20]), .B(n_39397), .Z(n_35108
		));
	notech_reg to_acu1_reg_21(.CP(n_62187), .D(n_35114), .CD(n_61637), .Q(to_acu1
		[21]));
	notech_mux2 i_42230(.S(n_58337), .A(to_acu1[21]), .B(n_39398), .Z(n_35114
		));
	notech_reg to_acu1_reg_22(.CP(n_62187), .D(n_35120), .CD(n_61637), .Q(to_acu1
		[22]));
	notech_mux2 i_42238(.S(n_58337), .A(to_acu1[22]), .B(n_39399), .Z(n_35120
		));
	notech_reg to_acu1_reg_23(.CP(n_62187), .D(n_35126), .CD(n_61639), .Q(to_acu1
		[23]));
	notech_mux2 i_42246(.S(n_58337), .A(to_acu1[23]), .B(n_39400), .Z(n_35126
		));
	notech_or4 i_2474130(.A(n_40479), .B(n_40490), .C(n_40741), .D(n_1643), 
		.Z(n_2144));
	notech_reg to_acu1_reg_24(.CP(n_62190), .D(n_35132), .CD(n_61639), .Q(to_acu1
		[24]));
	notech_mux2 i_42254(.S(n_58337), .A(to_acu1[24]), .B(n_39401), .Z(n_35132
		));
	notech_reg to_acu1_reg_25(.CP(n_62190), .D(n_35138), .CD(n_61639), .Q(to_acu1
		[25]));
	notech_mux2 i_42262(.S(n_58337), .A(to_acu1[25]), .B(n_39402), .Z(n_35138
		));
	notech_reg to_acu1_reg_26(.CP(n_62190), .D(n_35144), .CD(n_61639), .Q(to_acu1
		[26]));
	notech_mux2 i_42270(.S(n_58337), .A(to_acu1[26]), .B(n_39403), .Z(n_35144
		));
	notech_reg to_acu1_reg_27(.CP(n_62187), .D(n_35150), .CD(n_61639), .Q(to_acu1
		[27]));
	notech_mux2 i_42278(.S(n_58337), .A(to_acu1[27]), .B(n_39404), .Z(n_35150
		));
	notech_reg to_acu1_reg_28(.CP(n_62187), .D(n_35156), .CD(n_61642), .Q(to_acu1
		[28]));
	notech_mux2 i_42286(.S(n_58337), .A(to_acu1[28]), .B(n_39405), .Z(n_35156
		));
	notech_reg to_acu1_reg_29(.CP(n_62187), .D(n_35162), .CD(n_61642), .Q(to_acu1
		[29]));
	notech_mux2 i_42294(.S(n_58337), .A(to_acu1[29]), .B(n_39406), .Z(n_35162
		));
	notech_reg to_acu1_reg_30(.CP(n_62187), .D(n_35168), .CD(n_61639), .Q(to_acu1
		[30]));
	notech_mux2 i_42302(.S(n_58337), .A(to_acu1[30]), .B(n_39407), .Z(n_35168
		));
	notech_or2 i_2274132(.A(n_3053), .B(n_40735), .Z(n_2137));
	notech_reg to_acu1_reg_31(.CP(n_62187), .D(n_35174), .CD(n_61639), .Q(to_acu1
		[31]));
	notech_mux2 i_42310(.S(n_58337), .A(to_acu1[31]), .B(n_39408), .Z(n_35174
		));
	notech_reg to_acu1_reg_32(.CP(n_62187), .D(n_35180), .CD(n_61639), .Q(to_acu1
		[32]));
	notech_mux2 i_42318(.S(n_58337), .A(to_acu1[32]), .B(n_39409), .Z(n_35180
		));
	notech_reg to_acu1_reg_33(.CP(n_62187), .D(n_35186), .CD(n_61639), .Q(to_acu1
		[33]));
	notech_mux2 i_42326(.S(n_58337), .A(to_acu1[33]), .B(n_39411), .Z(n_35186
		));
	notech_reg to_acu1_reg_34(.CP(n_62187), .D(n_35192), .CD(n_61639), .Q(to_acu1
		[34]));
	notech_mux2 i_42334(.S(n_58269), .A(to_acu1[34]), .B(n_39414), .Z(n_35192
		));
	notech_reg to_acu1_reg_35(.CP(n_62187), .D(n_35198), .CD(n_61639), .Q(to_acu1
		[35]));
	notech_mux2 i_42342(.S(n_58269), .A(to_acu1[35]), .B(n_39416), .Z(n_35198
		));
	notech_reg to_acu1_reg_36(.CP(n_62187), .D(n_35204), .CD(n_61639), .Q(to_acu1
		[36]));
	notech_mux2 i_42350(.S(n_58269), .A(to_acu1[36]), .B(n_39421), .Z(n_35204
		));
	notech_reg to_acu1_reg_37(.CP(n_62187), .D(n_35210), .CD(n_61637), .Q(to_acu1
		[37]));
	notech_mux2 i_42358(.S(n_58269), .A(to_acu1[37]), .B(n_39424), .Z(n_35210
		));
	notech_or2 i_2374131(.A(n_253194488), .B(n_40752), .Z(n_2130));
	notech_reg to_acu1_reg_38(.CP(n_62187), .D(n_35216), .CD(n_61639), .Q(to_acu1
		[38]));
	notech_mux2 i_42366(.S(n_58269), .A(to_acu1[38]), .B(n_39427), .Z(n_35216
		));
	notech_reg to_acu1_reg_39(.CP(n_62187), .D(n_35222), .CD(n_61639), .Q(to_acu1
		[39]));
	notech_mux2 i_42374(.S(n_58269), .A(to_acu1[39]), .B(n_160996304), .Z(n_35222
		));
	notech_reg to_acu1_reg_40(.CP(n_62181), .D(n_35228), .CD(n_61639), .Q(to_acu1
		[40]));
	notech_mux2 i_42382(.S(n_58270), .A(to_acu1[40]), .B(n_39430), .Z(n_35228
		));
	notech_nor2 i_3779(.A(n_1644), .B(fpu), .Z(n_44046));
	notech_reg to_acu1_reg_41(.CP(n_62179), .D(n_35234), .CD(n_61639), .Q(to_acu1
		[41]));
	notech_mux2 i_42390(.S(n_58270), .A(to_acu1[41]), .B(n_39433), .Z(n_35234
		));
	notech_ao3 i_3315(.A(n_59969), .B(udeco[21]), .C(n_59657), .Z(n_43318)
		);
	notech_reg to_acu1_reg_42(.CP(n_62179), .D(n_35240), .CD(n_61639), .Q(to_acu1
		[42]));
	notech_mux2 i_42398(.S(n_58270), .A(to_acu1[42]), .B(n_39436), .Z(n_35240
		));
	notech_ao3 i_3313(.A(n_59969), .B(udeco[19]), .C(n_59657), .Z(n_43306)
		);
	notech_reg to_acu1_reg_43(.CP(n_62179), .D(n_35246), .CD(n_61639), .Q(to_acu1
		[43]));
	notech_mux2 i_42406(.S(n_58270), .A(to_acu1[43]), .B(n_39439), .Z(n_35246
		));
	notech_ao3 i_3311(.A(n_59969), .B(udeco[17]), .C(n_59653), .Z(n_43294)
		);
	notech_reg to_acu1_reg_44(.CP(n_62179), .D(n_35252), .CD(n_61631), .Q(to_acu1
		[44]));
	notech_mux2 i_42414(.S(n_58270), .A(to_acu1[44]), .B(n_39442), .Z(n_35252
		));
	notech_ao3 i_3309(.A(n_59969), .B(udeco[15]), .C(n_59653), .Z(n_43282)
		);
	notech_reg to_acu1_reg_45(.CP(n_62179), .D(n_35258), .CD(n_61631), .Q(to_acu1
		[45]));
	notech_mux2 i_42422(.S(n_58270), .A(to_acu1[45]), .B(n_39445), .Z(n_35258
		));
	notech_ao3 i_3308(.A(n_59975), .B(udeco[14]), .C(n_59657), .Z(n_43276)
		);
	notech_reg to_acu1_reg_46(.CP(n_62179), .D(n_35264), .CD(n_61631), .Q(to_acu1
		[46]));
	notech_mux2 i_42430(.S(n_58270), .A(to_acu1[46]), .B(n_39448), .Z(n_35264
		));
	notech_ao3 i_3307(.A(n_59980), .B(udeco[13]), .C(n_59657), .Z(n_43270)
		);
	notech_reg to_acu1_reg_47(.CP(n_62179), .D(n_35270), .CD(n_61631), .Q(to_acu1
		[47]));
	notech_mux2 i_42438(.S(n_58269), .A(to_acu1[47]), .B(n_39451), .Z(n_35270
		));
	notech_ao3 i_3305(.A(n_59980), .B(udeco[11]), .C(n_59657), .Z(n_43258)
		);
	notech_reg to_acu1_reg_48(.CP(n_62179), .D(n_35276), .CD(n_61631), .Q(to_acu1
		[48]));
	notech_mux2 i_42446(.S(n_58269), .A(to_acu1[48]), .B(n_39454), .Z(n_35276
		));
	notech_ao3 i_3304(.A(n_59980), .B(udeco[10]), .C(n_59657), .Z(n_43252)
		);
	notech_reg to_acu1_reg_49(.CP(n_62179), .D(n_35282), .CD(n_61631), .Q(to_acu1
		[49]));
	notech_mux2 i_42454(.S(n_58269), .A(to_acu1[49]), .B(n_39457), .Z(n_35282
		));
	notech_ao3 i_3303(.A(n_59980), .B(udeco[9]), .C(n_59657), .Z(n_43246));
	notech_reg to_acu1_reg_50(.CP(n_62179), .D(n_35288), .CD(n_61631), .Q(to_acu1
		[50]));
	notech_mux2 i_42462(.S(n_58264), .A(to_acu1[50]), .B(n_39460), .Z(n_35288
		));
	notech_ao3 i_3302(.A(n_59980), .B(udeco[8]), .C(n_59657), .Z(n_43240));
	notech_reg to_acu1_reg_51(.CP(n_62179), .D(n_35294), .CD(n_61631), .Q(to_acu1
		[51]));
	notech_mux2 i_42470(.S(n_58269), .A(to_acu1[51]), .B(n_39463), .Z(n_35294
		));
	notech_ao3 i_3301(.A(n_59980), .B(udeco[7]), .C(n_59653), .Z(n_43234));
	notech_reg to_acu1_reg_52(.CP(n_62176), .D(n_35300), .CD(n_61631), .Q(to_acu1
		[52]));
	notech_mux2 i_42478(.S(n_58269), .A(to_acu1[52]), .B(n_39466), .Z(n_35300
		));
	notech_ao3 i_3300(.A(n_59980), .B(udeco[6]), .C(n_59653), .Z(n_43228));
	notech_reg to_acu1_reg_53(.CP(n_62176), .D(n_35306), .CD(n_61631), .Q(to_acu1
		[53]));
	notech_mux2 i_42486(.S(n_58269), .A(to_acu1[53]), .B(n_39469), .Z(n_35306
		));
	notech_ao3 i_3299(.A(n_59980), .B(udeco[5]), .C(n_59653), .Z(n_43222));
	notech_reg to_acu1_reg_54(.CP(n_62176), .D(n_35312), .CD(n_61631), .Q(to_acu1
		[54]));
	notech_mux2 i_42494(.S(n_58269), .A(to_acu1[54]), .B(n_39472), .Z(n_35312
		));
	notech_ao3 i_3298(.A(n_59980), .B(udeco[4]), .C(n_59653), .Z(n_43216));
	notech_reg to_acu1_reg_55(.CP(n_62176), .D(n_35318), .CD(n_61628), .Q(to_acu1
		[55]));
	notech_mux2 i_42502(.S(n_58269), .A(to_acu1[55]), .B(n_39475), .Z(n_35318
		));
	notech_ao3 i_3297(.A(n_59980), .B(udeco[3]), .C(n_59653), .Z(n_43210));
	notech_reg to_acu1_reg_56(.CP(n_62176), .D(n_35324), .CD(n_61628), .Q(to_acu1
		[56]));
	notech_mux2 i_42510(.S(n_58269), .A(to_acu1[56]), .B(n_39478), .Z(n_35324
		));
	notech_ao3 i_3296(.A(n_59980), .B(udeco[2]), .C(n_59653), .Z(n_43204));
	notech_reg to_acu1_reg_57(.CP(n_62176), .D(n_35330), .CD(n_61628), .Q(to_acu1
		[57]));
	notech_mux2 i_42518(.S(n_58269), .A(to_acu1[57]), .B(n_39481), .Z(n_35330
		));
	notech_ao3 i_3295(.A(n_59980), .B(udeco[1]), .C(n_59653), .Z(n_43198));
	notech_reg to_acu1_reg_58(.CP(n_62176), .D(n_35336), .CD(n_61628), .Q(to_acu1
		[58]));
	notech_mux2 i_42526(.S(n_58269), .A(to_acu1[58]), .B(n_39484), .Z(n_35336
		));
	notech_ao3 i_3294(.A(n_59980), .B(udeco[0]), .C(n_59653), .Z(n_43192));
	notech_reg to_acu1_reg_59(.CP(n_62176), .D(n_35342), .CD(n_61628), .Q(to_acu1
		[59]));
	notech_mux2 i_42534(.S(n_58269), .A(to_acu1[59]), .B(n_39487), .Z(n_35342
		));
	notech_ao3 i_11774037(.A(n_59975), .B(in128[124]), .C(n_59653), .Z(n_48380
		));
	notech_reg to_acu1_reg_60(.CP(n_62176), .D(n_35348), .CD(n_61628), .Q(to_acu1
		[60]));
	notech_mux2 i_42542(.S(n_58270), .A(to_acu1[60]), .B(n_39490), .Z(n_35348
		));
	notech_ao3 i_11974035(.A(n_59975), .B(in128[122]), .C(n_59653), .Z(n_48368
		));
	notech_reg to_acu1_reg_61(.CP(n_62176), .D(n_35354), .CD(n_61628), .Q(to_acu1
		[61]));
	notech_mux2 i_42550(.S(n_58253), .A(to_acu1[61]), .B(n_39493), .Z(n_35354
		));
	notech_and2 i_72573439(.A(n_2168), .B(n_225896451), .Z(n_2127));
	notech_reg to_acu1_reg_62(.CP(n_62181), .D(n_35360), .CD(n_61628), .Q(to_acu1
		[62]));
	notech_mux2 i_42558(.S(n_58253), .A(to_acu1[62]), .B(n_39496), .Z(n_35360
		));
	notech_and4 i_72473440(.A(n_2154), .B(n_2151), .C(n_2150), .D(n_2144), .Z
		(n_2126));
	notech_reg to_acu1_reg_63(.CP(n_62181), .D(n_35366), .CD(n_61628), .Q(to_acu1
		[63]));
	notech_mux2 i_42566(.S(n_58253), .A(to_acu1[63]), .B(n_39499), .Z(n_35366
		));
	notech_and4 i_72373441(.A(n_2159), .B(n_2157), .C(n_2156), .D(n_2137), .Z
		(n_2125));
	notech_reg to_acu1_reg_64(.CP(n_62181), .D(n_35372), .CD(n_61628), .Q(to_acu1
		[64]));
	notech_mux2 i_42574(.S(n_58253), .A(to_acu1[64]), .B(n_39502), .Z(n_35372
		));
	notech_reg to_acu1_reg_65(.CP(n_62181), .D(n_35378), .CD(n_61633), .Q(to_acu1
		[65]));
	notech_mux2 i_42582(.S(n_58253), .A(to_acu1[65]), .B(n_39505), .Z(n_35378
		));
	notech_ao4 i_72273442(.A(n_40593), .B(n_2918), .C(n_254394500), .D(n_40534
		), .Z(n_2123));
	notech_reg to_acu1_reg_66(.CP(n_62181), .D(n_35384), .CD(n_61633), .Q(to_acu1
		[66]));
	notech_mux2 i_42590(.S(n_58253), .A(to_acu1[66]), .B(n_39508), .Z(n_35384
		));
	notech_and4 i_72173443(.A(n_2130), .B(n_2164), .C(n_2162), .D(n_2161), .Z
		(n_2122));
	notech_reg to_acu1_reg_67(.CP(n_62181), .D(n_35390), .CD(n_61633), .Q(to_acu1
		[67]));
	notech_mux2 i_42598(.S(n_58253), .A(to_acu1[67]), .B(n_39511), .Z(n_35390
		));
	notech_reg to_acu1_reg_68(.CP(n_62181), .D(n_35396), .CD(n_61633), .Q(to_acu1
		[68]));
	notech_mux2 i_42606(.S(n_58280), .A(to_acu1[68]), .B(n_39514), .Z(n_35396
		));
	notech_reg to_acu1_reg_69(.CP(n_62181), .D(n_35402), .CD(n_61633), .Q(to_acu1
		[69]));
	notech_mux2 i_42614(.S(n_58280), .A(to_acu1[69]), .B(n_39517), .Z(n_35402
		));
	notech_ao4 i_72073444(.A(n_40760), .B(n_40491), .C(n_40489), .D(n_40768)
		, .Z(n_2119));
	notech_reg to_acu1_reg_70(.CP(n_62181), .D(n_35408), .CD(n_61633), .Q(to_acu1
		[70]));
	notech_mux2 i_42622(.S(n_58280), .A(to_acu1[70]), .B(n_39520), .Z(n_35408
		));
	notech_reg to_acu1_reg_71(.CP(n_62181), .D(n_35414), .CD(n_61633), .Q(to_acu1
		[71]));
	notech_mux2 i_42630(.S(n_58253), .A(to_acu1[71]), .B(n_39523), .Z(n_35414
		));
	notech_reg to_acu1_reg_72(.CP(n_62181), .D(n_35420), .CD(n_61633), .Q(to_acu1
		[72]));
	notech_mux2 i_42638(.S(n_58253), .A(to_acu1[72]), .B(n_39526), .Z(n_35420
		));
	notech_ao4 i_71973445(.A(n_40764), .B(n_40491), .C(n_40772), .D(n_40489)
		, .Z(n_2116));
	notech_reg to_acu1_reg_73(.CP(n_62179), .D(n_35426), .CD(n_61633), .Q(to_acu1
		[73]));
	notech_mux2 i_42646(.S(n_58280), .A(to_acu1[73]), .B(n_39529), .Z(n_35426
		));
	notech_reg to_acu1_reg_74(.CP(n_62179), .D(n_35432), .CD(n_61633), .Q(to_acu1
		[74]));
	notech_mux2 i_42654(.S(n_58270), .A(to_acu1[74]), .B(n_39532), .Z(n_35432
		));
	notech_reg to_acu1_reg_75(.CP(n_62179), .D(n_35438), .CD(n_61633), .Q(to_acu1
		[75]));
	notech_mux2 i_42662(.S(n_58270), .A(to_acu1[75]), .B(n_39535), .Z(n_35438
		));
	notech_reg to_acu1_reg_76(.CP(n_62179), .D(n_35444), .CD(n_61631), .Q(to_acu1
		[76]));
	notech_mux2 i_42670(.S(n_58270), .A(to_acu1[76]), .B(n_39538), .Z(n_35444
		));
	notech_reg to_acu1_reg_77(.CP(n_62179), .D(n_35450), .CD(n_61631), .Q(to_acu1
		[77]));
	notech_mux2 i_42678(.S(n_58270), .A(to_acu1[77]), .B(n_39541), .Z(n_35450
		));
	notech_reg to_acu1_reg_78(.CP(n_62181), .D(n_35456), .CD(n_61631), .Q(to_acu1
		[78]));
	notech_mux2 i_42686(.S(n_58270), .A(to_acu1[78]), .B(n_39544), .Z(n_35456
		));
	notech_reg to_acu1_reg_79(.CP(n_62181), .D(n_35462), .CD(n_61631), .Q(to_acu1
		[79]));
	notech_mux2 i_42694(.S(n_58270), .A(to_acu1[79]), .B(n_39547), .Z(n_35462
		));
	notech_reg to_acu1_reg_80(.CP(n_62181), .D(n_35468), .CD(n_61631), .Q(to_acu1
		[80]));
	notech_mux2 i_42702(.S(n_58270), .A(to_acu1[80]), .B(n_39550), .Z(n_35468
		));
	notech_reg to_acu1_reg_81(.CP(n_62179), .D(n_35474), .CD(n_61633), .Q(to_acu1
		[81]));
	notech_mux2 i_42710(.S(n_58253), .A(to_acu1[81]), .B(n_39553), .Z(n_35474
		));
	notech_reg to_acu1_reg_82(.CP(n_62179), .D(n_35480), .CD(n_61633), .Q(to_acu1
		[82]));
	notech_mux2 i_42718(.S(n_58253), .A(to_acu1[82]), .B(n_39556), .Z(n_35480
		));
	notech_reg to_acu1_reg_83(.CP(n_62197), .D(n_35486), .CD(n_61633), .Q(to_acu1
		[83]));
	notech_mux2 i_42726(.S(n_58253), .A(to_acu1[83]), .B(n_39559), .Z(n_35486
		));
	notech_reg to_acu1_reg_84(.CP(n_62197), .D(n_35492), .CD(n_61631), .Q(to_acu1
		[84]));
	notech_mux2 i_42734(.S(n_58270), .A(to_acu1[84]), .B(n_40302), .Z(n_35492
		));
	notech_reg to_acu1_reg_85(.CP(n_62197), .D(n_35498), .CD(n_61631), .Q(to_acu1
		[85]));
	notech_mux2 i_42742(.S(n_58270), .A(to_acu1[85]), .B(n_39562), .Z(n_35498
		));
	notech_reg to_acu1_reg_86(.CP(n_62197), .D(n_35504), .CD(n_61642), .Q(to_acu1
		[86]));
	notech_mux2 i_42750(.S(n_58270), .A(to_acu1[86]), .B(n_39565), .Z(n_35504
		));
	notech_reg to_acu1_reg_87(.CP(n_62197), .D(n_35510), .CD(n_61649), .Q(to_acu1
		[87]));
	notech_mux2 i_42758(.S(n_58258), .A(to_acu1[87]), .B(n_39568), .Z(n_35510
		));
	notech_reg to_acu1_reg_88(.CP(n_62197), .D(n_35516), .CD(n_61649), .Q(to_acu1
		[88]));
	notech_mux2 i_42766(.S(n_58258), .A(to_acu1[88]), .B(n_39571), .Z(n_35516
		));
	notech_reg to_acu1_reg_89(.CP(n_62197), .D(n_35522), .CD(n_61649), .Q(to_acu1
		[89]));
	notech_mux2 i_42774(.S(n_58258), .A(to_acu1[89]), .B(n_39574), .Z(n_35522
		));
	notech_reg to_acu1_reg_90(.CP(n_62197), .D(n_35528), .CD(n_61649), .Q(to_acu1
		[90]));
	notech_mux2 i_42782(.S(n_58258), .A(to_acu1[90]), .B(n_40313), .Z(n_35528
		));
	notech_reg to_acu1_reg_91(.CP(n_62197), .D(n_35534), .CD(n_61649), .Q(to_acu1
		[91]));
	notech_mux2 i_42790(.S(n_58258), .A(to_acu1[91]), .B(n_40315), .Z(n_35534
		));
	notech_reg to_acu1_reg_92(.CP(n_62197), .D(n_35540), .CD(n_61649), .Q(to_acu1
		[92]));
	notech_mux2 i_42798(.S(n_58258), .A(to_acu1[92]), .B(n_40317), .Z(n_35540
		));
	notech_reg to_acu1_reg_93(.CP(n_62197), .D(n_35546), .CD(n_61649), .Q(to_acu1
		[93]));
	notech_mux2 i_42806(.S(n_58258), .A(to_acu1[93]), .B(n_40320), .Z(n_35546
		));
	notech_reg to_acu1_reg_94(.CP(n_62195), .D(n_35552), .CD(n_61649), .Q(to_acu1
		[94]));
	notech_mux2 i_42814(.S(n_58258), .A(to_acu1[94]), .B(n_40322), .Z(n_35552
		));
	notech_reg to_acu1_reg_95(.CP(n_62195), .D(n_35558), .CD(n_61649), .Q(to_acu1
		[95]));
	notech_mux2 i_42822(.S(n_58258), .A(to_acu1[95]), .B(n_40324), .Z(n_35558
		));
	notech_reg to_acu1_reg_96(.CP(n_62195), .D(n_35564), .CD(n_61649), .Q(to_acu1
		[96]));
	notech_mux2 i_42830(.S(n_58259), .A(to_acu1[96]), .B(n_40327), .Z(n_35564
		));
	notech_reg to_acu1_reg_97(.CP(n_62195), .D(n_35570), .CD(n_61649), .Q(to_acu1
		[97]));
	notech_mux2 i_42838(.S(n_58258), .A(to_acu1[97]), .B(n_40329), .Z(n_35570
		));
	notech_reg to_acu1_reg_98(.CP(n_62195), .D(n_35576), .CD(n_61647), .Q(to_acu1
		[98]));
	notech_mux2 i_42846(.S(n_58258), .A(to_acu1[98]), .B(n_40331), .Z(n_35576
		));
	notech_reg to_acu1_reg_99(.CP(n_62197), .D(n_35582), .CD(n_61647), .Q(to_acu1
		[99]));
	notech_mux2 i_42854(.S(n_58258), .A(to_acu1[99]), .B(n_40333), .Z(n_35582
		));
	notech_reg to_acu1_reg_100(.CP(n_62197), .D(n_35588), .CD(n_61647), .Q(to_acu1
		[100]));
	notech_mux2 i_42862(.S(n_58253), .A(to_acu1[100]), .B(n_40335), .Z(n_35588
		));
	notech_reg to_acu1_reg_101(.CP(n_62195), .D(n_35594), .CD(n_61647), .Q(to_acu1
		[101]));
	notech_mux2 i_42870(.S(n_58253), .A(to_acu1[101]), .B(n_40337), .Z(n_35594
		));
	notech_reg to_acu1_reg_102(.CP(n_62195), .D(n_35600), .CD(n_61647), .Q(to_acu1
		[102]));
	notech_mux2 i_42878(.S(n_58258), .A(to_acu1[102]), .B(n_40339), .Z(n_35600
		));
	notech_reg to_acu1_reg_103(.CP(n_62195), .D(n_35606), .CD(n_61647), .Q(to_acu1
		[103]));
	notech_mux2 i_42886(.S(n_58253), .A(to_acu1[103]), .B(n_40341), .Z(n_35606
		));
	notech_reg to_acu1_reg_104(.CP(n_62201), .D(n_35612), .CD(n_61649), .Q(to_acu1
		[104]));
	notech_mux2 i_42894(.S(n_58253), .A(to_acu1[104]), .B(n_40343), .Z(n_35612
		));
	notech_reg to_acu1_reg_105(.CP(n_62201), .D(n_35618), .CD(n_61647), .Q(to_acu1
		[105]));
	notech_mux2 i_42902(.S(n_58253), .A(to_acu1[105]), .B(n_40345), .Z(n_35618
		));
	notech_reg to_acu1_reg_106(.CP(n_62201), .D(n_35624), .CD(n_61647), .Q(to_acu1
		[106]));
	notech_mux2 i_42910(.S(n_58258), .A(to_acu1[106]), .B(n_40347), .Z(n_35624
		));
	notech_reg to_acu1_reg_107(.CP(n_62201), .D(n_35630), .CD(n_61647), .Q(to_acu1
		[107]));
	notech_mux2 i_42918(.S(n_58258), .A(to_acu1[107]), .B(n_39578), .Z(n_35630
		));
	notech_reg to_acu1_reg_108(.CP(n_62201), .D(n_35636), .CD(n_61653), .Q(to_acu1
		[108]));
	notech_mux2 i_42926(.S(n_58258), .A(to_acu1[108]), .B(n_40350), .Z(n_35636
		));
	notech_reg to_acu1_reg_109(.CP(n_62201), .D(n_35642), .CD(n_61653), .Q(to_acu1
		[109]));
	notech_mux2 i_42934(.S(n_58258), .A(to_acu1[109]), .B(n_39581), .Z(n_35642
		));
	notech_reg to_acu1_reg_110(.CP(n_62201), .D(n_35648), .CD(n_61653), .Q(to_acu1
		[110]));
	notech_mux2 i_42942(.S(n_58258), .A(to_acu1[110]), .B(n_39584), .Z(n_35648
		));
	notech_reg to_acu1_reg_111(.CP(n_62201), .D(n_35654), .CD(n_61653), .Q(to_acu1
		[111]));
	notech_mux2 i_42950(.S(n_58258), .A(to_acu1[111]), .B(n_39587), .Z(n_35654
		));
	notech_reg to_acu1_reg_112(.CP(n_62201), .D(n_35660), .CD(n_61653), .Q(to_acu1
		[112]));
	notech_mux2 i_42958(.S(n_58258), .A(to_acu1[112]), .B(n_39590), .Z(n_35660
		));
	notech_reg to_acu1_reg_113(.CP(n_62201), .D(n_35666), .CD(n_61653), .Q(to_acu1
		[113]));
	notech_mux2 i_42966(.S(n_58259), .A(to_acu1[113]), .B(n_39593), .Z(n_35666
		));
	notech_reg to_acu1_reg_114(.CP(n_62201), .D(n_35672), .CD(n_61653), .Q(to_acu1
		[114]));
	notech_mux2 i_42974(.S(n_58264), .A(to_acu1[114]), .B(n_40357), .Z(n_35672
		));
	notech_reg to_acu1_reg_115(.CP(n_62197), .D(n_35678), .CD(n_61653), .Q(to_acu1
		[115]));
	notech_mux2 i_42982(.S(n_58264), .A(to_acu1[115]), .B(n_40359), .Z(n_35678
		));
	notech_reg to_acu1_reg_116(.CP(n_62197), .D(n_35684), .CD(n_61653), .Q(to_acu1
		[116]));
	notech_mux2 i_42990(.S(n_58264), .A(to_acu1[116]), .B(n_40361), .Z(n_35684
		));
	notech_reg to_acu1_reg_117(.CP(n_62197), .D(n_35690), .CD(n_61653), .Q(to_acu1
		[117]));
	notech_mux2 i_42998(.S(n_58259), .A(to_acu1[117]), .B(n_40363), .Z(n_35690
		));
	notech_reg to_acu1_reg_118(.CP(n_62197), .D(n_35696), .CD(n_61653), .Q(to_acu1
		[118]));
	notech_mux2 i_43006(.S(n_58259), .A(to_acu1[118]), .B(n_40365), .Z(n_35696
		));
	notech_reg to_acu1_reg_119(.CP(n_62197), .D(n_35702), .CD(n_61649), .Q(to_acu1
		[119]));
	notech_mux2 i_43014(.S(n_58264), .A(to_acu1[119]), .B(n_39596), .Z(n_35702
		));
	notech_reg to_acu1_reg_120(.CP(n_62201), .D(n_35708), .CD(n_61649), .Q(to_acu1
		[120]));
	notech_mux2 i_43022(.S(n_58264), .A(to_acu1[120]), .B(n_40368), .Z(n_35708
		));
	notech_reg to_acu1_reg_121(.CP(n_62201), .D(n_35714), .CD(n_61649), .Q(to_acu1
		[121]));
	notech_mux2 i_43030(.S(n_58264), .A(to_acu1[121]), .B(n_39599), .Z(n_35714
		));
	notech_reg to_acu1_reg_122(.CP(n_62201), .D(n_35720), .CD(n_61649), .Q(to_acu1
		[122]));
	notech_mux2 i_43038(.S(n_58264), .A(to_acu1[122]), .B(n_39602), .Z(n_35720
		));
	notech_reg to_acu1_reg_123(.CP(n_62201), .D(n_35726), .CD(n_61649), .Q(to_acu1
		[123]));
	notech_mux2 i_43046(.S(n_58264), .A(to_acu1[123]), .B(n_39605), .Z(n_35726
		));
	notech_reg to_acu1_reg_124(.CP(n_62201), .D(n_35732), .CD(n_61653), .Q(to_acu1
		[124]));
	notech_mux2 i_43054(.S(n_58264), .A(to_acu1[124]), .B(n_40373), .Z(n_35732
		));
	notech_reg to_acu1_reg_125(.CP(n_62195), .D(n_35738), .CD(n_61653), .Q(to_acu1
		[125]));
	notech_mux2 i_43062(.S(n_58264), .A(to_acu1[125]), .B(n_39608), .Z(n_35738
		));
	notech_reg to_acu1_reg_126(.CP(n_62190), .D(n_35744), .CD(n_61653), .Q(to_acu1
		[126]));
	notech_mux2 i_43070(.S(n_58264), .A(to_acu1[126]), .B(n_39611), .Z(n_35744
		));
	notech_reg to_acu1_reg_127(.CP(n_62192), .D(n_35750), .CD(n_61649), .Q(to_acu1
		[127]));
	notech_mux2 i_43078(.S(n_58259), .A(to_acu1[127]), .B(n_39614), .Z(n_35750
		));
	notech_reg to_acu1_reg_128(.CP(n_62190), .D(n_35756), .CD(n_61653), .Q(to_acu1
		[128]));
	notech_mux2 i_43086(.S(n_58259), .A(to_acu1[128]), .B(n_39616), .Z(n_35756
		));
	notech_reg to_acu1_reg_129(.CP(n_62190), .D(n_35762), .CD(n_61642), .Q(to_acu1
		[129]));
	notech_mux2 i_43094(.S(n_58259), .A(to_acu1[129]), .B(n_39618), .Z(n_35762
		));
	notech_reg to_acu1_reg_130(.CP(n_62190), .D(n_35768), .CD(n_61644), .Q(to_acu1
		[130]));
	notech_mux2 i_43102(.S(n_58259), .A(to_acu1[130]), .B(n_39620), .Z(n_35768
		));
	notech_reg to_acu1_reg_131(.CP(n_62192), .D(n_35774), .CD(n_61642), .Q(to_acu1
		[131]));
	notech_mux2 i_43110(.S(n_58259), .A(to_acu1[131]), .B(n_39622), .Z(n_35774
		));
	notech_reg to_acu1_reg_132(.CP(n_62192), .D(n_35780), .CD(n_61642), .Q(to_acu1
		[132]));
	notech_mux2 i_43118(.S(n_58259), .A(to_acu1[132]), .B(n_39624), .Z(n_35780
		));
	notech_reg to_acu1_reg_133(.CP(n_62192), .D(n_35786), .CD(n_61642), .Q(to_acu1
		[133]));
	notech_mux2 i_43126(.S(n_58259), .A(to_acu1[133]), .B(n_39626), .Z(n_35786
		));
	notech_reg to_acu1_reg_134(.CP(n_62192), .D(n_35792), .CD(n_61644), .Q(to_acu1
		[134]));
	notech_mux2 i_43134(.S(n_58259), .A(to_acu1[134]), .B(n_39628), .Z(n_35792
		));
	notech_reg to_acu1_reg_135(.CP(n_62192), .D(n_35798), .CD(n_61644), .Q(to_acu1
		[135]));
	notech_mux2 i_43142(.S(n_58259), .A(to_acu1[135]), .B(n_39630), .Z(n_35798
		));
	notech_reg to_acu1_reg_136(.CP(n_62190), .D(n_35804), .CD(n_61644), .Q(to_acu1
		[136]));
	notech_mux2 i_43150(.S(n_58259), .A(to_acu1[136]), .B(n_39632), .Z(n_35804
		));
	notech_reg to_acu1_reg_137(.CP(n_62190), .D(n_35810), .CD(n_61644), .Q(to_acu1
		[137]));
	notech_mux2 i_43158(.S(n_58259), .A(to_acu1[137]), .B(n_39634), .Z(n_35810
		));
	notech_reg to_acu1_reg_138(.CP(n_62190), .D(n_35816), .CD(n_61644), .Q(to_acu1
		[138]));
	notech_mux2 i_43166(.S(n_58259), .A(to_acu1[138]), .B(n_39636), .Z(n_35816
		));
	notech_reg to_acu1_reg_139(.CP(n_62190), .D(n_35822), .CD(n_61642), .Q(to_acu1
		[139]));
	notech_mux2 i_43174(.S(n_58259), .A(to_acu1[139]), .B(n_39638), .Z(n_35822
		));
	notech_reg to_acu1_reg_140(.CP(n_62190), .D(n_35828), .CD(n_61642), .Q(to_acu1
		[140]));
	notech_mux2 i_43182(.S(n_58280), .A(to_acu1[140]), .B(n_39640), .Z(n_35828
		));
	notech_reg to_acu1_reg_141(.CP(n_62190), .D(n_35834), .CD(n_61642), .Q(to_acu1
		[141]));
	notech_mux2 i_43190(.S(n_58293), .A(to_acu1[141]), .B(n_39642), .Z(n_35834
		));
	notech_reg to_acu1_reg_142(.CP(n_62190), .D(n_35840), .CD(n_61642), .Q(to_acu1
		[142]));
	notech_mux2 i_43198(.S(n_58293), .A(to_acu1[142]), .B(n_39644), .Z(n_35840
		));
	notech_reg to_acu1_reg_143(.CP(n_62190), .D(n_35846), .CD(n_61642), .Q(to_acu1
		[143]));
	notech_mux2 i_43206(.S(n_58293), .A(to_acu1[143]), .B(n_39646), .Z(n_35846
		));
	notech_reg to_acu1_reg_144(.CP(n_62190), .D(n_35852), .CD(n_61642), .Q(to_acu1
		[144]));
	notech_mux2 i_43214(.S(n_58293), .A(to_acu1[144]), .B(n_39648), .Z(n_35852
		));
	notech_reg to_acu1_reg_145(.CP(n_62190), .D(n_35858), .CD(n_61642), .Q(to_acu1
		[145]));
	notech_mux2 i_43222(.S(n_58293), .A(to_acu1[145]), .B(n_39650), .Z(n_35858
		));
	notech_reg to_acu1_reg_146(.CP(n_62190), .D(n_35864), .CD(n_61642), .Q(to_acu1
		[146]));
	notech_mux2 i_43230(.S(n_58293), .A(to_acu1[146]), .B(n_39653), .Z(n_35864
		));
	notech_reg to_acu1_reg_147(.CP(n_62195), .D(n_35870), .CD(n_61642), .Q(to_acu1
		[147]));
	notech_mux2 i_43238(.S(n_58293), .A(to_acu1[147]), .B(n_39655), .Z(n_35870
		));
	notech_reg to_acu1_reg_148(.CP(n_62195), .D(n_35876), .CD(n_61642), .Q(to_acu1
		[148]));
	notech_mux2 i_43246(.S(n_58293), .A(to_acu1[148]), .B(n_39657), .Z(n_35876
		));
	notech_reg to_acu1_reg_149(.CP(n_62195), .D(n_35882), .CD(n_61642), .Q(to_acu1
		[149]));
	notech_mux2 i_43254(.S(n_58293), .A(to_acu1[149]), .B(n_39661), .Z(n_35882
		));
	notech_reg to_acu1_reg_150(.CP(n_62192), .D(n_35888), .CD(n_61647), .Q(to_acu1
		[150]));
	notech_mux2 i_43262(.S(n_58293), .A(to_acu1[150]), .B(n_40400), .Z(n_35888
		));
	notech_reg to_acu1_reg_151(.CP(n_62195), .D(n_35894), .CD(n_61647), .Q(to_acu1
		[151]));
	notech_mux2 i_43270(.S(n_58293), .A(to_acu1[151]), .B(n_40402), .Z(n_35894
		));
	notech_reg to_acu1_reg_152(.CP(n_62195), .D(n_35900), .CD(n_61647), .Q(to_acu1
		[152]));
	notech_mux2 i_43278(.S(n_58293), .A(to_acu1[152]), .B(n_40404), .Z(n_35900
		));
	notech_reg to_acu1_reg_153(.CP(n_62195), .D(n_35906), .CD(n_61644), .Q(to_acu1
		[153]));
	notech_mux2 i_43286(.S(n_58293), .A(to_acu1[153]), .B(n_39666), .Z(n_35906
		));
	notech_reg to_acu1_reg_154(.CP(n_62195), .D(n_35912), .CD(n_61647), .Q(to_acu1
		[154]));
	notech_mux2 i_43294(.S(n_58292), .A(to_acu1[154]), .B(n_39669), .Z(n_35912
		));
	notech_reg to_acu1_reg_155(.CP(n_62195), .D(n_35918), .CD(n_61647), .Q(to_acu1
		[155]));
	notech_mux2 i_43302(.S(n_58292), .A(to_acu1[155]), .B(n_39671), .Z(n_35918
		));
	notech_reg to_acu1_reg_156(.CP(n_62195), .D(n_35924), .CD(n_61647), .Q(to_acu1
		[156]));
	notech_mux2 i_43310(.S(n_58292), .A(to_acu1[156]), .B(n_40409), .Z(n_35924
		));
	notech_reg to_acu1_reg_157(.CP(n_62192), .D(n_35930), .CD(n_61647), .Q(to_acu1
		[157]));
	notech_mux2 i_43318(.S(n_58292), .A(to_acu1[157]), .B(n_39673), .Z(n_35930
		));
	notech_reg to_acu1_reg_158(.CP(n_62192), .D(n_35936), .CD(n_61647), .Q(to_acu1
		[158]));
	notech_mux2 i_43326(.S(n_58292), .A(to_acu1[158]), .B(n_39675), .Z(n_35936
		));
	notech_reg to_acu1_reg_159(.CP(n_62192), .D(n_35942), .CD(n_61647), .Q(to_acu1
		[159]));
	notech_mux2 i_43334(.S(n_58292), .A(to_acu1[159]), .B(n_39677), .Z(n_35942
		));
	notech_reg to_acu1_reg_160(.CP(n_62192), .D(n_35948), .CD(n_61644), .Q(to_acu1
		[160]));
	notech_mux2 i_43342(.S(n_58292), .A(to_acu1[160]), .B(n_39679), .Z(n_35948
		));
	notech_reg to_acu1_reg_161(.CP(n_62192), .D(n_35954), .CD(n_61644), .Q(to_acu1
		[161]));
	notech_mux2 i_43350(.S(n_58293), .A(to_acu1[161]), .B(n_39683), .Z(n_35954
		));
	notech_reg to_acu1_reg_162(.CP(n_62192), .D(n_35960), .CD(n_61644), .Q(to_acu1
		[162]));
	notech_mux2 i_43358(.S(n_58293), .A(to_acu1[162]), .B(n_39685), .Z(n_35960
		));
	notech_reg to_acu1_reg_163(.CP(n_62192), .D(n_35966), .CD(n_61644), .Q(to_acu1
		[163]));
	notech_mux2 i_43366(.S(n_58293), .A(to_acu1[163]), .B(n_40417), .Z(n_35966
		));
	notech_reg to_acu1_reg_164(.CP(n_62192), .D(n_35972), .CD(n_61644), .Q(to_acu1
		[164]));
	notech_mux2 i_43374(.S(n_58292), .A(to_acu1[164]), .B(n_40419), .Z(n_35972
		));
	notech_reg to_acu1_reg_165(.CP(n_62192), .D(n_35978), .CD(n_61644), .Q(to_acu1
		[165]));
	notech_mux2 i_43382(.S(n_58293), .A(to_acu1[165]), .B(n_39687), .Z(n_35978
		));
	notech_reg to_acu1_reg_166(.CP(n_62192), .D(n_35984), .CD(n_61644), .Q(to_acu1
		[166]));
	notech_mux2 i_43390(.S(n_58293), .A(to_acu1[166]), .B(n_39689), .Z(n_35984
		));
	notech_reg to_acu1_reg_167(.CP(n_62192), .D(n_35990), .CD(n_61644), .Q(to_acu1
		[167]));
	notech_mux2 i_43398(.S(n_58298), .A(to_acu1[167]), .B(n_39691), .Z(n_35990
		));
	notech_reg to_acu1_reg_168(.CP(n_62160), .D(n_35996), .CD(n_61644), .Q(to_acu1
		[168]));
	notech_mux2 i_43406(.S(n_58303), .A(to_acu1[168]), .B(n_39694), .Z(n_35996
		));
	notech_reg to_acu1_reg_169(.CP(n_62160), .D(n_36002), .CD(n_61644), .Q(to_acu1
		[169]));
	notech_mux2 i_43414(.S(n_58303), .A(to_acu1[169]), .B(n_39696), .Z(n_36002
		));
	notech_reg to_acu1_reg_170(.CP(n_62160), .D(n_36008), .CD(n_61644), .Q(to_acu1
		[170]));
	notech_mux2 i_43422(.S(n_58303), .A(to_acu1[170]), .B(n_39698), .Z(n_36008
		));
	notech_reg to_acu1_reg_171(.CP(n_62160), .D(n_36014), .CD(n_61628), .Q(to_acu1
		[171]));
	notech_mux2 i_43430(.S(n_58303), .A(to_acu1[171]), .B(n_39700), .Z(n_36014
		));
	notech_reg to_acu1_reg_172(.CP(n_62160), .D(n_36020), .CD(n_61612), .Q(to_acu1
		[172]));
	notech_mux2 i_43438(.S(n_58303), .A(to_acu1[172]), .B(n_39702), .Z(n_36020
		));
	notech_reg to_acu1_reg_173(.CP(n_62160), .D(n_36026), .CD(n_61612), .Q(to_acu1
		[173]));
	notech_mux2 i_43446(.S(n_58303), .A(to_acu1[173]), .B(n_39704), .Z(n_36026
		));
	notech_reg to_acu1_reg_174(.CP(n_62160), .D(n_36032), .CD(n_61612), .Q(to_acu1
		[174]));
	notech_mux2 i_43454(.S(n_58303), .A(to_acu1[174]), .B(n_39706), .Z(n_36032
		));
	notech_reg to_acu1_reg_175(.CP(n_62160), .D(n_36038), .CD(n_61610), .Q(to_acu1
		[175]));
	notech_mux2 i_43462(.S(n_58303), .A(to_acu1[175]), .B(n_39708), .Z(n_36038
		));
	notech_reg to_acu1_reg_176(.CP(n_62160), .D(n_36044), .CD(n_61612), .Q(to_acu1
		[176]));
	notech_mux2 i_43470(.S(n_58303), .A(to_acu1[176]), .B(n_39710), .Z(n_36044
		));
	notech_reg to_acu1_reg_177(.CP(n_62160), .D(n_36050), .CD(n_61612), .Q(to_acu1
		[177]));
	notech_mux2 i_43478(.S(n_58303), .A(to_acu1[177]), .B(n_39712), .Z(n_36050
		));
	notech_reg to_acu1_reg_178(.CP(n_62158), .D(n_36056), .CD(n_61612), .Q(to_acu1
		[178]));
	notech_mux2 i_43486(.S(n_58303), .A(to_acu1[178]), .B(n_39714), .Z(n_36056
		));
	notech_reg to_acu1_reg_179(.CP(n_62158), .D(n_36062), .CD(n_61612), .Q(to_acu1
		[179]));
	notech_mux2 i_43494(.S(n_58303), .A(to_acu1[179]), .B(n_39716), .Z(n_36062
		));
	notech_reg to_acu1_reg_180(.CP(n_62158), .D(n_36068), .CD(n_61612), .Q(to_acu1
		[180]));
	notech_mux2 i_43502(.S(n_58303), .A(to_acu1[180]), .B(n_39115), .Z(n_36068
		));
	notech_reg to_acu1_reg_181(.CP(n_62158), .D(n_36074), .CD(n_61612), .Q(to_acu1
		[181]));
	notech_mux2 i_43510(.S(n_58298), .A(to_acu1[181]), .B(n_39718), .Z(n_36074
		));
	notech_reg to_acu1_reg_182(.CP(n_62158), .D(n_36080), .CD(n_61610), .Q(to_acu1
		[182]));
	notech_mux2 i_43518(.S(n_58298), .A(to_acu1[182]), .B(n_39720), .Z(n_36080
		));
	notech_reg to_acu1_reg_183(.CP(n_62158), .D(n_36086), .CD(n_61610), .Q(to_acu1
		[183]));
	notech_mux2 i_43526(.S(n_58298), .A(to_acu1[183]), .B(n_39722), .Z(n_36086
		));
	notech_reg to_acu1_reg_184(.CP(n_62158), .D(n_36092), .CD(n_61610), .Q(to_acu1
		[184]));
	notech_mux2 i_43534(.S(n_58298), .A(to_acu1[184]), .B(n_39724), .Z(n_36092
		));
	notech_reg to_acu1_reg_185(.CP(n_62158), .D(n_36098), .CD(n_61610), .Q(to_acu1
		[185]));
	notech_mux2 i_43542(.S(n_58298), .A(to_acu1[185]), .B(n_39726), .Z(n_36098
		));
	notech_reg to_acu1_reg_186(.CP(n_62158), .D(n_36104), .CD(n_61610), .Q(to_acu1
		[186]));
	notech_mux2 i_43550(.S(n_58298), .A(to_acu1[186]), .B(n_39728), .Z(n_36104
		));
	notech_reg to_acu1_reg_187(.CP(n_62158), .D(n_36110), .CD(n_61610), .Q(to_acu1
		[187]));
	notech_mux2 i_43558(.S(n_58298), .A(to_acu1[187]), .B(n_39730), .Z(n_36110
		));
	notech_reg to_acu1_reg_188(.CP(n_62158), .D(n_36116), .CD(n_61610), .Q(to_acu1
		[188]));
	notech_mux2 i_43566(.S(n_58298), .A(to_acu1[188]), .B(n_39732), .Z(n_36116
		));
	notech_reg to_acu1_reg_189(.CP(n_62163), .D(n_36122), .CD(n_61610), .Q(to_acu1
		[189]));
	notech_mux2 i_43574(.S(n_58303), .A(to_acu1[189]), .B(n_39734), .Z(n_36122
		));
	notech_reg to_acu1_reg_190(.CP(n_62163), .D(n_36128), .CD(n_61610), .Q(to_acu1
		[190]));
	notech_mux2 i_43582(.S(n_58303), .A(to_acu1[190]), .B(n_39736), .Z(n_36128
		));
	notech_reg to_acu1_reg_191(.CP(n_62163), .D(n_36134), .CD(n_61610), .Q(to_acu1
		[191]));
	notech_mux2 i_43590(.S(n_58298), .A(to_acu1[191]), .B(n_39738), .Z(n_36134
		));
	notech_reg to_acu1_reg_192(.CP(n_62163), .D(n_36140), .CD(n_61610), .Q(to_acu1
		[192]));
	notech_mux2 i_43598(.S(n_58298), .A(to_acu1[192]), .B(n_39740), .Z(n_36140
		));
	notech_reg to_acu1_reg_193(.CP(n_62163), .D(n_36146), .CD(n_61615), .Q(to_acu1
		[193]));
	notech_mux2 i_43606(.S(n_58298), .A(to_acu1[193]), .B(n_39742), .Z(n_36146
		));
	notech_reg to_acu1_reg_194(.CP(n_62163), .D(n_36152), .CD(n_61615), .Q(to_acu1
		[194]));
	notech_mux2 i_43614(.S(n_58281), .A(to_acu1[194]), .B(n_39744), .Z(n_36152
		));
	notech_reg to_acu1_reg_195(.CP(n_62163), .D(n_36158), .CD(n_61615), .Q(to_acu1
		[195]));
	notech_mux2 i_43622(.S(n_58281), .A(to_acu1[195]), .B(n_40451), .Z(n_36158
		));
	notech_reg to_acu1_reg_196(.CP(n_62163), .D(n_36164), .CD(n_61615), .Q(to_acu1
		[196]));
	notech_mux2 i_43630(.S(n_58281), .A(to_acu1[196]), .B(n_39746), .Z(n_36164
		));
	notech_reg to_acu1_reg_197(.CP(n_62163), .D(n_36170), .CD(n_61615), .Q(to_acu1
		[197]));
	notech_mux2 i_43638(.S(n_58281), .A(to_acu1[197]), .B(n_39748), .Z(n_36170
		));
	notech_reg to_acu1_reg_198(.CP(n_62163), .D(n_36176), .CD(n_61615), .Q(to_acu1
		[198]));
	notech_mux2 i_43646(.S(n_58281), .A(to_acu1[198]), .B(n_39750), .Z(n_36176
		));
	notech_reg to_acu1_reg_199(.CP(n_62163), .D(n_36182), .CD(n_61615), .Q(to_acu1
		[199]));
	notech_mux2 i_43654(.S(n_58281), .A(to_acu1[199]), .B(n_39752), .Z(n_36182
		));
	notech_reg to_acu1_reg_200(.CP(n_62160), .D(n_36188), .CD(n_61615), .Q(to_acu1
		[200]));
	notech_mux2 i_43662(.S(n_58281), .A(to_acu1[200]), .B(n_39754), .Z(n_36188
		));
	notech_reg to_acu1_reg_201(.CP(n_62160), .D(n_36194), .CD(n_61615), .Q(to_acu1
		[201]));
	notech_mux2 i_43670(.S(n_58281), .A(to_acu1[201]), .B(n_39756), .Z(n_36194
		));
	notech_reg to_acu1_reg_202(.CP(n_62160), .D(n_36200), .CD(n_61615), .Q(to_acu1
		[202]));
	notech_mux2 i_43678(.S(n_58281), .A(to_acu1[202]), .B(n_39758), .Z(n_36200
		));
	notech_reg to_acu1_reg_203(.CP(n_62160), .D(n_36206), .CD(n_61615), .Q(to_acu1
		[203]));
	notech_mux2 i_43686(.S(n_58281), .A(to_acu1[203]), .B(n_39760), .Z(n_36206
		));
	notech_reg to_acu1_reg_204(.CP(n_62160), .D(n_36212), .CD(n_61612), .Q(to_acu1
		[204]));
	notech_mux2 i_43694(.S(n_58281), .A(to_acu1[204]), .B(n_39762), .Z(n_36212
		));
	notech_reg to_acu1_reg_205(.CP(n_62163), .D(n_36218), .CD(n_61612), .Q(to_acu1
		[205]));
	notech_mux2 i_43702(.S(n_58281), .A(to_acu1[205]), .B(n_39763), .Z(n_36218
		));
	notech_reg to_acu1_reg_206(.CP(n_62163), .D(n_36224), .CD(n_61612), .Q(to_acu1
		[206]));
	notech_mux2 i_43710(.S(n_58281), .A(to_acu1[206]), .B(n_39765), .Z(n_36224
		));
	notech_reg to_acu1_reg_207(.CP(n_62160), .D(n_36230), .CD(n_61612), .Q(to_acu1
		[207]));
	notech_mux2 i_43718(.S(n_58280), .A(to_acu1[207]), .B(n_39767), .Z(n_36230
		));
	notech_reg to_acu1_reg_208(.CP(n_62160), .D(n_36236), .CD(n_61612), .Q(to_acu1
		[208]));
	notech_mux2 i_43726(.S(n_58280), .A(to_acu1[208]), .B(n_39769), .Z(n_36236
		));
	notech_reg to_acu1_reg_209(.CP(n_62160), .D(n_36242), .CD(n_61612), .Q(to_acu1
		[209]));
	notech_mux2 i_43734(.S(n_58280), .A(to_acu1[209]), .B(n_39771), .Z(n_36242
		));
	notech_reg to_acu1_reg_210(.CP(n_62158), .D(n_36248), .CD(n_61615), .Q(to_acu1
		[210]));
	notech_mux2 i_43742(.S(n_58280), .A(to_acu1[210]), .B(n_39773), .Z(n_36248
		));
	notech_reg overgs_reg(.CP(n_62153), .D(n_36254), .CD(n_61612), .Q(overgs
		));
	notech_mux2 i_43750(.S(n_3183), .A(n_41563), .B(overgs), .Z(n_36254));
	notech_reg iack_reg(.CP(n_62153), .D(n_39128), .CD(n_61612), .Q(iack));
	notech_reg over_seg2_reg_5(.CP(n_62153), .D(n_36262), .CD(n_61612), .Q(\over_seg2[5] 
		));
	notech_mux2 i_43762(.S(n_55061), .A(\over_seg2[5] ), .B(n_45938), .Z(n_36262
		));
	notech_reg over_seg1_reg_5(.CP(n_62153), .D(n_36268), .CD(n_61605), .Q(\over_seg1[5] 
		));
	notech_mux2 i_43770(.S(n_58280), .A(\over_seg1[5] ), .B(n_40471), .Z(n_36268
		));
	notech_reg over_seg0_reg_5(.CP(n_62153), .D(n_36274), .CD(n_61605), .Q(\over_seg0[5] 
		));
	notech_mux2 i_43778(.S(n_55699), .A(\over_seg0[5] ), .B(n_39114), .Z(n_36274
		));
	notech_reg imm0_reg_0(.CP(n_62155), .D(n_36280), .CD(n_61605), .Q(\imm0[0] 
		));
	notech_mux2 i_43786(.S(n_55699), .A(\imm0[0] ), .B(n_40142), .Z(n_36280)
		);
	notech_reg imm0_reg_1(.CP(n_62155), .D(n_36286), .CD(n_61605), .Q(\imm0[1] 
		));
	notech_mux2 i_43794(.S(n_55669), .A(\imm0[1] ), .B(n_40145), .Z(n_36286)
		);
	notech_reg imm0_reg_2(.CP(n_62155), .D(n_36292), .CD(n_61605), .Q(\imm0[2] 
		));
	notech_mux2 i_43802(.S(n_55669), .A(\imm0[2] ), .B(n_40148), .Z(n_36292)
		);
	notech_reg imm0_reg_3(.CP(n_62153), .D(n_36298), .CD(n_61607), .Q(\imm0[3] 
		));
	notech_mux2 i_43810(.S(n_55699), .A(\imm0[3] ), .B(n_40151), .Z(n_36298)
		);
	notech_reg imm0_reg_4(.CP(n_62153), .D(n_36304), .CD(n_61607), .Q(\imm0[4] 
		));
	notech_mux2 i_43818(.S(n_55699), .A(\imm0[4] ), .B(n_40154), .Z(n_36304)
		);
	notech_reg imm0_reg_5(.CP(n_62153), .D(n_36310), .CD(n_61607), .Q(\imm0[5] 
		));
	notech_mux2 i_43826(.S(n_55699), .A(\imm0[5] ), .B(n_40157), .Z(n_36310)
		);
	notech_reg imm0_reg_6(.CP(n_62153), .D(n_36316), .CD(n_61605), .Q(\imm0[6] 
		));
	notech_mux2 i_43834(.S(n_55699), .A(\imm0[6] ), .B(n_40160), .Z(n_36316)
		);
	notech_reg imm0_reg_7(.CP(n_62153), .D(n_36322), .CD(n_61605), .Q(\imm0[7] 
		));
	notech_mux2 i_43842(.S(n_55669), .A(\imm0[7] ), .B(n_40163), .Z(n_36322)
		);
	notech_reg imm0_reg_8(.CP(n_62153), .D(n_36328), .CD(n_61605), .Q(\imm0[8] 
		));
	notech_mux2 i_43850(.S(n_55669), .A(\imm0[8] ), .B(n_40166), .Z(n_36328)
		);
	notech_reg imm0_reg_9(.CP(n_62153), .D(n_36334), .CD(n_61605), .Q(\imm0[9] 
		));
	notech_mux2 i_43858(.S(n_55669), .A(\imm0[9] ), .B(n_40169), .Z(n_36334)
		);
	notech_reg imm0_reg_10(.CP(n_62153), .D(n_36340), .CD(n_61605), .Q(\imm0[10] 
		));
	notech_mux2 i_43866(.S(n_55669), .A(\imm0[10] ), .B(n_40172), .Z(n_36340
		));
	notech_reg imm0_reg_11(.CP(n_62153), .D(n_36346), .CD(n_61605), .Q(\imm0[11] 
		));
	notech_mux2 i_43874(.S(n_55669), .A(\imm0[11] ), .B(n_40174), .Z(n_36346
		));
	notech_reg imm0_reg_12(.CP(n_62153), .D(n_36352), .CD(n_61605), .Q(\imm0[12] 
		));
	notech_mux2 i_43882(.S(n_55669), .A(\imm0[12] ), .B(n_40176), .Z(n_36352
		));
	notech_reg imm0_reg_13(.CP(n_62153), .D(n_36358), .CD(n_61605), .Q(\imm0[13] 
		));
	notech_mux2 i_43890(.S(n_55669), .A(\imm0[13] ), .B(n_40181), .Z(n_36358
		));
	notech_reg imm0_reg_14(.CP(n_62153), .D(n_36364), .CD(n_61605), .Q(\imm0[14] 
		));
	notech_mux2 i_43898(.S(n_55669), .A(\imm0[14] ), .B(n_39367), .Z(n_36364
		));
	notech_reg imm0_reg_15(.CP(n_62153), .D(n_36370), .CD(n_61605), .Q(\imm0[15] 
		));
	notech_mux2 i_43906(.S(n_55699), .A(\imm0[15] ), .B(n_40184), .Z(n_36370
		));
	notech_reg imm0_reg_16(.CP(n_62155), .D(n_36376), .CD(n_61605), .Q(\imm0[16] 
		));
	notech_mux2 i_43914(.S(n_55703), .A(\imm0[16] ), .B(n_39369), .Z(n_36376
		));
	notech_reg imm0_reg_17(.CP(n_62158), .D(n_36382), .CD(n_61605), .Q(\imm0[17] 
		));
	notech_mux2 i_43922(.S(n_55703), .A(\imm0[17] ), .B(n_40186), .Z(n_36382
		));
	notech_reg imm0_reg_18(.CP(n_62155), .D(n_36388), .CD(n_61605), .Q(\imm0[18] 
		));
	notech_mux2 i_43930(.S(n_55703), .A(\imm0[18] ), .B(n_40190), .Z(n_36388
		));
	notech_reg imm0_reg_19(.CP(n_62155), .D(n_36394), .CD(n_61607), .Q(\imm0[19] 
		));
	notech_mux2 i_43938(.S(n_55703), .A(\imm0[19] ), .B(n_39371), .Z(n_36394
		));
	notech_reg imm0_reg_20(.CP(n_62155), .D(n_36400), .CD(n_61610), .Q(\imm0[20] 
		));
	notech_mux2 i_43946(.S(n_55703), .A(\imm0[20] ), .B(n_40192), .Z(n_36400
		));
	notech_reg imm0_reg_21(.CP(n_62158), .D(n_36406), .CD(n_61607), .Q(\imm0[21] 
		));
	notech_mux2 i_43954(.S(n_55703), .A(\imm0[21] ), .B(n_40194), .Z(n_36406
		));
	notech_reg imm0_reg_22(.CP(n_62158), .D(n_36412), .CD(n_61607), .Q(\imm0[22] 
		));
	notech_mux2 i_43962(.S(n_55703), .A(\imm0[22] ), .B(n_40196), .Z(n_36412
		));
	notech_reg imm0_reg_23(.CP(n_62158), .D(n_36418), .CD(n_61607), .Q(\imm0[23] 
		));
	notech_mux2 i_43970(.S(n_55703), .A(\imm0[23] ), .B(n_40198), .Z(n_36418
		));
	notech_reg imm0_reg_24(.CP(n_62158), .D(n_36424), .CD(n_61610), .Q(\imm0[24] 
		));
	notech_mux2 i_43978(.S(n_55699), .A(\imm0[24] ), .B(n_40200), .Z(n_36424
		));
	notech_reg imm0_reg_25(.CP(n_62158), .D(n_36430), .CD(n_61610), .Q(\imm0[25] 
		));
	notech_mux2 i_43986(.S(n_55699), .A(\imm0[25] ), .B(n_39372), .Z(n_36430
		));
	notech_reg imm0_reg_26(.CP(n_62155), .D(n_36436), .CD(n_61610), .Q(\imm0[26] 
		));
	notech_mux2 i_43994(.S(n_55699), .A(\imm0[26] ), .B(n_40202), .Z(n_36436
		));
	notech_reg imm0_reg_27(.CP(n_62155), .D(n_36442), .CD(n_61610), .Q(\imm0[27] 
		));
	notech_mux2 i_44002(.S(n_55699), .A(\imm0[27] ), .B(n_40204), .Z(n_36442
		));
	notech_reg imm0_reg_28(.CP(n_62155), .D(n_36448), .CD(n_61610), .Q(\imm0[28] 
		));
	notech_mux2 i_44010(.S(n_55699), .A(\imm0[28] ), .B(n_40206), .Z(n_36448
		));
	notech_reg imm0_reg_29(.CP(n_62155), .D(n_36454), .CD(n_61607), .Q(\imm0[29] 
		));
	notech_mux2 i_44018(.S(n_55699), .A(\imm0[29] ), .B(n_40208), .Z(n_36454
		));
	notech_reg imm0_reg_30(.CP(n_62155), .D(n_36460), .CD(n_61607), .Q(\imm0[30] 
		));
	notech_mux2 i_44026(.S(n_55699), .A(\imm0[30] ), .B(n_40210), .Z(n_36460
		));
	notech_reg imm0_reg_31(.CP(n_62155), .D(n_36466), .CD(n_61607), .Q(\imm0[31] 
		));
	notech_mux2 i_44034(.S(n_55699), .A(\imm0[31] ), .B(n_40212), .Z(n_36466
		));
	notech_reg imm0_reg_32(.CP(n_62155), .D(n_36472), .CD(n_61607), .Q(\imm0[32] 
		));
	notech_mux2 i_44042(.S(n_55684), .A(\imm0[32] ), .B(n_40214), .Z(n_36472
		));
	notech_reg imm0_reg_33(.CP(n_62155), .D(n_36478), .CD(n_61607), .Q(\imm0[33] 
		));
	notech_mux2 i_44050(.S(n_55684), .A(\imm0[33] ), .B(n_40216), .Z(n_36478
		));
	notech_reg imm0_reg_34(.CP(n_62155), .D(n_36484), .CD(n_61607), .Q(\imm0[34] 
		));
	notech_mux2 i_44058(.S(n_55684), .A(\imm0[34] ), .B(n_39112), .Z(n_36484
		));
	notech_reg imm0_reg_35(.CP(n_62155), .D(n_36490), .CD(n_61607), .Q(\imm0[35] 
		));
	notech_mux2 i_44066(.S(n_55684), .A(\imm0[35] ), .B(n_40218), .Z(n_36490
		));
	notech_reg imm0_reg_36(.CP(n_62155), .D(n_36496), .CD(n_61607), .Q(\imm0[36] 
		));
	notech_mux2 i_44074(.S(n_55689), .A(\imm0[36] ), .B(n_40220), .Z(n_36496
		));
	notech_reg imm0_reg_37(.CP(n_62171), .D(n_36502), .CD(n_61607), .Q(\imm0[37] 
		));
	notech_mux2 i_44082(.S(n_55689), .A(\imm0[37] ), .B(n_40222), .Z(n_36502
		));
	notech_reg imm0_reg_38(.CP(n_62171), .D(n_36508), .CD(n_61607), .Q(\imm0[38] 
		));
	notech_mux2 i_44090(.S(n_55684), .A(\imm0[38] ), .B(n_40224), .Z(n_36508
		));
	notech_reg imm0_reg_39(.CP(n_62171), .D(n_36514), .CD(n_61607), .Q(\imm0[39] 
		));
	notech_mux2 i_44098(.S(n_55689), .A(\imm0[39] ), .B(n_40226), .Z(n_36514
		));
	notech_reg imm0_reg_40(.CP(n_62171), .D(n_36520), .CD(n_61615), .Q(\imm0[40] 
		));
	notech_mux2 i_44106(.S(n_55684), .A(\imm0[40] ), .B(n_40228), .Z(n_36520
		));
	notech_reg imm0_reg_41(.CP(n_62171), .D(n_36526), .CD(n_61623), .Q(\imm0[41] 
		));
	notech_mux2 i_44114(.S(n_55684), .A(\imm0[41] ), .B(n_39373), .Z(n_36526
		));
	notech_reg imm0_reg_42(.CP(n_62174), .D(n_36532), .CD(n_61623), .Q(\imm0[42] 
		));
	notech_mux2 i_44122(.S(n_55684), .A(\imm0[42] ), .B(n_40230), .Z(n_36532
		));
	notech_reg imm0_reg_43(.CP(n_62174), .D(n_36538), .CD(n_61623), .Q(\imm0[43] 
		));
	notech_mux2 i_44130(.S(n_55684), .A(\imm0[43] ), .B(n_40232), .Z(n_36538
		));
	notech_reg imm0_reg_44(.CP(n_62174), .D(n_36544), .CD(n_61623), .Q(\imm0[44] 
		));
	notech_mux2 i_44138(.S(n_55684), .A(\imm0[44] ), .B(n_39113), .Z(n_36544
		));
	notech_reg imm0_reg_45(.CP(n_62174), .D(n_36550), .CD(n_61623), .Q(\imm0[45] 
		));
	notech_mux2 i_44146(.S(n_55684), .A(\imm0[45] ), .B(n_39375), .Z(n_36550
		));
	notech_reg imm0_reg_46(.CP(n_62174), .D(n_36556), .CD(n_61626), .Q(\imm0[46] 
		));
	notech_mux2 i_44154(.S(n_55684), .A(\imm0[46] ), .B(n_40234), .Z(n_36556
		));
	notech_reg imm0_reg_47(.CP(n_62171), .D(n_36562), .CD(n_61626), .Q(\imm0[47] 
		));
	notech_mux2 i_44162(.S(n_55684), .A(\imm0[47] ), .B(n_40236), .Z(n_36562
		));
	notech_reg lenpc1_reg_0(.CP(n_62171), .D(n_36568), .CD(n_61626), .Q(lenpc1
		[0]));
	notech_mux2 i_44170(.S(n_58280), .A(lenpc1[0]), .B(n_40124), .Z(n_36568)
		);
	notech_reg lenpc1_reg_1(.CP(n_62171), .D(n_36574), .CD(n_61623), .Q(lenpc1
		[1]));
	notech_mux2 i_44178(.S(n_58280), .A(lenpc1[1]), .B(n_40127), .Z(n_36574)
		);
	notech_reg lenpc1_reg_2(.CP(n_62171), .D(n_36580), .CD(n_61626), .Q(lenpc1
		[2]));
	notech_mux2 i_44186(.S(n_58280), .A(lenpc1[2]), .B(n_40130), .Z(n_36580)
		);
	notech_reg lenpc1_reg_3(.CP(n_62171), .D(n_36586), .CD(n_61623), .Q(lenpc1
		[3]));
	notech_mux2 i_44194(.S(n_58280), .A(lenpc1[3]), .B(n_40133), .Z(n_36586)
		);
	notech_reg lenpc1_reg_4(.CP(n_62171), .D(n_36592), .CD(n_61623), .Q(lenpc1
		[4]));
	notech_mux2 i_44202(.S(n_58280), .A(lenpc1[4]), .B(n_40136), .Z(n_36592)
		);
	notech_reg lenpc1_reg_5(.CP(n_62171), .D(n_36598), .CD(n_61623), .Q(lenpc1
		[5]));
	notech_mux2 i_44210(.S(n_58280), .A(lenpc1[5]), .B(n_40139), .Z(n_36598)
		);
	notech_reg lenpc1_reg_6(.CP(n_62171), .D(n_36604), .CD(n_61623), .Q(lenpc1
		[6]));
	notech_mux2 i_44218(.S(n_58280), .A(lenpc1[6]), .B(n_133896033), .Z(n_36604
		));
	notech_reg lenpc1_reg_7(.CP(n_62171), .D(n_36610), .CD(n_61623), .Q(lenpc1
		[7]));
	notech_mux2 i_44226(.S(n_58280), .A(lenpc1[7]), .B(n_44145), .Z(n_36610)
		);
	notech_reg lenpc1_reg_8(.CP(n_62171), .D(n_36616), .CD(n_61623), .Q(lenpc1
		[8]));
	notech_mux2 i_44234(.S(n_58281), .A(lenpc1[8]), .B(n_133996034), .Z(n_36616
		));
	notech_reg lenpc1_reg_9(.CP(n_62171), .D(n_36622), .CD(n_61623), .Q(lenpc1
		[9]));
	notech_mux2 i_44242(.S(n_58292), .A(lenpc1[9]), .B(n_44157), .Z(n_36622)
		);
	notech_reg lenpc1_reg_10(.CP(n_62176), .D(n_36628), .CD(n_61623), .Q(lenpc1
		[10]));
	notech_mux2 i_44250(.S(n_58292), .A(lenpc1[10]), .B(n_44163), .Z(n_36628
		));
	notech_reg lenpc1_reg_11(.CP(n_62176), .D(n_36634), .CD(n_61623), .Q(lenpc1
		[11]));
	notech_mux2 i_44258(.S(n_58292), .A(lenpc1[11]), .B(n_44169), .Z(n_36634
		));
	notech_reg lenpc1_reg_12(.CP(n_62176), .D(n_36640), .CD(n_61623), .Q(lenpc1
		[12]));
	notech_mux2 i_44266(.S(n_58287), .A(lenpc1[12]), .B(n_44175), .Z(n_36640
		));
	notech_reg lenpc1_reg_13(.CP(n_62174), .D(n_36646), .CD(n_61623), .Q(lenpc1
		[13]));
	notech_mux2 i_44274(.S(n_58287), .A(lenpc1[13]), .B(n_134096035), .Z(n_36646
		));
	notech_reg lenpc1_reg_14(.CP(n_62174), .D(n_36652), .CD(n_61628), .Q(lenpc1
		[14]));
	notech_mux2 i_44282(.S(n_58287), .A(lenpc1[14]), .B(n_134196036), .Z(n_36652
		));
	notech_reg lenpc1_reg_15(.CP(n_62176), .D(n_36658), .CD(n_61628), .Q(lenpc1
		[15]));
	notech_mux2 i_44290(.S(n_58292), .A(lenpc1[15]), .B(n_134296037), .Z(n_36658
		));
	notech_reg lenpc1_reg_16(.CP(n_62176), .D(n_36664), .CD(n_61626), .Q(lenpc1
		[16]));
	notech_mux2 i_44298(.S(n_58292), .A(lenpc1[16]), .B(n_134396038), .Z(n_36664
		));
	notech_reg lenpc1_reg_17(.CP(n_62176), .D(n_36670), .CD(n_61626), .Q(lenpc1
		[17]));
	notech_mux2 i_44306(.S(n_58292), .A(lenpc1[17]), .B(n_134496039), .Z(n_36670
		));
	notech_reg lenpc1_reg_18(.CP(n_62176), .D(n_36676), .CD(n_61626), .Q(lenpc1
		[18]));
	notech_mux2 i_44314(.S(n_58292), .A(lenpc1[18]), .B(n_134596040), .Z(n_36676
		));
	notech_reg lenpc1_reg_19(.CP(n_62176), .D(n_36682), .CD(n_61628), .Q(lenpc1
		[19]));
	notech_mux2 i_44322(.S(n_58292), .A(lenpc1[19]), .B(n_44217), .Z(n_36682
		));
	notech_reg lenpc1_reg_20(.CP(n_62174), .D(n_36688), .CD(n_61628), .Q(lenpc1
		[20]));
	notech_mux2 i_44330(.S(n_58292), .A(lenpc1[20]), .B(n_134696041), .Z(n_36688
		));
	notech_reg lenpc1_reg_21(.CP(n_62174), .D(n_36694), .CD(n_61628), .Q(lenpc1
		[21]));
	notech_mux2 i_44338(.S(n_58292), .A(lenpc1[21]), .B(n_134796042), .Z(n_36694
		));
	notech_reg lenpc1_reg_22(.CP(n_62174), .D(n_36700), .CD(n_61628), .Q(lenpc1
		[22]));
	notech_mux2 i_44346(.S(n_58281), .A(lenpc1[22]), .B(n_134896043), .Z(n_36700
		));
	notech_reg lenpc1_reg_23(.CP(n_62174), .D(n_36706), .CD(n_61628), .Q(lenpc1
		[23]));
	notech_mux2 i_44354(.S(n_58287), .A(lenpc1[23]), .B(n_134996044), .Z(n_36706
		));
	notech_reg lenpc1_reg_24(.CP(n_62174), .D(n_36712), .CD(n_61626), .Q(lenpc1
		[24]));
	notech_mux2 i_44362(.S(n_58287), .A(lenpc1[24]), .B(n_44247), .Z(n_36712
		));
	notech_reg lenpc1_reg_25(.CP(n_62174), .D(n_36718), .CD(n_61626), .Q(lenpc1
		[25]));
	notech_mux2 i_44370(.S(n_58281), .A(lenpc1[25]), .B(n_135096045), .Z(n_36718
		));
	notech_reg lenpc1_reg_26(.CP(n_62174), .D(n_36724), .CD(n_61626), .Q(lenpc1
		[26]));
	notech_mux2 i_44378(.S(n_58281), .A(lenpc1[26]), .B(n_44259), .Z(n_36724
		));
	notech_reg lenpc1_reg_27(.CP(n_62174), .D(n_36730), .CD(n_61626), .Q(lenpc1
		[27]));
	notech_mux2 i_44386(.S(n_58281), .A(lenpc1[27]), .B(n_135196046), .Z(n_36730
		));
	notech_reg lenpc1_reg_28(.CP(n_62174), .D(n_36736), .CD(n_61626), .Q(lenpc1
		[28]));
	notech_mux2 i_44394(.S(n_58287), .A(lenpc1[28]), .B(n_135296047), .Z(n_36736
		));
	notech_reg lenpc1_reg_29(.CP(n_62174), .D(n_36742), .CD(n_61626), .Q(lenpc1
		[29]));
	notech_mux2 i_44402(.S(n_58287), .A(lenpc1[29]), .B(n_135396048), .Z(n_36742
		));
	notech_reg lenpc1_reg_30(.CP(n_62174), .D(n_36748), .CD(n_61626), .Q(lenpc1
		[30]));
	notech_mux2 i_44410(.S(n_58287), .A(lenpc1[30]), .B(n_135496049), .Z(n_36748
		));
	notech_reg lenpc1_reg_31(.CP(n_62171), .D(n_36754), .CD(n_61626), .Q(lenpc1
		[31]));
	notech_mux2 i_44418(.S(n_58287), .A(lenpc1[31]), .B(n_44289), .Z(n_36754
		));
	notech_reg lenpc_reg_0(.CP(n_62165), .D(n_36760), .CD(n_61626), .Q(lenpc
		[0]));
	notech_mux2 i_44426(.S(n_3185), .A(n_40480), .B(lenpc[0]), .Z(n_36760)
		);
	notech_reg lenpc_reg_1(.CP(n_62165), .D(n_36766), .CD(n_61626), .Q(lenpc
		[1]));
	notech_mux2 i_44434(.S(n_3185), .A(n_40481), .B(lenpc[1]), .Z(n_36766)
		);
	notech_reg lenpc_reg_2(.CP(n_62165), .D(n_36772), .CD(n_61626), .Q(lenpc
		[2]));
	notech_mux2 i_44442(.S(n_3185), .A(n_40482), .B(lenpc[2]), .Z(n_36772)
		);
	notech_reg lenpc_reg_3(.CP(n_62165), .D(n_36778), .CD(n_61617), .Q(lenpc
		[3]));
	notech_mux2 i_44450(.S(n_3185), .A(n_40483), .B(lenpc[3]), .Z(n_36778)
		);
	notech_reg lenpc_reg_4(.CP(n_62165), .D(n_36784), .CD(n_61617), .Q(lenpc
		[4]));
	notech_mux2 i_44458(.S(n_3185), .A(n_40484), .B(lenpc[4]), .Z(n_36784)
		);
	notech_reg lenpc_reg_5(.CP(n_62165), .D(n_36790), .CD(n_61617), .Q(lenpc
		[5]));
	notech_mux2 i_44466(.S(n_3185), .A(n_40485), .B(lenpc[5]), .Z(n_36790)
		);
	notech_reg lenpc_reg_6(.CP(n_62165), .D(n_36796), .CD(n_61617), .Q(lenpc
		[6]));
	notech_mux2 i_44474(.S(n_3185), .A(n_131296007), .B(lenpc[6]), .Z(n_36796
		));
	notech_reg lenpc_reg_7(.CP(n_62165), .D(n_36802), .CD(n_61617), .Q(lenpc
		[7]));
	notech_mux2 i_44482(.S(n_3185), .A(n_131396008), .B(lenpc[7]), .Z(n_36802
		));
	notech_reg lenpc_reg_8(.CP(n_62165), .D(n_36808), .CD(n_61617), .Q(lenpc
		[8]));
	notech_mux2 i_44490(.S(n_3185), .A(n_131496009), .B(lenpc[8]), .Z(n_36808
		));
	notech_reg lenpc_reg_9(.CP(n_62165), .D(n_36814), .CD(n_61617), .Q(lenpc
		[9]));
	notech_mux2 i_44498(.S(n_3185), .A(n_131596010), .B(lenpc[9]), .Z(n_36814
		));
	notech_reg lenpc_reg_10(.CP(n_62165), .D(n_36820), .CD(n_61617), .Q(lenpc
		[10]));
	notech_mux2 i_44506(.S(n_3185), .A(n_131696011), .B(lenpc[10]), .Z(n_36820
		));
	notech_reg lenpc_reg_11(.CP(n_62163), .D(n_36826), .CD(n_61617), .Q(lenpc
		[11]));
	notech_mux2 i_44514(.S(n_3185), .A(n_131796012), .B(lenpc[11]), .Z(n_36826
		));
	notech_reg lenpc_reg_12(.CP(n_62163), .D(n_36832), .CD(n_61617), .Q(lenpc
		[12]));
	notech_mux2 i_44522(.S(n_3185), .A(n_131896013), .B(lenpc[12]), .Z(n_36832
		));
	notech_reg lenpc_reg_13(.CP(n_62163), .D(n_36838), .CD(n_61617), .Q(lenpc
		[13]));
	notech_mux2 i_44530(.S(n_3185), .A(n_131996014), .B(lenpc[13]), .Z(n_36838
		));
	notech_reg lenpc_reg_14(.CP(n_62163), .D(n_36844), .CD(n_61615), .Q(lenpc
		[14]));
	notech_mux2 i_44538(.S(n_3185), .A(n_132096015), .B(lenpc[14]), .Z(n_36844
		));
	notech_reg lenpc_reg_15(.CP(n_62163), .D(n_36850), .CD(n_61615), .Q(lenpc
		[15]));
	notech_mux2 i_44546(.S(n_3185), .A(n_132196016), .B(lenpc[15]), .Z(n_36850
		));
	notech_reg lenpc_reg_16(.CP(n_62165), .D(n_36856), .CD(n_61615), .Q(lenpc
		[16]));
	notech_mux2 i_44554(.S(n_59067), .A(n_132296017), .B(lenpc[16]), .Z(n_36856
		));
	notech_reg lenpc_reg_17(.CP(n_62165), .D(n_36862), .CD(n_61615), .Q(lenpc
		[17]));
	notech_mux2 i_44562(.S(n_59067), .A(n_132396018), .B(lenpc[17]), .Z(n_36862
		));
	notech_reg lenpc_reg_18(.CP(n_62165), .D(n_36868), .CD(n_61615), .Q(lenpc
		[18]));
	notech_mux2 i_44570(.S(n_59067), .A(n_132496019), .B(lenpc[18]), .Z(n_36868
		));
	notech_reg lenpc_reg_19(.CP(n_62165), .D(n_36874), .CD(n_61617), .Q(lenpc
		[19]));
	notech_mux2 i_44578(.S(n_59067), .A(n_132596020), .B(lenpc[19]), .Z(n_36874
		));
	notech_reg lenpc_reg_20(.CP(n_62165), .D(n_36880), .CD(n_61617), .Q(lenpc
		[20]));
	notech_mux2 i_44586(.S(n_59067), .A(n_132696021), .B(lenpc[20]), .Z(n_36880
		));
	notech_reg lenpc_reg_21(.CP(n_62169), .D(n_36886), .CD(n_61617), .Q(lenpc
		[21]));
	notech_mux2 i_44594(.S(n_59067), .A(n_132796022), .B(lenpc[21]), .Z(n_36886
		));
	notech_reg lenpc_reg_22(.CP(n_62169), .D(n_36892), .CD(n_61617), .Q(lenpc
		[22]));
	notech_mux2 i_44602(.S(n_59067), .A(n_132896023), .B(lenpc[22]), .Z(n_36892
		));
	notech_reg lenpc_reg_23(.CP(n_62169), .D(n_36898), .CD(n_61617), .Q(lenpc
		[23]));
	notech_mux2 i_44610(.S(n_59067), .A(n_132996024), .B(lenpc[23]), .Z(n_36898
		));
	notech_reg lenpc_reg_24(.CP(n_62169), .D(n_36904), .CD(n_61621), .Q(lenpc
		[24]));
	notech_mux2 i_44618(.S(n_59067), .A(n_133096025), .B(lenpc[24]), .Z(n_36904
		));
	notech_reg lenpc_reg_25(.CP(n_62169), .D(n_36910), .CD(n_61621), .Q(lenpc
		[25]));
	notech_mux2 i_44626(.S(n_59067), .A(n_133196026), .B(lenpc[25]), .Z(n_36910
		));
	notech_reg lenpc_reg_26(.CP(n_62169), .D(n_36916), .CD(n_61621), .Q(lenpc
		[26]));
	notech_mux2 i_44634(.S(n_3185), .A(n_133296027), .B(lenpc[26]), .Z(n_36916
		));
	notech_reg lenpc_reg_27(.CP(n_62171), .D(n_36922), .CD(n_61621), .Q(lenpc
		[27]));
	notech_mux2 i_44642(.S(n_59067), .A(n_133396028), .B(lenpc[27]), .Z(n_36922
		));
	notech_reg lenpc_reg_28(.CP(n_62169), .D(n_36928), .CD(n_61621), .Q(lenpc
		[28]));
	notech_mux2 i_44650(.S(n_59067), .A(n_133496029), .B(lenpc[28]), .Z(n_36928
		));
	notech_reg lenpc_reg_29(.CP(n_62169), .D(n_36934), .CD(n_61621), .Q(lenpc
		[29]));
	notech_mux2 i_44658(.S(n_59067), .A(n_133596030), .B(lenpc[29]), .Z(n_36934
		));
	notech_reg lenpc_reg_30(.CP(n_62169), .D(n_36940), .CD(n_61623), .Q(lenpc
		[30]));
	notech_mux2 i_44666(.S(n_59067), .A(n_133696031), .B(lenpc[30]), .Z(n_36940
		));
	notech_reg lenpc_reg_31(.CP(n_62169), .D(n_36946), .CD(n_61621), .Q(lenpc
		[31]));
	notech_mux2 i_44674(.S(n_59067), .A(n_133796032), .B(lenpc[31]), .Z(n_36946
		));
	notech_reg opz2_reg_0(.CP(n_62169), .D(n_36952), .CD(n_61621), .Q(opz2[0
		]));
	notech_mux2 i_44682(.S(n_55061), .A(opz2[0]), .B(n_3239), .Z(n_36952));
	notech_reg opz2_reg_1(.CP(n_62169), .D(n_36958), .CD(n_61621), .Q(opz2[1
		]));
	notech_mux2 i_44690(.S(n_55061), .A(opz2[1]), .B(n_3237), .Z(n_36958));
	notech_reg_set opz2_reg_2(.CP(n_62169), .D(n_36964), .SD(n_61621), .Q(opz2
		[2]));
	notech_mux2 i_44698(.S(n_55061), .A(opz2[2]), .B(n_273394690), .Z(n_36964
		));
	notech_reg opz1_reg_0(.CP(n_62165), .D(n_36970), .CD(n_61621), .Q(opz1[0
		]));
	notech_mux2 i_44706(.S(n_58287), .A(opz1[0]), .B(n_40118), .Z(n_36970)
		);
	notech_reg opz1_reg_1(.CP(n_62165), .D(n_36976), .CD(n_61621), .Q(opz1[1
		]));
	notech_mux2 i_44714(.S(n_58287), .A(opz1[1]), .B(n_40121), .Z(n_36976)
		);
	notech_reg_set opz1_reg_2(.CP(n_62169), .D(n_36982), .SD(n_61621), .Q(opz1
		[2]));
	notech_mux2 i_44722(.S(n_58287), .A(opz1[2]), .B(n_273594692), .Z(n_36982
		));
	notech_reg opz0_reg_0(.CP(n_62169), .D(n_36988), .CD(n_61617), .Q(opz0[0
		]));
	notech_mux2 i_44730(.S(n_55689), .A(opz0[0]), .B(n_40112), .Z(n_36988)
		);
	notech_reg opz0_reg_1(.CP(n_62169), .D(n_36994), .CD(n_61617), .Q(opz0[1
		]));
	notech_mux2 i_44738(.S(n_55689), .A(opz0[1]), .B(n_40115), .Z(n_36994)
		);
	notech_reg_set opz0_reg_2(.CP(n_62169), .D(n_37000), .SD(n_61621), .Q(opz0
		[2]));
	notech_mux2 i_44746(.S(n_55669), .A(opz0[2]), .B(n_273794694), .Z(n_37000
		));
	notech_reg_set inst_deco_reg_0(.CP(n_62169), .D(n_37006), .SD(n_61621), 
		.Q(inst_deco[0]));
	notech_mux2 i_44754(.S(n_59058), .A(n_45072), .B(inst_deco[0]), .Z(n_37006
		));
	notech_reg_set inst_deco_reg_1(.CP(n_62201), .D(n_37012), .SD(n_61621), 
		.Q(inst_deco[1]));
	notech_mux2 i_44762(.S(n_59058), .A(n_45078), .B(inst_deco[1]), .Z(n_37012
		));
	notech_reg_set inst_deco_reg_2(.CP(n_62236), .D(n_37018), .SD(n_61621), 
		.Q(inst_deco[2]));
	notech_mux2 i_44770(.S(n_59058), .A(n_45084), .B(inst_deco[2]), .Z(n_37018
		));
	notech_reg_set inst_deco_reg_3(.CP(n_62236), .D(n_37024), .SD(n_61621), 
		.Q(inst_deco[3]));
	notech_mux2 i_44778(.S(n_59058), .A(n_45090), .B(inst_deco[3]), .Z(n_37024
		));
	notech_reg_set inst_deco_reg_4(.CP(n_62236), .D(n_37030), .SD(n_61688), 
		.Q(inst_deco[4]));
	notech_mux2 i_44786(.S(n_59058), .A(n_45096), .B(inst_deco[4]), .Z(n_37030
		));
	notech_reg_set inst_deco_reg_5(.CP(n_62236), .D(n_37036), .SD(n_61688), 
		.Q(inst_deco[5]));
	notech_mux2 i_44794(.S(n_59058), .A(n_45102), .B(inst_deco[5]), .Z(n_37036
		));
	notech_reg_set inst_deco_reg_6(.CP(n_62236), .D(n_37042), .SD(n_61688), 
		.Q(inst_deco[6]));
	notech_mux2 i_44802(.S(n_59058), .A(n_45108), .B(inst_deco[6]), .Z(n_37042
		));
	notech_reg_set inst_deco_reg_7(.CP(n_62236), .D(n_37048), .SD(n_61688), 
		.Q(inst_deco[7]));
	notech_mux2 i_44810(.S(n_59058), .A(n_45114), .B(inst_deco[7]), .Z(n_37048
		));
	notech_reg_set inst_deco_reg_8(.CP(n_62236), .D(n_37054), .SD(n_61688), 
		.Q(inst_deco[8]));
	notech_mux2 i_44818(.S(n_59058), .A(n_45120), .B(inst_deco[8]), .Z(n_37054
		));
	notech_reg_set inst_deco_reg_9(.CP(n_62236), .D(n_37060), .SD(n_61688), 
		.Q(inst_deco[9]));
	notech_mux2 i_44826(.S(n_59058), .A(n_45126), .B(inst_deco[9]), .Z(n_37060
		));
	notech_reg_set inst_deco_reg_10(.CP(n_62236), .D(n_37066), .SD(n_61688),
		 .Q(inst_deco[10]));
	notech_mux2 i_44834(.S(n_59058), .A(n_3270), .B(inst_deco[10]), .Z(n_37066
		));
	notech_reg_set inst_deco_reg_11(.CP(n_62236), .D(n_37072), .SD(n_61688),
		 .Q(inst_deco[11]));
	notech_mux2 i_44842(.S(n_59058), .A(n_45138), .B(inst_deco[11]), .Z(n_37072
		));
	notech_reg_set inst_deco_reg_12(.CP(n_62236), .D(n_37078), .SD(n_61688),
		 .Q(inst_deco[12]));
	notech_mux2 i_44850(.S(n_59058), .A(n_45144), .B(inst_deco[12]), .Z(n_37078
		));
	notech_reg_set inst_deco_reg_13(.CP(n_62234), .D(n_37084), .SD(n_61688),
		 .Q(inst_deco[13]));
	notech_mux2 i_44858(.S(n_59058), .A(n_3269), .B(inst_deco[13]), .Z(n_37084
		));
	notech_reg_set inst_deco_reg_14(.CP(n_62236), .D(n_37090), .SD(n_61688),
		 .Q(inst_deco[14]));
	notech_mux2 i_44866(.S(n_59058), .A(n_45156), .B(inst_deco[14]), .Z(n_37090
		));
	notech_reg_set inst_deco_reg_15(.CP(n_62234), .D(n_37096), .SD(n_61686),
		 .Q(inst_deco[15]));
	notech_mux2 i_44874(.S(n_59058), .A(n_45162), .B(inst_deco[15]), .Z(n_37096
		));
	notech_reg_set inst_deco_reg_16(.CP(n_62234), .D(n_37102), .SD(n_61686),
		 .Q(inst_deco[16]));
	notech_mux2 i_44882(.S(n_59056), .A(n_45168), .B(inst_deco[16]), .Z(n_37102
		));
	notech_reg_set inst_deco_reg_17(.CP(n_62234), .D(n_37108), .SD(n_61686),
		 .Q(inst_deco[17]));
	notech_mux2 i_44890(.S(n_59056), .A(n_45174), .B(inst_deco[17]), .Z(n_37108
		));
	notech_reg_set inst_deco_reg_18(.CP(n_62236), .D(n_37114), .SD(n_61686),
		 .Q(inst_deco[18]));
	notech_mux2 i_44898(.S(n_59056), .A(n_45180), .B(inst_deco[18]), .Z(n_37114
		));
	notech_reg_set inst_deco_reg_19(.CP(n_62236), .D(n_37120), .SD(n_61686),
		 .Q(inst_deco[19]));
	notech_mux2 i_44906(.S(n_59056), .A(n_45186), .B(inst_deco[19]), .Z(n_37120
		));
	notech_reg_set inst_deco_reg_20(.CP(n_62236), .D(n_37126), .SD(n_61688),
		 .Q(inst_deco[20]));
	notech_mux2 i_44914(.S(n_59056), .A(n_45192), .B(inst_deco[20]), .Z(n_37126
		));
	notech_reg_set inst_deco_reg_21(.CP(n_62236), .D(n_37132), .SD(n_61688),
		 .Q(inst_deco[21]));
	notech_mux2 i_44922(.S(n_59056), .A(n_45198), .B(inst_deco[21]), .Z(n_37132
		));
	notech_reg_set inst_deco_reg_22(.CP(n_62236), .D(n_37138), .SD(n_61688),
		 .Q(inst_deco[22]));
	notech_mux2 i_44930(.S(n_59056), .A(n_45204), .B(inst_deco[22]), .Z(n_37138
		));
	notech_reg_set inst_deco_reg_23(.CP(n_62239), .D(n_37144), .SD(n_61686),
		 .Q(inst_deco[23]));
	notech_mux2 i_44938(.S(n_59056), .A(n_45210), .B(inst_deco[23]), .Z(n_37144
		));
	notech_reg_set inst_deco_reg_24(.CP(n_62239), .D(n_37150), .SD(n_61688),
		 .Q(inst_deco[24]));
	notech_mux2 i_44946(.S(n_59056), .A(n_45216), .B(inst_deco[24]), .Z(n_37150
		));
	notech_reg_set inst_deco_reg_25(.CP(n_62239), .D(n_37156), .SD(n_61691),
		 .Q(inst_deco[25]));
	notech_mux2 i_44954(.S(n_59056), .A(n_45222), .B(inst_deco[25]), .Z(n_37156
		));
	notech_reg_set inst_deco_reg_26(.CP(n_62239), .D(n_37162), .SD(n_61691),
		 .Q(inst_deco[26]));
	notech_mux2 i_44962(.S(n_59056), .A(n_45228), .B(inst_deco[26]), .Z(n_37162
		));
	notech_reg_set inst_deco_reg_27(.CP(n_62239), .D(n_37168), .SD(n_61691),
		 .Q(inst_deco[27]));
	notech_mux2 i_44970(.S(n_59056), .A(n_45234), .B(inst_deco[27]), .Z(n_37168
		));
	notech_reg_set inst_deco_reg_28(.CP(n_62241), .D(n_37174), .SD(n_61691),
		 .Q(inst_deco[28]));
	notech_mux2 i_44978(.S(n_59056), .A(n_45240), .B(inst_deco[28]), .Z(n_37174
		));
	notech_reg_set inst_deco_reg_29(.CP(n_62241), .D(n_37181), .SD(n_61691),
		 .Q(inst_deco[29]));
	notech_mux2 i_44986(.S(n_59056), .A(n_45246), .B(inst_deco[29]), .Z(n_37181
		));
	notech_reg_set inst_deco_reg_30(.CP(n_62239), .D(n_37187), .SD(n_61691),
		 .Q(inst_deco[30]));
	notech_mux2 i_44994(.S(n_59056), .A(n_3268), .B(inst_deco[30]), .Z(n_37187
		));
	notech_reg_set inst_deco_reg_31(.CP(n_62239), .D(n_37193), .SD(n_61691),
		 .Q(inst_deco[31]));
	notech_mux2 i_45002(.S(n_59056), .A(n_45258), .B(inst_deco[31]), .Z(n_37193
		));
	notech_reg_set inst_deco_reg_32(.CP(n_62239), .D(n_37199), .SD(n_61691),
		 .Q(inst_deco[32]));
	notech_mux2 i_45010(.S(n_59063), .A(n_45264), .B(inst_deco[32]), .Z(n_37199
		));
	notech_reg_set inst_deco_reg_33(.CP(n_62239), .D(n_37205), .SD(n_61691),
		 .Q(inst_deco[33]));
	notech_mux2 i_45018(.S(n_59063), .A(n_45270), .B(inst_deco[33]), .Z(n_37205
		));
	notech_reg_set inst_deco_reg_34(.CP(n_62239), .D(n_37211), .SD(n_61691),
		 .Q(inst_deco[34]));
	notech_mux2 i_45026(.S(n_59063), .A(n_45276), .B(inst_deco[34]), .Z(n_37211
		));
	notech_reg_set inst_deco_reg_35(.CP(n_62239), .D(n_37217), .SD(n_61691),
		 .Q(inst_deco[35]));
	notech_mux2 i_45034(.S(n_59063), .A(n_45282), .B(inst_deco[35]), .Z(n_37217
		));
	notech_reg_set inst_deco_reg_36(.CP(n_62239), .D(n_37223), .SD(n_61691),
		 .Q(inst_deco[36]));
	notech_mux2 i_45042(.S(n_59063), .A(n_45288), .B(inst_deco[36]), .Z(n_37223
		));
	notech_reg_set inst_deco_reg_37(.CP(n_62236), .D(n_37229), .SD(n_61691),
		 .Q(inst_deco[37]));
	notech_mux2 i_45050(.S(n_59063), .A(n_45294), .B(inst_deco[37]), .Z(n_37229
		));
	notech_reg_set inst_deco_reg_38(.CP(n_62239), .D(n_37235), .SD(n_61688),
		 .Q(inst_deco[38]));
	notech_mux2 i_45058(.S(n_59063), .A(n_45300), .B(inst_deco[38]), .Z(n_37235
		));
	notech_reg_set inst_deco_reg_39(.CP(n_62239), .D(n_37241), .SD(n_61688),
		 .Q(inst_deco[39]));
	notech_mux2 i_45066(.S(n_59063), .A(n_45306), .B(inst_deco[39]), .Z(n_37241
		));
	notech_reg_set inst_deco_reg_40(.CP(n_62239), .D(n_37247), .SD(n_61688),
		 .Q(inst_deco[40]));
	notech_mux2 i_45074(.S(n_59063), .A(n_45312), .B(inst_deco[40]), .Z(n_37247
		));
	notech_reg_set inst_deco_reg_41(.CP(n_62239), .D(n_37253), .SD(n_61691),
		 .Q(inst_deco[41]));
	notech_mux2 i_45082(.S(n_59063), .A(n_45318), .B(inst_deco[41]), .Z(n_37253
		));
	notech_reg_set inst_deco_reg_42(.CP(n_62239), .D(n_37259), .SD(n_61691),
		 .Q(inst_deco[42]));
	notech_mux2 i_45090(.S(n_59063), .A(n_45324), .B(inst_deco[42]), .Z(n_37259
		));
	notech_reg_set inst_deco_reg_43(.CP(n_62239), .D(n_37265), .SD(n_61691),
		 .Q(inst_deco[43]));
	notech_mux2 i_45098(.S(n_59063), .A(n_45330), .B(inst_deco[43]), .Z(n_37265
		));
	notech_reg_set inst_deco_reg_44(.CP(n_62234), .D(n_37271), .SD(n_61691),
		 .Q(inst_deco[44]));
	notech_mux2 i_45106(.S(n_59063), .A(n_45336), .B(inst_deco[44]), .Z(n_37271
		));
	notech_reg_set inst_deco_reg_45(.CP(n_62230), .D(n_37277), .SD(n_61691),
		 .Q(inst_deco[45]));
	notech_mux2 i_45114(.S(n_59063), .A(n_45342), .B(inst_deco[45]), .Z(n_37277
		));
	notech_reg_set inst_deco_reg_46(.CP(n_62230), .D(n_37283), .SD(n_61682),
		 .Q(inst_deco[46]));
	notech_mux2 i_45122(.S(n_59063), .A(n_45348), .B(inst_deco[46]), .Z(n_37283
		));
	notech_reg_set inst_deco_reg_47(.CP(n_62230), .D(n_37289), .SD(n_61682),
		 .Q(inst_deco[47]));
	notech_mux2 i_45130(.S(n_59063), .A(n_45354), .B(inst_deco[47]), .Z(n_37289
		));
	notech_reg_set inst_deco_reg_48(.CP(n_62230), .D(n_37295), .SD(n_61682),
		 .Q(inst_deco[48]));
	notech_mux2 i_45138(.S(n_59061), .A(n_45360), .B(inst_deco[48]), .Z(n_37295
		));
	notech_reg_set inst_deco_reg_49(.CP(n_62230), .D(n_37301), .SD(n_61680),
		 .Q(inst_deco[49]));
	notech_mux2 i_45146(.S(n_59061), .A(n_45366), .B(inst_deco[49]), .Z(n_37301
		));
	notech_reg_set inst_deco_reg_50(.CP(n_62230), .D(n_37307), .SD(n_61682),
		 .Q(inst_deco[50]));
	notech_mux2 i_45154(.S(n_59061), .A(n_45372), .B(inst_deco[50]), .Z(n_37307
		));
	notech_reg_set inst_deco_reg_51(.CP(n_62230), .D(n_37313), .SD(n_61682),
		 .Q(inst_deco[51]));
	notech_mux2 i_45162(.S(n_59061), .A(n_3267), .B(inst_deco[51]), .Z(n_37313
		));
	notech_reg_set inst_deco_reg_52(.CP(n_62230), .D(n_37319), .SD(n_61682),
		 .Q(inst_deco[52]));
	notech_mux2 i_45170(.S(n_59061), .A(n_45384), .B(inst_deco[52]), .Z(n_37319
		));
	notech_reg_set inst_deco_reg_53(.CP(n_62230), .D(n_37325), .SD(n_61682),
		 .Q(inst_deco[53]));
	notech_mux2 i_45178(.S(n_59061), .A(n_45390), .B(inst_deco[53]), .Z(n_37325
		));
	notech_reg_set inst_deco_reg_54(.CP(n_62230), .D(n_37331), .SD(n_61682),
		 .Q(inst_deco[54]));
	notech_mux2 i_45186(.S(n_59061), .A(n_45396), .B(inst_deco[54]), .Z(n_37331
		));
	notech_reg_set inst_deco_reg_55(.CP(n_62228), .D(n_37337), .SD(n_61682),
		 .Q(inst_deco[55]));
	notech_mux2 i_45194(.S(n_59061), .A(n_45402), .B(inst_deco[55]), .Z(n_37337
		));
	notech_reg_set inst_deco_reg_56(.CP(n_62228), .D(n_37343), .SD(n_61680),
		 .Q(inst_deco[56]));
	notech_mux2 i_45202(.S(n_59061), .A(n_45408), .B(inst_deco[56]), .Z(n_37343
		));
	notech_reg_set inst_deco_reg_57(.CP(n_62228), .D(n_37349), .SD(n_61680),
		 .Q(inst_deco[57]));
	notech_mux2 i_45210(.S(n_59061), .A(n_45414), .B(inst_deco[57]), .Z(n_37349
		));
	notech_reg_set inst_deco_reg_58(.CP(n_62228), .D(n_37355), .SD(n_61680),
		 .Q(inst_deco[58]));
	notech_mux2 i_45218(.S(n_59061), .A(n_3266), .B(inst_deco[58]), .Z(n_37355
		));
	notech_reg_set inst_deco_reg_59(.CP(n_62228), .D(n_37361), .SD(n_61680),
		 .Q(inst_deco[59]));
	notech_mux2 i_45226(.S(n_59061), .A(n_3265), .B(inst_deco[59]), .Z(n_37361
		));
	notech_reg_set inst_deco_reg_60(.CP(n_62228), .D(n_37367), .SD(n_61680),
		 .Q(inst_deco[60]));
	notech_mux2 i_45234(.S(n_59061), .A(n_3264), .B(inst_deco[60]), .Z(n_37367
		));
	notech_reg_set inst_deco_reg_61(.CP(n_62228), .D(n_37373), .SD(n_61680),
		 .Q(inst_deco[61]));
	notech_mux2 i_45242(.S(n_59061), .A(n_45438), .B(inst_deco[61]), .Z(n_37373
		));
	notech_reg_set inst_deco_reg_62(.CP(n_62228), .D(n_37379), .SD(n_61680),
		 .Q(inst_deco[62]));
	notech_mux2 i_45250(.S(n_59061), .A(n_45444), .B(inst_deco[62]), .Z(n_37379
		));
	notech_reg_set inst_deco_reg_63(.CP(n_62228), .D(n_37385), .SD(n_61680),
		 .Q(inst_deco[63]));
	notech_mux2 i_45258(.S(n_59061), .A(n_45450), .B(inst_deco[63]), .Z(n_37385
		));
	notech_reg_set inst_deco_reg_64(.CP(n_62228), .D(n_37391), .SD(n_61680),
		 .Q(inst_deco[64]));
	notech_mux2 i_45266(.S(n_59048), .A(n_45456), .B(inst_deco[64]), .Z(n_37391
		));
	notech_reg_set inst_deco_reg_65(.CP(n_62228), .D(n_37397), .SD(n_61680),
		 .Q(inst_deco[65]));
	notech_mux2 i_45274(.S(n_59048), .A(n_3263), .B(inst_deco[65]), .Z(n_37397
		));
	notech_reg_set inst_deco_reg_66(.CP(n_62234), .D(n_37403), .SD(n_61680),
		 .Q(inst_deco[66]));
	notech_mux2 i_45282(.S(n_59048), .A(n_45468), .B(inst_deco[66]), .Z(n_37403
		));
	notech_reg_set inst_deco_reg_67(.CP(n_62234), .D(n_37409), .SD(n_61686),
		 .Q(inst_deco[67]));
	notech_mux2 i_45290(.S(n_59048), .A(n_45474), .B(inst_deco[67]), .Z(n_37409
		));
	notech_reg_set inst_deco_reg_68(.CP(n_62234), .D(n_37415), .SD(n_61686),
		 .Q(inst_deco[68]));
	notech_mux2 i_45298(.S(n_59048), .A(n_45480), .B(inst_deco[68]), .Z(n_37415
		));
	notech_reg_set inst_deco_reg_69(.CP(n_62234), .D(n_37421), .SD(n_61686),
		 .Q(inst_deco[69]));
	notech_mux2 i_45306(.S(n_59048), .A(n_45486), .B(inst_deco[69]), .Z(n_37421
		));
	notech_reg_set inst_deco_reg_70(.CP(n_62234), .D(n_37427), .SD(n_61686),
		 .Q(inst_deco[70]));
	notech_mux2 i_45314(.S(n_59048), .A(n_45492), .B(inst_deco[70]), .Z(n_37427
		));
	notech_reg_set inst_deco_reg_71(.CP(n_62234), .D(n_37433), .SD(n_61686),
		 .Q(inst_deco[71]));
	notech_mux2 i_45322(.S(n_59048), .A(n_45498), .B(inst_deco[71]), .Z(n_37433
		));
	notech_reg_set inst_deco_reg_72(.CP(n_62234), .D(n_37439), .SD(n_61686),
		 .Q(inst_deco[72]));
	notech_mux2 i_45330(.S(n_59048), .A(n_274494701), .B(inst_deco[72]), .Z(n_37439
		));
	notech_reg_set inst_deco_reg_73(.CP(n_62234), .D(n_37445), .SD(n_61686),
		 .Q(inst_deco[73]));
	notech_mux2 i_45338(.S(n_59048), .A(n_3262), .B(inst_deco[73]), .Z(n_37445
		));
	notech_reg_set inst_deco_reg_74(.CP(n_62234), .D(n_37451), .SD(n_61686),
		 .Q(inst_deco[74]));
	notech_mux2 i_45346(.S(n_59048), .A(n_45516), .B(inst_deco[74]), .Z(n_37451
		));
	notech_reg_set inst_deco_reg_75(.CP(n_62234), .D(n_37457), .SD(n_61686),
		 .Q(inst_deco[75]));
	notech_mux2 i_45354(.S(n_59048), .A(n_45522), .B(inst_deco[75]), .Z(n_37457
		));
	notech_reg_set inst_deco_reg_76(.CP(n_62234), .D(n_37463), .SD(n_61686),
		 .Q(inst_deco[76]));
	notech_mux2 i_45362(.S(n_59048), .A(n_45528), .B(inst_deco[76]), .Z(n_37463
		));
	notech_reg_set inst_deco_reg_77(.CP(n_62230), .D(n_37469), .SD(n_61686),
		 .Q(inst_deco[77]));
	notech_mux2 i_45370(.S(n_59048), .A(n_45534), .B(inst_deco[77]), .Z(n_37469
		));
	notech_reg_set inst_deco_reg_78(.CP(n_62230), .D(n_37475), .SD(n_61682),
		 .Q(inst_deco[78]));
	notech_mux2 i_45378(.S(n_59048), .A(n_45540), .B(inst_deco[78]), .Z(n_37475
		));
	notech_reg_set inst_deco_reg_79(.CP(n_62230), .D(n_37481), .SD(n_61682),
		 .Q(inst_deco[79]));
	notech_mux2 i_45386(.S(n_59048), .A(n_45546), .B(inst_deco[79]), .Z(n_37481
		));
	notech_reg_set inst_deco_reg_80(.CP(n_62230), .D(n_37487), .SD(n_61682),
		 .Q(inst_deco[80]));
	notech_mux2 i_45394(.S(n_59046), .A(n_3261), .B(inst_deco[80]), .Z(n_37487
		));
	notech_reg_set inst_deco_reg_81(.CP(n_62230), .D(n_37493), .SD(n_61682),
		 .Q(inst_deco[81]));
	notech_mux2 i_45402(.S(n_59046), .A(n_3260), .B(inst_deco[81]), .Z(n_37493
		));
	notech_reg_set inst_deco_reg_82(.CP(n_62234), .D(n_37499), .SD(n_61682),
		 .Q(inst_deco[82]));
	notech_mux2 i_45410(.S(n_59046), .A(n_3259), .B(inst_deco[82]), .Z(n_37499
		));
	notech_reg_set inst_deco_reg_83(.CP(n_62234), .D(n_37505), .SD(n_61682),
		 .Q(inst_deco[83]));
	notech_mux2 i_45418(.S(n_59046), .A(n_3258), .B(inst_deco[83]), .Z(n_37505
		));
	notech_reg_set inst_deco_reg_84(.CP(n_62230), .D(n_37511), .SD(n_61686),
		 .Q(inst_deco[84]));
	notech_mux2 i_45426(.S(n_59046), .A(n_3257), .B(inst_deco[84]), .Z(n_37511
		));
	notech_reg_set inst_deco_reg_85(.CP(n_62230), .D(n_37517), .SD(n_61682),
		 .Q(inst_deco[85]));
	notech_mux2 i_45434(.S(n_59046), .A(n_3256), .B(inst_deco[85]), .Z(n_37517
		));
	notech_reg_set inst_deco_reg_86(.CP(n_62230), .D(n_37523), .SD(n_61682),
		 .Q(inst_deco[86]));
	notech_mux2 i_45442(.S(n_59046), .A(n_3255), .B(inst_deco[86]), .Z(n_37523
		));
	notech_reg_set inst_deco_reg_87(.CP(n_62250), .D(n_37529), .SD(n_61682),
		 .Q(inst_deco[87]));
	notech_mux2 i_45450(.S(n_59046), .A(n_3254), .B(inst_deco[87]), .Z(n_37529
		));
	notech_reg_set inst_deco_reg_88(.CP(n_62250), .D(n_37535), .SD(n_61693),
		 .Q(inst_deco[88]));
	notech_mux2 i_45458(.S(n_59046), .A(n_3253), .B(inst_deco[88]), .Z(n_37535
		));
	notech_reg_set inst_deco_reg_89(.CP(n_62250), .D(n_37541), .SD(n_61702),
		 .Q(inst_deco[89]));
	notech_mux2 i_45466(.S(n_59046), .A(n_3252), .B(inst_deco[89]), .Z(n_37541
		));
	notech_reg_set inst_deco_reg_90(.CP(n_62250), .D(n_37547), .SD(n_61702),
		 .Q(inst_deco[90]));
	notech_mux2 i_45474(.S(n_59046), .A(n_3251), .B(inst_deco[90]), .Z(n_37547
		));
	notech_reg_set inst_deco_reg_91(.CP(n_62250), .D(n_37553), .SD(n_61702),
		 .Q(inst_deco[91]));
	notech_mux2 i_45482(.S(n_59046), .A(n_274094697), .B(inst_deco[91]), .Z(n_37553
		));
	notech_reg_set inst_deco_reg_92(.CP(n_62250), .D(n_37559), .SD(n_61702),
		 .Q(inst_deco[92]));
	notech_mux2 i_45490(.S(n_59046), .A(n_3250), .B(inst_deco[92]), .Z(n_37559
		));
	notech_reg_set inst_deco_reg_93(.CP(n_62250), .D(n_37565), .SD(n_61702),
		 .Q(inst_deco[93]));
	notech_mux2 i_45498(.S(n_59046), .A(n_3249), .B(inst_deco[93]), .Z(n_37565
		));
	notech_reg_set inst_deco_reg_94(.CP(n_62250), .D(n_37571), .SD(n_61702),
		 .Q(inst_deco[94]));
	notech_mux2 i_45506(.S(n_59046), .A(n_3248), .B(inst_deco[94]), .Z(n_37571
		));
	notech_reg_set inst_deco_reg_95(.CP(n_62250), .D(n_37577), .SD(n_61702),
		 .Q(inst_deco[95]));
	notech_mux2 i_45514(.S(n_59046), .A(n_3247), .B(inst_deco[95]), .Z(n_37577
		));
	notech_reg_set inst_deco_reg_96(.CP(n_62250), .D(n_37583), .SD(n_61702),
		 .Q(inst_deco[96]));
	notech_mux2 i_45522(.S(n_59053), .A(n_3246), .B(inst_deco[96]), .Z(n_37583
		));
	notech_reg_set inst_deco_reg_97(.CP(n_62250), .D(n_37589), .SD(n_61702),
		 .Q(inst_deco[97]));
	notech_mux2 i_45530(.S(n_59053), .A(n_3245), .B(inst_deco[97]), .Z(n_37589
		));
	notech_reg_set inst_deco_reg_98(.CP(n_62246), .D(n_37595), .SD(n_61702),
		 .Q(inst_deco[98]));
	notech_mux2 i_45538(.S(n_59053), .A(n_3244), .B(inst_deco[98]), .Z(n_37595
		));
	notech_reg_set inst_deco_reg_99(.CP(n_62246), .D(n_37601), .SD(n_61698),
		 .Q(inst_deco[99]));
	notech_mux2 i_45546(.S(n_59053), .A(n_3243), .B(inst_deco[99]), .Z(n_37601
		));
	notech_reg_set inst_deco_reg_100(.CP(n_62246), .D(n_37607), .SD(n_61698)
		, .Q(inst_deco[100]));
	notech_mux2 i_45554(.S(n_59053), .A(n_45672), .B(inst_deco[100]), .Z(n_37607
		));
	notech_reg_set inst_deco_reg_101(.CP(n_62246), .D(n_37613), .SD(n_61698)
		, .Q(inst_deco[101]));
	notech_mux2 i_45562(.S(n_59053), .A(n_45678), .B(inst_deco[101]), .Z(n_37613
		));
	notech_reg_set inst_deco_reg_102(.CP(n_62246), .D(n_37619), .SD(n_61698)
		, .Q(inst_deco[102]));
	notech_mux2 i_45570(.S(n_59053), .A(n_45684), .B(inst_deco[102]), .Z(n_37619
		));
	notech_reg_set inst_deco_reg_103(.CP(n_62246), .D(n_37625), .SD(n_61698)
		, .Q(inst_deco[103]));
	notech_mux2 i_45578(.S(n_59053), .A(n_45690), .B(inst_deco[103]), .Z(n_37625
		));
	notech_reg_set inst_deco_reg_104(.CP(n_62250), .D(n_37631), .SD(n_61698)
		, .Q(inst_deco[104]));
	notech_mux2 i_45586(.S(n_59053), .A(n_45696), .B(inst_deco[104]), .Z(n_37631
		));
	notech_reg_set inst_deco_reg_105(.CP(n_62246), .D(n_37637), .SD(n_61698)
		, .Q(inst_deco[105]));
	notech_mux2 i_45594(.S(n_59053), .A(n_45702), .B(inst_deco[105]), .Z(n_37637
		));
	notech_reg_set inst_deco_reg_106(.CP(n_62246), .D(n_37643), .SD(n_61698)
		, .Q(inst_deco[106]));
	notech_mux2 i_45602(.S(n_59053), .A(n_45708), .B(inst_deco[106]), .Z(n_37643
		));
	notech_reg_set inst_deco_reg_107(.CP(n_62246), .D(n_37649), .SD(n_61698)
		, .Q(inst_deco[107]));
	notech_mux2 i_45610(.S(n_59053), .A(n_45714), .B(inst_deco[107]), .Z(n_37649
		));
	notech_reg_set inst_deco_reg_108(.CP(n_62252), .D(n_37655), .SD(n_61698)
		, .Q(inst_deco[108]));
	notech_mux2 i_45618(.S(n_59053), .A(n_45720), .B(inst_deco[108]), .Z(n_37655
		));
	notech_reg_set inst_deco_reg_109(.CP(n_62252), .D(n_37661), .SD(n_61698)
		, .Q(inst_deco[109]));
	notech_mux2 i_45626(.S(n_59053), .A(n_45726), .B(inst_deco[109]), .Z(n_37661
		));
	notech_reg_set inst_deco_reg_110(.CP(n_62252), .D(n_37667), .SD(n_61704)
		, .Q(inst_deco[110]));
	notech_mux2 i_45634(.S(n_59053), .A(n_45732), .B(inst_deco[110]), .Z(n_37667
		));
	notech_reg_set inst_deco_reg_111(.CP(n_62252), .D(n_37673), .SD(n_61704)
		, .Q(inst_deco[111]));
	notech_mux2 i_45642(.S(n_59053), .A(n_45738), .B(inst_deco[111]), .Z(n_37673
		));
	notech_reg_set inst_deco_reg_112(.CP(n_62252), .D(n_37679), .SD(n_61704)
		, .Q(inst_deco[112]));
	notech_mux2 i_45650(.S(n_59051), .A(n_45744), .B(inst_deco[112]), .Z(n_37679
		));
	notech_reg_set inst_deco_reg_113(.CP(n_62252), .D(n_37685), .SD(n_61704)
		, .Q(inst_deco[113]));
	notech_mux2 i_45658(.S(n_59051), .A(n_45750), .B(inst_deco[113]), .Z(n_37685
		));
	notech_reg_set inst_deco_reg_114(.CP(n_62252), .D(n_37691), .SD(n_61704)
		, .Q(inst_deco[114]));
	notech_mux2 i_45666(.S(n_59051), .A(n_45756), .B(inst_deco[114]), .Z(n_37691
		));
	notech_reg_set inst_deco_reg_115(.CP(n_62252), .D(n_37697), .SD(n_61704)
		, .Q(inst_deco[115]));
	notech_mux2 i_45674(.S(n_59051), .A(n_45762), .B(inst_deco[115]), .Z(n_37697
		));
	notech_reg_set inst_deco_reg_116(.CP(n_62252), .D(n_37703), .SD(n_61704)
		, .Q(inst_deco[116]));
	notech_mux2 i_45682(.S(n_59051), .A(n_45768), .B(inst_deco[116]), .Z(n_37703
		));
	notech_reg_set inst_deco_reg_117(.CP(n_62252), .D(n_37709), .SD(n_61704)
		, .Q(inst_deco[117]));
	notech_mux2 i_45690(.S(n_59051), .A(n_45774), .B(inst_deco[117]), .Z(n_37709
		));
	notech_reg_set inst_deco_reg_118(.CP(n_62252), .D(n_37715), .SD(n_61704)
		, .Q(inst_deco[118]));
	notech_mux2 i_45698(.S(n_59051), .A(n_45780), .B(inst_deco[118]), .Z(n_37715
		));
	notech_reg_set inst_deco_reg_119(.CP(n_62250), .D(n_37721), .SD(n_61704)
		, .Q(inst_deco[119]));
	notech_mux2 i_45706(.S(n_59051), .A(n_45786), .B(inst_deco[119]), .Z(n_37721
		));
	notech_reg_set inst_deco_reg_120(.CP(n_62250), .D(n_37727), .SD(n_61704)
		, .Q(inst_deco[120]));
	notech_mux2 i_45714(.S(n_59051), .A(n_45792), .B(inst_deco[120]), .Z(n_37727
		));
	notech_reg_set inst_deco_reg_121(.CP(n_62250), .D(n_37733), .SD(n_61702)
		, .Q(inst_deco[121]));
	notech_mux2 i_45722(.S(n_59051), .A(n_45798), .B(inst_deco[121]), .Z(n_37733
		));
	notech_reg_set inst_deco_reg_122(.CP(n_62250), .D(n_37739), .SD(n_61702)
		, .Q(inst_deco[122]));
	notech_mux2 i_45730(.S(n_59051), .A(n_45804), .B(inst_deco[122]), .Z(n_37739
		));
	notech_reg_set inst_deco_reg_123(.CP(n_62250), .D(n_37745), .SD(n_61702)
		, .Q(inst_deco[123]));
	notech_mux2 i_45738(.S(n_59051), .A(n_45810), .B(inst_deco[123]), .Z(n_37745
		));
	notech_ao4 i_17473980(.A(n_40267), .B(n_3137), .C(n_40941), .D(n_3136), 
		.Z(n_1644));
	notech_reg_set inst_deco_reg_124(.CP(n_62252), .D(n_37751), .SD(n_61702)
		, .Q(inst_deco[124]));
	notech_mux2 i_45746(.S(n_59051), .A(n_45816), .B(inst_deco[124]), .Z(n_37751
		));
	notech_and2 i_2774127(.A(n_2149), .B(n_40534), .Z(n_1643));
	notech_reg_set inst_deco_reg_125(.CP(n_62252), .D(n_37757), .SD(n_61702)
		, .Q(inst_deco[125]));
	notech_mux2 i_45754(.S(n_59051), .A(n_45822), .B(inst_deco[125]), .Z(n_37757
		));
	notech_ao4 i_125474542(.A(n_59006), .B(n_39635), .C(n_59082), .D(n_40605
		), .Z(n_1642));
	notech_reg_set inst_deco_reg_126(.CP(n_62252), .D(n_37763), .SD(n_61704)
		, .Q(inst_deco[126]));
	notech_mux2 i_45762(.S(n_59051), .A(n_45828), .B(inst_deco[126]), .Z(n_37763
		));
	notech_ao4 i_125774539(.A(n_59006), .B(n_39641), .C(n_59082), .D(n_40608
		), .Z(n_1641));
	notech_reg_set inst_deco_reg_127(.CP(n_62250), .D(n_37769), .SD(n_61704)
		, .Q(inst_deco[127]));
	notech_mux2 i_45770(.S(n_59051), .A(n_45834), .B(inst_deco[127]), .Z(n_37769
		));
	notech_ao4 i_127474522(.A(n_59004), .B(n_39678), .C(n_59082), .D(n_40625
		), .Z(n_1640));
	notech_reg reps0_reg_0(.CP(n_62252), .D(n_37775), .CD(n_61702), .Q(reps0
		[0]));
	notech_mux2 i_45778(.S(n_55689), .A(reps0[0]), .B(n_40082), .Z(n_37775)
		);
	notech_ao4 i_129574501(.A(n_59004), .B(n_39721), .C(n_59082), .D(n_40646
		), .Z(n_1639));
	notech_reg reps0_reg_1(.CP(n_62246), .D(n_37781), .CD(n_61702), .Q(reps0
		[1]));
	notech_mux2 i_45786(.S(n_55689), .A(reps0[1]), .B(n_40085), .Z(n_37781)
		);
	notech_ao4 i_130274494(.A(n_59006), .B(n_39735), .C(n_59082), .D(n_40653
		), .Z(n_1638));
	notech_reg reps0_reg_2(.CP(n_62241), .D(n_37787), .CD(n_61702), .Q(reps0
		[2]));
	notech_mux2 i_45794(.S(n_55669), .A(reps0[2]), .B(n_39111), .Z(n_37787)
		);
	notech_ao4 i_130374493(.A(n_59004), .B(n_39737), .C(n_59084), .D(n_40654
		), .Z(n_1637));
	notech_reg to_acu0_reg_0(.CP(n_62241), .D(n_37793), .CD(n_61693), .Q(to_acu0
		[0]));
	notech_mux2 i_45802(.S(n_55669), .A(to_acu0[0]), .B(n_40507), .Z(n_37793
		));
	notech_ao4 i_130474492(.A(n_59001), .B(n_39739), .C(n_59084), .D(n_40655
		), .Z(n_1636));
	notech_reg to_acu0_reg_1(.CP(n_62241), .D(n_37799), .CD(n_61693), .Q(to_acu0
		[1]));
	notech_mux2 i_45810(.S(n_55669), .A(to_acu0[1]), .B(n_39066), .Z(n_37799
		));
	notech_ao4 i_130974487(.A(n_59001), .B(n_39749), .C(n_59084), .D(n_40660
		), .Z(n_1635));
	notech_reg to_acu0_reg_2(.CP(n_62241), .D(n_37805), .CD(n_61693), .Q(to_acu0
		[2]));
	notech_mux2 i_45818(.S(n_55669), .A(to_acu0[2]), .B(n_39067), .Z(n_37805
		));
	notech_ao4 i_131674480(.A(n_59001), .B(n_39764), .C(n_59084), .D(n_40668
		), .Z(n_1634));
	notech_reg to_acu0_reg_3(.CP(n_62241), .D(n_37811), .CD(n_61693), .Q(to_acu0
		[3]));
	notech_mux2 i_45826(.S(n_55689), .A(to_acu0[3]), .B(n_39068), .Z(n_37811
		));
	notech_reg to_acu0_reg_4(.CP(n_62244), .D(n_37817), .CD(n_61693), .Q(to_acu0
		[4]));
	notech_mux2 i_45834(.S(n_55689), .A(to_acu0[4]), .B(n_39069), .Z(n_37817
		));
	notech_ao4 i_132474472(.A(n_59082), .B(n_40675), .C(n_2025), .D(n_39339)
		, .Z(n_1632));
	notech_reg to_acu0_reg_5(.CP(n_62244), .D(n_37823), .CD(n_61696), .Q(to_acu0
		[5]));
	notech_mux2 i_45842(.S(n_55689), .A(to_acu0[5]), .B(n_40508), .Z(n_37823
		));
	notech_reg to_acu0_reg_6(.CP(n_62244), .D(n_37829), .CD(n_61696), .Q(to_acu0
		[6]));
	notech_mux2 i_45850(.S(n_55689), .A(to_acu0[6]), .B(n_39070), .Z(n_37829
		));
	notech_ao4 i_132674470(.A(n_59082), .B(n_40676), .C(n_2025), .D(n_39341)
		, .Z(n_1630));
	notech_reg to_acu0_reg_7(.CP(n_62244), .D(n_37835), .CD(n_61696), .Q(to_acu0
		[7]));
	notech_mux2 i_45858(.S(n_55689), .A(to_acu0[7]), .B(n_39071), .Z(n_37835
		));
	notech_reg to_acu0_reg_8(.CP(n_62244), .D(n_37841), .CD(n_61693), .Q(to_acu0
		[8]));
	notech_mux2 i_45866(.S(n_55689), .A(to_acu0[8]), .B(n_39072), .Z(n_37841
		));
	notech_ao4 i_132874468(.A(n_59084), .B(n_40677), .C(n_2025), .D(n_39342)
		, .Z(n_1628));
	notech_reg to_acu0_reg_9(.CP(n_62241), .D(n_37847), .CD(n_61696), .Q(to_acu0
		[9]));
	notech_mux2 i_45874(.S(n_55689), .A(to_acu0[9]), .B(n_40509), .Z(n_37847
		));
	notech_reg to_acu0_reg_10(.CP(n_62241), .D(n_37853), .CD(n_61693), .Q(to_acu0
		[10]));
	notech_mux2 i_45882(.S(n_55689), .A(to_acu0[10]), .B(n_39073), .Z(n_37853
		));
	notech_ao4 i_133074466(.A(n_59084), .B(n_40678), .C(n_2025), .D(n_39344)
		, .Z(n_1626));
	notech_reg to_acu0_reg_11(.CP(n_62241), .D(n_37859), .CD(n_61693), .Q(to_acu0
		[11]));
	notech_mux2 i_45890(.S(n_55703), .A(to_acu0[11]), .B(n_40510), .Z(n_37859
		));
	notech_reg to_acu0_reg_12(.CP(n_62241), .D(n_37865), .CD(n_61693), .Q(to_acu0
		[12]));
	notech_mux2 i_45898(.S(n_55717), .A(to_acu0[12]), .B(n_40511), .Z(n_37865
		));
	notech_ao4 i_133274464(.A(n_59079), .B(n_40679), .C(n_2025), .D(n_39345)
		, .Z(n_1624));
	notech_reg to_acu0_reg_13(.CP(n_62241), .D(n_37871), .CD(n_61693), .Q(to_acu0
		[13]));
	notech_mux2 i_45906(.S(n_55717), .A(to_acu0[13]), .B(n_40512), .Z(n_37871
		));
	notech_reg to_acu0_reg_14(.CP(n_62241), .D(n_37877), .CD(n_61693), .Q(to_acu0
		[14]));
	notech_mux2 i_45914(.S(n_55717), .A(to_acu0[14]), .B(n_40513), .Z(n_37877
		));
	notech_ao4 i_133474462(.A(n_59079), .B(n_40680), .C(n_2025), .D(n_39347)
		, .Z(n_1622));
	notech_reg to_acu0_reg_15(.CP(n_62241), .D(n_37883), .CD(n_61693), .Q(to_acu0
		[15]));
	notech_mux2 i_45922(.S(n_55717), .A(to_acu0[15]), .B(n_40514), .Z(n_37883
		));
	notech_reg to_acu0_reg_16(.CP(n_62241), .D(n_37889), .CD(n_61693), .Q(to_acu0
		[16]));
	notech_mux2 i_45930(.S(n_55717), .A(to_acu0[16]), .B(n_39197), .Z(n_37889
		));
	notech_ao4 i_133674460(.A(n_59079), .B(n_40681), .C(n_2025), .D(n_39348)
		, .Z(n_1620));
	notech_reg to_acu0_reg_17(.CP(n_62241), .D(n_37895), .CD(n_61693), .Q(to_acu0
		[17]));
	notech_mux2 i_45938(.S(n_55717), .A(to_acu0[17]), .B(n_39199), .Z(n_37895
		));
	notech_reg to_acu0_reg_18(.CP(n_62241), .D(n_37901), .CD(n_61693), .Q(to_acu0
		[18]));
	notech_mux2 i_45946(.S(n_55717), .A(to_acu0[18]), .B(n_40515), .Z(n_37901
		));
	notech_ao4 i_133874458(.A(n_59079), .B(n_40682), .C(n_2025), .D(n_39350)
		, .Z(n_1618));
	notech_reg to_acu0_reg_19(.CP(n_62241), .D(n_37907), .CD(n_61693), .Q(to_acu0
		[19]));
	notech_mux2 i_45954(.S(n_55717), .A(to_acu0[19]), .B(n_39201), .Z(n_37907
		));
	notech_ao4 i_133974457(.A(n_59001), .B(n_39786), .C(n_59079), .D(n_40683
		), .Z(n_1617));
	notech_reg to_acu0_reg_20(.CP(n_62246), .D(n_37913), .CD(n_61693), .Q(to_acu0
		[20]));
	notech_mux2 i_45962(.S(n_55712), .A(to_acu0[20]), .B(n_39203), .Z(n_37913
		));
	notech_ao4 i_134074456(.A(n_59001), .B(n_39788), .C(n_59079), .D(n_40684
		), .Z(n_1616));
	notech_reg to_acu0_reg_21(.CP(n_62246), .D(n_37919), .CD(n_61698), .Q(to_acu0
		[21]));
	notech_mux2 i_45970(.S(n_55717), .A(to_acu0[21]), .B(n_40516), .Z(n_37919
		));
	notech_ao4 i_134174455(.A(n_59001), .B(n_39790), .C(n_59079), .D(n_40685
		), .Z(n_1615));
	notech_reg to_acu0_reg_22(.CP(n_62246), .D(n_37925), .CD(n_61698), .Q(to_acu0
		[22]));
	notech_mux2 i_45978(.S(n_55712), .A(to_acu0[22]), .B(n_40517), .Z(n_37925
		));
	notech_ao4 i_134274454(.A(n_59001), .B(n_39793), .C(n_59079), .D(n_40687
		), .Z(n_1614));
	notech_reg to_acu0_reg_23(.CP(n_62244), .D(n_37931), .CD(n_61696), .Q(to_acu0
		[23]));
	notech_mux2 i_45986(.S(n_55712), .A(to_acu0[23]), .B(n_39205), .Z(n_37931
		));
	notech_ao4 i_134374453(.A(n_59004), .B(n_39795), .C(n_59082), .D(n_40688
		), .Z(n_1613));
	notech_reg to_acu0_reg_24(.CP(n_62244), .D(n_37937), .CD(n_61696), .Q(to_acu0
		[24]));
	notech_mux2 i_45994(.S(n_55717), .A(to_acu0[24]), .B(n_39207), .Z(n_37937
		));
	notech_ao4 i_134474452(.A(n_59004), .B(n_39797), .C(n_59082), .D(n_40689
		), .Z(n_1612));
	notech_reg to_acu0_reg_25(.CP(n_62246), .D(n_37943), .CD(n_61696), .Q(to_acu0
		[25]));
	notech_mux2 i_46002(.S(n_55717), .A(to_acu0[25]), .B(n_39209), .Z(n_37943
		));
	notech_ao4 i_134574451(.A(n_59004), .B(n_39799), .C(n_59082), .D(n_40690
		), .Z(n_1611));
	notech_reg to_acu0_reg_26(.CP(n_62246), .D(n_37949), .CD(n_61698), .Q(to_acu0
		[26]));
	notech_mux2 i_46010(.S(n_55717), .A(to_acu0[26]), .B(n_39211), .Z(n_37949
		));
	notech_ao4 i_134674450(.A(n_59004), .B(n_39801), .C(n_59082), .D(n_40691
		), .Z(n_1610));
	notech_reg to_acu0_reg_27(.CP(n_62246), .D(n_37955), .CD(n_61698), .Q(to_acu0
		[27]));
	notech_mux2 i_46018(.S(n_55717), .A(to_acu0[27]), .B(n_39213), .Z(n_37955
		));
	notech_ao4 i_134774449(.A(n_59001), .B(n_39803), .C(n_59082), .D(n_40692
		), .Z(n_1609));
	notech_reg to_acu0_reg_28(.CP(n_62246), .D(n_37961), .CD(n_61698), .Q(to_acu0
		[28]));
	notech_mux2 i_46026(.S(n_55717), .A(to_acu0[28]), .B(n_39215), .Z(n_37961
		));
	notech_ao4 i_134874448(.A(n_59004), .B(n_39805), .C(n_59082), .D(n_40693
		), .Z(n_1608));
	notech_reg to_acu0_reg_29(.CP(n_62246), .D(n_37967), .CD(n_61698), .Q(to_acu0
		[29]));
	notech_mux2 i_46034(.S(\nbus_13534[0] ), .A(to_acu0[29]), .B(n_39217), .Z
		(n_37967));
	notech_ao4 i_134974447(.A(n_59004), .B(n_39807), .C(n_59082), .D(n_40694
		), .Z(n_1607));
	notech_reg to_acu0_reg_30(.CP(n_62244), .D(n_37973), .CD(n_61698), .Q(to_acu0
		[30]));
	notech_mux2 i_46042(.S(\nbus_13534[0] ), .A(to_acu0[30]), .B(n_39219), .Z
		(n_37973));
	notech_reg to_acu0_reg_31(.CP(n_62244), .D(n_37979), .CD(n_61696), .Q(to_acu0
		[31]));
	notech_mux2 i_46050(.S(\nbus_13534[0] ), .A(to_acu0[31]), .B(n_39221), .Z
		(n_37979));
	notech_reg to_acu0_reg_32(.CP(n_62244), .D(n_37985), .CD(n_61696), .Q(to_acu0
		[32]));
	notech_mux2 i_46058(.S(\nbus_13534[0] ), .A(to_acu0[32]), .B(n_39223), .Z
		(n_37985));
	notech_reg to_acu0_reg_33(.CP(n_62244), .D(n_37991), .CD(n_61696), .Q(to_acu0
		[33]));
	notech_mux2 i_46066(.S(\nbus_13534[0] ), .A(to_acu0[33]), .B(n_39225), .Z
		(n_37991));
	notech_reg to_acu0_reg_34(.CP(n_62244), .D(n_37997), .CD(n_61696), .Q(to_acu0
		[34]));
	notech_mux2 i_46074(.S(\nbus_13534[0] ), .A(to_acu0[34]), .B(n_39227), .Z
		(n_37997));
	notech_reg to_acu0_reg_35(.CP(n_62244), .D(n_38003), .CD(n_61696), .Q(to_acu0
		[35]));
	notech_mux2 i_46082(.S(\nbus_13534[0] ), .A(to_acu0[35]), .B(n_39229), .Z
		(n_38003));
	notech_reg to_acu0_reg_36(.CP(n_62244), .D(n_38009), .CD(n_61696), .Q(to_acu0
		[36]));
	notech_mux2 i_46090(.S(\nbus_13534[0] ), .A(to_acu0[36]), .B(n_39231), .Z
		(n_38009));
	notech_reg to_acu0_reg_37(.CP(n_62244), .D(n_38015), .CD(n_61696), .Q(to_acu0
		[37]));
	notech_mux2 i_46098(.S(\nbus_13534[0] ), .A(to_acu0[37]), .B(n_39233), .Z
		(n_38015));
	notech_reg to_acu0_reg_38(.CP(n_62244), .D(n_38021), .CD(n_61696), .Q(to_acu0
		[38]));
	notech_mux2 i_46106(.S(\nbus_13534[0] ), .A(to_acu0[38]), .B(n_39235), .Z
		(n_38021));
	notech_and4 i_144274354(.A(n_60059), .B(n_2228), .C(n_1597), .D(n_1586),
		 .Z(n_1600));
	notech_reg to_acu0_reg_39(.CP(n_62244), .D(n_38027), .CD(n_61696), .Q(to_acu0
		[39]));
	notech_mux2 i_46114(.S(n_55717), .A(to_acu0[39]), .B(n_111395808), .Z(n_38027
		));
	notech_reg to_acu0_reg_40(.CP(n_62244), .D(n_38033), .CD(n_61696), .Q(to_acu0
		[40]));
	notech_mux2 i_46122(.S(\nbus_13534[0] ), .A(to_acu0[40]), .B(n_39237), .Z
		(n_38033));
	notech_reg to_acu0_reg_41(.CP(n_62211), .D(n_38039), .CD(n_61696), .Q(to_acu0
		[41]));
	notech_mux2 i_46130(.S(\nbus_13534[0] ), .A(to_acu0[41]), .B(n_39239), .Z
		(n_38039));
	notech_ao4 i_19375779(.A(n_224396466), .B(n_40501), .C(n_39195), .D(n_40502
		), .Z(n_1597));
	notech_reg to_acu0_reg_42(.CP(n_62211), .D(n_38045), .CD(n_61680), .Q(to_acu0
		[42]));
	notech_mux2 i_46138(.S(\nbus_13534[0] ), .A(to_acu0[42]), .B(n_39241), .Z
		(n_38045));
	notech_reg to_acu0_reg_43(.CP(n_62211), .D(n_38051), .CD(n_61660), .Q(to_acu0
		[43]));
	notech_mux2 i_46146(.S(\nbus_13534[0] ), .A(to_acu0[43]), .B(n_40518), .Z
		(n_38051));
	notech_and2 i_19075780(.A(n_40937), .B(n_59975), .Z(n_16151033));
	notech_reg to_acu0_reg_44(.CP(n_62208), .D(n_38057), .CD(n_61663), .Q(to_acu0
		[44]));
	notech_mux2 i_46154(.S(\nbus_13534[0] ), .A(to_acu0[44]), .B(n_40519), .Z
		(n_38057));
	notech_ao4 i_144574351(.A(n_3274), .B(n_1511), .C(n_1510), .D(n_18051052
		), .Z(n_1595));
	notech_reg to_acu0_reg_45(.CP(n_62211), .D(n_38063), .CD(n_61660), .Q(to_acu0
		[45]));
	notech_mux2 i_46162(.S(n_55708), .A(to_acu0[45]), .B(n_39243), .Z(n_38063
		));
	notech_reg to_acu0_reg_46(.CP(n_62211), .D(n_38069), .CD(n_61660), .Q(to_acu0
		[46]));
	notech_mux2 i_46170(.S(n_55708), .A(to_acu0[46]), .B(n_39245), .Z(n_38069
		));
	notech_nand2 i_144774349(.A(n_227296437), .B(n_2887), .Z(n_1593));
	notech_reg to_acu0_reg_47(.CP(n_62211), .D(n_38075), .CD(n_61660), .Q(to_acu0
		[47]));
	notech_mux2 i_46178(.S(n_55708), .A(to_acu0[47]), .B(n_39247), .Z(n_38075
		));
	notech_reg to_acu0_reg_48(.CP(n_62211), .D(n_38081), .CD(n_61663), .Q(to_acu0
		[48]));
	notech_mux2 i_46186(.S(n_55708), .A(to_acu0[48]), .B(n_40521), .Z(n_38081
		));
	notech_ao4 i_144974347(.A(pg_fault), .B(n_59975), .C(n_2870), .D(n_40502
		), .Z(n_1591));
	notech_reg to_acu0_reg_49(.CP(n_62211), .D(n_38087), .CD(n_61663), .Q(to_acu0
		[49]));
	notech_mux2 i_46194(.S(n_55708), .A(to_acu0[49]), .B(n_40522), .Z(n_38087
		));
	notech_or4 i_13575783(.A(n_59653), .B(pc_req), .C(pg_fault), .D(n_223996470
		), .Z(n_18051052));
	notech_reg to_acu0_reg_50(.CP(n_62211), .D(n_38093), .CD(n_61663), .Q(to_acu0
		[50]));
	notech_mux2 i_46202(.S(n_55708), .A(to_acu0[50]), .B(n_39250), .Z(n_38093
		));
	notech_and2 i_73646(.A(n_61663), .B(n_1445), .Z(\nbus_13559[0] ));
	notech_reg to_acu0_reg_51(.CP(n_62208), .D(n_38099), .CD(n_61663), .Q(to_acu0
		[51]));
	notech_mux2 i_46210(.S(n_55708), .A(to_acu0[51]), .B(n_39253), .Z(n_38099
		));
	notech_reg to_acu0_reg_52(.CP(n_62208), .D(n_38105), .CD(n_61660), .Q(to_acu0
		[52]));
	notech_mux2 i_46218(.S(n_55708), .A(to_acu0[52]), .B(n_40523), .Z(n_38105
		));
	notech_reg to_acu0_reg_53(.CP(n_62208), .D(n_38111), .CD(n_61660), .Q(to_acu0
		[53]));
	notech_mux2 i_46226(.S(n_55703), .A(to_acu0[53]), .B(n_39256), .Z(n_38111
		));
	notech_or2 i_123174565(.A(n_2025), .B(n_40501), .Z(n_1588));
	notech_reg to_acu0_reg_54(.CP(n_62208), .D(n_38117), .CD(n_61660), .Q(to_acu0
		[54]));
	notech_mux2 i_46234(.S(n_55703), .A(to_acu0[54]), .B(n_39259), .Z(n_38117
		));
	notech_reg to_acu0_reg_55(.CP(n_62208), .D(n_38123), .CD(n_61660), .Q(to_acu0
		[55]));
	notech_mux2 i_46242(.S(n_55703), .A(to_acu0[55]), .B(n_40524), .Z(n_38123
		));
	notech_or4 i_122574571(.A(n_57101), .B(pg_fault), .C(pc_req), .D(n_1507)
		, .Z(n_1586));
	notech_reg to_acu0_reg_56(.CP(n_62208), .D(n_38129), .CD(n_61660), .Q(to_acu0
		[56]));
	notech_mux2 i_46250(.S(n_55703), .A(to_acu0[56]), .B(n_40525), .Z(n_38129
		));
	notech_ao3 i_2881(.A(n_1504), .B(n_40498), .C(n_2876), .Z(useq_ptr[3])
		);
	notech_reg to_acu0_reg_57(.CP(n_62208), .D(n_38135), .CD(n_61660), .Q(to_acu0
		[57]));
	notech_mux2 i_46258(.S(n_55708), .A(to_acu0[57]), .B(n_40526), .Z(n_38135
		));
	notech_and3 i_2882(.A(n_40498), .B(n_1504), .C(n_2878), .Z(useq_ptr[2])
		);
	notech_reg to_acu0_reg_58(.CP(n_62208), .D(n_38141), .CD(n_61660), .Q(to_acu0
		[58]));
	notech_mux2 i_46266(.S(n_55708), .A(to_acu0[58]), .B(n_39074), .Z(n_38141
		));
	notech_and3 i_2883(.A(n_40498), .B(n_1504), .C(n_2880), .Z(useq_ptr[1])
		);
	notech_reg to_acu0_reg_59(.CP(n_62208), .D(n_38147), .CD(n_61660), .Q(to_acu0
		[59]));
	notech_mux2 i_46274(.S(n_55703), .A(to_acu0[59]), .B(n_40527), .Z(n_38147
		));
	notech_and3 i_2884(.A(n_40498), .B(n_1504), .C(n_2206), .Z(useq_ptr[0])
		);
	notech_reg to_acu0_reg_60(.CP(n_62208), .D(n_38153), .CD(n_61660), .Q(to_acu0
		[60]));
	notech_mux2 i_46282(.S(n_55703), .A(to_acu0[60]), .B(n_40528), .Z(n_38153
		));
	notech_and3 i_3075(.A(n_60042), .B(lenpc2[26]), .C(n_59975), .Z(n_44259)
		);
	notech_reg to_acu0_reg_61(.CP(n_62208), .D(n_38159), .CD(n_61660), .Q(to_acu0
		[61]));
	notech_mux2 i_46290(.S(n_55708), .A(to_acu0[61]), .B(n_40529), .Z(n_38159
		));
	notech_and3 i_3073(.A(n_60042), .B(lenpc2[24]), .C(n_59975), .Z(n_44247)
		);
	notech_reg to_acu0_reg_62(.CP(n_62213), .D(n_38165), .CD(n_61660), .Q(to_acu0
		[62]));
	notech_mux2 i_46298(.S(n_55712), .A(to_acu0[62]), .B(n_39262), .Z(n_38165
		));
	notech_and3 i_3068(.A(n_60042), .B(lenpc2[19]), .C(n_59980), .Z(n_44217)
		);
	notech_reg to_acu0_reg_63(.CP(n_62213), .D(n_38171), .CD(n_61665), .Q(to_acu0
		[63]));
	notech_mux2 i_46306(.S(n_55712), .A(to_acu0[63]), .B(n_40530), .Z(n_38171
		));
	notech_and3 i_3061(.A(n_60042), .B(lenpc2[12]), .C(n_59980), .Z(n_44175)
		);
	notech_reg to_acu0_reg_64(.CP(n_62213), .D(n_38177), .CD(n_61665), .Q(to_acu0
		[64]));
	notech_mux2 i_46314(.S(n_55712), .A(to_acu0[64]), .B(n_40531), .Z(n_38177
		));
	notech_and3 i_3060(.A(n_60042), .B(lenpc2[11]), .C(n_59980), .Z(n_44169)
		);
	notech_reg to_acu0_reg_65(.CP(n_62213), .D(n_38183), .CD(n_61665), .Q(to_acu0
		[65]));
	notech_mux2 i_46322(.S(n_55712), .A(to_acu0[65]), .B(n_40532), .Z(n_38183
		));
	notech_and3 i_3059(.A(n_60042), .B(lenpc2[10]), .C(n_59975), .Z(n_44163)
		);
	notech_reg to_acu0_reg_66(.CP(n_62213), .D(n_38189), .CD(n_61665), .Q(to_acu0
		[66]));
	notech_mux2 i_46330(.S(n_55712), .A(to_acu0[66]), .B(n_40533), .Z(n_38189
		));
	notech_and3 i_3058(.A(n_60042), .B(lenpc2[9]), .C(n_59975), .Z(n_44157)
		);
	notech_reg to_acu0_reg_67(.CP(n_62213), .D(n_38195), .CD(n_61665), .Q(to_acu0
		[67]));
	notech_mux2 i_46338(.S(n_55712), .A(to_acu0[67]), .B(n_40535), .Z(n_38195
		));
	notech_and3 i_3056(.A(n_60042), .B(lenpc2[7]), .C(n_59975), .Z(n_44145)
		);
	notech_reg to_acu0_reg_68(.CP(n_62213), .D(n_38201), .CD(n_61665), .Q(to_acu0
		[68]));
	notech_mux2 i_46346(.S(n_55712), .A(to_acu0[68]), .B(n_40536), .Z(n_38201
		));
	notech_reg to_acu0_reg_69(.CP(n_62213), .D(n_38207), .CD(n_61665), .Q(to_acu0
		[69]));
	notech_mux2 i_46354(.S(n_55712), .A(to_acu0[69]), .B(n_40537), .Z(n_38207
		));
	notech_reg to_acu0_reg_70(.CP(n_62213), .D(n_38213), .CD(n_61665), .Q(to_acu0
		[70]));
	notech_mux2 i_46362(.S(n_55708), .A(to_acu0[70]), .B(n_40538), .Z(n_38213
		));
	notech_reg to_acu0_reg_71(.CP(n_62213), .D(n_38219), .CD(n_61665), .Q(to_acu0
		[71]));
	notech_mux2 i_46370(.S(n_55708), .A(to_acu0[71]), .B(n_40539), .Z(n_38219
		));
	notech_reg to_acu0_reg_72(.CP(n_62213), .D(n_38225), .CD(n_61665), .Q(to_acu0
		[72]));
	notech_mux2 i_46378(.S(n_55708), .A(to_acu0[72]), .B(n_40540), .Z(n_38225
		));
	notech_reg to_acu0_reg_73(.CP(n_62211), .D(n_38231), .CD(n_61663), .Q(to_acu0
		[73]));
	notech_mux2 i_46386(.S(n_55708), .A(to_acu0[73]), .B(n_40541), .Z(n_38231
		));
	notech_reg to_acu0_reg_74(.CP(n_62211), .D(n_38237), .CD(n_61663), .Q(to_acu0
		[74]));
	notech_mux2 i_46394(.S(n_55712), .A(to_acu0[74]), .B(n_40542), .Z(n_38237
		));
	notech_reg to_acu0_reg_75(.CP(n_62211), .D(n_38243), .CD(n_61663), .Q(to_acu0
		[75]));
	notech_mux2 i_46402(.S(n_55712), .A(to_acu0[75]), .B(n_40543), .Z(n_38243
		));
	notech_reg to_acu0_reg_76(.CP(n_62211), .D(n_38249), .CD(n_61663), .Q(to_acu0
		[76]));
	notech_mux2 i_46410(.S(n_55712), .A(to_acu0[76]), .B(n_40544), .Z(n_38249
		));
	notech_reg to_acu0_reg_77(.CP(n_62211), .D(n_38255), .CD(n_61663), .Q(to_acu0
		[77]));
	notech_mux2 i_46418(.S(n_55712), .A(to_acu0[77]), .B(n_40545), .Z(n_38255
		));
	notech_reg to_acu0_reg_78(.CP(n_62211), .D(n_38261), .CD(n_61663), .Q(to_acu0
		[78]));
	notech_mux2 i_46426(.S(n_55656), .A(to_acu0[78]), .B(n_40546), .Z(n_38261
		));
	notech_reg to_acu0_reg_79(.CP(n_62213), .D(n_38267), .CD(n_61663), .Q(to_acu0
		[79]));
	notech_mux2 i_46434(.S(n_55656), .A(to_acu0[79]), .B(n_40547), .Z(n_38267
		));
	notech_reg to_acu0_reg_80(.CP(n_62211), .D(n_38273), .CD(n_61663), .Q(to_acu0
		[80]));
	notech_mux2 i_46442(.S(n_55656), .A(to_acu0[80]), .B(n_40548), .Z(n_38273
		));
	notech_reg to_acu0_reg_81(.CP(n_62211), .D(n_38279), .CD(n_61663), .Q(to_acu0
		[81]));
	notech_mux2 i_46450(.S(n_55656), .A(to_acu0[81]), .B(n_40549), .Z(n_38279
		));
	notech_reg to_acu0_reg_82(.CP(n_62211), .D(n_38285), .CD(n_61663), .Q(to_acu0
		[82]));
	notech_mux2 i_46458(.S(n_55656), .A(to_acu0[82]), .B(n_40550), .Z(n_38285
		));
	notech_reg to_acu0_reg_83(.CP(n_62208), .D(n_38291), .CD(n_61663), .Q(to_acu0
		[83]));
	notech_mux2 i_46466(.S(n_55656), .A(to_acu0[83]), .B(n_40551), .Z(n_38291
		));
	notech_reg to_acu0_reg_84(.CP(n_62203), .D(n_38297), .CD(n_61655), .Q(to_acu0
		[84]));
	notech_mux2 i_46474(.S(n_55656), .A(to_acu0[84]), .B(n_40552), .Z(n_38297
		));
	notech_reg to_acu0_reg_85(.CP(n_62203), .D(n_38303), .CD(n_61655), .Q(to_acu0
		[85]));
	notech_mux2 i_46482(.S(n_55656), .A(to_acu0[85]), .B(n_40553), .Z(n_38303
		));
	notech_reg to_acu0_reg_86(.CP(n_62203), .D(n_38309), .CD(n_61655), .Q(to_acu0
		[86]));
	notech_mux2 i_46490(.S(n_55652), .A(to_acu0[86]), .B(n_40554), .Z(n_38309
		));
	notech_reg to_acu0_reg_87(.CP(n_62203), .D(n_38315), .CD(n_61655), .Q(to_acu0
		[87]));
	notech_mux2 i_46498(.S(n_55652), .A(to_acu0[87]), .B(n_40555), .Z(n_38315
		));
	notech_reg to_acu0_reg_88(.CP(n_62203), .D(n_38321), .CD(n_61655), .Q(to_acu0
		[88]));
	notech_mux2 i_46506(.S(n_55652), .A(to_acu0[88]), .B(n_40556), .Z(n_38321
		));
	notech_reg to_acu0_reg_89(.CP(n_62206), .D(n_38327), .CD(n_61655), .Q(to_acu0
		[89]));
	notech_mux2 i_46514(.S(n_55652), .A(to_acu0[89]), .B(n_40557), .Z(n_38327
		));
	notech_reg to_acu0_reg_90(.CP(n_62206), .D(n_38333), .CD(n_61655), .Q(to_acu0
		[90]));
	notech_mux2 i_46522(.S(n_55652), .A(to_acu0[90]), .B(n_39265), .Z(n_38333
		));
	notech_reg to_acu0_reg_91(.CP(n_62203), .D(n_38339), .CD(n_61655), .Q(to_acu0
		[91]));
	notech_mux2 i_46530(.S(n_55652), .A(to_acu0[91]), .B(n_40558), .Z(n_38339
		));
	notech_reg to_acu0_reg_92(.CP(n_62203), .D(n_38345), .CD(n_61655), .Q(to_acu0
		[92]));
	notech_mux2 i_46538(.S(n_55652), .A(to_acu0[92]), .B(n_39268), .Z(n_38345
		));
	notech_nand3 i_20575584(.A(n_2885), .B(inst_deco1[87]), .C(n_59017), .Z(n_1561
		));
	notech_reg to_acu0_reg_93(.CP(n_62203), .D(n_38351), .CD(n_61655), .Q(to_acu0
		[93]));
	notech_mux2 i_46546(.S(n_55652), .A(to_acu0[93]), .B(n_40560), .Z(n_38351
		));
	notech_reg to_acu0_reg_94(.CP(n_62203), .D(n_38357), .CD(n_61655), .Q(to_acu0
		[94]));
	notech_mux2 i_46554(.S(n_55656), .A(to_acu0[94]), .B(n_39271), .Z(n_38357
		));
	notech_reg to_acu0_reg_95(.CP(n_62203), .D(n_38363), .CD(n_61655), .Q(to_acu0
		[95]));
	notech_mux2 i_46562(.S(n_55661), .A(to_acu0[95]), .B(n_39274), .Z(n_38363
		));
	notech_nand3 i_20175587(.A(n_2885), .B(inst_deco1[86]), .C(n_59017), .Z(n_1558
		));
	notech_reg to_acu0_reg_96(.CP(n_62203), .D(n_38369), .CD(n_61655), .Q(to_acu0
		[96]));
	notech_mux2 i_46570(.S(n_55661), .A(to_acu0[96]), .B(n_39277), .Z(n_38369
		));
	notech_reg to_acu0_reg_97(.CP(n_62203), .D(n_38375), .CD(n_61653), .Q(to_acu0
		[97]));
	notech_mux2 i_46578(.S(n_55661), .A(to_acu0[97]), .B(n_39280), .Z(n_38375
		));
	notech_reg to_acu0_reg_98(.CP(n_62201), .D(n_38381), .CD(n_61653), .Q(to_acu0
		[98]));
	notech_mux2 i_46586(.S(n_55661), .A(to_acu0[98]), .B(n_39283), .Z(n_38381
		));
	notech_nand3 i_19775590(.A(n_2885), .B(inst_deco1[85]), .C(n_59017), .Z(n_1555
		));
	notech_reg to_acu0_reg_99(.CP(n_62203), .D(n_38387), .CD(n_61653), .Q(to_acu0
		[99]));
	notech_mux2 i_46594(.S(n_55661), .A(to_acu0[99]), .B(n_39286), .Z(n_38387
		));
	notech_reg to_acu0_reg_100(.CP(n_62203), .D(n_38393), .CD(n_61655), .Q(to_acu0
		[100]));
	notech_mux2 i_46602(.S(n_55661), .A(to_acu0[100]), .B(n_39289), .Z(n_38393
		));
	notech_reg to_acu0_reg_101(.CP(n_62203), .D(n_38399), .CD(n_61655), .Q(to_acu0
		[101]));
	notech_mux2 i_46610(.S(n_55661), .A(to_acu0[101]), .B(n_39292), .Z(n_38399
		));
	notech_nand3 i_19475593(.A(n_2885), .B(inst_deco1[84]), .C(n_59017), .Z(n_1552
		));
	notech_reg to_acu0_reg_102(.CP(n_62203), .D(n_38405), .CD(n_61655), .Q(to_acu0
		[102]));
	notech_mux2 i_46618(.S(n_55661), .A(to_acu0[102]), .B(n_39295), .Z(n_38405
		));
	notech_reg to_acu0_reg_103(.CP(n_62203), .D(n_38411), .CD(n_61655), .Q(to_acu0
		[103]));
	notech_mux2 i_46626(.S(n_55656), .A(to_acu0[103]), .B(n_39298), .Z(n_38411
		));
	notech_reg to_acu0_reg_104(.CP(n_62203), .D(n_38417), .CD(n_61655), .Q(to_acu0
		[104]));
	notech_mux2 i_46634(.S(n_55656), .A(to_acu0[104]), .B(n_39301), .Z(n_38417
		));
	notech_nand3 i_18975596(.A(n_2885), .B(inst_deco1[83]), .C(n_59017), .Z(n_1549
		));
	notech_reg to_acu0_reg_105(.CP(n_62206), .D(n_38423), .CD(n_61658), .Q(to_acu0
		[105]));
	notech_mux2 i_46642(.S(n_55656), .A(to_acu0[105]), .B(n_39304), .Z(n_38423
		));
	notech_reg to_acu0_reg_106(.CP(n_62206), .D(n_38429), .CD(n_61658), .Q(to_acu0
		[106]));
	notech_mux2 i_46650(.S(n_55656), .A(to_acu0[106]), .B(n_39307), .Z(n_38429
		));
	notech_reg to_acu0_reg_107(.CP(n_62206), .D(n_38435), .CD(n_61658), .Q(to_acu0
		[107]));
	notech_mux2 i_46658(.S(n_55661), .A(to_acu0[107]), .B(n_39075), .Z(n_38435
		));
	notech_nand3 i_18675599(.A(n_2885), .B(inst_deco1[82]), .C(n_59017), .Z(n_1546
		));
	notech_reg to_acu0_reg_108(.CP(n_62206), .D(n_38441), .CD(n_61658), .Q(to_acu0
		[108]));
	notech_mux2 i_46666(.S(n_55661), .A(to_acu0[108]), .B(n_39310), .Z(n_38441
		));
	notech_reg to_acu0_reg_109(.CP(n_62206), .D(n_38447), .CD(n_61658), .Q(to_acu0
		[109]));
	notech_mux2 i_46674(.S(n_55656), .A(to_acu0[109]), .B(n_39076), .Z(n_38447
		));
	notech_reg to_acu0_reg_110(.CP(n_62208), .D(n_38453), .CD(n_61660), .Q(to_acu0
		[110]));
	notech_mux2 i_46682(.S(n_55656), .A(to_acu0[110]), .B(n_39077), .Z(n_38453
		));
	notech_nand3 i_18375602(.A(n_2885), .B(inst_deco1[81]), .C(n_59017), .Z(n_1543
		));
	notech_reg to_acu0_reg_111(.CP(n_62208), .D(n_38459), .CD(n_61660), .Q(to_acu0
		[111]));
	notech_mux2 i_46690(.S(n_55643), .A(to_acu0[111]), .B(n_39078), .Z(n_38459
		));
	notech_reg to_acu0_reg_112(.CP(n_62208), .D(n_38465), .CD(n_61660), .Q(to_acu0
		[112]));
	notech_mux2 i_46698(.S(n_55643), .A(to_acu0[112]), .B(n_39079), .Z(n_38465
		));
	notech_reg to_acu0_reg_113(.CP(n_62208), .D(n_38471), .CD(n_61658), .Q(to_acu0
		[113]));
	notech_mux2 i_46706(.S(n_55643), .A(to_acu0[113]), .B(n_39080), .Z(n_38471
		));
	notech_nand3 i_18075605(.A(n_2885), .B(inst_deco1[80]), .C(n_59017), .Z(n_1540
		));
	notech_reg to_acu0_reg_114(.CP(n_62208), .D(n_38477), .CD(n_61658), .Q(to_acu0
		[114]));
	notech_mux2 i_46714(.S(n_55643), .A(to_acu0[114]), .B(n_39081), .Z(n_38477
		));
	notech_reg to_acu0_reg_115(.CP(n_62206), .D(n_38483), .CD(n_61658), .Q(to_acu0
		[115]));
	notech_mux2 i_46722(.S(n_55647), .A(to_acu0[115]), .B(n_39082), .Z(n_38483
		));
	notech_reg to_acu0_reg_116(.CP(n_62206), .D(n_38489), .CD(n_61658), .Q(to_acu0
		[116]));
	notech_mux2 i_46730(.S(n_55647), .A(to_acu0[116]), .B(n_39083), .Z(n_38489
		));
	notech_reg to_acu0_reg_117(.CP(n_62206), .D(n_38495), .CD(n_61658), .Q(to_acu0
		[117]));
	notech_mux2 i_46738(.S(n_55647), .A(to_acu0[117]), .B(n_39084), .Z(n_38495
		));
	notech_reg to_acu0_reg_118(.CP(n_62206), .D(n_38501), .CD(n_61658), .Q(to_acu0
		[118]));
	notech_mux2 i_46746(.S(n_55647), .A(to_acu0[118]), .B(n_39085), .Z(n_38501
		));
	notech_reg to_acu0_reg_119(.CP(n_62206), .D(n_38507), .CD(n_61658), .Q(to_acu0
		[119]));
	notech_mux2 i_46754(.S(n_55643), .A(to_acu0[119]), .B(n_39086), .Z(n_38507
		));
	notech_reg to_acu0_reg_120(.CP(n_62206), .D(n_38513), .CD(n_61658), .Q(to_acu0
		[120]));
	notech_mux2 i_46762(.S(n_55643), .A(to_acu0[120]), .B(n_39087), .Z(n_38513
		));
	notech_reg to_acu0_reg_121(.CP(n_62206), .D(n_38519), .CD(n_61658), .Q(to_acu0
		[121]));
	notech_mux2 i_46770(.S(n_55643), .A(to_acu0[121]), .B(n_39088), .Z(n_38519
		));
	notech_reg to_acu0_reg_122(.CP(n_62206), .D(n_38525), .CD(n_61658), .Q(to_acu0
		[122]));
	notech_mux2 i_46778(.S(n_55643), .A(to_acu0[122]), .B(n_40561), .Z(n_38525
		));
	notech_reg to_acu0_reg_123(.CP(n_62206), .D(n_38531), .CD(n_61658), .Q(to_acu0
		[123]));
	notech_mux2 i_46786(.S(n_55643), .A(to_acu0[123]), .B(n_40562), .Z(n_38531
		));
	notech_reg to_acu0_reg_124(.CP(n_62206), .D(n_38537), .CD(n_61658), .Q(to_acu0
		[124]));
	notech_mux2 i_46794(.S(n_55643), .A(to_acu0[124]), .B(n_39089), .Z(n_38537
		));
	notech_reg to_acu0_reg_125(.CP(n_62206), .D(n_38543), .CD(n_61658), .Q(to_acu0
		[125]));
	notech_mux2 i_46802(.S(n_55643), .A(to_acu0[125]), .B(n_40563), .Z(n_38543
		));
	notech_reg to_acu0_reg_126(.CP(n_62223), .D(n_38549), .CD(n_61665), .Q(to_acu0
		[126]));
	notech_mux2 i_46810(.S(n_55643), .A(to_acu0[126]), .B(n_40564), .Z(n_38549
		));
	notech_reg to_acu0_reg_127(.CP(n_62223), .D(n_38555), .CD(n_61675), .Q(to_acu0
		[127]));
	notech_mux2 i_46818(.S(n_55647), .A(to_acu0[127]), .B(n_40565), .Z(n_38555
		));
	notech_reg to_acu0_reg_128(.CP(n_62223), .D(n_38561), .CD(n_61675), .Q(to_acu0
		[128]));
	notech_mux2 i_46826(.S(n_55652), .A(to_acu0[128]), .B(n_40566), .Z(n_38561
		));
	notech_reg to_acu0_reg_129(.CP(n_62223), .D(n_38567), .CD(n_61675), .Q(to_acu0
		[129]));
	notech_mux2 i_46834(.S(n_55652), .A(to_acu0[129]), .B(n_40567), .Z(n_38567
		));
	notech_reg to_acu0_reg_130(.CP(n_62223), .D(n_38573), .CD(n_61675), .Q(to_acu0
		[130]));
	notech_mux2 i_46842(.S(n_55647), .A(to_acu0[130]), .B(n_39090), .Z(n_38573
		));
	notech_reg to_acu0_reg_131(.CP(n_62225), .D(n_38579), .CD(n_61675), .Q(to_acu0
		[131]));
	notech_mux2 i_46850(.S(n_55652), .A(to_acu0[131]), .B(n_39091), .Z(n_38579
		));
	notech_reg to_acu0_reg_132(.CP(n_62225), .D(n_38585), .CD(n_61677), .Q(to_acu0
		[132]));
	notech_mux2 i_46858(.S(n_55652), .A(to_acu0[132]), .B(n_39092), .Z(n_38585
		));
	notech_or4 i_124174555(.A(n_2171), .B(n_40559), .C(n_2901), .D(n_40914),
		 .Z(n_1521));
	notech_reg to_acu0_reg_133(.CP(n_62225), .D(n_38591), .CD(n_61677), .Q(to_acu0
		[133]));
	notech_mux2 i_46866(.S(n_55652), .A(to_acu0[133]), .B(n_39093), .Z(n_38591
		));
	notech_or2 i_124074556(.A(n_2837), .B(n_268594642), .Z(n_1520));
	notech_reg to_acu0_reg_134(.CP(n_62223), .D(n_38597), .CD(n_61675), .Q(to_acu0
		[134]));
	notech_mux2 i_46874(.S(n_55652), .A(to_acu0[134]), .B(n_39094), .Z(n_38597
		));
	notech_reg to_acu0_reg_135(.CP(n_62225), .D(n_38603), .CD(n_61675), .Q(to_acu0
		[135]));
	notech_mux2 i_46882(.S(n_55652), .A(to_acu0[135]), .B(n_39095), .Z(n_38603
		));
	notech_reg to_acu0_reg_136(.CP(n_62223), .D(n_38609), .CD(n_61675), .Q(to_acu0
		[136]));
	notech_mux2 i_46890(.S(n_55647), .A(to_acu0[136]), .B(n_39096), .Z(n_38609
		));
	notech_ao4 i_175774(.A(n_2225), .B(n_39143), .C(n_2837), .D(n_2960), .Z(n_1517
		));
	notech_reg to_acu0_reg_137(.CP(n_62223), .D(n_38615), .CD(n_61675), .Q(to_acu0
		[137]));
	notech_mux2 i_46898(.S(n_55647), .A(to_acu0[137]), .B(n_39097), .Z(n_38615
		));
	notech_nand2 i_123774559(.A(db67), .B(n_40589), .Z(n_1516));
	notech_reg to_acu0_reg_138(.CP(n_62223), .D(n_38621), .CD(n_61675), .Q(to_acu0
		[138]));
	notech_mux2 i_46906(.S(n_55647), .A(to_acu0[138]), .B(n_39098), .Z(n_38621
		));
	notech_or2 i_123674560(.A(n_40559), .B(n_2227), .Z(n_1515));
	notech_reg to_acu0_reg_139(.CP(n_62223), .D(n_38627), .CD(n_61675), .Q(to_acu0
		[139]));
	notech_mux2 i_46914(.S(n_55647), .A(to_acu0[139]), .B(n_39099), .Z(n_38627
		));
	notech_or4 i_123574561(.A(n_40559), .B(n_2223), .C(n_2171), .D(n_2224), 
		.Z(n_1514));
	notech_reg to_acu0_reg_140(.CP(n_62223), .D(n_38633), .CD(n_61675), .Q(to_acu0
		[140]));
	notech_mux2 i_46922(.S(n_55647), .A(to_acu0[140]), .B(n_40568), .Z(n_38633
		));
	notech_reg to_acu0_reg_141(.CP(n_62223), .D(n_38639), .CD(n_61672), .Q(to_acu0
		[141]));
	notech_mux2 i_46930(.S(n_55647), .A(to_acu0[141]), .B(n_39100), .Z(n_38639
		));
	notech_ao4 i_123374563(.A(n_2871), .B(n_2865), .C(n_2870), .D(n_1593), .Z
		(n_1512));
	notech_reg to_acu0_reg_142(.CP(n_62223), .D(n_38645), .CD(n_61675), .Q(to_acu0
		[142]));
	notech_mux2 i_46938(.S(n_55647), .A(to_acu0[142]), .B(n_40569), .Z(n_38645
		));
	notech_nor2 i_375772(.A(idx_deco[1]), .B(idx_deco[0]), .Z(n_1511));
	notech_reg to_acu0_reg_143(.CP(n_62223), .D(n_38651), .CD(n_61675), .Q(to_acu0
		[143]));
	notech_mux2 i_46946(.S(n_55647), .A(to_acu0[143]), .B(n_40570), .Z(n_38651
		));
	notech_and2 i_275773(.A(n_1952), .B(n_39062), .Z(n_1510));
	notech_reg to_acu0_reg_144(.CP(n_62223), .D(n_38657), .CD(n_61675), .Q(to_acu0
		[144]));
	notech_mux2 i_46954(.S(n_55661), .A(to_acu0[144]), .B(n_40571), .Z(n_38657
		));
	notech_reg to_acu0_reg_145(.CP(n_62223), .D(n_38663), .CD(n_61675), .Q(to_acu0
		[145]));
	notech_mux2 i_46962(.S(n_55675), .A(to_acu0[145]), .B(n_39101), .Z(n_38663
		));
	notech_reg to_acu0_reg_146(.CP(n_62223), .D(n_38669), .CD(n_61675), .Q(to_acu0
		[146]));
	notech_mux2 i_46970(.S(n_55675), .A(to_acu0[146]), .B(n_39102), .Z(n_38669
		));
	notech_ao3 i_475771(.A(n_2219), .B(n_40501), .C(ipg_fault), .Z(n_1507)
		);
	notech_reg to_acu0_reg_147(.CP(n_62228), .D(n_38675), .CD(n_61675), .Q(to_acu0
		[147]));
	notech_mux2 i_46978(.S(n_55675), .A(to_acu0[147]), .B(n_39103), .Z(n_38675
		));
	notech_or4 i_122474572(.A(n_17551047), .B(in128[1]), .C(n_40916), .D(n_40839
		), .Z(n_1506));
	notech_reg to_acu0_reg_148(.CP(n_62228), .D(n_38681), .CD(n_61677), .Q(to_acu0
		[148]));
	notech_mux2 i_46986(.S(n_55675), .A(to_acu0[148]), .B(n_40572), .Z(n_38681
		));
	notech_or4 i_122374573(.A(idx_deco[1]), .B(n_59082), .C(idx_deco[0]), .D
		(n_223996470), .Z(n_1505));
	notech_reg to_acu0_reg_149(.CP(n_62225), .D(n_38687), .CD(n_61677), .Q(to_acu0
		[149]));
	notech_mux2 i_46994(.S(n_55675), .A(to_acu0[149]), .B(n_40573), .Z(n_38687
		));
	notech_or4 i_36475430(.A(i_ptr[1]), .B(i_ptr[0]), .C(i_ptr[3]), .D(i_ptr
		[2]), .Z(n_1504));
	notech_reg to_acu0_reg_150(.CP(n_62225), .D(n_38693), .CD(n_61677), .Q(to_acu0
		[150]));
	notech_mux2 i_47002(.S(n_55675), .A(to_acu0[150]), .B(n_39104), .Z(n_38693
		));
	notech_reg to_acu0_reg_151(.CP(n_62225), .D(n_38699), .CD(n_61677), .Q(to_acu0
		[151]));
	notech_mux2 i_47010(.S(n_55675), .A(to_acu0[151]), .B(n_39313), .Z(n_38699
		));
	notech_reg to_acu0_reg_152(.CP(n_62228), .D(n_38705), .CD(n_61677), .Q(to_acu0
		[152]));
	notech_mux2 i_47018(.S(n_55675), .A(to_acu0[152]), .B(n_39105), .Z(n_38705
		));
	notech_reg to_acu0_reg_153(.CP(n_62228), .D(n_38711), .CD(n_61680), .Q(to_acu0
		[153]));
	notech_mux2 i_47026(.S(n_55675), .A(to_acu0[153]), .B(n_39106), .Z(n_38711
		));
	notech_reg to_acu0_reg_154(.CP(n_62228), .D(n_38717), .CD(n_61680), .Q(to_acu0
		[154]));
	notech_mux2 i_47034(.S(n_55675), .A(to_acu0[154]), .B(n_40574), .Z(n_38717
		));
	notech_reg to_acu0_reg_155(.CP(n_62228), .D(n_38723), .CD(n_61680), .Q(to_acu0
		[155]));
	notech_mux2 i_47042(.S(n_55671), .A(to_acu0[155]), .B(n_40575), .Z(n_38723
		));
	notech_reg to_acu0_reg_156(.CP(n_62228), .D(n_38729), .CD(n_61680), .Q(to_acu0
		[156]));
	notech_mux2 i_47050(.S(n_55675), .A(to_acu0[156]), .B(n_39316), .Z(n_38729
		));
	notech_reg to_acu0_reg_157(.CP(n_62225), .D(n_38735), .CD(n_61680), .Q(to_acu0
		[157]));
	notech_mux2 i_47058(.S(n_55675), .A(to_acu0[157]), .B(n_40576), .Z(n_38735
		));
	notech_reg to_acu0_reg_158(.CP(n_62225), .D(n_38741), .CD(n_61677), .Q(to_acu0
		[158]));
	notech_mux2 i_47066(.S(n_55675), .A(to_acu0[158]), .B(n_39319), .Z(n_38741
		));
	notech_reg to_acu0_reg_159(.CP(n_62225), .D(n_38747), .CD(n_61677), .Q(to_acu0
		[159]));
	notech_mux2 i_47074(.S(n_55675), .A(to_acu0[159]), .B(n_40577), .Z(n_38747
		));
	notech_reg to_acu0_reg_160(.CP(n_62225), .D(n_38753), .CD(n_61677), .Q(to_acu0
		[160]));
	notech_mux2 i_47082(.S(n_55675), .A(to_acu0[160]), .B(n_40578), .Z(n_38753
		));
	notech_reg to_acu0_reg_161(.CP(n_62225), .D(n_38759), .CD(n_61677), .Q(to_acu0
		[161]));
	notech_mux2 i_47090(.S(n_55680), .A(to_acu0[161]), .B(n_40579), .Z(n_38759
		));
	notech_reg to_acu0_reg_162(.CP(n_62225), .D(n_38765), .CD(n_61677), .Q(to_acu0
		[162]));
	notech_mux2 i_47098(.S(n_55680), .A(to_acu0[162]), .B(n_39107), .Z(n_38765
		));
	notech_reg to_acu0_reg_163(.CP(n_62225), .D(n_38771), .CD(n_61677), .Q(to_acu0
		[163]));
	notech_mux2 i_47106(.S(n_55680), .A(to_acu0[163]), .B(n_39320), .Z(n_38771
		));
	notech_reg to_acu0_reg_164(.CP(n_62225), .D(n_38777), .CD(n_61677), .Q(to_acu0
		[164]));
	notech_mux2 i_47114(.S(n_55680), .A(to_acu0[164]), .B(n_39323), .Z(n_38777
		));
	notech_reg to_acu0_reg_165(.CP(n_62225), .D(n_38783), .CD(n_61677), .Q(to_acu0
		[165]));
	notech_mux2 i_47122(.S(n_55680), .A(to_acu0[165]), .B(n_39324), .Z(n_38783
		));
	notech_reg to_acu0_reg_166(.CP(n_62225), .D(n_38789), .CD(n_61677), .Q(to_acu0
		[166]));
	notech_mux2 i_47130(.S(n_55684), .A(to_acu0[166]), .B(n_39325), .Z(n_38789
		));
	notech_reg to_acu0_reg_167(.CP(n_62225), .D(n_38795), .CD(n_61677), .Q(to_acu0
		[167]));
	notech_mux2 i_47138(.S(n_55684), .A(to_acu0[167]), .B(n_39326), .Z(n_38795
		));
	notech_reg to_acu0_reg_168(.CP(n_62223), .D(n_38801), .CD(n_61677), .Q(to_acu0
		[168]));
	notech_mux2 i_47146(.S(n_55680), .A(to_acu0[168]), .B(n_40580), .Z(n_38801
		));
	notech_reg to_acu0_reg_169(.CP(n_62218), .D(n_38807), .CD(n_61670), .Q(to_acu0
		[169]));
	notech_mux2 i_47154(.S(n_55680), .A(to_acu0[169]), .B(n_39327), .Z(n_38807
		));
	notech_reg to_acu0_reg_170(.CP(n_62218), .D(n_38813), .CD(n_61670), .Q(to_acu0
		[170]));
	notech_mux2 i_47162(.S(n_55680), .A(to_acu0[170]), .B(n_39328), .Z(n_38813
		));
	notech_reg to_acu0_reg_171(.CP(n_62218), .D(n_38819), .CD(n_61670), .Q(to_acu0
		[171]));
	notech_mux2 i_47170(.S(n_55680), .A(to_acu0[171]), .B(n_39329), .Z(n_38819
		));
	notech_reg to_acu0_reg_172(.CP(n_62218), .D(n_38825), .CD(n_61670), .Q(to_acu0
		[172]));
	notech_mux2 i_47178(.S(n_55680), .A(to_acu0[172]), .B(n_39108), .Z(n_38825
		));
	notech_reg to_acu0_reg_173(.CP(n_62218), .D(n_38831), .CD(n_61670), .Q(to_acu0
		[173]));
	notech_mux2 i_47186(.S(n_55680), .A(to_acu0[173]), .B(n_39330), .Z(n_38831
		));
	notech_reg to_acu0_reg_174(.CP(n_62218), .D(n_38837), .CD(n_61670), .Q(to_acu0
		[174]));
	notech_mux2 i_47194(.S(n_55680), .A(to_acu0[174]), .B(n_39331), .Z(n_38837
		));
	notech_reg to_acu0_reg_175(.CP(n_62218), .D(n_38843), .CD(n_61670), .Q(to_acu0
		[175]));
	notech_mux2 i_47202(.S(n_55680), .A(to_acu0[175]), .B(n_39332), .Z(n_38843
		));
	notech_reg to_acu0_reg_176(.CP(n_62218), .D(n_38849), .CD(n_61670), .Q(to_acu0
		[176]));
	notech_mux2 i_47210(.S(n_55680), .A(to_acu0[176]), .B(n_39109), .Z(n_38849
		));
	notech_reg to_acu0_reg_177(.CP(n_62218), .D(n_38855), .CD(n_61670), .Q(to_acu0
		[177]));
	notech_mux2 i_47218(.S(n_55680), .A(to_acu0[177]), .B(n_39333), .Z(n_38855
		));
	notech_reg to_acu0_reg_178(.CP(n_62218), .D(n_38861), .CD(n_61670), .Q(to_acu0
		[178]));
	notech_mux2 i_47226(.S(n_55641), .A(to_acu0[178]), .B(n_39334), .Z(n_38861
		));
	notech_reg to_acu0_reg_179(.CP(n_62218), .D(n_38867), .CD(n_61670), .Q(to_acu0
		[179]));
	notech_mux2 i_47234(.S(n_55641), .A(to_acu0[179]), .B(n_39335), .Z(n_38867
		));
	notech_reg to_acu0_reg_180(.CP(n_62213), .D(n_38873), .CD(n_61665), .Q(to_acu0
		[180]));
	notech_mux2 i_47242(.S(n_55641), .A(to_acu0[180]), .B(n_39336), .Z(n_38873
		));
	notech_reg to_acu0_reg_181(.CP(n_62213), .D(n_38879), .CD(n_61665), .Q(to_acu0
		[181]));
	notech_mux2 i_47250(.S(n_55641), .A(to_acu0[181]), .B(n_39337), .Z(n_38879
		));
	notech_reg to_acu0_reg_182(.CP(n_62213), .D(n_38885), .CD(n_61665), .Q(to_acu0
		[182]));
	notech_mux2 i_47258(.S(n_55641), .A(to_acu0[182]), .B(n_39338), .Z(n_38885
		));
	notech_reg to_acu0_reg_183(.CP(n_62213), .D(n_38891), .CD(n_61665), .Q(to_acu0
		[183]));
	notech_mux2 i_47266(.S(n_55641), .A(to_acu0[183]), .B(n_39340), .Z(n_38891
		));
	notech_reg to_acu0_reg_184(.CP(n_62213), .D(n_38897), .CD(n_61665), .Q(to_acu0
		[184]));
	notech_mux2 i_47274(.S(n_55641), .A(to_acu0[184]), .B(n_39343), .Z(n_38897
		));
	notech_reg to_acu0_reg_185(.CP(n_62218), .D(n_38903), .CD(n_61670), .Q(to_acu0
		[185]));
	notech_mux2 i_47282(.S(n_55641), .A(to_acu0[185]), .B(n_39346), .Z(n_38903
		));
	notech_reg to_acu0_reg_186(.CP(n_62218), .D(n_38909), .CD(n_61670), .Q(to_acu0
		[186]));
	notech_mux2 i_47290(.S(n_55661), .A(to_acu0[186]), .B(n_39349), .Z(n_38909
		));
	notech_reg to_acu0_reg_187(.CP(n_62218), .D(n_38915), .CD(n_61670), .Q(to_acu0
		[187]));
	notech_mux2 i_47298(.S(n_55661), .A(to_acu0[187]), .B(n_39351), .Z(n_38915
		));
	notech_reg to_acu0_reg_188(.CP(n_62213), .D(n_38921), .CD(n_61665), .Q(to_acu0
		[188]));
	notech_mux2 i_47306(.S(n_55661), .A(to_acu0[188]), .B(n_39352), .Z(n_38921
		));
	notech_reg to_acu0_reg_189(.CP(n_62218), .D(n_38927), .CD(n_61665), .Q(to_acu0
		[189]));
	notech_mux2 i_47314(.S(n_55661), .A(to_acu0[189]), .B(n_39353), .Z(n_38927
		));
	notech_reg to_acu0_reg_190(.CP(n_62220), .D(n_38933), .CD(n_61672), .Q(to_acu0
		[190]));
	notech_mux2 i_47322(.S(n_55641), .A(to_acu0[190]), .B(n_39354), .Z(n_38933
		));
	notech_reg to_acu0_reg_191(.CP(n_62220), .D(n_38939), .CD(n_61672), .Q(to_acu0
		[191]));
	notech_mux2 i_47330(.S(n_55641), .A(to_acu0[191]), .B(n_39355), .Z(n_38939
		));
	notech_reg to_acu0_reg_192(.CP(n_62220), .D(n_38945), .CD(n_61672), .Q(to_acu0
		[192]));
	notech_mux2 i_47338(.S(n_55641), .A(to_acu0[192]), .B(n_39356), .Z(n_38945
		));
	notech_reg to_acu0_reg_193(.CP(n_62220), .D(n_38951), .CD(n_61672), .Q(to_acu0
		[193]));
	notech_mux2 i_47346(.S(n_55641), .A(to_acu0[193]), .B(n_39357), .Z(n_38951
		));
	notech_reg to_acu0_reg_194(.CP(n_62220), .D(n_38957), .CD(n_61672), .Q(to_acu0
		[194]));
	notech_mux2 i_47354(.S(n_55641), .A(to_acu0[194]), .B(n_39358), .Z(n_38957
		));
	notech_reg to_acu0_reg_195(.CP(n_62220), .D(n_38963), .CD(n_61672), .Q(to_acu0
		[195]));
	notech_mux2 i_47362(.S(n_55671), .A(to_acu0[195]), .B(n_39110), .Z(n_38963
		));
	notech_reg to_acu0_reg_196(.CP(n_62220), .D(n_38969), .CD(n_61672), .Q(to_acu0
		[196]));
	notech_mux2 i_47370(.S(n_55671), .A(to_acu0[196]), .B(n_39359), .Z(n_38969
		));
	notech_reg to_acu0_reg_197(.CP(n_62220), .D(n_38975), .CD(n_61672), .Q(to_acu0
		[197]));
	notech_mux2 i_47378(.S(n_55671), .A(to_acu0[197]), .B(n_39360), .Z(n_38975
		));
	notech_reg to_acu0_reg_198(.CP(n_62220), .D(n_38981), .CD(n_61672), .Q(to_acu0
		[198]));
	notech_mux2 i_47386(.S(n_55671), .A(to_acu0[198]), .B(n_39362), .Z(n_38981
		));
	notech_reg to_acu0_reg_199(.CP(n_62220), .D(n_38987), .CD(n_61672), .Q(to_acu0
		[199]));
	notech_mux2 i_47394(.S(n_55671), .A(to_acu0[199]), .B(n_40581), .Z(n_38987
		));
	notech_reg to_acu0_reg_200(.CP(n_62220), .D(n_38993), .CD(n_61672), .Q(to_acu0
		[200]));
	notech_mux2 i_47402(.S(n_55671), .A(to_acu0[200]), .B(n_39364), .Z(n_38993
		));
	notech_reg to_acu0_reg_201(.CP(n_62220), .D(n_38999), .CD(n_61670), .Q(to_acu0
		[201]));
	notech_mux2 i_47410(.S(n_55671), .A(to_acu0[201]), .B(n_40582), .Z(n_38999
		));
	notech_reg to_acu0_reg_202(.CP(n_62220), .D(n_39005), .CD(n_61672), .Q(to_acu0
		[202]));
	notech_mux2 i_47418(.S(n_55671), .A(to_acu0[202]), .B(n_40583), .Z(n_39005
		));
	notech_reg to_acu0_reg_203(.CP(n_62218), .D(n_39011), .CD(n_61670), .Q(to_acu0
		[203]));
	notech_mux2 i_47426(.S(n_55671), .A(to_acu0[203]), .B(n_40584), .Z(n_39011
		));
	notech_reg to_acu0_reg_204(.CP(n_62218), .D(n_39017), .CD(n_61670), .Q(to_acu0
		[204]));
	notech_mux2 i_47434(.S(n_55671), .A(to_acu0[204]), .B(n_40585), .Z(n_39017
		));
	notech_reg to_acu0_reg_205(.CP(n_62218), .D(n_39023), .CD(n_61670), .Q(to_acu0
		[205]));
	notech_mux2 i_47442(.S(n_55641), .A(to_acu0[205]), .B(n_39365), .Z(n_39023
		));
	notech_nao3 i_28375511(.A(cpl[0]), .B(cpl[1]), .C(n_59037), .Z(n_1448)
		);
	notech_reg to_acu0_reg_206(.CP(n_62220), .D(n_39029), .CD(n_61672), .Q(to_acu0
		[206]));
	notech_mux2 i_47450(.S(n_55641), .A(to_acu0[206]), .B(n_40586), .Z(n_39029
		));
	notech_reg to_acu0_reg_207(.CP(n_62220), .D(n_39035), .CD(n_61672), .Q(to_acu0
		[207]));
	notech_mux2 i_47458(.S(n_55671), .A(to_acu0[207]), .B(n_39366), .Z(n_39035
		));
	notech_reg to_acu0_reg_208(.CP(n_62220), .D(n_39041), .CD(n_61672), .Q(to_acu0
		[208]));
	notech_mux2 i_47466(.S(n_55671), .A(to_acu0[208]), .B(n_40587), .Z(n_39041
		));
	notech_nand3 i_075775(.A(n_18051052), .B(n_1591), .C(n_1521), .Z(n_1445)
		);
	notech_reg to_acu0_reg_209(.CP(n_62220), .D(n_39047), .CD(n_61672), .Q(to_acu0
		[209]));
	notech_mux2 i_47474(.S(n_55671), .A(to_acu0[209]), .B(n_40588), .Z(n_39047
		));
	notech_reg to_acu0_reg_210(.CP(n_62220), .D(n_39053), .CD(n_61672), .Q(to_acu0
		[210]));
	notech_mux2 i_47482(.S(n_55671), .A(to_acu0[210]), .B(n_40590), .Z(n_39053
		));
	notech_inv i_52668(.A(n_163996334), .Z(n_39059));
	notech_inv i_52669(.A(n_169996394), .Z(n_39060));
	notech_inv i_52670(.A(n_170196396), .Z(n_39061));
	notech_inv i_52671(.A(n_5414), .Z(n_39062));
	notech_inv i_52672(.A(n_14051012), .Z(n_39063));
	notech_inv i_52674(.A(n_1768), .Z(n_39065));
	notech_inv i_52675(.A(n_2836), .Z(n_39066));
	notech_inv i_52676(.A(n_2834), .Z(n_39067));
	notech_inv i_52677(.A(n_2832), .Z(n_39068));
	notech_inv i_52678(.A(n_2830), .Z(n_39069));
	notech_inv i_52679(.A(n_2828), .Z(n_39070));
	notech_inv i_52680(.A(n_2826), .Z(n_39071));
	notech_inv i_52681(.A(n_2824), .Z(n_39072));
	notech_inv i_52682(.A(n_2822), .Z(n_39073));
	notech_inv i_52683(.A(n_2820), .Z(n_39074));
	notech_inv i_52684(.A(n_2818), .Z(n_39075));
	notech_inv i_52685(.A(n_2816), .Z(n_39076));
	notech_inv i_52686(.A(n_2814), .Z(n_39077));
	notech_inv i_52687(.A(n_2812), .Z(n_39078));
	notech_inv i_52688(.A(n_2810), .Z(n_39079));
	notech_inv i_52689(.A(n_2808), .Z(n_39080));
	notech_inv i_52690(.A(n_2806), .Z(n_39081));
	notech_inv i_52691(.A(n_2804), .Z(n_39082));
	notech_inv i_52692(.A(n_2802), .Z(n_39083));
	notech_inv i_52693(.A(n_2800), .Z(n_39084));
	notech_inv i_52694(.A(n_2798), .Z(n_39085));
	notech_inv i_52695(.A(n_2796), .Z(n_39086));
	notech_inv i_52696(.A(n_2794), .Z(n_39087));
	notech_inv i_52697(.A(n_2792), .Z(n_39088));
	notech_inv i_52698(.A(n_2790), .Z(n_39089));
	notech_inv i_52699(.A(n_2788), .Z(n_39090));
	notech_inv i_52700(.A(n_2786), .Z(n_39091));
	notech_inv i_52701(.A(n_2784), .Z(n_39092));
	notech_inv i_52702(.A(n_2782), .Z(n_39093));
	notech_inv i_52703(.A(n_2780), .Z(n_39094));
	notech_inv i_52704(.A(n_2778), .Z(n_39095));
	notech_inv i_52705(.A(n_2776), .Z(n_39096));
	notech_inv i_52706(.A(n_2774), .Z(n_39097));
	notech_inv i_52707(.A(n_2772), .Z(n_39098));
	notech_inv i_52708(.A(n_2770), .Z(n_39099));
	notech_inv i_52709(.A(n_2768), .Z(n_39100));
	notech_inv i_52710(.A(n_2766), .Z(n_39101));
	notech_inv i_52711(.A(n_2764), .Z(n_39102));
	notech_inv i_52712(.A(n_2762), .Z(n_39103));
	notech_inv i_52713(.A(n_2760), .Z(n_39104));
	notech_inv i_52714(.A(n_2758), .Z(n_39105));
	notech_inv i_52715(.A(n_2756), .Z(n_39106));
	notech_inv i_52716(.A(n_2754), .Z(n_39107));
	notech_inv i_52717(.A(n_2752), .Z(n_39108));
	notech_inv i_52718(.A(n_275094707), .Z(n_39109));
	notech_inv i_52719(.A(n_274894705), .Z(n_39110));
	notech_inv i_52720(.A(n_274694703), .Z(n_39111));
	notech_inv i_52721(.A(n_273194688), .Z(n_39112));
	notech_inv i_52722(.A(n_272994686), .Z(n_39113));
	notech_inv i_52723(.A(n_272794684), .Z(n_39114));
	notech_inv i_52724(.A(n_272594682), .Z(n_39115));
	notech_inv i_52725(.A(n_272394680), .Z(n_39116));
	notech_inv i_52726(.A(n_272194678), .Z(n_39117));
	notech_inv i_52727(.A(n_271994676), .Z(n_39118));
	notech_inv i_52728(.A(n_271794674), .Z(n_39119));
	notech_inv i_52729(.A(n_271094667), .Z(n_39120));
	notech_inv i_52730(.A(n_270494661), .Z(n_39121));
	notech_inv i_52731(.A(n_269494651), .Z(n_39122));
	notech_inv i_52732(.A(n_268094637), .Z(n_39123));
	notech_inv i_52733(.A(n_267894635), .Z(n_39124));
	notech_inv i_52734(.A(n_267694633), .Z(n_39125));
	notech_inv i_52735(.A(n_267494631), .Z(n_39126));
	notech_inv i_52736(.A(n_267294629), .Z(n_39127));
	notech_inv i_52737(.A(n_146096155), .Z(n_39128));
	notech_inv i_52738(.A(n_267094627), .Z(n_39129));
	notech_inv i_52739(.A(n_266894625), .Z(n_39130));
	notech_inv i_52740(.A(n_172396417), .Z(n_39131));
	notech_inv i_52741(.A(n_266694623), .Z(n_39132));
	notech_inv i_52742(.A(n_227296437), .Z(n_39133));
	notech_inv i_52743(.A(n_266494621), .Z(n_39134));
	notech_inv i_52744(.A(n_2027), .Z(start));
	notech_inv i_52745(.A(n_266294619), .Z(n_39136));
	notech_inv i_52746(.A(n_266094617), .Z(n_39137));
	notech_inv i_52747(.A(n_265894615), .Z(n_39138));
	notech_inv i_52748(.A(term_f), .Z(n_39139));
	notech_inv i_52749(.A(n_265694613), .Z(n_39140));
	notech_inv i_52750(.A(n_265494611), .Z(n_39141));
	notech_inv i_52751(.A(n_265294609), .Z(n_39142));
	notech_inv i_52752(.A(\fpu_indrm[0] ), .Z(n_39143));
	notech_inv i_52753(.A(n_265094607), .Z(n_39144));
	notech_inv i_52754(.A(n_264894605), .Z(n_39145));
	notech_inv i_52755(.A(n_264694603), .Z(n_39146));
	notech_inv i_52756(.A(n_264494601), .Z(n_39147));
	notech_inv i_52757(.A(\fpu_indrm[3] ), .Z(n_39148));
	notech_inv i_52758(.A(n_264294599), .Z(n_39149));
	notech_inv i_52759(.A(n_264094597), .Z(n_39150));
	notech_inv i_52760(.A(n_263894595), .Z(n_39151));
	notech_inv i_52761(.A(n_263694593), .Z(n_39152));
	notech_inv i_52762(.A(n_263494591), .Z(n_39153));
	notech_inv i_52763(.A(n_263294589), .Z(n_39154));
	notech_inv i_52764(.A(n_263094587), .Z(n_39155));
	notech_inv i_52765(.A(n_262894585), .Z(n_39156));
	notech_inv i_52766(.A(n_262694583), .Z(n_39157));
	notech_inv i_52767(.A(n_262494581), .Z(n_39158));
	notech_inv i_52768(.A(n_262294579), .Z(n_39159));
	notech_inv i_52769(.A(n_262094577), .Z(n_39160));
	notech_inv i_52770(.A(n_261894575), .Z(n_39161));
	notech_inv i_52771(.A(n_261394570), .Z(n_39162));
	notech_inv i_52772(.A(n_261194568), .Z(n_39163));
	notech_inv i_52773(.A(n_260994566), .Z(n_39164));
	notech_inv i_52774(.A(n_260794564), .Z(n_39165));
	notech_inv i_52775(.A(n_260594562), .Z(n_39166));
	notech_inv i_52776(.A(n_260394560), .Z(n_39167));
	notech_inv i_52777(.A(n_260194558), .Z(n_39168));
	notech_inv i_52778(.A(n_259994556), .Z(n_39169));
	notech_inv i_52779(.A(n_259494551), .Z(n_39170));
	notech_inv i_52780(.A(n_259294549), .Z(n_39171));
	notech_inv i_52781(.A(\imm1[0] ), .Z(n_39172));
	notech_inv i_52782(.A(n_259094547), .Z(n_39173));
	notech_inv i_52783(.A(\imm1[1] ), .Z(n_39174));
	notech_inv i_52784(.A(\imm1[2] ), .Z(n_39175));
	notech_inv i_52785(.A(\imm1[3] ), .Z(n_39176));
	notech_inv i_52786(.A(\imm1[4] ), .Z(n_39177));
	notech_inv i_52787(.A(\imm1[5] ), .Z(n_39178));
	notech_inv i_52788(.A(\imm1[6] ), .Z(n_39179));
	notech_inv i_52789(.A(\imm1[7] ), .Z(n_39180));
	notech_inv i_52790(.A(\imm1[8] ), .Z(n_39181));
	notech_inv i_52791(.A(\imm1[9] ), .Z(n_39182));
	notech_inv i_52792(.A(\imm1[10] ), .Z(n_39183));
	notech_inv i_52793(.A(\imm1[11] ), .Z(n_39184));
	notech_inv i_52794(.A(\imm1[12] ), .Z(n_39185));
	notech_inv i_52795(.A(\imm1[13] ), .Z(n_39186));
	notech_inv i_52796(.A(\imm1[14] ), .Z(n_39187));
	notech_inv i_52797(.A(\imm1[15] ), .Z(n_39188));
	notech_inv i_52798(.A(\imm1[16] ), .Z(n_39189));
	notech_inv i_52799(.A(\imm1[17] ), .Z(n_39190));
	notech_inv i_52800(.A(\imm1[18] ), .Z(n_39191));
	notech_inv i_52801(.A(\imm1[19] ), .Z(n_39192));
	notech_inv i_52802(.A(\imm1[20] ), .Z(n_39193));
	notech_inv i_52803(.A(\imm1[21] ), .Z(n_39194));
	notech_inv i_52804(.A(n_223596474), .Z(n_39195));
	notech_inv i_52805(.A(\imm1[22] ), .Z(n_39196));
	notech_inv i_52806(.A(n_3819), .Z(n_39197));
	notech_inv i_52807(.A(\imm1[23] ), .Z(n_39198));
	notech_inv i_52808(.A(n_3818), .Z(n_39199));
	notech_inv i_52809(.A(\imm1[24] ), .Z(n_39200));
	notech_inv i_52810(.A(n_3817), .Z(n_39201));
	notech_inv i_52811(.A(\imm1[25] ), .Z(n_39202));
	notech_inv i_52812(.A(n_3816), .Z(n_39203));
	notech_inv i_52813(.A(\imm1[26] ), .Z(n_39204));
	notech_inv i_52814(.A(n_3815), .Z(n_39205));
	notech_inv i_52815(.A(\imm1[27] ), .Z(n_39206));
	notech_inv i_52816(.A(n_3814), .Z(n_39207));
	notech_inv i_52817(.A(\imm1[28] ), .Z(n_39208));
	notech_inv i_52818(.A(n_3813), .Z(n_39209));
	notech_inv i_52819(.A(\imm1[29] ), .Z(n_39210));
	notech_inv i_52820(.A(n_3812), .Z(n_39211));
	notech_inv i_52821(.A(\imm1[30] ), .Z(n_39212));
	notech_inv i_52822(.A(n_3811), .Z(n_39213));
	notech_inv i_52823(.A(\imm1[31] ), .Z(n_39214));
	notech_inv i_52824(.A(n_3810), .Z(n_39215));
	notech_inv i_52825(.A(\imm1[32] ), .Z(n_39216));
	notech_inv i_52826(.A(n_3809), .Z(n_39217));
	notech_inv i_52827(.A(\imm1[33] ), .Z(n_39218));
	notech_inv i_52828(.A(n_3808), .Z(n_39219));
	notech_inv i_52829(.A(\imm1[34] ), .Z(n_39220));
	notech_inv i_52830(.A(n_3807), .Z(n_39221));
	notech_inv i_52831(.A(\imm1[35] ), .Z(n_39222));
	notech_inv i_52832(.A(n_3806), .Z(n_39223));
	notech_inv i_52833(.A(\imm1[36] ), .Z(n_39224));
	notech_inv i_52834(.A(n_3805), .Z(n_39225));
	notech_inv i_52835(.A(\imm1[37] ), .Z(n_39226));
	notech_inv i_52836(.A(n_3804), .Z(n_39227));
	notech_inv i_52837(.A(\imm1[38] ), .Z(n_39228));
	notech_inv i_52838(.A(n_3803), .Z(n_39229));
	notech_inv i_52839(.A(\imm1[39] ), .Z(n_39230));
	notech_inv i_52840(.A(n_3802), .Z(n_39231));
	notech_inv i_52841(.A(\imm1[40] ), .Z(n_39232));
	notech_inv i_52842(.A(n_3801), .Z(n_39233));
	notech_inv i_52843(.A(\imm1[41] ), .Z(n_39234));
	notech_inv i_52844(.A(n_3800), .Z(n_39235));
	notech_inv i_52845(.A(\imm1[42] ), .Z(n_39236));
	notech_inv i_52846(.A(n_3799), .Z(n_39237));
	notech_inv i_52847(.A(\imm1[43] ), .Z(n_39238));
	notech_inv i_52848(.A(n_3798), .Z(n_39239));
	notech_inv i_52849(.A(\imm1[44] ), .Z(n_39240));
	notech_inv i_52850(.A(n_3797), .Z(n_39241));
	notech_inv i_52851(.A(\imm1[45] ), .Z(n_39242));
	notech_inv i_52852(.A(n_3796), .Z(n_39243));
	notech_inv i_52853(.A(\imm1[46] ), .Z(n_39244));
	notech_inv i_52854(.A(n_3795), .Z(n_39245));
	notech_inv i_52855(.A(\imm1[47] ), .Z(n_39246));
	notech_inv i_52856(.A(n_3794), .Z(n_39247));
	notech_inv i_52857(.A(\imm2[0] ), .Z(n_39248));
	notech_inv i_52858(.A(\imm2[1] ), .Z(n_39249));
	notech_inv i_52859(.A(n_3793), .Z(n_39250));
	notech_inv i_52860(.A(\imm2[2] ), .Z(n_39251));
	notech_inv i_52861(.A(\imm2[3] ), .Z(n_39252));
	notech_inv i_52862(.A(n_3792), .Z(n_39253));
	notech_inv i_52863(.A(\imm2[4] ), .Z(n_39254));
	notech_inv i_52864(.A(\imm2[5] ), .Z(n_39255));
	notech_inv i_52865(.A(n_3791), .Z(n_39256));
	notech_inv i_52866(.A(\imm2[6] ), .Z(n_39257));
	notech_inv i_52867(.A(\imm2[7] ), .Z(n_39258));
	notech_inv i_52868(.A(n_3790), .Z(n_39259));
	notech_inv i_52869(.A(\imm2[8] ), .Z(n_39260));
	notech_inv i_52870(.A(\imm2[9] ), .Z(n_39261));
	notech_inv i_52871(.A(n_3789), .Z(n_39262));
	notech_inv i_52872(.A(\imm2[10] ), .Z(n_39263));
	notech_inv i_52873(.A(\imm2[11] ), .Z(n_39264));
	notech_inv i_52874(.A(n_3788), .Z(n_39265));
	notech_inv i_52875(.A(\imm2[12] ), .Z(n_39266));
	notech_inv i_52876(.A(\imm2[13] ), .Z(n_39267));
	notech_inv i_52877(.A(n_3787), .Z(n_39268));
	notech_inv i_52878(.A(\imm2[14] ), .Z(n_39269));
	notech_inv i_52879(.A(\imm2[15] ), .Z(n_39270));
	notech_inv i_52880(.A(n_3786), .Z(n_39271));
	notech_inv i_52881(.A(\imm2[16] ), .Z(n_39272));
	notech_inv i_52882(.A(\imm2[17] ), .Z(n_39273));
	notech_inv i_52883(.A(n_3785), .Z(n_39274));
	notech_inv i_52884(.A(\imm2[18] ), .Z(n_39275));
	notech_inv i_52885(.A(\imm2[19] ), .Z(n_39276));
	notech_inv i_52886(.A(n_3784), .Z(n_39277));
	notech_inv i_52887(.A(\imm2[20] ), .Z(n_39278));
	notech_inv i_52888(.A(\imm2[21] ), .Z(n_39279));
	notech_inv i_52889(.A(n_3783), .Z(n_39280));
	notech_inv i_52890(.A(\imm2[22] ), .Z(n_39281));
	notech_inv i_52891(.A(\imm2[23] ), .Z(n_39282));
	notech_inv i_52892(.A(n_3782), .Z(n_39283));
	notech_inv i_52893(.A(\imm2[24] ), .Z(n_39284));
	notech_inv i_52894(.A(\imm2[25] ), .Z(n_39285));
	notech_inv i_52895(.A(n_3781), .Z(n_39286));
	notech_inv i_52896(.A(\imm2[26] ), .Z(n_39287));
	notech_inv i_52897(.A(\imm2[27] ), .Z(n_39288));
	notech_inv i_52898(.A(n_3780), .Z(n_39289));
	notech_inv i_52899(.A(\imm2[28] ), .Z(n_39290));
	notech_inv i_52900(.A(\imm2[29] ), .Z(n_39291));
	notech_inv i_52901(.A(n_3779), .Z(n_39292));
	notech_inv i_52902(.A(\imm2[30] ), .Z(n_39293));
	notech_inv i_52903(.A(\imm2[31] ), .Z(n_39294));
	notech_inv i_52904(.A(n_3778), .Z(n_39295));
	notech_inv i_52905(.A(\imm2[32] ), .Z(n_39296));
	notech_inv i_52906(.A(\imm2[33] ), .Z(n_39297));
	notech_inv i_52907(.A(n_3777), .Z(n_39298));
	notech_inv i_52908(.A(\imm2[34] ), .Z(n_39299));
	notech_inv i_52909(.A(\imm2[35] ), .Z(n_39300));
	notech_inv i_52910(.A(n_3776), .Z(n_39301));
	notech_inv i_52911(.A(\imm2[36] ), .Z(n_39302));
	notech_inv i_52912(.A(\imm2[37] ), .Z(n_39303));
	notech_inv i_52913(.A(n_3775), .Z(n_39304));
	notech_inv i_52914(.A(\imm2[38] ), .Z(n_39305));
	notech_inv i_52915(.A(\imm2[39] ), .Z(n_39306));
	notech_inv i_52916(.A(n_3774), .Z(n_39307));
	notech_inv i_52917(.A(\imm2[40] ), .Z(n_39308));
	notech_inv i_52918(.A(\imm2[41] ), .Z(n_39309));
	notech_inv i_52919(.A(n_3773), .Z(n_39310));
	notech_inv i_52920(.A(\imm2[42] ), .Z(n_39311));
	notech_inv i_52921(.A(\imm2[43] ), .Z(n_39312));
	notech_inv i_52922(.A(n_3772), .Z(n_39313));
	notech_inv i_52923(.A(\imm2[44] ), .Z(n_39314));
	notech_inv i_52924(.A(\imm2[45] ), .Z(n_39315));
	notech_inv i_52925(.A(n_3771), .Z(n_39316));
	notech_inv i_52926(.A(\imm2[46] ), .Z(n_39317));
	notech_inv i_52927(.A(\imm2[47] ), .Z(n_39318));
	notech_inv i_52928(.A(n_3770), .Z(n_39319));
	notech_inv i_52929(.A(n_3769), .Z(n_39320));
	notech_inv i_52930(.A(trig_itf), .Z(n_39321));
	notech_inv i_52931(.A(intf), .Z(n_39322));
	notech_inv i_52932(.A(n_3768), .Z(n_39323));
	notech_inv i_52933(.A(n_3767), .Z(n_39324));
	notech_inv i_52934(.A(n_3766), .Z(n_39325));
	notech_inv i_52935(.A(n_3765), .Z(n_39326));
	notech_inv i_52936(.A(n_3764), .Z(n_39327));
	notech_inv i_52937(.A(n_3763), .Z(n_39328));
	notech_inv i_52938(.A(n_3762), .Z(n_39329));
	notech_inv i_52939(.A(n_3761), .Z(n_39330));
	notech_inv i_52940(.A(n_3760), .Z(n_39331));
	notech_inv i_52941(.A(n_3759), .Z(n_39332));
	notech_inv i_52942(.A(n_3758), .Z(n_39333));
	notech_inv i_52943(.A(n_3757), .Z(n_39334));
	notech_inv i_52944(.A(n_3756), .Z(n_39335));
	notech_inv i_52945(.A(n_3755), .Z(n_39336));
	notech_inv i_52946(.A(n_3754), .Z(n_39337));
	notech_inv i_52947(.A(n_3753), .Z(n_39338));
	notech_inv i_52948(.A(ififo_rvect1[0]), .Z(n_39339));
	notech_inv i_52949(.A(n_3752), .Z(n_39340));
	notech_inv i_52950(.A(ififo_rvect1[1]), .Z(n_39341));
	notech_inv i_52951(.A(ififo_rvect1[2]), .Z(n_39342));
	notech_inv i_52952(.A(n_3751), .Z(n_39343));
	notech_inv i_52953(.A(ififo_rvect1[3]), .Z(n_39344));
	notech_inv i_52954(.A(ififo_rvect1[4]), .Z(n_39345));
	notech_inv i_52955(.A(n_3750), .Z(n_39346));
	notech_inv i_52956(.A(ififo_rvect1[5]), .Z(n_39347));
	notech_inv i_52957(.A(ififo_rvect1[6]), .Z(n_39348));
	notech_inv i_52958(.A(n_3749), .Z(n_39349));
	notech_inv i_52959(.A(ififo_rvect1[7]), .Z(n_39350));
	notech_inv i_52960(.A(n_3748), .Z(n_39351));
	notech_inv i_52961(.A(n_3747), .Z(n_39352));
	notech_inv i_52962(.A(n_3746), .Z(n_39353));
	notech_inv i_52963(.A(n_3745), .Z(n_39354));
	notech_inv i_52964(.A(n_3744), .Z(n_39355));
	notech_inv i_52965(.A(n_3743), .Z(n_39356));
	notech_inv i_52966(.A(n_3742), .Z(n_39357));
	notech_inv i_52967(.A(n_3741), .Z(n_39358));
	notech_inv i_52968(.A(n_3740), .Z(n_39359));
	notech_inv i_52969(.A(n_3739), .Z(n_39360));
	notech_inv i_52970(.A(n_44339), .Z(n_39361));
	notech_inv i_52971(.A(n_3738), .Z(n_39362));
	notech_inv i_52972(.A(n_49853), .Z(n_39363));
	notech_inv i_52973(.A(n_3737), .Z(n_39364));
	notech_inv i_52974(.A(n_3736), .Z(n_39365));
	notech_inv i_52975(.A(n_3735), .Z(n_39366));
	notech_inv i_52976(.A(n_3734), .Z(n_39367));
	notech_inv i_52977(.A(i_ptr[2]), .Z(n_39368));
	notech_inv i_52978(.A(n_3733), .Z(n_39369));
	notech_inv i_52979(.A(idx_deco[0]), .Z(n_39370));
	notech_inv i_52980(.A(n_3732), .Z(n_39371));
	notech_inv i_52981(.A(n_3731), .Z(n_39372));
	notech_inv i_52982(.A(n_3730), .Z(n_39373));
	notech_inv i_52983(.A(fsm[1]), .Z(n_39374));
	notech_inv i_52984(.A(n_3729), .Z(n_39375));
	notech_inv i_52985(.A(n_3728), .Z(n_39376));
	notech_inv i_52986(.A(fsm[4]), .Z(n_39377));
	notech_inv i_52987(.A(n_3727), .Z(n_39378));
	notech_inv i_52988(.A(n_3725), .Z(n_39379));
	notech_inv i_52989(.A(repz), .Z(n_39380));
	notech_inv i_52990(.A(rep), .Z(n_39381));
	notech_inv i_52991(.A(n_3723), .Z(n_39382));
	notech_inv i_52992(.A(n_3721), .Z(n_39383));
	notech_inv i_52993(.A(n_43076), .Z(n_39384));
	notech_inv i_52994(.A(n_3719), .Z(n_39385));
	notech_inv i_52995(.A(n_3717), .Z(n_39386));
	notech_inv i_52996(.A(n_3715), .Z(n_39387));
	notech_inv i_52997(.A(lenpc2[0]), .Z(n_39388));
	notech_inv i_52998(.A(n_3713), .Z(n_39389));
	notech_inv i_52999(.A(lenpc2[1]), .Z(n_39390));
	notech_inv i_53000(.A(lenpc2[2]), .Z(n_39391));
	notech_inv i_53001(.A(n_3711), .Z(n_39392));
	notech_inv i_53002(.A(lenpc2[3]), .Z(n_39393));
	notech_inv i_53003(.A(lenpc2[4]), .Z(n_39394));
	notech_inv i_53004(.A(n_3709), .Z(n_39395));
	notech_inv i_53005(.A(lenpc2[5]), .Z(n_39396));
	notech_inv i_53006(.A(n_3707), .Z(n_39397));
	notech_inv i_53007(.A(n_3705), .Z(n_39398));
	notech_inv i_53008(.A(n_3703), .Z(n_39399));
	notech_inv i_53009(.A(n_3701), .Z(n_39400));
	notech_inv i_53010(.A(n_3699), .Z(n_39401));
	notech_inv i_53011(.A(n_3697), .Z(n_39402));
	notech_inv i_53012(.A(n_3695), .Z(n_39403));
	notech_inv i_53013(.A(n_3693), .Z(n_39404));
	notech_inv i_53014(.A(n_3691), .Z(n_39405));
	notech_inv i_53015(.A(n_3689), .Z(n_39406));
	notech_inv i_53016(.A(n_3687), .Z(n_39407));
	notech_inv i_53017(.A(n_3685), .Z(n_39408));
	notech_inv i_53018(.A(n_3683), .Z(n_39409));
	notech_inv i_53019(.A(reps2[0]), .Z(n_39410));
	notech_inv i_53020(.A(n_3681), .Z(n_39411));
	notech_inv i_53021(.A(reps2[1]), .Z(n_39412));
	notech_inv i_53022(.A(reps2[2]), .Z(n_39413));
	notech_inv i_53023(.A(n_3679), .Z(n_39414));
	notech_inv i_53024(.A(reps1[0]), .Z(n_39415));
	notech_inv i_53025(.A(n_3677), .Z(n_39416));
	notech_inv i_53026(.A(n_50752), .Z(n_39417));
	notech_inv i_53027(.A(reps1[1]), .Z(n_39418));
	notech_inv i_53028(.A(n_50758), .Z(n_39419));
	notech_inv i_53029(.A(reps1[2]), .Z(n_39420));
	notech_inv i_53030(.A(n_3675), .Z(n_39421));
	notech_inv i_53031(.A(inst_deco2[0]), .Z(n_39422));
	notech_inv i_53032(.A(inst_deco2[1]), .Z(n_39423));
	notech_inv i_53033(.A(n_3673), .Z(n_39424));
	notech_inv i_53034(.A(inst_deco2[2]), .Z(n_39425));
	notech_inv i_53035(.A(inst_deco2[3]), .Z(n_39426));
	notech_inv i_53036(.A(n_3671), .Z(n_39427));
	notech_inv i_53037(.A(inst_deco2[4]), .Z(n_39428));
	notech_inv i_53038(.A(inst_deco2[5]), .Z(n_39429));
	notech_inv i_53039(.A(n_3669), .Z(n_39430));
	notech_inv i_53040(.A(inst_deco2[6]), .Z(n_39431));
	notech_inv i_53041(.A(inst_deco2[7]), .Z(n_39432));
	notech_inv i_53042(.A(n_3667), .Z(n_39433));
	notech_inv i_53043(.A(inst_deco2[8]), .Z(n_39434));
	notech_inv i_53044(.A(inst_deco2[9]), .Z(n_39435));
	notech_inv i_53045(.A(n_3665), .Z(n_39436));
	notech_inv i_53046(.A(inst_deco2[10]), .Z(n_39437));
	notech_inv i_53047(.A(inst_deco2[11]), .Z(n_39438));
	notech_inv i_53048(.A(n_3663), .Z(n_39439));
	notech_inv i_53049(.A(inst_deco2[12]), .Z(n_39440));
	notech_inv i_53050(.A(inst_deco2[13]), .Z(n_39441));
	notech_inv i_53051(.A(n_3661), .Z(n_39442));
	notech_inv i_53052(.A(inst_deco2[14]), .Z(n_39443));
	notech_inv i_53053(.A(inst_deco2[15]), .Z(n_39444));
	notech_inv i_53054(.A(n_3659), .Z(n_39445));
	notech_inv i_53055(.A(inst_deco2[16]), .Z(n_39446));
	notech_inv i_53056(.A(inst_deco2[17]), .Z(n_39447));
	notech_inv i_53057(.A(n_3657), .Z(n_39448));
	notech_inv i_53058(.A(inst_deco2[18]), .Z(n_39449));
	notech_inv i_53059(.A(inst_deco2[19]), .Z(n_39450));
	notech_inv i_53060(.A(n_3655), .Z(n_39451));
	notech_inv i_53061(.A(inst_deco2[20]), .Z(n_39452));
	notech_inv i_53062(.A(inst_deco2[21]), .Z(n_39453));
	notech_inv i_53063(.A(n_3653), .Z(n_39454));
	notech_inv i_53064(.A(inst_deco2[22]), .Z(n_39455));
	notech_inv i_53065(.A(inst_deco2[23]), .Z(n_39456));
	notech_inv i_53066(.A(n_3651), .Z(n_39457));
	notech_inv i_53067(.A(inst_deco2[24]), .Z(n_39458));
	notech_inv i_53068(.A(inst_deco2[25]), .Z(n_39459));
	notech_inv i_53069(.A(n_3649), .Z(n_39460));
	notech_inv i_53070(.A(inst_deco2[26]), .Z(n_39461));
	notech_inv i_53071(.A(inst_deco2[27]), .Z(n_39462));
	notech_inv i_53072(.A(n_3647), .Z(n_39463));
	notech_inv i_53073(.A(inst_deco2[28]), .Z(n_39464));
	notech_inv i_53074(.A(inst_deco2[29]), .Z(n_39465));
	notech_inv i_53075(.A(n_3645), .Z(n_39466));
	notech_inv i_53076(.A(inst_deco2[30]), .Z(n_39467));
	notech_inv i_53077(.A(inst_deco2[31]), .Z(n_39468));
	notech_inv i_53078(.A(n_3643), .Z(n_39469));
	notech_inv i_53079(.A(inst_deco2[32]), .Z(n_39470));
	notech_inv i_53080(.A(inst_deco2[33]), .Z(n_39471));
	notech_inv i_53081(.A(n_3641), .Z(n_39472));
	notech_inv i_53082(.A(inst_deco2[34]), .Z(n_39473));
	notech_inv i_53083(.A(inst_deco2[35]), .Z(n_39474));
	notech_inv i_53084(.A(n_3639), .Z(n_39475));
	notech_inv i_53085(.A(inst_deco2[36]), .Z(n_39476));
	notech_inv i_53086(.A(inst_deco2[37]), .Z(n_39477));
	notech_inv i_53087(.A(n_3637), .Z(n_39478));
	notech_inv i_53088(.A(inst_deco2[38]), .Z(n_39479));
	notech_inv i_53089(.A(inst_deco2[39]), .Z(n_39480));
	notech_inv i_53090(.A(n_3635), .Z(n_39481));
	notech_inv i_53091(.A(inst_deco2[40]), .Z(n_39482));
	notech_inv i_53092(.A(inst_deco2[41]), .Z(n_39483));
	notech_inv i_53093(.A(n_3634), .Z(n_39484));
	notech_inv i_53094(.A(inst_deco2[42]), .Z(n_39485));
	notech_inv i_53095(.A(inst_deco2[43]), .Z(n_39486));
	notech_inv i_53096(.A(n_3632), .Z(n_39487));
	notech_inv i_53097(.A(inst_deco2[44]), .Z(n_39488));
	notech_inv i_53098(.A(inst_deco2[45]), .Z(n_39489));
	notech_inv i_53099(.A(n_3630), .Z(n_39490));
	notech_inv i_53100(.A(inst_deco2[46]), .Z(n_39491));
	notech_inv i_53101(.A(inst_deco2[47]), .Z(n_39492));
	notech_inv i_53102(.A(n_3628), .Z(n_39493));
	notech_inv i_53103(.A(inst_deco2[48]), .Z(n_39494));
	notech_inv i_53104(.A(inst_deco2[49]), .Z(n_39495));
	notech_inv i_53105(.A(n_3626), .Z(n_39496));
	notech_inv i_53106(.A(inst_deco2[50]), .Z(n_39497));
	notech_inv i_53107(.A(inst_deco2[51]), .Z(n_39498));
	notech_inv i_53108(.A(n_3624), .Z(n_39499));
	notech_inv i_53109(.A(inst_deco2[52]), .Z(n_39500));
	notech_inv i_53110(.A(inst_deco2[53]), .Z(n_39501));
	notech_inv i_53111(.A(n_3622), .Z(n_39502));
	notech_inv i_53112(.A(inst_deco2[54]), .Z(n_39503));
	notech_inv i_53113(.A(inst_deco2[55]), .Z(n_39504));
	notech_inv i_53114(.A(n_3620), .Z(n_39505));
	notech_inv i_53115(.A(inst_deco2[56]), .Z(n_39506));
	notech_inv i_53116(.A(inst_deco2[57]), .Z(n_39507));
	notech_inv i_53117(.A(n_3618), .Z(n_39508));
	notech_inv i_53118(.A(inst_deco2[58]), .Z(n_39509));
	notech_inv i_53119(.A(inst_deco2[59]), .Z(n_39510));
	notech_inv i_53120(.A(n_3616), .Z(n_39511));
	notech_inv i_53121(.A(inst_deco2[60]), .Z(n_39512));
	notech_inv i_53122(.A(inst_deco2[61]), .Z(n_39513));
	notech_inv i_53123(.A(n_3614), .Z(n_39514));
	notech_inv i_53124(.A(inst_deco2[62]), .Z(n_39515));
	notech_inv i_53125(.A(inst_deco2[63]), .Z(n_39516));
	notech_inv i_53126(.A(n_3612), .Z(n_39517));
	notech_inv i_53127(.A(inst_deco2[64]), .Z(n_39518));
	notech_inv i_53128(.A(inst_deco2[65]), .Z(n_39519));
	notech_inv i_53129(.A(n_3610), .Z(n_39520));
	notech_inv i_53130(.A(inst_deco2[66]), .Z(n_39521));
	notech_inv i_53131(.A(inst_deco2[67]), .Z(n_39522));
	notech_inv i_53132(.A(n_3608), .Z(n_39523));
	notech_inv i_53133(.A(inst_deco2[68]), .Z(n_39524));
	notech_inv i_53134(.A(inst_deco2[69]), .Z(n_39525));
	notech_inv i_53135(.A(n_3606), .Z(n_39526));
	notech_inv i_53136(.A(inst_deco2[70]), .Z(n_39527));
	notech_inv i_53137(.A(inst_deco2[71]), .Z(n_39528));
	notech_inv i_53138(.A(n_3604), .Z(n_39529));
	notech_inv i_53139(.A(inst_deco2[72]), .Z(n_39530));
	notech_inv i_53140(.A(inst_deco2[73]), .Z(n_39531));
	notech_inv i_53141(.A(n_3602), .Z(n_39532));
	notech_inv i_53142(.A(inst_deco2[74]), .Z(n_39533));
	notech_inv i_53143(.A(inst_deco2[75]), .Z(n_39534));
	notech_inv i_53144(.A(n_3600), .Z(n_39535));
	notech_inv i_53145(.A(inst_deco2[76]), .Z(n_39536));
	notech_inv i_53146(.A(inst_deco2[77]), .Z(n_39537));
	notech_inv i_53147(.A(n_3598), .Z(n_39538));
	notech_inv i_53148(.A(inst_deco2[78]), .Z(n_39539));
	notech_inv i_53149(.A(inst_deco2[79]), .Z(n_39540));
	notech_inv i_53150(.A(n_3596), .Z(n_39541));
	notech_inv i_53151(.A(inst_deco2[80]), .Z(n_39542));
	notech_inv i_53152(.A(inst_deco2[81]), .Z(n_39543));
	notech_inv i_53153(.A(n_3594), .Z(n_39544));
	notech_inv i_53154(.A(inst_deco2[82]), .Z(n_39545));
	notech_inv i_53155(.A(inst_deco2[83]), .Z(n_39546));
	notech_inv i_53156(.A(n_3592), .Z(n_39547));
	notech_inv i_53157(.A(inst_deco2[84]), .Z(n_39548));
	notech_inv i_53158(.A(inst_deco2[85]), .Z(n_39549));
	notech_inv i_53159(.A(n_3590), .Z(n_39550));
	notech_inv i_53160(.A(inst_deco2[86]), .Z(n_39551));
	notech_inv i_53161(.A(inst_deco2[87]), .Z(n_39552));
	notech_inv i_53162(.A(n_3588), .Z(n_39553));
	notech_inv i_53163(.A(inst_deco2[88]), .Z(n_39554));
	notech_inv i_53164(.A(inst_deco2[89]), .Z(n_39555));
	notech_inv i_53165(.A(n_3586), .Z(n_39556));
	notech_inv i_53166(.A(inst_deco2[90]), .Z(n_39557));
	notech_inv i_53167(.A(inst_deco2[91]), .Z(n_39558));
	notech_inv i_53168(.A(n_3584), .Z(n_39559));
	notech_inv i_53169(.A(inst_deco2[92]), .Z(n_39560));
	notech_inv i_53170(.A(inst_deco2[93]), .Z(n_39561));
	notech_inv i_53171(.A(n_3582), .Z(n_39562));
	notech_inv i_53172(.A(inst_deco2[94]), .Z(n_39563));
	notech_inv i_53173(.A(inst_deco2[95]), .Z(n_39564));
	notech_inv i_53174(.A(n_3580), .Z(n_39565));
	notech_inv i_53175(.A(inst_deco2[96]), .Z(n_39566));
	notech_inv i_53176(.A(inst_deco2[97]), .Z(n_39567));
	notech_inv i_53177(.A(n_3578), .Z(n_39568));
	notech_inv i_53178(.A(inst_deco2[98]), .Z(n_39569));
	notech_inv i_53179(.A(inst_deco2[99]), .Z(n_39570));
	notech_inv i_53180(.A(n_3576), .Z(n_39571));
	notech_inv i_53181(.A(inst_deco2[100]), .Z(n_39572));
	notech_inv i_53182(.A(inst_deco2[101]), .Z(n_39573));
	notech_inv i_53183(.A(n_3574), .Z(n_39574));
	notech_inv i_53184(.A(inst_deco2[102]), .Z(n_39575));
	notech_inv i_53185(.A(n_43810), .Z(n_39576));
	notech_inv i_53186(.A(inst_deco2[103]), .Z(n_39577));
	notech_inv i_53187(.A(n_3573), .Z(n_39578));
	notech_inv i_53188(.A(inst_deco2[104]), .Z(n_39579));
	notech_inv i_53189(.A(inst_deco2[105]), .Z(n_39580));
	notech_inv i_53190(.A(n_3572), .Z(n_39581));
	notech_inv i_53191(.A(inst_deco2[106]), .Z(n_39582));
	notech_inv i_53192(.A(inst_deco2[107]), .Z(n_39583));
	notech_inv i_53193(.A(n_3571), .Z(n_39584));
	notech_inv i_53194(.A(inst_deco2[108]), .Z(n_39585));
	notech_inv i_53195(.A(inst_deco2[109]), .Z(n_39586));
	notech_inv i_53196(.A(n_3570), .Z(n_39587));
	notech_inv i_53197(.A(inst_deco2[110]), .Z(n_39588));
	notech_inv i_53198(.A(inst_deco2[111]), .Z(n_39589));
	notech_inv i_53199(.A(n_3569), .Z(n_39590));
	notech_inv i_53200(.A(inst_deco2[112]), .Z(n_39591));
	notech_inv i_53201(.A(inst_deco2[113]), .Z(n_39592));
	notech_inv i_53202(.A(n_3568), .Z(n_39593));
	notech_inv i_53203(.A(inst_deco2[114]), .Z(n_39594));
	notech_inv i_53204(.A(inst_deco2[115]), .Z(n_39595));
	notech_inv i_53205(.A(n_3567), .Z(n_39596));
	notech_inv i_53206(.A(inst_deco2[116]), .Z(n_39597));
	notech_inv i_53207(.A(inst_deco2[117]), .Z(n_39598));
	notech_inv i_53208(.A(n_3566), .Z(n_39599));
	notech_inv i_53209(.A(inst_deco2[118]), .Z(n_39600));
	notech_inv i_53210(.A(inst_deco2[119]), .Z(n_39601));
	notech_inv i_53211(.A(n_3565), .Z(n_39602));
	notech_inv i_53212(.A(inst_deco2[120]), .Z(n_39603));
	notech_inv i_53213(.A(inst_deco2[121]), .Z(n_39604));
	notech_inv i_53214(.A(n_3564), .Z(n_39605));
	notech_inv i_53215(.A(inst_deco2[122]), .Z(n_39606));
	notech_inv i_53216(.A(inst_deco2[123]), .Z(n_39607));
	notech_inv i_53217(.A(n_3563), .Z(n_39608));
	notech_inv i_53218(.A(inst_deco2[124]), .Z(n_39609));
	notech_inv i_53219(.A(inst_deco2[125]), .Z(n_39610));
	notech_inv i_53220(.A(n_3562), .Z(n_39611));
	notech_inv i_53221(.A(inst_deco2[126]), .Z(n_39612));
	notech_inv i_53222(.A(inst_deco2[127]), .Z(n_39613));
	notech_inv i_53223(.A(n_3561), .Z(n_39614));
	notech_inv i_53224(.A(inst_deco1[0]), .Z(n_39615));
	notech_inv i_53225(.A(n_3560), .Z(n_39616));
	notech_inv i_53226(.A(inst_deco1[1]), .Z(n_39617));
	notech_inv i_53227(.A(n_3559), .Z(n_39618));
	notech_inv i_53228(.A(inst_deco1[2]), .Z(n_39619));
	notech_inv i_53229(.A(n_3558), .Z(n_39620));
	notech_inv i_53230(.A(inst_deco1[3]), .Z(n_39621));
	notech_inv i_53231(.A(n_3557), .Z(n_39622));
	notech_inv i_53232(.A(inst_deco1[4]), .Z(n_39623));
	notech_inv i_53233(.A(n_3556), .Z(n_39624));
	notech_inv i_53234(.A(inst_deco1[5]), .Z(n_39625));
	notech_inv i_53235(.A(n_3555), .Z(n_39626));
	notech_inv i_53236(.A(inst_deco1[6]), .Z(n_39627));
	notech_inv i_53237(.A(n_3554), .Z(n_39628));
	notech_inv i_53238(.A(inst_deco1[7]), .Z(n_39629));
	notech_inv i_53239(.A(n_3553), .Z(n_39630));
	notech_inv i_53240(.A(inst_deco1[8]), .Z(n_39631));
	notech_inv i_53241(.A(n_3552), .Z(n_39632));
	notech_inv i_53242(.A(inst_deco1[9]), .Z(n_39633));
	notech_inv i_53243(.A(n_3551), .Z(n_39634));
	notech_inv i_53244(.A(inst_deco1[10]), .Z(n_39635));
	notech_inv i_53245(.A(n_3550), .Z(n_39636));
	notech_inv i_53246(.A(inst_deco1[11]), .Z(n_39637));
	notech_inv i_53247(.A(n_3549), .Z(n_39638));
	notech_inv i_53248(.A(inst_deco1[12]), .Z(n_39639));
	notech_inv i_53249(.A(n_3548), .Z(n_39640));
	notech_inv i_53250(.A(inst_deco1[13]), .Z(n_39641));
	notech_inv i_53251(.A(n_3547), .Z(n_39642));
	notech_inv i_53252(.A(inst_deco1[14]), .Z(n_39643));
	notech_inv i_53253(.A(n_3546), .Z(n_39644));
	notech_inv i_53254(.A(inst_deco1[15]), .Z(n_39645));
	notech_inv i_53255(.A(n_3545), .Z(n_39646));
	notech_inv i_53256(.A(inst_deco1[16]), .Z(n_39647));
	notech_inv i_53257(.A(n_3544), .Z(n_39648));
	notech_inv i_53258(.A(inst_deco1[17]), .Z(n_39649));
	notech_inv i_53259(.A(n_3543), .Z(n_39650));
	notech_inv i_53260(.A(n_50029), .Z(n_39651));
	notech_inv i_53261(.A(inst_deco1[18]), .Z(n_39652));
	notech_inv i_53262(.A(n_3542), .Z(n_39653));
	notech_inv i_53263(.A(inst_deco1[19]), .Z(n_39654));
	notech_inv i_53264(.A(n_3541), .Z(n_39655));
	notech_inv i_53265(.A(inst_deco1[20]), .Z(n_39656));
	notech_inv i_53266(.A(n_3540), .Z(n_39657));
	notech_inv i_53267(.A(inst_deco1[21]), .Z(n_39658));
	notech_inv i_53268(.A(n_50053), .Z(n_39659));
	notech_inv i_53269(.A(inst_deco1[22]), .Z(n_39660));
	notech_inv i_53270(.A(n_3539), .Z(n_39661));
	notech_inv i_53271(.A(n_50059), .Z(n_39662));
	notech_inv i_53272(.A(inst_deco1[23]), .Z(n_39663));
	notech_inv i_53273(.A(n_50065), .Z(n_39664));
	notech_inv i_53274(.A(inst_deco1[24]), .Z(n_39665));
	notech_inv i_53275(.A(n_3538), .Z(n_39666));
	notech_inv i_53276(.A(n_50071), .Z(n_39667));
	notech_inv i_53277(.A(inst_deco1[25]), .Z(n_39668));
	notech_inv i_53278(.A(n_3537), .Z(n_39669));
	notech_inv i_53279(.A(inst_deco1[26]), .Z(n_39670));
	notech_inv i_53280(.A(n_3536), .Z(n_39671));
	notech_inv i_53281(.A(inst_deco1[27]), .Z(n_39672));
	notech_inv i_53282(.A(n_3535), .Z(n_39673));
	notech_inv i_53283(.A(inst_deco1[28]), .Z(n_39674));
	notech_inv i_53284(.A(n_3533), .Z(n_39675));
	notech_inv i_53285(.A(inst_deco1[29]), .Z(n_39676));
	notech_inv i_53286(.A(n_3532), .Z(n_39677));
	notech_inv i_53287(.A(inst_deco1[30]), .Z(n_39678));
	notech_inv i_53288(.A(n_3531), .Z(n_39679));
	notech_inv i_53289(.A(inst_deco1[31]), .Z(n_39680));
	notech_inv i_53290(.A(n_50113), .Z(n_39681));
	notech_inv i_53291(.A(inst_deco1[32]), .Z(n_39682));
	notech_inv i_53292(.A(n_3530), .Z(n_39683));
	notech_inv i_53293(.A(inst_deco1[33]), .Z(n_39684));
	notech_inv i_53294(.A(n_3529), .Z(n_39685));
	notech_inv i_53295(.A(inst_deco1[34]), .Z(n_39686));
	notech_inv i_53296(.A(n_3528), .Z(n_39687));
	notech_inv i_53297(.A(inst_deco1[35]), .Z(n_39688));
	notech_inv i_53298(.A(n_3527), .Z(n_39689));
	notech_inv i_53299(.A(inst_deco1[36]), .Z(n_39690));
	notech_inv i_53300(.A(n_3525), .Z(n_39691));
	notech_inv i_53301(.A(n_50143), .Z(n_39692));
	notech_inv i_53302(.A(inst_deco1[37]), .Z(n_39693));
	notech_inv i_53303(.A(n_3524), .Z(n_39694));
	notech_inv i_53304(.A(inst_deco1[38]), .Z(n_39695));
	notech_inv i_53305(.A(n_3522), .Z(n_39696));
	notech_inv i_53306(.A(inst_deco1[39]), .Z(n_39697));
	notech_inv i_53307(.A(n_3520), .Z(n_39698));
	notech_inv i_53308(.A(inst_deco1[40]), .Z(n_39699));
	notech_inv i_53309(.A(n_3518), .Z(n_39700));
	notech_inv i_53310(.A(inst_deco1[41]), .Z(n_39701));
	notech_inv i_53311(.A(n_3517), .Z(n_39702));
	notech_inv i_53312(.A(inst_deco1[42]), .Z(n_39703));
	notech_inv i_53313(.A(n_3515), .Z(n_39704));
	notech_inv i_53314(.A(inst_deco1[43]), .Z(n_39705));
	notech_inv i_53315(.A(n_3513), .Z(n_39706));
	notech_inv i_53316(.A(inst_deco1[44]), .Z(n_39707));
	notech_inv i_53317(.A(n_3511), .Z(n_39708));
	notech_inv i_53318(.A(inst_deco1[45]), .Z(n_39709));
	notech_inv i_53319(.A(n_3510), .Z(n_39710));
	notech_inv i_53320(.A(inst_deco1[46]), .Z(n_39711));
	notech_inv i_53321(.A(n_3508), .Z(n_39712));
	notech_inv i_53322(.A(inst_deco1[47]), .Z(n_39713));
	notech_inv i_53323(.A(n_3506), .Z(n_39714));
	notech_inv i_53324(.A(inst_deco1[48]), .Z(n_39715));
	notech_inv i_53325(.A(n_3504), .Z(n_39716));
	notech_inv i_53326(.A(inst_deco1[49]), .Z(n_39717));
	notech_inv i_53327(.A(n_3502), .Z(n_39718));
	notech_inv i_53328(.A(inst_deco1[50]), .Z(n_39719));
	notech_inv i_53329(.A(n_3500), .Z(n_39720));
	notech_inv i_53330(.A(inst_deco1[51]), .Z(n_39721));
	notech_inv i_53331(.A(n_3498), .Z(n_39722));
	notech_inv i_53332(.A(inst_deco1[52]), .Z(n_39723));
	notech_inv i_53333(.A(n_3496), .Z(n_39724));
	notech_inv i_53334(.A(inst_deco1[53]), .Z(n_39725));
	notech_inv i_53335(.A(n_3494), .Z(n_39726));
	notech_inv i_53336(.A(inst_deco1[54]), .Z(n_39727));
	notech_inv i_53337(.A(n_3492), .Z(n_39728));
	notech_inv i_53338(.A(inst_deco1[55]), .Z(n_39729));
	notech_inv i_53339(.A(n_3490), .Z(n_39730));
	notech_inv i_53340(.A(inst_deco1[56]), .Z(n_39731));
	notech_inv i_53341(.A(n_3488), .Z(n_39732));
	notech_inv i_53342(.A(inst_deco1[57]), .Z(n_39733));
	notech_inv i_53343(.A(n_3486), .Z(n_39734));
	notech_inv i_53344(.A(inst_deco1[58]), .Z(n_39735));
	notech_inv i_53345(.A(n_3484), .Z(n_39736));
	notech_inv i_53346(.A(inst_deco1[59]), .Z(n_39737));
	notech_inv i_53347(.A(n_3482), .Z(n_39738));
	notech_inv i_53348(.A(inst_deco1[60]), .Z(n_39739));
	notech_inv i_53349(.A(n_3480), .Z(n_39740));
	notech_inv i_53350(.A(inst_deco1[61]), .Z(n_39741));
	notech_inv i_53351(.A(n_3478), .Z(n_39742));
	notech_inv i_53352(.A(inst_deco1[62]), .Z(n_39743));
	notech_inv i_53353(.A(n_3476), .Z(n_39744));
	notech_inv i_53354(.A(inst_deco1[63]), .Z(n_39745));
	notech_inv i_53355(.A(n_3474), .Z(n_39746));
	notech_inv i_53356(.A(inst_deco1[64]), .Z(n_39747));
	notech_inv i_53357(.A(n_3472), .Z(n_39748));
	notech_inv i_53358(.A(inst_deco1[65]), .Z(n_39749));
	notech_inv i_53359(.A(n_3470), .Z(n_39750));
	notech_inv i_53360(.A(inst_deco1[66]), .Z(n_39751));
	notech_inv i_53361(.A(n_3468), .Z(n_39752));
	notech_inv i_53362(.A(inst_deco1[67]), .Z(n_39753));
	notech_inv i_53363(.A(n_3466), .Z(n_39754));
	notech_inv i_53364(.A(inst_deco1[68]), .Z(n_39755));
	notech_inv i_53365(.A(n_3464), .Z(n_39756));
	notech_inv i_53366(.A(inst_deco1[69]), .Z(n_39757));
	notech_inv i_53367(.A(n_3462), .Z(n_39758));
	notech_inv i_53368(.A(inst_deco1[70]), .Z(n_39759));
	notech_inv i_53369(.A(n_3460), .Z(n_39760));
	notech_inv i_53370(.A(inst_deco1[71]), .Z(n_39761));
	notech_inv i_53371(.A(n_3459), .Z(n_39762));
	notech_inv i_53372(.A(n_3458), .Z(n_39763));
	notech_inv i_53373(.A(inst_deco1[73]), .Z(n_39764));
	notech_inv i_53374(.A(n_3457), .Z(n_39765));
	notech_inv i_53375(.A(inst_deco1[74]), .Z(n_39766));
	notech_inv i_53376(.A(n_3456), .Z(n_39767));
	notech_inv i_53377(.A(inst_deco1[75]), .Z(n_39768));
	notech_inv i_53378(.A(n_3455), .Z(n_39769));
	notech_inv i_53379(.A(inst_deco1[76]), .Z(n_39770));
	notech_inv i_53380(.A(n_3454), .Z(n_39771));
	notech_inv i_53381(.A(inst_deco1[77]), .Z(n_39772));
	notech_inv i_53382(.A(n_3453), .Z(n_39773));
	notech_inv i_53383(.A(inst_deco1[78]), .Z(n_39774));
	notech_inv i_53384(.A(n_3452), .Z(n_39775));
	notech_inv i_53385(.A(inst_deco1[79]), .Z(n_39776));
	notech_inv i_53386(.A(n_3451), .Z(n_39777));
	notech_inv i_53387(.A(n_3450), .Z(n_39778));
	notech_inv i_53388(.A(n_3449), .Z(n_39779));
	notech_inv i_53389(.A(n_3448), .Z(n_39780));
	notech_inv i_53390(.A(n_3447), .Z(n_39781));
	notech_inv i_53391(.A(n_3446), .Z(n_39782));
	notech_inv i_53392(.A(n_3445), .Z(n_39783));
	notech_inv i_53393(.A(n_3444), .Z(n_39784));
	notech_inv i_53394(.A(n_3443), .Z(n_39785));
	notech_inv i_53395(.A(inst_deco1[88]), .Z(n_39786));
	notech_inv i_53396(.A(n_3442), .Z(n_39787));
	notech_inv i_53397(.A(inst_deco1[89]), .Z(n_39788));
	notech_inv i_53398(.A(n_3441), .Z(n_39789));
	notech_inv i_53399(.A(inst_deco1[90]), .Z(n_39790));
	notech_inv i_53400(.A(n_3439), .Z(n_39791));
	notech_inv i_53401(.A(n_3438), .Z(n_39792));
	notech_inv i_53402(.A(inst_deco1[92]), .Z(n_39793));
	notech_inv i_53403(.A(n_3437), .Z(n_39794));
	notech_inv i_53404(.A(inst_deco1[93]), .Z(n_39795));
	notech_inv i_53405(.A(n_3436), .Z(n_39796));
	notech_inv i_53406(.A(inst_deco1[94]), .Z(n_39797));
	notech_inv i_53407(.A(n_3434), .Z(n_39798));
	notech_inv i_53408(.A(inst_deco1[95]), .Z(n_39799));
	notech_inv i_53409(.A(n_3433), .Z(n_39800));
	notech_inv i_53410(.A(inst_deco1[96]), .Z(n_39801));
	notech_inv i_53411(.A(n_3432), .Z(n_39802));
	notech_inv i_53412(.A(inst_deco1[97]), .Z(n_39803));
	notech_inv i_53413(.A(n_3430), .Z(n_39804));
	notech_inv i_53414(.A(inst_deco1[98]), .Z(n_39805));
	notech_inv i_53415(.A(n_3429), .Z(n_39806));
	notech_inv i_53416(.A(inst_deco1[99]), .Z(n_39807));
	notech_inv i_53417(.A(n_3427), .Z(n_39808));
	notech_inv i_53418(.A(inst_deco1[100]), .Z(n_39809));
	notech_inv i_53419(.A(n_3425), .Z(n_39810));
	notech_inv i_53420(.A(inst_deco1[101]), .Z(n_39811));
	notech_inv i_53421(.A(n_3423), .Z(n_39812));
	notech_inv i_53422(.A(inst_deco1[102]), .Z(n_39813));
	notech_inv i_53423(.A(n_3421), .Z(n_39814));
	notech_inv i_53424(.A(inst_deco1[103]), .Z(n_39815));
	notech_inv i_53425(.A(n_3419), .Z(n_39816));
	notech_inv i_53426(.A(inst_deco1[104]), .Z(n_39817));
	notech_inv i_53427(.A(n_3417), .Z(n_39818));
	notech_inv i_53428(.A(inst_deco1[105]), .Z(n_39819));
	notech_inv i_53429(.A(n_3415), .Z(n_39820));
	notech_inv i_53430(.A(n_3413), .Z(n_39821));
	notech_inv i_53431(.A(inst_deco1[107]), .Z(n_39822));
	notech_inv i_53432(.A(n_3411), .Z(n_39823));
	notech_inv i_53433(.A(inst_deco1[108]), .Z(n_39824));
	notech_inv i_53434(.A(n_3409), .Z(n_39825));
	notech_inv i_53435(.A(inst_deco1[109]), .Z(n_39826));
	notech_inv i_53436(.A(n_3407), .Z(n_39827));
	notech_inv i_53437(.A(inst_deco1[110]), .Z(n_39828));
	notech_inv i_53438(.A(n_3405), .Z(n_39829));
	notech_inv i_53439(.A(inst_deco1[111]), .Z(n_39830));
	notech_inv i_53440(.A(n_3403), .Z(n_39831));
	notech_inv i_53441(.A(inst_deco1[112]), .Z(n_39832));
	notech_inv i_53442(.A(n_3401), .Z(n_39833));
	notech_inv i_53443(.A(n_3399), .Z(n_39834));
	notech_inv i_53444(.A(inst_deco1[114]), .Z(n_39835));
	notech_inv i_53445(.A(n_3397), .Z(n_39836));
	notech_inv i_53446(.A(inst_deco1[115]), .Z(n_39837));
	notech_inv i_53447(.A(n_3395), .Z(n_39838));
	notech_inv i_53448(.A(inst_deco1[116]), .Z(n_39839));
	notech_inv i_53449(.A(n_3393), .Z(n_39840));
	notech_inv i_53450(.A(inst_deco1[117]), .Z(n_39841));
	notech_inv i_53451(.A(n_3391), .Z(n_39842));
	notech_inv i_53452(.A(inst_deco1[118]), .Z(n_39843));
	notech_inv i_53453(.A(n_3389), .Z(n_39844));
	notech_inv i_53454(.A(inst_deco1[119]), .Z(n_39845));
	notech_inv i_53455(.A(n_3387), .Z(n_39846));
	notech_inv i_53456(.A(inst_deco1[120]), .Z(n_39847));
	notech_inv i_53457(.A(n_3385), .Z(n_39848));
	notech_inv i_53458(.A(inst_deco1[121]), .Z(n_39849));
	notech_inv i_53459(.A(n_3383), .Z(n_39850));
	notech_inv i_53460(.A(inst_deco1[122]), .Z(n_39851));
	notech_inv i_53461(.A(n_3381), .Z(n_39852));
	notech_inv i_53462(.A(inst_deco1[123]), .Z(n_39853));
	notech_inv i_53463(.A(n_3379), .Z(n_39854));
	notech_inv i_53464(.A(inst_deco1[124]), .Z(n_39855));
	notech_inv i_53465(.A(n_3377), .Z(n_39856));
	notech_inv i_53466(.A(inst_deco1[125]), .Z(n_39857));
	notech_inv i_53467(.A(n_3375), .Z(n_39858));
	notech_inv i_53468(.A(inst_deco1[126]), .Z(n_39859));
	notech_inv i_53469(.A(n_3373), .Z(n_39860));
	notech_inv i_53470(.A(inst_deco1[127]), .Z(n_39861));
	notech_inv i_53471(.A(to_acu2[0]), .Z(n_39862));
	notech_inv i_53472(.A(n_3371), .Z(n_39863));
	notech_inv i_53473(.A(to_acu2[1]), .Z(n_39864));
	notech_inv i_53474(.A(to_acu2[2]), .Z(n_39865));
	notech_inv i_53475(.A(n_3369), .Z(n_39866));
	notech_inv i_53476(.A(to_acu2[3]), .Z(n_39867));
	notech_inv i_53477(.A(to_acu2[4]), .Z(n_39868));
	notech_inv i_53478(.A(n_3367), .Z(n_39869));
	notech_inv i_53479(.A(to_acu2[5]), .Z(n_39870));
	notech_inv i_53480(.A(to_acu2[6]), .Z(n_39871));
	notech_inv i_53481(.A(n_3365), .Z(n_39872));
	notech_inv i_53482(.A(to_acu2[7]), .Z(n_39873));
	notech_inv i_53483(.A(to_acu2[8]), .Z(n_39874));
	notech_inv i_53484(.A(n_3363), .Z(n_39875));
	notech_inv i_53485(.A(to_acu2[9]), .Z(n_39876));
	notech_inv i_53486(.A(to_acu2[10]), .Z(n_39877));
	notech_inv i_53487(.A(n_3361), .Z(n_39878));
	notech_inv i_53488(.A(to_acu2[11]), .Z(n_39879));
	notech_inv i_53489(.A(to_acu2[12]), .Z(n_39880));
	notech_inv i_53490(.A(n_3359), .Z(n_39881));
	notech_inv i_53491(.A(to_acu2[13]), .Z(n_39882));
	notech_inv i_53492(.A(to_acu2[14]), .Z(n_39883));
	notech_inv i_53493(.A(n_3357), .Z(n_39884));
	notech_inv i_53494(.A(to_acu2[15]), .Z(n_39885));
	notech_inv i_53495(.A(to_acu2[16]), .Z(n_39886));
	notech_inv i_53496(.A(n_3355), .Z(n_39887));
	notech_inv i_53497(.A(to_acu2[17]), .Z(n_39888));
	notech_inv i_53498(.A(to_acu2[18]), .Z(n_39889));
	notech_inv i_53499(.A(n_3353), .Z(n_39890));
	notech_inv i_53500(.A(to_acu2[19]), .Z(n_39891));
	notech_inv i_53501(.A(to_acu2[20]), .Z(n_39892));
	notech_inv i_53502(.A(n_3351), .Z(n_39893));
	notech_inv i_53503(.A(to_acu2[21]), .Z(n_39894));
	notech_inv i_53504(.A(to_acu2[22]), .Z(n_39895));
	notech_inv i_53505(.A(n_3349), .Z(n_39896));
	notech_inv i_53506(.A(to_acu2[23]), .Z(n_39897));
	notech_inv i_53507(.A(to_acu2[24]), .Z(n_39898));
	notech_inv i_53508(.A(n_3348), .Z(n_39899));
	notech_inv i_53509(.A(to_acu2[25]), .Z(n_39900));
	notech_inv i_53510(.A(to_acu2[26]), .Z(n_39901));
	notech_inv i_53511(.A(n_3347), .Z(n_39902));
	notech_inv i_53512(.A(to_acu2[27]), .Z(n_39903));
	notech_inv i_53513(.A(to_acu2[28]), .Z(n_39904));
	notech_inv i_53514(.A(n_3346), .Z(n_39905));
	notech_inv i_53515(.A(to_acu2[29]), .Z(n_39906));
	notech_inv i_53516(.A(to_acu2[30]), .Z(n_39907));
	notech_inv i_53517(.A(n_3345), .Z(n_39908));
	notech_inv i_53518(.A(to_acu2[31]), .Z(n_39909));
	notech_inv i_53519(.A(to_acu2[32]), .Z(n_39910));
	notech_inv i_53520(.A(n_3344), .Z(n_39911));
	notech_inv i_53521(.A(to_acu2[33]), .Z(n_39912));
	notech_inv i_53522(.A(to_acu2[34]), .Z(n_39913));
	notech_inv i_53523(.A(n_3343), .Z(n_39914));
	notech_inv i_53524(.A(to_acu2[35]), .Z(n_39915));
	notech_inv i_53525(.A(to_acu2[36]), .Z(n_39916));
	notech_inv i_53526(.A(n_3342), .Z(n_39917));
	notech_inv i_53527(.A(to_acu2[37]), .Z(n_39918));
	notech_inv i_53528(.A(to_acu2[38]), .Z(n_39919));
	notech_inv i_53529(.A(n_3341), .Z(n_39920));
	notech_inv i_53530(.A(to_acu2[40]), .Z(n_39921));
	notech_inv i_53531(.A(n_3340), .Z(n_39922));
	notech_inv i_53532(.A(to_acu2[41]), .Z(n_39923));
	notech_inv i_53533(.A(to_acu2[42]), .Z(n_39924));
	notech_inv i_53534(.A(n_3339), .Z(n_39925));
	notech_inv i_53535(.A(to_acu2[43]), .Z(n_39926));
	notech_inv i_53536(.A(to_acu2[44]), .Z(n_39927));
	notech_inv i_53537(.A(n_3338), .Z(n_39928));
	notech_inv i_53538(.A(to_acu2[45]), .Z(n_39929));
	notech_inv i_53539(.A(to_acu2[46]), .Z(n_39930));
	notech_inv i_53540(.A(n_3337), .Z(n_39931));
	notech_inv i_53541(.A(to_acu2[47]), .Z(n_39932));
	notech_inv i_53542(.A(to_acu2[48]), .Z(n_39933));
	notech_inv i_53543(.A(n_3336), .Z(n_39934));
	notech_inv i_53544(.A(to_acu2[49]), .Z(n_39935));
	notech_inv i_53545(.A(to_acu2[50]), .Z(n_39936));
	notech_inv i_53546(.A(n_3335), .Z(n_39937));
	notech_inv i_53547(.A(to_acu2[51]), .Z(n_39938));
	notech_inv i_53548(.A(to_acu2[52]), .Z(n_39939));
	notech_inv i_53549(.A(n_3334), .Z(n_39940));
	notech_inv i_53550(.A(to_acu2[53]), .Z(n_39941));
	notech_inv i_53551(.A(to_acu2[54]), .Z(n_39942));
	notech_inv i_53552(.A(n_3333), .Z(n_39943));
	notech_inv i_53553(.A(to_acu2[55]), .Z(n_39944));
	notech_inv i_53554(.A(to_acu2[56]), .Z(n_39945));
	notech_inv i_53555(.A(n_3331), .Z(n_39946));
	notech_inv i_53556(.A(to_acu2[57]), .Z(n_39947));
	notech_inv i_53557(.A(to_acu2[58]), .Z(n_39948));
	notech_inv i_53558(.A(n_3330), .Z(n_39949));
	notech_inv i_53559(.A(to_acu2[59]), .Z(n_39950));
	notech_inv i_53560(.A(to_acu2[60]), .Z(n_39951));
	notech_inv i_53561(.A(n_3328), .Z(n_39952));
	notech_inv i_53562(.A(to_acu2[61]), .Z(n_39953));
	notech_inv i_53563(.A(to_acu2[62]), .Z(n_39954));
	notech_inv i_53564(.A(n_3327), .Z(n_39955));
	notech_inv i_53565(.A(to_acu2[63]), .Z(n_39956));
	notech_inv i_53566(.A(to_acu2[64]), .Z(n_39957));
	notech_inv i_53567(.A(n_3325), .Z(n_39958));
	notech_inv i_53568(.A(to_acu2[65]), .Z(n_39959));
	notech_inv i_53569(.A(to_acu2[66]), .Z(n_39960));
	notech_inv i_53570(.A(n_3324), .Z(n_39961));
	notech_inv i_53571(.A(to_acu2[67]), .Z(n_39962));
	notech_inv i_53572(.A(to_acu2[68]), .Z(n_39963));
	notech_inv i_53573(.A(n_3323), .Z(n_39964));
	notech_inv i_53574(.A(to_acu2[69]), .Z(n_39965));
	notech_inv i_53575(.A(to_acu2[70]), .Z(n_39966));
	notech_inv i_53576(.A(n_3322), .Z(n_39967));
	notech_inv i_53577(.A(to_acu2[71]), .Z(n_39968));
	notech_inv i_53578(.A(to_acu2[72]), .Z(n_39969));
	notech_inv i_53579(.A(n_3321), .Z(n_39970));
	notech_inv i_53580(.A(to_acu2[73]), .Z(n_39971));
	notech_inv i_53581(.A(to_acu2[74]), .Z(n_39972));
	notech_inv i_53582(.A(n_3320), .Z(n_39973));
	notech_inv i_53583(.A(to_acu2[75]), .Z(n_39974));
	notech_inv i_53584(.A(to_acu2[76]), .Z(n_39975));
	notech_inv i_53585(.A(n_3319), .Z(n_39976));
	notech_inv i_53586(.A(to_acu2[77]), .Z(n_39977));
	notech_inv i_53587(.A(to_acu2[78]), .Z(n_39978));
	notech_inv i_53588(.A(n_3318), .Z(n_39979));
	notech_inv i_53589(.A(to_acu2[79]), .Z(n_39980));
	notech_inv i_53590(.A(to_acu2[80]), .Z(n_39981));
	notech_inv i_53591(.A(n_3317), .Z(n_39982));
	notech_inv i_53592(.A(to_acu2[81]), .Z(n_39983));
	notech_inv i_53593(.A(to_acu2[82]), .Z(n_39984));
	notech_inv i_53594(.A(n_3316), .Z(n_39985));
	notech_inv i_53595(.A(to_acu2[83]), .Z(n_39986));
	notech_inv i_53596(.A(n_47642), .Z(n_39987));
	notech_inv i_53597(.A(to_acu2[84]), .Z(n_39988));
	notech_inv i_53598(.A(n_3315), .Z(n_39989));
	notech_inv i_53599(.A(to_acu2[85]), .Z(n_39990));
	notech_inv i_53600(.A(to_acu2[86]), .Z(n_39991));
	notech_inv i_53601(.A(n_3314), .Z(n_39992));
	notech_inv i_53602(.A(to_acu2[87]), .Z(n_39993));
	notech_inv i_53603(.A(to_acu2[88]), .Z(n_39994));
	notech_inv i_53604(.A(n_3313), .Z(n_39995));
	notech_inv i_53605(.A(to_acu2[89]), .Z(n_39996));
	notech_inv i_53606(.A(n_3312), .Z(n_39997));
	notech_inv i_53607(.A(to_acu2[90]), .Z(n_39998));
	notech_inv i_53608(.A(n_3311), .Z(n_39999));
	notech_inv i_53609(.A(to_acu2[91]), .Z(n_40000));
	notech_inv i_53610(.A(n_3310), .Z(n_40001));
	notech_inv i_53611(.A(to_acu2[92]), .Z(n_40002));
	notech_inv i_53612(.A(n_3309), .Z(n_40003));
	notech_inv i_53613(.A(to_acu2[93]), .Z(n_40004));
	notech_inv i_53614(.A(n_3308), .Z(n_40005));
	notech_inv i_53615(.A(to_acu2[94]), .Z(n_40006));
	notech_inv i_53616(.A(n_3307), .Z(n_40007));
	notech_inv i_53617(.A(to_acu2[95]), .Z(n_40008));
	notech_inv i_53618(.A(n_3305), .Z(n_40009));
	notech_inv i_53619(.A(to_acu2[96]), .Z(n_40010));
	notech_inv i_53620(.A(n_3304), .Z(n_40011));
	notech_inv i_53621(.A(to_acu2[97]), .Z(n_40012));
	notech_inv i_53622(.A(n_3303), .Z(n_40013));
	notech_inv i_53623(.A(to_acu2[98]), .Z(n_40014));
	notech_inv i_53624(.A(n_3301), .Z(n_40015));
	notech_inv i_53625(.A(to_acu2[99]), .Z(n_40016));
	notech_inv i_53626(.A(n_3300), .Z(n_40017));
	notech_inv i_53627(.A(to_acu2[100]), .Z(n_40018));
	notech_inv i_53628(.A(n_3299), .Z(n_40019));
	notech_inv i_53629(.A(to_acu2[101]), .Z(n_40020));
	notech_inv i_53630(.A(n_3298), .Z(n_40021));
	notech_inv i_53631(.A(to_acu2[102]), .Z(n_40022));
	notech_inv i_53632(.A(n_3297), .Z(n_40023));
	notech_inv i_53633(.A(to_acu2[103]), .Z(n_40024));
	notech_inv i_53634(.A(n_3296), .Z(n_40025));
	notech_inv i_53635(.A(to_acu2[104]), .Z(n_40026));
	notech_inv i_53636(.A(n_3295), .Z(n_40027));
	notech_inv i_53637(.A(to_acu2[105]), .Z(n_40028));
	notech_inv i_53638(.A(n_3294), .Z(n_40029));
	notech_inv i_53639(.A(to_acu2[106]), .Z(n_40030));
	notech_inv i_53640(.A(to_acu2[107]), .Z(n_40031));
	notech_inv i_53641(.A(n_3293), .Z(n_40032));
	notech_inv i_53642(.A(to_acu2[108]), .Z(n_40033));
	notech_inv i_53643(.A(n_3292), .Z(n_40034));
	notech_inv i_53644(.A(to_acu2[109]), .Z(n_40035));
	notech_inv i_53645(.A(to_acu2[110]), .Z(n_40036));
	notech_inv i_53646(.A(n_3291), .Z(n_40037));
	notech_inv i_53647(.A(to_acu2[111]), .Z(n_40038));
	notech_inv i_53648(.A(to_acu2[112]), .Z(n_40039));
	notech_inv i_53649(.A(n_3290), .Z(n_40040));
	notech_inv i_53650(.A(to_acu2[113]), .Z(n_40041));
	notech_inv i_53651(.A(to_acu2[114]), .Z(n_40042));
	notech_inv i_53652(.A(n_3289), .Z(n_40043));
	notech_inv i_53653(.A(to_acu2[115]), .Z(n_40044));
	notech_inv i_53654(.A(to_acu2[116]), .Z(n_40045));
	notech_inv i_53655(.A(n_3288), .Z(n_40046));
	notech_inv i_53656(.A(to_acu2[117]), .Z(n_40047));
	notech_inv i_53657(.A(to_acu2[118]), .Z(n_40048));
	notech_inv i_53658(.A(n_3287), .Z(n_40049));
	notech_inv i_53659(.A(to_acu2[119]), .Z(n_40050));
	notech_inv i_53660(.A(to_acu2[120]), .Z(n_40051));
	notech_inv i_53661(.A(n_3286), .Z(n_40052));
	notech_inv i_53662(.A(to_acu2[121]), .Z(n_40053));
	notech_inv i_53663(.A(to_acu2[122]), .Z(n_40054));
	notech_inv i_53664(.A(n_3285), .Z(n_40055));
	notech_inv i_53665(.A(to_acu2[123]), .Z(n_40056));
	notech_inv i_53666(.A(to_acu2[124]), .Z(n_40057));
	notech_inv i_53667(.A(n_3284), .Z(n_40058));
	notech_inv i_53668(.A(to_acu2[125]), .Z(n_40059));
	notech_inv i_53669(.A(to_acu2[126]), .Z(n_40060));
	notech_inv i_53670(.A(n_3283), .Z(n_40061));
	notech_inv i_53671(.A(to_acu2[127]), .Z(n_40062));
	notech_inv i_53672(.A(to_acu2[128]), .Z(n_40063));
	notech_inv i_53673(.A(n_3282), .Z(n_40064));
	notech_inv i_53674(.A(to_acu2[129]), .Z(n_40065));
	notech_inv i_53675(.A(to_acu2[130]), .Z(n_40066));
	notech_inv i_53676(.A(n_3281), .Z(n_40067));
	notech_inv i_53677(.A(to_acu2[131]), .Z(n_40068));
	notech_inv i_53678(.A(to_acu2[132]), .Z(n_40069));
	notech_inv i_53679(.A(n_3280), .Z(n_40070));
	notech_inv i_53680(.A(to_acu2[133]), .Z(n_40071));
	notech_inv i_53681(.A(to_acu2[134]), .Z(n_40072));
	notech_inv i_53682(.A(n_3279), .Z(n_40073));
	notech_inv i_53683(.A(to_acu2[135]), .Z(n_40074));
	notech_inv i_53684(.A(to_acu2[136]), .Z(n_40075));
	notech_inv i_53685(.A(to_acu2[137]), .Z(n_40076));
	notech_inv i_53686(.A(to_acu2[138]), .Z(n_40077));
	notech_inv i_53687(.A(to_acu2[139]), .Z(n_40078));
	notech_inv i_53688(.A(to_acu2[140]), .Z(n_40079));
	notech_inv i_53689(.A(to_acu2[141]), .Z(n_40080));
	notech_inv i_53690(.A(to_acu2[142]), .Z(n_40081));
	notech_inv i_53691(.A(n_3272), .Z(n_40082));
	notech_inv i_53692(.A(to_acu2[143]), .Z(n_40083));
	notech_inv i_53693(.A(to_acu2[144]), .Z(n_40084));
	notech_inv i_53694(.A(n_3271), .Z(n_40085));
	notech_inv i_53695(.A(to_acu2[145]), .Z(n_40086));
	notech_inv i_53696(.A(to_acu2[146]), .Z(n_40087));
	notech_inv i_53697(.A(to_acu2[147]), .Z(n_40088));
	notech_inv i_53698(.A(to_acu2[148]), .Z(n_40089));
	notech_inv i_53699(.A(to_acu2[149]), .Z(n_40090));
	notech_inv i_53700(.A(to_acu2[150]), .Z(n_40091));
	notech_inv i_53701(.A(to_acu2[151]), .Z(n_40092));
	notech_inv i_53702(.A(to_acu2[152]), .Z(n_40093));
	notech_inv i_53703(.A(to_acu2[153]), .Z(n_40094));
	notech_inv i_53704(.A(to_acu2[154]), .Z(n_40095));
	notech_inv i_53705(.A(to_acu2[155]), .Z(n_40096));
	notech_inv i_53706(.A(to_acu2[156]), .Z(n_40097));
	notech_inv i_53707(.A(to_acu2[157]), .Z(n_40098));
	notech_inv i_53708(.A(to_acu2[158]), .Z(n_40099));
	notech_inv i_53709(.A(to_acu2[159]), .Z(n_40100));
	notech_inv i_53710(.A(to_acu2[160]), .Z(n_40101));
	notech_inv i_53711(.A(to_acu2[161]), .Z(n_40102));
	notech_inv i_53712(.A(to_acu2[162]), .Z(n_40103));
	notech_inv i_53713(.A(to_acu2[163]), .Z(n_40104));
	notech_inv i_53714(.A(to_acu2[164]), .Z(n_40105));
	notech_inv i_53715(.A(to_acu2[165]), .Z(n_40106));
	notech_inv i_53716(.A(to_acu2[166]), .Z(n_40107));
	notech_inv i_53717(.A(to_acu2[167]), .Z(n_40108));
	notech_inv i_53718(.A(to_acu2[168]), .Z(n_40109));
	notech_inv i_53719(.A(to_acu2[169]), .Z(n_40110));
	notech_inv i_53720(.A(to_acu2[170]), .Z(n_40111));
	notech_inv i_53721(.A(n_3242), .Z(n_40112));
	notech_inv i_53722(.A(to_acu2[171]), .Z(n_40113));
	notech_inv i_53723(.A(to_acu2[172]), .Z(n_40114));
	notech_inv i_53724(.A(n_3241), .Z(n_40115));
	notech_inv i_53725(.A(to_acu2[173]), .Z(n_40116));
	notech_inv i_53726(.A(to_acu2[174]), .Z(n_40117));
	notech_inv i_53727(.A(n_3240), .Z(n_40118));
	notech_inv i_53728(.A(to_acu2[175]), .Z(n_40119));
	notech_inv i_53729(.A(to_acu2[176]), .Z(n_40120));
	notech_inv i_53730(.A(n_3238), .Z(n_40121));
	notech_inv i_53731(.A(to_acu2[177]), .Z(n_40122));
	notech_inv i_53732(.A(to_acu2[178]), .Z(n_40123));
	notech_inv i_53733(.A(n_3236), .Z(n_40124));
	notech_inv i_53734(.A(to_acu2[179]), .Z(n_40125));
	notech_inv i_53735(.A(to_acu2[180]), .Z(n_40126));
	notech_inv i_53736(.A(n_3235), .Z(n_40127));
	notech_inv i_53737(.A(to_acu2[181]), .Z(n_40128));
	notech_inv i_53738(.A(to_acu2[182]), .Z(n_40129));
	notech_inv i_53739(.A(n_3234), .Z(n_40130));
	notech_inv i_53740(.A(to_acu2[183]), .Z(n_40131));
	notech_inv i_53741(.A(to_acu2[184]), .Z(n_40132));
	notech_inv i_53742(.A(n_3233), .Z(n_40133));
	notech_inv i_53743(.A(to_acu2[185]), .Z(n_40134));
	notech_inv i_53744(.A(to_acu2[186]), .Z(n_40135));
	notech_inv i_53745(.A(n_3232), .Z(n_40136));
	notech_inv i_53746(.A(to_acu2[187]), .Z(n_40137));
	notech_inv i_53747(.A(to_acu2[188]), .Z(n_40138));
	notech_inv i_53748(.A(n_3231), .Z(n_40139));
	notech_inv i_53749(.A(to_acu2[189]), .Z(n_40140));
	notech_inv i_53750(.A(to_acu2[190]), .Z(n_40141));
	notech_inv i_53751(.A(n_3230), .Z(n_40142));
	notech_inv i_53752(.A(to_acu2[191]), .Z(n_40143));
	notech_inv i_53753(.A(to_acu2[192]), .Z(n_40144));
	notech_inv i_53754(.A(n_3229), .Z(n_40145));
	notech_inv i_53755(.A(to_acu2[193]), .Z(n_40146));
	notech_inv i_53756(.A(to_acu2[194]), .Z(n_40147));
	notech_inv i_53757(.A(n_3228), .Z(n_40148));
	notech_inv i_53758(.A(to_acu2[195]), .Z(n_40149));
	notech_inv i_53759(.A(to_acu2[196]), .Z(n_40150));
	notech_inv i_53760(.A(n_3227), .Z(n_40151));
	notech_inv i_53761(.A(to_acu2[197]), .Z(n_40152));
	notech_inv i_53762(.A(to_acu2[198]), .Z(n_40153));
	notech_inv i_53763(.A(n_3226), .Z(n_40154));
	notech_inv i_53764(.A(to_acu2[199]), .Z(n_40155));
	notech_inv i_53765(.A(to_acu2[200]), .Z(n_40156));
	notech_inv i_53766(.A(n_3225), .Z(n_40157));
	notech_inv i_53767(.A(to_acu2[201]), .Z(n_40158));
	notech_inv i_53768(.A(to_acu2[202]), .Z(n_40159));
	notech_inv i_53769(.A(n_3224), .Z(n_40160));
	notech_inv i_53770(.A(to_acu2[203]), .Z(n_40161));
	notech_inv i_53771(.A(to_acu2[204]), .Z(n_40162));
	notech_inv i_53772(.A(n_3223), .Z(n_40163));
	notech_inv i_53773(.A(to_acu2[205]), .Z(n_40164));
	notech_inv i_53774(.A(to_acu2[206]), .Z(n_40165));
	notech_inv i_53775(.A(n_3222), .Z(n_40166));
	notech_inv i_53776(.A(to_acu2[207]), .Z(n_40167));
	notech_inv i_53777(.A(to_acu2[208]), .Z(n_40168));
	notech_inv i_53778(.A(n_3221), .Z(n_40169));
	notech_inv i_53779(.A(to_acu2[209]), .Z(n_40170));
	notech_inv i_53780(.A(to_acu2[210]), .Z(n_40171));
	notech_inv i_53781(.A(n_3220), .Z(n_40172));
	notech_inv i_53782(.A(to_acu1[0]), .Z(n_40173));
	notech_inv i_53783(.A(n_3219), .Z(n_40174));
	notech_inv i_53784(.A(to_acu1[1]), .Z(n_40175));
	notech_inv i_53785(.A(n_3218), .Z(n_40176));
	notech_inv i_53786(.A(n_48453), .Z(n_40177));
	notech_inv i_53787(.A(to_acu1[2]), .Z(n_40178));
	notech_inv i_53788(.A(n_48459), .Z(n_40179));
	notech_inv i_53789(.A(to_acu1[3]), .Z(n_40180));
	notech_inv i_53790(.A(n_3217), .Z(n_40181));
	notech_inv i_53791(.A(n_48465), .Z(n_40182));
	notech_inv i_53792(.A(to_acu1[4]), .Z(n_40183));
	notech_inv i_53793(.A(n_3216), .Z(n_40184));
	notech_inv i_53794(.A(to_acu1[5]), .Z(n_40185));
	notech_inv i_53795(.A(n_3215), .Z(n_40186));
	notech_inv i_53796(.A(to_acu1[6]), .Z(n_40187));
	notech_inv i_53797(.A(n_48483), .Z(n_40188));
	notech_inv i_53798(.A(to_acu1[7]), .Z(n_40189));
	notech_inv i_53799(.A(n_3214), .Z(n_40190));
	notech_inv i_53800(.A(to_acu1[8]), .Z(n_40191));
	notech_inv i_53801(.A(n_3213), .Z(n_40192));
	notech_inv i_53802(.A(to_acu1[9]), .Z(n_40193));
	notech_inv i_53803(.A(n_3212), .Z(n_40194));
	notech_inv i_53804(.A(to_acu1[10]), .Z(n_40195));
	notech_inv i_53805(.A(n_3211), .Z(n_40196));
	notech_inv i_53806(.A(to_acu1[11]), .Z(n_40197));
	notech_inv i_53807(.A(n_3210), .Z(n_40198));
	notech_inv i_53808(.A(to_acu1[12]), .Z(n_40199));
	notech_inv i_53809(.A(n_3209), .Z(n_40200));
	notech_inv i_53810(.A(to_acu1[13]), .Z(n_40201));
	notech_inv i_53811(.A(n_3208), .Z(n_40202));
	notech_inv i_53812(.A(to_acu1[14]), .Z(n_40203));
	notech_inv i_53813(.A(n_3207), .Z(n_40204));
	notech_inv i_53814(.A(to_acu1[15]), .Z(n_40205));
	notech_inv i_53815(.A(n_3206), .Z(n_40206));
	notech_inv i_53816(.A(to_acu1[16]), .Z(n_40207));
	notech_inv i_53817(.A(n_3205), .Z(n_40208));
	notech_inv i_53818(.A(to_acu1[17]), .Z(n_40209));
	notech_inv i_53819(.A(n_3204), .Z(n_40210));
	notech_inv i_53820(.A(to_acu1[18]), .Z(n_40211));
	notech_inv i_53821(.A(n_3203), .Z(n_40212));
	notech_inv i_53822(.A(to_acu1[19]), .Z(n_40213));
	notech_inv i_53823(.A(n_3202), .Z(n_40214));
	notech_inv i_53824(.A(to_acu1[20]), .Z(n_40215));
	notech_inv i_53825(.A(n_3201), .Z(n_40216));
	notech_inv i_53826(.A(to_acu1[21]), .Z(n_40217));
	notech_inv i_53827(.A(n_3200), .Z(n_40218));
	notech_inv i_53828(.A(to_acu1[22]), .Z(n_40219));
	notech_inv i_53829(.A(n_3199), .Z(n_40220));
	notech_inv i_53830(.A(to_acu1[23]), .Z(n_40221));
	notech_inv i_53831(.A(n_3198), .Z(n_40222));
	notech_inv i_53832(.A(to_acu1[24]), .Z(n_40223));
	notech_inv i_53833(.A(n_3197), .Z(n_40224));
	notech_inv i_53834(.A(to_acu1[25]), .Z(n_40225));
	notech_inv i_53835(.A(n_3196), .Z(n_40226));
	notech_inv i_53836(.A(to_acu1[26]), .Z(n_40227));
	notech_inv i_53837(.A(n_3195), .Z(n_40228));
	notech_inv i_53838(.A(to_acu1[27]), .Z(n_40229));
	notech_inv i_53839(.A(n_3194), .Z(n_40230));
	notech_inv i_53840(.A(to_acu1[28]), .Z(n_40231));
	notech_inv i_53841(.A(n_3193), .Z(n_40232));
	notech_inv i_53842(.A(to_acu1[29]), .Z(n_40233));
	notech_inv i_53843(.A(n_3192), .Z(n_40234));
	notech_inv i_53844(.A(to_acu1[30]), .Z(n_40235));
	notech_inv i_53845(.A(n_3191), .Z(n_40236));
	notech_inv i_53846(.A(to_acu1[31]), .Z(n_40237));
	notech_inv i_53847(.A(n_3190), .Z(n_40238));
	notech_inv i_53848(.A(to_acu1[32]), .Z(n_40239));
	notech_inv i_53849(.A(n_3189), .Z(n_40240));
	notech_inv i_53850(.A(to_acu1[33]), .Z(n_40241));
	notech_inv i_53851(.A(n_3188), .Z(n_40242));
	notech_inv i_53852(.A(to_acu1[34]), .Z(n_40243));
	notech_inv i_53853(.A(n_3187), .Z(n_40244));
	notech_inv i_53854(.A(to_acu1[35]), .Z(n_40245));
	notech_inv i_53855(.A(n_3186), .Z(n_40246));
	notech_inv i_53856(.A(to_acu1[36]), .Z(n_40247));
	notech_inv i_53857(.A(to_acu1[37]), .Z(n_40248));
	notech_inv i_53858(.A(to_acu1[38]), .Z(n_40249));
	notech_inv i_53859(.A(to_acu1[40]), .Z(n_40250));
	notech_inv i_53860(.A(to_acu1[41]), .Z(n_40251));
	notech_inv i_53861(.A(to_acu1[42]), .Z(n_40252));
	notech_inv i_53862(.A(to_acu1[43]), .Z(n_40253));
	notech_inv i_53863(.A(to_acu1[44]), .Z(n_40254));
	notech_inv i_53864(.A(to_acu1[45]), .Z(n_40255));
	notech_inv i_53865(.A(to_acu1[46]), .Z(n_40256));
	notech_inv i_53866(.A(to_acu1[47]), .Z(n_40257));
	notech_inv i_53867(.A(to_acu1[48]), .Z(n_40258));
	notech_inv i_53868(.A(to_acu1[49]), .Z(n_40259));
	notech_inv i_53869(.A(to_acu1[50]), .Z(n_40260));
	notech_inv i_53870(.A(to_acu1[51]), .Z(n_40261));
	notech_inv i_53871(.A(to_acu1[52]), .Z(n_40262));
	notech_inv i_53872(.A(to_acu1[53]), .Z(n_40263));
	notech_inv i_53873(.A(to_acu1[54]), .Z(n_40264));
	notech_inv i_53874(.A(to_acu1[55]), .Z(n_40265));
	notech_inv i_53875(.A(to_acu1[56]), .Z(n_40266));
	notech_inv i_53876(.A(n_2898), .Z(n_40267));
	notech_inv i_53877(.A(to_acu1[57]), .Z(n_40268));
	notech_inv i_53878(.A(to_acu1[58]), .Z(n_40269));
	notech_inv i_53879(.A(to_acu1[59]), .Z(n_40270));
	notech_inv i_53880(.A(to_acu1[60]), .Z(n_40271));
	notech_inv i_53881(.A(to_acu1[61]), .Z(n_40272));
	notech_inv i_53882(.A(to_acu1[62]), .Z(n_40273));
	notech_inv i_53883(.A(to_acu1[63]), .Z(n_40274));
	notech_inv i_53884(.A(to_acu1[64]), .Z(n_40275));
	notech_inv i_53885(.A(to_acu1[65]), .Z(n_40276));
	notech_inv i_53886(.A(to_acu1[66]), .Z(n_40277));
	notech_inv i_53887(.A(to_acu1[67]), .Z(n_40278));
	notech_inv i_53888(.A(n_3149), .Z(n_40279));
	notech_inv i_53889(.A(to_acu1[68]), .Z(n_40280));
	notech_inv i_53890(.A(n_3148), .Z(n_40281));
	notech_inv i_53891(.A(to_acu1[69]), .Z(n_40282));
	notech_inv i_53892(.A(to_acu1[70]), .Z(n_40283));
	notech_inv i_53893(.A(to_acu1[71]), .Z(n_40284));
	notech_inv i_53894(.A(to_acu1[72]), .Z(n_40285));
	notech_inv i_53895(.A(to_acu1[73]), .Z(n_40286));
	notech_inv i_53896(.A(to_acu1[74]), .Z(n_40287));
	notech_inv i_53897(.A(to_acu1[75]), .Z(n_40288));
	notech_inv i_53898(.A(to_acu1[76]), .Z(n_40289));
	notech_inv i_53899(.A(n_3134), .Z(n_40290));
	notech_inv i_53900(.A(to_acu1[77]), .Z(n_40291));
	notech_inv i_53901(.A(to_acu1[78]), .Z(n_40292));
	notech_inv i_53902(.A(n_3133), .Z(n_40293));
	notech_inv i_53903(.A(to_acu1[79]), .Z(n_40294));
	notech_inv i_53904(.A(n_3132), .Z(n_40295));
	notech_inv i_53905(.A(to_acu1[80]), .Z(n_40296));
	notech_inv i_53906(.A(to_acu1[81]), .Z(n_40297));
	notech_inv i_53907(.A(n_3131), .Z(n_40298));
	notech_inv i_53908(.A(to_acu1[82]), .Z(n_40299));
	notech_inv i_53909(.A(n_3130), .Z(n_40300));
	notech_inv i_53910(.A(to_acu1[83]), .Z(n_40301));
	notech_inv i_53911(.A(n_48945), .Z(n_40302));
	notech_inv i_53912(.A(to_acu1[84]), .Z(n_40303));
	notech_inv i_53913(.A(n_3129), .Z(n_40304));
	notech_inv i_53914(.A(to_acu1[85]), .Z(n_40305));
	notech_inv i_53915(.A(to_acu1[86]), .Z(n_40306));
	notech_inv i_53916(.A(n_3128), .Z(n_40307));
	notech_inv i_53917(.A(to_acu1[87]), .Z(n_40308));
	notech_inv i_53918(.A(n_3127), .Z(n_40309));
	notech_inv i_53919(.A(to_acu1[88]), .Z(n_40310));
	notech_inv i_53920(.A(to_acu1[89]), .Z(n_40311));
	notech_inv i_53921(.A(n_3126), .Z(n_40312));
	notech_inv i_53922(.A(n_48981), .Z(n_40313));
	notech_inv i_53923(.A(to_acu1[90]), .Z(n_40314));
	notech_inv i_53924(.A(n_48987), .Z(n_40315));
	notech_inv i_53925(.A(to_acu1[91]), .Z(n_40316));
	notech_inv i_53926(.A(n_48993), .Z(n_40317));
	notech_inv i_53927(.A(to_acu1[92]), .Z(n_40318));
	notech_inv i_53928(.A(n_3125), .Z(n_40319));
	notech_inv i_53929(.A(n_48999), .Z(n_40320));
	notech_inv i_53930(.A(to_acu1[93]), .Z(n_40321));
	notech_inv i_53931(.A(n_49005), .Z(n_40322));
	notech_inv i_53932(.A(to_acu1[94]), .Z(n_40323));
	notech_inv i_53933(.A(n_49011), .Z(n_40324));
	notech_inv i_53934(.A(to_acu1[95]), .Z(n_40325));
	notech_inv i_53935(.A(n_3124), .Z(n_40326));
	notech_inv i_53936(.A(n_49017), .Z(n_40327));
	notech_inv i_53937(.A(to_acu1[96]), .Z(n_40328));
	notech_inv i_53938(.A(n_49023), .Z(n_40329));
	notech_inv i_53939(.A(to_acu1[97]), .Z(n_40330));
	notech_inv i_53940(.A(n_49029), .Z(n_40331));
	notech_inv i_53941(.A(to_acu1[98]), .Z(n_40332));
	notech_inv i_53942(.A(n_49035), .Z(n_40333));
	notech_inv i_53943(.A(to_acu1[99]), .Z(n_40334));
	notech_inv i_53944(.A(n_49041), .Z(n_40335));
	notech_inv i_53945(.A(to_acu1[100]), .Z(n_40336));
	notech_inv i_53946(.A(n_49047), .Z(n_40337));
	notech_inv i_53947(.A(to_acu1[101]), .Z(n_40338));
	notech_inv i_53948(.A(n_49053), .Z(n_40339));
	notech_inv i_53949(.A(to_acu1[102]), .Z(n_40340));
	notech_inv i_53950(.A(n_49059), .Z(n_40341));
	notech_inv i_53951(.A(to_acu1[103]), .Z(n_40342));
	notech_inv i_53952(.A(n_49065), .Z(n_40343));
	notech_inv i_53953(.A(to_acu1[104]), .Z(n_40344));
	notech_inv i_53954(.A(n_49071), .Z(n_40345));
	notech_inv i_53955(.A(to_acu1[105]), .Z(n_40346));
	notech_inv i_53956(.A(n_49077), .Z(n_40347));
	notech_inv i_53957(.A(to_acu1[106]), .Z(n_40348));
	notech_inv i_53958(.A(to_acu1[107]), .Z(n_40349));
	notech_inv i_53959(.A(n_49089), .Z(n_40350));
	notech_inv i_53960(.A(to_acu1[108]), .Z(n_40351));
	notech_inv i_53961(.A(to_acu1[109]), .Z(n_40352));
	notech_inv i_53962(.A(to_acu1[110]), .Z(n_40353));
	notech_inv i_53963(.A(to_acu1[111]), .Z(n_40354));
	notech_inv i_53964(.A(to_acu1[112]), .Z(n_40355));
	notech_inv i_53965(.A(to_acu1[113]), .Z(n_40356));
	notech_inv i_53966(.A(n_49125), .Z(n_40357));
	notech_inv i_53967(.A(to_acu1[114]), .Z(n_40358));
	notech_inv i_53968(.A(n_49131), .Z(n_40359));
	notech_inv i_53969(.A(to_acu1[115]), .Z(n_40360));
	notech_inv i_53970(.A(n_49137), .Z(n_40361));
	notech_inv i_53971(.A(to_acu1[116]), .Z(n_40362));
	notech_inv i_53972(.A(n_49143), .Z(n_40363));
	notech_inv i_53973(.A(to_acu1[117]), .Z(n_40364));
	notech_inv i_53974(.A(n_49149), .Z(n_40365));
	notech_inv i_53975(.A(to_acu1[118]), .Z(n_40366));
	notech_inv i_53976(.A(to_acu1[119]), .Z(n_40367));
	notech_inv i_53977(.A(n_49161), .Z(n_40368));
	notech_inv i_53978(.A(to_acu1[120]), .Z(n_40369));
	notech_inv i_53979(.A(to_acu1[121]), .Z(n_40370));
	notech_inv i_53980(.A(to_acu1[122]), .Z(n_40371));
	notech_inv i_53981(.A(to_acu1[123]), .Z(n_40372));
	notech_inv i_53982(.A(n_49185), .Z(n_40373));
	notech_inv i_53983(.A(to_acu1[124]), .Z(n_40374));
	notech_inv i_53984(.A(to_acu1[125]), .Z(n_40375));
	notech_inv i_53985(.A(to_acu1[126]), .Z(n_40376));
	notech_inv i_53986(.A(to_acu1[127]), .Z(n_40377));
	notech_inv i_53987(.A(to_acu1[128]), .Z(n_40378));
	notech_inv i_53988(.A(to_acu1[129]), .Z(n_40379));
	notech_inv i_53989(.A(to_acu1[130]), .Z(n_40380));
	notech_inv i_53990(.A(to_acu1[131]), .Z(n_40381));
	notech_inv i_53991(.A(to_acu1[132]), .Z(n_40382));
	notech_inv i_53992(.A(to_acu1[133]), .Z(n_40383));
	notech_inv i_53993(.A(to_acu1[134]), .Z(n_40384));
	notech_inv i_53994(.A(to_acu1[135]), .Z(n_40385));
	notech_inv i_53995(.A(to_acu1[136]), .Z(n_40386));
	notech_inv i_53996(.A(to_acu1[137]), .Z(n_40387));
	notech_inv i_53997(.A(to_acu1[138]), .Z(n_40388));
	notech_inv i_53998(.A(to_acu1[139]), .Z(n_40389));
	notech_inv i_53999(.A(to_acu1[140]), .Z(n_40390));
	notech_inv i_54000(.A(to_acu1[141]), .Z(n_40391));
	notech_inv i_54001(.A(to_acu1[142]), .Z(n_40392));
	notech_inv i_54002(.A(to_acu1[143]), .Z(n_40393));
	notech_inv i_54003(.A(to_acu1[144]), .Z(n_40394));
	notech_inv i_54004(.A(to_acu1[145]), .Z(n_40395));
	notech_inv i_54005(.A(to_acu1[146]), .Z(n_40396));
	notech_inv i_54006(.A(to_acu1[147]), .Z(n_40397));
	notech_inv i_54007(.A(to_acu1[148]), .Z(n_40398));
	notech_inv i_54008(.A(to_acu1[149]), .Z(n_40399));
	notech_inv i_54009(.A(n_49341), .Z(n_40400));
	notech_inv i_54010(.A(to_acu1[150]), .Z(n_40401));
	notech_inv i_54011(.A(n_49347), .Z(n_40402));
	notech_inv i_54012(.A(to_acu1[151]), .Z(n_40403));
	notech_inv i_54013(.A(n_49353), .Z(n_40404));
	notech_inv i_54014(.A(to_acu1[152]), .Z(n_40405));
	notech_inv i_54015(.A(to_acu1[153]), .Z(n_40406));
	notech_inv i_54016(.A(to_acu1[154]), .Z(n_40407));
	notech_inv i_54017(.A(to_acu1[155]), .Z(n_40408));
	notech_inv i_54018(.A(n_49377), .Z(n_40409));
	notech_inv i_54019(.A(to_acu1[156]), .Z(n_40410));
	notech_inv i_54020(.A(to_acu1[157]), .Z(n_40411));
	notech_inv i_54021(.A(to_acu1[158]), .Z(n_40412));
	notech_inv i_54022(.A(to_acu1[159]), .Z(n_40413));
	notech_inv i_54023(.A(to_acu1[160]), .Z(n_40414));
	notech_inv i_54024(.A(to_acu1[161]), .Z(n_40415));
	notech_inv i_54025(.A(to_acu1[162]), .Z(n_40416));
	notech_inv i_54026(.A(n_49419), .Z(n_40417));
	notech_inv i_54027(.A(to_acu1[163]), .Z(n_40418));
	notech_inv i_54028(.A(n_49425), .Z(n_40419));
	notech_inv i_54029(.A(to_acu1[164]), .Z(n_40420));
	notech_inv i_54030(.A(to_acu1[165]), .Z(n_40421));
	notech_inv i_54031(.A(to_acu1[166]), .Z(n_40422));
	notech_inv i_54032(.A(to_acu1[167]), .Z(n_40423));
	notech_inv i_54033(.A(to_acu1[168]), .Z(n_40424));
	notech_inv i_54034(.A(to_acu1[169]), .Z(n_40425));
	notech_inv i_54035(.A(to_acu1[170]), .Z(n_40426));
	notech_inv i_54036(.A(to_acu1[171]), .Z(n_40427));
	notech_inv i_54037(.A(to_acu1[172]), .Z(n_40428));
	notech_inv i_54038(.A(to_acu1[173]), .Z(n_40429));
	notech_inv i_54039(.A(to_acu1[174]), .Z(n_40430));
	notech_inv i_54040(.A(to_acu1[175]), .Z(n_40431));
	notech_inv i_54041(.A(to_acu1[176]), .Z(n_40432));
	notech_inv i_54042(.A(to_acu1[177]), .Z(n_40433));
	notech_inv i_54043(.A(to_acu1[178]), .Z(n_40434));
	notech_inv i_54044(.A(to_acu1[179]), .Z(n_40435));
	notech_inv i_54045(.A(to_acu1[180]), .Z(n_40436));
	notech_inv i_54046(.A(to_acu1[181]), .Z(n_40437));
	notech_inv i_54047(.A(to_acu1[182]), .Z(n_40438));
	notech_inv i_54048(.A(to_acu1[183]), .Z(n_40439));
	notech_inv i_54049(.A(to_acu1[184]), .Z(n_40440));
	notech_inv i_54050(.A(to_acu1[185]), .Z(n_40441));
	notech_inv i_54051(.A(to_acu1[186]), .Z(n_40442));
	notech_inv i_54052(.A(to_acu1[187]), .Z(n_40443));
	notech_inv i_54053(.A(to_acu1[188]), .Z(n_40444));
	notech_inv i_54054(.A(to_acu1[189]), .Z(n_40445));
	notech_inv i_54055(.A(to_acu1[190]), .Z(n_40446));
	notech_inv i_54056(.A(to_acu1[191]), .Z(n_40447));
	notech_inv i_54057(.A(to_acu1[192]), .Z(n_40448));
	notech_inv i_54058(.A(to_acu1[193]), .Z(n_40449));
	notech_inv i_54059(.A(to_acu1[194]), .Z(n_40450));
	notech_inv i_54060(.A(n_49611), .Z(n_40451));
	notech_inv i_54061(.A(to_acu1[195]), .Z(n_40452));
	notech_inv i_54062(.A(to_acu1[196]), .Z(n_40453));
	notech_inv i_54063(.A(to_acu1[197]), .Z(n_40454));
	notech_inv i_54064(.A(to_acu1[198]), .Z(n_40455));
	notech_inv i_54065(.A(to_acu1[199]), .Z(n_40456));
	notech_inv i_54066(.A(to_acu1[200]), .Z(n_40457));
	notech_inv i_54067(.A(to_acu1[201]), .Z(n_40458));
	notech_inv i_54068(.A(to_acu1[202]), .Z(n_40459));
	notech_inv i_54069(.A(to_acu1[203]), .Z(n_40460));
	notech_inv i_54070(.A(to_acu1[204]), .Z(n_40461));
	notech_inv i_54071(.A(to_acu1[205]), .Z(n_40462));
	notech_inv i_54072(.A(to_acu1[206]), .Z(n_40463));
	notech_inv i_54073(.A(to_acu1[207]), .Z(n_40464));
	notech_inv i_54074(.A(to_acu1[208]), .Z(n_40465));
	notech_inv i_54075(.A(to_acu1[209]), .Z(n_40466));
	notech_inv i_54076(.A(to_acu1[210]), .Z(n_40467));
	notech_inv i_54077(.A(n_41563), .Z(n_40468));
	notech_inv i_54078(.A(overgs), .Z(n_40469));
	notech_inv i_54079(.A(\over_seg2[5] ), .Z(n_40470));
	notech_inv i_54080(.A(n_43160), .Z(n_40471));
	notech_inv i_54081(.A(\over_seg1[5] ), .Z(n_40472));
	notech_inv i_54082(.A(lenpc1[0]), .Z(n_40473));
	notech_inv i_54083(.A(lenpc1[1]), .Z(n_40474));
	notech_inv i_54084(.A(lenpc1[2]), .Z(n_40475));
	notech_inv i_54085(.A(lenpc1[3]), .Z(n_40476));
	notech_inv i_54086(.A(lenpc1[4]), .Z(n_40477));
	notech_inv i_54087(.A(lenpc1[5]), .Z(n_40478));
	notech_inv i_54088(.A(n_2933), .Z(n_40479));
	notech_inv i_54089(.A(n_46406), .Z(n_40480));
	notech_inv i_54090(.A(n_46412), .Z(n_40481));
	notech_inv i_54091(.A(n_46418), .Z(n_40482));
	notech_inv i_54092(.A(n_46424), .Z(n_40483));
	notech_inv i_54093(.A(n_46430), .Z(n_40484));
	notech_inv i_54094(.A(n_46436), .Z(n_40485));
	notech_inv i_54095(.A(n_227396436), .Z(n_40486));
	notech_inv i_54096(.A(n_2935), .Z(n_40487));
	notech_inv i_54097(.A(n_2949), .Z(n_40488));
	notech_inv i_54098(.A(n_2947), .Z(n_40489));
	notech_inv i_54099(.A(n_2942), .Z(n_40490));
	notech_inv i_54100(.A(n_2941), .Z(n_40491));
	notech_inv i_54101(.A(n_2940), .Z(n_40492));
	notech_inv i_54102(.A(n_2931), .Z(n_40493));
	notech_inv i_54103(.A(opz2[0]), .Z(n_40494));
	notech_inv i_54104(.A(opz2[1]), .Z(n_40495));
	notech_inv i_54105(.A(opz1[0]), .Z(n_40496));
	notech_inv i_54106(.A(opz1[1]), .Z(n_40497));
	notech_inv i_54107(.A(n_223996470), .Z(n_40498));
	notech_inv i_54108(.A(n_2905), .Z(n_40499));
	notech_inv i_54109(.A(n_2223), .Z(n_40500));
	notech_inv i_54110(.A(n_2887), .Z(n_40501));
	notech_inv i_54111(.A(n_2885), .Z(n_40502));
	notech_inv i_54112(.A(n_2880), .Z(n_40503));
	notech_inv i_54113(.A(n_2878), .Z(n_40504));
	notech_inv i_54114(.A(n_2874), .Z(n_40505));
	notech_inv i_54115(.A(n_2873), .Z(n_40506));
	notech_inv i_54116(.A(n_41603), .Z(n_40507));
	notech_inv i_54117(.A(n_41633), .Z(n_40508));
	notech_inv i_54118(.A(n_41657), .Z(n_40509));
	notech_inv i_54119(.A(n_41669), .Z(n_40510));
	notech_inv i_54120(.A(n_41675), .Z(n_40511));
	notech_inv i_54121(.A(n_41681), .Z(n_40512));
	notech_inv i_54122(.A(n_41687), .Z(n_40513));
	notech_inv i_54123(.A(n_41693), .Z(n_40514));
	notech_inv i_54124(.A(n_41711), .Z(n_40515));
	notech_inv i_54125(.A(n_41729), .Z(n_40516));
	notech_inv i_54126(.A(n_41735), .Z(n_40517));
	notech_inv i_54127(.A(n_41861), .Z(n_40518));
	notech_inv i_54128(.A(n_41867), .Z(n_40519));
	notech_inv i_54129(.A(n_254394500), .Z(n_40520));
	notech_inv i_54130(.A(n_41891), .Z(n_40521));
	notech_inv i_54131(.A(n_41897), .Z(n_40522));
	notech_inv i_54132(.A(n_41915), .Z(n_40523));
	notech_inv i_54133(.A(n_41933), .Z(n_40524));
	notech_inv i_54134(.A(n_41939), .Z(n_40525));
	notech_inv i_54135(.A(n_41945), .Z(n_40526));
	notech_inv i_54136(.A(n_41957), .Z(n_40527));
	notech_inv i_54137(.A(n_41963), .Z(n_40528));
	notech_inv i_54138(.A(n_41969), .Z(n_40529));
	notech_inv i_54139(.A(n_41981), .Z(n_40530));
	notech_inv i_54140(.A(n_41987), .Z(n_40531));
	notech_inv i_54141(.A(n_41993), .Z(n_40532));
	notech_inv i_54142(.A(n_41999), .Z(n_40533));
	notech_inv i_54143(.A(n_240094357), .Z(n_40534));
	notech_inv i_54144(.A(n_42005), .Z(n_40535));
	notech_inv i_54145(.A(n_42011), .Z(n_40536));
	notech_inv i_54146(.A(n_42017), .Z(n_40537));
	notech_inv i_54147(.A(n_42023), .Z(n_40538));
	notech_inv i_54148(.A(n_42029), .Z(n_40539));
	notech_inv i_54149(.A(n_42035), .Z(n_40540));
	notech_inv i_54150(.A(n_42041), .Z(n_40541));
	notech_inv i_54151(.A(n_42047), .Z(n_40542));
	notech_inv i_54152(.A(n_42053), .Z(n_40543));
	notech_inv i_54153(.A(n_42059), .Z(n_40544));
	notech_inv i_54154(.A(n_42065), .Z(n_40545));
	notech_inv i_54155(.A(n_42071), .Z(n_40546));
	notech_inv i_54156(.A(n_42077), .Z(n_40547));
	notech_inv i_54157(.A(n_42083), .Z(n_40548));
	notech_inv i_54158(.A(n_42089), .Z(n_40549));
	notech_inv i_54159(.A(n_42095), .Z(n_40550));
	notech_inv i_54160(.A(n_42101), .Z(n_40551));
	notech_inv i_54161(.A(n_42107), .Z(n_40552));
	notech_inv i_54162(.A(n_42113), .Z(n_40553));
	notech_inv i_54163(.A(n_42119), .Z(n_40554));
	notech_inv i_54164(.A(n_42125), .Z(n_40555));
	notech_inv i_54165(.A(n_42131), .Z(n_40556));
	notech_inv i_54166(.A(n_42137), .Z(n_40557));
	notech_inv i_54167(.A(n_42149), .Z(n_40558));
	notech_inv i_54168(.A(n_2222), .Z(n_40559));
	notech_inv i_54169(.A(n_42161), .Z(n_40560));
	notech_inv i_54170(.A(n_42335), .Z(n_40561));
	notech_inv i_54171(.A(n_42341), .Z(n_40562));
	notech_inv i_54172(.A(n_42353), .Z(n_40563));
	notech_inv i_54173(.A(n_42359), .Z(n_40564));
	notech_inv i_54174(.A(n_42365), .Z(n_40565));
	notech_inv i_54175(.A(n_42371), .Z(n_40566));
	notech_inv i_54176(.A(n_42377), .Z(n_40567));
	notech_inv i_54177(.A(n_42443), .Z(n_40568));
	notech_inv i_54178(.A(n_42455), .Z(n_40569));
	notech_inv i_54179(.A(n_42461), .Z(n_40570));
	notech_inv i_54180(.A(n_42467), .Z(n_40571));
	notech_inv i_54181(.A(n_42491), .Z(n_40572));
	notech_inv i_54182(.A(n_42497), .Z(n_40573));
	notech_inv i_54183(.A(n_42527), .Z(n_40574));
	notech_inv i_54184(.A(n_42533), .Z(n_40575));
	notech_inv i_54185(.A(n_42545), .Z(n_40576));
	notech_inv i_54186(.A(n_42557), .Z(n_40577));
	notech_inv i_54187(.A(n_42563), .Z(n_40578));
	notech_inv i_54188(.A(n_42569), .Z(n_40579));
	notech_inv i_54189(.A(n_42611), .Z(n_40580));
	notech_inv i_54190(.A(n_42797), .Z(n_40581));
	notech_inv i_54191(.A(n_42809), .Z(n_40582));
	notech_inv i_54192(.A(n_42815), .Z(n_40583));
	notech_inv i_54193(.A(n_42821), .Z(n_40584));
	notech_inv i_54194(.A(n_42827), .Z(n_40585));
	notech_inv i_54195(.A(n_42839), .Z(n_40586));
	notech_inv i_54196(.A(n_42851), .Z(n_40587));
	notech_inv i_54197(.A(n_42857), .Z(n_40588));
	notech_inv i_54198(.A(n_1517), .Z(n_40589));
	notech_inv i_54199(.A(n_42863), .Z(n_40590));
	notech_inv i_54200(.A(imm_sz[0]), .Z(n_40591));
	notech_inv i_54201(.A(imm_sz[1]), .Z(n_40592));
	notech_inv i_54202(.A(imm_sz[2]), .Z(n_40593));
	notech_inv i_54203(.A(displc[0]), .Z(n_40594));
	notech_inv i_54204(.A(udeco[0]), .Z(n_40595));
	notech_inv i_54205(.A(udeco[1]), .Z(n_40596));
	notech_inv i_54206(.A(udeco[2]), .Z(n_40597));
	notech_inv i_54207(.A(udeco[3]), .Z(n_40598));
	notech_inv i_54208(.A(udeco[4]), .Z(n_40599));
	notech_inv i_54209(.A(udeco[5]), .Z(n_40600));
	notech_inv i_54210(.A(udeco[6]), .Z(n_40601));
	notech_inv i_54211(.A(udeco[7]), .Z(n_40602));
	notech_inv i_54212(.A(udeco[8]), .Z(n_40603));
	notech_inv i_54213(.A(udeco[9]), .Z(n_40604));
	notech_inv i_54214(.A(udeco[10]), .Z(n_40605));
	notech_inv i_54215(.A(udeco[11]), .Z(n_40606));
	notech_inv i_54216(.A(udeco[12]), .Z(n_40607));
	notech_inv i_54217(.A(udeco[13]), .Z(n_40608));
	notech_inv i_54218(.A(udeco[14]), .Z(n_40609));
	notech_inv i_54219(.A(udeco[15]), .Z(n_40610));
	notech_inv i_54220(.A(udeco[16]), .Z(n_40611));
	notech_inv i_54221(.A(udeco[17]), .Z(n_40612));
	notech_inv i_54222(.A(udeco[18]), .Z(n_40613));
	notech_inv i_54223(.A(udeco[19]), .Z(n_40614));
	notech_inv i_54224(.A(udeco[20]), .Z(n_40615));
	notech_inv i_54225(.A(udeco[21]), .Z(n_40616));
	notech_inv i_54226(.A(udeco[22]), .Z(n_40617));
	notech_inv i_54227(.A(udeco[23]), .Z(n_40618));
	notech_inv i_54228(.A(udeco[24]), .Z(n_40619));
	notech_inv i_54229(.A(udeco[25]), .Z(n_40620));
	notech_inv i_54230(.A(udeco[26]), .Z(n_40621));
	notech_inv i_54231(.A(udeco[27]), .Z(n_40622));
	notech_inv i_54232(.A(udeco[28]), .Z(n_40623));
	notech_inv i_54233(.A(udeco[29]), .Z(n_40624));
	notech_inv i_54234(.A(udeco[30]), .Z(n_40625));
	notech_inv i_54235(.A(udeco[31]), .Z(n_40626));
	notech_inv i_54236(.A(udeco[32]), .Z(n_40627));
	notech_inv i_54237(.A(udeco[33]), .Z(n_40628));
	notech_inv i_54238(.A(udeco[34]), .Z(n_40629));
	notech_inv i_54239(.A(udeco[35]), .Z(n_40630));
	notech_inv i_54240(.A(udeco[36]), .Z(n_40631));
	notech_inv i_54241(.A(udeco[37]), .Z(n_40632));
	notech_inv i_54242(.A(udeco[38]), .Z(n_40633));
	notech_inv i_54243(.A(udeco[39]), .Z(n_40634));
	notech_inv i_54244(.A(udeco[40]), .Z(n_40635));
	notech_inv i_54245(.A(udeco[41]), .Z(n_40636));
	notech_inv i_54246(.A(udeco[42]), .Z(n_40637));
	notech_inv i_54247(.A(udeco[43]), .Z(n_40638));
	notech_inv i_54248(.A(udeco[44]), .Z(n_40639));
	notech_inv i_54249(.A(udeco[45]), .Z(n_40640));
	notech_inv i_54250(.A(udeco[46]), .Z(n_40641));
	notech_inv i_54251(.A(udeco[47]), .Z(n_40642));
	notech_inv i_54252(.A(udeco[48]), .Z(n_40643));
	notech_inv i_54253(.A(udeco[49]), .Z(n_40644));
	notech_inv i_54254(.A(udeco[50]), .Z(n_40645));
	notech_inv i_54255(.A(udeco[51]), .Z(n_40646));
	notech_inv i_54256(.A(udeco[52]), .Z(n_40647));
	notech_inv i_54257(.A(udeco[53]), .Z(n_40648));
	notech_inv i_54258(.A(udeco[54]), .Z(n_40649));
	notech_inv i_54259(.A(udeco[55]), .Z(n_40650));
	notech_inv i_54260(.A(udeco[56]), .Z(n_40651));
	notech_inv i_54261(.A(udeco[57]), .Z(n_40652));
	notech_inv i_54262(.A(udeco[58]), .Z(n_40653));
	notech_inv i_54263(.A(udeco[59]), .Z(n_40654));
	notech_inv i_54264(.A(udeco[60]), .Z(n_40655));
	notech_inv i_54265(.A(udeco[61]), .Z(n_40656));
	notech_inv i_54266(.A(udeco[62]), .Z(n_40657));
	notech_inv i_54267(.A(udeco[63]), .Z(n_40658));
	notech_inv i_54268(.A(udeco[64]), .Z(n_40659));
	notech_inv i_54269(.A(udeco[65]), .Z(n_40660));
	notech_inv i_54270(.A(udeco[66]), .Z(n_40661));
	notech_inv i_54271(.A(udeco[67]), .Z(n_40662));
	notech_inv i_54272(.A(udeco[68]), .Z(n_40663));
	notech_inv i_54273(.A(udeco[69]), .Z(n_40664));
	notech_inv i_54274(.A(udeco[70]), .Z(n_40665));
	notech_inv i_54275(.A(udeco[71]), .Z(n_40666));
	notech_inv i_54276(.A(udeco[72]), .Z(n_40667));
	notech_inv i_54277(.A(udeco[73]), .Z(n_40668));
	notech_inv i_54278(.A(udeco[74]), .Z(n_40669));
	notech_inv i_54279(.A(udeco[75]), .Z(n_40670));
	notech_inv i_54280(.A(udeco[76]), .Z(n_40671));
	notech_inv i_54281(.A(udeco[77]), .Z(n_40672));
	notech_inv i_54282(.A(udeco[78]), .Z(n_40673));
	notech_inv i_54283(.A(udeco[79]), .Z(n_40674));
	notech_inv i_54284(.A(udeco[80]), .Z(n_40675));
	notech_inv i_54285(.A(udeco[81]), .Z(n_40676));
	notech_inv i_54286(.A(udeco[82]), .Z(n_40677));
	notech_inv i_54287(.A(udeco[83]), .Z(n_40678));
	notech_inv i_54288(.A(udeco[84]), .Z(n_40679));
	notech_inv i_54289(.A(udeco[85]), .Z(n_40680));
	notech_inv i_54290(.A(udeco[86]), .Z(n_40681));
	notech_inv i_54291(.A(udeco[87]), .Z(n_40682));
	notech_inv i_54292(.A(udeco[88]), .Z(n_40683));
	notech_inv i_54293(.A(udeco[89]), .Z(n_40684));
	notech_inv i_54294(.A(udeco[90]), .Z(n_40685));
	notech_inv i_54295(.A(udeco[91]), .Z(n_40686));
	notech_inv i_54296(.A(udeco[92]), .Z(n_40687));
	notech_inv i_54297(.A(udeco[93]), .Z(n_40688));
	notech_inv i_54298(.A(udeco[94]), .Z(n_40689));
	notech_inv i_54299(.A(udeco[95]), .Z(n_40690));
	notech_inv i_54300(.A(udeco[96]), .Z(n_40691));
	notech_inv i_54301(.A(udeco[97]), .Z(n_40692));
	notech_inv i_54302(.A(udeco[98]), .Z(n_40693));
	notech_inv i_54303(.A(udeco[99]), .Z(n_40694));
	notech_inv i_54304(.A(udeco[100]), .Z(n_40695));
	notech_inv i_54305(.A(udeco[101]), .Z(n_40696));
	notech_inv i_54306(.A(udeco[102]), .Z(n_40697));
	notech_inv i_54307(.A(udeco[103]), .Z(n_40698));
	notech_inv i_54308(.A(udeco[104]), .Z(n_40699));
	notech_inv i_54309(.A(udeco[105]), .Z(n_40700));
	notech_inv i_54310(.A(udeco[106]), .Z(n_40701));
	notech_inv i_54311(.A(udeco[107]), .Z(n_40702));
	notech_inv i_54312(.A(udeco[108]), .Z(n_40703));
	notech_inv i_54313(.A(udeco[109]), .Z(n_40704));
	notech_inv i_54314(.A(udeco[110]), .Z(n_40705));
	notech_inv i_54315(.A(udeco[111]), .Z(n_40706));
	notech_inv i_54316(.A(udeco[112]), .Z(n_40707));
	notech_inv i_54317(.A(udeco[113]), .Z(n_40708));
	notech_inv i_54318(.A(udeco[114]), .Z(n_40709));
	notech_inv i_54319(.A(udeco[115]), .Z(n_40710));
	notech_inv i_54320(.A(udeco[116]), .Z(n_40711));
	notech_inv i_54321(.A(udeco[117]), .Z(n_40712));
	notech_inv i_54322(.A(udeco[118]), .Z(n_40713));
	notech_inv i_54323(.A(udeco[119]), .Z(n_40714));
	notech_inv i_54324(.A(udeco[120]), .Z(n_40715));
	notech_inv i_54325(.A(udeco[121]), .Z(n_40716));
	notech_inv i_54326(.A(udeco[122]), .Z(n_40717));
	notech_inv i_54327(.A(udeco[123]), .Z(n_40718));
	notech_inv i_54328(.A(udeco[124]), .Z(n_40719));
	notech_inv i_54329(.A(udeco[125]), .Z(n_40720));
	notech_inv i_54330(.A(udeco[126]), .Z(n_40721));
	notech_inv i_54331(.A(udeco[127]), .Z(n_40722));
	notech_inv i_54332(.A(valid_len[5]), .Z(n_40723));
	notech_inv i_54333(.A(pfx_sz[1]), .Z(n_40724));
	notech_inv i_54334(.A(opz[0]), .Z(n_40725));
	notech_inv i_54335(.A(opz[1]), .Z(n_40726));
	notech_inv i_54336(.A(in128[16]), .Z(n_40727));
	notech_inv i_54337(.A(in128[17]), .Z(n_40728));
	notech_inv i_54338(.A(in128[18]), .Z(n_40729));
	notech_inv i_54339(.A(in128[19]), .Z(n_40730));
	notech_inv i_54340(.A(in128[20]), .Z(n_40731));
	notech_inv i_54341(.A(in128[21]), .Z(n_40732));
	notech_inv i_54342(.A(in128[22]), .Z(n_40733));
	notech_inv i_54343(.A(in128[23]), .Z(n_40734));
	notech_inv i_54344(.A(in128[24]), .Z(n_40735));
	notech_inv i_54345(.A(in128[25]), .Z(n_40736));
	notech_inv i_54346(.A(in128[26]), .Z(n_40737));
	notech_inv i_54347(.A(in128[27]), .Z(n_40738));
	notech_inv i_54348(.A(in128[28]), .Z(n_40739));
	notech_inv i_54349(.A(in128[29]), .Z(n_40740));
	notech_inv i_54350(.A(in128[30]), .Z(n_40741));
	notech_inv i_54351(.A(in128[31]), .Z(n_40742));
	notech_inv i_54352(.A(in128[32]), .Z(n_40743));
	notech_inv i_54353(.A(in128[33]), .Z(n_40744));
	notech_inv i_54354(.A(in128[34]), .Z(n_40745));
	notech_inv i_54355(.A(in128[35]), .Z(n_40746));
	notech_inv i_54356(.A(in128[36]), .Z(n_40747));
	notech_inv i_54357(.A(in128[37]), .Z(n_40748));
	notech_inv i_54358(.A(in128[38]), .Z(n_40749));
	notech_inv i_54359(.A(in128[39]), .Z(n_40750));
	notech_inv i_54360(.A(in128[40]), .Z(n_40751));
	notech_inv i_54361(.A(in128[41]), .Z(n_40752));
	notech_inv i_54362(.A(in128[42]), .Z(n_40753));
	notech_inv i_54363(.A(in128[43]), .Z(n_40754));
	notech_inv i_54364(.A(in128[44]), .Z(n_40755));
	notech_inv i_54365(.A(in128[45]), .Z(n_40756));
	notech_inv i_54366(.A(in128[46]), .Z(n_40757));
	notech_inv i_54367(.A(in128[47]), .Z(n_40758));
	notech_inv i_54368(.A(in128[48]), .Z(n_40759));
	notech_inv i_54369(.A(in128[49]), .Z(n_40760));
	notech_inv i_54370(.A(in128[50]), .Z(n_40761));
	notech_inv i_54371(.A(in128[51]), .Z(n_40762));
	notech_inv i_54372(.A(in128[52]), .Z(n_40763));
	notech_inv i_54373(.A(in128[53]), .Z(n_40764));
	notech_inv i_54374(.A(in128[54]), .Z(n_40765));
	notech_inv i_54375(.A(in128[55]), .Z(n_40766));
	notech_inv i_54376(.A(in128[56]), .Z(n_40767));
	notech_inv i_54377(.A(in128[57]), .Z(n_40768));
	notech_inv i_54378(.A(in128[58]), .Z(n_40769));
	notech_inv i_54379(.A(in128[59]), .Z(n_40770));
	notech_inv i_54380(.A(in128[60]), .Z(n_40771));
	notech_inv i_54381(.A(in128[61]), .Z(n_40772));
	notech_inv i_54382(.A(in128[62]), .Z(n_40773));
	notech_inv i_54383(.A(in128[63]), .Z(n_40774));
	notech_inv i_54384(.A(in128[64]), .Z(n_40775));
	notech_inv i_54385(.A(in128[65]), .Z(n_40776));
	notech_inv i_54386(.A(in128[66]), .Z(n_40777));
	notech_inv i_54387(.A(in128[67]), .Z(n_40778));
	notech_inv i_54388(.A(in128[68]), .Z(n_40779));
	notech_inv i_54389(.A(in128[69]), .Z(n_40780));
	notech_inv i_54390(.A(in128[70]), .Z(n_40781));
	notech_inv i_54391(.A(in128[71]), .Z(n_40782));
	notech_inv i_54392(.A(in128[72]), .Z(n_40783));
	notech_inv i_54393(.A(in128[73]), .Z(n_40784));
	notech_inv i_54394(.A(in128[74]), .Z(n_40785));
	notech_inv i_54395(.A(in128[75]), .Z(n_40786));
	notech_inv i_54396(.A(in128[76]), .Z(n_40787));
	notech_inv i_54397(.A(in128[77]), .Z(n_40788));
	notech_inv i_54398(.A(in128[78]), .Z(n_40789));
	notech_inv i_54399(.A(in128[79]), .Z(n_40790));
	notech_inv i_54400(.A(in128[80]), .Z(n_40791));
	notech_inv i_54401(.A(in128[81]), .Z(n_40792));
	notech_inv i_54402(.A(in128[82]), .Z(n_40793));
	notech_inv i_54403(.A(in128[83]), .Z(n_40794));
	notech_inv i_54404(.A(in128[84]), .Z(n_40795));
	notech_inv i_54405(.A(in128[85]), .Z(n_40796));
	notech_inv i_54406(.A(in128[86]), .Z(n_40797));
	notech_inv i_54407(.A(in128[87]), .Z(n_40798));
	notech_inv i_54408(.A(in128[88]), .Z(n_40799));
	notech_inv i_54409(.A(in128[89]), .Z(n_40800));
	notech_inv i_54410(.A(in128[90]), .Z(n_40801));
	notech_inv i_54411(.A(in128[91]), .Z(n_40802));
	notech_inv i_54412(.A(in128[92]), .Z(n_40803));
	notech_inv i_54413(.A(in128[93]), .Z(n_40804));
	notech_inv i_54414(.A(in128[94]), .Z(n_40805));
	notech_inv i_54415(.A(in128[95]), .Z(n_40806));
	notech_inv i_54416(.A(in128[96]), .Z(n_40807));
	notech_inv i_54417(.A(in128[97]), .Z(n_40808));
	notech_inv i_54418(.A(in128[98]), .Z(n_40809));
	notech_inv i_54419(.A(in128[99]), .Z(n_40810));
	notech_inv i_54420(.A(in128[100]), .Z(n_40811));
	notech_inv i_54421(.A(in128[101]), .Z(n_40812));
	notech_inv i_54422(.A(in128[102]), .Z(n_40813));
	notech_inv i_54423(.A(in128[103]), .Z(n_40814));
	notech_inv i_54424(.A(in128[104]), .Z(n_40815));
	notech_inv i_54425(.A(in128[105]), .Z(n_40816));
	notech_inv i_54426(.A(in128[106]), .Z(n_40817));
	notech_inv i_54427(.A(in128[107]), .Z(n_40818));
	notech_inv i_54428(.A(in128[108]), .Z(n_40819));
	notech_inv i_54429(.A(in128[109]), .Z(n_40820));
	notech_inv i_54430(.A(in128[110]), .Z(n_40821));
	notech_inv i_54431(.A(in128[111]), .Z(n_40822));
	notech_inv i_54432(.A(in128[112]), .Z(n_40823));
	notech_inv i_54433(.A(in128[113]), .Z(n_40824));
	notech_inv i_54434(.A(in128[114]), .Z(n_40825));
	notech_inv i_54435(.A(in128[115]), .Z(n_40826));
	notech_inv i_54436(.A(in128[116]), .Z(n_40827));
	notech_inv i_54437(.A(in128[117]), .Z(n_40828));
	notech_inv i_54438(.A(in128[118]), .Z(n_40829));
	notech_inv i_54439(.A(in128[119]), .Z(n_40830));
	notech_inv i_54440(.A(in128[120]), .Z(n_40831));
	notech_inv i_54441(.A(in128[121]), .Z(n_40832));
	notech_inv i_54442(.A(in128[122]), .Z(n_40833));
	notech_inv i_54443(.A(in128[123]), .Z(n_40834));
	notech_inv i_54444(.A(in128[124]), .Z(n_40835));
	notech_inv i_54445(.A(in128[125]), .Z(n_40836));
	notech_inv i_54446(.A(in128[126]), .Z(n_40837));
	notech_inv i_54447(.A(in128[127]), .Z(n_40838));
	notech_inv i_54448(.A(in128[0]), .Z(n_40839));
	notech_inv i_54449(.A(\to_acu2_0[77] ), .Z(n_40840));
	notech_inv i_54450(.A(\to_acu2_0[67] ), .Z(n_40841));
	notech_inv i_54451(.A(\to_acu2_0[66] ), .Z(n_40842));
	notech_inv i_54452(.A(\to_acu2_0[65] ), .Z(n_40843));
	notech_inv i_54453(.A(\to_acu2_0[64] ), .Z(n_40844));
	notech_inv i_54454(.A(\to_acu2_0[63] ), .Z(n_40845));
	notech_inv i_54455(.A(\to_acu2_0[60] ), .Z(n_40846));
	notech_inv i_54456(.A(\to_acu2_0[49] ), .Z(n_40847));
	notech_inv i_54457(.A(\to_acu2_0[33] ), .Z(n_40848));
	notech_inv i_54458(.A(\to_acu2_0[32] ), .Z(n_40849));
	notech_inv i_54459(.A(\to_acu2_0[31] ), .Z(n_40850));
	notech_inv i_54460(.A(\to_acu2_0[30] ), .Z(n_40851));
	notech_inv i_54461(.A(\to_acu2_0[29] ), .Z(n_40852));
	notech_inv i_54462(.A(\to_acu2_0[71] ), .Z(n_40853));
	notech_inv i_54463(.A(\to_acu2_0[70] ), .Z(n_40854));
	notech_inv i_54464(.A(\to_acu2_0[75] ), .Z(n_40855));
	notech_inv i_54465(.A(in128[6]), .Z(n_40856));
	notech_inv i_54466(.A(in128[5]), .Z(n_40857));
	notech_inv i_54467(.A(in128[4]), .Z(n_40858));
	notech_inv i_54468(.A(in128[3]), .Z(n_40859));
	notech_inv i_54469(.A(\to_acu2_0[56] ), .Z(n_40860));
	notech_inv i_54470(.A(\to_acu2_0[50] ), .Z(n_40861));
	notech_inv i_54471(.A(\to_acu2_0[76] ), .Z(n_40862));
	notech_inv i_54472(.A(\to_acu2_0[72] ), .Z(n_40863));
	notech_inv i_54473(.A(\to_acu2_0[73] ), .Z(n_40864));
	notech_inv i_54474(.A(\to_acu2_0[74] ), .Z(n_40865));
	notech_inv i_54475(.A(\to_acu2_0[57] ), .Z(n_40866));
	notech_inv i_54476(.A(\to_acu2_0[52] ), .Z(n_40867));
	notech_inv i_54477(.A(\to_acu2_0[51] ), .Z(n_40868));
	notech_inv i_54478(.A(\to_acu2_0[53] ), .Z(n_40869));
	notech_inv i_54479(.A(\to_acu2_0[55] ), .Z(n_40870));
	notech_inv i_54480(.A(\to_acu2_0[54] ), .Z(n_40871));
	notech_inv i_54481(.A(\to_acu2_0[59] ), .Z(n_40872));
	notech_inv i_54482(.A(\to_acu2_0[80] ), .Z(n_40873));
	notech_inv i_54483(.A(\to_acu2_0[48] ), .Z(n_40874));
	notech_inv i_54484(.A(\to_acu2_0[5] ), .Z(n_40875));
	notech_inv i_54485(.A(\to_acu2_0[35] ), .Z(n_40876));
	notech_inv i_54486(.A(\to_acu2_0[34] ), .Z(n_40877));
	notech_inv i_54487(.A(\to_acu2_0[37] ), .Z(n_40878));
	notech_inv i_54488(.A(\to_acu2_0[36] ), .Z(n_40879));
	notech_inv i_54489(.A(\to_acu2_0[40] ), .Z(n_40880));
	notech_inv i_54490(.A(\to_acu2_0[38] ), .Z(n_40881));
	notech_inv i_54491(.A(\to_acu2_0[41] ), .Z(n_40882));
	notech_inv i_54492(.A(\to_acu2_0[43] ), .Z(n_40883));
	notech_inv i_54493(.A(\to_acu2_0[42] ), .Z(n_40884));
	notech_inv i_54494(.A(\to_acu2_0[44] ), .Z(n_40885));
	notech_inv i_54495(.A(\to_acu2_0[46] ), .Z(n_40886));
	notech_inv i_54496(.A(\to_acu2_0[45] ), .Z(n_40887));
	notech_inv i_54497(.A(\to_acu2_0[47] ), .Z(n_40888));
	notech_inv i_54498(.A(\to_acu2_0[79] ), .Z(n_40889));
	notech_inv i_54499(.A(\to_acu2_0[61] ), .Z(n_40890));
	notech_inv i_54500(.A(\to_acu2_0[78] ), .Z(n_40891));
	notech_inv i_54501(.A(in128[15]), .Z(n_40892));
	notech_inv i_54502(.A(in128[14]), .Z(n_40893));
	notech_inv i_54503(.A(in128[8]), .Z(n_40894));
	notech_inv i_54504(.A(\to_acu2_0[15] ), .Z(n_40895));
	notech_inv i_54505(.A(\to_acu2_0[14] ), .Z(n_40896));
	notech_inv i_54506(.A(\to_acu2_0[13] ), .Z(n_40897));
	notech_inv i_54507(.A(\to_acu2_0[17] ), .Z(n_40898));
	notech_inv i_54508(.A(\to_acu2_0[18] ), .Z(n_40899));
	notech_inv i_54509(.A(\to_acu2_0[12] ), .Z(n_40900));
	notech_inv i_54510(.A(\to_acu2_0[19] ), .Z(n_40901));
	notech_inv i_54511(.A(\to_acu2_0[20] ), .Z(n_40902));
	notech_inv i_54512(.A(\to_acu2_0[21] ), .Z(n_40903));
	notech_inv i_54513(.A(\to_acu2_0[23] ), .Z(n_40904));
	notech_inv i_54514(.A(\to_acu2_0[22] ), .Z(n_40905));
	notech_inv i_54515(.A(\to_acu2_0[68] ), .Z(n_40906));
	notech_inv i_54516(.A(\to_acu2_0[27] ), .Z(n_40907));
	notech_inv i_54517(.A(\to_acu2_0[26] ), .Z(n_40908));
	notech_inv i_54518(.A(\to_acu2_0[24] ), .Z(n_40909));
	notech_inv i_54519(.A(\to_acu2_0[25] ), .Z(n_40910));
	notech_inv i_54520(.A(\to_acu2_0[28] ), .Z(n_40911));
	notech_inv i_54521(.A(\to_acu2_0[16] ), .Z(n_40912));
	notech_inv i_54522(.A(\to_acu2_0[62] ), .Z(n_40913));
	notech_inv i_54523(.A(\to_acu2_0[69] ), .Z(n_40914));
	notech_inv i_54524(.A(\to_acu2_0[11] ), .Z(n_40915));
	notech_inv i_54525(.A(\to_acu2_0[9] ), .Z(n_40916));
	notech_inv i_54526(.A(in128[1]), .Z(n_40917));
	notech_inv i_54527(.A(in128[2]), .Z(n_40918));
	notech_inv i_54528(.A(sib_dec), .Z(n_40919));
	notech_inv i_54529(.A(mod_dec), .Z(n_40920));
	notech_inv i_54530(.A(\to_acu2_0[58] ), .Z(n_40921));
	notech_inv i_54531(.A(\to_acu2_0[10] ), .Z(n_40922));
	notech_inv i_54532(.A(\to_acu2_0[8] ), .Z(n_40923));
	notech_inv i_54533(.A(\to_acu2_0[6] ), .Z(n_40924));
	notech_inv i_54534(.A(\to_acu2_0[1] ), .Z(n_40925));
	notech_inv i_54535(.A(pc_req), .Z(n_40926));
	notech_inv i_54536(.A(n_58452), .Z(n_40927));
	notech_inv i_54537(.A(in128[9]), .Z(n_40928));
	notech_inv i_54538(.A(\nbus_12182[5] ), .Z(n_40929));
	notech_inv i_54539(.A(\nbus_12182[4] ), .Z(n_40930));
	notech_inv i_54540(.A(\nbus_12182[2] ), .Z(n_40931));
	notech_inv i_54541(.A(\nbus_12182[1] ), .Z(n_40932));
	notech_inv i_54542(.A(\nbus_12182[0] ), .Z(n_40933));
	notech_inv i_54543(.A(in128[11]), .Z(n_40934));
	notech_inv i_54544(.A(in128[12]), .Z(n_40935));
	notech_inv i_54545(.A(in128[13]), .Z(n_40936));
	notech_inv i_54546(.A(pg_fault), .Z(n_40937));
	notech_inv i_54547(.A(n_58991), .Z(n_40938));
	notech_inv i_54548(.A(twobyte), .Z(n_40939));
	notech_inv i_54549(.A(\to_acu2_0[4] ), .Z(n_40940));
	notech_inv i_54550(.A(\to_acu2_0[3] ), .Z(n_40941));
	notech_inv i_54551(.A(\to_acu2_0[0] ), .Z(n_40942));
	notech_inv i_54552(.A(\to_acu2_0[2] ), .Z(n_40943));
	notech_inv i_54553(.A(\to_acu2_0[7] ), .Z(n_40944));
	notech_inv i_54554(.A(int_main), .Z(n_40945));
	notech_inv i_54555(.A(\nbus_12182[3] ), .Z(n_40946));
	notech_inv i_54556(.A(in128[7]), .Z(n_40947));
	deco8 i_deco_1(.in8({in128[7], in128[6], in128[5], in128[4], in128[3], in128
		[2], in128[1], in128[0]}), .indic({\to_acu2_0[80] , \to_acu2_0[79] 
		, \to_acu2_0[78] , \to_acu2_0[77] , \to_acu2_0[76] , \to_acu2_0[75] 
		, \to_acu2_0[74] , \to_acu2_0[73] , \to_acu2_0[72] , \to_acu2_0[71] 
		, \to_acu2_0[70] , \to_acu2_0[69] , \to_acu2_0[68] , \to_acu2_0[67] 
		, \to_acu2_0[66] , \to_acu2_0[65] , \to_acu2_0[64] , \to_acu2_0[63] 
		, \to_acu2_0[62] , \to_acu2_0[61] , \to_acu2_0[60] , \to_acu2_0[59] 
		, \to_acu2_0[58] , \to_acu2_0[57] , \to_acu2_0[56] , \to_acu2_0[55] 
		, \to_acu2_0[54] , \to_acu2_0[53] , \to_acu2_0[52] , \to_acu2_0[51] 
		, \to_acu2_0[50] , \to_acu2_0[49] , \to_acu2_0[48] , \to_acu2_0[47] 
		, \to_acu2_0[46] , \to_acu2_0[45] , \to_acu2_0[44] , \to_acu2_0[43] 
		, \to_acu2_0[42] , \to_acu2_0[41] , \to_acu2_0[40] , 
		UNCONNECTED_000, \to_acu2_0[38] , \to_acu2_0[37] , \to_acu2_0[36] 
		, \to_acu2_0[35] , \to_acu2_0[34] , \to_acu2_0[33] , \to_acu2_0[32] 
		, \to_acu2_0[31] , \to_acu2_0[30] , \to_acu2_0[29] , \to_acu2_0[28] 
		, \to_acu2_0[27] , \to_acu2_0[26] , \to_acu2_0[25] , \to_acu2_0[24] 
		, \to_acu2_0[23] , \to_acu2_0[22] , \to_acu2_0[21] , \to_acu2_0[20] 
		, \to_acu2_0[19] , \to_acu2_0[18] , \to_acu2_0[17] , \to_acu2_0[16] 
		, \to_acu2_0[15] , \to_acu2_0[14] , \to_acu2_0[13] , \to_acu2_0[12] 
		, \to_acu2_0[11] , \to_acu2_0[10] , \to_acu2_0[9] , \to_acu2_0[8] 
		}));
	deco_rm i_deco_3(.in8({in128[15], in128[14], in128[13], in128[12], 
		UNCONNECTED_001, n_58451, in128[9], in128[8]}), .indic({\to_acu2_0[7] 
		, \to_acu2_0[6] , \to_acu2_0[5] , \to_acu2_0[4] , \to_acu2_0[3] 
		, \to_acu2_0[2] , \to_acu2_0[1] , \to_acu2_0[0] }));
	udecox i_udeco(.op({in128[7], in128[6], in128[5], in128[4], in128[3], in128
		[2], in128[1], in128[0]}), .modrm({in128[15], in128[14], in128[
		13], in128[12], in128[11], n_58452, in128[9], in128[8]}), .twobyte
		(twobyte), .cpl(cpl), .adz(adz), .opz(opz), .udeco(udeco), .fpu(n_58991
		), .emul(cr0[2]), .ipg_fault(ipg_fault));
	AWDP_partition_33 i_65708(.O0({\nbus_12182[5] , \nbus_12182[4] , \nbus_12182[3] 
		, \nbus_12182[2] , \nbus_12182[1] , \nbus_12182[0] }), .mod_dec(mod_dec
		), .sib_dec(sib_dec), .displc(displc), .imm_sz(imm_sz), .pfx_sz(pfx_sz
		), .twobyte(twobyte), .fpu(n_58991));
endmodule
module AWDP_ADD_0(O0, opb, I0);

	output [32:0] O0;
	input [31:0] opb;
	input [31:0] I0;




	notech_inv i_10541(.A(n_57226), .Z(n_57231));
	notech_inv i_10537(.A(n_57226), .Z(n_57227));
	notech_inv i_10536(.A(I0[18]), .Z(n_57226));
	notech_fa2 i_31(.A(n_57231), .B(n_354), .CI(opb[31]), .Z(O0[31]), .CO(O0
		[32]));
	notech_fa2 i_30(.A(n_57231), .B(n_352), .CI(opb[30]), .Z(O0[30]), .CO(n_354
		));
	notech_fa2 i_29(.A(n_57231), .B(n_350), .CI(opb[29]), .Z(O0[29]), .CO(n_352
		));
	notech_fa2 i_28(.A(n_57231), .B(n_348), .CI(opb[28]), .Z(O0[28]), .CO(n_350
		));
	notech_fa2 i_27(.A(n_57231), .B(n_346), .CI(opb[27]), .Z(O0[27]), .CO(n_348
		));
	notech_fa2 i_26(.A(n_57231), .B(n_344), .CI(opb[26]), .Z(O0[26]), .CO(n_346
		));
	notech_fa2 i_25(.A(n_57231), .B(n_342), .CI(opb[25]), .Z(O0[25]), .CO(n_344
		));
	notech_fa2 i_24(.A(n_57231), .B(n_340), .CI(opb[24]), .Z(O0[24]), .CO(n_342
		));
	notech_fa2 i_23(.A(n_57231), .B(n_338), .CI(opb[23]), .Z(O0[23]), .CO(n_340
		));
	notech_fa2 i_22(.A(n_57231), .B(n_336), .CI(opb[22]), .Z(O0[22]), .CO(n_338
		));
	notech_fa2 i_21(.A(n_57231), .B(n_334), .CI(opb[21]), .Z(O0[21]), .CO(n_336
		));
	notech_fa2 i_20(.A(n_57231), .B(n_332), .CI(opb[20]), .Z(O0[20]), .CO(n_334
		));
	notech_fa2 i_19(.A(n_57231), .B(n_330), .CI(opb[19]), .Z(O0[19]), .CO(n_332
		));
	notech_fa2 i_18(.A(n_57231), .B(n_328), .CI(opb[18]), .Z(O0[18]), .CO(n_330
		));
	notech_fa2 i_17(.A(n_57231), .B(n_326), .CI(opb[17]), .Z(O0[17]), .CO(n_328
		));
	notech_fa2 i_16(.A(n_57227), .B(n_324), .CI(opb[16]), .Z(O0[16]), .CO(n_326
		));
	notech_fa2 i_15(.A(n_57227), .B(n_322), .CI(opb[15]), .Z(O0[15]), .CO(n_324
		));
	notech_fa2 i_14(.A(n_57227), .B(n_320), .CI(opb[14]), .Z(O0[14]), .CO(n_322
		));
	notech_fa2 i_13(.A(n_57227), .B(n_318), .CI(opb[13]), .Z(O0[13]), .CO(n_320
		));
	notech_fa2 i_12(.A(n_57227), .B(n_316), .CI(opb[12]), .Z(O0[12]), .CO(n_318
		));
	notech_fa2 i_11(.A(n_57227), .B(n_314), .CI(opb[11]), .Z(O0[11]), .CO(n_316
		));
	notech_fa2 i_10(.A(n_57227), .B(n_312), .CI(opb[10]), .Z(O0[10]), .CO(n_314
		));
	notech_fa2 i_9(.A(n_57227), .B(n_310), .CI(opb[9]), .Z(O0[9]), .CO(n_312
		));
	notech_fa2 i_8(.A(n_57231), .B(n_308), .CI(opb[8]), .Z(O0[8]), .CO(n_310
		));
	notech_fa2 i_7(.A(n_57231), .B(n_306), .CI(opb[7]), .Z(O0[7]), .CO(n_308
		));
	notech_fa2 i_6(.A(n_57231), .B(n_304), .CI(opb[6]), .Z(O0[6]), .CO(n_306
		));
	notech_fa2 i_5(.A(n_57231), .B(n_302), .CI(opb[5]), .Z(O0[5]), .CO(n_304
		));
	notech_fa2 i_4(.A(n_57227), .B(n_300), .CI(opb[4]), .Z(O0[4]), .CO(n_302
		));
	notech_fa2 i_3(.A(n_57227), .B(n_298), .CI(opb[3]), .Z(O0[3]), .CO(n_300
		));
	notech_fa2 i_2(.A(n_57231), .B(n_296), .CI(opb[2]), .Z(O0[2]), .CO(n_298
		));
	notech_fa2 i_1(.A(I0[1]), .B(n_361), .CI(opb[1]), .Z(O0[1]), .CO(n_296)
		);
	notech_ha2 i_0(.A(opb[0]), .B(I0[0]), .Z(O0[0]), .CO(n_361));
endmodule
module AWDP_ADD_100(O0, opd, I0);

	output [32:0] O0;
	input [31:0] opd;
	input [31:0] I0;




	notech_inv i_10563(.A(n_57322), .Z(n_57327));
	notech_inv i_10559(.A(n_57322), .Z(n_57323));
	notech_inv i_10558(.A(I0[4]), .Z(n_57322));
	notech_fa2 i_31(.A(n_57327), .B(n_354), .CI(opd[31]), .Z(O0[31]), .CO(O0
		[32]));
	notech_fa2 i_30(.A(n_57327), .B(n_352), .CI(opd[30]), .Z(O0[30]), .CO(n_354
		));
	notech_fa2 i_29(.A(n_57327), .B(n_350), .CI(opd[29]), .Z(O0[29]), .CO(n_352
		));
	notech_fa2 i_28(.A(n_57327), .B(n_348), .CI(opd[28]), .Z(O0[28]), .CO(n_350
		));
	notech_fa2 i_27(.A(n_57327), .B(n_346), .CI(opd[27]), .Z(O0[27]), .CO(n_348
		));
	notech_fa2 i_26(.A(n_57327), .B(n_344), .CI(opd[26]), .Z(O0[26]), .CO(n_346
		));
	notech_fa2 i_25(.A(n_57327), .B(n_342), .CI(opd[25]), .Z(O0[25]), .CO(n_344
		));
	notech_fa2 i_24(.A(n_57327), .B(n_340), .CI(opd[24]), .Z(O0[24]), .CO(n_342
		));
	notech_fa2 i_23(.A(n_57327), .B(n_338), .CI(opd[23]), .Z(O0[23]), .CO(n_340
		));
	notech_fa2 i_22(.A(n_57327), .B(n_336), .CI(opd[22]), .Z(O0[22]), .CO(n_338
		));
	notech_fa2 i_21(.A(n_57327), .B(n_334), .CI(opd[21]), .Z(O0[21]), .CO(n_336
		));
	notech_fa2 i_20(.A(n_57327), .B(n_332), .CI(opd[20]), .Z(O0[20]), .CO(n_334
		));
	notech_fa2 i_19(.A(n_57327), .B(n_330), .CI(opd[19]), .Z(O0[19]), .CO(n_332
		));
	notech_fa2 i_18(.A(n_57327), .B(n_328), .CI(opd[18]), .Z(O0[18]), .CO(n_330
		));
	notech_fa2 i_17(.A(n_57327), .B(n_326), .CI(opd[17]), .Z(O0[17]), .CO(n_328
		));
	notech_fa2 i_16(.A(n_57323), .B(n_324), .CI(opd[16]), .Z(O0[16]), .CO(n_326
		));
	notech_fa2 i_15(.A(n_57323), .B(n_322), .CI(opd[15]), .Z(O0[15]), .CO(n_324
		));
	notech_fa2 i_14(.A(n_57323), .B(n_320), .CI(opd[14]), .Z(O0[14]), .CO(n_322
		));
	notech_fa2 i_13(.A(n_57323), .B(n_318), .CI(opd[13]), .Z(O0[13]), .CO(n_320
		));
	notech_fa2 i_12(.A(n_57323), .B(n_316), .CI(opd[12]), .Z(O0[12]), .CO(n_318
		));
	notech_fa2 i_11(.A(n_57323), .B(n_314), .CI(opd[11]), .Z(O0[11]), .CO(n_316
		));
	notech_fa2 i_10(.A(n_57323), .B(n_312), .CI(opd[10]), .Z(O0[10]), .CO(n_314
		));
	notech_fa2 i_9(.A(n_57323), .B(n_310), .CI(opd[9]), .Z(O0[9]), .CO(n_312
		));
	notech_fa2 i_8(.A(n_57327), .B(n_308), .CI(opd[8]), .Z(O0[8]), .CO(n_310
		));
	notech_fa2 i_7(.A(n_57327), .B(n_306), .CI(opd[7]), .Z(O0[7]), .CO(n_308
		));
	notech_fa2 i_6(.A(n_57327), .B(n_304), .CI(opd[6]), .Z(O0[6]), .CO(n_306
		));
	notech_fa2 i_5(.A(n_57327), .B(n_302), .CI(opd[5]), .Z(O0[5]), .CO(n_304
		));
	notech_fa2 i_4(.A(n_57323), .B(n_300), .CI(opd[4]), .Z(O0[4]), .CO(n_302
		));
	notech_fa2 i_3(.A(n_57323), .B(n_298), .CI(opd[3]), .Z(O0[3]), .CO(n_300
		));
	notech_fa2 i_2(.A(n_57327), .B(n_296), .CI(opd[2]), .Z(O0[2]), .CO(n_298
		));
	notech_fa2 i_1(.A(I0[1]), .B(n_361), .CI(opd[1]), .Z(O0[1]), .CO(n_296)
		);
	notech_ha2 i_0(.A(opd[0]), .B(I0[0]), .Z(O0[0]), .CO(n_361));
endmodule
module AWDP_ADD_102(O0, I0, I1);

	output [31:0] O0;
	input [31:0] I0;
	input [31:0] I1;

	wire \I0[4] ;
	wire \I0[5] ;
	wire \I0[6] ;
	wire \I0[7] ;
	wire \I0[8] ;
	wire \I0[9] ;
	wire \I0[10] ;
	wire \I0[11] ;
	wire \I0[12] ;
	wire \I0[13] ;
	wire \I0[14] ;
	wire \I0[15] ;


	assign O0[0] = I0[0];
	assign O0[1] = I0[1];
	assign O0[2] = I0[2];
	assign O0[3] = I0[3];
	assign \I0[4]  = I0[4];
	assign \I0[5]  = I0[5];
	assign \I0[6]  = I0[6];
	assign \I0[7]  = I0[7];
	assign \I0[8]  = I0[8];
	assign \I0[9]  = I0[9];
	assign \I0[10]  = I0[10];
	assign \I0[11]  = I0[11];
	assign \I0[12]  = I0[12];
	assign \I0[13]  = I0[13];
	assign \I0[14]  = I0[14];
	assign \I0[15]  = I0[15];

	notech_ha2 i_27(.A(I1[31]), .B(n_376), .Z(O0[31]));
	notech_ha2 i_26(.A(I1[30]), .B(n_374), .Z(O0[30]), .CO(n_376));
	notech_ha2 i_25(.A(I1[29]), .B(n_372), .Z(O0[29]), .CO(n_374));
	notech_ha2 i_24(.A(I1[28]), .B(n_370), .Z(O0[28]), .CO(n_372));
	notech_ha2 i_23(.A(I1[27]), .B(n_368), .Z(O0[27]), .CO(n_370));
	notech_ha2 i_22(.A(I1[26]), .B(n_366), .Z(O0[26]), .CO(n_368));
	notech_ha2 i_21(.A(I1[25]), .B(n_364), .Z(O0[25]), .CO(n_366));
	notech_ha2 i_20(.A(I1[24]), .B(n_362), .Z(O0[24]), .CO(n_364));
	notech_ha2 i_19(.A(I1[23]), .B(n_360), .Z(O0[23]), .CO(n_362));
	notech_ha2 i_18(.A(I1[22]), .B(n_358), .Z(O0[22]), .CO(n_360));
	notech_ha2 i_17(.A(I1[21]), .B(n_356), .Z(O0[21]), .CO(n_358));
	notech_ha2 i_16(.A(I1[20]), .B(n_354), .Z(O0[20]), .CO(n_356));
	notech_ha2 i_15(.A(I1[19]), .B(n_352), .Z(O0[19]), .CO(n_354));
	notech_ha2 i_14(.A(I1[18]), .B(n_350), .Z(O0[18]), .CO(n_352));
	notech_ha2 i_13(.A(I1[17]), .B(n_348), .Z(O0[17]), .CO(n_350));
	notech_ha2 i_12(.A(I1[16]), .B(n_311), .Z(O0[16]), .CO(n_348));
	notech_fa2 i_11(.A(\I0[15] ), .B(n_309), .CI(I1[15]), .Z(O0[15]), .CO(n_311
		));
	notech_fa2 i_10(.A(\I0[14] ), .B(n_307), .CI(I1[14]), .Z(O0[14]), .CO(n_309
		));
	notech_fa2 i_9(.A(\I0[13] ), .B(n_305), .CI(I1[13]), .Z(O0[13]), .CO(n_307
		));
	notech_fa2 i_8(.A(\I0[12] ), .B(n_303), .CI(I1[12]), .Z(O0[12]), .CO(n_305
		));
	notech_fa2 i_7(.A(\I0[11] ), .B(n_301), .CI(I1[11]), .Z(O0[11]), .CO(n_303
		));
	notech_fa2 i_6(.A(\I0[10] ), .B(n_299), .CI(I1[10]), .Z(O0[10]), .CO(n_301
		));
	notech_fa2 i_5(.A(\I0[9] ), .B(n_297), .CI(I1[9]), .Z(O0[9]), .CO(n_299)
		);
	notech_fa2 i_4(.A(\I0[8] ), .B(n_295), .CI(I1[8]), .Z(O0[8]), .CO(n_297)
		);
	notech_fa2 i_3(.A(\I0[7] ), .B(n_293), .CI(I1[7]), .Z(O0[7]), .CO(n_295)
		);
	notech_fa2 i_2(.A(\I0[6] ), .B(n_291), .CI(I1[6]), .Z(O0[6]), .CO(n_293)
		);
	notech_fa2 i_1(.A(\I0[5] ), .B(n_346), .CI(I1[5]), .Z(O0[5]), .CO(n_291)
		);
	notech_ha2 i_0(.A(\I0[4] ), .B(I1[4]), .Z(O0[4]), .CO(n_346));
endmodule
module AWDP_ADD_109(O0, opb, I0);

	output [16:0] O0;
	input [15:0] opb;
	input [15:0] I0;




	notech_fa2 i_15(.A(I0[15]), .B(n_178), .CI(opb[15]), .Z(O0[15]), .CO(O0[
		16]));
	notech_fa2 i_14(.A(I0[15]), .B(n_176), .CI(opb[14]), .Z(O0[14]), .CO(n_178
		));
	notech_fa2 i_13(.A(I0[15]), .B(n_174), .CI(opb[13]), .Z(O0[13]), .CO(n_176
		));
	notech_fa2 i_12(.A(I0[15]), .B(n_172), .CI(opb[12]), .Z(O0[12]), .CO(n_174
		));
	notech_fa2 i_11(.A(I0[15]), .B(n_170), .CI(opb[11]), .Z(O0[11]), .CO(n_172
		));
	notech_fa2 i_10(.A(I0[15]), .B(n_168), .CI(opb[10]), .Z(O0[10]), .CO(n_170
		));
	notech_fa2 i_9(.A(I0[15]), .B(n_166), .CI(opb[9]), .Z(O0[9]), .CO(n_168)
		);
	notech_fa2 i_8(.A(I0[15]), .B(n_164), .CI(opb[8]), .Z(O0[8]), .CO(n_166)
		);
	notech_fa2 i_7(.A(I0[15]), .B(n_162), .CI(opb[7]), .Z(O0[7]), .CO(n_164)
		);
	notech_fa2 i_6(.A(I0[15]), .B(n_160), .CI(opb[6]), .Z(O0[6]), .CO(n_162)
		);
	notech_fa2 i_5(.A(I0[15]), .B(n_158), .CI(opb[5]), .Z(O0[5]), .CO(n_160)
		);
	notech_fa2 i_4(.A(I0[15]), .B(n_156), .CI(opb[4]), .Z(O0[4]), .CO(n_158)
		);
	notech_fa2 i_3(.A(I0[15]), .B(n_154), .CI(opb[3]), .Z(O0[3]), .CO(n_156)
		);
	notech_fa2 i_2(.A(I0[15]), .B(n_152), .CI(opb[2]), .Z(O0[2]), .CO(n_154)
		);
	notech_fa2 i_1(.A(I0[1]), .B(n_185), .CI(opb[1]), .Z(O0[1]), .CO(n_152)
		);
	notech_ha2 i_0(.A(opb[0]), .B(I0[0]), .Z(O0[0]), .CO(n_185));
endmodule
module AWDP_ADD_114(O0, regs_4, calc_sz);
    output [31:0] O0;
    input [31:0] regs_4;
    input [2:0] calc_sz;
    // Line 470
    wire [31:0] N104;
    // Line 348
    wire [31:0] O0;

    // Line 470
    assign N104 = calc_sz + regs_4;
    // Line 348
    assign O0 = N104;
endmodule

module AWDP_ADD_116(O0, opa, I0);

	output [32:0] O0;
	input [31:0] opa;
	input [31:0] I0;




	notech_inv i_10551(.A(n_57284), .Z(n_57285));
	notech_inv i_10550(.A(I0[19]), .Z(n_57284));
	notech_fa2 i_31(.A(I0[19]), .B(n_354), .CI(opa[31]), .Z(O0[31]), .CO(O0[
		32]));
	notech_fa2 i_30(.A(I0[19]), .B(n_352), .CI(opa[30]), .Z(O0[30]), .CO(n_354
		));
	notech_fa2 i_29(.A(I0[19]), .B(n_350), .CI(opa[29]), .Z(O0[29]), .CO(n_352
		));
	notech_fa2 i_28(.A(I0[19]), .B(n_348), .CI(opa[28]), .Z(O0[28]), .CO(n_350
		));
	notech_fa2 i_27(.A(I0[19]), .B(n_346), .CI(opa[27]), .Z(O0[27]), .CO(n_348
		));
	notech_fa2 i_26(.A(I0[19]), .B(n_344), .CI(opa[26]), .Z(O0[26]), .CO(n_346
		));
	notech_fa2 i_25(.A(I0[19]), .B(n_342), .CI(opa[25]), .Z(O0[25]), .CO(n_344
		));
	notech_fa2 i_24(.A(I0[19]), .B(n_340), .CI(opa[24]), .Z(O0[24]), .CO(n_342
		));
	notech_fa2 i_23(.A(I0[19]), .B(n_338), .CI(opa[23]), .Z(O0[23]), .CO(n_340
		));
	notech_fa2 i_22(.A(I0[19]), .B(n_336), .CI(opa[22]), .Z(O0[22]), .CO(n_338
		));
	notech_fa2 i_21(.A(I0[19]), .B(n_334), .CI(opa[21]), .Z(O0[21]), .CO(n_336
		));
	notech_fa2 i_20(.A(I0[19]), .B(n_332), .CI(opa[20]), .Z(O0[20]), .CO(n_334
		));
	notech_fa2 i_19(.A(I0[19]), .B(n_330), .CI(opa[19]), .Z(O0[19]), .CO(n_332
		));
	notech_fa2 i_18(.A(I0[19]), .B(n_328), .CI(opa[18]), .Z(O0[18]), .CO(n_330
		));
	notech_fa2 i_17(.A(I0[19]), .B(n_326), .CI(opa[17]), .Z(O0[17]), .CO(n_328
		));
	notech_fa2 i_16(.A(n_57285), .B(n_324), .CI(opa[16]), .Z(O0[16]), .CO(n_326
		));
	notech_fa2 i_15(.A(n_57285), .B(n_322), .CI(opa[15]), .Z(O0[15]), .CO(n_324
		));
	notech_fa2 i_14(.A(n_57285), .B(n_320), .CI(opa[14]), .Z(O0[14]), .CO(n_322
		));
	notech_fa2 i_13(.A(n_57285), .B(n_318), .CI(opa[13]), .Z(O0[13]), .CO(n_320
		));
	notech_fa2 i_12(.A(n_57285), .B(n_316), .CI(opa[12]), .Z(O0[12]), .CO(n_318
		));
	notech_fa2 i_11(.A(n_57285), .B(n_314), .CI(opa[11]), .Z(O0[11]), .CO(n_316
		));
	notech_fa2 i_10(.A(n_57285), .B(n_312), .CI(opa[10]), .Z(O0[10]), .CO(n_314
		));
	notech_fa2 i_9(.A(n_57285), .B(n_310), .CI(opa[9]), .Z(O0[9]), .CO(n_312
		));
	notech_fa2 i_8(.A(n_57285), .B(n_308), .CI(opa[8]), .Z(O0[8]), .CO(n_310
		));
	notech_fa2 i_7(.A(n_57285), .B(n_306), .CI(opa[7]), .Z(O0[7]), .CO(n_308
		));
	notech_fa2 i_6(.A(n_57285), .B(n_304), .CI(opa[6]), .Z(O0[6]), .CO(n_306
		));
	notech_fa2 i_5(.A(n_57285), .B(n_302), .CI(opa[5]), .Z(O0[5]), .CO(n_304
		));
	notech_fa2 i_4(.A(n_57285), .B(n_300), .CI(opa[4]), .Z(O0[4]), .CO(n_302
		));
	notech_fa2 i_3(.A(n_57285), .B(n_298), .CI(opa[3]), .Z(O0[3]), .CO(n_300
		));
	notech_fa2 i_2(.A(n_57285), .B(n_296), .CI(opa[2]), .Z(O0[2]), .CO(n_298
		));
	notech_fa2 i_1(.A(I0[1]), .B(n_361), .CI(opa[1]), .Z(O0[1]), .CO(n_296)
		);
	notech_ha2 i_0(.A(opa[0]), .B(I0[0]), .Z(O0[0]), .CO(n_361));
endmodule
module AWDP_ADD_121(O0, opa, opd);
    output [8:0] O0;
    input [7:0] opa;
    input [7:0] opd;
    // Line 601
    wire [8:0] N124;
    // Line 601
    wire [8:0] O0;

    // Line 601
    assign N124 = opa + opd;
    // Line 601
    assign O0 = N124;
endmodule

module AWDP_ADD_123(O0, opd);

	output [31:0] O0;
	input [31:0] opd;

	wire \opd[2] ;
	wire \opd[3] ;
	wire \opd[4] ;
	wire \opd[5] ;
	wire \opd[6] ;
	wire \opd[7] ;
	wire \opd[8] ;
	wire \opd[9] ;
	wire \opd[10] ;
	wire \opd[11] ;
	wire \opd[12] ;
	wire \opd[13] ;
	wire \opd[14] ;
	wire \opd[15] ;
	wire \opd[16] ;
	wire \opd[17] ;
	wire \opd[18] ;
	wire \opd[19] ;
	wire \opd[20] ;
	wire \opd[21] ;
	wire \opd[22] ;
	wire \opd[23] ;
	wire \opd[24] ;
	wire \opd[25] ;
	wire \opd[26] ;
	wire \opd[27] ;
	wire \opd[28] ;
	wire \opd[29] ;
	wire \opd[30] ;
	wire \opd[31] ;


	assign O0[0] = opd[0];
	assign O0[1] = opd[1];
	assign \opd[2]  = opd[2];
	assign \opd[3]  = opd[3];
	assign \opd[4]  = opd[4];
	assign \opd[5]  = opd[5];
	assign \opd[6]  = opd[6];
	assign \opd[7]  = opd[7];
	assign \opd[8]  = opd[8];
	assign \opd[9]  = opd[9];
	assign \opd[10]  = opd[10];
	assign \opd[11]  = opd[11];
	assign \opd[12]  = opd[12];
	assign \opd[13]  = opd[13];
	assign \opd[14]  = opd[14];
	assign \opd[15]  = opd[15];
	assign \opd[16]  = opd[16];
	assign \opd[17]  = opd[17];
	assign \opd[18]  = opd[18];
	assign \opd[19]  = opd[19];
	assign \opd[20]  = opd[20];
	assign \opd[21]  = opd[21];
	assign \opd[22]  = opd[22];
	assign \opd[23]  = opd[23];
	assign \opd[24]  = opd[24];
	assign \opd[25]  = opd[25];
	assign \opd[26]  = opd[26];
	assign \opd[27]  = opd[27];
	assign \opd[28]  = opd[28];
	assign \opd[29]  = opd[29];
	assign \opd[30]  = opd[30];
	assign \opd[31]  = opd[31];

	notech_ha2 i_29(.A(\opd[31] ), .B(n_308), .Z(O0[31]));
	notech_ha2 i_28(.A(\opd[30] ), .B(n_306), .Z(O0[30]), .CO(n_308));
	notech_ha2 i_27(.A(\opd[29] ), .B(n_304), .Z(O0[29]), .CO(n_306));
	notech_ha2 i_26(.A(\opd[28] ), .B(n_302), .Z(O0[28]), .CO(n_304));
	notech_ha2 i_25(.A(\opd[27] ), .B(n_300), .Z(O0[27]), .CO(n_302));
	notech_ha2 i_24(.A(\opd[26] ), .B(n_298), .Z(O0[26]), .CO(n_300));
	notech_ha2 i_23(.A(\opd[25] ), .B(n_296), .Z(O0[25]), .CO(n_298));
	notech_ha2 i_22(.A(\opd[24] ), .B(n_294), .Z(O0[24]), .CO(n_296));
	notech_ha2 i_21(.A(\opd[23] ), .B(n_292), .Z(O0[23]), .CO(n_294));
	notech_ha2 i_20(.A(\opd[22] ), .B(n_290), .Z(O0[22]), .CO(n_292));
	notech_ha2 i_19(.A(\opd[21] ), .B(n_288), .Z(O0[21]), .CO(n_290));
	notech_ha2 i_18(.A(\opd[20] ), .B(n_286), .Z(O0[20]), .CO(n_288));
	notech_ha2 i_17(.A(\opd[19] ), .B(n_284), .Z(O0[19]), .CO(n_286));
	notech_ha2 i_16(.A(\opd[18] ), .B(n_282), .Z(O0[18]), .CO(n_284));
	notech_ha2 i_15(.A(\opd[17] ), .B(n_280), .Z(O0[17]), .CO(n_282));
	notech_ha2 i_14(.A(\opd[16] ), .B(n_278), .Z(O0[16]), .CO(n_280));
	notech_ha2 i_13(.A(\opd[15] ), .B(n_276), .Z(O0[15]), .CO(n_278));
	notech_ha2 i_12(.A(\opd[14] ), .B(n_274), .Z(O0[14]), .CO(n_276));
	notech_ha2 i_11(.A(\opd[13] ), .B(n_272), .Z(O0[13]), .CO(n_274));
	notech_ha2 i_10(.A(\opd[12] ), .B(n_270), .Z(O0[12]), .CO(n_272));
	notech_ha2 i_9(.A(\opd[11] ), .B(n_268), .Z(O0[11]), .CO(n_270));
	notech_ha2 i_8(.A(\opd[10] ), .B(n_266), .Z(O0[10]), .CO(n_268));
	notech_ha2 i_7(.A(\opd[9] ), .B(n_264), .Z(O0[9]), .CO(n_266));
	notech_ha2 i_6(.A(\opd[8] ), .B(n_262), .Z(O0[8]), .CO(n_264));
	notech_ha2 i_5(.A(\opd[7] ), .B(n_260), .Z(O0[7]), .CO(n_262));
	notech_ha2 i_4(.A(\opd[6] ), .B(n_258), .Z(O0[6]), .CO(n_260));
	notech_ha2 i_3(.A(\opd[5] ), .B(n_256), .Z(O0[5]), .CO(n_258));
	notech_ha2 i_2(.A(\opd[4] ), .B(n_254), .Z(O0[4]), .CO(n_256));
	notech_ha2 i_1(.A(\opd[3] ), .B(\opd[2] ), .Z(O0[3]), .CO(n_254));
	notech_inv i_0(.A(\opd[2] ), .Z(O0[2]));
endmodule
module AWDP_ADD_149(O0, opd, I0);

	output [16:0] O0;
	input [15:0] opd;
	input [15:0] I0;




	notech_fa2 i_15(.A(I0[4]), .B(n_178), .CI(opd[15]), .Z(O0[15]), .CO(O0[
		16]));
	notech_fa2 i_14(.A(I0[4]), .B(n_176), .CI(opd[14]), .Z(O0[14]), .CO(n_178
		));
	notech_fa2 i_13(.A(I0[4]), .B(n_174), .CI(opd[13]), .Z(O0[13]), .CO(n_176
		));
	notech_fa2 i_12(.A(I0[4]), .B(n_172), .CI(opd[12]), .Z(O0[12]), .CO(n_174
		));
	notech_fa2 i_11(.A(I0[4]), .B(n_170), .CI(opd[11]), .Z(O0[11]), .CO(n_172
		));
	notech_fa2 i_10(.A(I0[4]), .B(n_168), .CI(opd[10]), .Z(O0[10]), .CO(n_170
		));
	notech_fa2 i_9(.A(I0[4]), .B(n_166), .CI(opd[9]), .Z(O0[9]), .CO(n_168)
		);
	notech_fa2 i_8(.A(I0[4]), .B(n_164), .CI(opd[8]), .Z(O0[8]), .CO(n_166)
		);
	notech_fa2 i_7(.A(I0[4]), .B(n_162), .CI(opd[7]), .Z(O0[7]), .CO(n_164)
		);
	notech_fa2 i_6(.A(I0[4]), .B(n_160), .CI(opd[6]), .Z(O0[6]), .CO(n_162)
		);
	notech_fa2 i_5(.A(I0[4]), .B(n_158), .CI(opd[5]), .Z(O0[5]), .CO(n_160)
		);
	notech_fa2 i_4(.A(I0[4]), .B(n_156), .CI(opd[4]), .Z(O0[4]), .CO(n_158)
		);
	notech_fa2 i_3(.A(I0[4]), .B(n_154), .CI(opd[3]), .Z(O0[3]), .CO(n_156)
		);
	notech_fa2 i_2(.A(I0[4]), .B(n_152), .CI(opd[2]), .Z(O0[2]), .CO(n_154)
		);
	notech_fa2 i_1(.A(I0[1]), .B(n_185), .CI(opd[1]), .Z(O0[1]), .CO(n_152)
		);
	notech_ha2 i_0(.A(opd[0]), .B(I0[0]), .Z(O0[0]), .CO(n_185));
endmodule
module AWDP_ADD_166(O0, ldtr, I0);

	output [31:0] O0;
	input [31:0] ldtr;
	input [31:0] I0;

	wire \ldtr[1] ;
	wire \ldtr[2] ;
	wire \ldtr[3] ;
	wire \ldtr[4] ;
	wire \ldtr[5] ;
	wire \ldtr[6] ;
	wire \ldtr[7] ;
	wire \ldtr[8] ;
	wire \ldtr[9] ;
	wire \ldtr[10] ;
	wire \ldtr[11] ;
	wire \ldtr[12] ;
	wire \ldtr[13] ;
	wire \ldtr[14] ;
	wire \ldtr[15] ;
	wire \ldtr[16] ;
	wire \ldtr[17] ;
	wire \ldtr[18] ;
	wire \ldtr[19] ;
	wire \ldtr[20] ;
	wire \ldtr[21] ;
	wire \ldtr[22] ;
	wire \ldtr[23] ;
	wire \ldtr[24] ;
	wire \ldtr[25] ;
	wire \ldtr[26] ;
	wire \ldtr[27] ;
	wire \ldtr[28] ;
	wire \ldtr[29] ;
	wire \ldtr[30] ;
	wire \ldtr[31] ;


	assign O0[0] = ldtr[0];
	assign \ldtr[1]  = ldtr[1];
	assign \ldtr[2]  = ldtr[2];
	assign \ldtr[3]  = ldtr[3];
	assign \ldtr[4]  = ldtr[4];
	assign \ldtr[5]  = ldtr[5];
	assign \ldtr[6]  = ldtr[6];
	assign \ldtr[7]  = ldtr[7];
	assign \ldtr[8]  = ldtr[8];
	assign \ldtr[9]  = ldtr[9];
	assign \ldtr[10]  = ldtr[10];
	assign \ldtr[11]  = ldtr[11];
	assign \ldtr[12]  = ldtr[12];
	assign \ldtr[13]  = ldtr[13];
	assign \ldtr[14]  = ldtr[14];
	assign \ldtr[15]  = ldtr[15];
	assign \ldtr[16]  = ldtr[16];
	assign \ldtr[17]  = ldtr[17];
	assign \ldtr[18]  = ldtr[18];
	assign \ldtr[19]  = ldtr[19];
	assign \ldtr[20]  = ldtr[20];
	assign \ldtr[21]  = ldtr[21];
	assign \ldtr[22]  = ldtr[22];
	assign \ldtr[23]  = ldtr[23];
	assign \ldtr[24]  = ldtr[24];
	assign \ldtr[25]  = ldtr[25];
	assign \ldtr[26]  = ldtr[26];
	assign \ldtr[27]  = ldtr[27];
	assign \ldtr[28]  = ldtr[28];
	assign \ldtr[29]  = ldtr[29];
	assign \ldtr[30]  = ldtr[30];
	assign \ldtr[31]  = ldtr[31];

	notech_fa2 i_30(.A(I0[31]), .B(n_347), .CI(\ldtr[31] ), .Z(O0[31]));
	notech_fa2 i_29(.A(I0[30]), .B(n_345), .CI(\ldtr[30] ), .Z(O0[30]), .CO(n_347
		));
	notech_fa2 i_28(.A(I0[29]), .B(n_343), .CI(\ldtr[29] ), .Z(O0[29]), .CO(n_345
		));
	notech_fa2 i_27(.A(I0[28]), .B(n_341), .CI(\ldtr[28] ), .Z(O0[28]), .CO(n_343
		));
	notech_fa2 i_26(.A(I0[27]), .B(n_339), .CI(\ldtr[27] ), .Z(O0[27]), .CO(n_341
		));
	notech_fa2 i_25(.A(I0[26]), .B(n_337), .CI(\ldtr[26] ), .Z(O0[26]), .CO(n_339
		));
	notech_fa2 i_24(.A(I0[25]), .B(n_335), .CI(\ldtr[25] ), .Z(O0[25]), .CO(n_337
		));
	notech_fa2 i_23(.A(I0[24]), .B(n_333), .CI(\ldtr[24] ), .Z(O0[24]), .CO(n_335
		));
	notech_fa2 i_22(.A(I0[23]), .B(n_331), .CI(\ldtr[23] ), .Z(O0[23]), .CO(n_333
		));
	notech_fa2 i_21(.A(I0[22]), .B(n_329), .CI(\ldtr[22] ), .Z(O0[22]), .CO(n_331
		));
	notech_fa2 i_20(.A(I0[21]), .B(n_327), .CI(\ldtr[21] ), .Z(O0[21]), .CO(n_329
		));
	notech_fa2 i_19(.A(I0[20]), .B(n_325), .CI(\ldtr[20] ), .Z(O0[20]), .CO(n_327
		));
	notech_fa2 i_18(.A(I0[19]), .B(n_323), .CI(\ldtr[19] ), .Z(O0[19]), .CO(n_325
		));
	notech_fa2 i_17(.A(I0[18]), .B(n_321), .CI(\ldtr[18] ), .Z(O0[18]), .CO(n_323
		));
	notech_fa2 i_16(.A(I0[17]), .B(n_319), .CI(\ldtr[17] ), .Z(O0[17]), .CO(n_321
		));
	notech_fa2 i_15(.A(I0[16]), .B(n_317), .CI(\ldtr[16] ), .Z(O0[16]), .CO(n_319
		));
	notech_fa2 i_14(.A(I0[15]), .B(n_315), .CI(\ldtr[15] ), .Z(O0[15]), .CO(n_317
		));
	notech_fa2 i_13(.A(I0[14]), .B(n_313), .CI(\ldtr[14] ), .Z(O0[14]), .CO(n_315
		));
	notech_fa2 i_12(.A(I0[13]), .B(n_311), .CI(\ldtr[13] ), .Z(O0[13]), .CO(n_313
		));
	notech_fa2 i_11(.A(I0[12]), .B(n_309), .CI(\ldtr[12] ), .Z(O0[12]), .CO(n_311
		));
	notech_fa2 i_10(.A(I0[11]), .B(n_307), .CI(\ldtr[11] ), .Z(O0[11]), .CO(n_309
		));
	notech_fa2 i_9(.A(I0[10]), .B(n_305), .CI(\ldtr[10] ), .Z(O0[10]), .CO(n_307
		));
	notech_fa2 i_8(.A(I0[9]), .B(n_303), .CI(\ldtr[9] ), .Z(O0[9]), .CO(n_305
		));
	notech_fa2 i_7(.A(I0[8]), .B(n_301), .CI(\ldtr[8] ), .Z(O0[8]), .CO(n_303
		));
	notech_fa2 i_6(.A(I0[7]), .B(n_299), .CI(\ldtr[7] ), .Z(O0[7]), .CO(n_301
		));
	notech_fa2 i_5(.A(I0[6]), .B(n_297), .CI(\ldtr[6] ), .Z(O0[6]), .CO(n_299
		));
	notech_fa2 i_4(.A(I0[5]), .B(n_295), .CI(\ldtr[5] ), .Z(O0[5]), .CO(n_297
		));
	notech_fa2 i_3(.A(I0[4]), .B(n_293), .CI(\ldtr[4] ), .Z(O0[4]), .CO(n_295
		));
	notech_fa2 i_2(.A(I0[3]), .B(n_354), .CI(\ldtr[3] ), .Z(O0[3]), .CO(n_293
		));
	notech_ha2 i_1(.A(\ldtr[2] ), .B(\ldtr[1] ), .Z(O0[2]), .CO(n_354));
	notech_inv i_0(.A(\ldtr[1] ), .Z(O0[1]));
endmodule
module AWDP_ADD_168(O0, opa, opd);
    output [32:0] O0;
    input [31:0] opa;
    input [31:0] opd;
    // Line 599
    wire [32:0] O0;
    // Line 599
    wire [32:0] N172;

    // Line 599
    assign O0 = N172;
    // Line 599
    assign N172 = opa + opd;
endmodule

module AWDP_ADD_169(O0, gdtr, I0);

	output [31:0] O0;
	input [31:0] gdtr;
	input [31:0] I0;

	wire \gdtr[1] ;
	wire \gdtr[2] ;
	wire \gdtr[3] ;
	wire \gdtr[4] ;
	wire \gdtr[5] ;
	wire \gdtr[6] ;
	wire \gdtr[7] ;
	wire \gdtr[8] ;
	wire \gdtr[9] ;
	wire \gdtr[10] ;
	wire \gdtr[11] ;
	wire \gdtr[12] ;
	wire \gdtr[13] ;
	wire \gdtr[14] ;
	wire \gdtr[15] ;
	wire \gdtr[16] ;
	wire \gdtr[17] ;
	wire \gdtr[18] ;
	wire \gdtr[19] ;
	wire \gdtr[20] ;
	wire \gdtr[21] ;
	wire \gdtr[22] ;
	wire \gdtr[23] ;
	wire \gdtr[24] ;
	wire \gdtr[25] ;
	wire \gdtr[26] ;
	wire \gdtr[27] ;
	wire \gdtr[28] ;
	wire \gdtr[29] ;
	wire \gdtr[30] ;
	wire \gdtr[31] ;


	assign O0[0] = gdtr[0];
	assign \gdtr[1]  = gdtr[1];
	assign \gdtr[2]  = gdtr[2];
	assign \gdtr[3]  = gdtr[3];
	assign \gdtr[4]  = gdtr[4];
	assign \gdtr[5]  = gdtr[5];
	assign \gdtr[6]  = gdtr[6];
	assign \gdtr[7]  = gdtr[7];
	assign \gdtr[8]  = gdtr[8];
	assign \gdtr[9]  = gdtr[9];
	assign \gdtr[10]  = gdtr[10];
	assign \gdtr[11]  = gdtr[11];
	assign \gdtr[12]  = gdtr[12];
	assign \gdtr[13]  = gdtr[13];
	assign \gdtr[14]  = gdtr[14];
	assign \gdtr[15]  = gdtr[15];
	assign \gdtr[16]  = gdtr[16];
	assign \gdtr[17]  = gdtr[17];
	assign \gdtr[18]  = gdtr[18];
	assign \gdtr[19]  = gdtr[19];
	assign \gdtr[20]  = gdtr[20];
	assign \gdtr[21]  = gdtr[21];
	assign \gdtr[22]  = gdtr[22];
	assign \gdtr[23]  = gdtr[23];
	assign \gdtr[24]  = gdtr[24];
	assign \gdtr[25]  = gdtr[25];
	assign \gdtr[26]  = gdtr[26];
	assign \gdtr[27]  = gdtr[27];
	assign \gdtr[28]  = gdtr[28];
	assign \gdtr[29]  = gdtr[29];
	assign \gdtr[30]  = gdtr[30];
	assign \gdtr[31]  = gdtr[31];

	notech_fa2 i_30(.A(I0[31]), .B(n_347), .CI(\gdtr[31] ), .Z(O0[31]));
	notech_fa2 i_29(.A(I0[30]), .B(n_345), .CI(\gdtr[30] ), .Z(O0[30]), .CO(n_347
		));
	notech_fa2 i_28(.A(I0[29]), .B(n_343), .CI(\gdtr[29] ), .Z(O0[29]), .CO(n_345
		));
	notech_fa2 i_27(.A(I0[28]), .B(n_341), .CI(\gdtr[28] ), .Z(O0[28]), .CO(n_343
		));
	notech_fa2 i_26(.A(I0[27]), .B(n_339), .CI(\gdtr[27] ), .Z(O0[27]), .CO(n_341
		));
	notech_fa2 i_25(.A(I0[26]), .B(n_337), .CI(\gdtr[26] ), .Z(O0[26]), .CO(n_339
		));
	notech_fa2 i_24(.A(I0[25]), .B(n_335), .CI(\gdtr[25] ), .Z(O0[25]), .CO(n_337
		));
	notech_fa2 i_23(.A(I0[24]), .B(n_333), .CI(\gdtr[24] ), .Z(O0[24]), .CO(n_335
		));
	notech_fa2 i_22(.A(I0[23]), .B(n_331), .CI(\gdtr[23] ), .Z(O0[23]), .CO(n_333
		));
	notech_fa2 i_21(.A(I0[22]), .B(n_329), .CI(\gdtr[22] ), .Z(O0[22]), .CO(n_331
		));
	notech_fa2 i_20(.A(I0[21]), .B(n_327), .CI(\gdtr[21] ), .Z(O0[21]), .CO(n_329
		));
	notech_fa2 i_19(.A(I0[20]), .B(n_325), .CI(\gdtr[20] ), .Z(O0[20]), .CO(n_327
		));
	notech_fa2 i_18(.A(I0[19]), .B(n_323), .CI(\gdtr[19] ), .Z(O0[19]), .CO(n_325
		));
	notech_fa2 i_17(.A(I0[18]), .B(n_321), .CI(\gdtr[18] ), .Z(O0[18]), .CO(n_323
		));
	notech_fa2 i_16(.A(I0[17]), .B(n_319), .CI(\gdtr[17] ), .Z(O0[17]), .CO(n_321
		));
	notech_fa2 i_15(.A(I0[16]), .B(n_317), .CI(\gdtr[16] ), .Z(O0[16]), .CO(n_319
		));
	notech_fa2 i_14(.A(I0[15]), .B(n_315), .CI(\gdtr[15] ), .Z(O0[15]), .CO(n_317
		));
	notech_fa2 i_13(.A(I0[14]), .B(n_313), .CI(\gdtr[14] ), .Z(O0[14]), .CO(n_315
		));
	notech_fa2 i_12(.A(I0[13]), .B(n_311), .CI(\gdtr[13] ), .Z(O0[13]), .CO(n_313
		));
	notech_fa2 i_11(.A(I0[12]), .B(n_309), .CI(\gdtr[12] ), .Z(O0[12]), .CO(n_311
		));
	notech_fa2 i_10(.A(I0[11]), .B(n_307), .CI(\gdtr[11] ), .Z(O0[11]), .CO(n_309
		));
	notech_fa2 i_9(.A(I0[10]), .B(n_305), .CI(\gdtr[10] ), .Z(O0[10]), .CO(n_307
		));
	notech_fa2 i_8(.A(I0[9]), .B(n_303), .CI(\gdtr[9] ), .Z(O0[9]), .CO(n_305
		));
	notech_fa2 i_7(.A(I0[8]), .B(n_301), .CI(\gdtr[8] ), .Z(O0[8]), .CO(n_303
		));
	notech_fa2 i_6(.A(I0[7]), .B(n_299), .CI(\gdtr[7] ), .Z(O0[7]), .CO(n_301
		));
	notech_fa2 i_5(.A(I0[6]), .B(n_297), .CI(\gdtr[6] ), .Z(O0[6]), .CO(n_299
		));
	notech_fa2 i_4(.A(I0[5]), .B(n_295), .CI(\gdtr[5] ), .Z(O0[5]), .CO(n_297
		));
	notech_fa2 i_3(.A(I0[4]), .B(n_293), .CI(\gdtr[4] ), .Z(O0[4]), .CO(n_295
		));
	notech_fa2 i_2(.A(I0[3]), .B(n_354), .CI(\gdtr[3] ), .Z(O0[3]), .CO(n_293
		));
	notech_ha2 i_1(.A(\gdtr[2] ), .B(\gdtr[1] ), .Z(O0[2]), .CO(n_354));
	notech_inv i_0(.A(\gdtr[1] ), .Z(O0[1]));
endmodule
module AWDP_ADD_179(add_len_pc16, regs_14, lenpc);
    output [15:0] add_len_pc16;
    input [15:0] regs_14;
    input [15:0] lenpc;
    // Line 156
    wire [15:0] add_len_pc16;
    // Line 154
    wire [15:0] N206;

    // Line 156
    assign add_len_pc16 = N206;
    // Line 154
    assign N206 = lenpc + regs_14;
endmodule

module AWDP_ADD_21(O0, opa, opd);
    output [16:0] O0;
    input [15:0] opa;
    input [15:0] opd;
    // Line 600
    wire [16:0] N215;
    // Line 600
    wire [16:0] O0;

    // Line 600
    assign N215 = opa + opd;
    // Line 600
    assign O0 = N215;
endmodule

module AWDP_ADD_234(O0, opa, I0);

	output [16:0] O0;
	input [15:0] opa;
	input [15:0] I0;




	notech_fa2 i_15(.A(I0[13]), .B(n_178), .CI(opa[15]), .Z(O0[15]), .CO(O0[
		16]));
	notech_fa2 i_14(.A(I0[13]), .B(n_176), .CI(opa[14]), .Z(O0[14]), .CO(n_178
		));
	notech_fa2 i_13(.A(I0[13]), .B(n_174), .CI(opa[13]), .Z(O0[13]), .CO(n_176
		));
	notech_fa2 i_12(.A(I0[13]), .B(n_172), .CI(opa[12]), .Z(O0[12]), .CO(n_174
		));
	notech_fa2 i_11(.A(I0[13]), .B(n_170), .CI(opa[11]), .Z(O0[11]), .CO(n_172
		));
	notech_fa2 i_10(.A(I0[13]), .B(n_168), .CI(opa[10]), .Z(O0[10]), .CO(n_170
		));
	notech_fa2 i_9(.A(I0[13]), .B(n_166), .CI(opa[9]), .Z(O0[9]), .CO(n_168)
		);
	notech_fa2 i_8(.A(I0[13]), .B(n_164), .CI(opa[8]), .Z(O0[8]), .CO(n_166)
		);
	notech_fa2 i_7(.A(I0[13]), .B(n_162), .CI(opa[7]), .Z(O0[7]), .CO(n_164)
		);
	notech_fa2 i_6(.A(I0[13]), .B(n_160), .CI(opa[6]), .Z(O0[6]), .CO(n_162)
		);
	notech_fa2 i_5(.A(I0[13]), .B(n_158), .CI(opa[5]), .Z(O0[5]), .CO(n_160)
		);
	notech_fa2 i_4(.A(I0[13]), .B(n_156), .CI(opa[4]), .Z(O0[4]), .CO(n_158)
		);
	notech_fa2 i_3(.A(I0[13]), .B(n_154), .CI(opa[3]), .Z(O0[3]), .CO(n_156)
		);
	notech_fa2 i_2(.A(I0[13]), .B(n_152), .CI(opa[2]), .Z(O0[2]), .CO(n_154)
		);
	notech_fa2 i_1(.A(I0[1]), .B(n_185), .CI(opa[1]), .Z(O0[1]), .CO(n_152)
		);
	notech_ha2 i_0(.A(opa[0]), .B(I0[0]), .Z(O0[0]), .CO(n_185));
endmodule
module AWDP_ADD_24(O0, opd, desc);
    output [31:0] O0;
    input [31:0] opd;
    input [31:0] desc;
    // Line 1144
    wire [31:0] O0;
    // Line 1146
    wire [31:0] N235;

    // Line 1144
    assign O0 = N235;
    // Line 1146
    assign N235 = desc + opd;
endmodule

module AWDP_ADD_26(O0, opd, I0);

	output [31:0] O0;
	input [31:0] opd;
	input [31:0] I0;

	wire \opd[2] ;
	wire \opd[3] ;
	wire \opd[4] ;
	wire \opd[5] ;
	wire \opd[6] ;
	wire \opd[7] ;
	wire \opd[8] ;
	wire \opd[9] ;
	wire \opd[10] ;
	wire \opd[11] ;
	wire \opd[12] ;
	wire \opd[13] ;
	wire \opd[14] ;
	wire \opd[15] ;
	wire \opd[16] ;
	wire \opd[17] ;
	wire \opd[18] ;
	wire \opd[19] ;
	wire \opd[20] ;
	wire \opd[21] ;
	wire \opd[22] ;
	wire \opd[23] ;
	wire \opd[24] ;
	wire \opd[25] ;
	wire \opd[26] ;
	wire \opd[27] ;
	wire \opd[28] ;
	wire \opd[29] ;
	wire \opd[30] ;
	wire \opd[31] ;


	assign O0[0] = opd[0];
	assign O0[1] = opd[1];
	assign \opd[2]  = opd[2];
	assign \opd[3]  = opd[3];
	assign \opd[4]  = opd[4];
	assign \opd[5]  = opd[5];
	assign \opd[6]  = opd[6];
	assign \opd[7]  = opd[7];
	assign \opd[8]  = opd[8];
	assign \opd[9]  = opd[9];
	assign \opd[10]  = opd[10];
	assign \opd[11]  = opd[11];
	assign \opd[12]  = opd[12];
	assign \opd[13]  = opd[13];
	assign \opd[14]  = opd[14];
	assign \opd[15]  = opd[15];
	assign \opd[16]  = opd[16];
	assign \opd[17]  = opd[17];
	assign \opd[18]  = opd[18];
	assign \opd[19]  = opd[19];
	assign \opd[20]  = opd[20];
	assign \opd[21]  = opd[21];
	assign \opd[22]  = opd[22];
	assign \opd[23]  = opd[23];
	assign \opd[24]  = opd[24];
	assign \opd[25]  = opd[25];
	assign \opd[26]  = opd[26];
	assign \opd[27]  = opd[27];
	assign \opd[28]  = opd[28];
	assign \opd[29]  = opd[29];
	assign \opd[30]  = opd[30];
	assign \opd[31]  = opd[31];

	notech_ha2 i_29(.A(\opd[31] ), .B(n_354), .Z(O0[31]));
	notech_ha2 i_28(.A(\opd[30] ), .B(n_352), .Z(O0[30]), .CO(n_354));
	notech_ha2 i_27(.A(\opd[29] ), .B(n_341), .Z(O0[29]), .CO(n_352));
	notech_fa2 i_26(.A(I0[28]), .B(n_339), .CI(\opd[28] ), .Z(O0[28]), .CO(n_341
		));
	notech_fa2 i_25(.A(I0[27]), .B(n_337), .CI(\opd[27] ), .Z(O0[27]), .CO(n_339
		));
	notech_fa2 i_24(.A(I0[26]), .B(n_335), .CI(\opd[26] ), .Z(O0[26]), .CO(n_337
		));
	notech_fa2 i_23(.A(I0[25]), .B(n_333), .CI(\opd[25] ), .Z(O0[25]), .CO(n_335
		));
	notech_fa2 i_22(.A(I0[24]), .B(n_331), .CI(\opd[24] ), .Z(O0[24]), .CO(n_333
		));
	notech_fa2 i_21(.A(I0[23]), .B(n_329), .CI(\opd[23] ), .Z(O0[23]), .CO(n_331
		));
	notech_fa2 i_20(.A(I0[22]), .B(n_327), .CI(\opd[22] ), .Z(O0[22]), .CO(n_329
		));
	notech_fa2 i_19(.A(I0[21]), .B(n_325), .CI(\opd[21] ), .Z(O0[21]), .CO(n_327
		));
	notech_fa2 i_18(.A(I0[20]), .B(n_323), .CI(\opd[20] ), .Z(O0[20]), .CO(n_325
		));
	notech_fa2 i_17(.A(I0[19]), .B(n_321), .CI(\opd[19] ), .Z(O0[19]), .CO(n_323
		));
	notech_fa2 i_16(.A(I0[18]), .B(n_319), .CI(\opd[18] ), .Z(O0[18]), .CO(n_321
		));
	notech_fa2 i_15(.A(I0[17]), .B(n_317), .CI(\opd[17] ), .Z(O0[17]), .CO(n_319
		));
	notech_fa2 i_14(.A(I0[16]), .B(n_315), .CI(\opd[16] ), .Z(O0[16]), .CO(n_317
		));
	notech_fa2 i_13(.A(I0[15]), .B(n_313), .CI(\opd[15] ), .Z(O0[15]), .CO(n_315
		));
	notech_fa2 i_12(.A(I0[14]), .B(n_311), .CI(\opd[14] ), .Z(O0[14]), .CO(n_313
		));
	notech_fa2 i_11(.A(I0[13]), .B(n_309), .CI(\opd[13] ), .Z(O0[13]), .CO(n_311
		));
	notech_fa2 i_10(.A(I0[12]), .B(n_307), .CI(\opd[12] ), .Z(O0[12]), .CO(n_309
		));
	notech_fa2 i_9(.A(I0[11]), .B(n_305), .CI(\opd[11] ), .Z(O0[11]), .CO(n_307
		));
	notech_fa2 i_8(.A(I0[10]), .B(n_303), .CI(\opd[10] ), .Z(O0[10]), .CO(n_305
		));
	notech_fa2 i_7(.A(I0[9]), .B(n_301), .CI(\opd[9] ), .Z(O0[9]), .CO(n_303
		));
	notech_fa2 i_6(.A(I0[8]), .B(n_299), .CI(\opd[8] ), .Z(O0[8]), .CO(n_301
		));
	notech_fa2 i_5(.A(I0[7]), .B(n_297), .CI(\opd[7] ), .Z(O0[7]), .CO(n_299
		));
	notech_fa2 i_4(.A(I0[6]), .B(n_295), .CI(\opd[6] ), .Z(O0[6]), .CO(n_297
		));
	notech_fa2 i_3(.A(I0[5]), .B(n_293), .CI(\opd[5] ), .Z(O0[5]), .CO(n_295
		));
	notech_fa2 i_2(.A(I0[4]), .B(n_291), .CI(\opd[4] ), .Z(O0[4]), .CO(n_293
		));
	notech_fa2 i_1(.A(I0[3]), .B(n_350), .CI(\opd[3] ), .Z(O0[3]), .CO(n_291
		));
	notech_ha2 i_0(.A(I0[2]), .B(\opd[2] ), .Z(O0[2]), .CO(n_350));
endmodule
module AWDP_ADD_40(O0, opb, I0);

	output [31:0] O0;
	input [31:0] opb;
	input [31:0] I0;




	notech_ha2 i_31(.A(opb[31]), .B(n_400), .Z(O0[31]));
	notech_ha2 i_30(.A(opb[30]), .B(n_398), .Z(O0[30]), .CO(n_400));
	notech_ha2 i_29(.A(opb[29]), .B(n_396), .Z(O0[29]), .CO(n_398));
	notech_ha2 i_28(.A(opb[28]), .B(n_394), .Z(O0[28]), .CO(n_396));
	notech_ha2 i_27(.A(opb[27]), .B(n_392), .Z(O0[27]), .CO(n_394));
	notech_ha2 i_26(.A(opb[26]), .B(n_390), .Z(O0[26]), .CO(n_392));
	notech_ha2 i_25(.A(opb[25]), .B(n_388), .Z(O0[25]), .CO(n_390));
	notech_ha2 i_24(.A(opb[24]), .B(n_386), .Z(O0[24]), .CO(n_388));
	notech_ha2 i_23(.A(opb[23]), .B(n_384), .Z(O0[23]), .CO(n_386));
	notech_ha2 i_22(.A(opb[22]), .B(n_382), .Z(O0[22]), .CO(n_384));
	notech_ha2 i_21(.A(opb[21]), .B(n_380), .Z(O0[21]), .CO(n_382));
	notech_ha2 i_20(.A(opb[20]), .B(n_378), .Z(O0[20]), .CO(n_380));
	notech_ha2 i_19(.A(opb[19]), .B(n_376), .Z(O0[19]), .CO(n_378));
	notech_ha2 i_18(.A(opb[18]), .B(n_374), .Z(O0[18]), .CO(n_376));
	notech_ha2 i_17(.A(opb[17]), .B(n_372), .Z(O0[17]), .CO(n_374));
	notech_ha2 i_16(.A(opb[16]), .B(n_370), .Z(O0[16]), .CO(n_372));
	notech_ha2 i_15(.A(opb[15]), .B(n_368), .Z(O0[15]), .CO(n_370));
	notech_ha2 i_14(.A(opb[14]), .B(n_366), .Z(O0[14]), .CO(n_368));
	notech_ha2 i_13(.A(opb[13]), .B(n_364), .Z(O0[13]), .CO(n_366));
	notech_ha2 i_12(.A(opb[12]), .B(n_362), .Z(O0[12]), .CO(n_364));
	notech_ha2 i_11(.A(opb[11]), .B(n_360), .Z(O0[11]), .CO(n_362));
	notech_ha2 i_10(.A(opb[10]), .B(n_358), .Z(O0[10]), .CO(n_360));
	notech_ha2 i_9(.A(opb[9]), .B(n_356), .Z(O0[9]), .CO(n_358));
	notech_ha2 i_8(.A(opb[8]), .B(n_303), .Z(O0[8]), .CO(n_356));
	notech_fa2 i_7(.A(I0[7]), .B(n_301), .CI(opb[7]), .Z(O0[7]), .CO(n_303)
		);
	notech_fa2 i_6(.A(I0[6]), .B(n_299), .CI(opb[6]), .Z(O0[6]), .CO(n_301)
		);
	notech_fa2 i_5(.A(I0[5]), .B(n_297), .CI(opb[5]), .Z(O0[5]), .CO(n_299)
		);
	notech_fa2 i_4(.A(I0[4]), .B(n_295), .CI(opb[4]), .Z(O0[4]), .CO(n_297)
		);
	notech_fa2 i_3(.A(I0[3]), .B(n_293), .CI(opb[3]), .Z(O0[3]), .CO(n_295)
		);
	notech_fa2 i_2(.A(I0[2]), .B(n_291), .CI(opb[2]), .Z(O0[2]), .CO(n_293)
		);
	notech_fa2 i_1(.A(I0[1]), .B(n_354), .CI(opb[1]), .Z(O0[1]), .CO(n_291)
		);
	notech_ha2 i_0(.A(I0[0]), .B(opb[0]), .Z(O0[0]), .CO(n_354));
endmodule
module AWDP_ADD_44(O0, I0, add_len_pc);
    output [31:0] O0;
    input [31:0] I0;
    input [31:0] add_len_pc;
    // Line 879
    wire [31:0] N263;
    // Line 386
    wire [31:0] O0;

    // Line 879
    assign N263 = I0 + add_len_pc;
    // Line 386
    assign O0 = N263;
endmodule

module AWDP_ADD_47(O0, Daddrs);

	output [31:0] O0;
	input [31:0] Daddrs;

	wire \Daddrs[2] ;
	wire \Daddrs[3] ;
	wire \Daddrs[4] ;
	wire \Daddrs[5] ;
	wire \Daddrs[6] ;
	wire \Daddrs[7] ;
	wire \Daddrs[8] ;
	wire \Daddrs[9] ;
	wire \Daddrs[10] ;
	wire \Daddrs[11] ;
	wire \Daddrs[12] ;
	wire \Daddrs[13] ;
	wire \Daddrs[14] ;
	wire \Daddrs[15] ;
	wire \Daddrs[16] ;
	wire \Daddrs[17] ;
	wire \Daddrs[18] ;
	wire \Daddrs[19] ;
	wire \Daddrs[20] ;
	wire \Daddrs[21] ;
	wire \Daddrs[22] ;
	wire \Daddrs[23] ;
	wire \Daddrs[24] ;
	wire \Daddrs[25] ;
	wire \Daddrs[26] ;
	wire \Daddrs[27] ;
	wire \Daddrs[28] ;
	wire \Daddrs[29] ;
	wire \Daddrs[30] ;
	wire \Daddrs[31] ;


	assign O0[0] = Daddrs[0];
	assign O0[1] = Daddrs[1];
	assign \Daddrs[2]  = Daddrs[2];
	assign \Daddrs[3]  = Daddrs[3];
	assign \Daddrs[4]  = Daddrs[4];
	assign \Daddrs[5]  = Daddrs[5];
	assign \Daddrs[6]  = Daddrs[6];
	assign \Daddrs[7]  = Daddrs[7];
	assign \Daddrs[8]  = Daddrs[8];
	assign \Daddrs[9]  = Daddrs[9];
	assign \Daddrs[10]  = Daddrs[10];
	assign \Daddrs[11]  = Daddrs[11];
	assign \Daddrs[12]  = Daddrs[12];
	assign \Daddrs[13]  = Daddrs[13];
	assign \Daddrs[14]  = Daddrs[14];
	assign \Daddrs[15]  = Daddrs[15];
	assign \Daddrs[16]  = Daddrs[16];
	assign \Daddrs[17]  = Daddrs[17];
	assign \Daddrs[18]  = Daddrs[18];
	assign \Daddrs[19]  = Daddrs[19];
	assign \Daddrs[20]  = Daddrs[20];
	assign \Daddrs[21]  = Daddrs[21];
	assign \Daddrs[22]  = Daddrs[22];
	assign \Daddrs[23]  = Daddrs[23];
	assign \Daddrs[24]  = Daddrs[24];
	assign \Daddrs[25]  = Daddrs[25];
	assign \Daddrs[26]  = Daddrs[26];
	assign \Daddrs[27]  = Daddrs[27];
	assign \Daddrs[28]  = Daddrs[28];
	assign \Daddrs[29]  = Daddrs[29];
	assign \Daddrs[30]  = Daddrs[30];
	assign \Daddrs[31]  = Daddrs[31];

	notech_ha2 i_29(.A(\Daddrs[31] ), .B(n_308), .Z(O0[31]));
	notech_ha2 i_28(.A(\Daddrs[30] ), .B(n_306), .Z(O0[30]), .CO(n_308));
	notech_ha2 i_27(.A(\Daddrs[29] ), .B(n_304), .Z(O0[29]), .CO(n_306));
	notech_ha2 i_26(.A(\Daddrs[28] ), .B(n_302), .Z(O0[28]), .CO(n_304));
	notech_ha2 i_25(.A(\Daddrs[27] ), .B(n_300), .Z(O0[27]), .CO(n_302));
	notech_ha2 i_24(.A(\Daddrs[26] ), .B(n_298), .Z(O0[26]), .CO(n_300));
	notech_ha2 i_23(.A(\Daddrs[25] ), .B(n_296), .Z(O0[25]), .CO(n_298));
	notech_ha2 i_22(.A(\Daddrs[24] ), .B(n_294), .Z(O0[24]), .CO(n_296));
	notech_ha2 i_21(.A(\Daddrs[23] ), .B(n_292), .Z(O0[23]), .CO(n_294));
	notech_ha2 i_20(.A(\Daddrs[22] ), .B(n_290), .Z(O0[22]), .CO(n_292));
	notech_ha2 i_19(.A(\Daddrs[21] ), .B(n_288), .Z(O0[21]), .CO(n_290));
	notech_ha2 i_18(.A(\Daddrs[20] ), .B(n_286), .Z(O0[20]), .CO(n_288));
	notech_ha2 i_17(.A(\Daddrs[19] ), .B(n_284), .Z(O0[19]), .CO(n_286));
	notech_ha2 i_16(.A(\Daddrs[18] ), .B(n_282), .Z(O0[18]), .CO(n_284));
	notech_ha2 i_15(.A(\Daddrs[17] ), .B(n_280), .Z(O0[17]), .CO(n_282));
	notech_ha2 i_14(.A(\Daddrs[16] ), .B(n_278), .Z(O0[16]), .CO(n_280));
	notech_ha2 i_13(.A(\Daddrs[15] ), .B(n_276), .Z(O0[15]), .CO(n_278));
	notech_ha2 i_12(.A(\Daddrs[14] ), .B(n_274), .Z(O0[14]), .CO(n_276));
	notech_ha2 i_11(.A(\Daddrs[13] ), .B(n_272), .Z(O0[13]), .CO(n_274));
	notech_ha2 i_10(.A(\Daddrs[12] ), .B(n_270), .Z(O0[12]), .CO(n_272));
	notech_ha2 i_9(.A(\Daddrs[11] ), .B(n_268), .Z(O0[11]), .CO(n_270));
	notech_ha2 i_8(.A(\Daddrs[10] ), .B(n_266), .Z(O0[10]), .CO(n_268));
	notech_ha2 i_7(.A(\Daddrs[9] ), .B(n_264), .Z(O0[9]), .CO(n_266));
	notech_ha2 i_6(.A(\Daddrs[8] ), .B(n_262), .Z(O0[8]), .CO(n_264));
	notech_ha2 i_5(.A(\Daddrs[7] ), .B(n_260), .Z(O0[7]), .CO(n_262));
	notech_ha2 i_4(.A(\Daddrs[6] ), .B(n_258), .Z(O0[6]), .CO(n_260));
	notech_ha2 i_3(.A(\Daddrs[5] ), .B(n_256), .Z(O0[5]), .CO(n_258));
	notech_ha2 i_2(.A(\Daddrs[4] ), .B(n_254), .Z(O0[4]), .CO(n_256));
	notech_ha2 i_1(.A(\Daddrs[3] ), .B(\Daddrs[2] ), .Z(O0[3]), .CO(n_254)
		);
	notech_inv i_0(.A(\Daddrs[2] ), .Z(O0[2]));
endmodule
module AWDP_ADD_5(add_len_pc32, regs_14, lenpc);
    output [31:0] add_len_pc32;
    input [31:0] regs_14;
    input [31:0] lenpc;
    // Line 156
    wire [31:0] add_len_pc32;
    // Line 155
    wire [31:0] N355;

    // Line 156
    assign add_len_pc32 = N355;
    // Line 155
    assign N355 = lenpc + regs_14;
endmodule

module AWDP_ADD_61(O0, gdtr, I0);

	output [31:0] O0;
	input [31:0] gdtr;
	input [15:0] I0;

	wire \gdtr[1] ;
	wire \gdtr[2] ;
	wire \gdtr[3] ;
	wire \gdtr[4] ;
	wire \gdtr[5] ;
	wire \gdtr[6] ;
	wire \gdtr[7] ;
	wire \gdtr[8] ;
	wire \gdtr[9] ;
	wire \gdtr[10] ;
	wire \gdtr[11] ;
	wire \gdtr[12] ;
	wire \gdtr[13] ;
	wire \gdtr[14] ;
	wire \gdtr[15] ;
	wire \gdtr[16] ;
	wire \gdtr[17] ;
	wire \gdtr[18] ;
	wire \gdtr[19] ;
	wire \gdtr[20] ;
	wire \gdtr[21] ;
	wire \gdtr[22] ;
	wire \gdtr[23] ;
	wire \gdtr[24] ;
	wire \gdtr[25] ;
	wire \gdtr[26] ;
	wire \gdtr[27] ;
	wire \gdtr[28] ;
	wire \gdtr[29] ;
	wire \gdtr[30] ;
	wire \gdtr[31] ;


	assign O0[0] = gdtr[0];
	assign \gdtr[1]  = gdtr[1];
	assign \gdtr[2]  = gdtr[2];
	assign \gdtr[3]  = gdtr[3];
	assign \gdtr[4]  = gdtr[4];
	assign \gdtr[5]  = gdtr[5];
	assign \gdtr[6]  = gdtr[6];
	assign \gdtr[7]  = gdtr[7];
	assign \gdtr[8]  = gdtr[8];
	assign \gdtr[9]  = gdtr[9];
	assign \gdtr[10]  = gdtr[10];
	assign \gdtr[11]  = gdtr[11];
	assign \gdtr[12]  = gdtr[12];
	assign \gdtr[13]  = gdtr[13];
	assign \gdtr[14]  = gdtr[14];
	assign \gdtr[15]  = gdtr[15];
	assign \gdtr[16]  = gdtr[16];
	assign \gdtr[17]  = gdtr[17];
	assign \gdtr[18]  = gdtr[18];
	assign \gdtr[19]  = gdtr[19];
	assign \gdtr[20]  = gdtr[20];
	assign \gdtr[21]  = gdtr[21];
	assign \gdtr[22]  = gdtr[22];
	assign \gdtr[23]  = gdtr[23];
	assign \gdtr[24]  = gdtr[24];
	assign \gdtr[25]  = gdtr[25];
	assign \gdtr[26]  = gdtr[26];
	assign \gdtr[27]  = gdtr[27];
	assign \gdtr[28]  = gdtr[28];
	assign \gdtr[29]  = gdtr[29];
	assign \gdtr[30]  = gdtr[30];
	assign \gdtr[31]  = gdtr[31];

	notech_ha2 i_30(.A(\gdtr[31] ), .B(n_352), .Z(O0[31]));
	notech_ha2 i_29(.A(\gdtr[30] ), .B(n_350), .Z(O0[30]), .CO(n_352));
	notech_ha2 i_28(.A(\gdtr[29] ), .B(n_348), .Z(O0[29]), .CO(n_350));
	notech_ha2 i_27(.A(\gdtr[28] ), .B(n_346), .Z(O0[28]), .CO(n_348));
	notech_ha2 i_26(.A(\gdtr[27] ), .B(n_344), .Z(O0[27]), .CO(n_346));
	notech_ha2 i_25(.A(\gdtr[26] ), .B(n_342), .Z(O0[26]), .CO(n_344));
	notech_ha2 i_24(.A(\gdtr[25] ), .B(n_340), .Z(O0[25]), .CO(n_342));
	notech_ha2 i_23(.A(\gdtr[24] ), .B(n_338), .Z(O0[24]), .CO(n_340));
	notech_ha2 i_22(.A(\gdtr[23] ), .B(n_336), .Z(O0[23]), .CO(n_338));
	notech_ha2 i_21(.A(\gdtr[22] ), .B(n_334), .Z(O0[22]), .CO(n_336));
	notech_ha2 i_20(.A(\gdtr[21] ), .B(n_332), .Z(O0[21]), .CO(n_334));
	notech_ha2 i_19(.A(\gdtr[20] ), .B(n_330), .Z(O0[20]), .CO(n_332));
	notech_ha2 i_18(.A(\gdtr[19] ), .B(n_328), .Z(O0[19]), .CO(n_330));
	notech_ha2 i_17(.A(\gdtr[18] ), .B(n_326), .Z(O0[18]), .CO(n_328));
	notech_ha2 i_16(.A(\gdtr[17] ), .B(n_324), .Z(O0[17]), .CO(n_326));
	notech_ha2 i_15(.A(\gdtr[16] ), .B(n_285), .Z(O0[16]), .CO(n_324));
	notech_fa2 i_14(.A(I0[15]), .B(n_283), .CI(\gdtr[15] ), .Z(O0[15]), .CO(n_285
		));
	notech_fa2 i_13(.A(I0[14]), .B(n_281), .CI(\gdtr[14] ), .Z(O0[14]), .CO(n_283
		));
	notech_fa2 i_12(.A(I0[13]), .B(n_279), .CI(\gdtr[13] ), .Z(O0[13]), .CO(n_281
		));
	notech_fa2 i_11(.A(I0[12]), .B(n_277), .CI(\gdtr[12] ), .Z(O0[12]), .CO(n_279
		));
	notech_fa2 i_10(.A(I0[11]), .B(n_275), .CI(\gdtr[11] ), .Z(O0[11]), .CO(n_277
		));
	notech_fa2 i_9(.A(I0[10]), .B(n_273), .CI(\gdtr[10] ), .Z(O0[10]), .CO(n_275
		));
	notech_fa2 i_8(.A(I0[9]), .B(n_271), .CI(\gdtr[9] ), .Z(O0[9]), .CO(n_273
		));
	notech_fa2 i_7(.A(I0[8]), .B(n_269), .CI(\gdtr[8] ), .Z(O0[8]), .CO(n_271
		));
	notech_fa2 i_6(.A(I0[7]), .B(n_267), .CI(\gdtr[7] ), .Z(O0[7]), .CO(n_269
		));
	notech_fa2 i_5(.A(I0[6]), .B(n_265), .CI(\gdtr[6] ), .Z(O0[6]), .CO(n_267
		));
	notech_fa2 i_4(.A(I0[5]), .B(n_263), .CI(\gdtr[5] ), .Z(O0[5]), .CO(n_265
		));
	notech_fa2 i_3(.A(I0[4]), .B(n_261), .CI(\gdtr[4] ), .Z(O0[4]), .CO(n_263
		));
	notech_fa2 i_2(.A(I0[3]), .B(n_322), .CI(\gdtr[3] ), .Z(O0[3]), .CO(n_261
		));
	notech_ha2 i_1(.A(\gdtr[2] ), .B(\gdtr[1] ), .Z(O0[2]), .CO(n_322));
	notech_inv i_0(.A(\gdtr[1] ), .Z(O0[1]));
endmodule
module AWDP_ADD_62(O0, Daddrs);

	output [31:0] O0;
	input [31:0] Daddrs;

	wire \Daddrs[1] ;
	wire \Daddrs[2] ;
	wire \Daddrs[3] ;
	wire \Daddrs[4] ;
	wire \Daddrs[5] ;
	wire \Daddrs[6] ;
	wire \Daddrs[7] ;
	wire \Daddrs[8] ;
	wire \Daddrs[9] ;
	wire \Daddrs[10] ;
	wire \Daddrs[11] ;
	wire \Daddrs[12] ;
	wire \Daddrs[13] ;
	wire \Daddrs[14] ;
	wire \Daddrs[15] ;
	wire \Daddrs[16] ;
	wire \Daddrs[17] ;
	wire \Daddrs[18] ;
	wire \Daddrs[19] ;
	wire \Daddrs[20] ;
	wire \Daddrs[21] ;
	wire \Daddrs[22] ;
	wire \Daddrs[23] ;
	wire \Daddrs[24] ;
	wire \Daddrs[25] ;
	wire \Daddrs[26] ;
	wire \Daddrs[27] ;
	wire \Daddrs[28] ;
	wire \Daddrs[29] ;
	wire \Daddrs[30] ;
	wire \Daddrs[31] ;


	assign O0[0] = Daddrs[0];
	assign \Daddrs[1]  = Daddrs[1];
	assign \Daddrs[2]  = Daddrs[2];
	assign \Daddrs[3]  = Daddrs[3];
	assign \Daddrs[4]  = Daddrs[4];
	assign \Daddrs[5]  = Daddrs[5];
	assign \Daddrs[6]  = Daddrs[6];
	assign \Daddrs[7]  = Daddrs[7];
	assign \Daddrs[8]  = Daddrs[8];
	assign \Daddrs[9]  = Daddrs[9];
	assign \Daddrs[10]  = Daddrs[10];
	assign \Daddrs[11]  = Daddrs[11];
	assign \Daddrs[12]  = Daddrs[12];
	assign \Daddrs[13]  = Daddrs[13];
	assign \Daddrs[14]  = Daddrs[14];
	assign \Daddrs[15]  = Daddrs[15];
	assign \Daddrs[16]  = Daddrs[16];
	assign \Daddrs[17]  = Daddrs[17];
	assign \Daddrs[18]  = Daddrs[18];
	assign \Daddrs[19]  = Daddrs[19];
	assign \Daddrs[20]  = Daddrs[20];
	assign \Daddrs[21]  = Daddrs[21];
	assign \Daddrs[22]  = Daddrs[22];
	assign \Daddrs[23]  = Daddrs[23];
	assign \Daddrs[24]  = Daddrs[24];
	assign \Daddrs[25]  = Daddrs[25];
	assign \Daddrs[26]  = Daddrs[26];
	assign \Daddrs[27]  = Daddrs[27];
	assign \Daddrs[28]  = Daddrs[28];
	assign \Daddrs[29]  = Daddrs[29];
	assign \Daddrs[30]  = Daddrs[30];
	assign \Daddrs[31]  = Daddrs[31];

	notech_ha2 i_30(.A(\Daddrs[31] ), .B(n_312), .Z(O0[31]));
	notech_ha2 i_29(.A(\Daddrs[30] ), .B(n_310), .Z(O0[30]), .CO(n_312));
	notech_ha2 i_28(.A(\Daddrs[29] ), .B(n_308), .Z(O0[29]), .CO(n_310));
	notech_ha2 i_27(.A(\Daddrs[28] ), .B(n_306), .Z(O0[28]), .CO(n_308));
	notech_ha2 i_26(.A(\Daddrs[27] ), .B(n_304), .Z(O0[27]), .CO(n_306));
	notech_ha2 i_25(.A(\Daddrs[26] ), .B(n_302), .Z(O0[26]), .CO(n_304));
	notech_ha2 i_24(.A(\Daddrs[25] ), .B(n_300), .Z(O0[25]), .CO(n_302));
	notech_ha2 i_23(.A(\Daddrs[24] ), .B(n_298), .Z(O0[24]), .CO(n_300));
	notech_ha2 i_22(.A(\Daddrs[23] ), .B(n_296), .Z(O0[23]), .CO(n_298));
	notech_ha2 i_21(.A(\Daddrs[22] ), .B(n_294), .Z(O0[22]), .CO(n_296));
	notech_ha2 i_20(.A(\Daddrs[21] ), .B(n_292), .Z(O0[21]), .CO(n_294));
	notech_ha2 i_19(.A(\Daddrs[20] ), .B(n_290), .Z(O0[20]), .CO(n_292));
	notech_ha2 i_18(.A(\Daddrs[19] ), .B(n_288), .Z(O0[19]), .CO(n_290));
	notech_ha2 i_17(.A(\Daddrs[18] ), .B(n_286), .Z(O0[18]), .CO(n_288));
	notech_ha2 i_16(.A(\Daddrs[17] ), .B(n_284), .Z(O0[17]), .CO(n_286));
	notech_ha2 i_15(.A(\Daddrs[16] ), .B(n_282), .Z(O0[16]), .CO(n_284));
	notech_ha2 i_14(.A(\Daddrs[15] ), .B(n_280), .Z(O0[15]), .CO(n_282));
	notech_ha2 i_13(.A(\Daddrs[14] ), .B(n_278), .Z(O0[14]), .CO(n_280));
	notech_ha2 i_12(.A(\Daddrs[13] ), .B(n_276), .Z(O0[13]), .CO(n_278));
	notech_ha2 i_11(.A(\Daddrs[12] ), .B(n_274), .Z(O0[12]), .CO(n_276));
	notech_ha2 i_10(.A(\Daddrs[11] ), .B(n_272), .Z(O0[11]), .CO(n_274));
	notech_ha2 i_9(.A(\Daddrs[10] ), .B(n_270), .Z(O0[10]), .CO(n_272));
	notech_ha2 i_8(.A(\Daddrs[9] ), .B(n_268), .Z(O0[9]), .CO(n_270));
	notech_ha2 i_7(.A(\Daddrs[8] ), .B(n_266), .Z(O0[8]), .CO(n_268));
	notech_ha2 i_6(.A(\Daddrs[7] ), .B(n_264), .Z(O0[7]), .CO(n_266));
	notech_ha2 i_5(.A(\Daddrs[6] ), .B(n_262), .Z(O0[6]), .CO(n_264));
	notech_ha2 i_4(.A(\Daddrs[5] ), .B(n_260), .Z(O0[5]), .CO(n_262));
	notech_ha2 i_3(.A(\Daddrs[4] ), .B(n_258), .Z(O0[4]), .CO(n_260));
	notech_ha2 i_2(.A(\Daddrs[3] ), .B(n_256), .Z(O0[3]), .CO(n_258));
	notech_ha2 i_1(.A(\Daddrs[2] ), .B(\Daddrs[1] ), .Z(O0[2]), .CO(n_256)
		);
	notech_inv i_0(.A(\Daddrs[1] ), .Z(O0[1]));
endmodule
module AWDP_ADD_67(O0, regs_7, opd);
    output [31:0] O0;
    input [31:0] regs_7;
    input [31:0] opd;
    // Line 348
    wire [31:0] O0;
    // Line 520
    wire [31:0] N385;

    // Line 348
    assign O0 = N385;
    // Line 520
    assign N385 = regs_7 + opd;
endmodule

module AWDP_ADD_69(O0, regs_6, opd);
    output [31:0] O0;
    input [31:0] regs_6;
    input [31:0] opd;
    // Line 348
    wire [31:0] O0;
    // Line 520
    wire [31:0] N397;

    // Line 348
    assign O0 = N397;
    // Line 520
    assign N397 = regs_6 + opd;
endmodule

module AWDP_ADD_8(O0, opc, I0);
    output [31:0] O0;
    input [31:0] opc;
    input [31:0] I0;
    // Line 1006
    wire [31:0] O0;
    // Line 1006
    wire [31:0] N404;

    // Line 1006
    assign O0 = N404;
    // Line 1006
    assign N404 = opc + I0;
endmodule

module AWDP_ADD_92(O0, idtr, I0);

	output [31:0] O0;
	input [31:0] idtr;
	input [18:0] I0;

	wire \idtr[3] ;
	wire \idtr[4] ;
	wire \idtr[5] ;
	wire \idtr[6] ;
	wire \idtr[7] ;
	wire \idtr[8] ;
	wire \idtr[9] ;
	wire \idtr[10] ;
	wire \idtr[11] ;
	wire \idtr[12] ;
	wire \idtr[13] ;
	wire \idtr[14] ;
	wire \idtr[15] ;
	wire \idtr[16] ;
	wire \idtr[17] ;
	wire \idtr[18] ;
	wire \idtr[19] ;
	wire \idtr[20] ;
	wire \idtr[21] ;
	wire \idtr[22] ;
	wire \idtr[23] ;
	wire \idtr[24] ;
	wire \idtr[25] ;
	wire \idtr[26] ;
	wire \idtr[27] ;
	wire \idtr[28] ;
	wire \idtr[29] ;
	wire \idtr[30] ;
	wire \idtr[31] ;


	assign O0[0] = idtr[0];
	assign O0[1] = idtr[1];
	assign O0[2] = idtr[2];
	assign \idtr[3]  = idtr[3];
	assign \idtr[4]  = idtr[4];
	assign \idtr[5]  = idtr[5];
	assign \idtr[6]  = idtr[6];
	assign \idtr[7]  = idtr[7];
	assign \idtr[8]  = idtr[8];
	assign \idtr[9]  = idtr[9];
	assign \idtr[10]  = idtr[10];
	assign \idtr[11]  = idtr[11];
	assign \idtr[12]  = idtr[12];
	assign \idtr[13]  = idtr[13];
	assign \idtr[14]  = idtr[14];
	assign \idtr[15]  = idtr[15];
	assign \idtr[16]  = idtr[16];
	assign \idtr[17]  = idtr[17];
	assign \idtr[18]  = idtr[18];
	assign \idtr[19]  = idtr[19];
	assign \idtr[20]  = idtr[20];
	assign \idtr[21]  = idtr[21];
	assign \idtr[22]  = idtr[22];
	assign \idtr[23]  = idtr[23];
	assign \idtr[24]  = idtr[24];
	assign \idtr[25]  = idtr[25];
	assign \idtr[26]  = idtr[26];
	assign \idtr[27]  = idtr[27];
	assign \idtr[28]  = idtr[28];
	assign \idtr[29]  = idtr[29];
	assign \idtr[30]  = idtr[30];
	assign \idtr[31]  = idtr[31];

	notech_ha2 i_28(.A(\idtr[31] ), .B(n_346), .Z(O0[31]));
	notech_ha2 i_27(.A(\idtr[30] ), .B(n_344), .Z(O0[30]), .CO(n_346));
	notech_ha2 i_26(.A(\idtr[29] ), .B(n_342), .Z(O0[29]), .CO(n_344));
	notech_ha2 i_25(.A(\idtr[28] ), .B(n_340), .Z(O0[28]), .CO(n_342));
	notech_ha2 i_24(.A(\idtr[27] ), .B(n_338), .Z(O0[27]), .CO(n_340));
	notech_ha2 i_23(.A(\idtr[26] ), .B(n_336), .Z(O0[26]), .CO(n_338));
	notech_ha2 i_22(.A(\idtr[25] ), .B(n_334), .Z(O0[25]), .CO(n_336));
	notech_ha2 i_21(.A(\idtr[24] ), .B(n_332), .Z(O0[24]), .CO(n_334));
	notech_ha2 i_20(.A(\idtr[23] ), .B(n_330), .Z(O0[23]), .CO(n_332));
	notech_ha2 i_19(.A(\idtr[22] ), .B(n_328), .Z(O0[22]), .CO(n_330));
	notech_ha2 i_18(.A(\idtr[21] ), .B(n_326), .Z(O0[21]), .CO(n_328));
	notech_ha2 i_17(.A(\idtr[20] ), .B(n_324), .Z(O0[20]), .CO(n_326));
	notech_ha2 i_16(.A(\idtr[19] ), .B(n_293), .Z(O0[19]), .CO(n_324));
	notech_fa2 i_15(.A(I0[18]), .B(n_291), .CI(\idtr[18] ), .Z(O0[18]), .CO(n_293
		));
	notech_fa2 i_14(.A(I0[17]), .B(n_289), .CI(\idtr[17] ), .Z(O0[17]), .CO(n_291
		));
	notech_fa2 i_13(.A(I0[16]), .B(n_287), .CI(\idtr[16] ), .Z(O0[16]), .CO(n_289
		));
	notech_fa2 i_12(.A(I0[15]), .B(n_285), .CI(\idtr[15] ), .Z(O0[15]), .CO(n_287
		));
	notech_fa2 i_11(.A(I0[14]), .B(n_283), .CI(\idtr[14] ), .Z(O0[14]), .CO(n_285
		));
	notech_fa2 i_10(.A(I0[13]), .B(n_281), .CI(\idtr[13] ), .Z(O0[13]), .CO(n_283
		));
	notech_fa2 i_9(.A(I0[12]), .B(n_279), .CI(\idtr[12] ), .Z(O0[12]), .CO(n_281
		));
	notech_fa2 i_8(.A(I0[11]), .B(n_277), .CI(\idtr[11] ), .Z(O0[11]), .CO(n_279
		));
	notech_fa2 i_7(.A(I0[10]), .B(n_275), .CI(\idtr[10] ), .Z(O0[10]), .CO(n_277
		));
	notech_fa2 i_6(.A(I0[9]), .B(n_273), .CI(\idtr[9] ), .Z(O0[9]), .CO(n_275
		));
	notech_fa2 i_5(.A(I0[8]), .B(n_271), .CI(\idtr[8] ), .Z(O0[8]), .CO(n_273
		));
	notech_fa2 i_4(.A(I0[7]), .B(n_269), .CI(\idtr[7] ), .Z(O0[7]), .CO(n_271
		));
	notech_fa2 i_3(.A(I0[6]), .B(n_267), .CI(\idtr[6] ), .Z(O0[6]), .CO(n_269
		));
	notech_fa2 i_2(.A(I0[5]), .B(n_265), .CI(\idtr[5] ), .Z(O0[5]), .CO(n_267
		));
	notech_fa2 i_1(.A(I0[4]), .B(n_322), .CI(\idtr[4] ), .Z(O0[4]), .CO(n_265
		));
	notech_ha2 i_0(.A(\idtr[3] ), .B(I0[3]), .Z(O0[3]), .CO(n_322));
endmodule
module AWDP_DEC_155(O0, opc);

	output [7:0] O0;
	input [7:0] opc;




	notech_ha2 i_8(.A(n_48), .B(n_62), .Z(O0[7]));
	notech_inv i_1(.A(opc[0]), .Z(O0[0]));
	notech_inv i_0(.A(opc[7]), .Z(n_48));
	notech_xor2 i_61089(.A(opc[6]), .B(n_60), .Z(n_43632));
	notech_inv i_61090(.A(n_43632), .Z(O0[6]));
	notech_or2 i_61088(.A(opc[6]), .B(n_60), .Z(n_62));
	notech_xor2 i_27(.A(opc[5]), .B(n_58), .Z(n_43659));
	notech_inv i_28(.A(n_43659), .Z(O0[5]));
	notech_or2 i_26(.A(opc[5]), .B(n_58), .Z(n_60));
	notech_xor2 i_2795652(.A(opc[4]), .B(n_56), .Z(n_43686));
	notech_inv i_2895653(.A(n_43686), .Z(O0[4]));
	notech_or2 i_2695654(.A(opc[4]), .B(n_56), .Z(n_58));
	notech_xor2 i_2795655(.A(opc[3]), .B(n_54), .Z(n_43713));
	notech_inv i_2895656(.A(n_43713), .Z(O0[3]));
	notech_or2 i_2695657(.A(opc[3]), .B(n_54), .Z(n_56));
	notech_xor2 i_2795658(.A(opc[2]), .B(n_52), .Z(n_43740));
	notech_inv i_2895659(.A(n_43740), .Z(O0[2]));
	notech_or2 i_2695660(.A(opc[2]), .B(n_52), .Z(n_54));
	notech_xor2 i_2795661(.A(opc[1]), .B(opc[0]), .Z(n_43768));
	notech_inv i_2895662(.A(n_43768), .Z(O0[1]));
	notech_or2 i_2695663(.A(opc[1]), .B(opc[0]), .Z(n_52));
endmodule
module AWDP_DEC_2(O0, cx);

	output [15:0] O0;
	input [15:0] cx;




	notech_ha2 i_16(.A(n_96), .B(n_126), .Z(O0[15]));
	notech_inv i_1(.A(cx[0]), .Z(O0[0]));
	notech_inv i_0(.A(cx[15]), .Z(n_96));
	notech_xor2 i_33(.A(cx[14]), .B(n_124), .Z(n_43795));
	notech_inv i_34(.A(n_43795), .Z(O0[14]));
	notech_or2 i_32(.A(cx[14]), .B(n_124), .Z(n_126));
	notech_xor2 i_3295664(.A(cx[13]), .B(n_122), .Z(n_43822));
	notech_inv i_3395665(.A(n_43822), .Z(O0[13]));
	notech_or2 i_31(.A(cx[13]), .B(n_122), .Z(n_124));
	notech_xor2 i_30(.A(cx[12]), .B(n_120), .Z(n_43849));
	notech_inv i_3195666(.A(n_43849), .Z(O0[12]));
	notech_or2 i_29(.A(cx[12]), .B(n_120), .Z(n_122));
	notech_xor2 i_2995667(.A(cx[11]), .B(n_118), .Z(n_43876));
	notech_inv i_3095668(.A(n_43876), .Z(O0[11]));
	notech_or2 i_28(.A(cx[11]), .B(n_118), .Z(n_120));
	notech_xor2 i_2895669(.A(cx[10]), .B(n_116), .Z(n_43903));
	notech_inv i_2995670(.A(n_43903), .Z(O0[10]));
	notech_or2 i_27(.A(cx[10]), .B(n_116), .Z(n_118));
	notech_xor2 i_2795671(.A(cx[9]), .B(n_114), .Z(n_43930));
	notech_inv i_2895672(.A(n_43930), .Z(O0[9]));
	notech_or2 i_26(.A(cx[9]), .B(n_114), .Z(n_116));
	notech_xor2 i_2795673(.A(cx[8]), .B(n_112), .Z(n_43957));
	notech_inv i_2895674(.A(n_43957), .Z(O0[8]));
	notech_or2 i_2695675(.A(cx[8]), .B(n_112), .Z(n_114));
	notech_xor2 i_2795676(.A(cx[7]), .B(n_110), .Z(n_43984));
	notech_inv i_2895677(.A(n_43984), .Z(O0[7]));
	notech_or2 i_2695678(.A(cx[7]), .B(n_110), .Z(n_112));
	notech_xor2 i_2795679(.A(cx[6]), .B(n_108), .Z(n_44011));
	notech_inv i_2895680(.A(n_44011), .Z(O0[6]));
	notech_or2 i_2695681(.A(cx[6]), .B(n_108), .Z(n_110));
	notech_xor2 i_2795682(.A(cx[5]), .B(n_106), .Z(n_44038));
	notech_inv i_2895683(.A(n_44038), .Z(O0[5]));
	notech_or2 i_2695684(.A(cx[5]), .B(n_106), .Z(n_108));
	notech_xor2 i_2795685(.A(cx[4]), .B(n_104), .Z(n_44065));
	notech_inv i_2895686(.A(n_44065), .Z(O0[4]));
	notech_or2 i_2695687(.A(cx[4]), .B(n_104), .Z(n_106));
	notech_xor2 i_2795688(.A(cx[3]), .B(n_102), .Z(n_44092));
	notech_inv i_2895689(.A(n_44092), .Z(O0[3]));
	notech_or2 i_2695690(.A(cx[3]), .B(n_102), .Z(n_104));
	notech_xor2 i_2795691(.A(cx[2]), .B(n_100), .Z(n_44119));
	notech_inv i_2895692(.A(n_44119), .Z(O0[2]));
	notech_or2 i_2695693(.A(cx[2]), .B(n_100), .Z(n_102));
	notech_xor2 i_2795694(.A(cx[1]), .B(cx[0]), .Z(n_44147));
	notech_inv i_2895695(.A(n_44147), .Z(O0[1]));
	notech_or2 i_2695696(.A(cx[1]), .B(cx[0]), .Z(n_100));
endmodule
module AWDP_DEC_7(O0, ecx);

	output [31:0] O0;
	input [31:0] ecx;




	notech_ha2 i_32(.A(n_192), .B(n_254), .Z(O0[31]));
	notech_inv i_1(.A(ecx[0]), .Z(O0[0]));
	notech_inv i_0(.A(ecx[31]), .Z(n_192));
	notech_xor2 i_49(.A(ecx[30]), .B(n_252), .Z(n_44174));
	notech_inv i_50(.A(n_44174), .Z(O0[30]));
	notech_or2 i_48(.A(ecx[30]), .B(n_252), .Z(n_254));
	notech_xor2 i_4895697(.A(ecx[29]), .B(n_250), .Z(n_44201));
	notech_inv i_4995698(.A(n_44201), .Z(O0[29]));
	notech_or2 i_47(.A(ecx[29]), .B(n_250), .Z(n_252));
	notech_xor2 i_46(.A(ecx[28]), .B(n_248), .Z(n_44228));
	notech_inv i_4795699(.A(n_44228), .Z(O0[28]));
	notech_or2 i_45(.A(ecx[28]), .B(n_248), .Z(n_250));
	notech_xor2 i_4595700(.A(ecx[27]), .B(n_246), .Z(n_44255));
	notech_inv i_4695701(.A(n_44255), .Z(O0[27]));
	notech_or2 i_44(.A(ecx[27]), .B(n_246), .Z(n_248));
	notech_xor2 i_4495702(.A(ecx[26]), .B(n_244), .Z(n_44282));
	notech_inv i_4595703(.A(n_44282), .Z(O0[26]));
	notech_or2 i_43(.A(ecx[26]), .B(n_244), .Z(n_246));
	notech_xor2 i_4395704(.A(ecx[25]), .B(n_242), .Z(n_44309));
	notech_inv i_4495705(.A(n_44309), .Z(O0[25]));
	notech_or2 i_42(.A(ecx[25]), .B(n_242), .Z(n_244));
	notech_xor2 i_4295706(.A(ecx[24]), .B(n_240), .Z(n_44336));
	notech_inv i_4395707(.A(n_44336), .Z(O0[24]));
	notech_or2 i_41(.A(ecx[24]), .B(n_240), .Z(n_242));
	notech_xor2 i_4195708(.A(ecx[23]), .B(n_238), .Z(n_44363));
	notech_inv i_4295709(.A(n_44363), .Z(O0[23]));
	notech_or2 i_40(.A(ecx[23]), .B(n_238), .Z(n_240));
	notech_xor2 i_4095710(.A(ecx[22]), .B(n_236), .Z(n_44390));
	notech_inv i_4195711(.A(n_44390), .Z(O0[22]));
	notech_or2 i_39(.A(ecx[22]), .B(n_236), .Z(n_238));
	notech_xor2 i_3995712(.A(ecx[21]), .B(n_234), .Z(n_44417));
	notech_inv i_4095713(.A(n_44417), .Z(O0[21]));
	notech_or2 i_38(.A(ecx[21]), .B(n_234), .Z(n_236));
	notech_xor2 i_3895714(.A(ecx[20]), .B(n_232), .Z(n_44444));
	notech_inv i_3995715(.A(n_44444), .Z(O0[20]));
	notech_or2 i_37(.A(ecx[20]), .B(n_232), .Z(n_234));
	notech_xor2 i_3795716(.A(ecx[19]), .B(n_230), .Z(n_44471));
	notech_inv i_3895717(.A(n_44471), .Z(O0[19]));
	notech_or2 i_36(.A(ecx[19]), .B(n_230), .Z(n_232));
	notech_xor2 i_3695718(.A(ecx[18]), .B(n_228), .Z(n_44498));
	notech_inv i_3795719(.A(n_44498), .Z(O0[18]));
	notech_or2 i_35(.A(ecx[18]), .B(n_228), .Z(n_230));
	notech_xor2 i_3595720(.A(ecx[17]), .B(n_226), .Z(n_44525));
	notech_inv i_3695721(.A(n_44525), .Z(O0[17]));
	notech_or2 i_34(.A(ecx[17]), .B(n_226), .Z(n_228));
	notech_xor2 i_3495722(.A(ecx[16]), .B(n_224), .Z(n_44552));
	notech_inv i_3595723(.A(n_44552), .Z(O0[16]));
	notech_or2 i_33(.A(ecx[16]), .B(n_224), .Z(n_226));
	notech_xor2 i_3395724(.A(ecx[15]), .B(n_222), .Z(n_44579));
	notech_inv i_3495725(.A(n_44579), .Z(O0[15]));
	notech_or2 i_3295726(.A(ecx[15]), .B(n_222), .Z(n_224));
	notech_xor2 i_3295727(.A(ecx[14]), .B(n_220), .Z(n_44606));
	notech_inv i_3395728(.A(n_44606), .Z(O0[14]));
	notech_or2 i_31(.A(ecx[14]), .B(n_220), .Z(n_222));
	notech_xor2 i_3195729(.A(ecx[13]), .B(n_218), .Z(n_44633));
	notech_inv i_3295730(.A(n_44633), .Z(O0[13]));
	notech_or2 i_30(.A(ecx[13]), .B(n_218), .Z(n_220));
	notech_xor2 i_3095731(.A(ecx[12]), .B(n_216), .Z(n_44660));
	notech_inv i_3195732(.A(n_44660), .Z(O0[12]));
	notech_or2 i_29(.A(ecx[12]), .B(n_216), .Z(n_218));
	notech_xor2 i_2995733(.A(ecx[11]), .B(n_214), .Z(n_44687));
	notech_inv i_3095734(.A(n_44687), .Z(O0[11]));
	notech_or2 i_28(.A(ecx[11]), .B(n_214), .Z(n_216));
	notech_xor2 i_2895735(.A(ecx[10]), .B(n_212), .Z(n_44714));
	notech_inv i_2995736(.A(n_44714), .Z(O0[10]));
	notech_or2 i_27(.A(ecx[10]), .B(n_212), .Z(n_214));
	notech_xor2 i_2795737(.A(ecx[9]), .B(n_210), .Z(n_44741));
	notech_inv i_2895738(.A(n_44741), .Z(O0[9]));
	notech_or2 i_26(.A(ecx[9]), .B(n_210), .Z(n_212));
	notech_xor2 i_2795739(.A(ecx[8]), .B(n_208), .Z(n_44768));
	notech_inv i_2895740(.A(n_44768), .Z(O0[8]));
	notech_or2 i_2695741(.A(ecx[8]), .B(n_208), .Z(n_210));
	notech_xor2 i_2795742(.A(ecx[7]), .B(n_206), .Z(n_44795));
	notech_inv i_2895743(.A(n_44795), .Z(O0[7]));
	notech_or2 i_2695744(.A(ecx[7]), .B(n_206), .Z(n_208));
	notech_xor2 i_2795745(.A(ecx[6]), .B(n_204), .Z(n_44822));
	notech_inv i_2895746(.A(n_44822), .Z(O0[6]));
	notech_or2 i_2695747(.A(ecx[6]), .B(n_204), .Z(n_206));
	notech_xor2 i_2795748(.A(ecx[5]), .B(n_202), .Z(n_44849));
	notech_inv i_2895749(.A(n_44849), .Z(O0[5]));
	notech_or2 i_2695750(.A(ecx[5]), .B(n_202), .Z(n_204));
	notech_xor2 i_2795751(.A(ecx[4]), .B(n_200), .Z(n_44876));
	notech_inv i_2895752(.A(n_44876), .Z(O0[4]));
	notech_or2 i_2695753(.A(ecx[4]), .B(n_200), .Z(n_202));
	notech_xor2 i_2795754(.A(ecx[3]), .B(n_198), .Z(n_44903));
	notech_inv i_2895755(.A(n_44903), .Z(O0[3]));
	notech_or2 i_2695756(.A(ecx[3]), .B(n_198), .Z(n_200));
	notech_xor2 i_2795757(.A(ecx[2]), .B(n_196), .Z(n_44930));
	notech_inv i_2895758(.A(n_44930), .Z(O0[2]));
	notech_or2 i_2695759(.A(ecx[2]), .B(n_196), .Z(n_198));
	notech_xor2 i_2795760(.A(ecx[1]), .B(ecx[0]), .Z(n_44958));
	notech_inv i_2895761(.A(n_44958), .Z(O0[1]));
	notech_or2 i_2695762(.A(ecx[1]), .B(ecx[0]), .Z(n_196));
endmodule
module AWDP_DEC_83(O0, opc);

	output [31:0] O0;
	input [31:0] opc;




	notech_ha2 i_32(.A(n_192), .B(n_254), .Z(O0[31]));
	notech_inv i_1(.A(opc[0]), .Z(O0[0]));
	notech_inv i_0(.A(opc[31]), .Z(n_192));
	notech_xor2 i_49(.A(opc[30]), .B(n_252), .Z(n_44985));
	notech_inv i_50(.A(n_44985), .Z(O0[30]));
	notech_or2 i_48(.A(opc[30]), .B(n_252), .Z(n_254));
	notech_xor2 i_4895763(.A(opc[29]), .B(n_250), .Z(n_45012));
	notech_inv i_4995764(.A(n_45012), .Z(O0[29]));
	notech_or2 i_47(.A(opc[29]), .B(n_250), .Z(n_252));
	notech_xor2 i_46(.A(opc[28]), .B(n_248), .Z(n_45039));
	notech_inv i_4795765(.A(n_45039), .Z(O0[28]));
	notech_or2 i_45(.A(opc[28]), .B(n_248), .Z(n_250));
	notech_xor2 i_4595766(.A(opc[27]), .B(n_246), .Z(n_45066));
	notech_inv i_4695767(.A(n_45066), .Z(O0[27]));
	notech_or2 i_44(.A(opc[27]), .B(n_246), .Z(n_248));
	notech_xor2 i_4495768(.A(opc[26]), .B(n_244), .Z(n_45093));
	notech_inv i_4595769(.A(n_45093), .Z(O0[26]));
	notech_or2 i_43(.A(opc[26]), .B(n_244), .Z(n_246));
	notech_xor2 i_4395770(.A(opc[25]), .B(n_242), .Z(n_45120));
	notech_inv i_4495771(.A(n_45120), .Z(O0[25]));
	notech_or2 i_42(.A(opc[25]), .B(n_242), .Z(n_244));
	notech_xor2 i_4295772(.A(opc[24]), .B(n_240), .Z(n_45147));
	notech_inv i_4395773(.A(n_45147), .Z(O0[24]));
	notech_or2 i_41(.A(opc[24]), .B(n_240), .Z(n_242));
	notech_xor2 i_4195774(.A(opc[23]), .B(n_238), .Z(n_45174));
	notech_inv i_4295775(.A(n_45174), .Z(O0[23]));
	notech_or2 i_40(.A(opc[23]), .B(n_238), .Z(n_240));
	notech_xor2 i_4095776(.A(opc[22]), .B(n_236), .Z(n_45201));
	notech_inv i_4195777(.A(n_45201), .Z(O0[22]));
	notech_or2 i_39(.A(opc[22]), .B(n_236), .Z(n_238));
	notech_xor2 i_3995778(.A(opc[21]), .B(n_234), .Z(n_45228));
	notech_inv i_4095779(.A(n_45228), .Z(O0[21]));
	notech_or2 i_38(.A(opc[21]), .B(n_234), .Z(n_236));
	notech_xor2 i_3895780(.A(opc[20]), .B(n_232), .Z(n_45255));
	notech_inv i_3995781(.A(n_45255), .Z(O0[20]));
	notech_or2 i_37(.A(opc[20]), .B(n_232), .Z(n_234));
	notech_xor2 i_3795782(.A(opc[19]), .B(n_230), .Z(n_45282));
	notech_inv i_3895783(.A(n_45282), .Z(O0[19]));
	notech_or2 i_36(.A(opc[19]), .B(n_230), .Z(n_232));
	notech_xor2 i_3695784(.A(opc[18]), .B(n_228), .Z(n_45309));
	notech_inv i_3795785(.A(n_45309), .Z(O0[18]));
	notech_or2 i_35(.A(opc[18]), .B(n_228), .Z(n_230));
	notech_xor2 i_3595786(.A(opc[17]), .B(n_226), .Z(n_45336));
	notech_inv i_3695787(.A(n_45336), .Z(O0[17]));
	notech_or2 i_34(.A(opc[17]), .B(n_226), .Z(n_228));
	notech_xor2 i_3495788(.A(opc[16]), .B(n_224), .Z(n_45363));
	notech_inv i_3595789(.A(n_45363), .Z(O0[16]));
	notech_or2 i_33(.A(opc[16]), .B(n_224), .Z(n_226));
	notech_xor2 i_3395790(.A(opc[15]), .B(n_222), .Z(n_45390));
	notech_inv i_3495791(.A(n_45390), .Z(O0[15]));
	notech_or2 i_3295792(.A(opc[15]), .B(n_222), .Z(n_224));
	notech_xor2 i_3295793(.A(opc[14]), .B(n_220), .Z(n_45417));
	notech_inv i_3395794(.A(n_45417), .Z(O0[14]));
	notech_or2 i_31(.A(opc[14]), .B(n_220), .Z(n_222));
	notech_xor2 i_3195795(.A(opc[13]), .B(n_218), .Z(n_45444));
	notech_inv i_3295796(.A(n_45444), .Z(O0[13]));
	notech_or2 i_30(.A(opc[13]), .B(n_218), .Z(n_220));
	notech_xor2 i_3095797(.A(opc[12]), .B(n_216), .Z(n_45471));
	notech_inv i_3195798(.A(n_45471), .Z(O0[12]));
	notech_or2 i_29(.A(opc[12]), .B(n_216), .Z(n_218));
	notech_xor2 i_2995799(.A(opc[11]), .B(n_214), .Z(n_45498));
	notech_inv i_3095800(.A(n_45498), .Z(O0[11]));
	notech_or2 i_28(.A(opc[11]), .B(n_214), .Z(n_216));
	notech_xor2 i_2895801(.A(opc[10]), .B(n_212), .Z(n_45525));
	notech_inv i_2995802(.A(n_45525), .Z(O0[10]));
	notech_or2 i_27(.A(opc[10]), .B(n_212), .Z(n_214));
	notech_xor2 i_2795803(.A(opc[9]), .B(n_210), .Z(n_45552));
	notech_inv i_2895804(.A(n_45552), .Z(O0[9]));
	notech_or2 i_26(.A(opc[9]), .B(n_210), .Z(n_212));
	notech_xor2 i_2795805(.A(opc[8]), .B(n_208), .Z(n_45579));
	notech_inv i_2895806(.A(n_45579), .Z(O0[8]));
	notech_or2 i_2695807(.A(opc[8]), .B(n_208), .Z(n_210));
	notech_xor2 i_2795808(.A(opc[7]), .B(n_206), .Z(n_45606));
	notech_inv i_2895809(.A(n_45606), .Z(O0[7]));
	notech_or2 i_2695810(.A(opc[7]), .B(n_206), .Z(n_208));
	notech_xor2 i_2795811(.A(opc[6]), .B(n_204), .Z(n_45633));
	notech_inv i_2895812(.A(n_45633), .Z(O0[6]));
	notech_or2 i_2695813(.A(opc[6]), .B(n_204), .Z(n_206));
	notech_xor2 i_2795814(.A(opc[5]), .B(n_202), .Z(n_45660));
	notech_inv i_2895815(.A(n_45660), .Z(O0[5]));
	notech_or2 i_2695816(.A(opc[5]), .B(n_202), .Z(n_204));
	notech_xor2 i_2795817(.A(opc[4]), .B(n_200), .Z(n_45687));
	notech_inv i_2895818(.A(n_45687), .Z(O0[4]));
	notech_or2 i_2695819(.A(opc[4]), .B(n_200), .Z(n_202));
	notech_xor2 i_2795820(.A(opc[3]), .B(n_198), .Z(n_45714));
	notech_inv i_2895821(.A(n_45714), .Z(O0[3]));
	notech_or2 i_2695822(.A(opc[3]), .B(n_198), .Z(n_200));
	notech_xor2 i_2795823(.A(opc[2]), .B(n_196), .Z(n_45741));
	notech_inv i_2895824(.A(n_45741), .Z(O0[2]));
	notech_or2 i_2695825(.A(opc[2]), .B(n_196), .Z(n_198));
	notech_xor2 i_2795826(.A(opc[1]), .B(opc[0]), .Z(n_45769));
	notech_inv i_2895827(.A(n_45769), .Z(O0[1]));
	notech_or2 i_2695828(.A(opc[1]), .B(opc[0]), .Z(n_196));
endmodule
module AWDP_EQ_111(O0, mul64);
    output [0:0] O0;
    input [63:8] mul64;
    // Line 125
    wire [0:0] N554;
    // Line 125
    wire [0:0] O0;

    // Line 125
    assign N554 = mul64 == 56'h0;
    // Line 125
    assign O0 = N554;
endmodule

module AWDP_EQ_124(O0, mul64);
    output [0:0] O0;
    input [63:16] mul64;
    // Line 130
    wire [0:0] N564;
    // Line 130
    wire [0:0] O0;

    // Line 130
    assign N564 = mul64 == 48'hffffffff;
    // Line 130
    assign O0 = N564;
endmodule

module AWDP_EQ_128(O0, mul64);
    output [0:0] O0;
    input [63:16] mul64;
    // Line 126
    wire [0:0] N577;
    // Line 126
    wire [0:0] O0;

    // Line 126
    assign N577 = mul64 == 48'h0;
    // Line 126
    assign O0 = N577;
endmodule

module AWDP_EQ_158(O0, I0, I1);
    output [0:0] O0;
    input [63:0] I0;
    input [63:0] I1;
    // Line 790
    wire [0:0] N596;
    // Line 790
    wire [0:0] O0;

    // Line 790
    assign N596 = I0 == I1;
    // Line 790
    assign O0 = N596;
endmodule

module AWDP_EQ_222(O0, mul64);
    output [0:0] O0;
    input [63:32] mul64;
    // Line 131
    wire [0:0] N616;
    // Line 131
    wire [0:0] O0;

    // Line 131
    assign N616 = mul64 == 32'hffffffff;
    // Line 131
    assign O0 = N616;
endmodule

module AWDP_EQ_231(O0, mul64);
    output [0:0] O0;
    input [63:8] mul64;
    // Line 129
    wire [0:0] N625;
    // Line 129
    wire [0:0] O0;

    // Line 129
    assign N625 = mul64 == 56'hffffffff;
    // Line 129
    assign O0 = N625;
endmodule

module AWDP_GE_13(O0, divr, divq);
    output [0:0] O0;
    input [63:0] divr;
    input [63:0] divq;
    // Line 1006
    wire [0:0] N635;
    // Line 1006
    wire [0:0] O0;

    // Line 1006
    assign N635 = divr >= divq;
    // Line 1006
    assign O0 = N635;
endmodule

module AWDP_INC_11111286(O0, I0);

	output [63:0] O0;
	input [63:0] I0;




	notech_ha2 i_31(.A(I0[31]), .B(n_573), .Z(O0[31]), .CO(O0[32]));
	notech_ha2 i_30(.A(I0[30]), .B(n_571), .Z(O0[30]), .CO(n_573));
	notech_ha2 i_29(.A(I0[29]), .B(n_569), .Z(O0[29]), .CO(n_571));
	notech_ha2 i_28(.A(I0[28]), .B(n_567), .Z(O0[28]), .CO(n_569));
	notech_ha2 i_27(.A(I0[27]), .B(n_565), .Z(O0[27]), .CO(n_567));
	notech_ha2 i_26(.A(I0[26]), .B(n_563), .Z(O0[26]), .CO(n_565));
	notech_ha2 i_25(.A(I0[25]), .B(n_561), .Z(O0[25]), .CO(n_563));
	notech_ha2 i_24(.A(I0[24]), .B(n_559), .Z(O0[24]), .CO(n_561));
	notech_ha2 i_23(.A(I0[23]), .B(n_557), .Z(O0[23]), .CO(n_559));
	notech_ha2 i_22(.A(I0[22]), .B(n_555), .Z(O0[22]), .CO(n_557));
	notech_ha2 i_21(.A(I0[21]), .B(n_553), .Z(O0[21]), .CO(n_555));
	notech_ha2 i_20(.A(I0[20]), .B(n_551), .Z(O0[20]), .CO(n_553));
	notech_ha2 i_19(.A(I0[19]), .B(n_549), .Z(O0[19]), .CO(n_551));
	notech_ha2 i_18(.A(I0[18]), .B(n_547), .Z(O0[18]), .CO(n_549));
	notech_ha2 i_17(.A(I0[17]), .B(n_545), .Z(O0[17]), .CO(n_547));
	notech_ha2 i_16(.A(I0[16]), .B(n_543), .Z(O0[16]), .CO(n_545));
	notech_ha2 i_15(.A(I0[15]), .B(n_541), .Z(O0[15]), .CO(n_543));
	notech_ha2 i_14(.A(I0[14]), .B(n_539), .Z(O0[14]), .CO(n_541));
	notech_ha2 i_13(.A(I0[13]), .B(n_537), .Z(O0[13]), .CO(n_539));
	notech_ha2 i_12(.A(I0[12]), .B(n_535), .Z(O0[12]), .CO(n_537));
	notech_ha2 i_11(.A(I0[11]), .B(n_533), .Z(O0[11]), .CO(n_535));
	notech_ha2 i_10(.A(I0[10]), .B(n_531), .Z(O0[10]), .CO(n_533));
	notech_ha2 i_9(.A(I0[9]), .B(n_529), .Z(O0[9]), .CO(n_531));
	notech_ha2 i_8(.A(I0[8]), .B(n_527), .Z(O0[8]), .CO(n_529));
	notech_ha2 i_7(.A(I0[7]), .B(n_525), .Z(O0[7]), .CO(n_527));
	notech_ha2 i_6(.A(I0[6]), .B(n_523), .Z(O0[6]), .CO(n_525));
	notech_ha2 i_5(.A(I0[5]), .B(n_521), .Z(O0[5]), .CO(n_523));
	notech_ha2 i_4(.A(I0[4]), .B(n_519), .Z(O0[4]), .CO(n_521));
	notech_ha2 i_3(.A(I0[3]), .B(n_517), .Z(O0[3]), .CO(n_519));
	notech_ha2 i_2(.A(I0[2]), .B(n_515), .Z(O0[2]), .CO(n_517));
	notech_ha2 i_1(.A(I0[1]), .B(I0[0]), .Z(O0[1]), .CO(n_515));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_INC_167(O0, I0);

	output [15:0] O0;
	input [15:0] I0;




	notech_ha2 i_15(.A(I0[15]), .B(n_156), .Z(O0[15]));
	notech_ha2 i_14(.A(I0[14]), .B(n_154), .Z(O0[14]), .CO(n_156));
	notech_ha2 i_13(.A(I0[13]), .B(n_152), .Z(O0[13]), .CO(n_154));
	notech_ha2 i_12(.A(I0[12]), .B(n_150), .Z(O0[12]), .CO(n_152));
	notech_ha2 i_11(.A(I0[11]), .B(n_148), .Z(O0[11]), .CO(n_150));
	notech_ha2 i_10(.A(I0[10]), .B(n_146), .Z(O0[10]), .CO(n_148));
	notech_ha2 i_9(.A(I0[9]), .B(n_144), .Z(O0[9]), .CO(n_146));
	notech_ha2 i_8(.A(I0[8]), .B(n_142), .Z(O0[8]), .CO(n_144));
	notech_ha2 i_7(.A(I0[7]), .B(n_140), .Z(O0[7]), .CO(n_142));
	notech_ha2 i_6(.A(I0[6]), .B(n_138), .Z(O0[6]), .CO(n_140));
	notech_ha2 i_5(.A(I0[5]), .B(n_136), .Z(O0[5]), .CO(n_138));
	notech_ha2 i_4(.A(I0[4]), .B(n_134), .Z(O0[4]), .CO(n_136));
	notech_ha2 i_3(.A(I0[3]), .B(n_132), .Z(O0[3]), .CO(n_134));
	notech_ha2 i_2(.A(I0[2]), .B(n_130), .Z(O0[2]), .CO(n_132));
	notech_ha2 i_1(.A(I0[1]), .B(I0[0]), .Z(O0[1]), .CO(n_130));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_INC_183(O0, I0);

	output [31:0] O0;
	input [31:0] I0;




	notech_ha2 i_31(.A(I0[31]), .B(n_316), .Z(O0[31]));
	notech_ha2 i_30(.A(I0[30]), .B(n_314), .Z(O0[30]), .CO(n_316));
	notech_ha2 i_29(.A(I0[29]), .B(n_312), .Z(O0[29]), .CO(n_314));
	notech_ha2 i_28(.A(I0[28]), .B(n_310), .Z(O0[28]), .CO(n_312));
	notech_ha2 i_27(.A(I0[27]), .B(n_308), .Z(O0[27]), .CO(n_310));
	notech_ha2 i_26(.A(I0[26]), .B(n_306), .Z(O0[26]), .CO(n_308));
	notech_ha2 i_25(.A(I0[25]), .B(n_304), .Z(O0[25]), .CO(n_306));
	notech_ha2 i_24(.A(I0[24]), .B(n_302), .Z(O0[24]), .CO(n_304));
	notech_ha2 i_23(.A(I0[23]), .B(n_300), .Z(O0[23]), .CO(n_302));
	notech_ha2 i_22(.A(I0[22]), .B(n_298), .Z(O0[22]), .CO(n_300));
	notech_ha2 i_21(.A(I0[21]), .B(n_296), .Z(O0[21]), .CO(n_298));
	notech_ha2 i_20(.A(I0[20]), .B(n_294), .Z(O0[20]), .CO(n_296));
	notech_ha2 i_19(.A(I0[19]), .B(n_292), .Z(O0[19]), .CO(n_294));
	notech_ha2 i_18(.A(I0[18]), .B(n_290), .Z(O0[18]), .CO(n_292));
	notech_ha2 i_17(.A(I0[17]), .B(n_288), .Z(O0[17]), .CO(n_290));
	notech_ha2 i_16(.A(I0[16]), .B(n_286), .Z(O0[16]), .CO(n_288));
	notech_ha2 i_15(.A(I0[15]), .B(n_284), .Z(O0[15]), .CO(n_286));
	notech_ha2 i_14(.A(I0[14]), .B(n_282), .Z(O0[14]), .CO(n_284));
	notech_ha2 i_13(.A(I0[13]), .B(n_280), .Z(O0[13]), .CO(n_282));
	notech_ha2 i_12(.A(I0[12]), .B(n_278), .Z(O0[12]), .CO(n_280));
	notech_ha2 i_11(.A(I0[11]), .B(n_276), .Z(O0[11]), .CO(n_278));
	notech_ha2 i_10(.A(I0[10]), .B(n_274), .Z(O0[10]), .CO(n_276));
	notech_ha2 i_9(.A(I0[9]), .B(n_272), .Z(O0[9]), .CO(n_274));
	notech_ha2 i_8(.A(I0[8]), .B(n_270), .Z(O0[8]), .CO(n_272));
	notech_ha2 i_7(.A(I0[7]), .B(n_268), .Z(O0[7]), .CO(n_270));
	notech_ha2 i_6(.A(I0[6]), .B(n_266), .Z(O0[6]), .CO(n_268));
	notech_ha2 i_5(.A(I0[5]), .B(n_264), .Z(O0[5]), .CO(n_266));
	notech_ha2 i_4(.A(I0[4]), .B(n_262), .Z(O0[4]), .CO(n_264));
	notech_ha2 i_3(.A(I0[3]), .B(n_260), .Z(O0[3]), .CO(n_262));
	notech_ha2 i_2(.A(I0[2]), .B(n_258), .Z(O0[2]), .CO(n_260));
	notech_ha2 i_1(.A(I0[1]), .B(I0[0]), .Z(O0[1]), .CO(n_258));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_INC_212(O0, I0);

	output [63:0] O0;
	input [63:0] I0;




	notech_ha2 i_63(.A(I0[63]), .B(n_636), .Z(O0[63]));
	notech_ha2 i_62(.A(I0[62]), .B(n_634), .Z(O0[62]), .CO(n_636));
	notech_ha2 i_61(.A(I0[61]), .B(n_632), .Z(O0[61]), .CO(n_634));
	notech_ha2 i_60(.A(I0[60]), .B(n_630), .Z(O0[60]), .CO(n_632));
	notech_ha2 i_59(.A(I0[59]), .B(n_628), .Z(O0[59]), .CO(n_630));
	notech_ha2 i_58(.A(I0[58]), .B(n_626), .Z(O0[58]), .CO(n_628));
	notech_ha2 i_57(.A(I0[57]), .B(n_624), .Z(O0[57]), .CO(n_626));
	notech_ha2 i_56(.A(I0[56]), .B(n_622), .Z(O0[56]), .CO(n_624));
	notech_ha2 i_55(.A(I0[55]), .B(n_620), .Z(O0[55]), .CO(n_622));
	notech_ha2 i_54(.A(I0[54]), .B(n_618), .Z(O0[54]), .CO(n_620));
	notech_ha2 i_53(.A(I0[53]), .B(n_616), .Z(O0[53]), .CO(n_618));
	notech_ha2 i_52(.A(I0[52]), .B(n_614), .Z(O0[52]), .CO(n_616));
	notech_ha2 i_51(.A(I0[51]), .B(n_612), .Z(O0[51]), .CO(n_614));
	notech_ha2 i_50(.A(I0[50]), .B(n_610), .Z(O0[50]), .CO(n_612));
	notech_ha2 i_49(.A(I0[49]), .B(n_608), .Z(O0[49]), .CO(n_610));
	notech_ha2 i_48(.A(I0[48]), .B(n_606), .Z(O0[48]), .CO(n_608));
	notech_ha2 i_47(.A(I0[47]), .B(n_604), .Z(O0[47]), .CO(n_606));
	notech_ha2 i_46(.A(I0[46]), .B(n_602), .Z(O0[46]), .CO(n_604));
	notech_ha2 i_45(.A(I0[45]), .B(n_600), .Z(O0[45]), .CO(n_602));
	notech_ha2 i_44(.A(I0[44]), .B(n_598), .Z(O0[44]), .CO(n_600));
	notech_ha2 i_43(.A(I0[43]), .B(n_596), .Z(O0[43]), .CO(n_598));
	notech_ha2 i_42(.A(I0[42]), .B(n_594), .Z(O0[42]), .CO(n_596));
	notech_ha2 i_41(.A(I0[41]), .B(n_592), .Z(O0[41]), .CO(n_594));
	notech_ha2 i_40(.A(I0[40]), .B(n_590), .Z(O0[40]), .CO(n_592));
	notech_ha2 i_39(.A(I0[39]), .B(n_588), .Z(O0[39]), .CO(n_590));
	notech_ha2 i_38(.A(I0[38]), .B(n_586), .Z(O0[38]), .CO(n_588));
	notech_ha2 i_37(.A(I0[37]), .B(n_584), .Z(O0[37]), .CO(n_586));
	notech_ha2 i_36(.A(I0[36]), .B(n_582), .Z(O0[36]), .CO(n_584));
	notech_ha2 i_35(.A(I0[35]), .B(n_580), .Z(O0[35]), .CO(n_582));
	notech_ha2 i_34(.A(I0[34]), .B(n_578), .Z(O0[34]), .CO(n_580));
	notech_ha2 i_33(.A(I0[33]), .B(n_576), .Z(O0[33]), .CO(n_578));
	notech_ha2 i_32(.A(I0[32]), .B(n_574), .Z(O0[32]), .CO(n_576));
	notech_ha2 i_31(.A(I0[31]), .B(n_572), .Z(O0[31]), .CO(n_574));
	notech_ha2 i_30(.A(I0[30]), .B(n_570), .Z(O0[30]), .CO(n_572));
	notech_ha2 i_29(.A(I0[29]), .B(n_568), .Z(O0[29]), .CO(n_570));
	notech_ha2 i_28(.A(I0[28]), .B(n_566), .Z(O0[28]), .CO(n_568));
	notech_ha2 i_27(.A(I0[27]), .B(n_564), .Z(O0[27]), .CO(n_566));
	notech_ha2 i_26(.A(I0[26]), .B(n_562), .Z(O0[26]), .CO(n_564));
	notech_ha2 i_25(.A(I0[25]), .B(n_560), .Z(O0[25]), .CO(n_562));
	notech_ha2 i_24(.A(I0[24]), .B(n_558), .Z(O0[24]), .CO(n_560));
	notech_ha2 i_23(.A(I0[23]), .B(n_556), .Z(O0[23]), .CO(n_558));
	notech_ha2 i_22(.A(I0[22]), .B(n_554), .Z(O0[22]), .CO(n_556));
	notech_ha2 i_21(.A(I0[21]), .B(n_552), .Z(O0[21]), .CO(n_554));
	notech_ha2 i_20(.A(I0[20]), .B(n_550), .Z(O0[20]), .CO(n_552));
	notech_ha2 i_19(.A(I0[19]), .B(n_548), .Z(O0[19]), .CO(n_550));
	notech_ha2 i_18(.A(I0[18]), .B(n_546), .Z(O0[18]), .CO(n_548));
	notech_ha2 i_17(.A(I0[17]), .B(n_544), .Z(O0[17]), .CO(n_546));
	notech_ha2 i_16(.A(I0[16]), .B(n_542), .Z(O0[16]), .CO(n_544));
	notech_ha2 i_15(.A(I0[15]), .B(n_540), .Z(O0[15]), .CO(n_542));
	notech_ha2 i_14(.A(I0[14]), .B(n_538), .Z(O0[14]), .CO(n_540));
	notech_ha2 i_13(.A(I0[13]), .B(n_536), .Z(O0[13]), .CO(n_538));
	notech_ha2 i_12(.A(I0[12]), .B(n_534), .Z(O0[12]), .CO(n_536));
	notech_ha2 i_11(.A(I0[11]), .B(n_532), .Z(O0[11]), .CO(n_534));
	notech_ha2 i_10(.A(I0[10]), .B(n_530), .Z(O0[10]), .CO(n_532));
	notech_ha2 i_9(.A(I0[9]), .B(n_528), .Z(O0[9]), .CO(n_530));
	notech_ha2 i_8(.A(I0[8]), .B(n_526), .Z(O0[8]), .CO(n_528));
	notech_ha2 i_7(.A(I0[7]), .B(n_524), .Z(O0[7]), .CO(n_526));
	notech_ha2 i_6(.A(I0[6]), .B(n_522), .Z(O0[6]), .CO(n_524));
	notech_ha2 i_5(.A(I0[5]), .B(n_520), .Z(O0[5]), .CO(n_522));
	notech_ha2 i_4(.A(I0[4]), .B(n_518), .Z(O0[4]), .CO(n_520));
	notech_ha2 i_3(.A(I0[3]), .B(n_516), .Z(O0[3]), .CO(n_518));
	notech_ha2 i_2(.A(I0[2]), .B(n_514), .Z(O0[2]), .CO(n_516));
	notech_ha2 i_1(.A(I0[1]), .B(I0[0]), .Z(O0[1]), .CO(n_514));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_INC_232(O0, tsc);

	output [63:0] O0;
	input [63:0] tsc;




	notech_ha2 i_63(.A(tsc[63]), .B(n_636), .Z(O0[63]));
	notech_ha2 i_62(.A(tsc[62]), .B(n_634), .Z(O0[62]), .CO(n_636));
	notech_ha2 i_61(.A(tsc[61]), .B(n_632), .Z(O0[61]), .CO(n_634));
	notech_ha2 i_60(.A(tsc[60]), .B(n_630), .Z(O0[60]), .CO(n_632));
	notech_ha2 i_59(.A(tsc[59]), .B(n_628), .Z(O0[59]), .CO(n_630));
	notech_ha2 i_58(.A(tsc[58]), .B(n_626), .Z(O0[58]), .CO(n_628));
	notech_ha2 i_57(.A(tsc[57]), .B(n_624), .Z(O0[57]), .CO(n_626));
	notech_ha2 i_56(.A(tsc[56]), .B(n_622), .Z(O0[56]), .CO(n_624));
	notech_ha2 i_55(.A(tsc[55]), .B(n_620), .Z(O0[55]), .CO(n_622));
	notech_ha2 i_54(.A(tsc[54]), .B(n_618), .Z(O0[54]), .CO(n_620));
	notech_ha2 i_53(.A(tsc[53]), .B(n_616), .Z(O0[53]), .CO(n_618));
	notech_ha2 i_52(.A(tsc[52]), .B(n_614), .Z(O0[52]), .CO(n_616));
	notech_ha2 i_51(.A(tsc[51]), .B(n_612), .Z(O0[51]), .CO(n_614));
	notech_ha2 i_50(.A(tsc[50]), .B(n_610), .Z(O0[50]), .CO(n_612));
	notech_ha2 i_49(.A(tsc[49]), .B(n_608), .Z(O0[49]), .CO(n_610));
	notech_ha2 i_48(.A(tsc[48]), .B(n_606), .Z(O0[48]), .CO(n_608));
	notech_ha2 i_47(.A(tsc[47]), .B(n_604), .Z(O0[47]), .CO(n_606));
	notech_ha2 i_46(.A(tsc[46]), .B(n_602), .Z(O0[46]), .CO(n_604));
	notech_ha2 i_45(.A(tsc[45]), .B(n_600), .Z(O0[45]), .CO(n_602));
	notech_ha2 i_44(.A(tsc[44]), .B(n_598), .Z(O0[44]), .CO(n_600));
	notech_ha2 i_43(.A(tsc[43]), .B(n_596), .Z(O0[43]), .CO(n_598));
	notech_ha2 i_42(.A(tsc[42]), .B(n_594), .Z(O0[42]), .CO(n_596));
	notech_ha2 i_41(.A(tsc[41]), .B(n_592), .Z(O0[41]), .CO(n_594));
	notech_ha2 i_40(.A(tsc[40]), .B(n_590), .Z(O0[40]), .CO(n_592));
	notech_ha2 i_39(.A(tsc[39]), .B(n_588), .Z(O0[39]), .CO(n_590));
	notech_ha2 i_38(.A(tsc[38]), .B(n_586), .Z(O0[38]), .CO(n_588));
	notech_ha2 i_37(.A(tsc[37]), .B(n_584), .Z(O0[37]), .CO(n_586));
	notech_ha2 i_36(.A(tsc[36]), .B(n_582), .Z(O0[36]), .CO(n_584));
	notech_ha2 i_35(.A(tsc[35]), .B(n_580), .Z(O0[35]), .CO(n_582));
	notech_ha2 i_34(.A(tsc[34]), .B(n_578), .Z(O0[34]), .CO(n_580));
	notech_ha2 i_33(.A(tsc[33]), .B(n_576), .Z(O0[33]), .CO(n_578));
	notech_ha2 i_32(.A(tsc[32]), .B(n_574), .Z(O0[32]), .CO(n_576));
	notech_ha2 i_31(.A(tsc[31]), .B(n_572), .Z(O0[31]), .CO(n_574));
	notech_ha2 i_30(.A(tsc[30]), .B(n_570), .Z(O0[30]), .CO(n_572));
	notech_ha2 i_29(.A(tsc[29]), .B(n_568), .Z(O0[29]), .CO(n_570));
	notech_ha2 i_28(.A(tsc[28]), .B(n_566), .Z(O0[28]), .CO(n_568));
	notech_ha2 i_27(.A(tsc[27]), .B(n_564), .Z(O0[27]), .CO(n_566));
	notech_ha2 i_26(.A(tsc[26]), .B(n_562), .Z(O0[26]), .CO(n_564));
	notech_ha2 i_25(.A(tsc[25]), .B(n_560), .Z(O0[25]), .CO(n_562));
	notech_ha2 i_24(.A(tsc[24]), .B(n_558), .Z(O0[24]), .CO(n_560));
	notech_ha2 i_23(.A(tsc[23]), .B(n_556), .Z(O0[23]), .CO(n_558));
	notech_ha2 i_22(.A(tsc[22]), .B(n_554), .Z(O0[22]), .CO(n_556));
	notech_ha2 i_21(.A(tsc[21]), .B(n_552), .Z(O0[21]), .CO(n_554));
	notech_ha2 i_20(.A(tsc[20]), .B(n_550), .Z(O0[20]), .CO(n_552));
	notech_ha2 i_19(.A(tsc[19]), .B(n_548), .Z(O0[19]), .CO(n_550));
	notech_ha2 i_18(.A(tsc[18]), .B(n_546), .Z(O0[18]), .CO(n_548));
	notech_ha2 i_17(.A(tsc[17]), .B(n_544), .Z(O0[17]), .CO(n_546));
	notech_ha2 i_16(.A(tsc[16]), .B(n_542), .Z(O0[16]), .CO(n_544));
	notech_ha2 i_15(.A(tsc[15]), .B(n_540), .Z(O0[15]), .CO(n_542));
	notech_ha2 i_14(.A(tsc[14]), .B(n_538), .Z(O0[14]), .CO(n_540));
	notech_ha2 i_13(.A(tsc[13]), .B(n_536), .Z(O0[13]), .CO(n_538));
	notech_ha2 i_12(.A(tsc[12]), .B(n_534), .Z(O0[12]), .CO(n_536));
	notech_ha2 i_11(.A(tsc[11]), .B(n_532), .Z(O0[11]), .CO(n_534));
	notech_ha2 i_10(.A(tsc[10]), .B(n_530), .Z(O0[10]), .CO(n_532));
	notech_ha2 i_9(.A(tsc[9]), .B(n_528), .Z(O0[9]), .CO(n_530));
	notech_ha2 i_8(.A(tsc[8]), .B(n_526), .Z(O0[8]), .CO(n_528));
	notech_ha2 i_7(.A(tsc[7]), .B(n_524), .Z(O0[7]), .CO(n_526));
	notech_ha2 i_6(.A(tsc[6]), .B(n_522), .Z(O0[6]), .CO(n_524));
	notech_ha2 i_5(.A(tsc[5]), .B(n_520), .Z(O0[5]), .CO(n_522));
	notech_ha2 i_4(.A(tsc[4]), .B(n_518), .Z(O0[4]), .CO(n_520));
	notech_ha2 i_3(.A(tsc[3]), .B(n_516), .Z(O0[3]), .CO(n_518));
	notech_ha2 i_2(.A(tsc[2]), .B(n_514), .Z(O0[2]), .CO(n_516));
	notech_ha2 i_1(.A(tsc[1]), .B(tsc[0]), .Z(O0[1]), .CO(n_514));
	notech_inv i_0(.A(tsc[0]), .Z(O0[0]));
endmodule
module AWDP_INC_28(O0, I0);

	output [31:0] O0;
	input [31:0] I0;




	notech_ha2 i_31(.A(I0[31]), .B(n_316), .Z(O0[31]));
	notech_ha2 i_30(.A(I0[30]), .B(n_314), .Z(O0[30]), .CO(n_316));
	notech_ha2 i_29(.A(I0[29]), .B(n_312), .Z(O0[29]), .CO(n_314));
	notech_ha2 i_28(.A(I0[28]), .B(n_310), .Z(O0[28]), .CO(n_312));
	notech_ha2 i_27(.A(I0[27]), .B(n_308), .Z(O0[27]), .CO(n_310));
	notech_ha2 i_26(.A(I0[26]), .B(n_306), .Z(O0[26]), .CO(n_308));
	notech_ha2 i_25(.A(I0[25]), .B(n_304), .Z(O0[25]), .CO(n_306));
	notech_ha2 i_24(.A(I0[24]), .B(n_302), .Z(O0[24]), .CO(n_304));
	notech_ha2 i_23(.A(I0[23]), .B(n_300), .Z(O0[23]), .CO(n_302));
	notech_ha2 i_22(.A(I0[22]), .B(n_298), .Z(O0[22]), .CO(n_300));
	notech_ha2 i_21(.A(I0[21]), .B(n_296), .Z(O0[21]), .CO(n_298));
	notech_ha2 i_20(.A(I0[20]), .B(n_294), .Z(O0[20]), .CO(n_296));
	notech_ha2 i_19(.A(I0[19]), .B(n_292), .Z(O0[19]), .CO(n_294));
	notech_ha2 i_18(.A(I0[18]), .B(n_290), .Z(O0[18]), .CO(n_292));
	notech_ha2 i_17(.A(I0[17]), .B(n_288), .Z(O0[17]), .CO(n_290));
	notech_ha2 i_16(.A(I0[16]), .B(n_286), .Z(O0[16]), .CO(n_288));
	notech_ha2 i_15(.A(I0[15]), .B(n_284), .Z(O0[15]), .CO(n_286));
	notech_ha2 i_14(.A(I0[14]), .B(n_282), .Z(O0[14]), .CO(n_284));
	notech_ha2 i_13(.A(I0[13]), .B(n_280), .Z(O0[13]), .CO(n_282));
	notech_ha2 i_12(.A(I0[12]), .B(n_278), .Z(O0[12]), .CO(n_280));
	notech_ha2 i_11(.A(I0[11]), .B(n_276), .Z(O0[11]), .CO(n_278));
	notech_ha2 i_10(.A(I0[10]), .B(n_274), .Z(O0[10]), .CO(n_276));
	notech_ha2 i_9(.A(I0[9]), .B(n_272), .Z(O0[9]), .CO(n_274));
	notech_ha2 i_8(.A(I0[8]), .B(n_270), .Z(O0[8]), .CO(n_272));
	notech_ha2 i_7(.A(I0[7]), .B(n_268), .Z(O0[7]), .CO(n_270));
	notech_ha2 i_6(.A(I0[6]), .B(n_266), .Z(O0[6]), .CO(n_268));
	notech_ha2 i_5(.A(I0[5]), .B(n_264), .Z(O0[5]), .CO(n_266));
	notech_ha2 i_4(.A(I0[4]), .B(n_262), .Z(O0[4]), .CO(n_264));
	notech_ha2 i_3(.A(I0[3]), .B(n_260), .Z(O0[3]), .CO(n_262));
	notech_ha2 i_2(.A(I0[2]), .B(n_258), .Z(O0[2]), .CO(n_260));
	notech_ha2 i_1(.A(I0[1]), .B(I0[0]), .Z(O0[1]), .CO(n_258));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_INC_91(O0, I0);

	output [31:0] O0;
	input [31:0] I0;




	notech_ha2 i_31(.A(I0[31]), .B(n_316), .Z(O0[31]));
	notech_ha2 i_30(.A(I0[30]), .B(n_314), .Z(O0[30]), .CO(n_316));
	notech_ha2 i_29(.A(I0[29]), .B(n_312), .Z(O0[29]), .CO(n_314));
	notech_ha2 i_28(.A(I0[28]), .B(n_310), .Z(O0[28]), .CO(n_312));
	notech_ha2 i_27(.A(I0[27]), .B(n_308), .Z(O0[27]), .CO(n_310));
	notech_ha2 i_26(.A(I0[26]), .B(n_306), .Z(O0[26]), .CO(n_308));
	notech_ha2 i_25(.A(I0[25]), .B(n_304), .Z(O0[25]), .CO(n_306));
	notech_ha2 i_24(.A(I0[24]), .B(n_302), .Z(O0[24]), .CO(n_304));
	notech_ha2 i_23(.A(I0[23]), .B(n_300), .Z(O0[23]), .CO(n_302));
	notech_ha2 i_22(.A(I0[22]), .B(n_298), .Z(O0[22]), .CO(n_300));
	notech_ha2 i_21(.A(I0[21]), .B(n_296), .Z(O0[21]), .CO(n_298));
	notech_ha2 i_20(.A(I0[20]), .B(n_294), .Z(O0[20]), .CO(n_296));
	notech_ha2 i_19(.A(I0[19]), .B(n_292), .Z(O0[19]), .CO(n_294));
	notech_ha2 i_18(.A(I0[18]), .B(n_290), .Z(O0[18]), .CO(n_292));
	notech_ha2 i_17(.A(I0[17]), .B(n_288), .Z(O0[17]), .CO(n_290));
	notech_ha2 i_16(.A(I0[16]), .B(n_286), .Z(O0[16]), .CO(n_288));
	notech_ha2 i_15(.A(I0[15]), .B(n_284), .Z(O0[15]), .CO(n_286));
	notech_ha2 i_14(.A(I0[14]), .B(n_282), .Z(O0[14]), .CO(n_284));
	notech_ha2 i_13(.A(I0[13]), .B(n_280), .Z(O0[13]), .CO(n_282));
	notech_ha2 i_12(.A(I0[12]), .B(n_278), .Z(O0[12]), .CO(n_280));
	notech_ha2 i_11(.A(I0[11]), .B(n_276), .Z(O0[11]), .CO(n_278));
	notech_ha2 i_10(.A(I0[10]), .B(n_274), .Z(O0[10]), .CO(n_276));
	notech_ha2 i_9(.A(I0[9]), .B(n_272), .Z(O0[9]), .CO(n_274));
	notech_ha2 i_8(.A(I0[8]), .B(n_270), .Z(O0[8]), .CO(n_272));
	notech_ha2 i_7(.A(I0[7]), .B(n_268), .Z(O0[7]), .CO(n_270));
	notech_ha2 i_6(.A(I0[6]), .B(n_266), .Z(O0[6]), .CO(n_268));
	notech_ha2 i_5(.A(I0[5]), .B(n_264), .Z(O0[5]), .CO(n_266));
	notech_ha2 i_4(.A(I0[4]), .B(n_262), .Z(O0[4]), .CO(n_264));
	notech_ha2 i_3(.A(I0[3]), .B(n_260), .Z(O0[3]), .CO(n_262));
	notech_ha2 i_2(.A(I0[2]), .B(n_258), .Z(O0[2]), .CO(n_260));
	notech_ha2 i_1(.A(I0[1]), .B(I0[0]), .Z(O0[1]), .CO(n_258));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_LE_215(O0, divq, I0);

	output [0:0] O0;
	input [63:0] divq;
	input [63:0] I0;




	notech_inv i_320(.A(n_710), .Z(O0[0]));
	notech_nand2 i_317(.A(n_703), .B(n_709), .Z(n_710));
	notech_inv i_506(.A(n_835), .Z(n_703));
	notech_or2 i_505(.A(n_834), .B(n_701), .Z(n_835));
	notech_and2 i_504(.A(n_702), .B(n_700), .Z(n_834));
	notech_inv i_315(.A(n_512), .Z(n_702));
	notech_inv i_314(.A(n_577), .Z(n_701));
	notech_inv i_503(.A(n_928), .Z(n_700));
	notech_nor2 i_502(.A(n_927), .B(n_866), .Z(n_928));
	notech_nor2 i_501(.A(n_699), .B(n_511), .Z(n_927));
	notech_inv i_500(.A(n_831), .Z(n_699));
	notech_or2 i_499(.A(n_830), .B(n_697), .Z(n_831));
	notech_and2 i_498(.A(n_698), .B(n_696), .Z(n_830));
	notech_inv i_311(.A(n_510), .Z(n_698));
	notech_inv i_310(.A(n_575), .Z(n_697));
	notech_inv i_497(.A(n_926), .Z(n_696));
	notech_nor2 i_496(.A(n_925), .B(n_865), .Z(n_926));
	notech_nor2 i_495(.A(n_695), .B(n_509), .Z(n_925));
	notech_inv i_494(.A(n_827), .Z(n_695));
	notech_or2 i_493(.A(n_826), .B(n_693), .Z(n_827));
	notech_and2 i_492(.A(n_694), .B(n_692), .Z(n_826));
	notech_inv i_307(.A(n_508), .Z(n_694));
	notech_inv i_306(.A(n_573), .Z(n_693));
	notech_inv i_491(.A(n_924), .Z(n_692));
	notech_nor2 i_490(.A(n_923), .B(n_864), .Z(n_924));
	notech_nor2 i_489(.A(n_691), .B(n_507), .Z(n_923));
	notech_inv i_488(.A(n_823), .Z(n_691));
	notech_or2 i_487(.A(n_822), .B(n_689), .Z(n_823));
	notech_and2 i_486(.A(n_690), .B(n_688), .Z(n_822));
	notech_inv i_303(.A(n_506), .Z(n_690));
	notech_inv i_302(.A(n_571), .Z(n_689));
	notech_inv i_485(.A(n_922), .Z(n_688));
	notech_nor2 i_484(.A(n_921), .B(n_863), .Z(n_922));
	notech_nor2 i_483(.A(n_687), .B(n_505), .Z(n_921));
	notech_inv i_482(.A(n_819), .Z(n_687));
	notech_or2 i_481(.A(n_818), .B(n_685), .Z(n_819));
	notech_and2 i_480(.A(n_686), .B(n_684), .Z(n_818));
	notech_inv i_299(.A(n_504), .Z(n_686));
	notech_inv i_298(.A(n_569), .Z(n_685));
	notech_inv i_479(.A(n_920), .Z(n_684));
	notech_nor2 i_478(.A(n_919), .B(n_862), .Z(n_920));
	notech_nor2 i_477(.A(n_683), .B(n_503), .Z(n_919));
	notech_inv i_476(.A(n_815), .Z(n_683));
	notech_or2 i_475(.A(n_814), .B(n_681), .Z(n_815));
	notech_and2 i_474(.A(n_682), .B(n_680), .Z(n_814));
	notech_inv i_295(.A(n_502), .Z(n_682));
	notech_inv i_294(.A(n_567), .Z(n_681));
	notech_inv i_473(.A(n_918), .Z(n_680));
	notech_nor2 i_472(.A(n_917), .B(n_861), .Z(n_918));
	notech_nor2 i_471(.A(n_679), .B(n_501), .Z(n_917));
	notech_inv i_470(.A(n_811), .Z(n_679));
	notech_or2 i_469(.A(n_810), .B(n_677), .Z(n_811));
	notech_and2 i_468(.A(n_678), .B(n_676), .Z(n_810));
	notech_inv i_291(.A(n_500), .Z(n_678));
	notech_inv i_290(.A(n_565), .Z(n_677));
	notech_inv i_467(.A(n_916), .Z(n_676));
	notech_nor2 i_466(.A(n_915), .B(n_860), .Z(n_916));
	notech_nor2 i_465(.A(n_675), .B(n_499), .Z(n_915));
	notech_inv i_464(.A(n_807), .Z(n_675));
	notech_or2 i_463(.A(n_806), .B(n_673), .Z(n_807));
	notech_and2 i_462(.A(n_674), .B(n_672), .Z(n_806));
	notech_inv i_287(.A(n_498), .Z(n_674));
	notech_inv i_286(.A(n_563), .Z(n_673));
	notech_inv i_461(.A(n_914), .Z(n_672));
	notech_nor2 i_460(.A(n_913), .B(n_859), .Z(n_914));
	notech_nor2 i_459(.A(n_671), .B(n_497), .Z(n_913));
	notech_inv i_458(.A(n_803), .Z(n_671));
	notech_or2 i_457(.A(n_802), .B(n_669), .Z(n_803));
	notech_and2 i_456(.A(n_670), .B(n_668), .Z(n_802));
	notech_inv i_283(.A(n_496), .Z(n_670));
	notech_inv i_282(.A(n_561), .Z(n_669));
	notech_inv i_455(.A(n_912), .Z(n_668));
	notech_nor2 i_454(.A(n_911), .B(n_858), .Z(n_912));
	notech_nor2 i_453(.A(n_667), .B(n_495), .Z(n_911));
	notech_inv i_452(.A(n_799), .Z(n_667));
	notech_or2 i_451(.A(n_798), .B(n_665), .Z(n_799));
	notech_and2 i_450(.A(n_666), .B(n_664), .Z(n_798));
	notech_inv i_279(.A(n_494), .Z(n_666));
	notech_inv i_278(.A(n_559), .Z(n_665));
	notech_inv i_449(.A(n_910), .Z(n_664));
	notech_nor2 i_448(.A(n_909), .B(n_857), .Z(n_910));
	notech_nor2 i_447(.A(n_663), .B(n_493), .Z(n_909));
	notech_inv i_446(.A(n_795), .Z(n_663));
	notech_or2 i_445(.A(n_794), .B(n_661), .Z(n_795));
	notech_and2 i_444(.A(n_662), .B(n_660), .Z(n_794));
	notech_inv i_275(.A(n_492), .Z(n_662));
	notech_inv i_274(.A(n_557), .Z(n_661));
	notech_inv i_443(.A(n_908), .Z(n_660));
	notech_nor2 i_442(.A(n_907), .B(n_856), .Z(n_908));
	notech_nor2 i_441(.A(n_659), .B(n_491), .Z(n_907));
	notech_inv i_440(.A(n_791), .Z(n_659));
	notech_or2 i_439(.A(n_790), .B(n_657), .Z(n_791));
	notech_and2 i_438(.A(n_658), .B(n_656), .Z(n_790));
	notech_inv i_271(.A(n_490), .Z(n_658));
	notech_inv i_270(.A(n_555), .Z(n_657));
	notech_inv i_437(.A(n_906), .Z(n_656));
	notech_nor2 i_436(.A(n_905), .B(n_855), .Z(n_906));
	notech_nor2 i_435(.A(n_655), .B(n_489), .Z(n_905));
	notech_inv i_434(.A(n_787), .Z(n_655));
	notech_or2 i_433(.A(n_786), .B(n_653), .Z(n_787));
	notech_and2 i_432(.A(n_654), .B(n_652), .Z(n_786));
	notech_inv i_267(.A(n_488), .Z(n_654));
	notech_inv i_266(.A(n_553), .Z(n_653));
	notech_inv i_431(.A(n_904), .Z(n_652));
	notech_nor2 i_430(.A(n_903), .B(n_854), .Z(n_904));
	notech_nor2 i_429(.A(n_651), .B(n_487), .Z(n_903));
	notech_inv i_428(.A(n_783), .Z(n_651));
	notech_or2 i_427(.A(n_782), .B(n_649), .Z(n_783));
	notech_and2 i_426(.A(n_650), .B(n_648), .Z(n_782));
	notech_inv i_263(.A(n_486), .Z(n_650));
	notech_inv i_262(.A(n_551), .Z(n_649));
	notech_inv i_425(.A(n_902), .Z(n_648));
	notech_nor2 i_424(.A(n_901), .B(n_853), .Z(n_902));
	notech_nor2 i_423(.A(n_647), .B(n_485), .Z(n_901));
	notech_inv i_422(.A(n_779), .Z(n_647));
	notech_or2 i_421(.A(n_778), .B(n_645), .Z(n_779));
	notech_and2 i_420(.A(n_646), .B(n_644), .Z(n_778));
	notech_inv i_259(.A(n_484), .Z(n_646));
	notech_inv i_258(.A(n_549), .Z(n_645));
	notech_inv i_419(.A(n_900), .Z(n_644));
	notech_nor2 i_418(.A(n_899), .B(n_852), .Z(n_900));
	notech_nor2 i_417(.A(n_643), .B(n_483), .Z(n_899));
	notech_inv i_416(.A(n_775), .Z(n_643));
	notech_or2 i_415(.A(n_774), .B(n_641), .Z(n_775));
	notech_and2 i_414(.A(n_642), .B(n_640), .Z(n_774));
	notech_inv i_255(.A(n_482), .Z(n_642));
	notech_inv i_254(.A(n_547), .Z(n_641));
	notech_inv i_413(.A(n_898), .Z(n_640));
	notech_nor2 i_412(.A(n_897), .B(n_851), .Z(n_898));
	notech_nor2 i_411(.A(n_639), .B(n_481), .Z(n_897));
	notech_inv i_410(.A(n_771), .Z(n_639));
	notech_or2 i_409(.A(n_770), .B(n_637), .Z(n_771));
	notech_and2 i_408(.A(n_638), .B(n_636), .Z(n_770));
	notech_inv i_251(.A(n_480), .Z(n_638));
	notech_inv i_250(.A(n_545), .Z(n_637));
	notech_inv i_407(.A(n_896), .Z(n_636));
	notech_nor2 i_406(.A(n_895), .B(n_850), .Z(n_896));
	notech_nor2 i_405(.A(n_635), .B(n_479), .Z(n_895));
	notech_inv i_404(.A(n_767), .Z(n_635));
	notech_or2 i_403(.A(n_766), .B(n_633), .Z(n_767));
	notech_and2 i_402(.A(n_634), .B(n_632), .Z(n_766));
	notech_inv i_247(.A(n_478), .Z(n_634));
	notech_inv i_246(.A(n_543), .Z(n_633));
	notech_inv i_401(.A(n_894), .Z(n_632));
	notech_nor2 i_400(.A(n_893), .B(n_849), .Z(n_894));
	notech_nor2 i_399(.A(n_631), .B(n_477), .Z(n_893));
	notech_inv i_398(.A(n_763), .Z(n_631));
	notech_or2 i_397(.A(n_762), .B(n_629), .Z(n_763));
	notech_and2 i_396(.A(n_630), .B(n_628), .Z(n_762));
	notech_inv i_243(.A(n_476), .Z(n_630));
	notech_inv i_242(.A(n_541), .Z(n_629));
	notech_inv i_395(.A(n_892), .Z(n_628));
	notech_nor2 i_394(.A(n_891), .B(n_848), .Z(n_892));
	notech_nor2 i_393(.A(n_627), .B(n_475), .Z(n_891));
	notech_inv i_392(.A(n_759), .Z(n_627));
	notech_or2 i_391(.A(n_758), .B(n_625), .Z(n_759));
	notech_and2 i_390(.A(n_626), .B(n_624), .Z(n_758));
	notech_inv i_239(.A(n_474), .Z(n_626));
	notech_inv i_238(.A(n_539), .Z(n_625));
	notech_inv i_389(.A(n_890), .Z(n_624));
	notech_nor2 i_388(.A(n_889), .B(n_847), .Z(n_890));
	notech_nor2 i_387(.A(n_623), .B(n_473), .Z(n_889));
	notech_inv i_386(.A(n_755), .Z(n_623));
	notech_or2 i_385(.A(n_754), .B(n_621), .Z(n_755));
	notech_and2 i_384(.A(n_622), .B(n_620), .Z(n_754));
	notech_inv i_235(.A(n_472), .Z(n_622));
	notech_inv i_234(.A(n_537), .Z(n_621));
	notech_inv i_383(.A(n_888), .Z(n_620));
	notech_nor2 i_382(.A(n_887), .B(n_846), .Z(n_888));
	notech_nor2 i_381(.A(n_619), .B(n_471), .Z(n_887));
	notech_inv i_380(.A(n_751), .Z(n_619));
	notech_or2 i_379(.A(n_750), .B(n_617), .Z(n_751));
	notech_and2 i_378(.A(n_618), .B(n_616), .Z(n_750));
	notech_inv i_231(.A(n_470), .Z(n_618));
	notech_inv i_230(.A(n_535), .Z(n_617));
	notech_inv i_377(.A(n_886), .Z(n_616));
	notech_nor2 i_376(.A(n_885), .B(n_845), .Z(n_886));
	notech_nor2 i_375(.A(n_615), .B(n_469), .Z(n_885));
	notech_inv i_374(.A(n_747), .Z(n_615));
	notech_or2 i_373(.A(n_746), .B(n_613), .Z(n_747));
	notech_and2 i_372(.A(n_614), .B(n_612), .Z(n_746));
	notech_inv i_227(.A(n_468), .Z(n_614));
	notech_inv i_226(.A(n_533), .Z(n_613));
	notech_inv i_371(.A(n_884), .Z(n_612));
	notech_nor2 i_370(.A(n_883), .B(n_844), .Z(n_884));
	notech_nor2 i_369(.A(n_611), .B(n_467), .Z(n_883));
	notech_inv i_368(.A(n_743), .Z(n_611));
	notech_or2 i_367(.A(n_742), .B(n_609), .Z(n_743));
	notech_and2 i_366(.A(n_610), .B(n_608), .Z(n_742));
	notech_inv i_223(.A(n_466), .Z(n_610));
	notech_inv i_222(.A(n_531), .Z(n_609));
	notech_inv i_365(.A(n_882), .Z(n_608));
	notech_nor2 i_364(.A(n_881), .B(n_843), .Z(n_882));
	notech_nor2 i_363(.A(n_607), .B(n_465), .Z(n_881));
	notech_inv i_362(.A(n_739), .Z(n_607));
	notech_or2 i_361(.A(n_738), .B(n_605), .Z(n_739));
	notech_and2 i_360(.A(n_606), .B(n_604), .Z(n_738));
	notech_inv i_219(.A(n_464), .Z(n_606));
	notech_inv i_218(.A(n_529), .Z(n_605));
	notech_inv i_359(.A(n_880), .Z(n_604));
	notech_nor2 i_358(.A(n_879), .B(n_842), .Z(n_880));
	notech_nor2 i_357(.A(n_603), .B(n_463), .Z(n_879));
	notech_inv i_356(.A(n_735), .Z(n_603));
	notech_or2 i_355(.A(n_734), .B(n_601), .Z(n_735));
	notech_and2 i_354(.A(n_602), .B(n_600), .Z(n_734));
	notech_inv i_215(.A(n_462), .Z(n_602));
	notech_inv i_214(.A(n_527), .Z(n_601));
	notech_inv i_353(.A(n_878), .Z(n_600));
	notech_nor2 i_352(.A(n_877), .B(n_841), .Z(n_878));
	notech_nor2 i_351(.A(n_599), .B(n_461), .Z(n_877));
	notech_inv i_350(.A(n_731), .Z(n_599));
	notech_or2 i_349(.A(n_730), .B(n_597), .Z(n_731));
	notech_and2 i_348(.A(n_598), .B(n_596), .Z(n_730));
	notech_inv i_211(.A(n_460), .Z(n_598));
	notech_inv i_210(.A(n_525), .Z(n_597));
	notech_inv i_347(.A(n_876), .Z(n_596));
	notech_nor2 i_346(.A(n_875), .B(n_840), .Z(n_876));
	notech_nor2 i_345(.A(n_595), .B(n_459), .Z(n_875));
	notech_inv i_344(.A(n_727), .Z(n_595));
	notech_or2 i_343(.A(n_726), .B(n_593), .Z(n_727));
	notech_and2 i_342(.A(n_594), .B(n_592), .Z(n_726));
	notech_inv i_207(.A(n_458), .Z(n_594));
	notech_inv i_206(.A(n_523), .Z(n_593));
	notech_inv i_341(.A(n_874), .Z(n_592));
	notech_nor2 i_340(.A(n_873), .B(n_839), .Z(n_874));
	notech_nor2 i_339(.A(n_591), .B(n_457), .Z(n_873));
	notech_inv i_338(.A(n_723), .Z(n_591));
	notech_or2 i_337(.A(n_722), .B(n_589), .Z(n_723));
	notech_and2 i_336(.A(n_590), .B(n_588), .Z(n_722));
	notech_inv i_203(.A(n_456), .Z(n_590));
	notech_inv i_202(.A(n_521), .Z(n_589));
	notech_inv i_335(.A(n_872), .Z(n_588));
	notech_nor2 i_334(.A(n_871), .B(n_838), .Z(n_872));
	notech_nor2 i_333(.A(n_587), .B(n_455), .Z(n_871));
	notech_inv i_332(.A(n_719), .Z(n_587));
	notech_or2 i_331(.A(n_718), .B(n_585), .Z(n_719));
	notech_and2 i_330(.A(n_586), .B(n_584), .Z(n_718));
	notech_inv i_199(.A(n_454), .Z(n_586));
	notech_inv i_198(.A(n_519), .Z(n_585));
	notech_inv i_329(.A(n_870), .Z(n_584));
	notech_nor2 i_328(.A(n_869), .B(n_837), .Z(n_870));
	notech_nor2 i_327(.A(n_583), .B(n_453), .Z(n_869));
	notech_inv i_326(.A(n_715), .Z(n_583));
	notech_or2 i_325(.A(n_714), .B(n_581), .Z(n_715));
	notech_and2 i_324(.A(n_582), .B(n_580), .Z(n_714));
	notech_inv i_195(.A(n_452), .Z(n_582));
	notech_inv i_194(.A(n_517), .Z(n_581));
	notech_inv i_323(.A(n_868), .Z(n_580));
	notech_nor2 i_322(.A(n_867), .B(n_836), .Z(n_868));
	notech_nor2 i_321(.A(n_451), .B(n_515), .Z(n_867));
	notech_inv i_191(.A(divq[63]), .Z(n_709));
	notech_nand2 i_190(.A(n_449), .B(divq[62]), .Z(n_577));
	notech_and2 i_189(.A(n_448), .B(divq[61]), .Z(n_866));
	notech_nand2 i_188(.A(n_447), .B(divq[60]), .Z(n_575));
	notech_and2 i_187(.A(n_446), .B(divq[59]), .Z(n_865));
	notech_nand2 i_186(.A(n_445), .B(divq[58]), .Z(n_573));
	notech_and2 i_185(.A(n_444), .B(divq[57]), .Z(n_864));
	notech_nand2 i_184(.A(n_443), .B(divq[56]), .Z(n_571));
	notech_and2 i_183(.A(n_442), .B(divq[55]), .Z(n_863));
	notech_nand2 i_182(.A(n_441), .B(divq[54]), .Z(n_569));
	notech_and2 i_181(.A(n_440), .B(divq[53]), .Z(n_862));
	notech_nand2 i_180(.A(n_439), .B(divq[52]), .Z(n_567));
	notech_and2 i_179(.A(n_438), .B(divq[51]), .Z(n_861));
	notech_nand2 i_178(.A(n_437), .B(divq[50]), .Z(n_565));
	notech_and2 i_177(.A(n_436), .B(divq[49]), .Z(n_860));
	notech_nand2 i_176(.A(n_435), .B(divq[48]), .Z(n_563));
	notech_and2 i_175(.A(n_434), .B(divq[47]), .Z(n_859));
	notech_nand2 i_174(.A(n_433), .B(divq[46]), .Z(n_561));
	notech_and2 i_173(.A(n_432), .B(divq[45]), .Z(n_858));
	notech_nand2 i_172(.A(n_431), .B(divq[44]), .Z(n_559));
	notech_and2 i_171(.A(n_430), .B(divq[43]), .Z(n_857));
	notech_nand2 i_170(.A(n_429), .B(divq[42]), .Z(n_557));
	notech_and2 i_169(.A(n_428), .B(divq[41]), .Z(n_856));
	notech_nand2 i_168(.A(n_427), .B(divq[40]), .Z(n_555));
	notech_and2 i_167(.A(n_426), .B(divq[39]), .Z(n_855));
	notech_nand2 i_166(.A(n_425), .B(divq[38]), .Z(n_553));
	notech_and2 i_165(.A(n_424), .B(divq[37]), .Z(n_854));
	notech_nand2 i_164(.A(n_423), .B(divq[36]), .Z(n_551));
	notech_and2 i_163(.A(n_422), .B(divq[35]), .Z(n_853));
	notech_nand2 i_162(.A(n_421), .B(divq[34]), .Z(n_549));
	notech_and2 i_161(.A(n_420), .B(divq[33]), .Z(n_852));
	notech_nand2 i_160(.A(n_419), .B(divq[32]), .Z(n_547));
	notech_and2 i_159(.A(n_418), .B(divq[31]), .Z(n_851));
	notech_nand2 i_158(.A(n_417), .B(divq[30]), .Z(n_545));
	notech_and2 i_157(.A(n_416), .B(divq[29]), .Z(n_850));
	notech_nand2 i_156(.A(n_415), .B(divq[28]), .Z(n_543));
	notech_and2 i_155(.A(n_414), .B(divq[27]), .Z(n_849));
	notech_nand2 i_154(.A(n_413), .B(divq[26]), .Z(n_541));
	notech_and2 i_153(.A(n_412), .B(divq[25]), .Z(n_848));
	notech_nand2 i_152(.A(n_411), .B(divq[24]), .Z(n_539));
	notech_and2 i_151(.A(n_410), .B(divq[23]), .Z(n_847));
	notech_nand2 i_150(.A(n_409), .B(divq[22]), .Z(n_537));
	notech_and2 i_149(.A(n_408), .B(divq[21]), .Z(n_846));
	notech_nand2 i_148(.A(n_407), .B(divq[20]), .Z(n_535));
	notech_and2 i_147(.A(n_406), .B(divq[19]), .Z(n_845));
	notech_nand2 i_146(.A(n_405), .B(divq[18]), .Z(n_533));
	notech_and2 i_145(.A(n_404), .B(divq[17]), .Z(n_844));
	notech_nand2 i_144(.A(n_403), .B(divq[16]), .Z(n_531));
	notech_and2 i_143(.A(n_402), .B(divq[15]), .Z(n_843));
	notech_nand2 i_142(.A(n_401), .B(divq[14]), .Z(n_529));
	notech_and2 i_141(.A(n_400), .B(divq[13]), .Z(n_842));
	notech_nand2 i_140(.A(n_399), .B(divq[12]), .Z(n_527));
	notech_and2 i_139(.A(n_398), .B(divq[11]), .Z(n_841));
	notech_nand2 i_138(.A(n_397), .B(divq[10]), .Z(n_525));
	notech_and2 i_137(.A(n_396), .B(divq[9]), .Z(n_840));
	notech_nand2 i_136(.A(n_395), .B(divq[8]), .Z(n_523));
	notech_and2 i_135(.A(n_394), .B(divq[7]), .Z(n_839));
	notech_nand2 i_134(.A(n_393), .B(divq[6]), .Z(n_521));
	notech_and2 i_133(.A(n_392), .B(divq[5]), .Z(n_838));
	notech_nand2 i_132(.A(n_391), .B(divq[4]), .Z(n_519));
	notech_and2 i_131(.A(n_390), .B(divq[3]), .Z(n_837));
	notech_nand2 i_130(.A(n_389), .B(divq[2]), .Z(n_517));
	notech_and2 i_129(.A(n_388), .B(divq[1]), .Z(n_836));
	notech_nand2 i_128(.A(n_387), .B(divq[0]), .Z(n_515));
	notech_nor2 i_125(.A(n_449), .B(divq[62]), .Z(n_512));
	notech_nor2 i_124(.A(n_448), .B(divq[61]), .Z(n_511));
	notech_nor2 i_123(.A(n_447), .B(divq[60]), .Z(n_510));
	notech_nor2 i_122(.A(n_446), .B(divq[59]), .Z(n_509));
	notech_nor2 i_121(.A(n_445), .B(divq[58]), .Z(n_508));
	notech_nor2 i_120(.A(n_444), .B(divq[57]), .Z(n_507));
	notech_nor2 i_119(.A(n_443), .B(divq[56]), .Z(n_506));
	notech_nor2 i_118(.A(n_442), .B(divq[55]), .Z(n_505));
	notech_nor2 i_117(.A(n_441), .B(divq[54]), .Z(n_504));
	notech_nor2 i_116(.A(n_440), .B(divq[53]), .Z(n_503));
	notech_nor2 i_115(.A(n_439), .B(divq[52]), .Z(n_502));
	notech_nor2 i_114(.A(n_438), .B(divq[51]), .Z(n_501));
	notech_nor2 i_113(.A(n_437), .B(divq[50]), .Z(n_500));
	notech_nor2 i_112(.A(n_436), .B(divq[49]), .Z(n_499));
	notech_nor2 i_111(.A(n_435), .B(divq[48]), .Z(n_498));
	notech_nor2 i_110(.A(n_434), .B(divq[47]), .Z(n_497));
	notech_nor2 i_109(.A(n_433), .B(divq[46]), .Z(n_496));
	notech_nor2 i_108(.A(n_432), .B(divq[45]), .Z(n_495));
	notech_nor2 i_107(.A(n_431), .B(divq[44]), .Z(n_494));
	notech_nor2 i_106(.A(n_430), .B(divq[43]), .Z(n_493));
	notech_nor2 i_105(.A(n_429), .B(divq[42]), .Z(n_492));
	notech_nor2 i_104(.A(n_428), .B(divq[41]), .Z(n_491));
	notech_nor2 i_103(.A(n_427), .B(divq[40]), .Z(n_490));
	notech_nor2 i_102(.A(n_426), .B(divq[39]), .Z(n_489));
	notech_nor2 i_101(.A(n_425), .B(divq[38]), .Z(n_488));
	notech_nor2 i_100(.A(n_424), .B(divq[37]), .Z(n_487));
	notech_nor2 i_99(.A(n_423), .B(divq[36]), .Z(n_486));
	notech_nor2 i_98(.A(n_422), .B(divq[35]), .Z(n_485));
	notech_nor2 i_97(.A(n_421), .B(divq[34]), .Z(n_484));
	notech_nor2 i_96(.A(n_420), .B(divq[33]), .Z(n_483));
	notech_nor2 i_95(.A(n_419), .B(divq[32]), .Z(n_482));
	notech_nor2 i_94(.A(n_418), .B(divq[31]), .Z(n_481));
	notech_nor2 i_93(.A(n_417), .B(divq[30]), .Z(n_480));
	notech_nor2 i_92(.A(n_416), .B(divq[29]), .Z(n_479));
	notech_nor2 i_91(.A(n_415), .B(divq[28]), .Z(n_478));
	notech_nor2 i_90(.A(n_414), .B(divq[27]), .Z(n_477));
	notech_nor2 i_89(.A(n_413), .B(divq[26]), .Z(n_476));
	notech_nor2 i_88(.A(n_412), .B(divq[25]), .Z(n_475));
	notech_nor2 i_87(.A(n_411), .B(divq[24]), .Z(n_474));
	notech_nor2 i_86(.A(n_410), .B(divq[23]), .Z(n_473));
	notech_nor2 i_85(.A(n_409), .B(divq[22]), .Z(n_472));
	notech_nor2 i_84(.A(n_408), .B(divq[21]), .Z(n_471));
	notech_nor2 i_83(.A(n_407), .B(divq[20]), .Z(n_470));
	notech_nor2 i_82(.A(n_406), .B(divq[19]), .Z(n_469));
	notech_nor2 i_81(.A(n_405), .B(divq[18]), .Z(n_468));
	notech_nor2 i_80(.A(n_404), .B(divq[17]), .Z(n_467));
	notech_nor2 i_79(.A(n_403), .B(divq[16]), .Z(n_466));
	notech_nor2 i_78(.A(n_402), .B(divq[15]), .Z(n_465));
	notech_nor2 i_77(.A(n_401), .B(divq[14]), .Z(n_464));
	notech_nor2 i_76(.A(n_400), .B(divq[13]), .Z(n_463));
	notech_nor2 i_75(.A(n_399), .B(divq[12]), .Z(n_462));
	notech_nor2 i_74(.A(n_398), .B(divq[11]), .Z(n_461));
	notech_nor2 i_73(.A(n_397), .B(divq[10]), .Z(n_460));
	notech_nor2 i_72(.A(n_396), .B(divq[9]), .Z(n_459));
	notech_nor2 i_71(.A(n_395), .B(divq[8]), .Z(n_458));
	notech_nor2 i_70(.A(n_394), .B(divq[7]), .Z(n_457));
	notech_nor2 i_69(.A(n_393), .B(divq[6]), .Z(n_456));
	notech_nor2 i_68(.A(n_392), .B(divq[5]), .Z(n_455));
	notech_nor2 i_67(.A(n_391), .B(divq[4]), .Z(n_454));
	notech_nor2 i_66(.A(n_390), .B(divq[3]), .Z(n_453));
	notech_nor2 i_65(.A(n_389), .B(divq[2]), .Z(n_452));
	notech_nor2 i_64(.A(n_388), .B(divq[1]), .Z(n_451));
	notech_inv i_62(.A(I0[62]), .Z(n_449));
	notech_inv i_61(.A(I0[61]), .Z(n_448));
	notech_inv i_60(.A(I0[60]), .Z(n_447));
	notech_inv i_59(.A(I0[59]), .Z(n_446));
	notech_inv i_58(.A(I0[58]), .Z(n_445));
	notech_inv i_57(.A(I0[57]), .Z(n_444));
	notech_inv i_56(.A(I0[56]), .Z(n_443));
	notech_inv i_55(.A(I0[55]), .Z(n_442));
	notech_inv i_54(.A(I0[54]), .Z(n_441));
	notech_inv i_53(.A(I0[53]), .Z(n_440));
	notech_inv i_52(.A(I0[52]), .Z(n_439));
	notech_inv i_51(.A(I0[51]), .Z(n_438));
	notech_inv i_50(.A(I0[50]), .Z(n_437));
	notech_inv i_49(.A(I0[49]), .Z(n_436));
	notech_inv i_48(.A(I0[48]), .Z(n_435));
	notech_inv i_47(.A(I0[47]), .Z(n_434));
	notech_inv i_46(.A(I0[46]), .Z(n_433));
	notech_inv i_45(.A(I0[45]), .Z(n_432));
	notech_inv i_44(.A(I0[44]), .Z(n_431));
	notech_inv i_43(.A(I0[43]), .Z(n_430));
	notech_inv i_42(.A(I0[42]), .Z(n_429));
	notech_inv i_41(.A(I0[41]), .Z(n_428));
	notech_inv i_40(.A(I0[40]), .Z(n_427));
	notech_inv i_39(.A(I0[39]), .Z(n_426));
	notech_inv i_38(.A(I0[38]), .Z(n_425));
	notech_inv i_37(.A(I0[37]), .Z(n_424));
	notech_inv i_36(.A(I0[36]), .Z(n_423));
	notech_inv i_35(.A(I0[35]), .Z(n_422));
	notech_inv i_34(.A(I0[34]), .Z(n_421));
	notech_inv i_33(.A(I0[33]), .Z(n_420));
	notech_inv i_32(.A(I0[32]), .Z(n_419));
	notech_inv i_31(.A(I0[31]), .Z(n_418));
	notech_inv i_30(.A(I0[30]), .Z(n_417));
	notech_inv i_29(.A(I0[29]), .Z(n_416));
	notech_inv i_28(.A(I0[28]), .Z(n_415));
	notech_inv i_27(.A(I0[27]), .Z(n_414));
	notech_inv i_26(.A(I0[26]), .Z(n_413));
	notech_inv i_25(.A(I0[25]), .Z(n_412));
	notech_inv i_24(.A(I0[24]), .Z(n_411));
	notech_inv i_23(.A(I0[23]), .Z(n_410));
	notech_inv i_22(.A(I0[22]), .Z(n_409));
	notech_inv i_21(.A(I0[21]), .Z(n_408));
	notech_inv i_20(.A(I0[20]), .Z(n_407));
	notech_inv i_19(.A(I0[19]), .Z(n_406));
	notech_inv i_18(.A(I0[18]), .Z(n_405));
	notech_inv i_17(.A(I0[17]), .Z(n_404));
	notech_inv i_16(.A(I0[16]), .Z(n_403));
	notech_inv i_15(.A(I0[15]), .Z(n_402));
	notech_inv i_14(.A(I0[14]), .Z(n_401));
	notech_inv i_13(.A(I0[13]), .Z(n_400));
	notech_inv i_12(.A(I0[12]), .Z(n_399));
	notech_inv i_11(.A(I0[11]), .Z(n_398));
	notech_inv i_10(.A(I0[10]), .Z(n_397));
	notech_inv i_9(.A(I0[9]), .Z(n_396));
	notech_inv i_8(.A(I0[8]), .Z(n_395));
	notech_inv i_7(.A(I0[7]), .Z(n_394));
	notech_inv i_6(.A(I0[6]), .Z(n_393));
	notech_inv i_5(.A(I0[5]), .Z(n_392));
	notech_inv i_4(.A(I0[4]), .Z(n_391));
	notech_inv i_3(.A(I0[3]), .Z(n_390));
	notech_inv i_2(.A(I0[2]), .Z(n_389));
	notech_inv i_1(.A(I0[1]), .Z(n_388));
	notech_inv i_0(.A(I0[0]), .Z(n_387));
endmodule
module AWDP_LSH_38(O0, opb);
    output [31:0] O0;
    input [4:0] opb;
    // Line 636
    wire [31:0] N745;
    // Line 348
    wire [31:0] O0;

    // Line 636
    assign N745 = 5'h1 << opb;
    // Line 348
    assign O0 = N745;
endmodule

module AWDP_LSH_9(O0, opd);
    output [31:0] O0;
    input [5:0] opd;
    // Line 1006
    wire [31:0] N760;
    wire [31:0] O0;

    // Line 1006
    assign N760 = 6'h1 << opd;
    assign O0 = N760;
endmodule

module AWDP_SUB_129(O0, opa, I0);

	output [16:0] O0;
	input [15:0] opa;
	input [15:0] I0;




	notech_inv i_10544(.A(I0[13]), .Z(n_57264));
	notech_inv i_32(.A(n_230), .Z(O0[16]));
	notech_fa2 i_31(.A(n_57264), .B(n_228), .CI(opa[15]), .Z(O0[15]), .CO(n_230
		));
	notech_fa2 i_30(.A(n_57264), .B(n_226), .CI(opa[14]), .Z(O0[14]), .CO(n_228
		));
	notech_fa2 i_29(.A(n_57264), .B(n_224), .CI(opa[13]), .Z(O0[13]), .CO(n_226
		));
	notech_fa2 i_28(.A(n_57264), .B(n_222), .CI(opa[12]), .Z(O0[12]), .CO(n_224
		));
	notech_fa2 i_27(.A(n_57264), .B(n_220), .CI(opa[11]), .Z(O0[11]), .CO(n_222
		));
	notech_fa2 i_26(.A(n_57264), .B(n_218), .CI(opa[10]), .Z(O0[10]), .CO(n_220
		));
	notech_fa2 i_25(.A(n_57264), .B(n_216), .CI(opa[9]), .Z(O0[9]), .CO(n_218
		));
	notech_fa2 i_24(.A(n_57264), .B(n_214), .CI(opa[8]), .Z(O0[8]), .CO(n_216
		));
	notech_fa2 i_23(.A(n_57264), .B(n_212), .CI(opa[7]), .Z(O0[7]), .CO(n_214
		));
	notech_fa2 i_22(.A(n_57264), .B(n_210), .CI(opa[6]), .Z(O0[6]), .CO(n_212
		));
	notech_fa2 i_21(.A(n_57264), .B(n_208), .CI(opa[5]), .Z(O0[5]), .CO(n_210
		));
	notech_fa2 i_20(.A(n_57264), .B(n_206), .CI(opa[4]), .Z(O0[4]), .CO(n_208
		));
	notech_fa2 i_19(.A(n_57264), .B(n_204), .CI(opa[3]), .Z(O0[3]), .CO(n_206
		));
	notech_fa2 i_18(.A(n_57264), .B(n_202), .CI(opa[2]), .Z(O0[2]), .CO(n_204
		));
	notech_fa2 i_17(.A(n_184), .B(n_200), .CI(opa[1]), .Z(O0[1]), .CO(n_202)
		);
	notech_inv i_1(.A(I0[1]), .Z(n_184));
	notech_inv i_0(.A(I0[0]), .Z(n_183));
	notech_xor2 i_60(.A(opa[0]), .B(n_183), .Z(n_45796));
	notech_inv i_61(.A(n_45796), .Z(O0[0]));
	notech_or2 i_59(.A(opa[0]), .B(n_183), .Z(n_200));
endmodule
module AWDP_SUB_177(O0, opd);

	output [31:0] O0;
	input [31:0] opd;

	wire \opd[2] ;
	wire \opd[3] ;
	wire \opd[4] ;
	wire \opd[5] ;
	wire \opd[6] ;
	wire \opd[7] ;
	wire \opd[8] ;
	wire \opd[9] ;
	wire \opd[10] ;
	wire \opd[11] ;
	wire \opd[12] ;
	wire \opd[13] ;
	wire \opd[14] ;
	wire \opd[15] ;
	wire \opd[16] ;
	wire \opd[17] ;
	wire \opd[18] ;
	wire \opd[19] ;
	wire \opd[20] ;
	wire \opd[21] ;
	wire \opd[22] ;
	wire \opd[23] ;
	wire \opd[24] ;
	wire \opd[25] ;
	wire \opd[26] ;
	wire \opd[27] ;
	wire \opd[28] ;
	wire \opd[29] ;
	wire \opd[30] ;
	wire \opd[31] ;


	assign O0[0] = opd[0];
	assign O0[1] = opd[1];
	assign \opd[2]  = opd[2];
	assign \opd[3]  = opd[3];
	assign \opd[4]  = opd[4];
	assign \opd[5]  = opd[5];
	assign \opd[6]  = opd[6];
	assign \opd[7]  = opd[7];
	assign \opd[8]  = opd[8];
	assign \opd[9]  = opd[9];
	assign \opd[10]  = opd[10];
	assign \opd[11]  = opd[11];
	assign \opd[12]  = opd[12];
	assign \opd[13]  = opd[13];
	assign \opd[14]  = opd[14];
	assign \opd[15]  = opd[15];
	assign \opd[16]  = opd[16];
	assign \opd[17]  = opd[17];
	assign \opd[18]  = opd[18];
	assign \opd[19]  = opd[19];
	assign \opd[20]  = opd[20];
	assign \opd[21]  = opd[21];
	assign \opd[22]  = opd[22];
	assign \opd[23]  = opd[23];
	assign \opd[24]  = opd[24];
	assign \opd[25]  = opd[25];
	assign \opd[26]  = opd[26];
	assign \opd[27]  = opd[27];
	assign \opd[28]  = opd[28];
	assign \opd[29]  = opd[29];
	assign \opd[30]  = opd[30];
	assign \opd[31]  = opd[31];

	notech_ha2 i_30(.A(n_192), .B(n_250), .Z(O0[31]));
	notech_inv i_1(.A(\opd[2] ), .Z(O0[2]));
	notech_inv i_0(.A(\opd[31] ), .Z(n_192));
	notech_xor2 i_47(.A(\opd[30] ), .B(n_248), .Z(n_45823));
	notech_inv i_48(.A(n_45823), .Z(O0[30]));
	notech_or2 i_46(.A(\opd[30] ), .B(n_248), .Z(n_250));
	notech_xor2 i_4695829(.A(\opd[29] ), .B(n_246), .Z(n_45850));
	notech_inv i_4795830(.A(n_45850), .Z(O0[29]));
	notech_or2 i_45(.A(\opd[29] ), .B(n_246), .Z(n_248));
	notech_xor2 i_44(.A(\opd[28] ), .B(n_244), .Z(n_45877));
	notech_inv i_4595831(.A(n_45877), .Z(O0[28]));
	notech_or2 i_43(.A(\opd[28] ), .B(n_244), .Z(n_246));
	notech_xor2 i_4395832(.A(\opd[27] ), .B(n_242), .Z(n_45904));
	notech_inv i_4495833(.A(n_45904), .Z(O0[27]));
	notech_or2 i_42(.A(\opd[27] ), .B(n_242), .Z(n_244));
	notech_xor2 i_4295834(.A(\opd[26] ), .B(n_240), .Z(n_45931));
	notech_inv i_4395835(.A(n_45931), .Z(O0[26]));
	notech_or2 i_41(.A(\opd[26] ), .B(n_240), .Z(n_242));
	notech_xor2 i_4195836(.A(\opd[25] ), .B(n_238), .Z(n_45958));
	notech_inv i_4295837(.A(n_45958), .Z(O0[25]));
	notech_or2 i_40(.A(\opd[25] ), .B(n_238), .Z(n_240));
	notech_xor2 i_4095838(.A(\opd[24] ), .B(n_236), .Z(n_45985));
	notech_inv i_4195839(.A(n_45985), .Z(O0[24]));
	notech_or2 i_39(.A(\opd[24] ), .B(n_236), .Z(n_238));
	notech_xor2 i_3995840(.A(\opd[23] ), .B(n_234), .Z(n_46012));
	notech_inv i_4095841(.A(n_46012), .Z(O0[23]));
	notech_or2 i_38(.A(\opd[23] ), .B(n_234), .Z(n_236));
	notech_xor2 i_3895842(.A(\opd[22] ), .B(n_232), .Z(n_46039));
	notech_inv i_3995843(.A(n_46039), .Z(O0[22]));
	notech_or2 i_37(.A(\opd[22] ), .B(n_232), .Z(n_234));
	notech_xor2 i_3795844(.A(\opd[21] ), .B(n_230), .Z(n_46066));
	notech_inv i_3895845(.A(n_46066), .Z(O0[21]));
	notech_or2 i_36(.A(\opd[21] ), .B(n_230), .Z(n_232));
	notech_xor2 i_3695846(.A(\opd[20] ), .B(n_228), .Z(n_46093));
	notech_inv i_3795847(.A(n_46093), .Z(O0[20]));
	notech_or2 i_35(.A(\opd[20] ), .B(n_228), .Z(n_230));
	notech_xor2 i_3595848(.A(\opd[19] ), .B(n_226), .Z(n_46120));
	notech_inv i_3695849(.A(n_46120), .Z(O0[19]));
	notech_or2 i_34(.A(\opd[19] ), .B(n_226), .Z(n_228));
	notech_xor2 i_3495850(.A(\opd[18] ), .B(n_224), .Z(n_46147));
	notech_inv i_3595851(.A(n_46147), .Z(O0[18]));
	notech_or2 i_33(.A(\opd[18] ), .B(n_224), .Z(n_226));
	notech_xor2 i_3395852(.A(\opd[17] ), .B(n_222), .Z(n_46174));
	notech_inv i_3495853(.A(n_46174), .Z(O0[17]));
	notech_or2 i_32(.A(\opd[17] ), .B(n_222), .Z(n_224));
	notech_xor2 i_3295854(.A(\opd[16] ), .B(n_220), .Z(n_46201));
	notech_inv i_3395855(.A(n_46201), .Z(O0[16]));
	notech_or2 i_31(.A(\opd[16] ), .B(n_220), .Z(n_222));
	notech_xor2 i_3195856(.A(\opd[15] ), .B(n_218), .Z(n_46228));
	notech_inv i_3295857(.A(n_46228), .Z(O0[15]));
	notech_or2 i_3095858(.A(\opd[15] ), .B(n_218), .Z(n_220));
	notech_xor2 i_3095859(.A(\opd[14] ), .B(n_216), .Z(n_46255));
	notech_inv i_3195860(.A(n_46255), .Z(O0[14]));
	notech_or2 i_29(.A(\opd[14] ), .B(n_216), .Z(n_218));
	notech_xor2 i_2995861(.A(\opd[13] ), .B(n_214), .Z(n_46282));
	notech_inv i_3095862(.A(n_46282), .Z(O0[13]));
	notech_or2 i_28(.A(\opd[13] ), .B(n_214), .Z(n_216));
	notech_xor2 i_2895863(.A(\opd[12] ), .B(n_212), .Z(n_46309));
	notech_inv i_2995864(.A(n_46309), .Z(O0[12]));
	notech_or2 i_27(.A(\opd[12] ), .B(n_212), .Z(n_214));
	notech_xor2 i_2795865(.A(\opd[11] ), .B(n_210), .Z(n_46336));
	notech_inv i_2895866(.A(n_46336), .Z(O0[11]));
	notech_or2 i_26(.A(\opd[11] ), .B(n_210), .Z(n_212));
	notech_xor2 i_2795867(.A(\opd[10] ), .B(n_208), .Z(n_46363));
	notech_inv i_2895868(.A(n_46363), .Z(O0[10]));
	notech_or2 i_2695869(.A(\opd[10] ), .B(n_208), .Z(n_210));
	notech_xor2 i_2795870(.A(\opd[9] ), .B(n_206), .Z(n_46390));
	notech_inv i_2895871(.A(n_46390), .Z(O0[9]));
	notech_or2 i_2695872(.A(\opd[9] ), .B(n_206), .Z(n_208));
	notech_xor2 i_2795873(.A(\opd[8] ), .B(n_204), .Z(n_46417));
	notech_inv i_2895874(.A(n_46417), .Z(O0[8]));
	notech_or2 i_2695875(.A(\opd[8] ), .B(n_204), .Z(n_206));
	notech_xor2 i_2795876(.A(\opd[7] ), .B(n_202), .Z(n_46444));
	notech_inv i_2895877(.A(n_46444), .Z(O0[7]));
	notech_or2 i_2695878(.A(\opd[7] ), .B(n_202), .Z(n_204));
	notech_xor2 i_2795879(.A(\opd[6] ), .B(n_200), .Z(n_46471));
	notech_inv i_2895880(.A(n_46471), .Z(O0[6]));
	notech_or2 i_2695881(.A(\opd[6] ), .B(n_200), .Z(n_202));
	notech_xor2 i_2795882(.A(\opd[5] ), .B(n_198), .Z(n_46498));
	notech_inv i_2895883(.A(n_46498), .Z(O0[5]));
	notech_or2 i_2695884(.A(\opd[5] ), .B(n_198), .Z(n_200));
	notech_xor2 i_2795885(.A(\opd[4] ), .B(n_196), .Z(n_46525));
	notech_inv i_2895886(.A(n_46525), .Z(O0[4]));
	notech_or2 i_2695887(.A(\opd[4] ), .B(n_196), .Z(n_198));
	notech_xor2 i_2795888(.A(\opd[3] ), .B(\opd[2] ), .Z(n_46553));
	notech_inv i_2895889(.A(n_46553), .Z(O0[3]));
	notech_or2 i_2695890(.A(\opd[3] ), .B(\opd[2] ), .Z(n_196));
endmodule
module AWDP_SUB_197(O0, regs_7, opd);
    output [31:0] O0;
    input [31:0] regs_7;
    input [31:0] opd;
    // Line 521
    wire [31:0] N800;
    // Line 348
    wire [31:0] O0;

    // Line 521
    assign N800 = regs_7 - opd;
    // Line 348
    assign O0 = N800;
endmodule

module AWDP_SUB_200(O0, regs_6, opd);
    output [31:0] O0;
    input [31:0] regs_6;
    input [31:0] opd;
    // Line 521
    wire [31:0] N815;
    // Line 348
    wire [31:0] O0;

    // Line 521
    assign N815 = regs_6 - opd;
    // Line 348
    assign O0 = N815;
endmodule

module AWDP_SUB_206(O0, opa, I0);

	output [32:0] O0;
	input [31:0] opa;
	input [31:0] I0;




	notech_inv i_10529(.A(n_57188), .Z(n_57189));
	notech_inv i_10528(.A(I0[19]), .Z(n_57188));
	notech_inv i_64(.A(n_454), .Z(O0[32]));
	notech_fa2 i_63(.A(n_57188), .B(n_452), .CI(opa[31]), .Z(O0[31]), .CO(n_454
		));
	notech_fa2 i_62(.A(n_57188), .B(n_450), .CI(opa[30]), .Z(O0[30]), .CO(n_452
		));
	notech_fa2 i_61(.A(n_57188), .B(n_448), .CI(opa[29]), .Z(O0[29]), .CO(n_450
		));
	notech_fa2 i_60(.A(n_57188), .B(n_446), .CI(opa[28]), .Z(O0[28]), .CO(n_448
		));
	notech_fa2 i_59(.A(n_57188), .B(n_444), .CI(opa[27]), .Z(O0[27]), .CO(n_446
		));
	notech_fa2 i_58(.A(n_57188), .B(n_442), .CI(opa[26]), .Z(O0[26]), .CO(n_444
		));
	notech_fa2 i_57(.A(n_57188), .B(n_440), .CI(opa[25]), .Z(O0[25]), .CO(n_442
		));
	notech_fa2 i_56(.A(n_57188), .B(n_438), .CI(opa[24]), .Z(O0[24]), .CO(n_440
		));
	notech_fa2 i_55(.A(n_57188), .B(n_436), .CI(opa[23]), .Z(O0[23]), .CO(n_438
		));
	notech_fa2 i_54(.A(n_57188), .B(n_434), .CI(opa[22]), .Z(O0[22]), .CO(n_436
		));
	notech_fa2 i_53(.A(n_57188), .B(n_432), .CI(opa[21]), .Z(O0[21]), .CO(n_434
		));
	notech_fa2 i_52(.A(n_57188), .B(n_430), .CI(opa[20]), .Z(O0[20]), .CO(n_432
		));
	notech_fa2 i_51(.A(n_57188), .B(n_428), .CI(opa[19]), .Z(O0[19]), .CO(n_430
		));
	notech_fa2 i_50(.A(n_57188), .B(n_426), .CI(opa[18]), .Z(O0[18]), .CO(n_428
		));
	notech_fa2 i_49(.A(n_57188), .B(n_424), .CI(opa[17]), .Z(O0[17]), .CO(n_426
		));
	notech_fa2 i_48(.A(n_361), .B(n_422), .CI(opa[16]), .Z(O0[16]), .CO(n_424
		));
	notech_fa2 i_47(.A(n_361), .B(n_420), .CI(opa[15]), .Z(O0[15]), .CO(n_422
		));
	notech_fa2 i_46(.A(n_361), .B(n_418), .CI(opa[14]), .Z(O0[14]), .CO(n_420
		));
	notech_fa2 i_45(.A(n_361), .B(n_416), .CI(opa[13]), .Z(O0[13]), .CO(n_418
		));
	notech_fa2 i_44(.A(n_361), .B(n_414), .CI(opa[12]), .Z(O0[12]), .CO(n_416
		));
	notech_fa2 i_43(.A(n_361), .B(n_412), .CI(opa[11]), .Z(O0[11]), .CO(n_414
		));
	notech_fa2 i_42(.A(n_361), .B(n_410), .CI(opa[10]), .Z(O0[10]), .CO(n_412
		));
	notech_fa2 i_41(.A(n_361), .B(n_408), .CI(opa[9]), .Z(O0[9]), .CO(n_410)
		);
	notech_fa2 i_40(.A(n_361), .B(n_406), .CI(opa[8]), .Z(O0[8]), .CO(n_408)
		);
	notech_fa2 i_39(.A(n_361), .B(n_404), .CI(opa[7]), .Z(O0[7]), .CO(n_406)
		);
	notech_fa2 i_38(.A(n_361), .B(n_402), .CI(opa[6]), .Z(O0[6]), .CO(n_404)
		);
	notech_fa2 i_37(.A(n_361), .B(n_400), .CI(opa[5]), .Z(O0[5]), .CO(n_402)
		);
	notech_fa2 i_36(.A(n_361), .B(n_398), .CI(opa[4]), .Z(O0[4]), .CO(n_400)
		);
	notech_fa2 i_35(.A(n_361), .B(n_396), .CI(opa[3]), .Z(O0[3]), .CO(n_398)
		);
	notech_fa2 i_34(.A(n_361), .B(n_394), .CI(opa[2]), .Z(O0[2]), .CO(n_396)
		);
	notech_fa2 i_33(.A(n_360), .B(n_392), .CI(opa[1]), .Z(O0[1]), .CO(n_394)
		);
	notech_inv i_2(.A(n_57189), .Z(n_361));
	notech_inv i_1(.A(I0[1]), .Z(n_360));
	notech_inv i_0(.A(I0[0]), .Z(n_359));
	notech_xor2 i_81(.A(opa[0]), .B(n_359), .Z(n_46634));
	notech_inv i_82(.A(n_46634), .Z(O0[0]));
	notech_or2 i_80(.A(opa[0]), .B(n_359), .Z(n_392));
endmodule
module AWDP_SUB_237(O0, divr, divq);
    output [63:0] O0;
    input [63:0] divr;
    input [63:0] divq;
    // Line 1006
    wire [63:0] N835;
    // Line 1006
    wire [63:0] O0;

    // Line 1006
    assign N835 = divr - divq;
    // Line 1006
    assign O0 = N835;
endmodule

module AWDP_SUB_81(O0, regs_4, calc_sz);
    output [31:0] O0;
    input [31:0] regs_4;
    input [2:0] calc_sz;
    // Line 348
    wire [31:0] O0;
    // Line 456
    wire [31:0] N848;

    // Line 348
    assign O0 = N848;
    // Line 456
    assign N848 = regs_4 - calc_sz;
endmodule

module AWMUX_16_1(I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14
		, I15, S, O0);

	input I0;
	input I1;
	input I2;
	input I3;
	input I4;
	input I5;
	input I6;
	input I7;
	input I8;
	input I9;
	input I10;
	input I11;
	input I12;
	input I13;
	input I14;
	input I15;
	input [3:0] S;
	output O0;




	notech_inv i_16118(.A(n_62871), .Z(n_62872));
	notech_inv i_16117(.A(S[0]), .Z(n_62871));
	notech_mux4 i_14(.S0(S[2]), .S1(S[3]), .A(n_23), .B(n_26), .C(n_29), .D(n_32
		), .Z(O0));
	notech_mux4 i_11(.S0(n_62872), .S1(S[1]), .A(I12), .B(n_14531), .C(I14),
		 .D(n_14530), .Z(n_32));
	notech_mux4 i_8(.S0(n_62872), .S1(S[1]), .A(I8), .B(n_14533), .C(I10), .D
		(n_14532), .Z(n_29));
	notech_mux4 i_5(.S0(n_62872), .S1(S[1]), .A(I4), .B(n_14535), .C(I6), .D
		(n_14534), .Z(n_26));
	notech_mux4 i_2(.S0(n_62872), .S1(S[1]), .A(I0), .B(n_14537), .C(I2), .D
		(n_14536), .Z(n_23));
	notech_inv i_41(.A(I14), .Z(n_14530));
	notech_inv i_42(.A(I12), .Z(n_14531));
	notech_inv i_43(.A(I10), .Z(n_14532));
	notech_inv i_44(.A(I8), .Z(n_14533));
	notech_inv i_45(.A(I6), .Z(n_14534));
	notech_inv i_46(.A(I4), .Z(n_14535));
	notech_inv i_47(.A(I2), .Z(n_14536));
	notech_inv i_48(.A(I0), .Z(n_14537));
endmodule
module AWMUX_16_32_0(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_1(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_2(I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13,
		 I14, I15, S, O0);

	input [31:0] I0;
	input [31:0] I1;
	input [31:0] I2;
	input [31:0] I3;
	input [31:0] I4;
	input [31:0] I5;
	input [31:0] I6;
	input [31:0] I7;
	input [31:0] I8;
	input [31:0] I9;
	input [31:0] I10;
	input [31:0] I11;
	input [31:0] I12;
	input [31:0] I13;
	input [31:0] I14;
	input [31:0] I15;
	input [3:0] S;
	output [31:0] O0;




	notech_inv i_7707(.A(n_53849), .Z(n_54140));
	notech_inv i_7702(.A(n_53849), .Z(n_54135));
	notech_inv i_7697(.A(n_53838), .Z(n_54129));
	notech_inv i_7692(.A(n_53838), .Z(n_54124));
	notech_inv i_7447(.A(n_53871), .Z(n_53872));
	notech_inv i_7446(.A(n_14529), .Z(n_53871));
	notech_inv i_7444(.A(n_723), .Z(n_53868));
	notech_inv i_7442(.A(n_723), .Z(n_53866));
	notech_inv i_7439(.A(n_723), .Z(n_53863));
	notech_inv i_7437(.A(n_723), .Z(n_53861));
	notech_inv i_7427(.A(n_53849), .Z(n_53850));
	notech_inv i_7426(.A(n_548), .Z(n_53849));
	notech_inv i_7417(.A(n_53838), .Z(n_53839));
	notech_inv i_7416(.A(n_549), .Z(n_53838));
	notech_inv i_180(.A(S[3]), .Z(n_723));
	notech_inv i_179(.A(n_722), .Z(n_684));
	notech_inv i_178(.A(S[2]), .Z(n_722));
	notech_mux4 i_67(.S0(n_548), .S1(n_549), .A(I4[31]), .B(I5[31]), .C(I6[
		31]), .D(I7[31]), .Z(n_615));
	notech_mux4 i_66(.S0(n_548), .S1(n_549), .A(I4[30]), .B(I5[30]), .C(I6[
		30]), .D(I7[30]), .Z(n_614));
	notech_mux4 i_65(.S0(n_548), .S1(n_549), .A(I4[29]), .B(I5[29]), .C(I6[
		29]), .D(I7[29]), .Z(n_613));
	notech_mux4 i_64(.S0(n_548), .S1(n_549), .A(I4[28]), .B(I5[28]), .C(I6[
		28]), .D(I7[28]), .Z(n_612));
	notech_mux4 i_63(.S0(n_548), .S1(n_549), .A(I4[27]), .B(I5[27]), .C(I6[
		27]), .D(I7[27]), .Z(n_611));
	notech_mux4 i_62(.S0(n_548), .S1(n_549), .A(I4[26]), .B(I5[26]), .C(I6[
		26]), .D(I7[26]), .Z(n_610));
	notech_mux4 i_61(.S0(n_548), .S1(n_549), .A(I4[25]), .B(I5[25]), .C(I6[
		25]), .D(I7[25]), .Z(n_609));
	notech_mux4 i_60(.S0(n_548), .S1(n_549), .A(I4[24]), .B(I5[24]), .C(I6[
		24]), .D(I7[24]), .Z(n_608));
	notech_mux4 i_59(.S0(n_548), .S1(n_549), .A(I4[23]), .B(I5[23]), .C(I6[
		23]), .D(I7[23]), .Z(n_607));
	notech_mux4 i_58(.S0(n_548), .S1(n_549), .A(I4[22]), .B(I5[22]), .C(I6[
		22]), .D(I7[22]), .Z(n_606));
	notech_mux4 i_57(.S0(n_548), .S1(n_549), .A(I4[21]), .B(I5[21]), .C(I6[
		21]), .D(I7[21]), .Z(n_605));
	notech_mux4 i_56(.S0(n_548), .S1(n_549), .A(I4[20]), .B(I5[20]), .C(I6[
		20]), .D(I7[20]), .Z(n_604));
	notech_mux4 i_55(.S0(n_548), .S1(n_549), .A(I4[19]), .B(I5[19]), .C(I6[
		19]), .D(I7[19]), .Z(n_603));
	notech_mux4 i_54(.S0(n_548), .S1(n_549), .A(I4[18]), .B(I5[18]), .C(I6[
		18]), .D(I7[18]), .Z(n_602));
	notech_mux4 i_53(.S0(n_548), .S1(n_549), .A(I4[17]), .B(I5[17]), .C(I6[
		17]), .D(I7[17]), .Z(n_601));
	notech_mux4 i_52(.S0(n_548), .S1(n_549), .A(I4[16]), .B(I5[16]), .C(I6[
		16]), .D(I7[16]), .Z(n_600));
	notech_mux4 i_51(.S0(n_53850), .S1(n_53839), .A(I4[15]), .B(I5[15]), .C(I6
		[15]), .D(I7[15]), .Z(n_599));
	notech_mux4 i_50(.S0(n_53850), .S1(n_53839), .A(I4[14]), .B(I5[14]), .C(I6
		[14]), .D(I7[14]), .Z(n_598));
	notech_mux4 i_49(.S0(n_53850), .S1(n_53839), .A(I4[13]), .B(I5[13]), .C(I6
		[13]), .D(I7[13]), .Z(n_597));
	notech_mux4 i_48(.S0(n_53850), .S1(n_53839), .A(I4[12]), .B(I5[12]), .C(I6
		[12]), .D(I7[12]), .Z(n_596));
	notech_mux4 i_47(.S0(n_53850), .S1(n_53839), .A(I4[11]), .B(I5[11]), .C(I6
		[11]), .D(I7[11]), .Z(n_595));
	notech_mux4 i_46(.S0(n_53850), .S1(n_53839), .A(I4[10]), .B(I5[10]), .C(I6
		[10]), .D(I7[10]), .Z(n_594));
	notech_mux4 i_45(.S0(n_53850), .S1(n_53839), .A(I4[9]), .B(I5[9]), .C(I6
		[9]), .D(I7[9]), .Z(n_593));
	notech_mux4 i_44(.S0(n_53850), .S1(n_53839), .A(I4[8]), .B(I5[8]), .C(I6
		[8]), .D(I7[8]), .Z(n_592));
	notech_mux4 i_43(.S0(n_53850), .S1(n_53839), .A(I4[7]), .B(I5[7]), .C(I6
		[7]), .D(I7[7]), .Z(n_591));
	notech_mux4 i_42(.S0(n_53850), .S1(n_53839), .A(I4[6]), .B(I5[6]), .C(I6
		[6]), .D(I7[6]), .Z(n_590));
	notech_mux4 i_41(.S0(n_53850), .S1(n_53839), .A(I4[5]), .B(I5[5]), .C(I6
		[5]), .D(I7[5]), .Z(n_589));
	notech_mux4 i_40(.S0(n_53850), .S1(n_53839), .A(I4[4]), .B(I5[4]), .C(I6
		[4]), .D(I7[4]), .Z(n_588));
	notech_mux4 i_39(.S0(n_53850), .S1(n_53839), .A(I4[3]), .B(I5[3]), .C(I6
		[3]), .D(I7[3]), .Z(n_587));
	notech_mux4 i_38(.S0(n_53850), .S1(n_53839), .A(I4[2]), .B(I5[2]), .C(I6
		[2]), .D(I7[2]), .Z(n_586));
	notech_mux4 i_37(.S0(n_53850), .S1(n_53839), .A(I4[1]), .B(I5[1]), .C(I6
		[1]), .D(I7[1]), .Z(n_585));
	notech_mux4 i_36(.S0(n_53850), .S1(n_53839), .A(I4[0]), .B(I5[0]), .C(I6
		[0]), .D(I7[0]), .Z(n_584));
	notech_mux4 i_33(.S0(n_54135), .S1(n_54124), .A(I0[31]), .B(I1[31]), .C(I2
		[31]), .D(I3[31]), .Z(n_581));
	notech_mux4 i_32(.S0(n_54135), .S1(n_54124), .A(I0[30]), .B(I1[30]), .C(I2
		[30]), .D(I3[30]), .Z(n_580));
	notech_mux4 i_31(.S0(n_54135), .S1(n_54124), .A(I0[29]), .B(I1[29]), .C(I2
		[29]), .D(I3[29]), .Z(n_579));
	notech_mux4 i_30(.S0(n_54135), .S1(n_54124), .A(I0[28]), .B(I1[28]), .C(I2
		[28]), .D(I3[28]), .Z(n_578));
	notech_mux4 i_29(.S0(n_54135), .S1(n_54124), .A(I0[27]), .B(I1[27]), .C(I2
		[27]), .D(I3[27]), .Z(n_577));
	notech_mux4 i_28(.S0(n_54135), .S1(n_54124), .A(I0[26]), .B(I1[26]), .C(I2
		[26]), .D(I3[26]), .Z(n_576));
	notech_mux4 i_27(.S0(n_54135), .S1(n_54124), .A(I0[25]), .B(I1[25]), .C(I2
		[25]), .D(I3[25]), .Z(n_575));
	notech_mux4 i_26(.S0(n_54135), .S1(n_54124), .A(I0[24]), .B(I1[24]), .C(I2
		[24]), .D(I3[24]), .Z(n_574));
	notech_mux4 i_25(.S0(n_54135), .S1(n_54124), .A(I0[23]), .B(I1[23]), .C(I2
		[23]), .D(I3[23]), .Z(n_573));
	notech_mux4 i_24(.S0(n_54135), .S1(n_54124), .A(I0[22]), .B(I1[22]), .C(I2
		[22]), .D(I3[22]), .Z(n_572));
	notech_mux4 i_23(.S0(n_54135), .S1(n_54124), .A(I0[21]), .B(I1[21]), .C(I2
		[21]), .D(I3[21]), .Z(n_571));
	notech_mux4 i_22(.S0(n_54135), .S1(n_54124), .A(I0[20]), .B(I1[20]), .C(I2
		[20]), .D(I3[20]), .Z(n_570));
	notech_mux4 i_21(.S0(n_54135), .S1(n_54124), .A(I0[19]), .B(I1[19]), .C(I2
		[19]), .D(I3[19]), .Z(n_569));
	notech_mux4 i_20(.S0(n_54135), .S1(n_54124), .A(I0[18]), .B(I1[18]), .C(I2
		[18]), .D(I3[18]), .Z(n_568));
	notech_mux4 i_19(.S0(n_54135), .S1(n_54124), .A(I0[17]), .B(I1[17]), .C(I2
		[17]), .D(I3[17]), .Z(n_567));
	notech_mux4 i_18(.S0(n_54135), .S1(n_54124), .A(I0[16]), .B(I1[16]), .C(I2
		[16]), .D(I3[16]), .Z(n_566));
	notech_mux4 i_17(.S0(n_54140), .S1(n_54129), .A(I0[15]), .B(I1[15]), .C(I2
		[15]), .D(I3[15]), .Z(n_565));
	notech_mux4 i_16(.S0(n_54140), .S1(n_54129), .A(I0[14]), .B(I1[14]), .C(I2
		[14]), .D(I3[14]), .Z(n_564));
	notech_mux4 i_15(.S0(n_54140), .S1(n_54129), .A(I0[13]), .B(I1[13]), .C(I2
		[13]), .D(I3[13]), .Z(n_563));
	notech_mux4 i_14(.S0(n_54140), .S1(n_54129), .A(I0[12]), .B(I1[12]), .C(I2
		[12]), .D(I3[12]), .Z(n_562));
	notech_mux4 i_13(.S0(n_54140), .S1(n_54129), .A(I0[11]), .B(I1[11]), .C(I2
		[11]), .D(I3[11]), .Z(n_561));
	notech_mux4 i_12(.S0(n_54140), .S1(n_54129), .A(I0[10]), .B(I1[10]), .C(I2
		[10]), .D(I3[10]), .Z(n_560));
	notech_mux4 i_11(.S0(n_54140), .S1(n_54129), .A(I0[9]), .B(I1[9]), .C(I2
		[9]), .D(I3[9]), .Z(n_559));
	notech_mux4 i_10(.S0(n_54140), .S1(n_54129), .A(I0[8]), .B(I1[8]), .C(I2
		[8]), .D(I3[8]), .Z(n_558));
	notech_mux4 i_9(.S0(n_54140), .S1(n_54129), .A(I0[7]), .B(I1[7]), .C(I2[
		7]), .D(I3[7]), .Z(n_557));
	notech_mux4 i_8(.S0(n_54140), .S1(n_54129), .A(I0[6]), .B(I1[6]), .C(I2[
		6]), .D(I3[6]), .Z(n_556));
	notech_mux4 i_7(.S0(n_54140), .S1(n_54129), .A(I0[5]), .B(I1[5]), .C(I2[
		5]), .D(I3[5]), .Z(n_555));
	notech_mux4 i_6(.S0(n_54140), .S1(n_54129), .A(I0[4]), .B(I1[4]), .C(I2[
		4]), .D(I3[4]), .Z(n_554));
	notech_mux4 i_5(.S0(n_54140), .S1(n_54129), .A(I0[3]), .B(I1[3]), .C(I2[
		3]), .D(I3[3]), .Z(n_553));
	notech_mux4 i_4(.S0(n_54140), .S1(n_54129), .A(I0[2]), .B(I1[2]), .C(I2[
		2]), .D(I3[2]), .Z(n_552));
	notech_mux4 i_3(.S0(n_54140), .S1(n_54129), .A(I0[1]), .B(I1[1]), .C(I2[
		1]), .D(I3[1]), .Z(n_551));
	notech_mux4 i_2(.S0(n_54140), .S1(n_54129), .A(I0[0]), .B(I1[0]), .C(I2[
		0]), .D(I3[0]), .Z(n_550));
	notech_inv i_173(.A(n_719), .Z(n_549));
	notech_inv i_172(.A(S[1]), .Z(n_719));
	notech_inv i_171(.A(n_718), .Z(n_548));
	notech_inv i_170(.A(S[0]), .Z(n_718));
	notech_nand2 i_21807(.A(n_13767), .B(n_13770), .Z(O0[0]));
	notech_nao3 i_21799(.A(n_53871), .B(n_584), .C(n_53863), .Z(n_13770));
	notech_nao3 i_21796(.A(n_550), .B(n_14529), .C(n_53863), .Z(n_13767));
	notech_nand2 i_5095227(.A(n_13791), .B(n_13794), .Z(O0[1]));
	notech_nao3 i_4295228(.A(n_53871), .B(n_585), .C(n_53863), .Z(n_13794)
		);
	notech_nao3 i_3995229(.A(n_551), .B(n_53872), .C(n_53863), .Z(n_13791)
		);
	notech_nand2 i_5095231(.A(n_13815), .B(n_13818), .Z(O0[2]));
	notech_nao3 i_4295232(.A(n_53871), .B(n_586), .C(n_53863), .Z(n_13818)
		);
	notech_nao3 i_3995233(.A(n_552), .B(n_14529), .C(n_53863), .Z(n_13815)
		);
	notech_nand2 i_5095235(.A(n_13839), .B(n_13842), .Z(O0[3]));
	notech_nao3 i_4295236(.A(n_53871), .B(n_587), .C(n_53863), .Z(n_13842)
		);
	notech_nao3 i_3995237(.A(n_553), .B(n_53872), .C(n_53863), .Z(n_13839)
		);
	notech_nand2 i_5095239(.A(n_13863), .B(n_13866), .Z(O0[4]));
	notech_nao3 i_4295240(.A(n_53871), .B(n_588), .C(n_53863), .Z(n_13866)
		);
	notech_nao3 i_3995241(.A(n_554), .B(n_14529), .C(n_53863), .Z(n_13863)
		);
	notech_nand2 i_5095243(.A(n_13887), .B(n_13890), .Z(O0[5]));
	notech_nao3 i_4295244(.A(n_684), .B(n_589), .C(n_53863), .Z(n_13890));
	notech_nao3 i_3995245(.A(n_555), .B(n_53872), .C(n_53863), .Z(n_13887)
		);
	notech_nand2 i_5095247(.A(n_13911), .B(n_13914), .Z(O0[6]));
	notech_nao3 i_4295248(.A(n_53871), .B(n_590), .C(n_53863), .Z(n_13914)
		);
	notech_nao3 i_3995249(.A(n_556), .B(n_14529), .C(n_53863), .Z(n_13911)
		);
	notech_nand2 i_5095251(.A(n_13935), .B(n_13938), .Z(O0[7]));
	notech_nao3 i_4295252(.A(n_53871), .B(n_591), .C(n_53863), .Z(n_13938)
		);
	notech_nao3 i_3995253(.A(n_557), .B(n_53872), .C(n_53863), .Z(n_13935)
		);
	notech_nand2 i_5095255(.A(n_13959), .B(n_13962), .Z(O0[8]));
	notech_nao3 i_4295256(.A(n_53871), .B(n_592), .C(n_53861), .Z(n_13962)
		);
	notech_nao3 i_3995257(.A(n_558), .B(n_14529), .C(n_53861), .Z(n_13959)
		);
	notech_nand2 i_5095259(.A(n_13983), .B(n_13986), .Z(O0[9]));
	notech_nao3 i_4295260(.A(n_53871), .B(n_593), .C(n_53861), .Z(n_13986)
		);
	notech_nao3 i_3995261(.A(n_559), .B(n_53872), .C(n_53861), .Z(n_13983)
		);
	notech_nand2 i_5095263(.A(n_14007), .B(n_14010), .Z(O0[10]));
	notech_nao3 i_4295264(.A(n_53871), .B(n_594), .C(n_53861), .Z(n_14010)
		);
	notech_nao3 i_3995265(.A(n_560), .B(n_14529), .C(n_53861), .Z(n_14007)
		);
	notech_nand2 i_5095267(.A(n_14031), .B(n_14034), .Z(O0[11]));
	notech_nao3 i_4295268(.A(n_53871), .B(n_595), .C(n_53861), .Z(n_14034)
		);
	notech_nao3 i_3995269(.A(n_561), .B(n_53872), .C(n_53861), .Z(n_14031)
		);
	notech_nand2 i_5095271(.A(n_14055), .B(n_14058), .Z(O0[12]));
	notech_nao3 i_4295272(.A(n_53871), .B(n_596), .C(n_53861), .Z(n_14058)
		);
	notech_nao3 i_3995273(.A(n_562), .B(n_14529), .C(n_53861), .Z(n_14055)
		);
	notech_nand2 i_5095275(.A(n_14079), .B(n_14082), .Z(O0[13]));
	notech_nao3 i_4295276(.A(n_53871), .B(n_597), .C(n_53861), .Z(n_14082)
		);
	notech_nao3 i_3995277(.A(n_563), .B(n_53872), .C(n_53861), .Z(n_14079)
		);
	notech_nand2 i_5095279(.A(n_14103), .B(n_14106), .Z(O0[14]));
	notech_nao3 i_4295280(.A(n_53871), .B(n_598), .C(n_53861), .Z(n_14106)
		);
	notech_nao3 i_3995281(.A(n_564), .B(n_14529), .C(n_53861), .Z(n_14103)
		);
	notech_nand2 i_5095283(.A(n_14127), .B(n_14130), .Z(O0[15]));
	notech_nao3 i_4295284(.A(n_53871), .B(n_599), .C(n_53861), .Z(n_14130)
		);
	notech_nao3 i_3995285(.A(n_565), .B(n_53872), .C(n_53861), .Z(n_14127)
		);
	notech_nand2 i_5095287(.A(n_14151), .B(n_14154), .Z(O0[16]));
	notech_nao3 i_4295288(.A(n_684), .B(n_600), .C(n_53868), .Z(n_14154));
	notech_nao3 i_3995289(.A(n_566), .B(n_14529), .C(n_53868), .Z(n_14151)
		);
	notech_nand2 i_5095291(.A(n_14175), .B(n_14178), .Z(O0[17]));
	notech_nao3 i_4295292(.A(n_684), .B(n_601), .C(n_53868), .Z(n_14178));
	notech_nao3 i_3995293(.A(n_567), .B(n_53872), .C(n_53868), .Z(n_14175)
		);
	notech_nand2 i_5095295(.A(n_14199), .B(n_14202), .Z(O0[18]));
	notech_nao3 i_4295296(.A(n_684), .B(n_602), .C(n_53868), .Z(n_14202));
	notech_nao3 i_3995297(.A(n_568), .B(n_14529), .C(n_53868), .Z(n_14199)
		);
	notech_nand2 i_5095299(.A(n_14223), .B(n_14226), .Z(O0[19]));
	notech_nao3 i_4295300(.A(n_684), .B(n_603), .C(n_53868), .Z(n_14226));
	notech_nao3 i_3995301(.A(n_569), .B(n_53872), .C(n_53868), .Z(n_14223)
		);
	notech_nand2 i_5095303(.A(n_14247), .B(n_14250), .Z(O0[20]));
	notech_nao3 i_4295304(.A(n_684), .B(n_604), .C(n_53868), .Z(n_14250));
	notech_nao3 i_3995305(.A(n_570), .B(n_14529), .C(n_53868), .Z(n_14247)
		);
	notech_nand2 i_5095307(.A(n_14271), .B(n_14274), .Z(O0[21]));
	notech_nao3 i_4295308(.A(n_684), .B(n_605), .C(n_53868), .Z(n_14274));
	notech_nao3 i_3995309(.A(n_571), .B(n_14529), .C(n_53868), .Z(n_14271)
		);
	notech_nand2 i_5095311(.A(n_14295), .B(n_14298), .Z(O0[22]));
	notech_nao3 i_4295312(.A(n_684), .B(n_606), .C(n_53868), .Z(n_14298));
	notech_nao3 i_3995313(.A(n_572), .B(n_14529), .C(n_53868), .Z(n_14295)
		);
	notech_nand2 i_5095315(.A(n_14319), .B(n_14322), .Z(O0[23]));
	notech_nao3 i_4295316(.A(n_684), .B(n_607), .C(n_53868), .Z(n_14322));
	notech_nao3 i_3995317(.A(n_573), .B(n_53872), .C(n_53868), .Z(n_14319)
		);
	notech_nand2 i_5095319(.A(n_14343), .B(n_14346), .Z(O0[24]));
	notech_nao3 i_4295320(.A(n_684), .B(n_608), .C(n_53866), .Z(n_14346));
	notech_nao3 i_3995321(.A(n_574), .B(n_14529), .C(n_53866), .Z(n_14343)
		);
	notech_nand2 i_5095323(.A(n_14367), .B(n_14370), .Z(O0[25]));
	notech_nao3 i_4295324(.A(n_684), .B(n_609), .C(n_53866), .Z(n_14370));
	notech_nao3 i_3995325(.A(n_575), .B(n_53872), .C(n_53866), .Z(n_14367)
		);
	notech_nand2 i_5095327(.A(n_14391), .B(n_14394), .Z(O0[26]));
	notech_nao3 i_4295328(.A(n_684), .B(n_610), .C(n_53866), .Z(n_14394));
	notech_nao3 i_3995329(.A(n_576), .B(n_14529), .C(n_53866), .Z(n_14391)
		);
	notech_nand2 i_5095331(.A(n_14415), .B(n_14418), .Z(O0[27]));
	notech_nao3 i_4295332(.A(n_684), .B(n_611), .C(n_53866), .Z(n_14418));
	notech_nao3 i_3995333(.A(n_577), .B(n_53872), .C(n_53866), .Z(n_14415)
		);
	notech_nand2 i_5095335(.A(n_14439), .B(n_14442), .Z(O0[28]));
	notech_nao3 i_4295336(.A(n_684), .B(n_612), .C(n_53866), .Z(n_14442));
	notech_nao3 i_3995337(.A(n_578), .B(n_14529), .C(n_53866), .Z(n_14439)
		);
	notech_nand2 i_5095339(.A(n_14463), .B(n_14466), .Z(O0[29]));
	notech_nao3 i_4295340(.A(n_684), .B(n_613), .C(n_53866), .Z(n_14466));
	notech_nao3 i_3995341(.A(n_579), .B(n_53872), .C(n_53866), .Z(n_14463)
		);
	notech_nand2 i_5095343(.A(n_14487), .B(n_14490), .Z(O0[30]));
	notech_nao3 i_4295344(.A(n_684), .B(n_614), .C(n_53866), .Z(n_14490));
	notech_nao3 i_3995345(.A(n_580), .B(n_14529), .C(n_53866), .Z(n_14487)
		);
	notech_inv i_395346(.A(n_684), .Z(n_14529));
	notech_nand2 i_5095347(.A(n_14511), .B(n_14514), .Z(O0[31]));
	notech_nao3 i_4295348(.A(n_684), .B(n_615), .C(n_53866), .Z(n_14514));
	notech_nao3 i_3995349(.A(n_581), .B(n_53872), .C(n_53866), .Z(n_14511)
		);
endmodule
module AWMUX_16_32_3(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_4(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_5(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_6(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_7(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module vliw(clk, rstn, instrc, ie, readio_data, io_add, writeio_data, writeio_req
		, readio_req, writeio_ack, readio_ack, read_reqs, read_ack, read_data
		, over_seg, cr3, cr2, icr2, cr1, cr0, write_reqs, write_ack, write_data
		, Daddr, write_sz, read_sz, cs, add_src, from_acu, to_acu, seg_src
		, pg_en, ready_vliw, valid_op, imm, lenpc, pc_out, pc_req, opz, reps
		, adz, flush_tlb, flush_Dtlb, terminate, start_up, pg_fault, ipg_fault
		, wr_fault, pt_fault, repbytecache);

	input clk;
	input rstn;
	input [127:0] instrc;
	output ie;
	input [31:0] readio_data;
	output [31:0] io_add;
	output [31:0] writeio_data;
	output writeio_req;
	output readio_req;
	input writeio_ack;
	input readio_ack;
	output read_reqs;
	input read_ack;
	input [31:0] read_data;
	input [5:0] over_seg;
	output [31:0] cr3;
	input [31:0] cr2;
	input [31:0] icr2;
	output [31:0] cr1;
	output [31:0] cr0;
	output write_reqs;
	input write_ack;
	output [31:0] write_data;
	output [31:0] Daddr;
	output [1:0] write_sz;
	output [1:0] read_sz;
	output [31:0] cs;
	input [31:0] add_src;
	input [7:0] from_acu;
	output [63:0] to_acu;
	input [2:0] seg_src;
	output pg_en;
	output ready_vliw;
	input valid_op;
	input [63:0] imm;
	input [31:0] lenpc;
	output [31:0] pc_out;
	output pc_req;
	input [2:0] opz;
	input [2:0] reps;
	input adz;
	output flush_tlb;
	output flush_Dtlb;
	output terminate;
	input start_up;
	input pg_fault;
	input ipg_fault;
	input wr_fault;
	input pt_fault;
	output repbytecache;

	wire [4:0] fsm;
	wire [31:0] opa;
	wire [31:0] opc;
	wire [31:0] nbus_11295;
	wire [31:0] opd;
	wire [3:0] calc_sz;
	wire [31:0] gs;
	wire [31:0] sav_edi;
	wire [31:0] sav_esi;
	wire [31:0] sav_epc;
	wire [31:0] sav_esp;
	wire [31:0] sav_ecx;
	wire [31:0] temp_sp;
	wire [1:0] sav_cs;
	wire [31:0] cr2_reg;
	wire [31:0] nbus_14521;
	wire [4:0] vliw_pc;
	wire [31:0] Daddrgs;
	wire [2:0] mask8b;
	wire [4:0] fsmf;
	wire [31:0] temp_ss;
	wire [31:0] errco;
	wire [1:0] pipe_mul;
	wire [63:0] to_acu100236;
	wire [31:0] nbus_11360;
	wire [31:0] nbus_11328;
	wire [31:0] nbus_11310;
	wire [31:0] Daddrs_8;
	wire [31:0] write_data_33;
	wire [31:0] write_data_32;
	wire [31:0] write_data_31;
	wire [31:0] write_data_30;
	wire [31:0] write_data_29;
	wire [31:0] write_data_28;
	wire [31:0] write_data_27;
	wire [31:0] write_data_26;
	wire [31:0] write_data_25;
	wire [31:0] opc_14;
	wire [31:0] opc_10;
	wire [31:0] Daddrs_3;
	wire [31:0] Daddrs_1;
	wire [63:0] divr_1;
	wire [31:0] regs_4_2;
	wire [31:0] add_len_pc;
	wire [31:0] opa_0;
	wire [31:0] resa_arithbox;
	wire [16:0] nbus_167;
	wire [32:0] nbus_166;
	wire [16:0] nbus_165;
	wire [32:0] nbus_164;
	wire [16:0] nbus_163;
	wire [32:0] nbus_162;
	wire [16:0] nbus_161;
	wire [32:0] nbus_160;
	wire [8:0] nbus_159;
	wire [16:0] nbus_158;
	wire [32:0] nbus_157;
	wire [63:0] mul64;
	wire [31:0] add_len_pc32;
	wire [31:0] resb_shift4box;
	wire [31:0] resa_shift4box;
	wire [31:0] resb_shiftbox;
	wire [31:0] resa_shiftbox;
	wire [63:0] tsc;
	wire [3:0] all_cnt;
	wire [31:0] regs_14;
	wire [31:0] regs_12;
	wire [31:0] regs_11;
	wire [31:0] regs_10;
	wire [31:0] regs_8;
	wire [31:0] regs_7;
	wire [31:0] regs_6;
	wire [31:0] regs_5;
	wire [31:0] regs_4;
	wire [31:0] regs_3;
	wire [31:0] opb;
	wire [31:0] regs_2;
	wire [31:0] ecx;
	wire [63:0] divq;
	wire [63:0] divr;
	wire [31:0] regs_0;
	wire [31:0] ldtr;
	wire [31:0] gdtr;
	wire [31:0] idtr;
	wire [31:0] desc;



	notech_inv i_16138(.A(n_62891), .Z(n_62892));
	notech_inv i_16137(.A(\opcode[3] ), .Z(n_62891));
	notech_inv i_16116(.A(n_62869), .Z(n_62870));
	notech_inv i_16115(.A(\opcode[0] ), .Z(n_62869));
	notech_inv i_16114(.A(n_62867), .Z(n_62868));
	notech_inv i_16113(.A(n_62870), .Z(n_62867));
	notech_inv i_16110(.A(n_62863), .Z(n_62864));
	notech_inv i_16109(.A(n_62854), .Z(n_62863));
	notech_inv i_16106(.A(n_62859), .Z(n_62860));
	notech_inv i_16105(.A(n_62846), .Z(n_62859));
	notech_inv i_16104(.A(n_62857), .Z(n_62858));
	notech_inv i_16103(.A(n_62842), .Z(n_62857));
	notech_inv i_16102(.A(n_62855), .Z(n_62856));
	notech_inv i_16101(.A(n_62840), .Z(n_62855));
	notech_inv i_16100(.A(n_62853), .Z(n_62854));
	notech_inv i_16099(.A(n_62856), .Z(n_62853));
	notech_inv i_16096(.A(n_62849), .Z(n_62850));
	notech_inv i_16095(.A(n_62834), .Z(n_62849));
	notech_inv i_16094(.A(n_62847), .Z(n_62848));
	notech_inv i_16093(.A(n_62832), .Z(n_62847));
	notech_inv i_16092(.A(n_62845), .Z(n_62846));
	notech_inv i_16091(.A(n_62848), .Z(n_62845));
	notech_inv i_16090(.A(n_62843), .Z(n_62844));
	notech_inv i_16089(.A(n_62830), .Z(n_62843));
	notech_inv i_16088(.A(n_62841), .Z(n_62842));
	notech_inv i_16087(.A(n_62844), .Z(n_62841));
	notech_inv i_16086(.A(n_62839), .Z(n_62840));
	notech_inv i_16085(.A(n_62858), .Z(n_62839));
	notech_inv i_16082(.A(n_62835), .Z(n_62836));
	notech_inv i_16081(.A(\opcode[1] ), .Z(n_62835));
	notech_inv i_16080(.A(n_62833), .Z(n_62834));
	notech_inv i_16079(.A(n_62836), .Z(n_62833));
	notech_inv i_16078(.A(n_62831), .Z(n_62832));
	notech_inv i_16077(.A(n_62850), .Z(n_62831));
	notech_inv i_16076(.A(n_62829), .Z(n_62830));
	notech_inv i_16075(.A(n_62860), .Z(n_62829));
	notech_inv i_16072(.A(n_62825), .Z(n_62826));
	notech_inv i_16071(.A(n_62818), .Z(n_62825));
	notech_inv i_16070(.A(n_62823), .Z(n_62824));
	notech_inv i_16069(.A(n_62810), .Z(n_62823));
	notech_inv i_16068(.A(n_62821), .Z(n_62822));
	notech_inv i_16067(.A(n_62804), .Z(n_62821));
	notech_inv i_16066(.A(n_62819), .Z(n_62820));
	notech_inv i_16065(.A(n_62802), .Z(n_62819));
	notech_inv i_16064(.A(n_62817), .Z(n_62818));
	notech_inv i_16063(.A(n_62798), .Z(n_62817));
	notech_inv i_16062(.A(n_62815), .Z(n_62816));
	notech_inv i_16061(.A(n_62790), .Z(n_62815));
	notech_inv i_16060(.A(n_62813), .Z(n_62814));
	notech_inv i_16059(.A(n_62786), .Z(n_62813));
	notech_inv i_16058(.A(n_62811), .Z(n_62812));
	notech_inv i_16057(.A(n_62784), .Z(n_62811));
	notech_inv i_16056(.A(n_62809), .Z(n_62810));
	notech_inv i_16055(.A(n_62812), .Z(n_62809));
	notech_inv i_16054(.A(n_62807), .Z(n_62808));
	notech_inv i_16053(.A(n_62780), .Z(n_62807));
	notech_inv i_16052(.A(n_62805), .Z(n_62806));
	notech_inv i_16051(.A(n_62778), .Z(n_62805));
	notech_inv i_16050(.A(n_62803), .Z(n_62804));
	notech_inv i_16049(.A(n_62806), .Z(n_62803));
	notech_inv i_16048(.A(n_62801), .Z(n_62802));
	notech_inv i_16047(.A(n_62776), .Z(n_62801));
	notech_inv i_16044(.A(n_62797), .Z(n_62798));
	notech_inv i_16043(.A(n_62820), .Z(n_62797));
	notech_inv i_16040(.A(n_62793), .Z(n_62794));
	notech_inv i_16039(.A(n_62772), .Z(n_62793));
	notech_inv i_16038(.A(n_62791), .Z(n_62792));
	notech_inv i_16037(.A(n_62770), .Z(n_62791));
	notech_inv i_16036(.A(n_62789), .Z(n_62790));
	notech_inv i_16035(.A(n_62792), .Z(n_62789));
	notech_inv i_16034(.A(n_62787), .Z(n_62788));
	notech_inv i_16033(.A(n_62768), .Z(n_62787));
	notech_inv i_16032(.A(n_62785), .Z(n_62786));
	notech_inv i_16031(.A(n_62788), .Z(n_62785));
	notech_inv i_16030(.A(n_62783), .Z(n_62784));
	notech_inv i_16029(.A(n_62814), .Z(n_62783));
	notech_inv i_16028(.A(n_62781), .Z(n_62782));
	notech_inv i_16027(.A(n_62766), .Z(n_62781));
	notech_inv i_16026(.A(n_62779), .Z(n_62780));
	notech_inv i_16025(.A(n_62782), .Z(n_62779));
	notech_inv i_16024(.A(n_62777), .Z(n_62778));
	notech_inv i_16023(.A(n_62808), .Z(n_62777));
	notech_inv i_16022(.A(n_62775), .Z(n_62776));
	notech_inv i_16021(.A(n_62822), .Z(n_62775));
	notech_inv i_16018(.A(n_62771), .Z(n_62772));
	notech_inv i_16017(.A(\opcode[2] ), .Z(n_62771));
	notech_inv i_16016(.A(n_62769), .Z(n_62770));
	notech_inv i_16015(.A(n_62794), .Z(n_62769));
	notech_inv i_16014(.A(n_62767), .Z(n_62768));
	notech_inv i_16013(.A(n_62816), .Z(n_62767));
	notech_inv i_16012(.A(n_62765), .Z(n_62766));
	notech_inv i_16011(.A(n_62824), .Z(n_62765));
	notech_inv i_16008(.A(n_62761), .Z(n_62762));
	notech_inv i_16007(.A(n_62748), .Z(n_62761));
	notech_inv i_16006(.A(n_62759), .Z(n_62760));
	notech_inv i_16005(.A(n_62736), .Z(n_62759));
	notech_inv i_16004(.A(n_62757), .Z(n_62758));
	notech_inv i_16003(.A(n_62726), .Z(n_62757));
	notech_inv i_16002(.A(n_62755), .Z(n_62756));
	notech_inv i_16001(.A(n_62718), .Z(n_62755));
	notech_inv i_16000(.A(n_62753), .Z(n_62754));
	notech_inv i_15999(.A(n_62712), .Z(n_62753));
	notech_inv i_15998(.A(n_62751), .Z(n_62752));
	notech_inv i_15997(.A(n_62708), .Z(n_62751));
	notech_inv i_15996(.A(n_62749), .Z(n_62750));
	notech_inv i_15995(.A(n_62706), .Z(n_62749));
	notech_inv i_15994(.A(n_62747), .Z(n_62748));
	notech_inv i_15993(.A(n_62750), .Z(n_62747));
	notech_inv i_15990(.A(n_62743), .Z(n_62744));
	notech_inv i_15989(.A(n_62688), .Z(n_62743));
	notech_inv i_15988(.A(n_62741), .Z(n_62742));
	notech_inv i_15987(.A(n_62682), .Z(n_62741));
	notech_inv i_15986(.A(n_62739), .Z(n_62740));
	notech_inv i_15985(.A(n_62678), .Z(n_62739));
	notech_inv i_15984(.A(n_62737), .Z(n_62738));
	notech_inv i_15983(.A(n_62676), .Z(n_62737));
	notech_inv i_15982(.A(n_62735), .Z(n_62736));
	notech_inv i_15981(.A(n_62738), .Z(n_62735));
	notech_inv i_15980(.A(n_62733), .Z(n_62734));
	notech_inv i_15979(.A(n_62668), .Z(n_62733));
	notech_inv i_15978(.A(n_62731), .Z(n_62732));
	notech_inv i_15977(.A(n_62662), .Z(n_62731));
	notech_inv i_15976(.A(n_62729), .Z(n_62730));
	notech_inv i_15975(.A(n_62658), .Z(n_62729));
	notech_inv i_15974(.A(n_62727), .Z(n_62728));
	notech_inv i_15973(.A(n_62656), .Z(n_62727));
	notech_inv i_15972(.A(n_62725), .Z(n_62726));
	notech_inv i_15971(.A(n_62728), .Z(n_62725));
	notech_inv i_15970(.A(n_62723), .Z(n_62724));
	notech_inv i_15969(.A(n_62650), .Z(n_62723));
	notech_inv i_15968(.A(n_62721), .Z(n_62722));
	notech_inv i_15967(.A(n_62646), .Z(n_62721));
	notech_inv i_15966(.A(n_62719), .Z(n_62720));
	notech_inv i_15965(.A(n_62644), .Z(n_62719));
	notech_inv i_15964(.A(n_62717), .Z(n_62718));
	notech_inv i_15963(.A(n_62720), .Z(n_62717));
	notech_inv i_15962(.A(n_62715), .Z(n_62716));
	notech_inv i_15961(.A(n_62640), .Z(n_62715));
	notech_inv i_15960(.A(n_62713), .Z(n_62714));
	notech_inv i_15959(.A(n_62638), .Z(n_62713));
	notech_inv i_15958(.A(n_62711), .Z(n_62712));
	notech_inv i_15957(.A(n_62714), .Z(n_62711));
	notech_inv i_15956(.A(n_62709), .Z(n_62710));
	notech_inv i_15955(.A(n_62636), .Z(n_62709));
	notech_inv i_15954(.A(n_62707), .Z(n_62708));
	notech_inv i_15953(.A(n_62710), .Z(n_62707));
	notech_inv i_15952(.A(n_62705), .Z(n_62706));
	notech_inv i_15951(.A(n_62752), .Z(n_62705));
	notech_inv i_15940(.A(n_62693), .Z(n_62694));
	notech_inv i_15939(.A(n_62610), .Z(n_62693));
	notech_inv i_15938(.A(n_62691), .Z(n_62692));
	notech_inv i_15937(.A(n_62606), .Z(n_62691));
	notech_inv i_15936(.A(n_62689), .Z(n_62690));
	notech_inv i_15935(.A(n_62604), .Z(n_62689));
	notech_inv i_15934(.A(n_62687), .Z(n_62688));
	notech_inv i_15933(.A(n_62690), .Z(n_62687));
	notech_inv i_15932(.A(n_62685), .Z(n_62686));
	notech_inv i_15931(.A(n_62600), .Z(n_62685));
	notech_inv i_15930(.A(n_62683), .Z(n_62684));
	notech_inv i_15929(.A(n_62598), .Z(n_62683));
	notech_inv i_15928(.A(n_62681), .Z(n_62682));
	notech_inv i_15927(.A(n_62684), .Z(n_62681));
	notech_inv i_15926(.A(n_62679), .Z(n_62680));
	notech_inv i_15925(.A(n_62596), .Z(n_62679));
	notech_inv i_15924(.A(n_62677), .Z(n_62678));
	notech_inv i_15923(.A(n_62680), .Z(n_62677));
	notech_inv i_15922(.A(n_62675), .Z(n_62676));
	notech_inv i_15921(.A(n_62740), .Z(n_62675));
	notech_inv i_15920(.A(n_62673), .Z(n_62674));
	notech_inv i_15919(.A(n_62590), .Z(n_62673));
	notech_inv i_15918(.A(n_62671), .Z(n_62672));
	notech_inv i_15917(.A(n_62586), .Z(n_62671));
	notech_inv i_15916(.A(n_62669), .Z(n_62670));
	notech_inv i_15915(.A(n_62584), .Z(n_62669));
	notech_inv i_15914(.A(n_62667), .Z(n_62668));
	notech_inv i_15913(.A(n_62670), .Z(n_62667));
	notech_inv i_15912(.A(n_62665), .Z(n_62666));
	notech_inv i_15911(.A(n_62580), .Z(n_62665));
	notech_inv i_15910(.A(n_62663), .Z(n_62664));
	notech_inv i_15909(.A(n_62578), .Z(n_62663));
	notech_inv i_15908(.A(n_62661), .Z(n_62662));
	notech_inv i_15907(.A(n_62664), .Z(n_62661));
	notech_inv i_15906(.A(n_62659), .Z(n_62660));
	notech_inv i_15905(.A(n_62576), .Z(n_62659));
	notech_inv i_15904(.A(n_62657), .Z(n_62658));
	notech_inv i_15903(.A(n_62660), .Z(n_62657));
	notech_inv i_15902(.A(n_62655), .Z(n_62656));
	notech_inv i_15901(.A(n_62730), .Z(n_62655));
	notech_inv i_15900(.A(n_62653), .Z(n_62654));
	notech_inv i_15899(.A(n_62572), .Z(n_62653));
	notech_inv i_15898(.A(n_62651), .Z(n_62652));
	notech_inv i_15897(.A(n_62570), .Z(n_62651));
	notech_inv i_15896(.A(n_62649), .Z(n_62650));
	notech_inv i_15895(.A(n_62652), .Z(n_62649));
	notech_inv i_15894(.A(n_62647), .Z(n_62648));
	notech_inv i_15893(.A(n_62568), .Z(n_62647));
	notech_inv i_15892(.A(n_62645), .Z(n_62646));
	notech_inv i_15891(.A(n_62648), .Z(n_62645));
	notech_inv i_15890(.A(n_62643), .Z(n_62644));
	notech_inv i_15889(.A(n_62722), .Z(n_62643));
	notech_inv i_15888(.A(n_62641), .Z(n_62642));
	notech_inv i_15887(.A(n_62566), .Z(n_62641));
	notech_inv i_15886(.A(n_62639), .Z(n_62640));
	notech_inv i_15885(.A(n_62642), .Z(n_62639));
	notech_inv i_15884(.A(n_62637), .Z(n_62638));
	notech_inv i_15883(.A(n_62716), .Z(n_62637));
	notech_inv i_15882(.A(n_62635), .Z(n_62636));
	notech_inv i_15881(.A(n_62754), .Z(n_62635));
	notech_inv i_15880(.A(n_62633), .Z(n_62634));
	notech_inv i_15879(.A(n_62560), .Z(n_62633));
	notech_inv i_15860(.A(n_62613), .Z(n_62614));
	notech_inv i_15859(.A(n_62542), .Z(n_62613));
	notech_inv i_15858(.A(n_62611), .Z(n_62612));
	notech_inv i_15857(.A(n_62540), .Z(n_62611));
	notech_inv i_15856(.A(n_62609), .Z(n_62610));
	notech_inv i_15855(.A(n_62612), .Z(n_62609));
	notech_inv i_15854(.A(n_62607), .Z(n_62608));
	notech_inv i_15853(.A(n_62538), .Z(n_62607));
	notech_inv i_15852(.A(n_62605), .Z(n_62606));
	notech_inv i_15851(.A(n_62608), .Z(n_62605));
	notech_inv i_15850(.A(n_62603), .Z(n_62604));
	notech_inv i_15849(.A(n_62692), .Z(n_62603));
	notech_inv i_15848(.A(n_62601), .Z(n_62602));
	notech_inv i_15847(.A(n_62536), .Z(n_62601));
	notech_inv i_15846(.A(n_62599), .Z(n_62600));
	notech_inv i_15845(.A(n_62602), .Z(n_62599));
	notech_inv i_15844(.A(n_62597), .Z(n_62598));
	notech_inv i_15843(.A(n_62686), .Z(n_62597));
	notech_inv i_15842(.A(n_62595), .Z(n_62596));
	notech_inv i_15841(.A(n_62742), .Z(n_62595));
	notech_inv i_15840(.A(n_62593), .Z(n_62594));
	notech_inv i_15839(.A(n_62532), .Z(n_62593));
	notech_inv i_15838(.A(n_62591), .Z(n_62592));
	notech_inv i_15837(.A(n_62530), .Z(n_62591));
	notech_inv i_15836(.A(n_62589), .Z(n_62590));
	notech_inv i_15835(.A(n_62592), .Z(n_62589));
	notech_inv i_15834(.A(n_62587), .Z(n_62588));
	notech_inv i_15833(.A(n_62528), .Z(n_62587));
	notech_inv i_15832(.A(n_62585), .Z(n_62586));
	notech_inv i_15831(.A(n_62588), .Z(n_62585));
	notech_inv i_15830(.A(n_62583), .Z(n_62584));
	notech_inv i_15829(.A(n_62672), .Z(n_62583));
	notech_inv i_15828(.A(n_62581), .Z(n_62582));
	notech_inv i_15827(.A(n_62526), .Z(n_62581));
	notech_inv i_15826(.A(n_62579), .Z(n_62580));
	notech_inv i_15825(.A(n_62582), .Z(n_62579));
	notech_inv i_15824(.A(n_62577), .Z(n_62578));
	notech_inv i_15823(.A(n_62666), .Z(n_62577));
	notech_inv i_15822(.A(n_62575), .Z(n_62576));
	notech_inv i_15821(.A(n_62732), .Z(n_62575));
	notech_inv i_15820(.A(n_62573), .Z(n_62574));
	notech_inv i_15819(.A(n_62524), .Z(n_62573));
	notech_inv i_15818(.A(n_62571), .Z(n_62572));
	notech_inv i_15817(.A(n_62574), .Z(n_62571));
	notech_inv i_15816(.A(n_62569), .Z(n_62570));
	notech_inv i_15815(.A(n_62654), .Z(n_62569));
	notech_inv i_15814(.A(n_62567), .Z(n_62568));
	notech_inv i_15813(.A(n_62724), .Z(n_62567));
	notech_inv i_15812(.A(n_62565), .Z(n_62566));
	notech_inv i_15811(.A(n_62756), .Z(n_62565));
	notech_inv i_15810(.A(n_62563), .Z(n_62564));
	notech_inv i_15809(.A(n_62518), .Z(n_62563));
	notech_inv i_15808(.A(n_62561), .Z(n_62562));
	notech_inv i_15807(.A(n_62490), .Z(n_62561));
	notech_inv i_15806(.A(n_62559), .Z(n_62560));
	notech_inv i_15805(.A(n_62562), .Z(n_62559));
	notech_inv i_15790(.A(n_62543), .Z(n_62544));
	notech_inv i_15789(.A(n_62448), .Z(n_62543));
	notech_inv i_15788(.A(n_62541), .Z(n_62542));
	notech_inv i_15787(.A(n_62544), .Z(n_62541));
	notech_inv i_15786(.A(n_62539), .Z(n_62540));
	notech_inv i_15785(.A(n_62614), .Z(n_62539));
	notech_inv i_15784(.A(n_62537), .Z(n_62538));
	notech_inv i_15783(.A(n_62694), .Z(n_62537));
	notech_inv i_15782(.A(n_62535), .Z(n_62536));
	notech_inv i_15781(.A(n_62744), .Z(n_62535));
	notech_inv i_15780(.A(n_62533), .Z(n_62534));
	notech_inv i_15779(.A(n_62432), .Z(n_62533));
	notech_inv i_15778(.A(n_62531), .Z(n_62532));
	notech_inv i_15777(.A(n_62534), .Z(n_62531));
	notech_inv i_15776(.A(n_62529), .Z(n_62530));
	notech_inv i_15775(.A(n_62594), .Z(n_62529));
	notech_inv i_15774(.A(n_62527), .Z(n_62528));
	notech_inv i_15773(.A(n_62674), .Z(n_62527));
	notech_inv i_15772(.A(n_62525), .Z(n_62526));
	notech_inv i_15771(.A(n_62734), .Z(n_62525));
	notech_inv i_15770(.A(n_62523), .Z(n_62524));
	notech_inv i_15769(.A(n_62758), .Z(n_62523));
	notech_inv i_15764(.A(n_62517), .Z(n_62518));
	notech_inv i_15763(.A(clk), .Z(n_62517));
	notech_inv i_15735(.A(n_62489), .Z(n_62490));
	notech_inv i_15734(.A(n_62564), .Z(n_62489));
	notech_inv i_15693(.A(n_62447), .Z(n_62448));
	notech_inv i_15692(.A(n_62634), .Z(n_62447));
	notech_inv i_15677(.A(n_62431), .Z(n_62432));
	notech_inv i_15676(.A(n_62760), .Z(n_62431));
	notech_inv i_14548(.A(n_61466), .Z(n_61600));
	notech_inv i_14547(.A(n_61466), .Z(n_61599));
	notech_inv i_14546(.A(n_61466), .Z(n_61598));
	notech_inv i_14545(.A(n_61466), .Z(n_61597));
	notech_inv i_14543(.A(n_61466), .Z(n_61595));
	notech_inv i_14542(.A(n_61466), .Z(n_61594));
	notech_inv i_14541(.A(n_61466), .Z(n_61593));
	notech_inv i_14540(.A(n_61466), .Z(n_61592));
	notech_inv i_14537(.A(n_61466), .Z(n_61589));
	notech_inv i_14536(.A(n_61466), .Z(n_61588));
	notech_inv i_14535(.A(n_61466), .Z(n_61587));
	notech_inv i_14534(.A(n_61466), .Z(n_61586));
	notech_inv i_14532(.A(n_61466), .Z(n_61584));
	notech_inv i_14531(.A(n_61466), .Z(n_61583));
	notech_inv i_14530(.A(n_61466), .Z(n_61582));
	notech_inv i_14529(.A(n_61466), .Z(n_61581));
	notech_inv i_14526(.A(n_61569), .Z(n_61578));
	notech_inv i_14525(.A(n_61569), .Z(n_61577));
	notech_inv i_14524(.A(n_61569), .Z(n_61576));
	notech_inv i_14523(.A(n_61569), .Z(n_61575));
	notech_inv i_14521(.A(n_61569), .Z(n_61573));
	notech_inv i_14520(.A(n_61569), .Z(n_61572));
	notech_inv i_14519(.A(n_61569), .Z(n_61571));
	notech_inv i_14518(.A(n_61569), .Z(n_61570));
	notech_inv i_14517(.A(n_61586), .Z(n_61569));
	notech_inv i_14515(.A(n_61569), .Z(n_61567));
	notech_inv i_14514(.A(n_61569), .Z(n_61566));
	notech_inv i_14513(.A(n_61569), .Z(n_61565));
	notech_inv i_14512(.A(n_61569), .Z(n_61564));
	notech_inv i_14510(.A(n_61569), .Z(n_61562));
	notech_inv i_14509(.A(n_61569), .Z(n_61561));
	notech_inv i_14508(.A(n_61569), .Z(n_61560));
	notech_inv i_14507(.A(n_61569), .Z(n_61559));
	notech_inv i_14503(.A(n_61546), .Z(n_61555));
	notech_inv i_14502(.A(n_61546), .Z(n_61554));
	notech_inv i_14501(.A(n_61546), .Z(n_61553));
	notech_inv i_14500(.A(n_61546), .Z(n_61552));
	notech_inv i_14498(.A(n_61546), .Z(n_61550));
	notech_inv i_14497(.A(n_61546), .Z(n_61549));
	notech_inv i_14496(.A(n_61546), .Z(n_61548));
	notech_inv i_14495(.A(n_61546), .Z(n_61547));
	notech_inv i_14494(.A(n_61592), .Z(n_61546));
	notech_inv i_14492(.A(n_61546), .Z(n_61544));
	notech_inv i_14491(.A(n_61546), .Z(n_61543));
	notech_inv i_14490(.A(n_61546), .Z(n_61542));
	notech_inv i_14489(.A(n_61546), .Z(n_61541));
	notech_inv i_14487(.A(n_61546), .Z(n_61539));
	notech_inv i_14486(.A(n_61546), .Z(n_61538));
	notech_inv i_14485(.A(n_61546), .Z(n_61537));
	notech_inv i_14484(.A(n_61546), .Z(n_61536));
	notech_inv i_14480(.A(n_61524), .Z(n_61533));
	notech_inv i_14479(.A(n_61524), .Z(n_61532));
	notech_inv i_14478(.A(n_61524), .Z(n_61531));
	notech_inv i_14477(.A(n_61524), .Z(n_61530));
	notech_inv i_14475(.A(n_61524), .Z(n_61528));
	notech_inv i_14474(.A(n_61524), .Z(n_61527));
	notech_inv i_14473(.A(n_61524), .Z(n_61526));
	notech_inv i_14472(.A(n_61524), .Z(n_61525));
	notech_inv i_14471(.A(n_61592), .Z(n_61524));
	notech_inv i_14469(.A(n_61524), .Z(n_61522));
	notech_inv i_14468(.A(n_61524), .Z(n_61521));
	notech_inv i_14467(.A(n_61524), .Z(n_61520));
	notech_inv i_14466(.A(n_61524), .Z(n_61519));
	notech_inv i_14464(.A(n_61524), .Z(n_61517));
	notech_inv i_14463(.A(n_61524), .Z(n_61516));
	notech_inv i_14462(.A(n_61524), .Z(n_61515));
	notech_inv i_14461(.A(n_61524), .Z(n_61514));
	notech_inv i_14457(.A(n_61501), .Z(n_61510));
	notech_inv i_14456(.A(n_61501), .Z(n_61509));
	notech_inv i_14455(.A(n_61501), .Z(n_61508));
	notech_inv i_14454(.A(n_61501), .Z(n_61507));
	notech_inv i_14452(.A(n_61501), .Z(n_61505));
	notech_inv i_14451(.A(n_61501), .Z(n_61504));
	notech_inv i_14450(.A(n_61501), .Z(n_61503));
	notech_inv i_14449(.A(n_61501), .Z(n_61502));
	notech_inv i_14448(.A(n_61586), .Z(n_61501));
	notech_inv i_14446(.A(n_61501), .Z(n_61499));
	notech_inv i_14445(.A(n_61501), .Z(n_61498));
	notech_inv i_14444(.A(n_61501), .Z(n_61497));
	notech_inv i_14443(.A(n_61501), .Z(n_61496));
	notech_inv i_14441(.A(n_61501), .Z(n_61494));
	notech_inv i_14440(.A(n_61501), .Z(n_61493));
	notech_inv i_14439(.A(n_61501), .Z(n_61492));
	notech_inv i_14438(.A(n_61501), .Z(n_61491));
	notech_inv i_14435(.A(n_61479), .Z(n_61488));
	notech_inv i_14434(.A(n_61479), .Z(n_61487));
	notech_inv i_14433(.A(n_61479), .Z(n_61486));
	notech_inv i_14432(.A(n_61479), .Z(n_61485));
	notech_inv i_14430(.A(n_61479), .Z(n_61483));
	notech_inv i_14429(.A(n_61479), .Z(n_61482));
	notech_inv i_14428(.A(n_61479), .Z(n_61481));
	notech_inv i_14427(.A(n_61479), .Z(n_61480));
	notech_inv i_14426(.A(n_61586), .Z(n_61479));
	notech_inv i_14424(.A(n_61479), .Z(n_61477));
	notech_inv i_14423(.A(n_61479), .Z(n_61476));
	notech_inv i_14422(.A(n_61479), .Z(n_61475));
	notech_inv i_14421(.A(n_61479), .Z(n_61474));
	notech_inv i_14419(.A(n_61479), .Z(n_61472));
	notech_inv i_14418(.A(n_61479), .Z(n_61471));
	notech_inv i_14417(.A(n_61479), .Z(n_61470));
	notech_inv i_14416(.A(n_61479), .Z(n_61469));
	notech_inv i_14413(.A(rstn), .Z(n_61466));
	notech_inv i_14133(.A(n_61170), .Z(n_61175));
	notech_inv i_14128(.A(n_61170), .Z(n_61171));
	notech_inv i_14127(.A(fsm[2]), .Z(n_61170));
	notech_inv i_14125(.A(n_61159), .Z(n_61167));
	notech_inv i_14123(.A(n_61159), .Z(n_61165));
	notech_inv i_14118(.A(n_61159), .Z(n_61161));
	notech_inv i_14117(.A(n_61159), .Z(n_61160));
	notech_inv i_14116(.A(fsm[4]), .Z(n_61159));
	notech_inv i_14114(.A(n_272491901), .Z(n_61156));
	notech_inv i_14111(.A(n_272491901), .Z(n_61154));
	notech_inv i_14108(.A(n_272491901), .Z(n_61151));
	notech_inv i_14106(.A(n_272491901), .Z(n_61149));
	notech_inv i_14102(.A(n_61129), .Z(n_61145));
	notech_inv i_14100(.A(n_61129), .Z(n_61143));
	notech_inv i_14099(.A(n_61129), .Z(n_61142));
	notech_inv i_14094(.A(n_61129), .Z(n_61138));
	notech_inv i_14092(.A(n_61129), .Z(n_61136));
	notech_inv i_14088(.A(n_61129), .Z(n_61133));
	notech_inv i_14086(.A(n_61129), .Z(n_61131));
	notech_inv i_14085(.A(n_61129), .Z(n_61130));
	notech_inv i_14084(.A(pg_fault), .Z(n_61129));
	notech_inv i_14075(.A(n_61102), .Z(n_61117));
	notech_inv i_14072(.A(n_61102), .Z(n_61115));
	notech_inv i_14067(.A(n_61102), .Z(n_61110));
	notech_inv i_14066(.A(n_61102), .Z(n_61109));
	notech_inv i_14059(.A(n_61102), .Z(n_61103));
	notech_inv i_14058(.A(n_32855), .Z(n_61102));
	notech_inv i_13944(.A(n_60985), .Z(n_60986));
	notech_inv i_13943(.A(n_32730), .Z(n_60985));
	notech_inv i_13933(.A(n_60974), .Z(n_60975));
	notech_inv i_13932(.A(instrc[122]), .Z(n_60974));
	notech_inv i_13928(.A(n_60963), .Z(n_60970));
	notech_inv i_13927(.A(n_60963), .Z(n_60969));
	notech_inv i_13922(.A(n_60963), .Z(n_60964));
	notech_inv i_13920(.A(n_2547), .Z(n_60963));
	notech_inv i_13917(.A(n_60952), .Z(n_60959));
	notech_inv i_13916(.A(n_60952), .Z(n_60958));
	notech_inv i_13910(.A(n_60952), .Z(n_60953));
	notech_inv i_13909(.A(n_2788), .Z(n_60952));
	notech_inv i_13907(.A(n_60923), .Z(n_60949));
	notech_inv i_13904(.A(n_60923), .Z(n_60947));
	notech_inv i_13902(.A(n_60923), .Z(n_60945));
	notech_inv i_13899(.A(n_60923), .Z(n_60942));
	notech_inv i_13896(.A(n_60923), .Z(n_60940));
	notech_inv i_13894(.A(n_60923), .Z(n_60938));
	notech_inv i_13891(.A(n_60923), .Z(n_60935));
	notech_inv i_13888(.A(n_60923), .Z(n_60933));
	notech_inv i_13886(.A(n_60923), .Z(n_60931));
	notech_inv i_13883(.A(n_60923), .Z(n_60928));
	notech_inv i_13880(.A(n_60923), .Z(n_60926));
	notech_inv i_13878(.A(n_60923), .Z(n_60924));
	notech_inv i_13877(.A(n_2561), .Z(n_60923));
	notech_inv i_13869(.A(n_60914), .Z(n_60915));
	notech_inv i_13868(.A(instrc[121]), .Z(n_60914));
	notech_inv i_13864(.A(n_60898), .Z(n_60910));
	notech_inv i_13863(.A(n_60898), .Z(n_60909));
	notech_inv i_13858(.A(n_60898), .Z(n_60904));
	notech_inv i_13852(.A(n_60898), .Z(n_60899));
	notech_inv i_13851(.A(n_2546), .Z(n_60898));
	notech_inv i_13847(.A(n_60882), .Z(n_60894));
	notech_inv i_13846(.A(n_60882), .Z(n_60893));
	notech_inv i_13840(.A(n_60882), .Z(n_60888));
	notech_inv i_13835(.A(n_60882), .Z(n_60883));
	notech_inv i_13834(.A(n_32467), .Z(n_60882));
	notech_inv i_13826(.A(n_60873), .Z(n_60874));
	notech_inv i_13824(.A(n_32747), .Z(n_60873));
	notech_inv i_13820(.A(n_60862), .Z(n_60868));
	notech_inv i_13814(.A(n_60862), .Z(n_60863));
	notech_inv i_13813(.A(n_32448), .Z(n_60862));
	notech_inv i_13805(.A(n_60853), .Z(n_60854));
	notech_inv i_13804(.A(n_32326), .Z(n_60853));
	notech_inv i_13796(.A(n_60840), .Z(n_60845));
	notech_inv i_13791(.A(n_60840), .Z(n_60841));
	notech_inv i_13790(.A(n_27104), .Z(n_60840));
	notech_inv i_13780(.A(n_60829), .Z(n_60830));
	notech_inv i_13779(.A(n_328290780), .Z(n_60829));
	notech_inv i_13730(.A(n_60764), .Z(n_60774));
	notech_inv i_13728(.A(n_60764), .Z(n_60773));
	notech_inv i_13724(.A(n_60764), .Z(n_60769));
	notech_inv i_13719(.A(n_60764), .Z(n_60765));
	notech_inv i_13718(.A(ipg_fault), .Z(n_60764));
	notech_inv i_13603(.A(n_60535), .Z(n_60550));
	notech_inv i_13601(.A(n_60535), .Z(n_60548));
	notech_inv i_13594(.A(n_60535), .Z(n_60542));
	notech_inv i_13588(.A(n_60535), .Z(n_60537));
	notech_inv i_13587(.A(n_60535), .Z(cr0[0]));
	notech_inv i_13586(.A(\nbus_14526[0] ), .Z(n_60535));
	notech_inv i_13450(.A(n_60386), .Z(n_60387));
	notech_inv i_13449(.A(n_60123), .Z(n_60386));
	notech_inv i_13441(.A(n_60377), .Z(n_60378));
	notech_inv i_13440(.A(n_2885), .Z(n_60377));
	notech_inv i_13436(.A(n_19101), .Z(n_60373));
	notech_inv i_13435(.A(n_19101), .Z(n_60372));
	notech_inv i_13429(.A(n_19101), .Z(n_60367));
	notech_inv i_13420(.A(n_60357), .Z(n_60358));
	notech_inv i_13419(.A(n_60356), .Z(n_60357));
	notech_inv i_13418(.A(n_60291), .Z(n_60356));
	notech_inv i_13410(.A(n_60348), .Z(n_60349));
	notech_inv i_13409(.A(n_60347), .Z(n_60348));
	notech_inv i_13408(.A(n_60291), .Z(n_60347));
	notech_inv i_13400(.A(n_60339), .Z(n_60340));
	notech_inv i_13399(.A(n_60338), .Z(n_60339));
	notech_inv i_13397(.A(n_60291), .Z(n_60338));
	notech_inv i_13389(.A(n_60330), .Z(n_60331));
	notech_inv i_13388(.A(n_60329), .Z(n_60330));
	notech_inv i_13387(.A(n_60291), .Z(n_60329));
	notech_inv i_13378(.A(n_60320), .Z(n_60321));
	notech_inv i_13377(.A(n_60319), .Z(n_60320));
	notech_inv i_13376(.A(n_60291), .Z(n_60319));
	notech_inv i_13375(.A(n_60291), .Z(n_60318));
	notech_inv i_13372(.A(n_60291), .Z(n_60316));
	notech_inv i_13368(.A(n_60291), .Z(n_60312));
	notech_inv i_13357(.A(n_60302), .Z(n_60303));
	notech_inv i_13356(.A(n_60292), .Z(n_60302));
	notech_inv i_13352(.A(n_60302), .Z(n_60298));
	notech_inv i_13347(.A(n_60302), .Z(n_60294));
	notech_inv i_13345(.A(n_60291), .Z(n_60292));
	notech_inv i_13344(.A(n_1914992224), .Z(n_60291));
	notech_inv i_13336(.A(n_60282), .Z(n_60283));
	notech_inv i_13335(.A(n_19086), .Z(n_60282));
	notech_inv i_13327(.A(n_60273), .Z(n_60274));
	notech_inv i_13325(.A(n_2875), .Z(n_60273));
	notech_inv i_13321(.A(n_60318), .Z(n_60268));
	notech_inv i_13315(.A(n_60318), .Z(n_60263));
	notech_inv i_13308(.A(n_60318), .Z(n_60257));
	notech_inv i_13302(.A(n_60318), .Z(n_60252));
	notech_inv i_13295(.A(n_60318), .Z(n_60246));
	notech_inv i_13289(.A(n_60318), .Z(n_60241));
	notech_inv i_13281(.A(n_60318), .Z(n_60234));
	notech_inv i_13275(.A(n_60318), .Z(n_60229));
	notech_inv i_13268(.A(n_60318), .Z(n_60223));
	notech_inv i_13263(.A(n_60318), .Z(n_60218));
	notech_inv i_13256(.A(n_60318), .Z(n_60212));
	notech_inv i_13250(.A(n_60318), .Z(n_60207));
	notech_inv i_13236(.A(n_60194), .Z(n_60195));
	notech_inv i_13235(.A(n_60193), .Z(n_60194));
	notech_inv i_13234(.A(n_60318), .Z(n_60193));
	notech_inv i_13224(.A(n_60183), .Z(n_60184));
	notech_inv i_13223(.A(n_60171), .Z(n_60183));
	notech_inv i_13217(.A(n_60183), .Z(n_60178));
	notech_inv i_13211(.A(n_60183), .Z(n_60173));
	notech_inv i_13209(.A(n_60318), .Z(n_60171));
	notech_inv i_13206(.A(n_60110), .Z(n_60167));
	notech_inv i_13204(.A(n_60110), .Z(n_60166));
	notech_inv i_13200(.A(n_60110), .Z(n_60162));
	notech_inv i_13195(.A(n_60110), .Z(n_60158));
	notech_inv i_13194(.A(n_60110), .Z(n_60157));
	notech_inv i_13190(.A(n_60110), .Z(n_60153));
	notech_inv i_13185(.A(n_60110), .Z(n_60149));
	notech_inv i_13184(.A(n_60110), .Z(n_60148));
	notech_inv i_13179(.A(n_60110), .Z(n_60144));
	notech_inv i_13174(.A(n_60110), .Z(n_60139));
	notech_inv i_13172(.A(n_60110), .Z(n_60138));
	notech_inv i_13168(.A(n_60110), .Z(n_60133));
	notech_inv i_13163(.A(n_60110), .Z(n_60128));
	notech_inv i_13162(.A(n_60110), .Z(n_60127));
	notech_inv i_13158(.A(n_60110), .Z(n_60122));
	notech_inv i_13152(.A(n_60110), .Z(n_60117));
	notech_inv i_13147(.A(n_60110), .Z(n_60113));
	notech_inv i_13144(.A(n_29654), .Z(n_60110));
	notech_inv i_13136(.A(n_60101), .Z(n_60102));
	notech_inv i_13135(.A(opa[15]), .Z(n_60101));
	notech_inv i_13127(.A(n_60090), .Z(n_60091));
	notech_inv i_13126(.A(opa[7]), .Z(n_60090));
	notech_inv i_13118(.A(n_60081), .Z(n_60082));
	notech_inv i_13116(.A(opa[6]), .Z(n_60081));
	notech_inv i_13108(.A(n_60071), .Z(n_60072));
	notech_inv i_13107(.A(opa[0]), .Z(n_60071));
	notech_inv i_12819(.A(n_59750), .Z(n_59766));
	notech_inv i_12817(.A(n_59750), .Z(n_59764));
	notech_inv i_12816(.A(n_59750), .Z(n_59763));
	notech_inv i_12810(.A(n_59750), .Z(n_59758));
	notech_inv i_12802(.A(n_59750), .Z(n_59751));
	notech_inv i_12801(.A(n_58215), .Z(n_59750));
	notech_inv i_12793(.A(n_59741), .Z(n_59742));
	notech_inv i_12792(.A(\nbus_11307[0] ), .Z(n_59741));
	notech_inv i_12786(.A(n_59734), .Z(n_59735));
	notech_inv i_12785(.A(opc[0]), .Z(n_59734));
	notech_inv i_12777(.A(n_59725), .Z(n_59726));
	notech_inv i_12776(.A(\nbus_11365[31] ), .Z(n_59725));
	notech_inv i_12768(.A(n_59716), .Z(n_59717));
	notech_inv i_12767(.A(nbus_11295[0]), .Z(n_59716));
	notech_inv i_12759(.A(n_59707), .Z(n_59708));
	notech_inv i_12758(.A(n_26602), .Z(n_59707));
	notech_inv i_12531(.A(n_59477), .Z(n_59478));
	notech_inv i_12529(.A(n_25617), .Z(n_59477));
	notech_inv i_12521(.A(n_59468), .Z(n_59469));
	notech_inv i_12520(.A(n_24989), .Z(n_59468));
	notech_inv i_12512(.A(n_59459), .Z(n_59460));
	notech_inv i_12511(.A(n_27917), .Z(n_59459));
	notech_inv i_12503(.A(n_59450), .Z(n_59451));
	notech_inv i_12502(.A(n_27907), .Z(n_59450));
	notech_inv i_12497(.A(n_59439), .Z(n_59445));
	notech_inv i_12493(.A(n_59439), .Z(n_59441));
	notech_inv i_12492(.A(n_59439), .Z(n_59440));
	notech_inv i_12491(.A(n_32763), .Z(n_59439));
	notech_inv i_12487(.A(n_59441), .Z(n_59435));
	notech_inv i_12486(.A(n_59441), .Z(n_59434));
	notech_inv i_12480(.A(n_59441), .Z(n_59429));
	notech_inv i_12475(.A(n_59441), .Z(n_59424));
	notech_inv i_12470(.A(n_59412), .Z(n_59419));
	notech_inv i_12469(.A(n_59412), .Z(n_59418));
	notech_inv i_12463(.A(n_59412), .Z(n_59413));
	notech_inv i_12462(.A(n_32650), .Z(n_59412));
	notech_inv i_12459(.A(n_59401), .Z(n_59408));
	notech_inv i_12457(.A(n_59401), .Z(n_59407));
	notech_inv i_12452(.A(n_59401), .Z(n_59402));
	notech_inv i_12451(.A(instrc[113]), .Z(n_59401));
	notech_inv i_12448(.A(n_59392), .Z(n_59398));
	notech_inv i_12447(.A(n_59392), .Z(n_59397));
	notech_inv i_12443(.A(n_59392), .Z(n_59393));
	notech_inv i_12441(.A(instrc[114]), .Z(n_59392));
	notech_inv i_12437(.A(n_59381), .Z(n_59387));
	notech_inv i_12431(.A(n_59381), .Z(n_59382));
	notech_inv i_12430(.A(instrc[112]), .Z(n_59381));
	notech_inv i_12422(.A(n_59372), .Z(n_59373));
	notech_inv i_12421(.A(instrc[115]), .Z(n_59372));
	notech_inv i_12413(.A(n_59363), .Z(n_59364));
	notech_inv i_12412(.A(n_29178), .Z(n_59363));
	notech_inv i_12404(.A(n_59354), .Z(n_59355));
	notech_inv i_12403(.A(n_2479), .Z(n_59354));
	notech_inv i_12398(.A(n_32612), .Z(n_59349));
	notech_inv i_12392(.A(n_32612), .Z(n_59344));
	notech_inv i_12383(.A(n_59334), .Z(n_59335));
	notech_inv i_12382(.A(n_27065), .Z(n_59334));
	notech_inv i_12374(.A(n_59321), .Z(n_59326));
	notech_inv i_12369(.A(n_59321), .Z(n_59322));
	notech_inv i_12368(.A(n_32270), .Z(n_59321));
	notech_inv i_12336(.A(n_59285), .Z(n_59286));
	notech_inv i_12335(.A(n_246991940), .Z(n_59285));
	notech_inv i_12324(.A(n_59274), .Z(n_59275));
	notech_inv i_12323(.A(n_246891941), .Z(n_59274));
	notech_inv i_12308(.A(n_59258), .Z(n_59259));
	notech_inv i_12307(.A(n_27984), .Z(n_59258));
	notech_inv i_12290(.A(n_59240), .Z(n_59241));
	notech_inv i_12287(.A(n_27983), .Z(n_59240));
	notech_inv i_12270(.A(n_59222), .Z(n_59223));
	notech_inv i_12269(.A(n_27985), .Z(n_59222));
	notech_inv i_12261(.A(n_27986), .Z(n_59214));
	notech_inv i_12251(.A(n_59204), .Z(n_59205));
	notech_inv i_12250(.A(n_27987), .Z(n_59204));
	notech_inv i_12233(.A(n_59186), .Z(n_59187));
	notech_inv i_12232(.A(n_27981), .Z(n_59186));
	notech_inv i_12221(.A(n_59175), .Z(n_59176));
	notech_inv i_12220(.A(n_330563522), .Z(n_59175));
	notech_inv i_12212(.A(n_59166), .Z(n_59167));
	notech_inv i_12211(.A(n_1887), .Z(n_59166));
	notech_inv i_12202(.A(n_59157), .Z(n_59158));
	notech_inv i_12201(.A(n_58662), .Z(n_59157));
	notech_inv i_12197(.A(n_59141), .Z(n_59153));
	notech_inv i_12196(.A(n_59141), .Z(n_59152));
	notech_inv i_12191(.A(n_59141), .Z(n_59147));
	notech_inv i_12185(.A(n_59141), .Z(n_59142));
	notech_inv i_12184(.A(n_315491669), .Z(n_59141));
	notech_inv i_12176(.A(n_59132), .Z(n_59133));
	notech_inv i_12175(.A(n_315391670), .Z(n_59132));
	notech_inv i_12167(.A(n_59123), .Z(n_59124));
	notech_inv i_12165(.A(n_151028787), .Z(n_59123));
	notech_inv i_12157(.A(n_59114), .Z(n_59115));
	notech_inv i_12156(.A(n_318391640), .Z(n_59114));
	notech_inv i_12148(.A(n_59105), .Z(n_59106));
	notech_inv i_12147(.A(n_318291641), .Z(n_59105));
	notech_inv i_12143(.A(n_59094), .Z(n_59100));
	notech_inv i_12137(.A(n_59094), .Z(n_59095));
	notech_inv i_12136(.A(n_32269), .Z(n_59094));
	notech_inv i_11204(.A(n_58096), .Z(n_58101));
	notech_inv i_11202(.A(calc_sz[1]), .Z(n_58096));
	notech_inv i_11194(.A(n_58083), .Z(n_58086));
	notech_inv i_11193(.A(n_25625), .Z(n_58083));
	notech_inv i_11185(.A(n_58070), .Z(n_58072));
	notech_inv i_11184(.A(n_2941), .Z(n_58070));
	notech_inv i_11176(.A(n_58061), .Z(n_58062));
	notech_inv i_11175(.A(n_2938), .Z(n_58061));
	notech_inv i_11167(.A(n_58045), .Z(n_58046));
	notech_inv i_11166(.A(n_25385), .Z(n_58045));
	notech_inv i_11158(.A(n_58032), .Z(n_58033));
	notech_inv i_11157(.A(n_26965), .Z(n_58032));
	notech_inv i_11149(.A(n_58019), .Z(n_58024));
	notech_inv i_11144(.A(n_58019), .Z(n_58020));
	notech_inv i_11143(.A(n_27089), .Z(n_58019));
	notech_inv i_11138(.A(n_32316), .Z(n_58014));
	notech_inv i_11133(.A(n_32316), .Z(n_58009));
	notech_inv i_11124(.A(n_57991), .Z(n_57992));
	notech_inv i_11122(.A(n_32341), .Z(n_57991));
	notech_inv i_11118(.A(n_57992), .Z(n_57985));
	notech_inv i_11112(.A(n_57992), .Z(n_57976));
	notech_inv i_11103(.A(n_57965), .Z(n_57967));
	notech_inv i_11102(.A(n_27896), .Z(n_57965));
	notech_inv i_11094(.A(n_57956), .Z(n_57957));
	notech_inv i_11093(.A(\nbus_11307[7] ), .Z(n_57956));
	notech_inv i_11085(.A(n_57946), .Z(n_57948));
	notech_inv i_11084(.A(n_3901), .Z(n_57946));
	notech_inv i_11076(.A(n_57932), .Z(n_57933));
	notech_inv i_11074(.A(n_2949), .Z(n_57932));
	notech_inv i_11066(.A(n_57919), .Z(n_57920));
	notech_inv i_11065(.A(n_23029), .Z(n_57919));
	notech_inv i_11057(.A(n_57908), .Z(n_57909));
	notech_inv i_11056(.A(nbus_11295[3]), .Z(n_57908));
	notech_inv i_11048(.A(n_57898), .Z(n_57899));
	notech_inv i_11047(.A(n_27877), .Z(n_57898));
	notech_inv i_11039(.A(n_57880), .Z(n_57881));
	notech_inv i_11038(.A(nbus_11295[27]), .Z(n_57880));
	notech_inv i_11028(.A(n_57858), .Z(n_57859));
	notech_inv i_11026(.A(n_23019), .Z(n_57858));
	notech_inv i_11016(.A(n_57847), .Z(n_57848));
	notech_inv i_11015(.A(n_23003), .Z(n_57847));
	notech_inv i_11007(.A(n_57836), .Z(n_57837));
	notech_inv i_11006(.A(\nbus_11358[31] ), .Z(n_57836));
	notech_inv i_10998(.A(n_57826), .Z(n_57828));
	notech_inv i_10997(.A(\nbus_11365[30] ), .Z(n_57826));
	notech_inv i_10989(.A(n_57814), .Z(n_57815));
	notech_inv i_10988(.A(\nbus_11365[29] ), .Z(n_57814));
	notech_inv i_10980(.A(n_57801), .Z(n_57802));
	notech_inv i_10978(.A(\nbus_11365[28] ), .Z(n_57801));
	notech_inv i_10970(.A(n_57791), .Z(n_57792));
	notech_inv i_10969(.A(\nbus_11365[27] ), .Z(n_57791));
	notech_inv i_10961(.A(n_57782), .Z(n_57783));
	notech_inv i_10960(.A(\nbus_11365[26] ), .Z(n_57782));
	notech_inv i_10952(.A(n_57770), .Z(n_57771));
	notech_inv i_10951(.A(\nbus_11365[25] ), .Z(n_57770));
	notech_inv i_10943(.A(n_57760), .Z(n_57761));
	notech_inv i_10942(.A(\nbus_11365[24] ), .Z(n_57760));
	notech_inv i_10934(.A(n_57750), .Z(n_57751));
	notech_inv i_10933(.A(\nbus_11365[23] ), .Z(n_57750));
	notech_inv i_10925(.A(n_57741), .Z(n_57742));
	notech_inv i_10924(.A(\nbus_11365[22] ), .Z(n_57741));
	notech_inv i_10916(.A(n_57732), .Z(n_57733));
	notech_inv i_10914(.A(\nbus_11365[21] ), .Z(n_57732));
	notech_inv i_10906(.A(n_57719), .Z(n_57720));
	notech_inv i_10905(.A(\nbus_11365[20] ), .Z(n_57719));
	notech_inv i_10897(.A(n_57706), .Z(n_57707));
	notech_inv i_10896(.A(\nbus_11365[19] ), .Z(n_57706));
	notech_inv i_10888(.A(n_57697), .Z(n_57698));
	notech_inv i_10887(.A(\nbus_11365[18] ), .Z(n_57697));
	notech_inv i_10879(.A(n_57688), .Z(n_57689));
	notech_inv i_10878(.A(\nbus_11365[17] ), .Z(n_57688));
	notech_inv i_10870(.A(n_57679), .Z(n_57680));
	notech_inv i_10869(.A(\nbus_11365[16] ), .Z(n_57679));
	notech_inv i_10861(.A(n_57670), .Z(n_57671));
	notech_inv i_10860(.A(\nbus_11307[15] ), .Z(n_57670));
	notech_inv i_10852(.A(n_57661), .Z(n_57662));
	notech_inv i_10850(.A(\nbus_11307[14] ), .Z(n_57661));
	notech_inv i_10842(.A(n_57652), .Z(n_57653));
	notech_inv i_10841(.A(\nbus_11307[13] ), .Z(n_57652));
	notech_inv i_10833(.A(n_57643), .Z(n_57644));
	notech_inv i_10832(.A(\nbus_11307[12] ), .Z(n_57643));
	notech_inv i_10824(.A(n_57634), .Z(n_57635));
	notech_inv i_10823(.A(\nbus_11307[11] ), .Z(n_57634));
	notech_inv i_10815(.A(n_57624), .Z(n_57625));
	notech_inv i_10814(.A(\nbus_11307[10] ), .Z(n_57624));
	notech_inv i_10806(.A(n_57612), .Z(n_57613));
	notech_inv i_10805(.A(\nbus_11307[9] ), .Z(n_57612));
	notech_inv i_10797(.A(n_57603), .Z(n_57604));
	notech_inv i_10796(.A(\nbus_11307[8] ), .Z(n_57603));
	notech_inv i_10788(.A(n_57591), .Z(n_57592));
	notech_inv i_10786(.A(\nbus_11307[6] ), .Z(n_57591));
	notech_inv i_10778(.A(n_57582), .Z(n_57583));
	notech_inv i_10777(.A(\nbus_11307[5] ), .Z(n_57582));
	notech_inv i_10769(.A(n_57572), .Z(n_57574));
	notech_inv i_10768(.A(\nbus_11307[4] ), .Z(n_57572));
	notech_inv i_10760(.A(n_57562), .Z(n_57563));
	notech_inv i_10759(.A(\nbus_11307[3] ), .Z(n_57562));
	notech_inv i_10754(.A(opa[2]), .Z(n_57557));
	notech_inv i_10749(.A(opa[2]), .Z(n_57552));
	notech_inv i_10740(.A(n_57541), .Z(n_57542));
	notech_inv i_10738(.A(\nbus_11307[1] ), .Z(n_57541));
	notech_inv i_10736(.A(n_57532), .Z(n_57538));
	notech_inv i_10735(.A(n_57532), .Z(n_57537));
	notech_inv i_10730(.A(n_57532), .Z(n_57533));
	notech_inv i_10729(.A(n_23947), .Z(n_57532));
	notech_inv i_10721(.A(n_57523), .Z(n_57524));
	notech_inv i_10720(.A(n_23059), .Z(n_57523));
	notech_inv i_10710(.A(n_57511), .Z(n_57512));
	notech_inv i_10709(.A(n_1877), .Z(n_57511));
	notech_inv i_10699(.A(n_57497), .Z(n_57498));
	notech_inv i_10697(.A(n_1876), .Z(n_57497));
	notech_inv i_10586(.A(n_57374), .Z(n_57379));
	notech_inv i_10581(.A(n_57374), .Z(n_57375));
	notech_inv i_10580(.A(n_227976218), .Z(n_57374));
	notech_inv i_10576(.A(n_57360), .Z(n_57369));
	notech_inv i_10575(.A(n_57360), .Z(n_57368));
	notech_inv i_10570(.A(n_57360), .Z(n_57363));
	notech_inv i_10569(.A(n_57360), .Z(n_57362));
	notech_inv i_10568(.A(n_57360), .Z(n_57361));
	notech_inv i_10567(.A(instrc[106]), .Z(n_57360));
	notech_inv i_10520(.A(n_57176), .Z(n_57177));
	notech_inv i_10519(.A(n_296376902), .Z(n_57176));
	notech_inv i_10508(.A(n_57164), .Z(n_57165));
	notech_inv i_10507(.A(n_23052), .Z(n_57164));
	notech_inv i_10499(.A(n_57153), .Z(n_57155));
	notech_inv i_10498(.A(n_23049), .Z(n_57153));
	notech_inv i_10488(.A(n_57142), .Z(n_57143));
	notech_inv i_10487(.A(n_23045), .Z(n_57142));
	notech_inv i_10479(.A(n_57131), .Z(n_57132));
	notech_inv i_10477(.A(n_303747815), .Z(n_57131));
	notech_inv i_10467(.A(n_57120), .Z(n_57121));
	notech_inv i_10466(.A(n_18756873), .Z(n_57120));
	notech_inv i_10440(.A(n_57091), .Z(n_57092));
	notech_inv i_10439(.A(n_3918), .Z(n_57091));
	notech_inv i_10436(.A(n_57077), .Z(n_57088));
	notech_inv i_10435(.A(n_57077), .Z(n_57087));
	notech_inv i_10431(.A(n_57077), .Z(n_57082));
	notech_inv i_10426(.A(n_57077), .Z(n_57078));
	notech_inv i_10425(.A(instrc[117]), .Z(n_57077));
	notech_inv i_10417(.A(n_57063), .Z(n_57068));
	notech_inv i_10412(.A(n_57063), .Z(n_57064));
	notech_inv i_10411(.A(instrc[116]), .Z(n_57063));
	notech_inv i_10403(.A(n_57050), .Z(n_57055));
	notech_inv i_10399(.A(n_57050), .Z(n_57051));
	notech_inv i_10397(.A(n_29652), .Z(n_57050));
	notech_inv i_10389(.A(n_57041), .Z(n_57042));
	notech_inv i_10388(.A(instrc[119]), .Z(n_57041));
	notech_inv i_10378(.A(n_57032), .Z(n_57033));
	notech_inv i_10377(.A(n_29653), .Z(n_57032));
	notech_inv i_10373(.A(n_57019), .Z(n_57026));
	notech_inv i_10367(.A(n_57019), .Z(n_57020));
	notech_inv i_10366(.A(instrc[118]), .Z(n_57019));
	notech_inv i_10358(.A(n_57010), .Z(n_57011));
	notech_inv i_10357(.A(n_29658), .Z(n_57010));
	notech_inv i_10349(.A(n_57001), .Z(n_57002));
	notech_inv i_10347(.A(n_27090), .Z(n_57001));
	notech_inv i_10339(.A(n_56991), .Z(n_56992));
	notech_inv i_10338(.A(n_3921), .Z(n_56991));
	notech_inv i_10330(.A(n_56978), .Z(n_56983));
	notech_inv i_10326(.A(n_56978), .Z(n_56979));
	notech_inv i_10325(.A(n_26610), .Z(n_56978));
	notech_inv i_10317(.A(n_56969), .Z(n_56970));
	notech_inv i_10315(.A(n_246691943), .Z(n_56969));
	notech_inv i_10305(.A(n_56958), .Z(n_56959));
	notech_inv i_10304(.A(n_32382), .Z(n_56958));
	notech_inv i_10296(.A(n_56939), .Z(n_56950));
	notech_inv i_10293(.A(n_32380), .Z(n_56946));
	notech_inv i_10290(.A(n_32380), .Z(n_56944));
	notech_inv i_10287(.A(n_32380), .Z(n_56941));
	notech_inv i_10285(.A(n_32380), .Z(n_56939));
	notech_inv i_10280(.A(n_32380), .Z(n_56935));
	notech_inv i_10270(.A(n_56924), .Z(n_56925));
	notech_inv i_10269(.A(n_319191632), .Z(n_56924));
	notech_inv i_10266(.A(n_32299), .Z(n_56921));
	notech_inv i_10264(.A(n_32299), .Z(n_56919));
	notech_inv i_10261(.A(n_32299), .Z(n_56916));
	notech_inv i_10258(.A(n_32299), .Z(n_56914));
	notech_inv i_10254(.A(n_32325), .Z(n_56909));
	notech_inv i_10253(.A(n_32325), .Z(n_56908));
	notech_inv i_10247(.A(n_32325), .Z(n_56903));
	notech_inv i_10238(.A(n_56893), .Z(n_56894));
	notech_inv i_10237(.A(n_3914), .Z(n_56893));
	notech_inv i_10232(.A(n_56882), .Z(n_56888));
	notech_inv i_10226(.A(n_56882), .Z(n_56883));
	notech_inv i_10225(.A(n_3920), .Z(n_56882));
	notech_inv i_10215(.A(n_56871), .Z(n_56872));
	notech_inv i_10214(.A(\nbus_11335[0] ), .Z(n_56871));
	notech_inv i_10206(.A(n_56862), .Z(n_56863));
	notech_inv i_10205(.A(n_30854), .Z(n_56862));
	notech_inv i_10202(.A(n_56853), .Z(n_56859));
	notech_inv i_10201(.A(n_56853), .Z(n_56858));
	notech_inv i_10197(.A(n_56853), .Z(n_56854));
	notech_inv i_10195(.A(n_32376), .Z(n_56853));
	notech_inv i_10191(.A(n_56842), .Z(n_56848));
	notech_inv i_10185(.A(n_56842), .Z(n_56843));
	notech_inv i_10184(.A(n_308691737), .Z(n_56842));
	notech_inv i_10182(.A(n_56821), .Z(n_56839));
	notech_inv i_10179(.A(n_56821), .Z(n_56837));
	notech_inv i_10176(.A(n_56821), .Z(n_56834));
	notech_inv i_10174(.A(n_56821), .Z(n_56832));
	notech_inv i_10170(.A(n_56821), .Z(n_56829));
	notech_inv i_10168(.A(n_56821), .Z(n_56827));
	notech_inv i_10165(.A(n_56821), .Z(n_56824));
	notech_inv i_10162(.A(n_56821), .Z(n_56822));
	notech_inv i_10161(.A(n_32372), .Z(n_56821));
	notech_inv i_10153(.A(n_56812), .Z(n_56813));
	notech_inv i_10152(.A(n_32348), .Z(n_56812));
	notech_inv i_10144(.A(n_56802), .Z(n_56803));
	notech_inv i_10143(.A(n_58477), .Z(n_56802));
	notech_inv i_10041(.A(n_56683), .Z(n_56689));
	notech_inv i_10040(.A(n_56683), .Z(n_56688));
	notech_inv i_10035(.A(n_56683), .Z(n_56684));
	notech_inv i_10034(.A(n_32371), .Z(n_56683));
	notech_inv i_10026(.A(n_56674), .Z(n_56675));
	notech_inv i_10025(.A(n_32356), .Z(n_56674));
	notech_inv i_10017(.A(n_56661), .Z(n_56666));
	notech_inv i_10013(.A(n_56661), .Z(n_56662));
	notech_inv i_10011(.A(n_26924), .Z(n_56661));
	notech_inv i_10003(.A(n_56648), .Z(n_56653));
	notech_inv i_9999(.A(n_56648), .Z(n_56649));
	notech_inv i_9998(.A(n_26922), .Z(n_56648));
	notech_inv i_9990(.A(n_56635), .Z(n_56640));
	notech_inv i_9985(.A(n_56635), .Z(n_56636));
	notech_inv i_9984(.A(n_26969), .Z(n_56635));
	notech_inv i_9982(.A(n_32287), .Z(n_56632));
	notech_inv i_9979(.A(n_32287), .Z(n_56630));
	notech_inv i_9976(.A(n_32287), .Z(n_56627));
	notech_inv i_9974(.A(n_32287), .Z(n_56625));
	notech_inv i_9968(.A(n_32286), .Z(n_56619));
	notech_inv i_9962(.A(n_32286), .Z(n_56614));
	notech_inv i_9953(.A(n_56600), .Z(n_56605));
	notech_inv i_9949(.A(n_56600), .Z(n_56601));
	notech_inv i_9947(.A(n_26928), .Z(n_56600));
	notech_inv i_9939(.A(n_56591), .Z(n_56592));
	notech_inv i_9938(.A(n_26651), .Z(n_56591));
	notech_inv i_9930(.A(n_56578), .Z(n_56583));
	notech_inv i_9926(.A(n_56578), .Z(n_56579));
	notech_inv i_9925(.A(n_26925), .Z(n_56578));
	notech_inv i_9917(.A(n_56565), .Z(n_56570));
	notech_inv i_9912(.A(n_56565), .Z(n_56566));
	notech_inv i_9911(.A(n_27036), .Z(n_56565));
	notech_inv i_9903(.A(n_56552), .Z(n_56557));
	notech_inv i_9898(.A(n_56552), .Z(n_56553));
	notech_inv i_9897(.A(n_26721), .Z(n_56552));
	notech_inv i_9894(.A(n_32279), .Z(n_56548));
	notech_inv i_9893(.A(n_32279), .Z(n_56547));
	notech_inv i_9887(.A(n_32279), .Z(n_56542));
	notech_inv i_9878(.A(n_56526), .Z(n_56532));
	notech_inv i_9873(.A(n_56526), .Z(n_56527));
	notech_inv i_9872(.A(n_26927), .Z(n_56526));
	notech_inv i_9864(.A(n_56511), .Z(n_56518));
	notech_inv i_9859(.A(n_56511), .Z(n_56513));
	notech_inv i_9858(.A(n_26649), .Z(n_56511));
	notech_inv i_9848(.A(n_56497), .Z(n_56502));
	notech_inv i_9844(.A(n_56497), .Z(n_56498));
	notech_inv i_9843(.A(n_26920), .Z(n_56497));
	notech_inv i_9834(.A(n_56484), .Z(n_56489));
	notech_inv i_9829(.A(n_56484), .Z(n_56485));
	notech_inv i_9828(.A(n_26933), .Z(n_56484));
	notech_inv i_9820(.A(n_56474), .Z(n_56475));
	notech_inv i_9819(.A(\nbus_11358[24] ), .Z(n_56474));
	notech_inv i_9814(.A(n_32327), .Z(n_56468));
	notech_inv i_9808(.A(n_32327), .Z(n_56463));
	notech_inv i_9803(.A(n_32338), .Z(n_56457));
	notech_inv i_9797(.A(n_32338), .Z(n_56452));
	notech_inv i_9794(.A(n_32332), .Z(n_56448));
	notech_inv i_9792(.A(n_32332), .Z(n_56447));
	notech_inv i_9788(.A(n_32332), .Z(n_56443));
	notech_inv i_9782(.A(n_32331), .Z(n_56437));
	notech_inv i_9776(.A(n_32331), .Z(n_56432));
	notech_inv i_9773(.A(n_32322), .Z(n_56428));
	notech_inv i_9772(.A(n_32322), .Z(n_56427));
	notech_inv i_9767(.A(n_32322), .Z(n_56423));
	notech_inv i_9758(.A(n_56413), .Z(n_56414));
	notech_inv i_9757(.A(n_27094), .Z(n_56413));
	notech_inv i_9749(.A(n_56404), .Z(n_56405));
	notech_inv i_9748(.A(n_26950), .Z(n_56404));
	notech_inv i_9746(.A(n_32365), .Z(n_56401));
	notech_inv i_9744(.A(n_32365), .Z(n_56400));
	notech_inv i_9740(.A(n_32365), .Z(n_56396));
	notech_inv i_9735(.A(n_32334), .Z(n_56391));
	notech_inv i_9734(.A(n_32334), .Z(n_56390));
	notech_inv i_9728(.A(n_32334), .Z(n_56385));
	notech_inv i_9723(.A(n_32334), .Z(n_56380));
	notech_inv i_9714(.A(n_56366), .Z(n_56371));
	notech_inv i_9709(.A(n_56366), .Z(n_56367));
	notech_inv i_9708(.A(n_26664), .Z(n_56366));
	notech_inv i_9698(.A(n_56355), .Z(n_56356));
	notech_inv i_9696(.A(n_154331958), .Z(n_56355));
	notech_inv i_9688(.A(n_56346), .Z(n_56347));
	notech_inv i_9687(.A(\nbus_11358[23] ), .Z(n_56346));
	notech_inv i_9679(.A(n_56337), .Z(n_56338));
	notech_inv i_9678(.A(\nbus_11358[22] ), .Z(n_56337));
	notech_inv i_9670(.A(n_56328), .Z(n_56329));
	notech_inv i_9669(.A(\nbus_11358[21] ), .Z(n_56328));
	notech_inv i_9661(.A(n_56319), .Z(n_56320));
	notech_inv i_9660(.A(\nbus_11358[20] ), .Z(n_56319));
	notech_inv i_9652(.A(n_56310), .Z(n_56311));
	notech_inv i_9651(.A(\nbus_11358[19] ), .Z(n_56310));
	notech_inv i_9643(.A(n_56301), .Z(n_56302));
	notech_inv i_9642(.A(\nbus_11358[18] ), .Z(n_56301));
	notech_inv i_9634(.A(n_56292), .Z(n_56293));
	notech_inv i_9632(.A(\nbus_11358[17] ), .Z(n_56292));
	notech_inv i_9624(.A(n_56283), .Z(n_56284));
	notech_inv i_9623(.A(\nbus_11358[16] ), .Z(n_56283));
	notech_inv i_9615(.A(n_56274), .Z(n_56275));
	notech_inv i_9614(.A(\nbus_11358[15] ), .Z(n_56274));
	notech_inv i_9606(.A(n_56265), .Z(n_56266));
	notech_inv i_9605(.A(n_29754), .Z(n_56265));
	notech_inv i_9597(.A(n_56256), .Z(n_56257));
	notech_inv i_9596(.A(n_29680), .Z(n_56256));
	notech_inv i_9588(.A(n_56247), .Z(n_56248));
	notech_inv i_9587(.A(\nbus_11358[14] ), .Z(n_56247));
	notech_inv i_9579(.A(n_56238), .Z(n_56239));
	notech_inv i_9578(.A(n_29592), .Z(n_56238));
	notech_inv i_9570(.A(n_56229), .Z(n_56230));
	notech_inv i_9568(.A(\nbus_11358[13] ), .Z(n_56229));
	notech_inv i_9560(.A(n_56220), .Z(n_56221));
	notech_inv i_9559(.A(\nbus_11358[12] ), .Z(n_56220));
	notech_inv i_9549(.A(n_56209), .Z(n_56210));
	notech_inv i_9548(.A(n_3906), .Z(n_56209));
	notech_inv i_9544(.A(n_56198), .Z(n_56205));
	notech_inv i_9543(.A(n_56198), .Z(n_56204));
	notech_inv i_9537(.A(n_56198), .Z(n_56199));
	notech_inv i_9535(.A(n_81541430), .Z(n_56198));
	notech_inv i_9527(.A(n_56189), .Z(n_56190));
	notech_inv i_9526(.A(n_29596), .Z(n_56189));
	notech_inv i_9518(.A(n_56180), .Z(n_56181));
	notech_inv i_9517(.A(\nbus_11358[11] ), .Z(n_56180));
	notech_inv i_9509(.A(n_56171), .Z(n_56172));
	notech_inv i_9508(.A(\eflags[10] ), .Z(n_56171));
	notech_inv i_9500(.A(n_56162), .Z(n_56163));
	notech_inv i_9499(.A(n_29601), .Z(n_56162));
	notech_inv i_9491(.A(n_56153), .Z(n_56154));
	notech_inv i_9490(.A(\nbus_11358[10] ), .Z(n_56153));
	notech_inv i_9482(.A(n_56144), .Z(n_56145));
	notech_inv i_9481(.A(n_29684), .Z(n_56144));
	notech_inv i_9473(.A(n_56135), .Z(n_56136));
	notech_inv i_9471(.A(\nbus_11358[9] ), .Z(n_56135));
	notech_inv i_9463(.A(n_56126), .Z(n_56127));
	notech_inv i_9462(.A(n_29743), .Z(n_56126));
	notech_inv i_9454(.A(n_56117), .Z(n_56118));
	notech_inv i_9453(.A(\nbus_11358[8] ), .Z(n_56117));
	notech_inv i_9445(.A(n_56108), .Z(n_56109));
	notech_inv i_9444(.A(\nbus_11358[7] ), .Z(n_56108));
	notech_inv i_9436(.A(n_56099), .Z(n_56100));
	notech_inv i_9435(.A(n_27990), .Z(n_56099));
	notech_inv i_9427(.A(n_56090), .Z(n_56091));
	notech_inv i_9426(.A(n_309191732), .Z(n_56090));
	notech_inv i_9418(.A(n_56081), .Z(n_56082));
	notech_inv i_9417(.A(\nbus_11358[6] ), .Z(n_56081));
	notech_inv i_9409(.A(n_56072), .Z(n_56073));
	notech_inv i_9407(.A(\nbus_11358[5] ), .Z(n_56072));
	notech_inv i_9399(.A(n_56063), .Z(n_56064));
	notech_inv i_9398(.A(\nbus_11358[4] ), .Z(n_56063));
	notech_inv i_9390(.A(n_56054), .Z(n_56055));
	notech_inv i_9389(.A(n_29725), .Z(n_56054));
	notech_inv i_9381(.A(n_56045), .Z(n_56046));
	notech_inv i_9380(.A(n_60025), .Z(n_56045));
	notech_inv i_9371(.A(n_56036), .Z(n_56037));
	notech_inv i_9370(.A(n_29742), .Z(n_56036));
	notech_inv i_9362(.A(n_56027), .Z(n_56028));
	notech_inv i_9361(.A(\nbus_11358[0] ), .Z(n_56027));
	notech_inv i_9353(.A(n_56018), .Z(n_56019));
	notech_inv i_9352(.A(n_29678), .Z(n_56018));
	notech_inv i_9344(.A(n_56009), .Z(n_56010));
	notech_inv i_9342(.A(\nbus_11358[1] ), .Z(n_56009));
	notech_inv i_9340(.A(n_56000), .Z(n_56006));
	notech_inv i_9339(.A(n_56000), .Z(n_56005));
	notech_inv i_9334(.A(n_56000), .Z(n_56001));
	notech_inv i_9333(.A(gs[2]), .Z(n_56000));
	notech_inv i_9325(.A(n_55991), .Z(n_55992));
	notech_inv i_9324(.A(\nbus_11358[2] ), .Z(n_55991));
	notech_inv i_9316(.A(n_55982), .Z(n_55983));
	notech_inv i_9315(.A(\nbus_11358[3] ), .Z(n_55982));
	notech_inv i_9307(.A(n_55973), .Z(n_55974));
	notech_inv i_9306(.A(\nbus_11358[28] ), .Z(n_55973));
	notech_inv i_9298(.A(n_55964), .Z(n_55965));
	notech_inv i_9297(.A(\nbus_11358[25] ), .Z(n_55964));
	notech_inv i_9289(.A(n_55955), .Z(n_55956));
	notech_inv i_9288(.A(\nbus_11358[29] ), .Z(n_55955));
	notech_inv i_9280(.A(n_55946), .Z(n_55947));
	notech_inv i_9278(.A(\nbus_11358[26] ), .Z(n_55946));
	notech_inv i_9269(.A(n_55937), .Z(n_55938));
	notech_inv i_9268(.A(\nbus_11358[27] ), .Z(n_55937));
	notech_inv i_9260(.A(n_55928), .Z(n_55929));
	notech_inv i_9259(.A(\nbus_11358[30] ), .Z(n_55928));
	notech_inv i_9249(.A(n_55917), .Z(n_55918));
	notech_inv i_9248(.A(n_328090778), .Z(n_55917));
	notech_inv i_9240(.A(n_55908), .Z(n_55909));
	notech_inv i_9239(.A(n_54912649), .Z(n_55908));
	notech_inv i_9231(.A(n_55899), .Z(n_55900));
	notech_inv i_9229(.A(n_3892), .Z(n_55899));
	notech_inv i_9221(.A(n_55890), .Z(n_55891));
	notech_inv i_9220(.A(n_3882), .Z(n_55890));
	notech_inv i_9217(.A(n_55879), .Z(n_55886));
	notech_inv i_9216(.A(n_55879), .Z(n_55885));
	notech_inv i_9210(.A(n_55879), .Z(n_55880));
	notech_inv i_9209(.A(n_25329), .Z(n_55879));
	notech_inv i_9199(.A(n_55868), .Z(n_55869));
	notech_inv i_9197(.A(n_54212642), .Z(n_55868));
	notech_inv i_9189(.A(n_55859), .Z(n_55860));
	notech_inv i_9188(.A(n_54012640), .Z(n_55859));
	notech_inv i_9178(.A(n_55848), .Z(n_55849));
	notech_inv i_9176(.A(n_53612636), .Z(n_55848));
	notech_inv i_9166(.A(n_55837), .Z(n_55838));
	notech_inv i_9164(.A(n_53412634), .Z(n_55837));
	notech_inv i_9156(.A(n_55828), .Z(n_55829));
	notech_inv i_9155(.A(n_53512635), .Z(n_55828));
	notech_inv i_9147(.A(n_55819), .Z(n_55820));
	notech_inv i_9146(.A(n_27855), .Z(n_55819));
	notech_inv i_9136(.A(n_55808), .Z(n_55809));
	notech_inv i_9135(.A(n_388360286), .Z(n_55808));
	notech_inv i_9127(.A(n_55799), .Z(n_55800));
	notech_inv i_9126(.A(n_3887), .Z(n_55799));
	notech_inv i_9118(.A(n_55790), .Z(n_55791));
	notech_inv i_9116(.A(n_276383754), .Z(n_55790));
	notech_inv i_9108(.A(n_55781), .Z(n_55782));
	notech_inv i_9107(.A(n_3888), .Z(n_55781));
	notech_inv i_9099(.A(n_55772), .Z(n_55773));
	notech_inv i_9098(.A(n_23940), .Z(n_55772));
	notech_inv i_9090(.A(n_55763), .Z(n_55764));
	notech_inv i_9089(.A(n_23023), .Z(n_55763));
	notech_inv i_9063(.A(n_55734), .Z(n_55735));
	notech_inv i_9062(.A(n_27761), .Z(n_55734));
	notech_inv i_9054(.A(n_55725), .Z(n_55726));
	notech_inv i_9052(.A(n_308091743), .Z(n_55725));
	notech_inv i_8960(.A(n_55631), .Z(n_55632));
	notech_inv i_8959(.A(n_58768), .Z(n_55631));
	notech_inv i_8951(.A(n_55622), .Z(n_55623));
	notech_inv i_8950(.A(n_308084071), .Z(n_55622));
	notech_inv i_8939(.A(n_55611), .Z(n_55612));
	notech_inv i_8938(.A(n_307884069), .Z(n_55611));
	notech_inv i_8920(.A(n_55591), .Z(n_55592));
	notech_inv i_8919(.A(n_57367), .Z(n_55591));
	notech_inv i_8909(.A(n_55580), .Z(n_55581));
	notech_inv i_8907(.A(n_26062), .Z(n_55580));
	notech_inv i_8905(.A(\nbus_11353[0] ), .Z(n_55577));
	notech_inv i_8903(.A(\nbus_11353[0] ), .Z(n_55575));
	notech_inv i_8899(.A(\nbus_11353[0] ), .Z(n_55572));
	notech_inv i_8897(.A(\nbus_11353[0] ), .Z(n_55570));
	notech_inv i_8893(.A(n_55553), .Z(n_55565));
	notech_inv i_8891(.A(n_55553), .Z(n_55564));
	notech_inv i_8886(.A(n_55553), .Z(n_55559));
	notech_inv i_8880(.A(n_55553), .Z(n_55554));
	notech_inv i_8879(.A(n_148482485), .Z(n_55553));
	notech_inv i_8877(.A(n_55540), .Z(n_55550));
	notech_inv i_8875(.A(n_55540), .Z(n_55549));
	notech_inv i_8871(.A(n_55540), .Z(n_55545));
	notech_inv i_8867(.A(n_55540), .Z(n_55542));
	notech_inv i_8866(.A(n_55540), .Z(n_55541));
	notech_inv i_8865(.A(n_255640574), .Z(n_55540));
	notech_inv i_8863(.A(\nbus_11301[0] ), .Z(n_55537));
	notech_inv i_8861(.A(\nbus_11301[0] ), .Z(n_55535));
	notech_inv i_8857(.A(\nbus_11301[0] ), .Z(n_55532));
	notech_inv i_8855(.A(\nbus_11301[0] ), .Z(n_55530));
	notech_inv i_8850(.A(n_55513), .Z(n_55525));
	notech_inv i_8849(.A(n_55513), .Z(n_55524));
	notech_inv i_8843(.A(n_55513), .Z(n_55519));
	notech_inv i_8838(.A(n_55513), .Z(n_55514));
	notech_inv i_8837(.A(n_67341288), .Z(n_55513));
	notech_inv i_8833(.A(n_55497), .Z(n_55509));
	notech_inv i_8832(.A(n_55497), .Z(n_55508));
	notech_inv i_8826(.A(n_55497), .Z(n_55503));
	notech_inv i_8821(.A(n_55497), .Z(n_55498));
	notech_inv i_8819(.A(n_188810100), .Z(n_55497));
	notech_inv i_8811(.A(n_55488), .Z(n_55489));
	notech_inv i_8810(.A(n_148382484), .Z(n_55488));
	notech_inv i_8802(.A(n_55479), .Z(n_55480));
	notech_inv i_8801(.A(n_167885955), .Z(n_55479));
	notech_inv i_8762(.A(n_55437), .Z(n_55438));
	notech_inv i_8761(.A(\nbus_11377[0] ), .Z(n_55437));
	notech_inv i_8753(.A(n_55428), .Z(n_55429));
	notech_inv i_8752(.A(n_58751), .Z(n_55428));
	notech_inv i_8744(.A(n_55419), .Z(n_55420));
	notech_inv i_8743(.A(n_310447752), .Z(n_55419));
	notech_inv i_8733(.A(n_55408), .Z(n_55409));
	notech_inv i_8732(.A(n_310247754), .Z(n_55408));
	notech_inv i_8724(.A(n_55399), .Z(n_55400));
	notech_inv i_8722(.A(n_58750), .Z(n_55399));
	notech_inv i_8712(.A(n_55388), .Z(n_55389));
	notech_inv i_8711(.A(n_58789), .Z(n_55388));
	notech_inv i_8701(.A(n_55377), .Z(n_55378));
	notech_inv i_8700(.A(n_58791), .Z(n_55377));
	notech_inv i_8689(.A(n_55366), .Z(n_55367));
	notech_inv i_8688(.A(n_58788), .Z(n_55366));
	notech_inv i_8670(.A(n_55346), .Z(n_55347));
	notech_inv i_8669(.A(n_310347753), .Z(n_55346));
	notech_inv i_8569(.A(n_55228), .Z(n_55229));
	notech_inv i_8568(.A(n_53341148), .Z(n_55228));
	notech_inv i_8560(.A(n_55219), .Z(n_55220));
	notech_inv i_8559(.A(n_53641151), .Z(n_55219));
	notech_inv i_8549(.A(n_55208), .Z(n_55209));
	notech_inv i_8548(.A(n_53841153), .Z(n_55208));
	notech_inv i_8540(.A(n_55199), .Z(n_55200));
	notech_inv i_8538(.A(n_54141156), .Z(n_55199));
	notech_inv i_8530(.A(n_55190), .Z(n_55191));
	notech_inv i_8529(.A(n_26781), .Z(n_55190));
	notech_inv i_8359(.A(n_55015), .Z(n_55016));
	notech_inv i_8358(.A(\nbus_11297[0] ), .Z(n_55015));
	notech_inv i_8348(.A(n_55004), .Z(n_55005));
	notech_inv i_8347(.A(n_328084271), .Z(n_55004));
	notech_inv i_8326(.A(n_54982), .Z(n_54983));
	notech_inv i_8325(.A(n_27652), .Z(n_54982));
	notech_inv i_8317(.A(n_54973), .Z(n_54974));
	notech_inv i_8316(.A(n_316491659), .Z(n_54973));
	notech_inv i_8305(.A(n_54962), .Z(n_54963));
	notech_inv i_8304(.A(n_27575), .Z(n_54962));
	notech_inv i_8296(.A(n_54953), .Z(n_54954));
	notech_inv i_8295(.A(n_3854), .Z(n_54953));
	notech_inv i_8285(.A(n_54942), .Z(n_54943));
	notech_inv i_8284(.A(n_3816), .Z(n_54942));
	notech_inv i_8276(.A(n_54933), .Z(n_54934));
	notech_inv i_8275(.A(n_26054), .Z(n_54933));
	notech_inv i_8272(.A(n_17107), .Z(n_54930));
	notech_inv i_8271(.A(n_17107), .Z(n_54929));
	notech_inv i_8267(.A(n_17107), .Z(n_54925));
	notech_inv i_8257(.A(n_54915), .Z(n_54916));
	notech_inv i_8256(.A(n_26770), .Z(n_54915));
	notech_inv i_8246(.A(n_54904), .Z(n_54905));
	notech_inv i_8245(.A(n_177458870), .Z(n_54904));
	notech_inv i_8235(.A(n_54893), .Z(n_54894));
	notech_inv i_8233(.A(n_310191722), .Z(n_54893));
	notech_inv i_8223(.A(n_54882), .Z(n_54883));
	notech_inv i_8222(.A(n_146328740), .Z(n_54882));
	notech_inv i_8214(.A(n_54873), .Z(n_54874));
	notech_inv i_8213(.A(n_310291721), .Z(n_54873));
	notech_inv i_8205(.A(n_54864), .Z(n_54865));
	notech_inv i_8204(.A(n_146228739), .Z(n_54864));
	notech_inv i_8193(.A(n_54853), .Z(n_54854));
	notech_inv i_8192(.A(\nbus_11332[0] ), .Z(n_54853));
	notech_inv i_8182(.A(n_54842), .Z(n_54843));
	notech_inv i_8181(.A(n_3815), .Z(n_54842));
	notech_inv i_8173(.A(n_54833), .Z(n_54834));
	notech_inv i_8172(.A(n_1429), .Z(n_54833));
	notech_inv i_8161(.A(n_54822), .Z(n_54823));
	notech_inv i_8159(.A(\nbus_11350[0] ), .Z(n_54822));
	notech_inv i_8151(.A(n_54813), .Z(n_54814));
	notech_inv i_8150(.A(n_58810), .Z(n_54813));
	notech_inv i_8140(.A(n_54802), .Z(n_54803));
	notech_inv i_8139(.A(n_27365), .Z(n_54802));
	notech_inv i_8131(.A(n_54793), .Z(n_54794));
	notech_inv i_8130(.A(n_174962032), .Z(n_54793));
	notech_inv i_8119(.A(n_54782), .Z(n_54783));
	notech_inv i_8118(.A(\nbus_11302[0] ), .Z(n_54782));
	notech_inv i_8110(.A(n_54773), .Z(n_54774));
	notech_inv i_8109(.A(n_286463131), .Z(n_54773));
	notech_inv i_8101(.A(n_54764), .Z(n_54765));
	notech_inv i_8100(.A(n_58805), .Z(n_54764));
	notech_inv i_8092(.A(n_54755), .Z(n_54756));
	notech_inv i_8091(.A(n_58099), .Z(n_54755));
	notech_inv i_8080(.A(n_54744), .Z(n_54745));
	notech_inv i_8079(.A(\nbus_11372[0] ), .Z(n_54744));
	notech_inv i_8071(.A(n_54735), .Z(n_54736));
	notech_inv i_8070(.A(n_58478), .Z(n_54735));
	notech_inv i_8062(.A(n_54726), .Z(n_54727));
	notech_inv i_8061(.A(n_245362720), .Z(n_54726));
	notech_inv i_8053(.A(n_54717), .Z(n_54718));
	notech_inv i_8052(.A(n_58817), .Z(n_54717));
	notech_inv i_8044(.A(n_54708), .Z(n_54709));
	notech_inv i_8043(.A(n_58100), .Z(n_54708));
	notech_inv i_8032(.A(n_54697), .Z(n_54698));
	notech_inv i_8031(.A(\nbus_11373[0] ), .Z(n_54697));
	notech_inv i_8021(.A(n_54686), .Z(n_54687));
	notech_inv i_8020(.A(\nbus_11374[0] ), .Z(n_54686));
	notech_inv i_8012(.A(n_54677), .Z(n_54678));
	notech_inv i_8011(.A(n_58480), .Z(n_54677));
	notech_inv i_8000(.A(n_54666), .Z(n_54667));
	notech_inv i_7999(.A(n_125828535), .Z(n_54666));
	notech_inv i_7991(.A(n_54657), .Z(n_54658));
	notech_inv i_7990(.A(n_27335), .Z(n_54657));
	notech_inv i_7982(.A(n_54648), .Z(n_54649));
	notech_inv i_7981(.A(n_28530), .Z(n_54648));
	notech_inv i_7976(.A(n_54637), .Z(n_54643));
	notech_inv i_7971(.A(n_54637), .Z(n_54638));
	notech_inv i_7970(.A(n_310591718), .Z(n_54637));
	notech_inv i_7951(.A(n_54617), .Z(n_54618));
	notech_inv i_7950(.A(n_27270), .Z(n_54617));
	notech_inv i_7932(.A(n_54545), .Z(n_54546));
	notech_inv i_7931(.A(n_327790775), .Z(n_54545));
	notech_inv i_7920(.A(n_54534), .Z(n_54535));
	notech_inv i_7919(.A(n_327890776), .Z(n_54534));
	notech_inv i_7863(.A(n_54430), .Z(n_54431));
	notech_inv i_7862(.A(n_27107), .Z(n_54430));
	notech_inv i_7852(.A(n_54419), .Z(n_54420));
	notech_inv i_7851(.A(\nbus_11363[0] ), .Z(n_54419));
	notech_inv i_7840(.A(n_54408), .Z(n_54409));
	notech_inv i_7839(.A(n_62041235), .Z(n_54408));
	notech_inv i_7831(.A(n_54399), .Z(n_54400));
	notech_inv i_7830(.A(n_317887452), .Z(n_54399));
	notech_inv i_7820(.A(n_54388), .Z(n_54389));
	notech_inv i_7819(.A(n_328390781), .Z(n_54388));
	notech_inv i_7808(.A(n_54377), .Z(n_54378));
	notech_inv i_7807(.A(n_327990777), .Z(n_54377));
	notech_inv i_7712(.A(n_54145), .Z(n_54146));
	notech_inv i_7711(.A(\nbus_11378[0] ), .Z(n_54145));
	notech_inv i_7681(.A(n_54112), .Z(n_54113));
	notech_inv i_7680(.A(n_154179045), .Z(n_54112));
	notech_inv i_7672(.A(n_54103), .Z(n_54104));
	notech_inv i_7671(.A(n_154279046), .Z(n_54103));
	notech_inv i_7659(.A(n_54092), .Z(n_54093));
	notech_inv i_7658(.A(n_154379047), .Z(n_54092));
	notech_inv i_7647(.A(n_54081), .Z(n_54082));
	notech_inv i_7646(.A(n_326790765), .Z(n_54081));
	notech_inv i_7638(.A(n_54072), .Z(n_54073));
	notech_inv i_7637(.A(n_326890766), .Z(n_54072));
	notech_inv i_7626(.A(n_54061), .Z(n_54062));
	notech_inv i_7625(.A(n_326990767), .Z(n_54061));
	notech_inv i_7615(.A(n_54050), .Z(n_54051));
	notech_inv i_7614(.A(n_136861651), .Z(n_54050));
	notech_inv i_7606(.A(n_54041), .Z(n_54042));
	notech_inv i_7605(.A(n_136761650), .Z(n_54041));
	notech_inv i_7594(.A(n_54030), .Z(n_54031));
	notech_inv i_7593(.A(n_136661649), .Z(n_54030));
	notech_inv i_7583(.A(n_54019), .Z(n_54020));
	notech_inv i_7582(.A(n_349981000), .Z(n_54019));
	notech_inv i_7474(.A(n_53900), .Z(n_53901));
	notech_inv i_7473(.A(n_349780998), .Z(n_53900));
	notech_inv i_7463(.A(n_53889), .Z(n_53890));
	notech_inv i_7462(.A(n_349880999), .Z(n_53889));
	notech_inv i_7408(.A(n_53829), .Z(n_53830));
	notech_inv i_7407(.A(n_152689025), .Z(n_53829));
	notech_inv i_7297(.A(n_53708), .Z(n_53709));
	notech_inv i_7296(.A(n_152789026), .Z(n_53708));
	notech_inv i_7288(.A(n_53699), .Z(n_53700));
	notech_inv i_7287(.A(n_152889027), .Z(n_53699));
	notech_inv i_7279(.A(n_53690), .Z(n_53691));
	notech_inv i_7278(.A(n_140088899), .Z(n_53690));
	notech_inv i_7268(.A(n_53679), .Z(n_53680));
	notech_inv i_7266(.A(n_139788896), .Z(n_53679));
	notech_inv i_7158(.A(n_53560), .Z(n_53561));
	notech_inv i_7157(.A(n_139488893), .Z(n_53560));
	notech_inv i_7146(.A(n_53549), .Z(n_53550));
	notech_inv i_7145(.A(n_324290740), .Z(n_53549));
	notech_inv i_7037(.A(n_53430), .Z(n_53431));
	notech_inv i_7036(.A(n_324190739), .Z(n_53430));
	notech_inv i_7025(.A(n_53419), .Z(n_53420));
	notech_inv i_7024(.A(n_324090738), .Z(n_53419));
	notech_inv i_7016(.A(n_53410), .Z(n_53411));
	notech_inv i_7015(.A(n_315290650), .Z(n_53410));
	notech_inv i_7005(.A(n_53399), .Z(n_53400));
	notech_inv i_7004(.A(n_314990647), .Z(n_53399));
	notech_inv i_6895(.A(n_53280), .Z(n_53281));
	notech_inv i_6894(.A(n_314690644), .Z(n_53280));
	notech_inv i_6884(.A(n_53269), .Z(n_53270));
	notech_inv i_6882(.A(\nbus_11346[0] ), .Z(n_53269));
	notech_inv i_6872(.A(n_53258), .Z(n_53259));
	notech_inv i_6871(.A(n_161285889), .Z(n_53258));
	notech_inv i_6870(.A(n_53253), .Z(n_53256));
	notech_inv i_6869(.A(n_53253), .Z(n_53255));
	notech_inv i_6868(.A(n_53253), .Z(n_53254));
	notech_inv i_6866(.A(n_276490263), .Z(n_53253));
	notech_inv i_6865(.A(n_53249), .Z(n_53252));
	notech_inv i_6864(.A(n_53249), .Z(n_53251));
	notech_inv i_6863(.A(n_53249), .Z(n_53250));
	notech_inv i_6862(.A(n_276490263), .Z(n_53249));
	notech_inv i_6861(.A(n_53244), .Z(n_53247));
	notech_inv i_6860(.A(n_53244), .Z(n_53246));
	notech_inv i_6858(.A(n_53244), .Z(n_53245));
	notech_inv i_6857(.A(n_276990268), .Z(n_53244));
	notech_inv i_6856(.A(n_53240), .Z(n_53243));
	notech_inv i_6855(.A(n_53240), .Z(n_53242));
	notech_inv i_6854(.A(n_53240), .Z(n_53241));
	notech_inv i_6853(.A(n_276990268), .Z(n_53240));
	notech_inv i_6852(.A(n_53234), .Z(n_53238));
	notech_inv i_6850(.A(n_53234), .Z(n_53237));
	notech_inv i_6849(.A(n_53234), .Z(n_53236));
	notech_inv i_6848(.A(n_53234), .Z(n_53235));
	notech_inv i_6847(.A(n_276790266), .Z(n_53234));
	notech_inv i_6846(.A(n_53229), .Z(n_53233));
	notech_inv i_6845(.A(n_53229), .Z(n_53232));
	notech_inv i_6844(.A(n_53229), .Z(n_53231));
	notech_inv i_6842(.A(n_53229), .Z(n_53230));
	notech_inv i_6841(.A(n_276790266), .Z(n_53229));
	notech_inv i_6840(.A(n_53224), .Z(n_53227));
	notech_inv i_6839(.A(n_53224), .Z(n_53226));
	notech_inv i_6838(.A(n_53224), .Z(n_53225));
	notech_inv i_6837(.A(n_276690265), .Z(n_53224));
	notech_inv i_6836(.A(n_53220), .Z(n_53223));
	notech_inv i_6834(.A(n_53220), .Z(n_53222));
	notech_inv i_6833(.A(n_53220), .Z(n_53221));
	notech_inv i_6832(.A(n_276690265), .Z(n_53220));
	notech_inv i_6831(.A(n_53214), .Z(n_53218));
	notech_inv i_6830(.A(n_53214), .Z(n_53217));
	notech_inv i_6829(.A(n_53214), .Z(n_53216));
	notech_inv i_6828(.A(n_53214), .Z(n_53215));
	notech_inv i_6826(.A(n_276090259), .Z(n_53214));
	notech_inv i_6825(.A(n_53209), .Z(n_53213));
	notech_inv i_6824(.A(n_53209), .Z(n_53212));
	notech_inv i_6823(.A(n_53209), .Z(n_53211));
	notech_inv i_6822(.A(n_53209), .Z(n_53210));
	notech_inv i_6821(.A(n_276090259), .Z(n_53209));
	notech_inv i_6820(.A(n_53204), .Z(n_53207));
	notech_inv i_6818(.A(n_53204), .Z(n_53206));
	notech_inv i_6817(.A(n_53204), .Z(n_53205));
	notech_inv i_6816(.A(n_275990258), .Z(n_53204));
	notech_inv i_6815(.A(n_53200), .Z(n_53203));
	notech_inv i_6814(.A(n_53200), .Z(n_53202));
	notech_inv i_6813(.A(n_53200), .Z(n_53201));
	notech_inv i_6812(.A(n_275990258), .Z(n_53200));
	notech_inv i_6810(.A(n_53194), .Z(n_53198));
	notech_inv i_6809(.A(n_53194), .Z(n_53197));
	notech_inv i_6808(.A(n_53194), .Z(n_53196));
	notech_inv i_6807(.A(n_53194), .Z(n_53195));
	notech_inv i_6806(.A(n_275690255), .Z(n_53194));
	notech_inv i_6805(.A(n_53189), .Z(n_53193));
	notech_inv i_6804(.A(n_53189), .Z(n_53192));
	notech_inv i_6802(.A(n_53189), .Z(n_53191));
	notech_inv i_6801(.A(n_53189), .Z(n_53190));
	notech_inv i_6800(.A(n_275690255), .Z(n_53189));
	notech_inv i_6799(.A(n_53184), .Z(n_53187));
	notech_inv i_6798(.A(n_53184), .Z(n_53186));
	notech_inv i_6797(.A(n_53184), .Z(n_53185));
	notech_inv i_6796(.A(n_275390252), .Z(n_53184));
	notech_inv i_6794(.A(n_53180), .Z(n_53183));
	notech_inv i_6793(.A(n_53180), .Z(n_53182));
	notech_inv i_6792(.A(n_53180), .Z(n_53181));
	notech_inv i_6791(.A(n_275390252), .Z(n_53180));
	notech_inv i_6790(.A(n_53175), .Z(n_53178));
	notech_inv i_6789(.A(n_53175), .Z(n_53177));
	notech_inv i_6788(.A(n_53175), .Z(n_53176));
	notech_inv i_6786(.A(n_255190050), .Z(n_53175));
	notech_inv i_6785(.A(n_53171), .Z(n_53174));
	notech_inv i_6784(.A(n_53171), .Z(n_53173));
	notech_inv i_6783(.A(n_53171), .Z(n_53172));
	notech_inv i_6782(.A(n_255190050), .Z(n_53171));
	notech_inv i_6781(.A(n_53166), .Z(n_53169));
	notech_inv i_6780(.A(n_53166), .Z(n_53168));
	notech_inv i_6778(.A(n_53166), .Z(n_53167));
	notech_inv i_6777(.A(n_27078), .Z(n_53166));
	notech_inv i_6776(.A(n_53162), .Z(n_53165));
	notech_inv i_6775(.A(n_53162), .Z(n_53164));
	notech_inv i_6774(.A(n_53162), .Z(n_53163));
	notech_inv i_6773(.A(n_27078), .Z(n_53162));
	notech_inv i_6772(.A(n_53156), .Z(n_53160));
	notech_inv i_6770(.A(n_53156), .Z(n_53159));
	notech_inv i_6769(.A(n_53156), .Z(n_53158));
	notech_inv i_6768(.A(n_53156), .Z(n_53157));
	notech_inv i_6767(.A(n_256090059), .Z(n_53156));
	notech_inv i_6766(.A(n_53151), .Z(n_53155));
	notech_inv i_6765(.A(n_53151), .Z(n_53154));
	notech_inv i_6764(.A(n_53151), .Z(n_53153));
	notech_inv i_6762(.A(n_53151), .Z(n_53152));
	notech_inv i_6761(.A(n_256090059), .Z(n_53151));
	notech_inv i_6760(.A(n_53146), .Z(n_53149));
	notech_inv i_6759(.A(n_53146), .Z(n_53148));
	notech_inv i_6758(.A(n_53146), .Z(n_53147));
	notech_inv i_6757(.A(n_255990058), .Z(n_53146));
	notech_inv i_6756(.A(n_53142), .Z(n_53145));
	notech_inv i_6754(.A(n_53142), .Z(n_53144));
	notech_inv i_6753(.A(n_53142), .Z(n_53143));
	notech_inv i_6752(.A(n_255990058), .Z(n_53142));
	notech_inv i_6751(.A(n_53136), .Z(n_53140));
	notech_inv i_6750(.A(n_53136), .Z(n_53139));
	notech_inv i_6749(.A(n_53136), .Z(n_53138));
	notech_inv i_6748(.A(n_53136), .Z(n_53137));
	notech_inv i_6746(.A(n_255690055), .Z(n_53136));
	notech_inv i_6745(.A(n_53131), .Z(n_53135));
	notech_inv i_6744(.A(n_53131), .Z(n_53134));
	notech_inv i_6743(.A(n_53131), .Z(n_53133));
	notech_inv i_6742(.A(n_53131), .Z(n_53132));
	notech_inv i_6741(.A(n_255690055), .Z(n_53131));
	notech_inv i_6740(.A(n_53126), .Z(n_53129));
	notech_inv i_6738(.A(n_53126), .Z(n_53128));
	notech_inv i_6737(.A(n_53126), .Z(n_53127));
	notech_inv i_6736(.A(n_255390052), .Z(n_53126));
	notech_inv i_6735(.A(n_53122), .Z(n_53125));
	notech_inv i_6734(.A(n_53122), .Z(n_53124));
	notech_inv i_6733(.A(n_53122), .Z(n_53123));
	notech_inv i_6732(.A(n_255390052), .Z(n_53122));
	notech_inv i_6730(.A(n_53116), .Z(n_53120));
	notech_inv i_6729(.A(n_53116), .Z(n_53119));
	notech_inv i_6728(.A(n_53116), .Z(n_53118));
	notech_inv i_6727(.A(n_53116), .Z(n_53117));
	notech_inv i_6726(.A(n_254890047), .Z(n_53116));
	notech_inv i_6725(.A(n_53111), .Z(n_53115));
	notech_inv i_6724(.A(n_53111), .Z(n_53114));
	notech_inv i_6722(.A(n_53111), .Z(n_53113));
	notech_inv i_6721(.A(n_53111), .Z(n_53112));
	notech_inv i_6720(.A(n_254890047), .Z(n_53111));
	notech_inv i_6719(.A(n_52998), .Z(n_53001));
	notech_inv i_6718(.A(n_52998), .Z(n_53000));
	notech_inv i_6717(.A(n_52998), .Z(n_52999));
	notech_inv i_6716(.A(n_254690045), .Z(n_52998));
	notech_inv i_6714(.A(n_52994), .Z(n_52997));
	notech_inv i_6713(.A(n_52994), .Z(n_52996));
	notech_inv i_6712(.A(n_52994), .Z(n_52995));
	notech_inv i_6711(.A(n_254690045), .Z(n_52994));
	notech_and4 i_1021343(.A(n_167665205), .B(n_168465213), .C(n_141964948),
		 .D(n_167565204), .Z(n_21390));
	notech_nand2 i_521338(.A(n_169765226), .B(n_169165220), .Z(n_21360));
	notech_nand2 i_221335(.A(n_171065239), .B(n_170465233), .Z(n_21342));
	notech_and4 i_2221387(.A(n_137764906), .B(n_171565244), .C(n_171765246),
		 .D(n_171465243), .Z(n_25372));
	notech_and4 i_1621381(.A(n_172465253), .B(n_172665255), .C(n_136764896),
		 .D(n_172365252), .Z(n_25336));
	notech_nand2 i_2221547(.A(n_173865267), .B(n_173365262), .Z(n_18258));
	notech_nand2 i_1621541(.A(n_174865277), .B(n_174465273), .Z(n_18222));
	notech_and4 i_1521540(.A(n_175665285), .B(n_175565284), .C(n_175465283),
		 .D(n_175965288), .Z(n_18216));
	notech_nand2 i_1021535(.A(n_176965298), .B(n_176565294), .Z(n_18186));
	notech_and4 i_821533(.A(n_177665305), .B(n_177565304), .C(n_130964838), 
		.D(n_177965308), .Z(n_18174));
	notech_and4 i_2221643(.A(n_178165310), .B(n_178365312), .C(n_178865317),
		 .D(n_130464833), .Z(n_17906));
	notech_nand2 i_3121812(.A(n_179965328), .B(n_179465323), .Z(n_21164));
	notech_nand2 i_2221803(.A(n_181165340), .B(n_180565334), .Z(n_21110));
	notech_nand2 i_1621797(.A(n_182265351), .B(n_181765346), .Z(n_21074));
	notech_and4 i_1521796(.A(n_183165360), .B(n_183065359), .C(n_182965358),
		 .D(n_183565364), .Z(n_21068));
	notech_nand2 i_1321794(.A(n_184865377), .B(n_184265371), .Z(n_21056));
	notech_and4 i_1221793(.A(n_185765386), .B(n_185665385), .C(n_185565384),
		 .D(n_186165390), .Z(n_21050));
	notech_nand2 i_1021791(.A(n_187365402), .B(n_186865397), .Z(n_21038));
	notech_nand2 i_821789(.A(n_188765416), .B(n_188165410), .Z(n_21026));
	notech_nand2 i_2221931(.A(n_189765426), .B(n_189265421), .Z(n_17558));
	notech_nand2 i_2217611(.A(n_190765436), .B(n_190265431), .Z(n_16832));
	notech_and4 i_143841315(.A(n_307766606), .B(n_307666605), .C(n_307266601
		), .D(n_307566604), .Z(n_59962));
	notech_ao4 i_106461762(.A(n_32347), .B(n_59962), .C(n_114464673), .D(n_28000
		), .Z(n_320137996));
	notech_and2 i_061723(.A(n_115964688), .B(n_155565084), .Z(n_316137956)
		);
	notech_and4 i_1221345(.A(n_166865197), .B(n_166765196), .C(n_166665195),
		 .D(n_167165200), .Z(n_21402));
	notech_ao4 i_5947640(.A(n_30821), .B(n_61115), .C(n_303791786), .D(n_299691827
		), .Z(n_57160));
	notech_ao4 i_94461783(.A(n_32348), .B(n_59962), .C(n_58186), .D(n_28000)
		, .Z(n_58105));
	notech_or4 i_160455549(.A(n_306491759), .B(n_308391740), .C(n_48163), .D
		(n_304791776), .Z(n_57481));
	notech_ao4 i_142255547(.A(n_306891755), .B(n_27761), .C(n_306291761), .D
		(n_32382), .Z(n_57627));
	notech_ao4 i_127455546(.A(n_27761), .B(n_27746), .C(n_27754), .D(n_207265601
		), .Z(n_57775));
	notech_and3 i_159555548(.A(n_308291741), .B(n_306691757), .C(n_207365602
		), .Z(n_57490));
	notech_and4 i_133455550(.A(n_56848), .B(n_1441), .C(n_304991774), .D(n_305191772
		), .Z(n_57715));
	notech_and4 i_1421347(.A(n_165565184), .B(n_165465183), .C(n_165365182),
		 .D(n_165965188), .Z(n_21414));
	notech_and4 i_1521348(.A(n_164165170), .B(n_164065169), .C(n_163965168),
		 .D(n_164665175), .Z(n_21420));
	notech_and4 i_1621349(.A(n_162165150), .B(n_162965158), .C(n_146864997),
		 .D(n_162065149), .Z(n_21426));
	notech_nand2 i_2221355(.A(n_161765146), .B(n_161265141), .Z(n_21462));
	notech_nand2 i_1321346(.A(n_201465543), .B(n_200965538), .Z(n_21408));
	notech_nand2 i_1121344(.A(n_202565554), .B(n_202065549), .Z(n_21396));
	notech_and4 i_121334(.A(n_203465563), .B(n_203765566), .C(n_203365562), 
		.D(n_196265491), .Z(n_21336));
	notech_nand2 i_1121792(.A(n_205065579), .B(n_204465573), .Z(n_21044));
	notech_and4 i_121782(.A(n_206465593), .B(n_206665595), .C(n_193365462), 
		.D(n_206365592), .Z(n_20984));
	notech_and3 i_69955544(.A(n_58432), .B(n_304691777), .C(n_207465603), .Z
		(n_58318));
	notech_nand2 i_3121364(.A(n_160665135), .B(n_160165130), .Z(n_21516));
	notech_nand2 i_2621359(.A(n_226765796), .B(n_226265791), .Z(n_21486));
	notech_nand2 i_2521358(.A(n_227765806), .B(n_227265801), .Z(n_21480));
	notech_nand2 i_2421357(.A(n_228765816), .B(n_228265811), .Z(n_21474));
	notech_nand2 i_2321356(.A(n_229765826), .B(n_229265821), .Z(n_21468));
	notech_and4 i_321336(.A(n_230665835), .B(n_230565834), .C(n_230465833), 
		.D(n_231165840), .Z(n_21348));
	notech_nand2 i_2621807(.A(n_232365852), .B(n_231865847), .Z(n_21134));
	notech_nand3 i_29983(.A(n_62826), .B(n_62848), .C(\opa_12[2] ), .Z(n_312347735
		));
	notech_nao3 i_29982(.A(n_62776), .B(\opcode[1] ), .C(n_60023), .Z(n_312447734
		));
	notech_and2 i_850641(.A(n_58717), .B(n_312447734), .Z(n_284927231));
	notech_and2 i_750642(.A(n_58717), .B(n_312347735), .Z(n_285027232));
	notech_and4 i_144550676(.A(n_225265781), .B(n_225165780), .C(n_224765776
		), .D(n_225065779), .Z(n_289227274));
	notech_and4 i_144650675(.A(n_223765766), .B(n_223665765), .C(n_223265761
		), .D(n_223565764), .Z(n_289127273));
	notech_and4 i_144750674(.A(n_222265751), .B(n_222165750), .C(n_221765746
		), .D(n_222065749), .Z(n_289027272));
	notech_and4 i_2221195(.A(n_158965118), .B(n_159165120), .C(n_150465033),
		 .D(n_159665125), .Z(n_18606));
	notech_or4 i_2221099(.A(n_111264641), .B(n_150565034), .C(n_158665115), 
		.D(n_26746), .Z(n_18955));
	notech_and4 i_2221003(.A(n_157265101), .B(n_157465103), .C(n_157965108),
		 .D(n_152365052), .Z(n_23860));
	notech_or4 i_2220875(.A(n_152465053), .B(n_111264641), .C(n_156765096), 
		.D(n_26747), .Z(n_24208));
	notech_and4 i_2220779(.A(n_154065069), .B(n_155665085), .C(n_155865087),
		 .D(n_156365092), .Z(n_24556));
	notech_or4 i_76461766(.A(calc_sz[1]), .B(n_246691943), .C(n_56834), .D(n_59962
		), .Z(n_320538000));
	notech_ao4 i_105061815(.A(n_61115), .B(n_30825), .C(n_26614), .D(n_319291631
		), .Z(n_57999));
	notech_and4 i_144447720(.A(n_252666055), .B(n_252566054), .C(n_252166050
		), .D(n_252466053), .Z(n_59980));
	notech_nand2 i_2121354(.A(n_255466083), .B(n_254966078), .Z(n_21456));
	notech_nand2 i_2021353(.A(n_256566094), .B(n_256066089), .Z(n_21450));
	notech_nand2 i_1921352(.A(n_257666105), .B(n_257166100), .Z(n_21444));
	notech_nand2 i_1821351(.A(n_258766116), .B(n_258266111), .Z(n_21438));
	notech_and4 i_1721350(.A(n_259266121), .B(n_259966128), .C(n_242565954),
		 .D(n_259066119), .Z(n_21432));
	notech_nand2 i_2121802(.A(n_261066139), .B(n_260566134), .Z(n_21104));
	notech_nand2 i_2021801(.A(n_262266151), .B(n_261666145), .Z(n_21098));
	notech_nand2 i_1921800(.A(n_263466163), .B(n_262866157), .Z(n_21092));
	notech_nand2 i_1821799(.A(n_264666175), .B(n_264066169), .Z(n_21086));
	notech_nand2 i_1721798(.A(n_265966188), .B(n_265366182), .Z(n_21080));
	notech_nand2 i_2221867(.A(n_266866197), .B(n_266466193), .Z(n_20744));
	notech_or4 i_30747697(.A(n_60970), .B(n_60959), .C(\opcode[1] ), .D(\nbus_11365[16] 
		), .Z(n_312324377));
	notech_ao4 i_3747662(.A(n_30821), .B(\nbus_11365[16] ), .C(n_30822), .D(\nbus_11358[16] 
		), .Z(n_307624340));
	notech_and2 i_104961816(.A(n_2991), .B(n_347066999), .Z(n_58000));
	notech_and4 i_143947711(.A(n_254166070), .B(n_254066069), .C(n_253666065
		), .D(n_253966068), .Z(n_313747721));
	notech_and3 i_65061829(.A(n_313191692), .B(n_154865077), .C(n_310391720)
		, .Z(n_58367));
	notech_and2 i_2964424(.A(n_58106), .B(n_109364622), .Z(n_252740545));
	notech_and4 i_1020767(.A(n_200065529), .B(n_110664635), .C(n_109464623),
		 .D(n_110564634), .Z(n_24484));
	notech_and3 i_116444550(.A(n_312991694), .B(n_28222), .C(n_270466233), .Z
		(n_57885));
	notech_and2 i_116344549(.A(n_298991830), .B(n_270366232), .Z(n_57886));
	notech_and4 i_3221365(.A(n_283766366), .B(n_283966368), .C(n_284466373),
		 .D(n_279866327), .Z(n_21522));
	notech_and4 i_721340(.A(n_284766376), .B(n_285066379), .C(n_285666385), 
		.D(n_26673), .Z(n_21372));
	notech_nand2 i_621339(.A(n_286966398), .B(n_286366392), .Z(n_21366));
	notech_nand2 i_421337(.A(n_288266411), .B(n_287666405), .Z(n_21354));
	notech_nand2 i_3221813(.A(n_289466423), .B(n_288966418), .Z(n_21170));
	notech_nand2 i_721788(.A(n_290666435), .B(n_290166430), .Z(n_21020));
	notech_nand2 i_621787(.A(n_292066449), .B(n_291366442), .Z(n_21014));
	notech_nand3 i_12203(.A(n_60153), .B(n_60340), .C(n_269266221), .Z(n_306121225
		));
	notech_and2 i_4644448(.A(n_284966378), .B(n_269766226), .Z(n_303221196)
		);
	notech_nand2 i_2218027(.A(n_109264621), .B(n_109164620), .Z(write_data_26
		[21]));
	notech_and4 i_142844500(.A(n_283466363), .B(n_283366362), .C(n_282966358
		), .D(n_283266361), .Z(n_308621250));
	notech_and3 i_85032005(.A(n_111364642), .B(n_348467013), .C(n_345166980)
		, .Z(n_348667015));
	notech_ao4 i_84932006(.A(n_345066979), .B(\nbus_11358[13] ), .C(n_344966978
		), .D(\nbus_11307[13] ), .Z(n_348467013));
	notech_and4 i_142441325(.A(n_304966578), .B(n_304866577), .C(n_304466573
		), .D(n_304766576), .Z(n_59992));
	notech_and4 i_143741316(.A(n_306366592), .B(n_306266591), .C(n_305866587
		), .D(n_306166590), .Z(n_59963));
	notech_or4 i_39541310(.A(n_60970), .B(n_60959), .C(n_62836), .D(n_29754)
		, .Z(n_58622));
	notech_ao4 i_85132004(.A(n_31540), .B(n_26616), .C(n_27998), .D(n_344866977
		), .Z(n_348267011));
	notech_nand2 i_921342(.A(n_310766636), .B(n_310266631), .Z(n_21384));
	notech_nand2 i_921790(.A(n_311966648), .B(n_311366642), .Z(n_21032));
	notech_and4 i_143141289(.A(n_309366622), .B(n_309266621), .C(n_308866617
		), .D(n_309166620), .Z(n_293018129));
	notech_ao4 i_85232003(.A(n_146328740), .B(n_28606), .C(n_146228739), .D(n_29870
		), .Z(n_348167010));
	notech_and4 i_86731994(.A(n_347867007), .B(n_347767006), .C(n_347567004)
		, .D(n_347467003), .Z(n_348067009));
	notech_ao4 i_85532000(.A(n_31560), .B(n_344666975), .C(n_310291721), .D(n_28102
		), .Z(n_347867007));
	notech_ao4 i_85631999(.A(n_310191722), .B(n_27449), .C(n_313191692), .D(n_301691807
		), .Z(n_347767006));
	notech_ao4 i_85831997(.A(n_30109), .B(n_346866997), .C(n_346766996), .D(n_31576
		), .Z(n_347567004));
	notech_ao4 i_86331996(.A(n_302091803), .B(n_267466203), .C(n_346666995),
		 .D(n_29592), .Z(n_347467003));
	notech_or2 i_10383(.A(n_26611), .B(n_26614), .Z(n_347066999));
	notech_and4 i_91238299(.A(n_330366832), .B(n_330266831), .C(n_329866827)
		, .D(n_330166830), .Z(n_60024));
	notech_and4 i_91638295(.A(n_331766846), .B(n_331666845), .C(n_331266841)
		, .D(n_331566844), .Z(n_60020));
	notech_and4 i_91938292(.A(n_333166860), .B(n_333066859), .C(n_332666855)
		, .D(n_332966858), .Z(n_5933));
	notech_and4 i_92538287(.A(n_334566874), .B(n_334466873), .C(n_334066869)
		, .D(n_334366872), .Z(n_60011));
	notech_and4 i_92638285(.A(n_335966888), .B(n_335866887), .C(n_335466883)
		, .D(n_335766886), .Z(n_60010));
	notech_and4 i_92738284(.A(n_337366902), .B(n_337266901), .C(n_336866897)
		, .D(n_337166900), .Z(n_60009));
	notech_and4 i_93238279(.A(n_338766916), .B(n_338666915), .C(n_338266911)
		, .D(n_338566914), .Z(n_60004));
	notech_and4 i_93338278(.A(n_340166930), .B(n_340066929), .C(n_339666925)
		, .D(n_339966928), .Z(n_60003));
	notech_and4 i_93438277(.A(n_341566944), .B(n_341466943), .C(n_341066939)
		, .D(n_341366942), .Z(n_60002));
	notech_and4 i_93538276(.A(n_342966958), .B(n_342866957), .C(n_342466953)
		, .D(n_342766956), .Z(n_60001));
	notech_nand2 i_2216235(.A(n_344266971), .B(n_343766966), .Z(n_19232));
	notech_nand3 i_30035145(.A(n_60909), .B(\opcode[2] ), .C(\opa_12[2] ), .Z
		(n_58717));
	notech_or4 i_30335124(.A(n_60970), .B(n_60959), .C(n_62836), .D(n_29733)
		, .Z(n_58714));
	notech_or4 i_29986(.A(n_60970), .B(n_60959), .C(n_60909), .D(n_29733), .Z
		(n_312147737));
	notech_or2 i_10385(.A(n_26614), .B(n_312091703), .Z(n_346966998));
	notech_or4 i_33601(.A(n_344766976), .B(n_57087), .C(instrc[116]), .D(n_26770
		), .Z(n_346866997));
	notech_or2 i_33613(.A(n_26616), .B(n_17107), .Z(n_346766996));
	notech_and4 i_1421795(.A(n_348267011), .B(n_348167010), .C(n_348067009),
		 .D(n_348667015), .Z(n_21062));
	notech_or2 i_33617(.A(n_26616), .B(n_317191652), .Z(n_346666995));
	notech_nand2 i_45432353(.A(sav_esp[13]), .B(n_61142), .Z(n_345166980));
	notech_and4 i_109632891(.A(n_312991694), .B(n_299591828), .C(n_347066999
		), .D(n_116164690), .Z(n_345066979));
	notech_and3 i_109532890(.A(n_2993), .B(n_346966998), .C(n_344566974), .Z
		(n_344966978));
	notech_and2 i_63732888(.A(n_310391720), .B(n_313091693), .Z(n_344866977)
		);
	notech_and3 i_21632554(.A(n_26613), .B(n_312191702), .C(n_26614), .Z(n_344766976
		));
	notech_or4 i_166032760(.A(n_26616), .B(n_57087), .C(n_57068), .D(n_26770
		), .Z(n_344666975));
	notech_nand2 i_114732860(.A(n_27109), .B(n_281666345), .Z(n_344566974)
		);
	notech_or2 i_29985(.A(n_60023), .B(n_60868), .Z(n_344466973));
	notech_nand2 i_29991(.A(opc_10[2]), .B(\opcode[2] ), .Z(n_344366972));
	notech_and4 i_158336722(.A(n_277183762), .B(n_344066969), .C(n_343866967
		), .D(n_312466653), .Z(n_344266971));
	notech_ao4 i_157936726(.A(n_3882), .B(n_29238), .C(n_52112621), .D(n_29202
		), .Z(n_344066969));
	notech_ao4 i_158136724(.A(n_53412634), .B(n_29636), .C(n_53512635), .D(n_28006
		), .Z(n_343866967));
	notech_and4 i_158936716(.A(n_343566964), .B(n_343366962), .C(n_343266961
		), .D(n_312766656), .Z(n_343766966));
	notech_ao4 i_158436721(.A(n_54012640), .B(n_29273), .C(n_388360286), .D(nbus_11295
		[21]), .Z(n_343566964));
	notech_ao4 i_158636719(.A(n_310315179), .B(\nbus_11358[21] ), .C(n_3887)
		, .D(n_29075), .Z(n_343366962));
	notech_ao4 i_158736718(.A(n_276383754), .B(n_29012), .C(n_3888), .D(n_28110
		), .Z(n_343266961));
	notech_ao4 i_177836529(.A(n_57985), .B(n_28314), .C(n_27104), .D(n_28508
		), .Z(n_342966958));
	notech_ao4 i_177936528(.A(n_58014), .B(n_27886), .C(n_56468), .D(n_29841
		), .Z(n_342866957));
	notech_and2 i_178336524(.A(n_342666955), .B(n_342566954), .Z(n_342766956
		));
	notech_ao4 i_178136526(.A(n_56401), .B(n_28182), .C(n_28411), .D(n_56390
		), .Z(n_342666955));
	notech_ao4 i_178236525(.A(n_59349), .B(n_28550), .C(n_26664), .D(n_28347
		), .Z(n_342566954));
	notech_and4 i_179136516(.A(n_342266951), .B(n_342166950), .C(n_341966948
		), .D(n_341866947), .Z(n_342466953));
	notech_ao4 i_178536522(.A(n_56457), .B(n_28281), .C(n_27089), .D(n_28475
		), .Z(n_342266951));
	notech_ao4 i_178636521(.A(n_56448), .B(n_28249), .C(n_56437), .D(n_28214
		), .Z(n_342166950));
	notech_ao4 i_178836519(.A(n_56909), .B(n_29840), .C(n_56428), .D(n_28379
		), .Z(n_341966948));
	notech_ao4 i_178936518(.A(n_27094), .B(n_28443), .C(n_26950), .D(n_28585
		), .Z(n_341866947));
	notech_ao4 i_179236515(.A(n_57985), .B(n_28313), .C(n_60845), .D(n_28507
		), .Z(n_341566944));
	notech_ao4 i_179336514(.A(n_58014), .B(n_27884), .C(n_56468), .D(n_29839
		), .Z(n_341466943));
	notech_and2 i_179736510(.A(n_341266941), .B(n_341166940), .Z(n_341366942
		));
	notech_ao4 i_179536512(.A(n_56400), .B(n_28181), .C(n_28410), .D(n_56390
		), .Z(n_341266941));
	notech_ao4 i_179636511(.A(n_59349), .B(n_28549), .C(n_56371), .D(n_28346
		), .Z(n_341166940));
	notech_and4 i_180536502(.A(n_340866937), .B(n_340766936), .C(n_340566934
		), .D(n_340466933), .Z(n_341066939));
	notech_ao4 i_179936508(.A(n_56457), .B(n_28280), .C(n_58024), .D(n_28474
		), .Z(n_340866937));
	notech_ao4 i_180036507(.A(n_56447), .B(n_28248), .C(n_56437), .D(n_28213
		), .Z(n_340766936));
	notech_ao4 i_180236505(.A(n_56909), .B(n_29838), .C(n_56427), .D(n_28378
		), .Z(n_340566934));
	notech_ao4 i_180336504(.A(n_27094), .B(n_28442), .C(n_26950), .D(n_28584
		), .Z(n_340466933));
	notech_ao4 i_180636501(.A(n_57985), .B(n_28312), .C(n_27104), .D(n_28506
		), .Z(n_340166930));
	notech_ao4 i_180736500(.A(n_58014), .B(n_27883), .C(n_56468), .D(n_29837
		), .Z(n_340066929));
	notech_and2 i_181236496(.A(n_339866927), .B(n_339766926), .Z(n_339966928
		));
	notech_ao4 i_181036498(.A(n_56401), .B(n_28180), .C(n_28409), .D(n_56390
		), .Z(n_339866927));
	notech_ao4 i_181136497(.A(n_59349), .B(n_28548), .C(n_26664), .D(n_28345
		), .Z(n_339766926));
	notech_and4 i_182036488(.A(n_339466923), .B(n_339366922), .C(n_339166920
		), .D(n_339066919), .Z(n_339666925));
	notech_ao4 i_181436494(.A(n_56457), .B(n_28279), .C(n_27089), .D(n_28473
		), .Z(n_339466923));
	notech_ao4 i_181536493(.A(n_56448), .B(n_28247), .C(n_56437), .D(n_28212
		), .Z(n_339366922));
	notech_ao4 i_181736491(.A(n_56909), .B(n_29835), .C(n_56428), .D(n_28377
		), .Z(n_339166920));
	notech_ao4 i_181836490(.A(n_27094), .B(n_28441), .C(n_26950), .D(n_28583
		), .Z(n_339066919));
	notech_ao4 i_182136487(.A(n_57985), .B(n_28311), .C(n_27104), .D(n_28505
		), .Z(n_338766916));
	notech_ao4 i_182236486(.A(n_58014), .B(n_27882), .C(n_56468), .D(n_29855
		), .Z(n_338666915));
	notech_and2 i_182636482(.A(n_338466913), .B(n_338366912), .Z(n_338566914
		));
	notech_ao4 i_182436484(.A(n_56401), .B(n_28179), .C(n_56390), .D(n_28408
		), .Z(n_338466913));
	notech_ao4 i_182536483(.A(n_28547), .B(n_59349), .C(n_26664), .D(n_28344
		), .Z(n_338366912));
	notech_and4 i_183436474(.A(n_338066909), .B(n_337966908), .C(n_337766906
		), .D(n_337666905), .Z(n_338266911));
	notech_ao4 i_182836480(.A(n_56457), .B(n_28278), .C(n_27089), .D(n_28472
		), .Z(n_338066909));
	notech_ao4 i_182936479(.A(n_56448), .B(n_28246), .C(n_56437), .D(n_28211
		), .Z(n_337966908));
	notech_ao4 i_183136477(.A(n_56909), .B(n_29854), .C(n_56428), .D(n_28376
		), .Z(n_337766906));
	notech_ao4 i_183236476(.A(n_27094), .B(n_28440), .C(n_26950), .D(n_28582
		), .Z(n_337666905));
	notech_ao4 i_187736431(.A(n_57985), .B(n_28306), .C(n_27104), .D(n_28499
		), .Z(n_337366902));
	notech_ao4 i_187836430(.A(n_58014), .B(n_27874), .C(n_56468), .D(n_29853
		), .Z(n_337266901));
	notech_and2 i_188236426(.A(n_337066899), .B(n_336966898), .Z(n_337166900
		));
	notech_ao4 i_188036428(.A(n_56401), .B(n_28174), .C(n_56390), .D(n_28403
		), .Z(n_337066899));
	notech_ao4 i_188136427(.A(n_28537), .B(n_59349), .C(n_26664), .D(n_28339
		), .Z(n_336966898));
	notech_and4 i_189036418(.A(n_336666895), .B(n_336566894), .C(n_336366892
		), .D(n_336266891), .Z(n_336866897));
	notech_ao4 i_188436424(.A(n_56457), .B(n_28273), .C(n_27089), .D(n_28467
		), .Z(n_336666895));
	notech_ao4 i_188536423(.A(n_56448), .B(n_28241), .C(n_56437), .D(n_28206
		), .Z(n_336566894));
	notech_ao4 i_188736421(.A(n_56909), .B(n_29852), .C(n_56428), .D(n_28371
		), .Z(n_336366892));
	notech_ao4 i_188836420(.A(n_27094), .B(n_28435), .C(n_26950), .D(n_28577
		), .Z(n_336266891));
	notech_ao4 i_189136417(.A(n_57985), .B(n_28305), .C(n_60845), .D(n_28498
		), .Z(n_335966888));
	notech_ao4 i_189236416(.A(n_58014), .B(n_27873), .C(n_56468), .D(n_29866
		), .Z(n_335866887));
	notech_and2 i_189636412(.A(n_335666885), .B(n_335566884), .Z(n_335766886
		));
	notech_ao4 i_189436414(.A(n_56400), .B(n_28173), .C(n_28402), .D(n_56390
		), .Z(n_335666885));
	notech_ao4 i_189536413(.A(n_59349), .B(n_28536), .C(n_56371), .D(n_28338
		), .Z(n_335566884));
	notech_and4 i_190436404(.A(n_335266881), .B(n_335166880), .C(n_334966878
		), .D(n_334866877), .Z(n_335466883));
	notech_ao4 i_189836410(.A(n_56457), .B(n_28272), .C(n_58024), .D(n_28466
		), .Z(n_335266881));
	notech_ao4 i_189936409(.A(n_56447), .B(n_28240), .C(n_56437), .D(n_28205
		), .Z(n_335166880));
	notech_ao4 i_190136407(.A(n_56909), .B(n_29865), .C(n_56427), .D(n_28370
		), .Z(n_334966878));
	notech_ao4 i_190236406(.A(n_27094), .B(n_28434), .C(n_26950), .D(n_28576
		), .Z(n_334866877));
	notech_ao4 i_190536403(.A(n_57985), .B(n_28304), .C(n_60845), .D(n_28497
		), .Z(n_334566874));
	notech_ao4 i_190636402(.A(n_58014), .B(n_27872), .C(n_56468), .D(n_29868
		), .Z(n_334466873));
	notech_and2 i_191036398(.A(n_334266871), .B(n_334166870), .Z(n_334366872
		));
	notech_ao4 i_190836400(.A(n_56400), .B(n_28172), .C(n_28401), .D(n_56390
		), .Z(n_334266871));
	notech_ao4 i_190936399(.A(n_28535), .B(n_59349), .C(n_56371), .D(n_28337
		), .Z(n_334166870));
	notech_and4 i_191836390(.A(n_333866867), .B(n_333766866), .C(n_333566864
		), .D(n_333466863), .Z(n_334066869));
	notech_ao4 i_191236396(.A(n_56457), .B(n_28271), .C(n_58024), .D(n_28465
		), .Z(n_333866867));
	notech_ao4 i_191336395(.A(n_56447), .B(n_28239), .C(n_56437), .D(n_28204
		), .Z(n_333766866));
	notech_ao4 i_191536393(.A(n_56908), .B(n_29867), .C(n_56427), .D(n_28369
		), .Z(n_333566864));
	notech_ao4 i_191636392(.A(n_27094), .B(n_28433), .C(n_26950), .D(n_28575
		), .Z(n_333466863));
	notech_ao4 i_197536333(.A(n_57985), .B(n_28297), .C(n_60845), .D(n_28491
		), .Z(n_333166860));
	notech_ao4 i_197636332(.A(n_58014), .B(n_27866), .C(n_56468), .D(n_29864
		), .Z(n_333066859));
	notech_and2 i_198036328(.A(n_332866857), .B(n_332766856), .Z(n_332966858
		));
	notech_ao4 i_197836330(.A(n_56400), .B(n_28166), .C(n_28395), .D(n_56390
		), .Z(n_332866857));
	notech_ao4 i_197936329(.A(n_59349), .B(n_28525), .C(n_56371), .D(n_28330
		), .Z(n_332766856));
	notech_and4 i_198836320(.A(n_332466853), .B(n_332366852), .C(n_332166850
		), .D(n_332066849), .Z(n_332666855));
	notech_ao4 i_198236326(.A(n_56457), .B(n_28265), .C(n_58024), .D(n_28459
		), .Z(n_332466853));
	notech_ao4 i_198336325(.A(n_56447), .B(n_28231), .C(n_56437), .D(n_28198
		), .Z(n_332366852));
	notech_ao4 i_198536323(.A(n_56908), .B(n_29863), .C(n_56427), .D(n_28363
		), .Z(n_332166850));
	notech_ao4 i_198636322(.A(n_27094), .B(n_28427), .C(n_26950), .D(n_28568
		), .Z(n_332066849));
	notech_ao4 i_201736291(.A(n_57985), .B(n_28294), .C(n_60845), .D(n_28488
		), .Z(n_331766846));
	notech_ao4 i_201836290(.A(n_58014), .B(n_27863), .C(n_56468), .D(n_29860
		), .Z(n_331666845));
	notech_and2 i_202236286(.A(n_331466843), .B(n_331366842), .Z(n_331566844
		));
	notech_ao4 i_202036288(.A(n_56400), .B(n_28163), .C(n_28392), .D(n_56390
		), .Z(n_331466843));
	notech_ao4 i_202136287(.A(n_59349), .B(n_28521), .C(n_56371), .D(n_28327
		), .Z(n_331366842));
	notech_and4 i_203036278(.A(n_331066839), .B(n_330966838), .C(n_330766836
		), .D(n_330666835), .Z(n_331266841));
	notech_ao4 i_202436284(.A(n_56457), .B(n_28262), .C(n_58024), .D(n_28456
		), .Z(n_331066839));
	notech_ao4 i_202536283(.A(n_56447), .B(n_28228), .C(n_56437), .D(n_28195
		), .Z(n_330966838));
	notech_ao4 i_202736281(.A(n_56908), .B(n_29859), .C(n_56427), .D(n_28360
		), .Z(n_330766836));
	notech_ao4 i_202836280(.A(n_27094), .B(n_28424), .C(n_26950), .D(n_28565
		), .Z(n_330666835));
	notech_ao4 i_205936249(.A(n_57985), .B(n_28290), .C(n_60845), .D(n_28484
		), .Z(n_330366832));
	notech_ao4 i_206036248(.A(n_58014), .B(n_27859), .C(n_56468), .D(n_29869
		), .Z(n_330266831));
	notech_and2 i_206436244(.A(n_330066829), .B(n_329966828), .Z(n_330166830
		));
	notech_ao4 i_206236246(.A(n_56400), .B(n_28159), .C(n_28388), .D(n_56390
		), .Z(n_330066829));
	notech_ao4 i_206336245(.A(n_59349), .B(n_28517), .C(n_56371), .D(n_28323
		), .Z(n_329966828));
	notech_and4 i_207236236(.A(n_329666825), .B(n_329566824), .C(n_329366822
		), .D(n_329266821), .Z(n_329866827));
	notech_ao4 i_206636242(.A(n_56457), .B(n_28258), .C(n_58024), .D(n_28452
		), .Z(n_329666825));
	notech_ao4 i_206736241(.A(n_56447), .B(n_28224), .C(n_56437), .D(n_28191
		), .Z(n_329566824));
	notech_ao4 i_206936239(.A(n_56908), .B(n_27851), .C(n_56427), .D(n_28356
		), .Z(n_329366822));
	notech_ao4 i_207036238(.A(n_27094), .B(n_28420), .C(n_26950), .D(n_28561
		), .Z(n_329266821));
	notech_or2 i_49137775(.A(n_54212642), .B(\nbus_11365[21] ), .Z(n_312766656
		));
	notech_or2 i_49437772(.A(n_53612636), .B(n_60004), .Z(n_312466653));
	notech_and4 i_156639815(.A(n_311766646), .B(n_311566644), .C(n_311466643
		), .D(n_293366462), .Z(n_311966648));
	notech_ao4 i_156139820(.A(n_146328740), .B(n_28601), .C(n_146228739), .D
		(n_29861), .Z(n_311766646));
	notech_ao4 i_156339818(.A(n_5933), .B(n_292366452), .C(n_292266451), .D(n_29787
		), .Z(n_311566644));
	notech_ao4 i_156439817(.A(n_345066979), .B(\nbus_11358[8] ), .C(n_344866977
		), .D(n_27991), .Z(n_311466643));
	notech_and4 i_157239809(.A(n_311166640), .B(n_310966638), .C(n_310866637
		), .D(n_294066469), .Z(n_311366642));
	notech_ao4 i_156739814(.A(n_344966978), .B(\nbus_11307[8] ), .C(n_60153)
		, .D(n_27164), .Z(n_311166640));
	notech_ao4 i_156939812(.A(n_293018129), .B(n_313191692), .C(n_346866997)
		, .D(n_309666625), .Z(n_310966638));
	notech_ao4 i_157039811(.A(n_308066609), .B(n_344666975), .C(n_26616), .D
		(n_308166610), .Z(n_310866637));
	notech_and4 i_160839775(.A(n_294766476), .B(n_310566634), .C(n_310366632
		), .D(n_295066479), .Z(n_310766636));
	notech_ao4 i_160439779(.A(n_28530), .B(n_29862), .C(n_32270), .D(n_28097
		), .Z(n_310566634));
	notech_ao4 i_160639777(.A(n_292866457), .B(n_29787), .C(n_5933), .D(n_292766456
		), .Z(n_310366632));
	notech_and4 i_161539769(.A(n_310066629), .B(n_309866627), .C(n_309766626
		), .D(n_295366482), .Z(n_310266631));
	notech_ao4 i_161039774(.A(n_292566454), .B(\nbus_11307[8] ), .C(n_292466453
		), .D(n_27991), .Z(n_310066629));
	notech_ao4 i_161239772(.A(n_293018129), .B(n_297466503), .C(n_308066609)
		, .D(n_297566504), .Z(n_309866627));
	notech_ao4 i_161339771(.A(n_308166610), .B(n_28545), .C(n_309666625), .D
		(n_292166450), .Z(n_309766626));
	notech_nand2 i_3441288(.A(opc[8]), .B(\opcode[2] ), .Z(n_309666625));
	notech_ao4 i_172139666(.A(n_26924), .B(n_28231), .C(n_26922), .D(n_28198
		), .Z(n_309366622));
	notech_ao4 i_172239665(.A(n_56919), .B(n_29863), .C(n_26969), .D(n_28265
		), .Z(n_309266621));
	notech_and2 i_172639661(.A(n_309066619), .B(n_308966618), .Z(n_309166620
		));
	notech_ao4 i_172439663(.A(n_26927), .B(n_28297), .C(n_26649), .D(n_29864
		), .Z(n_309066619));
	notech_ao4 i_172539662(.A(n_26920), .B(n_28363), .C(n_26933), .D(n_28330
		), .Z(n_308966618));
	notech_and4 i_173439653(.A(n_308666615), .B(n_308566614), .C(n_308366612
		), .D(n_308266611), .Z(n_308866617));
	notech_ao4 i_172839659(.A(n_56630), .B(n_28427), .C(n_56619), .D(n_28395
		), .Z(n_308666615));
	notech_ao4 i_172939658(.A(n_26928), .B(n_28459), .C(n_26651), .D(n_28166
		), .Z(n_308566614));
	notech_ao4 i_173139656(.A(n_26925), .B(n_28491), .C(n_27036), .D(n_28525
		), .Z(n_308366612));
	notech_ao4 i_173239655(.A(n_26721), .B(n_27866), .C(n_56548), .D(n_28568
		), .Z(n_308266611));
	notech_or4 i_40841283(.A(n_60970), .B(n_60959), .C(n_62836), .D(n_29787)
		, .Z(n_308166610));
	notech_nand2 i_39241284(.A(opc_10[8]), .B(\opcode[2] ), .Z(n_308066609)
		);
	notech_ao4 i_186939524(.A(n_26924), .B(n_28240), .C(n_26922), .D(n_28205
		), .Z(n_307766606));
	notech_ao4 i_187039523(.A(n_56919), .B(n_29865), .C(n_56640), .D(n_28272
		), .Z(n_307666605));
	notech_and2 i_187439519(.A(n_307466603), .B(n_307366602), .Z(n_307566604
		));
	notech_ao4 i_187239521(.A(n_26927), .B(n_28305), .C(n_56518), .D(n_29866
		), .Z(n_307466603));
	notech_ao4 i_187339520(.A(n_26920), .B(n_28370), .C(n_26933), .D(n_28338
		), .Z(n_307366602));
	notech_and4 i_188239511(.A(n_307066599), .B(n_306966598), .C(n_306766596
		), .D(n_306666595), .Z(n_307266601));
	notech_ao4 i_187639517(.A(n_56630), .B(n_28434), .C(n_56619), .D(n_28402
		), .Z(n_307066599));
	notech_ao4 i_187739516(.A(n_26928), .B(n_28466), .C(n_26651), .D(n_28173
		), .Z(n_306966598));
	notech_ao4 i_187939514(.A(n_26925), .B(n_28498), .C(n_56570), .D(n_28536
		), .Z(n_306766596));
	notech_ao4 i_188039513(.A(n_56557), .B(n_27873), .C(n_56548), .D(n_28576
		), .Z(n_306666595));
	notech_ao4 i_188339510(.A(n_56666), .B(n_28239), .C(n_56653), .D(n_28204
		), .Z(n_306366592));
	notech_ao4 i_188439509(.A(n_56919), .B(n_29867), .C(n_56640), .D(n_28271
		), .Z(n_306266591));
	notech_and2 i_188839505(.A(n_306066589), .B(n_305966588), .Z(n_306166590
		));
	notech_ao4 i_188639507(.A(n_56532), .B(n_28304), .C(n_56518), .D(n_29868
		), .Z(n_306066589));
	notech_ao4 i_188739506(.A(n_56502), .B(n_28369), .C(n_56489), .D(n_28337
		), .Z(n_305966588));
	notech_and4 i_189739497(.A(n_305666585), .B(n_305566584), .C(n_305366582
		), .D(n_305266581), .Z(n_305866587));
	notech_ao4 i_189039503(.A(n_56630), .B(n_28433), .C(n_56619), .D(n_28401
		), .Z(n_305666585));
	notech_ao4 i_189139502(.A(n_56605), .B(n_28465), .C(n_26651), .D(n_28172
		), .Z(n_305566584));
	notech_ao4 i_189439500(.A(n_56583), .B(n_28497), .C(n_56570), .D(n_28535
		), .Z(n_305366582));
	notech_ao4 i_189539499(.A(n_26721), .B(n_27872), .C(n_56548), .D(n_28575
		), .Z(n_305266581));
	notech_ao4 i_198039420(.A(n_28224), .B(n_26924), .C(n_28191), .D(n_26922
		), .Z(n_304966578));
	notech_ao4 i_198139419(.A(n_56919), .B(n_27851), .C(n_28258), .D(n_26969
		), .Z(n_304866577));
	notech_and2 i_198539415(.A(n_304666575), .B(n_304566574), .Z(n_304766576
		));
	notech_ao4 i_198339417(.A(n_28290), .B(n_26927), .C(n_26649), .D(n_29869
		), .Z(n_304666575));
	notech_ao4 i_198439416(.A(n_26920), .B(n_28356), .C(n_26933), .D(n_28323
		), .Z(n_304566574));
	notech_and4 i_199439407(.A(n_304266571), .B(n_304166570), .C(n_303966568
		), .D(n_303866567), .Z(n_304466573));
	notech_ao4 i_198739413(.A(n_28420), .B(n_56630), .C(n_56619), .D(n_28388
		), .Z(n_304266571));
	notech_ao4 i_198839412(.A(n_26928), .B(n_28452), .C(n_26651), .D(n_28159
		), .Z(n_304166570));
	notech_ao4 i_199039410(.A(n_28484), .B(n_26925), .C(n_27036), .D(n_28517
		), .Z(n_303966568));
	notech_ao4 i_199139409(.A(n_26721), .B(n_27859), .C(n_56548), .D(n_28561
		), .Z(n_303866567));
	notech_or2 i_99640330(.A(n_28544), .B(n_299891825), .Z(n_303466563));
	notech_or4 i_99140331(.A(n_56834), .B(n_26962), .C(n_61142), .D(n_27036)
		, .Z(n_303366562));
	notech_nand2 i_28324(.A(opc_10[15]), .B(\opcode[2] ), .Z(n_298466513));
	notech_nand3 i_28352(.A(n_60909), .B(n_62794), .C(\opa_12[14] ), .Z(n_298366512
		));
	notech_nand2 i_28372(.A(opc_10[14]), .B(n_62794), .Z(n_298266511));
	notech_or4 i_28392(.A(n_60970), .B(n_60959), .C(n_62836), .D(n_29680), .Z
		(n_298166510));
	notech_nand2 i_28956(.A(opc_10[1]), .B(n_62794), .Z(n_298066509));
	notech_nand2 i_28957(.A(opc[1]), .B(n_62794), .Z(n_297966508));
	notech_nao3 i_28960(.A(n_62776), .B(opa[1]), .C(n_62836), .Z(n_297866507
		));
	notech_or4 i_28962(.A(n_60969), .B(n_60958), .C(n_62850), .D(\nbus_11307[1] 
		), .Z(n_297766506));
	notech_or4 i_28980(.A(n_60969), .B(n_60958), .C(n_62850), .D(n_29678), .Z
		(n_297666505));
	notech_or4 i_31628(.A(n_29652), .B(n_29658), .C(n_26770), .D(n_28545), .Z
		(n_297566504));
	notech_or4 i_31649(.A(n_56834), .B(n_32382), .C(n_61142), .D(n_27036), .Z
		(n_297466503));
	notech_nand2 i_52940756(.A(opb[8]), .B(n_292666455), .Z(n_295366482));
	notech_nand2 i_53240753(.A(sav_edi[8]), .B(n_61142), .Z(n_295066479));
	notech_nand3 i_53540750(.A(n_6365), .B(n_29601), .C(n_1430), .Z(n_294766476
		));
	notech_or4 i_47440805(.A(n_32555), .B(n_61142), .C(n_60340), .D(n_28097)
		, .Z(n_294066469));
	notech_or2 i_48140798(.A(n_310191722), .B(n_27439), .Z(n_293366462));
	notech_and3 i_79340511(.A(n_28543), .B(n_28544), .C(n_301091813), .Z(n_292966458
		));
	notech_ao4 i_122541349(.A(n_61115), .B(n_30594), .C(n_300491819), .D(n_28545
		), .Z(n_292866457));
	notech_and2 i_122441348(.A(n_301891805), .B(n_102135817), .Z(n_292766456
		));
	notech_nand3 i_110041347(.A(n_299591828), .B(n_299991824), .C(n_300191822
		), .Z(n_292666455));
	notech_and3 i_109941346(.A(n_2993), .B(n_299791826), .C(n_303466563), .Z
		(n_292566454));
	notech_and3 i_64941345(.A(n_28502), .B(n_303366562), .C(n_303591788), .Z
		(n_292466453));
	notech_and2 i_122061801(.A(n_102135817), .B(n_312791696), .Z(n_292366452
		));
	notech_ao4 i_122161800(.A(n_61115), .B(n_30594), .C(n_26616), .D(n_319291631
		), .Z(n_292266451));
	notech_or4 i_140941256(.A(n_29652), .B(n_29658), .C(n_26770), .D(n_292966458
		), .Z(n_292166450));
	notech_and4 i_147643101(.A(n_291866447), .B(n_291766446), .C(n_291566444
		), .D(n_291466443), .Z(n_292066449));
	notech_ao4 i_146843107(.A(n_310191722), .B(n_27432), .C(n_146328740), .D
		(n_28598), .Z(n_291866447));
	notech_ao4 i_146943106(.A(n_146228739), .B(n_29856), .C(n_60020), .D(n_58000
		), .Z(n_291766446));
	notech_ao4 i_147143104(.A(n_57999), .B(n_29651), .C(n_58367), .D(n_27987
		), .Z(n_291566444));
	notech_ao4 i_147243103(.A(n_310291721), .B(n_28094), .C(n_60149), .D(n_27160
		), .Z(n_291466443));
	notech_and4 i_148743094(.A(n_291166440), .B(n_291066439), .C(n_290866437
		), .D(n_290766436), .Z(n_291366442));
	notech_ao4 i_147743100(.A(\nbus_11358[5] ), .B(n_57885), .C(\nbus_11307[5] 
		), .D(n_57886), .Z(n_291166440));
	notech_ao4 i_147843099(.A(n_308621250), .B(n_111564644), .C(n_26614), .D
		(n_282266351), .Z(n_291066439));
	notech_ao4 i_148043097(.A(n_282166350), .B(n_236065889), .C(n_282066349)
		, .D(n_111464643), .Z(n_290866437));
	notech_ao4 i_148343096(.A(n_281966348), .B(n_56512), .C(n_281866347), .D
		(n_281566344), .Z(n_290766436));
	notech_and4 i_149343089(.A(n_290466433), .B(n_290266431), .C(n_306121225
		), .D(n_272566254), .Z(n_290666435));
	notech_ao4 i_148943093(.A(n_310191722), .B(n_27434), .C(n_146328740), .D
		(n_28599), .Z(n_290466433));
	notech_ao4 i_149143091(.A(n_310291721), .B(n_28095), .C(n_60153), .D(n_27161
		), .Z(n_290266431));
	notech_and4 i_149843084(.A(n_289966428), .B(n_289566424), .C(n_272866257
		), .D(n_273166260), .Z(n_290166430));
	notech_ao4 i_149443088(.A(n_56619), .B(n_303221196), .C(n_26614), .D(n_267266201
		), .Z(n_289966428));
	notech_ao4 i_150043082(.A(n_317191652), .B(n_29723), .C(n_92519107), .D(n_17107
		), .Z(n_289766426));
	notech_ao4 i_149643086(.A(\nbus_11358[6] ), .B(n_267066199), .C(\nbus_11307[6] 
		), .D(n_266966198), .Z(n_289566424));
	notech_and4 i_150743077(.A(n_38618568), .B(n_289266421), .C(n_289066419)
		, .D(n_273966268), .Z(n_289466423));
	notech_ao4 i_150143081(.A(n_310191722), .B(n_27487), .C(n_146328740), .D
		(n_28624), .Z(n_289266421));
	notech_ao4 i_150443079(.A(n_310291721), .B(n_28123), .C(n_60153), .D(n_27188
		), .Z(n_289066419));
	notech_and4 i_151343071(.A(n_288766416), .B(n_288566414), .C(n_288466413
		), .D(n_274266271), .Z(n_288966418));
	notech_ao4 i_150843076(.A(n_314591678), .B(n_56619), .C(n_83019012), .D(n_267966208
		), .Z(n_288766416));
	notech_ao4 i_151043074(.A(n_314791676), .B(n_267866207), .C(n_267766206)
		, .D(\nbus_11358[31] ), .Z(n_288566414));
	notech_ao4 i_151143073(.A(n_29619), .B(n_267666205), .C(\nbus_11365[31] 
		), .D(n_288366412), .Z(n_288466413));
	notech_or2 i_151443070(.A(n_312191702), .B(n_312091703), .Z(n_288366412)
		);
	notech_and4 i_164042947(.A(n_274966278), .B(n_288066409), .C(n_287866407
		), .D(n_287766406), .Z(n_288266411));
	notech_ao4 i_163542952(.A(n_28530), .B(n_29857), .C(n_60022), .D(n_300091823
		), .Z(n_288066409));
	notech_ao4 i_163742950(.A(n_300291821), .B(n_29728), .C(n_268366212), .D
		(\nbus_11307[3] ), .Z(n_287866407));
	notech_ao4 i_163842949(.A(n_268266211), .B(\nbus_11358[3] ), .C(n_303291791
		), .D(n_27985), .Z(n_287766406));
	notech_and4 i_164742940(.A(n_287466403), .B(n_287366402), .C(n_287166400
		), .D(n_287066399), .Z(n_287666405));
	notech_ao4 i_164142946(.A(n_32270), .B(n_28092), .C(n_60153), .D(n_27219
		), .Z(n_287466403));
	notech_ao4 i_164242945(.A(n_308721251), .B(n_28502), .C(n_306970080), .D
		(n_28544), .Z(n_287366402));
	notech_ao4 i_164442943(.A(n_306870079), .B(n_28236), .C(n_306770078), .D
		(n_28234), .Z(n_287166400));
	notech_ao4 i_164542942(.A(n_306670077), .B(n_111664645), .C(n_306570076)
		, .D(n_303891785), .Z(n_287066399));
	notech_and4 i_165342934(.A(n_276466293), .B(n_286766396), .C(n_286566394
		), .D(n_286466393), .Z(n_286966398));
	notech_ao4 i_164842939(.A(n_28530), .B(n_29858), .C(n_300091823), .D(n_60020
		), .Z(n_286766396));
	notech_ao4 i_165042937(.A(n_300291821), .B(n_29651), .C(\nbus_11307[5] )
		, .D(n_268366212), .Z(n_286566394));
	notech_ao4 i_165142936(.A(n_268266211), .B(\nbus_11358[5] ), .C(n_303291791
		), .D(n_27987), .Z(n_286466393));
	notech_and4 i_166142927(.A(n_286166390), .B(n_286066389), .C(n_285866387
		), .D(n_285766386), .Z(n_286366392));
	notech_ao4 i_165442933(.A(n_59326), .B(n_28094), .C(n_60153), .D(n_27222
		), .Z(n_286166390));
	notech_ao4 i_165642932(.A(n_308621250), .B(n_28502), .C(n_282266351), .D
		(n_28544), .Z(n_286066389));
	notech_ao4 i_165842930(.A(n_28236), .B(n_282166350), .C(n_282066349), .D
		(n_28234), .Z(n_285866387));
	notech_ao4 i_165942929(.A(n_303891785), .B(n_281966348), .C(n_281866347)
		, .D(n_111664645), .Z(n_285766386));
	notech_and4 i_166542923(.A(n_308470095), .B(n_277766306), .C(n_285266381
		), .D(n_278066309), .Z(n_285666385));
	notech_ao4 i_167042918(.A(\nbus_11358[6] ), .B(n_27306), .C(n_3852), .D(\nbus_11307[6] 
		), .Z(n_285466383));
	notech_ao4 i_166342925(.A(n_60149), .B(n_27223), .C(n_92019102), .D(n_28236
		), .Z(n_285266381));
	notech_ao4 i_166642922(.A(n_92519107), .B(n_199965528), .C(n_56570), .D(n_303221196
		), .Z(n_285066379));
	notech_ao4 i_4244452(.A(n_32370), .B(n_27989), .C(n_3868), .D(n_32355), 
		.Z(n_284966378));
	notech_ao4 i_166742921(.A(n_268566214), .B(n_59349), .C(n_268466213), .D
		(n_284666375), .Z(n_284766376));
	notech_nand2 i_167242916(.A(n_59349), .B(n_26668), .Z(n_284666375));
	notech_ao4 i_167142917(.A(n_299891825), .B(\nbus_11307[6] ), .C(n_26802)
		, .D(n_26890), .Z(n_284566374));
	notech_and4 i_167642912(.A(n_284166370), .B(n_297680477), .C(n_279066319
		), .D(n_279366322), .Z(n_284466373));
	notech_ao4 i_167442914(.A(n_29619), .B(n_26700), .C(n_314791676), .D(n_104922313
		), .Z(n_284166370));
	notech_ao4 i_167742911(.A(n_60149), .B(n_27245), .C(n_83019012), .D(n_309691727
		), .Z(n_283966368));
	notech_ao4 i_167842910(.A(n_314591678), .B(n_56570), .C(n_301091813), .D
		(n_270066229), .Z(n_283766366));
	notech_ao4 i_205642534(.A(n_26924), .B(n_28228), .C(n_26922), .D(n_28195
		), .Z(n_283466363));
	notech_ao4 i_205742533(.A(n_56919), .B(n_29859), .C(n_26969), .D(n_28262
		), .Z(n_283366362));
	notech_and2 i_206142529(.A(n_283166360), .B(n_283066359), .Z(n_283266361
		));
	notech_ao4 i_205942531(.A(n_26927), .B(n_28294), .C(n_26920), .D(n_28360
		), .Z(n_283166360));
	notech_ao4 i_206042530(.A(n_26933), .B(n_28327), .C(n_56630), .D(n_28424
		), .Z(n_283066359));
	notech_and4 i_206942521(.A(n_282766356), .B(n_282666355), .C(n_282466353
		), .D(n_282366352), .Z(n_282966358));
	notech_ao4 i_206342527(.A(n_56619), .B(n_28392), .C(n_26928), .D(n_28456
		), .Z(n_282766356));
	notech_ao4 i_206442526(.A(n_26651), .B(n_28163), .C(n_26925), .D(n_28488
		), .Z(n_282666355));
	notech_ao4 i_206642524(.A(n_56570), .B(n_28521), .C(n_26721), .D(n_27863
		), .Z(n_282466353));
	notech_ao4 i_206742523(.A(n_56548), .B(n_28565), .C(n_26649), .D(n_29860
		), .Z(n_282366352));
	notech_or4 i_61544490(.A(n_60969), .B(n_60958), .C(n_62834), .D(n_29651)
		, .Z(n_282266351));
	notech_nand2 i_61844489(.A(opc_10[5]), .B(n_62794), .Z(n_282166350));
	notech_nand2 i_70244487(.A(opc[5]), .B(n_62794), .Z(n_282066349));
	notech_or4 i_70744485(.A(n_60969), .B(n_60958), .C(n_62850), .D(\nbus_11307[5] 
		), .Z(n_281966348));
	notech_nao3 i_71544482(.A(n_62776), .B(opa[5]), .C(n_62850), .Z(n_281866347
		));
	notech_nand2 i_217642414(.A(n_26613), .B(n_312191702), .Z(n_281666345)
		);
	notech_or2 i_10044394(.A(n_56512), .B(n_17107), .Z(n_281566344));
	notech_nand3 i_65443862(.A(n_309791726), .B(n_62790), .C(opc[31]), .Z(n_279866327
		));
	notech_nand3 i_65943857(.A(n_1430), .B(n_6412), .C(\eflags[10] ), .Z(n_279366322
		));
	notech_nand3 i_66043856(.A(n_1430), .B(n_6411), .C(n_29601), .Z(n_279066319
		));
	notech_ao4 i_63343883(.A(n_269066219), .B(n_26674), .C(n_28332), .D(n_26683
		), .Z(n_278566314));
	notech_nand3 i_63843878(.A(n_1430), .B(n_6362), .C(\eflags[10] ), .Z(n_278066309
		));
	notech_nand3 i_63943877(.A(n_1430), .B(n_6361), .C(n_29601), .Z(n_277766306
		));
	notech_nand3 i_63043886(.A(n_1430), .B(n_6359), .C(n_29601), .Z(n_276466293
		));
	notech_nand3 i_60943901(.A(n_1430), .B(n_6355), .C(n_29601), .Z(n_274966278
		));
	notech_or4 i_42544072(.A(n_312191702), .B(n_60942), .C(nbus_11295[31]), 
		.D(n_54929), .Z(n_274266271));
	notech_nand2 i_42844069(.A(n_7380), .B(n_26986), .Z(n_273966268));
	notech_or2 i_41844079(.A(n_3874), .B(n_26611), .Z(n_273266261));
	notech_nand3 i_40344093(.A(n_62776), .B(opc[6]), .C(n_267166200), .Z(n_273166260
		));
	notech_or4 i_40644090(.A(n_26614), .B(n_60942), .C(n_28131), .D(n_54929)
		, .Z(n_272866257));
	notech_nand2 i_40944087(.A(n_7355), .B(n_26986), .Z(n_272566254));
	notech_and3 i_10544390(.A(n_26613), .B(n_312191702), .C(n_26616), .Z(n_56512
		));
	notech_or2 i_125243310(.A(n_26611), .B(n_56512), .Z(n_270466233));
	notech_or2 i_125143311(.A(n_56512), .B(n_317191652), .Z(n_270366232));
	notech_ao4 i_13244364(.A(\nbus_11358[31] ), .B(n_26681), .C(n_299891825)
		, .D(\nbus_11365[31] ), .Z(n_270066229));
	notech_nand2 i_64943867(.A(n_304491779), .B(opd[6]), .Z(n_269766226));
	notech_ao4 i_64843868(.A(n_3874), .B(n_26602), .C(n_29723), .D(n_308891735
		), .Z(n_269466223));
	notech_or2 i_8944405(.A(n_26610), .B(n_269466223), .Z(n_269366222));
	notech_nand2 i_64743869(.A(n_285466383), .B(n_269366222), .Z(n_269266221
		));
	notech_or4 i_64543871(.A(n_60942), .B(n_60909), .C(n_29723), .D(n_28551)
		, .Z(n_269166220));
	notech_and2 i_64443872(.A(opb[6]), .B(n_28546), .Z(n_269066219));
	notech_nor2 i_232361787(.A(n_28332), .B(n_26683), .Z(n_268666215));
	notech_ao4 i_13344363(.A(n_305621220), .B(n_28544), .C(n_199965528), .D(n_310073580
		), .Z(n_268566214));
	notech_and2 i_8544409(.A(n_305721221), .B(n_269166220), .Z(n_268466213)
		);
	notech_and2 i_116661802(.A(n_298991830), .B(n_116264691), .Z(n_268366212
		));
	notech_ao4 i_116561803(.A(n_61115), .B(n_27306), .C(n_26681), .D(n_268666215
		), .Z(n_268266211));
	notech_nand2 i_43444063(.A(n_303491789), .B(n_17107), .Z(n_268166210));
	notech_and2 i_15244344(.A(n_344666975), .B(n_268166210), .Z(n_267966208)
		);
	notech_and2 i_15144345(.A(n_312691697), .B(n_267466203), .Z(n_267866207)
		);
	notech_ao4 i_15044346(.A(n_1895), .B(n_61115), .C(n_312191702), .D(n_26611
		), .Z(n_267766206));
	notech_and2 i_14944347(.A(n_312591698), .B(n_312891695), .Z(n_267666205)
		);
	notech_nand2 i_41444082(.A(n_281666345), .B(n_17107), .Z(n_267566204));
	notech_or2 i_41344083(.A(n_26611), .B(n_26616), .Z(n_267466203));
	notech_and3 i_15644340(.A(n_92619108), .B(n_289766426), .C(n_273266261),
		 .Z(n_267266201));
	notech_nand2 i_15544341(.A(n_344666975), .B(n_267566204), .Z(n_267166200
		));
	notech_and3 i_15444342(.A(n_312991694), .B(n_116164690), .C(n_267466203)
		, .Z(n_267066199));
	notech_and2 i_15344343(.A(n_344566974), .B(n_312891695), .Z(n_266966198)
		);
	notech_and4 i_138046364(.A(n_125828535), .B(n_266566194), .C(n_233965868
		), .D(n_26754), .Z(n_266866197));
	notech_ao4 i_137846366(.A(n_3845), .B(n_111164640), .C(n_3877), .D(\nbus_11358[21] 
		), .Z(n_266566194));
	notech_and4 i_138546359(.A(n_266266191), .B(n_266066189), .C(n_234265871
		), .D(n_234565874), .Z(n_266466193));
	notech_ao4 i_138146363(.A(n_26642), .B(n_29681), .C(n_3857), .D(n_28006)
		, .Z(n_266266191));
	notech_ao4 i_138346361(.A(n_263180132), .B(\nbus_11365[21] ), .C(n_3858)
		, .D(n_249866027), .Z(n_266066189));
	notech_and4 i_139146353(.A(n_265766186), .B(n_265566184), .C(n_265466183
		), .D(n_234865877), .Z(n_265966188));
	notech_ao4 i_138646358(.A(n_146328740), .B(n_28609), .C(n_146228739), .D
		(n_29842), .Z(n_265766186));
	notech_ao4 i_138846356(.A(n_310291721), .B(n_28105), .C(n_310391720), .D
		(n_28001), .Z(n_265566184));
	notech_ao4 i_138946355(.A(n_60149), .B(n_27171), .C(n_232565854), .D(\nbus_11365[16] 
		), .Z(n_265466183));
	notech_and4 i_139746347(.A(n_265166180), .B(n_264966178), .C(n_264866177
		), .D(n_235565884), .Z(n_265366182));
	notech_ao4 i_139246352(.A(n_147128748), .B(n_29710), .C(n_147028747), .D
		(\nbus_11358[16] ), .Z(n_265166180));
	notech_ao4 i_139446350(.A(n_313747721), .B(n_146428741), .C(n_312191702)
		, .D(n_312324377), .Z(n_264966178));
	notech_ao4 i_139546349(.A(n_252966058), .B(n_310491719), .C(n_254466073)
		, .D(n_232465853), .Z(n_264866177));
	notech_and4 i_140446340(.A(n_264466173), .B(n_264266171), .C(n_264166170
		), .D(n_236465893), .Z(n_264666175));
	notech_ao4 i_139946345(.A(n_146328740), .B(n_28610), .C(n_146228739), .D
		(n_29843), .Z(n_264466173));
	notech_ao4 i_140146343(.A(n_310291721), .B(n_28106), .C(n_310391720), .D
		(n_28002), .Z(n_264266171));
	notech_ao4 i_140246342(.A(n_60149), .B(n_27172), .C(n_232565854), .D(\nbus_11365[17] 
		), .Z(n_264166170));
	notech_and4 i_141046334(.A(n_263866167), .B(n_263666165), .C(n_263566164
		), .D(n_237165900), .Z(n_264066169));
	notech_ao4 i_140546339(.A(n_147128748), .B(n_29772), .C(n_147028747), .D
		(\nbus_11358[17] ), .Z(n_263866167));
	notech_ao4 i_140746337(.A(n_313647722), .B(n_146428741), .C(n_249672976)
		, .D(n_301791806), .Z(n_263666165));
	notech_ao4 i_140846336(.A(n_254673026), .B(n_312191702), .C(n_245572935)
		, .D(n_310491719), .Z(n_263566164));
	notech_and4 i_141646328(.A(n_263266161), .B(n_263066159), .C(n_262966158
		), .D(n_237865907), .Z(n_263466163));
	notech_ao4 i_141146333(.A(n_146328740), .B(n_28611), .C(n_146228739), .D
		(n_29844), .Z(n_263266161));
	notech_ao4 i_141346331(.A(n_310291721), .B(n_28107), .C(n_310391720), .D
		(n_28003), .Z(n_263066159));
	notech_ao4 i_141446330(.A(n_60149), .B(n_27173), .C(n_232565854), .D(\nbus_11365[18] 
		), .Z(n_262966158));
	notech_and4 i_142246322(.A(n_262666155), .B(n_262466153), .C(n_262366152
		), .D(n_238565914), .Z(n_262866157));
	notech_ao4 i_141746327(.A(n_147128748), .B(n_29711), .C(n_147028747), .D
		(\nbus_11358[18] ), .Z(n_262666155));
	notech_ao4 i_141946325(.A(n_3861), .B(n_146428741), .C(n_77522039), .D(n_301791806
		), .Z(n_262466153));
	notech_ao4 i_142046324(.A(n_60121865), .B(n_312191702), .C(n_95222216), 
		.D(n_310491719), .Z(n_262366152));
	notech_and4 i_142846316(.A(n_262066149), .B(n_261866147), .C(n_261766146
		), .D(n_239265921), .Z(n_262266151));
	notech_ao4 i_142346321(.A(n_146328740), .B(n_28612), .C(n_146228739), .D
		(n_29845), .Z(n_262066149));
	notech_ao4 i_142546319(.A(n_310291721), .B(n_28108), .C(n_310391720), .D
		(n_28004), .Z(n_261866147));
	notech_ao4 i_142646318(.A(n_60149), .B(n_27175), .C(n_232565854), .D(\nbus_11365[19] 
		), .Z(n_261766146));
	notech_and4 i_143446310(.A(n_261466143), .B(n_261266141), .C(n_261166140
		), .D(n_239965928), .Z(n_261666145));
	notech_ao4 i_142946315(.A(n_147128748), .B(n_29773), .C(n_147028747), .D
		(\nbus_11358[19] ), .Z(n_261466143));
	notech_ao4 i_143146313(.A(n_313447724), .B(n_146428741), .C(n_247972959)
		, .D(n_301791806), .Z(n_261266141));
	notech_ao4 i_143246312(.A(n_253773017), .B(n_312191702), .C(n_243072910)
		, .D(n_310491719), .Z(n_261166140));
	notech_and4 i_144546305(.A(n_260866137), .B(n_260666135), .C(n_240665935
		), .D(n_240965938), .Z(n_261066139));
	notech_ao4 i_143546309(.A(n_146328740), .B(n_28613), .C(n_146228739), .D
		(n_29846), .Z(n_260866137));
	notech_ao4 i_143746307(.A(n_310291721), .B(n_28109), .C(n_310391720), .D
		(n_28005), .Z(n_260666135));
	notech_and4 i_145146299(.A(n_260366132), .B(n_260166130), .C(n_260066129
		), .D(n_241265941), .Z(n_260566134));
	notech_ao4 i_144646304(.A(n_60005), .B(n_147228749), .C(n_29775), .D(n_147128748
		), .Z(n_260366132));
	notech_ao4 i_144846302(.A(\nbus_11358[20] ), .B(n_147028747), .C(n_313347725
		), .D(n_146428741), .Z(n_260166130));
	notech_ao4 i_144946301(.A(n_247072950), .B(n_301791806), .C(n_241572895)
		, .D(n_310491719), .Z(n_260066129));
	notech_and4 i_159446161(.A(n_259766126), .B(n_259566124), .C(n_241965948
		), .D(n_242265951), .Z(n_259966128));
	notech_ao4 i_159046165(.A(n_28530), .B(n_29847), .C(n_32270), .D(n_28105
		), .Z(n_259766126));
	notech_ao4 i_159246163(.A(n_60149), .B(n_27232), .C(n_254466073), .D(n_309691727
		), .Z(n_259566124));
	notech_ao4 i_159546160(.A(n_252966058), .B(n_26678), .C(n_301091813), .D
		(n_232865857), .Z(n_259266121));
	notech_ao4 i_160146155(.A(n_300491819), .B(\nbus_11365[16] ), .C(\nbus_11358[16] 
		), .D(n_26681), .Z(n_259166120));
	notech_ao3 i_159946157(.A(n_242665955), .B(n_242865957), .C(n_242765956)
		, .Z(n_259066119));
	notech_and4 i_160846149(.A(n_258566114), .B(n_258366112), .C(n_243365962
		), .D(n_243665965), .Z(n_258766116));
	notech_ao4 i_160446153(.A(n_28530), .B(n_29848), .C(n_32270), .D(n_28106
		), .Z(n_258566114));
	notech_ao4 i_160646151(.A(n_60149), .B(n_27234), .C(n_233165860), .D(\nbus_11365[17] 
		), .Z(n_258366112));
	notech_and4 i_161446143(.A(n_258066109), .B(n_257866107), .C(n_257766106
		), .D(n_243965968), .Z(n_258266111));
	notech_ao4 i_160946148(.A(n_140328680), .B(n_29772), .C(n_140228679), .D
		(\nbus_11358[17] ), .Z(n_258066109));
	notech_ao4 i_161146146(.A(n_313647722), .B(n_139728674), .C(n_254673026)
		, .D(n_301091813), .Z(n_257866107));
	notech_ao4 i_161246145(.A(n_249672976), .B(n_309691727), .C(n_245572935)
		, .D(n_26678), .Z(n_257766106));
	notech_and4 i_162046138(.A(n_257466103), .B(n_257266101), .C(n_244665975
		), .D(n_244965978), .Z(n_257666105));
	notech_ao4 i_161646142(.A(n_28530), .B(n_29849), .C(n_32270), .D(n_28107
		), .Z(n_257466103));
	notech_ao4 i_161846140(.A(n_60153), .B(n_27235), .C(n_233165860), .D(\nbus_11365[18] 
		), .Z(n_257266101));
	notech_and4 i_162646132(.A(n_256966098), .B(n_256766096), .C(n_256666095
		), .D(n_245265981), .Z(n_257166100));
	notech_ao4 i_162146137(.A(n_140328680), .B(n_29711), .C(n_140228679), .D
		(\nbus_11358[18] ), .Z(n_256966098));
	notech_ao4 i_162346135(.A(n_3861), .B(n_139728674), .C(n_60121865), .D(n_301091813
		), .Z(n_256766096));
	notech_ao4 i_162446134(.A(n_77522039), .B(n_309691727), .C(n_95222216), 
		.D(n_26678), .Z(n_256666095));
	notech_and4 i_163146127(.A(n_256366092), .B(n_256166090), .C(n_245965988
		), .D(n_246265991), .Z(n_256566094));
	notech_ao4 i_162746131(.A(n_28530), .B(n_29850), .C(n_59326), .D(n_28108
		), .Z(n_256366092));
	notech_ao4 i_162946129(.A(n_60157), .B(n_27236), .C(n_233165860), .D(\nbus_11365[19] 
		), .Z(n_256166090));
	notech_and4 i_163746121(.A(n_255866087), .B(n_255666085), .C(n_255566084
		), .D(n_246565994), .Z(n_256066089));
	notech_ao4 i_163246126(.A(n_140328680), .B(n_29773), .C(n_140228679), .D
		(\nbus_11358[19] ), .Z(n_255866087));
	notech_ao4 i_163446124(.A(n_313447724), .B(n_139728674), .C(n_253773017)
		, .D(n_301091813), .Z(n_255666085));
	notech_ao4 i_163546123(.A(n_247972959), .B(n_309691727), .C(n_243072910)
		, .D(n_26678), .Z(n_255566084));
	notech_and4 i_164246116(.A(n_255266081), .B(n_255066079), .C(n_247266001
		), .D(n_247566004), .Z(n_255466083));
	notech_ao4 i_163846120(.A(n_28530), .B(n_29851), .C(n_59326), .D(n_28109
		), .Z(n_255266081));
	notech_ao4 i_164046118(.A(n_60157), .B(n_27237), .C(n_60005), .D(n_140428681
		), .Z(n_255066079));
	notech_and4 i_164746111(.A(n_254766076), .B(n_254566074), .C(n_247866007
		), .D(n_248166010), .Z(n_254966078));
	notech_ao4 i_164346115(.A(n_140228679), .B(\nbus_11358[20] ), .C(n_140128678
		), .D(\nbus_11365[20] ), .Z(n_254766076));
	notech_ao4 i_164546113(.A(n_247072950), .B(n_309691727), .C(n_241572895)
		, .D(n_26678), .Z(n_254566074));
	notech_nand2 i_1547706(.A(opc_10[16]), .B(n_62816), .Z(n_254466073));
	notech_ao4 i_200245780(.A(n_28241), .B(n_26924), .C(n_28206), .D(n_26922
		), .Z(n_254166070));
	notech_ao4 i_200345779(.A(n_56919), .B(n_29852), .C(n_28273), .D(n_26969
		), .Z(n_254066069));
	notech_and2 i_200745775(.A(n_253866067), .B(n_253766066), .Z(n_253966068
		));
	notech_ao4 i_200545777(.A(n_28306), .B(n_26927), .C(n_26649), .D(n_29853
		), .Z(n_253866067));
	notech_ao4 i_200645776(.A(n_26920), .B(n_28371), .C(n_26933), .D(n_28339
		), .Z(n_253766066));
	notech_and4 i_201545767(.A(n_253466063), .B(n_253366062), .C(n_253166060
		), .D(n_253066059), .Z(n_253666065));
	notech_ao4 i_200945773(.A(n_28435), .B(n_56630), .C(n_56619), .D(n_28403
		), .Z(n_253466063));
	notech_ao4 i_201045772(.A(n_26928), .B(n_28467), .C(n_26651), .D(n_28174
		), .Z(n_253366062));
	notech_ao4 i_201245770(.A(n_28499), .B(n_26925), .C(n_56557), .D(n_27874
		), .Z(n_253166060));
	notech_ao4 i_201345769(.A(n_56548), .B(n_28577), .C(n_56570), .D(n_28537
		), .Z(n_253066059));
	notech_nand2 i_29247699(.A(opc[16]), .B(n_62816), .Z(n_252966058));
	notech_ao4 i_213745646(.A(n_28246), .B(n_56666), .C(n_28211), .D(n_56653
		), .Z(n_252666055));
	notech_ao4 i_213845645(.A(n_56919), .B(n_29854), .C(n_28278), .D(n_56640
		), .Z(n_252566054));
	notech_and2 i_214245641(.A(n_252366052), .B(n_252266051), .Z(n_252466053
		));
	notech_ao4 i_214045643(.A(n_28311), .B(n_56532), .C(n_56518), .D(n_29855
		), .Z(n_252366052));
	notech_ao4 i_214145642(.A(n_56502), .B(n_28376), .C(n_56489), .D(n_28344
		), .Z(n_252266051));
	notech_and4 i_215045633(.A(n_251966048), .B(n_251866047), .C(n_251666045
		), .D(n_251566044), .Z(n_252166050));
	notech_ao4 i_214445639(.A(n_28440), .B(n_56630), .C(n_56619), .D(n_28408
		), .Z(n_251966048));
	notech_ao4 i_214545638(.A(n_56605), .B(n_28472), .C(n_28505), .D(n_56583
		), .Z(n_251866047));
	notech_ao4 i_214745636(.A(n_56557), .B(n_27882), .C(n_56547), .D(n_28582
		), .Z(n_251666045));
	notech_ao4 i_214845635(.A(n_26651), .B(n_28179), .C(n_56570), .D(n_28547
		), .Z(n_251566044));
	notech_nand2 i_6947630(.A(opc[21]), .B(n_62816), .Z(n_249866027));
	notech_or2 i_62247097(.A(n_313347725), .B(n_139728674), .Z(n_248166010)
		);
	notech_or2 i_62547094(.A(n_140328680), .B(n_29775), .Z(n_247866007));
	notech_or4 i_62847091(.A(n_56689), .B(n_56570), .C(n_61142), .D(n_28005)
		, .Z(n_247566004));
	notech_nand3 i_63147088(.A(n_1430), .B(n_6389), .C(n_29601), .Z(n_247266001
		));
	notech_or2 i_61347106(.A(n_60006), .B(n_140428681), .Z(n_246565994));
	notech_or4 i_61647103(.A(n_56688), .B(n_56570), .C(n_61142), .D(n_28004)
		, .Z(n_246265991));
	notech_nand3 i_61947100(.A(n_1430), .B(n_6387), .C(n_29601), .Z(n_245965988
		));
	notech_or2 i_60047119(.A(n_3864), .B(n_140428681), .Z(n_245265981));
	notech_or4 i_60347116(.A(n_56689), .B(n_27036), .C(n_61142), .D(n_28003)
		, .Z(n_244965978));
	notech_nand3 i_60647113(.A(n_1430), .B(n_6385), .C(n_29601), .Z(n_244665975
		));
	notech_or2 i_58647132(.A(n_60008), .B(n_140428681), .Z(n_243965968));
	notech_or4 i_58947129(.A(n_56689), .B(n_27036), .C(n_61142), .D(n_28002)
		, .Z(n_243665965));
	notech_nand3 i_59247126(.A(n_1430), .B(n_6383), .C(n_29601), .Z(n_243365962
		));
	notech_nand2 i_56647152(.A(\regs_13_14[16] ), .B(n_232765856), .Z(n_242865957
		));
	notech_nor2 i_56547153(.A(n_60009), .B(n_232665855), .Z(n_242765956));
	notech_or4 i_56447154(.A(n_2479), .B(n_313747721), .C(n_246791942), .D(n_314091683
		), .Z(n_242665955));
	notech_nao3 i_56947149(.A(n_60157), .B(n_60340), .C(n_307624340), .Z(n_242565954
		));
	notech_or4 i_57247146(.A(n_56689), .B(n_27036), .C(n_61143), .D(n_28001)
		, .Z(n_242265951));
	notech_nand3 i_57547143(.A(n_1430), .B(n_6381), .C(n_29601), .Z(n_241965948
		));
	notech_nand2 i_38747322(.A(sav_esp[20]), .B(n_61142), .Z(n_241265941));
	notech_or2 i_39047319(.A(n_146928746), .B(\nbus_11365[20] ), .Z(n_240965938
		));
	notech_or2 i_39347316(.A(n_310191722), .B(n_27463), .Z(n_240665935));
	notech_or2 i_37247336(.A(n_60006), .B(n_147228749), .Z(n_239965928));
	notech_ao4 i_131468548(.A(n_326990767), .B(n_60013), .C(n_56390), .D(n_27447
		), .Z(n_113268149));
	notech_ao4 i_131368549(.A(n_326790765), .B(n_27741), .C(n_326890766), .D
		(n_27780), .Z(n_113368150));
	notech_ao4 i_129068572(.A(n_326990767), .B(n_60000), .C(n_56390), .D(n_27475
		), .Z(n_113468151));
	notech_ao4 i_128968573(.A(n_326790765), .B(n_27758), .C(n_326890766), .D
		(n_27797), .Z(n_113568152));
	notech_nao3 i_10367299(.A(n_60157), .B(n_60340), .C(n_113768154), .Z(n_113668153
		));
	notech_ao4 i_5867343(.A(n_26702), .B(n_3911), .C(n_343570446), .D(n_343770448
		), .Z(n_113768154));
	notech_and4 i_56144(.A(n_343370444), .B(n_114368160), .C(n_114168158), .D
		(n_113668153), .Z(\nbus_11376[9] ));
	notech_nand3 i_56139(.A(n_114568162), .B(n_114368160), .C(n_221669228), 
		.Z(\nbus_11376[0] ));
	notech_ao4 i_10567297(.A(n_280634762), .B(n_3916), .C(n_27509), .D(n_32263
		), .Z(n_114168158));
	notech_ao4 i_28664455(.A(n_251540533), .B(n_116368180), .C(n_61115), .D(n_3603
		), .Z(n_114368160));
	notech_or2 i_47896(.A(n_252140539), .B(n_117368190), .Z(n_114468161));
	notech_nao3 i_9664357(.A(n_60157), .B(n_60338), .C(n_3917), .Z(n_114568162
		));
	notech_or4 i_9864355(.A(n_61115), .B(n_2839), .C(n_2888), .D(n_59434), .Z
		(n_114668163));
	notech_ao4 i_14764307(.A(n_32384), .B(n_26782), .C(n_27903), .D(n_27906)
		, .Z(n_114768164));
	notech_or4 i_98063497(.A(n_32446), .B(n_57772), .C(n_61143), .D(n_60241)
		, .Z(n_115268169));
	notech_or4 i_98663491(.A(calc_sz[1]), .B(n_246691943), .C(n_61115), .D(n_32446
		), .Z(n_115568172));
	notech_nand3 i_98963489(.A(n_60157), .B(n_60338), .C(n_115768174), .Z(n_115668173
		));
	notech_nand3 i_14064314(.A(n_32656), .B(n_1869), .C(n_115868175), .Z(n_115768174
		));
	notech_nand2 i_99063488(.A(n_252140539), .B(n_1891), .Z(n_115868175));
	notech_nand3 i_88963587(.A(n_114768164), .B(n_60157), .C(n_60340), .Z(n_116068177
		));
	notech_or4 i_97763500(.A(n_57823), .B(n_116468181), .C(n_61143), .D(n_60241
		), .Z(n_116168178));
	notech_or4 i_97863499(.A(n_56939), .B(n_61115), .C(n_116468181), .D(n_26782
		), .Z(n_116268179));
	notech_or4 i_12464330(.A(n_32581), .B(n_26900), .C(n_61142), .D(n_60338)
		, .Z(n_116368180));
	notech_or4 i_32472(.A(n_27125), .B(n_27580), .C(n_2869), .D(n_59434), .Z
		(n_116468181));
	notech_or4 i_172862775(.A(n_27988), .B(n_60868), .C(n_61142), .D(n_60241
		), .Z(n_116568182));
	notech_and2 i_6464389(.A(n_114568162), .B(n_115268169), .Z(n_116968186)
		);
	notech_nand3 i_162362878(.A(n_1891), .B(n_60157), .C(n_60340), .Z(n_117368190
		));
	notech_ao4 i_9464359(.A(n_27917), .B(n_125461537), .C(n_252140539), .D(n_117368190
		), .Z(n_117468191));
	notech_nao3 i_68661767(.A(n_138768404), .B(n_138968406), .C(n_138568402)
		, .Z(n_117868195));
	notech_or2 i_152361748(.A(n_297369985), .B(n_27353), .Z(n_117968196));
	notech_ao4 i_132961752(.A(n_306291761), .B(n_32382), .C(n_27761), .D(n_306991754
		), .Z(n_118068197));
	notech_or2 i_121760574(.A(n_118468201), .B(n_1393), .Z(n_118268199));
	notech_and3 i_260261724(.A(n_27346), .B(n_303791786), .C(n_27349), .Z(n_118468201
		));
	notech_nao3 i_6361665(.A(tsc[14]), .B(n_27855), .C(n_24989), .Z(n_118668203
		));
	notech_or4 i_6261666(.A(n_28140), .B(n_60942), .C(n_26942), .D(n_23512),
		 .Z(n_118968206));
	notech_nand2 i_5961669(.A(n_58097), .B(opb[14]), .Z(n_119268209));
	notech_nao3 i_5461674(.A(n_26941), .B(\opa_12[14] ), .C(n_316191662), .Z
		(n_119368210));
	notech_nao3 i_5561673(.A(n_318791636), .B(n_246991940), .C(n_139068407),
		 .Z(n_119468211));
	notech_nao3 i_5661672(.A(opc[14]), .B(n_62816), .C(n_312970140), .Z(n_119568212
		));
	notech_nao3 i_25561473(.A(tsc[45]), .B(n_27855), .C(n_24989), .Z(n_119668213
		));
	notech_or4 i_25461474(.A(n_62844), .B(n_183768854), .C(n_60942), .D(n_29592
		), .Z(n_119968216));
	notech_or4 i_25161477(.A(n_62844), .B(n_62816), .C(n_29592), .D(n_25010)
		, .Z(n_120268219));
	notech_ao3 i_26661462(.A(tsc[46]), .B(n_27855), .C(n_24989), .Z(n_120768224
		));
	notech_or4 i_26561463(.A(n_62844), .B(n_183768854), .C(n_60942), .D(n_29680
		), .Z(n_121068227));
	notech_or4 i_26261466(.A(n_62844), .B(n_62816), .C(n_29680), .D(n_25010)
		, .Z(n_121368230));
	notech_nao3 i_30561423(.A(n_26767), .B(n_26669), .C(n_298366512), .Z(n_121868235
		));
	notech_or4 i_30461424(.A(n_26062), .B(n_298266511), .C(n_27119), .D(n_26054
		), .Z(n_122168238));
	notech_or2 i_30161427(.A(n_302291801), .B(\nbus_11358[14] ), .Z(n_122468241
		));
	notech_or4 i_29861430(.A(n_3854), .B(n_26054), .C(n_32335), .D(n_29680),
		 .Z(n_122768244));
	notech_or4 i_48761243(.A(n_30854), .B(n_298266511), .C(n_26770), .D(n_58482
		), .Z(n_122868245));
	notech_nand2 i_48661244(.A(n_58378), .B(opd[14]), .Z(n_123168248));
	notech_nand2 i_48361247(.A(n_58055), .B(opa[14]), .Z(n_123468251));
	notech_or4 i_47961250(.A(n_58184), .B(n_58482), .C(n_60011), .D(n_56371)
		, .Z(n_123768254));
	notech_nand3 i_52161210(.A(n_1429), .B(n_7284), .C(\eflags[10] ), .Z(n_124068257
		));
	notech_nand3 i_53661195(.A(n_1429), .B(n_7290), .C(\eflags[10] ), .Z(n_125568272
		));
	notech_or4 i_59161148(.A(n_32348), .B(n_56547), .C(n_59965), .D(n_61142)
		, .Z(n_127268289));
	notech_or2 i_58761151(.A(n_302591798), .B(n_27997), .Z(n_127568292));
	notech_nand2 i_60161139(.A(n_27289), .B(opb[13]), .Z(n_128868305));
	notech_nand2 i_67561075(.A(opd[13]), .B(n_26640), .Z(n_129768314));
	notech_nand2 i_67261078(.A(opa[13]), .B(n_313870149), .Z(n_130068317));
	notech_nao3 i_66961081(.A(n_62820), .B(opc[13]), .C(n_4009), .Z(n_130368320
		));
	notech_nand2 i_68861064(.A(n_26640), .B(opd[14]), .Z(n_130868325));
	notech_nand2 i_68461067(.A(n_313870149), .B(opa[14]), .Z(n_131168328));
	notech_nao3 i_68161070(.A(opc[14]), .B(n_62816), .C(n_4009), .Z(n_131468331
		));
	notech_or2 i_71461038(.A(n_142828705), .B(\nbus_11358[30] ), .Z(n_132368340
		));
	notech_or4 i_89460864(.A(n_62844), .B(n_62816), .C(n_29680), .D(n_58481)
		, .Z(n_132468341));
	notech_nand2 i_89360865(.A(n_58377), .B(opd[14]), .Z(n_132768344));
	notech_or4 i_89060868(.A(n_58810), .B(n_58481), .C(n_28140), .D(n_60940)
		, .Z(n_133068347));
	notech_nao3 i_88660871(.A(n_58810), .B(n_26821), .C(n_298366512), .Z(n_133368350
		));
	notech_or2 i_94260818(.A(n_154331958), .B(nbus_11295[14]), .Z(n_133868355
		));
	notech_nand2 i_93960821(.A(n_58050), .B(opb[14]), .Z(n_134168358));
	notech_or4 i_93660824(.A(n_58477), .B(n_58132), .C(n_32325), .D(n_29680)
		, .Z(n_134468361));
	notech_or4 i_103460730(.A(n_62844), .B(n_184468861), .C(n_60940), .D(n_29680
		), .Z(n_134568362));
	notech_or4 i_103360731(.A(n_58805), .B(n_28140), .C(n_60940), .D(n_58478
		), .Z(n_134868365));
	notech_or2 i_103060734(.A(n_57181), .B(\nbus_11358[14] ), .Z(n_135168368
		));
	notech_or4 i_102760737(.A(n_58099), .B(n_58478), .C(n_32331), .D(n_29680
		), .Z(n_135468371));
	notech_or4 i_109760684(.A(n_58817), .B(n_58495), .C(n_60940), .D(nbus_11295
		[14]), .Z(n_135968376));
	notech_nand2 i_109460687(.A(n_57179), .B(opb[14]), .Z(n_136268379));
	notech_or4 i_109160690(.A(n_58100), .B(n_58479), .C(n_32332), .D(n_29680
		), .Z(n_136568382));
	notech_or4 i_115660631(.A(n_62844), .B(n_184768864), .C(n_60940), .D(n_29680
		), .Z(n_136668383));
	notech_nao3 i_115560632(.A(opc_10[14]), .B(n_62816), .C(n_57473), .Z(n_136968386
		));
	notech_or4 i_115160635(.A(n_62844), .B(n_58480), .C(n_62792), .D(n_29680
		), .Z(n_137268389));
	notech_or4 i_114860638(.A(n_58087), .B(n_58480), .C(n_60011), .D(n_56457
		), .Z(n_137568392));
	notech_or2 i_115960628(.A(n_30565), .B(n_60011), .Z(n_138068397));
	notech_nand2 i_31193(.A(n_26921), .B(n_26813), .Z(n_138168398));
	notech_ao3 i_120760584(.A(n_60340), .B(opb[30]), .C(n_30822), .Z(n_138568402
		));
	notech_ao4 i_224759591(.A(n_30803), .B(n_302991794), .C(n_309491729), .D
		(\nbus_11365[30] ), .Z(n_138768404));
	notech_ao4 i_224659592(.A(n_60340), .B(n_28121), .C(n_309591728), .D(n_29591
		), .Z(n_138968406));
	notech_or4 i_65661772(.A(calc_sz[1]), .B(n_246691943), .C(n_56834), .D(n_59963
		), .Z(n_139068407));
	notech_ao4 i_221159627(.A(n_184868865), .B(n_29680), .C(n_56640), .D(n_139068407
		), .Z(n_139168408));
	notech_ao4 i_220959629(.A(n_57807), .B(\nbus_11358[14] ), .C(n_57809), .D
		(\nbus_11307[14] ), .Z(n_139368410));
	notech_and4 i_221359625(.A(n_139368410), .B(n_137568392), .C(n_139168408
		), .D(n_137268389), .Z(n_139568412));
	notech_ao4 i_220659632(.A(nbus_11295[14]), .B(n_26823), .C(n_58376), .D(n_27999
		), .Z(n_139668413));
	notech_ao4 i_221559623(.A(n_28103), .B(n_60340), .C(n_30570), .D(n_29680
		), .Z(n_139868415));
	notech_ao4 i_221459624(.A(n_30569), .B(\nbus_11358[14] ), .C(n_30568), .D
		(\nbus_11307[14] ), .Z(n_140068417));
	notech_and3 i_66461769(.A(n_139868415), .B(n_140068417), .C(n_138068397)
		, .Z(n_140168418));
	notech_and4 i_220859630(.A(n_140168418), .B(n_136968386), .C(n_139668413
		), .D(n_136668383), .Z(n_140368420));
	notech_ao4 i_216759671(.A(n_323080731), .B(n_157165100), .C(n_56666), .D
		(n_139068407), .Z(n_140468421));
	notech_ao4 i_216559673(.A(n_26856), .B(\nbus_11307[14] ), .C(n_228579786
		), .D(n_60011), .Z(n_140668423));
	notech_and4 i_216959669(.A(n_140668423), .B(n_140468421), .C(n_136268379
		), .D(n_136568382), .Z(n_140868425));
	notech_ao4 i_216259676(.A(n_58375), .B(n_27999), .C(n_58479), .D(n_298166510
		), .Z(n_140968426));
	notech_ao4 i_216059678(.A(n_298366512), .B(n_228779788), .C(n_322780728)
		, .D(n_298266511), .Z(n_141168428));
	notech_and4 i_216459674(.A(n_140168418), .B(n_141168428), .C(n_140968426
		), .D(n_135968376), .Z(n_141368430));
	notech_ao4 i_212459714(.A(n_157165100), .B(n_313270143), .C(n_56653), .D
		(n_139068407), .Z(n_141468431));
	notech_ao4 i_212259716(.A(\nbus_11307[14] ), .B(n_26607), .C(n_60011), .D
		(n_184368860), .Z(n_141668433));
	notech_and4 i_212659712(.A(n_141668433), .B(n_141468431), .C(n_135168368
		), .D(n_135468371), .Z(n_141868435));
	notech_ao4 i_211959719(.A(n_58374), .B(n_27999), .C(n_58478), .D(n_298166510
		), .Z(n_141968436));
	notech_and4 i_212159717(.A(n_140168418), .B(n_141968436), .C(n_134568362
		), .D(n_134868365), .Z(n_142268439));
	notech_ao4 i_204759791(.A(n_58041), .B(n_157165100), .C(n_56919), .D(n_139068407
		), .Z(n_142368440));
	notech_ao4 i_204459793(.A(\nbus_11307[14] ), .B(n_26854), .C(n_228479785
		), .D(n_60011), .Z(n_142568442));
	notech_and4 i_204959789(.A(n_142568442), .B(n_142368440), .C(n_134168358
		), .D(n_134468361), .Z(n_142768444));
	notech_ao4 i_204159796(.A(n_58372), .B(n_27999), .C(n_58477), .D(n_298166510
		), .Z(n_142868445));
	notech_ao4 i_203859798(.A(n_228379784), .B(n_298366512), .C(n_322580726)
		, .D(n_298266511), .Z(n_143068447));
	notech_and4 i_204359794(.A(n_140168418), .B(n_143068447), .C(n_142868445
		), .D(n_133868355), .Z(n_143268449));
	notech_ao4 i_200259834(.A(n_181679320), .B(n_29680), .C(n_181779321), .D
		(n_60011), .Z(n_143368450));
	notech_ao4 i_200059836(.A(n_58038), .B(n_157165100), .C(n_56502), .D(n_139068407
		), .Z(n_143568452));
	notech_and4 i_200459832(.A(n_133068347), .B(n_143568452), .C(n_143368450
		), .D(n_133368350), .Z(n_143768454));
	notech_ao4 i_199759839(.A(n_26851), .B(\nbus_11307[14] ), .C(n_58052), .D
		(\nbus_11358[14] ), .Z(n_143868455));
	notech_and4 i_199959837(.A(n_140168418), .B(n_143868455), .C(n_132468341
		), .D(n_132768344), .Z(n_144168458));
	notech_ao4 i_185959969(.A(n_302991794), .B(n_143028707), .C(n_142728704)
		, .D(\nbus_11365[30] ), .Z(n_144268459));
	notech_ao4 i_185859970(.A(n_303091793), .B(n_309891725), .C(n_142928706)
		, .D(n_29591), .Z(n_144468461));
	notech_and3 i_186159967(.A(n_144268459), .B(n_144468461), .C(n_132368340
		), .Z(n_144568462));
	notech_ao4 i_185659972(.A(n_32252), .B(n_26595), .C(n_4014), .D(n_28015)
		, .Z(n_144668463));
	notech_ao4 i_185559973(.A(n_308091743), .B(n_28121), .C(n_30809), .D(n_295269964
		), .Z(n_144768464));
	notech_ao4 i_183459993(.A(n_56518), .B(n_139068407), .C(n_118068197), .D
		(n_56257), .Z(n_144968466));
	notech_ao4 i_183259995(.A(n_60011), .B(n_4007), .C(n_308091743), .D(n_28103
		), .Z(n_145168468));
	notech_and4 i_183659991(.A(n_145168468), .B(n_144968466), .C(n_131168328
		), .D(n_131468331), .Z(n_145368470));
	notech_ao4 i_182959998(.A(n_27761), .B(n_298166510), .C(n_4008), .D(\nbus_11358[14] 
		), .Z(n_145468471));
	notech_ao4 i_182859999(.A(n_27604), .B(n_298366512), .C(n_298266511), .D
		(n_307991744), .Z(n_145668473));
	notech_ao4 i_182560002(.A(n_56518), .B(n_94935745), .C(n_118068197), .D(n_29592
		), .Z(n_145868475));
	notech_ao4 i_182360004(.A(n_302091803), .B(n_4007), .C(n_308091743), .D(n_28102
		), .Z(n_146068477));
	notech_and4 i_182760000(.A(n_146068477), .B(n_145868475), .C(n_130068317
		), .D(n_130368320), .Z(n_146268479));
	notech_ao4 i_182060007(.A(n_27761), .B(n_31540), .C(n_4008), .D(\nbus_11358[13] 
		), .Z(n_146368480));
	notech_ao4 i_181960008(.A(n_27604), .B(n_31576), .C(n_31560), .D(n_307991744
		), .Z(n_146568482));
	notech_ao4 i_176860055(.A(n_52135317), .B(n_29592), .C(n_52335319), .D(n_302091803
		), .Z(n_146768484));
	notech_ao4 i_176760056(.A(n_60153), .B(n_27202), .C(n_30109), .D(n_27157
		), .Z(n_146868485));
	notech_ao4 i_176560058(.A(n_302691797), .B(\nbus_11307[13] ), .C(n_51735313
		), .D(n_31576), .Z(n_147068487));
	notech_and4 i_177060053(.A(n_147068487), .B(n_146868485), .C(n_146768484
		), .D(n_128868305), .Z(n_147268489));
	notech_ao4 i_176260061(.A(n_302591798), .B(n_27998), .C(n_27349), .D(n_31540
		), .Z(n_147368490));
	notech_ao4 i_176160062(.A(n_301691807), .B(n_27142), .C(n_27348), .D(n_31560
		), .Z(n_147468491));
	notech_ao4 i_175860064(.A(n_27334), .B(n_29876), .C(n_27335), .D(n_29875
		), .Z(n_147668493));
	notech_and3 i_175960063(.A(n_111364642), .B(n_147668493), .C(n_114664675
		), .Z(n_147768494));
	notech_ao4 i_175560067(.A(n_27335), .B(n_29874), .C(n_60153), .D(n_27201
		), .Z(n_147968496));
	notech_ao4 i_175460068(.A(n_27157), .B(n_156768584), .C(n_27334), .D(n_29873
		), .Z(n_148068497));
	notech_ao4 i_175260070(.A(n_320070211), .B(n_27349), .C(n_27348), .D(n_320170212
		), .Z(n_148268499));
	notech_and4 i_175760065(.A(n_148268499), .B(n_148068497), .C(n_147968496
		), .D(n_127568292), .Z(n_148468501));
	notech_ao4 i_174860073(.A(\nbus_11358[12] ), .B(n_302791796), .C(n_302691797
		), .D(\nbus_11307[12] ), .Z(n_148568502));
	notech_ao4 i_174660075(.A(n_313770148), .B(n_29679), .C(n_60013), .D(n_313670147
		), .Z(n_148768504));
	notech_and4 i_175160071(.A(n_148768504), .B(n_148568502), .C(n_47649), .D
		(n_127268289), .Z(n_148968506));
	notech_ao4 i_170260110(.A(n_297569987), .B(\nbus_11307[4] ), .C(n_291663183
		), .D(n_117968196), .Z(n_149068507));
	notech_ao4 i_170060111(.A(n_58001), .B(n_29725), .C(n_297469986), .D(\nbus_11358[4] 
		), .Z(n_149168508));
	notech_ao4 i_169860113(.A(n_60153), .B(n_27191), .C(n_5743), .D(n_58002)
		, .Z(n_149368510));
	notech_ao4 i_169760114(.A(n_58383), .B(n_27986), .C(n_59326), .D(n_28093
		), .Z(n_149468511));
	notech_and4 i_170460108(.A(n_149468511), .B(n_149368510), .C(n_149168508
		), .D(n_149068507), .Z(n_149668513));
	notech_ao4 i_169460117(.A(n_291463181), .B(n_300891815), .C(n_5723), .D(n_303691787
		), .Z(n_149768514));
	notech_ao4 i_169360118(.A(n_291763184), .B(n_185068867), .C(n_291563182)
		, .D(n_297369985), .Z(n_149868515));
	notech_ao4 i_169160120(.A(n_27335), .B(n_29872), .C(n_291863185), .D(n_274369755
		), .Z(n_150068517));
	notech_and4 i_169660115(.A(n_150068517), .B(n_149868515), .C(n_149768514
		), .D(n_125568272), .Z(n_150268519));
	notech_ao4 i_168860123(.A(n_297569987), .B(\nbus_11307[1] ), .C(n_297866507
		), .D(n_117968196), .Z(n_150368520));
	notech_ao4 i_168760124(.A(n_58001), .B(n_29678), .C(n_297469986), .D(\nbus_11358[1] 
		), .Z(n_150468521));
	notech_ao4 i_168560126(.A(n_60153), .B(n_27189), .C(n_60024), .D(n_58002
		), .Z(n_150668523));
	notech_ao4 i_168460127(.A(n_58383), .B(n_27983), .C(n_59326), .D(n_28090
		), .Z(n_150768524));
	notech_and4 i_169060121(.A(n_150768524), .B(n_150668523), .C(n_150468521
		), .D(n_150368520), .Z(n_150968526));
	notech_ao4 i_168160130(.A(n_297666505), .B(n_300891815), .C(n_59992), .D
		(n_303691787), .Z(n_151068527));
	notech_ao4 i_168060131(.A(n_297966508), .B(n_185068867), .C(n_297369985)
		, .D(n_297766506), .Z(n_151168528));
	notech_ao4 i_167860133(.A(n_27335), .B(n_29871), .C(n_298066509), .D(n_274369755
		), .Z(n_151368530));
	notech_and4 i_168360128(.A(n_151368530), .B(n_151168528), .C(n_151068527
		), .D(n_124068257), .Z(n_151568532));
	notech_ao4 i_165960152(.A(n_298366512), .B(n_128371763), .C(n_128471764)
		, .D(n_56257), .Z(n_151668533));
	notech_ao4 i_165760154(.A(n_58040), .B(n_157165100), .C(n_56489), .D(n_139068407
		), .Z(n_151868535));
	notech_and4 i_166160150(.A(n_151868535), .B(n_123768254), .C(n_151668533
		), .D(n_123468251), .Z(n_152068537));
	notech_ao4 i_165460157(.A(n_58482), .B(n_298166510), .C(n_58054), .D(\nbus_11358[14] 
		), .Z(n_152168538));
	notech_and4 i_165660155(.A(n_140168418), .B(n_122868245), .C(n_152168538
		), .D(n_123168248), .Z(n_152468541));
	notech_ao4 i_149060313(.A(n_301991804), .B(n_157165100), .C(n_56605), .D
		(n_139068407), .Z(n_152568542));
	notech_ao4 i_148860315(.A(\nbus_11307[14] ), .B(n_27293), .C(n_25875), .D
		(n_60011), .Z(n_152768544));
	notech_and4 i_149260311(.A(n_152768544), .B(n_152568542), .C(n_122468241
		), .D(n_122768244), .Z(n_152968546));
	notech_ao4 i_148560318(.A(n_302391800), .B(n_27999), .C(n_26054), .D(n_298166510
		), .Z(n_153068547));
	notech_and3 i_148460319(.A(n_140168418), .B(n_125828535), .C(n_121868235
		), .Z(n_153368550));
	notech_ao4 i_144960352(.A(n_157165100), .B(n_313070141), .C(n_56532), .D
		(n_139068407), .Z(n_153568552));
	notech_ao4 i_144860353(.A(n_60011), .B(n_312391700), .C(n_56257), .D(n_183868855
		), .Z(n_153668553));
	notech_ao4 i_144660355(.A(n_313570146), .B(\nbus_11358[14] ), .C(\nbus_11307[14] 
		), .D(n_26597), .Z(n_153868555));
	notech_and4 i_145160350(.A(n_153868555), .B(n_153668553), .C(n_153568552
		), .D(n_121368230), .Z(n_154068557));
	notech_ao4 i_144360358(.A(n_298266511), .B(n_319770208), .C(n_313370144)
		, .D(n_27999), .Z(n_154168558));
	notech_ao3 i_144260359(.A(n_140168418), .B(n_125828535), .C(n_120768224)
		, .Z(n_154468561));
	notech_ao4 i_143860363(.A(n_30109), .B(n_313070141), .C(n_94935745), .D(n_56532
		), .Z(n_154668563));
	notech_ao4 i_143760364(.A(n_302091803), .B(n_312391700), .C(n_183868855)
		, .D(n_29592), .Z(n_154768564));
	notech_ao4 i_143560366(.A(\nbus_11358[13] ), .B(n_313570146), .C(\nbus_11307[13] 
		), .D(n_26597), .Z(n_154968566));
	notech_and4 i_144060361(.A(n_154968566), .B(n_154768564), .C(n_154668563
		), .D(n_120268219), .Z(n_155168568));
	notech_ao4 i_143260369(.A(n_31560), .B(n_319770208), .C(n_313370144), .D
		(n_27998), .Z(n_155268569));
	notech_and3 i_143160370(.A(n_93835734), .B(n_125828535), .C(n_119668213)
		, .Z(n_155568572));
	notech_and3 i_125460541(.A(n_119468211), .B(n_119368210), .C(n_119568212
		), .Z(n_155968576));
	notech_ao4 i_125160544(.A(n_26819), .B(\nbus_11307[14] ), .C(n_60011), .D
		(n_316691657), .Z(n_156068577));
	notech_ao4 i_124860547(.A(n_151028787), .B(nbus_11295[14]), .C(n_58408),
		 .D(n_27999), .Z(n_156368580));
	notech_and4 i_125060545(.A(n_118968206), .B(n_156368580), .C(n_140168418
		), .D(n_118668203), .Z(n_156668583));
	notech_nand2 i_3858483(.A(opc[12]), .B(n_62792), .Z(n_156768584));
	notech_ao4 i_10058391(.A(n_30594), .B(n_60241), .C(n_315191672), .D(n_25010
		), .Z(n_157268589));
	notech_ao4 i_15858335(.A(n_26770), .B(n_27712), .C(n_27163), .D(n_26591)
		, .Z(n_157368590));
	notech_and2 i_15958334(.A(n_199669008), .B(n_58610), .Z(n_157468591));
	notech_and2 i_16058333(.A(n_58646), .B(n_199869010), .Z(n_157568592));
	notech_and2 i_9958392(.A(n_3894), .B(n_307091753), .Z(n_157868595));
	notech_ao4 i_9058401(.A(n_26625), .B(n_26789), .C(n_306991754), .D(n_56508
		), .Z(n_157968596));
	notech_and2 i_15658337(.A(n_26606), .B(n_193668949), .Z(n_158268599));
	notech_nand3 i_72757783(.A(n_60153), .B(n_60241), .C(read_data[0]), .Z(n_158668603
		));
	notech_or2 i_105457473(.A(n_304291781), .B(n_56518), .Z(n_159168608));
	notech_or2 i_29058203(.A(n_151028787), .B(nbus_11295[12]), .Z(n_159668613
		));
	notech_nand2 i_28758206(.A(opb[12]), .B(n_58097), .Z(n_159968616));
	notech_or2 i_28458209(.A(n_60013), .B(n_316691657), .Z(n_160268619));
	notech_ao3 i_37158123(.A(tsc[41]), .B(n_27855), .C(n_24989), .Z(n_160568622
		));
	notech_or2 i_36858126(.A(n_313370144), .B(n_27992), .Z(n_160868625));
	notech_ao3 i_38558109(.A(tsc[42]), .B(n_27855), .C(n_24989), .Z(n_161368630
		));
	notech_or4 i_38458110(.A(n_26939), .B(n_60940), .C(n_28136), .D(n_25010)
		, .Z(n_161668633));
	notech_or2 i_38158113(.A(n_313570146), .B(\nbus_11358[10] ), .Z(n_161968636
		));
	notech_or2 i_37858116(.A(n_3850), .B(n_312391700), .Z(n_162268639));
	notech_nao3 i_39658098(.A(tsc[43]), .B(n_27855), .C(n_24989), .Z(n_162368640
		));
	notech_nao3 i_39558099(.A(n_62820), .B(opc[11]), .C(n_313070141), .Z(n_162668643
		));
	notech_or2 i_39258102(.A(n_313370144), .B(n_27996), .Z(n_162968646));
	notech_ao3 i_40658088(.A(tsc[44]), .B(n_27855), .C(n_24989), .Z(n_163468651
		));
	notech_or4 i_40558089(.A(n_26939), .B(n_28138), .C(n_60940), .D(n_25010)
		, .Z(n_163768654));
	notech_or2 i_40258092(.A(n_313570146), .B(\nbus_11358[12] ), .Z(n_164068657
		));
	notech_or2 i_39958095(.A(n_60013), .B(n_312391700), .Z(n_164368660));
	notech_ao3 i_41658078(.A(tsc[47]), .B(n_27855), .C(n_24989), .Z(n_164668663
		));
	notech_or4 i_41358081(.A(n_26939), .B(n_28141), .C(n_60942), .D(n_25010)
		, .Z(n_164968666));
	notech_or4 i_48658008(.A(n_26062), .B(n_320170212), .C(n_27119), .D(n_26054
		), .Z(n_165468671));
	notech_or2 i_48558009(.A(n_302391800), .B(n_27997), .Z(n_165768674));
	notech_or4 i_48058014(.A(n_3854), .B(n_26054), .C(n_60013), .D(n_58024),
		 .Z(n_166268679));
	notech_or4 i_56157933(.A(n_30854), .B(n_320170212), .C(n_26770), .D(n_58482
		), .Z(n_166368680));
	notech_nand2 i_56057934(.A(n_58378), .B(opd[12]), .Z(n_166668683));
	notech_or2 i_55557939(.A(n_57329), .B(n_60013), .Z(n_167168688));
	notech_nand2 i_57357922(.A(sav_esi[0]), .B(n_61142), .Z(n_167268689));
	notech_or2 i_57257923(.A(n_58383), .B(n_27981), .Z(n_167568692));
	notech_nao3 i_56857926(.A(opc[0]), .B(n_62812), .C(n_185068867), .Z(n_167868695
		));
	notech_or4 i_61357886(.A(n_32348), .B(n_56547), .C(n_3851), .D(n_61142),
		 .Z(n_168968706));
	notech_nand2 i_61057889(.A(opb[10]), .B(n_27289), .Z(n_169268709));
	notech_or2 i_60757892(.A(n_3850), .B(n_313670147), .Z(n_169568712));
	notech_nand3 i_62657873(.A(n_26983), .B(n_60241), .C(read_data[0]), .Z(n_170268719
		));
	notech_or2 i_62357876(.A(n_58370), .B(n_27981), .Z(n_170568722));
	notech_or2 i_62057879(.A(n_57812), .B(\nbus_11358[0] ), .Z(n_170868725)
		);
	notech_or4 i_61457885(.A(n_32459), .B(n_26610), .C(n_27754), .D(n_29742)
		, .Z(n_171168728));
	notech_ao4 i_61557884(.A(n_1448), .B(n_305291771), .C(n_26905), .D(n_26592
		), .Z(n_171268729));
	notech_or2 i_63757864(.A(n_57821), .B(n_29678), .Z(n_172368740));
	notech_or4 i_66557843(.A(n_56834), .B(n_56983), .C(n_5723), .D(n_56518),
		 .Z(n_173068747));
	notech_nand3 i_65957846(.A(n_26983), .B(n_60241), .C(read_data[4]), .Z(n_173368750
		));
	notech_or4 i_65557849(.A(n_62844), .B(n_56508), .C(n_62812), .D(\nbus_11307[4] 
		), .Z(n_173668753));
	notech_or4 i_68057830(.A(n_60942), .B(n_28133), .C(n_305191772), .D(n_26601
		), .Z(n_174368760));
	notech_nand3 i_67757833(.A(n_26983), .B(n_60241), .C(read_data[7]), .Z(n_174668763
		));
	notech_or2 i_67457836(.A(n_303191792), .B(n_58071), .Z(n_174968766));
	notech_or4 i_67157839(.A(n_56834), .B(n_26610), .C(n_303391790), .D(n_56518
		), .Z(n_175268769));
	notech_or2 i_69357817(.A(n_4008), .B(\nbus_11358[10] ), .Z(n_175868775)
		);
	notech_or2 i_69057820(.A(n_3850), .B(n_4007), .Z(n_176168778));
	notech_nand2 i_68757823(.A(\eflags[10] ), .B(n_26593), .Z(n_176468781)
		);
	notech_or2 i_70357807(.A(n_4008), .B(\nbus_11358[12] ), .Z(n_176968786)
		);
	notech_or4 i_69857812(.A(n_62842), .B(n_27761), .C(n_62812), .D(n_29679)
		, .Z(n_177468791));
	notech_or4 i_82757690(.A(n_58810), .B(n_58481), .C(n_28138), .D(n_60942)
		, .Z(n_177568792));
	notech_nand2 i_82657691(.A(n_58377), .B(opd[12]), .Z(n_177868795));
	notech_or2 i_82157696(.A(n_181779321), .B(n_60013), .Z(n_178368800));
	notech_or4 i_86357659(.A(n_58806), .B(n_58477), .C(n_28138), .D(n_60945)
		, .Z(n_178468801));
	notech_or2 i_86257660(.A(n_154331958), .B(nbus_11295[12]), .Z(n_178768804
		));
	notech_nand2 i_85957663(.A(n_58050), .B(opb[12]), .Z(n_179068807));
	notech_or4 i_85557666(.A(n_58132), .B(n_58477), .C(n_60013), .D(n_56908)
		, .Z(n_179368810));
	notech_or4 i_93357590(.A(n_58805), .B(n_28138), .C(n_60942), .D(n_58478)
		, .Z(n_179468811));
	notech_or2 i_93257591(.A(n_58374), .B(n_27997), .Z(n_179768814));
	notech_or2 i_92757596(.A(n_60013), .B(n_57025), .Z(n_180268819));
	notech_or4 i_98057547(.A(n_58817), .B(n_58479), .C(n_28138), .D(n_60942)
		, .Z(n_180368820));
	notech_or4 i_97957548(.A(n_58817), .B(n_58495), .C(n_60942), .D(nbus_11295
		[12]), .Z(n_180668823));
	notech_nand2 i_97557551(.A(n_57179), .B(opb[12]), .Z(n_180968826));
	notech_or2 i_97257554(.A(n_228579786), .B(n_60013), .Z(n_181268829));
	notech_nand3 i_99257535(.A(n_60340), .B(n_299491829), .C(opa[10]), .Z(n_181768834
		));
	notech_or2 i_100757520(.A(n_30568), .B(\nbus_11307[11] ), .Z(n_182268839
		));
	notech_nao3 i_101857509(.A(opc_10[12]), .B(n_62824), .C(n_57473), .Z(n_182368840
		));
	notech_nand2 i_101757510(.A(opc[12]), .B(n_57808), .Z(n_182668843));
	notech_nao3 i_101257515(.A(n_26829), .B(\opa_12[12] ), .C(n_58480), .Z(n_183168848
		));
	notech_ao3 i_102157506(.A(n_60340), .B(\opa_12[12] ), .C(n_30594), .Z(n_183668853
		));
	notech_nand2 i_35027(.A(n_26939), .B(n_26938), .Z(n_183768854));
	notech_nand3 i_35026(.A(n_27221), .B(n_26938), .C(n_57985), .Z(n_183868855
		));
	notech_or2 i_32927(.A(n_300891815), .B(n_27353), .Z(n_184068857));
	notech_or2 i_10758384(.A(n_56508), .B(n_27757), .Z(n_184168858));
	notech_nao3 i_9758394(.A(n_246591944), .B(n_57068), .C(n_56508), .Z(n_184268859
		));
	notech_nao3 i_30209(.A(n_26884), .B(n_32331), .C(n_58099), .Z(n_184368860
		));
	notech_nand2 i_30208(.A(n_58805), .B(n_26884), .Z(n_184468861));
	notech_nao3 i_29393(.A(n_26731), .B(n_32338), .C(n_58480), .Z(n_184668863
		));
	notech_or2 i_29392(.A(n_58480), .B(n_58815), .Z(n_184768864));
	notech_nao3 i_29391(.A(n_26731), .B(n_56457), .C(n_58480), .Z(n_184868865
		));
	notech_or4 i_32359(.A(n_27037), .B(n_3790), .C(n_19086), .D(n_60340), .Z
		(n_184968866));
	notech_or4 i_32911(.A(n_297369985), .B(instrc[116]), .C(n_29658), .D(n_26770
		), .Z(n_185068867));
	notech_ao4 i_192756623(.A(n_304891775), .B(n_314291681), .C(n_306991754)
		, .D(n_56508), .Z(n_185268869));
	notech_or4 i_65158482(.A(calc_sz[1]), .B(n_246691943), .C(n_56834), .D(n_59965
		), .Z(n_185668873));
	notech_ao4 i_185756692(.A(n_57299), .B(n_60013), .C(n_56640), .D(n_185668873
		), .Z(n_185768874));
	notech_ao4 i_185656693(.A(n_57807), .B(\nbus_11358[12] ), .C(n_57809), .D
		(\nbus_11307[12] ), .Z(n_185968876));
	notech_ao4 i_185356696(.A(n_58376), .B(n_27997), .C(n_58480), .D(n_320070211
		), .Z(n_186168878));
	notech_ao4 i_186156688(.A(n_30565), .B(n_60013), .C(n_60340), .D(n_28101
		), .Z(n_186368880));
	notech_ao4 i_186056689(.A(n_30569), .B(\nbus_11358[12] ), .C(n_30568), .D
		(\nbus_11307[12] ), .Z(n_186668882));
	notech_nao3 i_66258477(.A(n_186368880), .B(n_186668882), .C(n_183668853)
		, .Z(n_186768883));
	notech_and4 i_185556694(.A(n_182368840), .B(n_186168878), .C(n_26609), .D
		(n_182668843), .Z(n_186968885));
	notech_ao4 i_185056699(.A(n_30570), .B(n_29596), .C(n_302491799), .D(n_30565
		), .Z(n_187068886));
	notech_ao4 i_184956700(.A(n_28100), .B(n_60340), .C(n_30569), .D(\nbus_11358[11] 
		), .Z(n_187268888));
	notech_and3 i_66158478(.A(n_187068886), .B(n_187268888), .C(n_182268839)
		, .Z(n_187368889));
	notech_or4 i_65358481(.A(calc_sz[1]), .B(n_246691943), .C(n_56834), .D(n_3851
		), .Z(n_187568890));
	notech_ao4 i_183856711(.A(n_30570), .B(n_29684), .C(n_3850), .D(n_30565)
		, .Z(n_187668891));
	notech_ao4 i_183756712(.A(n_28099), .B(n_60338), .C(n_30569), .D(\nbus_11358[10] 
		), .Z(n_187868893));
	notech_and3 i_66058479(.A(n_187668891), .B(n_187868893), .C(n_181768834)
		, .Z(n_187968894));
	notech_ao4 i_182656723(.A(n_323080731), .B(n_156768584), .C(n_56666), .D
		(n_185668873), .Z(n_188068895));
	notech_ao4 i_182456725(.A(n_26856), .B(\nbus_11307[12] ), .C(n_322980730
		), .D(n_29679), .Z(n_188268897));
	notech_and4 i_182856721(.A(n_188268897), .B(n_188068895), .C(n_180968826
		), .D(n_181268829), .Z(n_188468899));
	notech_ao4 i_182156728(.A(n_58375), .B(n_27997), .C(n_58479), .D(n_320070211
		), .Z(n_188568900));
	notech_and4 i_182356726(.A(n_180368820), .B(n_188568900), .C(n_26609), .D
		(n_180668823), .Z(n_188868903));
	notech_ao4 i_178756761(.A(n_156768584), .B(n_313270143), .C(n_56653), .D
		(n_185668873), .Z(n_188968904));
	notech_ao4 i_178656762(.A(\nbus_11307[12] ), .B(n_26607), .C(n_319970210
		), .D(n_29679), .Z(n_189268906));
	notech_ao4 i_178356765(.A(n_320070211), .B(n_58478), .C(n_57181), .D(\nbus_11358[12] 
		), .Z(n_189468908));
	notech_and4 i_178556763(.A(n_189468908), .B(n_26609), .C(n_179468811), .D
		(n_179768814), .Z(n_189768911));
	notech_ao4 i_172756821(.A(n_58041), .B(n_156768584), .C(n_56919), .D(n_185668873
		), .Z(n_189868912));
	notech_ao4 i_172556823(.A(n_26854), .B(\nbus_11307[12] ), .C(n_322680727
		), .D(n_29679), .Z(n_190068914));
	notech_and4 i_172956819(.A(n_190068914), .B(n_179368810), .C(n_189868912
		), .D(n_179068807), .Z(n_190268916));
	notech_ao4 i_172256826(.A(n_58372), .B(n_27997), .C(n_58477), .D(n_320070211
		), .Z(n_190368917));
	notech_and4 i_172456824(.A(n_178468801), .B(n_190368917), .C(n_26609), .D
		(n_178768804), .Z(n_190768920));
	notech_ao4 i_169956849(.A(n_58038), .B(n_156768584), .C(n_56502), .D(n_185668873
		), .Z(n_190868921));
	notech_ao4 i_169856850(.A(n_26851), .B(\nbus_11307[12] ), .C(n_197279473
		), .D(n_29679), .Z(n_191068923));
	notech_ao4 i_169556853(.A(n_58481), .B(n_320070211), .C(n_58052), .D(\nbus_11358[12] 
		), .Z(n_191268925));
	notech_and4 i_169756851(.A(n_177568792), .B(n_191268925), .C(n_26609), .D
		(n_177868795), .Z(n_191568928));
	notech_ao4 i_155456991(.A(n_156768584), .B(n_4009), .C(n_56518), .D(n_185668873
		), .Z(n_191768930));
	notech_ao4 i_155356992(.A(n_60013), .B(n_4007), .C(n_308091743), .D(n_28101
		), .Z(n_191968932));
	notech_and3 i_155656989(.A(n_191768930), .B(n_191968932), .C(n_177468791
		), .Z(n_192068933));
	notech_ao4 i_155056995(.A(\nbus_11307[12] ), .B(n_26598), .C(n_313970150
		), .D(n_29679), .Z(n_192168934));
	notech_ao4 i_154956996(.A(n_320170212), .B(n_307991744), .C(n_27997), .D
		(n_4013), .Z(n_192368936));
	notech_ao4 i_154656999(.A(n_87532846), .B(n_4009), .C(n_26649), .D(n_187568890
		), .Z(n_192568938));
	notech_ao4 i_154457001(.A(n_308091743), .B(n_28099), .C(n_31411), .D(n_27761
		), .Z(n_192768940));
	notech_and4 i_154856997(.A(n_192768940), .B(n_192568938), .C(n_176168778
		), .D(n_176468781), .Z(n_192968942));
	notech_ao4 i_154157004(.A(\nbus_11307[10] ), .B(n_26598), .C(n_313970150
		), .D(n_29684), .Z(n_193068943));
	notech_ao4 i_154057005(.A(n_31433), .B(n_307991744), .C(n_27993), .D(n_4013
		), .Z(n_193268945));
	notech_nao3 i_153957006(.A(n_27377), .B(n_60338), .C(n_26610), .Z(n_193468947
		));
	notech_ao4 i_7858413(.A(n_306891755), .B(n_305191772), .C(n_32459), .D(n_193468947
		), .Z(n_193568948));
	notech_ao4 i_153857007(.A(n_26789), .B(n_26625), .C(n_304591778), .D(n_56508
		), .Z(n_193668949));
	notech_ao4 i_153557010(.A(\nbus_11307[7] ), .B(n_158268599), .C(n_193568948
		), .D(n_29614), .Z(n_193768950));
	notech_ao4 i_153257012(.A(n_57812), .B(\nbus_11358[7] ), .C(n_31307), .D
		(n_184268859), .Z(n_193968952));
	notech_and4 i_153757008(.A(n_193968952), .B(n_175268769), .C(n_193768950
		), .D(n_174968766), .Z(n_194168954));
	notech_ao4 i_152957015(.A(n_307091753), .B(n_27383), .C(n_58370), .D(n_27990
		), .Z(n_194268955));
	notech_ao4 i_152757017(.A(n_3997), .B(n_3996), .C(n_31279), .D(n_305191772
		), .Z(n_194468957));
	notech_and4 i_153157013(.A(n_194468957), .B(n_194268955), .C(n_174368760
		), .D(n_174668763), .Z(n_194668959));
	notech_ao4 i_152457020(.A(n_157868595), .B(n_27382), .C(n_184168858), .D
		(n_291663183), .Z(n_194768960));
	notech_ao4 i_152357021(.A(n_157968596), .B(\nbus_11307[4] ), .C(n_291763184
		), .D(n_184268859), .Z(n_194868961));
	notech_ao4 i_152157023(.A(n_57812), .B(\nbus_11358[4] ), .C(n_193568948)
		, .D(n_29725), .Z(n_195068963));
	notech_and4 i_152657018(.A(n_195068963), .B(n_194868961), .C(n_194768960
		), .D(n_173668753), .Z(n_195268965));
	notech_ao4 i_151857026(.A(n_27986), .B(n_58370), .C(n_5743), .D(n_58071)
		, .Z(n_195368966));
	notech_ao4 i_151657028(.A(n_291863185), .B(n_343270443), .C(n_291463181)
		, .D(n_305191772), .Z(n_195568968));
	notech_and4 i_152057024(.A(n_195568968), .B(n_195368966), .C(n_173068747
		), .D(n_173368750), .Z(n_195768970));
	notech_ao4 i_150657037(.A(n_297966508), .B(n_184268859), .C(n_297866507)
		, .D(n_184168858), .Z(n_195868971));
	notech_ao4 i_150557038(.A(n_184968866), .B(n_28090), .C(n_57812), .D(\nbus_11358[1] 
		), .Z(n_195968972));
	notech_ao4 i_150357040(.A(n_57711), .B(\nbus_11307[1] ), .C(n_297766506)
		, .D(n_56508), .Z(n_196168974));
	notech_and4 i_150857035(.A(n_196168974), .B(n_195968972), .C(n_195868971
		), .D(n_172368740), .Z(n_196368976));
	notech_ao4 i_150057043(.A(n_58370), .B(n_27983), .C(n_60024), .D(n_58071
		), .Z(n_196468977));
	notech_ao4 i_149957044(.A(n_297666505), .B(n_305191772), .C(n_308091743)
		, .D(n_19014), .Z(n_196568978));
	notech_ao4 i_149757046(.A(n_59992), .B(n_211169123), .C(n_298066509), .D
		(n_343270443), .Z(n_196768980));
	notech_and4 i_150257041(.A(n_196768980), .B(n_196568978), .C(n_196468977
		), .D(n_307091753), .Z(n_196968982));
	notech_ao4 i_149457049(.A(n_291363180), .B(n_27757), .C(n_306991754), .D
		(n_29742), .Z(n_197268985));
	notech_ao4 i_149057053(.A(n_157868595), .B(n_27381), .C(n_175062033), .D
		(n_184168858), .Z(n_197468987));
	notech_ao3 i_149257051(.A(n_171168728), .B(n_197468987), .C(n_171268729)
		, .Z(n_197568988));
	notech_ao4 i_148857055(.A(n_157968596), .B(\nbus_11307[0] ), .C(n_291263179
		), .D(n_184268859), .Z(n_197668989));
	notech_ao4 i_148557058(.A(n_60025), .B(n_58071), .C(n_58646), .D(n_56508
		), .Z(n_198068992));
	notech_ao4 i_148357060(.A(n_291163178), .B(n_343270443), .C(n_59993), .D
		(n_211169123), .Z(n_198268994));
	notech_and4 i_148757056(.A(n_198268994), .B(n_198068992), .C(n_170268719
		), .D(n_170568722), .Z(n_198468996));
	notech_ao4 i_148057063(.A(n_27334), .B(n_29880), .C(n_27335), .D(n_29879
		), .Z(n_198568997));
	notech_ao4 i_147957064(.A(n_31411), .B(n_27349), .C(n_87532846), .D(n_27157
		), .Z(n_198668998));
	notech_ao4 i_147757066(.A(n_59326), .B(n_28099), .C(n_60153), .D(n_27199
		), .Z(n_198869000));
	notech_and4 i_148257061(.A(n_198869000), .B(n_198668998), .C(n_198568997
		), .D(n_169568712), .Z(n_199069002));
	notech_ao4 i_147457069(.A(n_302691797), .B(\nbus_11307[10] ), .C(n_313770148
		), .D(n_29684), .Z(n_199169003));
	notech_ao4 i_147257071(.A(n_31433), .B(n_27348), .C(n_302591798), .D(n_27993
		), .Z(n_199369005));
	notech_and4 i_147657067(.A(n_199369005), .B(n_199169003), .C(n_168968706
		), .D(n_169268709), .Z(n_199569007));
	notech_ao4 i_143157111(.A(n_29742), .B(n_1393), .C(n_60025), .D(n_26815)
		, .Z(n_199669008));
	notech_ao4 i_142757115(.A(n_300891815), .B(n_157468591), .C(n_175062033)
		, .D(n_26605), .Z(n_199769009));
	notech_ao4 i_143057112(.A(n_1393), .B(\nbus_11307[0] ), .C(\nbus_11358[0] 
		), .D(n_26815), .Z(n_199869010));
	notech_ao4 i_142657116(.A(n_27335), .B(n_29878), .C(n_297369985), .D(n_157568592
		), .Z(n_199969011));
	notech_ao4 i_142457118(.A(n_291363180), .B(n_184068857), .C(n_27334), .D
		(n_29877), .Z(n_200169013));
	notech_and4 i_142957113(.A(n_200169013), .B(n_199969011), .C(n_199769009
		), .D(n_167868695), .Z(n_200369015));
	notech_ao4 i_142157121(.A(n_59993), .B(n_303691787), .C(n_291163178), .D
		(n_274369755), .Z(n_200469016));
	notech_and4 i_142057122(.A(n_185362136), .B(n_158668603), .C(n_185262135
		), .D(n_167268689), .Z(n_200769019));
	notech_ao4 i_141657126(.A(n_58040), .B(n_156768584), .C(n_56489), .D(n_185668873
		), .Z(n_200969021));
	notech_ao4 i_141557127(.A(\nbus_11307[12] ), .B(n_26679), .C(n_325273732
		), .D(n_29679), .Z(n_201169023));
	notech_ao4 i_141157130(.A(n_320070211), .B(n_58482), .C(n_58054), .D(\nbus_11358[12] 
		), .Z(n_201369025));
	notech_and4 i_141357128(.A(n_166368680), .B(n_201369025), .C(n_26609), .D
		(n_166668683), .Z(n_201669028));
	notech_ao4 i_135657185(.A(n_301991804), .B(n_156768584), .C(n_56605), .D
		(n_185668873), .Z(n_201769029));
	notech_ao4 i_135557186(.A(\nbus_11307[12] ), .B(n_27293), .C(n_322480725
		), .D(n_29679), .Z(n_201969031));
	notech_ao4 i_135257189(.A(n_26054), .B(n_320070211), .C(n_302291801), .D
		(\nbus_11358[12] ), .Z(n_202169033));
	notech_and4 i_135457187(.A(n_202169033), .B(n_26609), .C(n_165468671), .D
		(n_165768674), .Z(n_202469036));
	notech_ao4 i_128857248(.A(n_58622), .B(n_25010), .C(n_157268589), .D(n_29754
		), .Z(n_202569037));
	notech_ao4 i_128757249(.A(n_320538000), .B(n_56532), .C(n_313370144), .D
		(n_28000), .Z(n_202669038));
	notech_ao4 i_128557251(.A(n_313570146), .B(\nbus_11358[15] ), .C(\nbus_11307[15] 
		), .D(n_26597), .Z(n_202869040));
	notech_and4 i_129057246(.A(n_164968666), .B(n_202869040), .C(n_202669038
		), .D(n_202569037), .Z(n_203069042));
	notech_ao4 i_128257254(.A(n_60010), .B(n_312391700), .C(n_111064639), .D
		(n_313070141), .Z(n_203169043));
	notech_nand3 i_128157255(.A(n_3849), .B(n_115075094), .C(n_115175095), .Z
		(n_203469046));
	notech_ao4 i_127757259(.A(n_156768584), .B(n_313070141), .C(n_56532), .D
		(n_185668873), .Z(n_203669048));
	notech_ao4 i_127557261(.A(\nbus_11307[12] ), .B(n_26597), .C(n_29679), .D
		(n_312870139), .Z(n_203869050));
	notech_and4 i_127957257(.A(n_203869050), .B(n_203669048), .C(n_164068657
		), .D(n_164368660), .Z(n_204069052));
	notech_ao4 i_127257264(.A(n_313370144), .B(n_27997), .C(n_25010), .D(n_320070211
		), .Z(n_204169053));
	notech_nand2 i_127357263(.A(n_204169053), .B(n_163768654), .Z(n_204269054
		));
	notech_ao4 i_126857268(.A(n_183868855), .B(n_29596), .C(n_31492), .D(n_183768854
		), .Z(n_204569057));
	notech_ao4 i_126757269(.A(\nbus_11307[11] ), .B(n_26597), .C(n_302491799
		), .D(n_312391700), .Z(n_204669058));
	notech_ao4 i_126557271(.A(n_31456), .B(n_25010), .C(n_313570146), .D(\nbus_11358[11] 
		), .Z(n_204869060));
	notech_and4 i_127057266(.A(n_204869060), .B(n_204669058), .C(n_204569057
		), .D(n_162968646), .Z(n_205069062));
	notech_ao4 i_126257274(.A(n_31476), .B(n_319770208), .C(n_30528), .D(n_56532
		), .Z(n_205169063));
	notech_and3 i_126157275(.A(n_187368889), .B(n_125828535), .C(n_162368640
		), .Z(n_205469066));
	notech_ao4 i_125757279(.A(n_87532846), .B(n_313070141), .C(n_56532), .D(n_187568890
		), .Z(n_205669068));
	notech_ao4 i_125557281(.A(\nbus_11307[10] ), .B(n_26597), .C(n_312870139
		), .D(n_29684), .Z(n_205869070));
	notech_and4 i_125957277(.A(n_205869070), .B(n_205669068), .C(n_161968636
		), .D(n_162268639), .Z(n_206069072));
	notech_ao4 i_125157284(.A(n_313370144), .B(n_27993), .C(n_31411), .D(n_25010
		), .Z(n_206169073));
	notech_ao3 i_125057285(.A(n_187968894), .B(n_125828535), .C(n_161368630)
		, .Z(n_206469076));
	notech_ao4 i_124657289(.A(n_208969101), .B(n_26927), .C(n_157268589), .D
		(n_29743), .Z(n_206669078));
	notech_ao4 i_124557290(.A(n_60016), .B(n_312391700), .C(\nbus_11307[9] )
		, .D(n_26597), .Z(n_206769079));
	notech_ao4 i_124357292(.A(n_58608), .B(n_25010), .C(n_313570146), .D(\nbus_11358[9] 
		), .Z(n_206969081));
	notech_and4 i_124857287(.A(n_206969081), .B(n_206769079), .C(n_206669078
		), .D(n_160868625), .Z(n_207169083));
	notech_ao4 i_124057295(.A(n_189962171), .B(n_313070141), .C(n_291963186)
		, .D(n_319770208), .Z(n_207269084));
	notech_ao4 i_10158390(.A(n_28098), .B(n_60338), .C(n_30569), .D(\nbus_11358[9] 
		), .Z(n_207469086));
	notech_ao4 i_10258389(.A(\nbus_11307[9] ), .B(n_30568), .C(n_60016), .D(n_30565
		), .Z(n_207569087));
	notech_nand3 i_123957296(.A(n_207569087), .B(n_207469086), .C(n_125828535
		), .Z(n_207769089));
	notech_ao4 i_116757363(.A(n_156768584), .B(n_312970140), .C(n_56583), .D
		(n_185668873), .Z(n_207969091));
	notech_ao4 i_116557365(.A(n_26819), .B(\nbus_11307[12] ), .C(n_57415), .D
		(n_29679), .Z(n_208169093));
	notech_and4 i_116957361(.A(n_208169093), .B(n_207969091), .C(n_159968616
		), .D(n_160268619), .Z(n_208369095));
	notech_ao4 i_116257368(.A(n_58408), .B(n_27997), .C(n_23512), .D(n_320070211
		), .Z(n_208469096));
	notech_ao4 i_116057370(.A(n_54643), .B(n_28952), .C(n_320170212), .D(n_319670207
		), .Z(n_208669098));
	notech_and4 i_116457366(.A(n_208669098), .B(n_208469096), .C(n_159668613
		), .D(n_26609), .Z(n_208869100));
	notech_or4 i_76555593(.A(calc_sz[1]), .B(n_246691943), .C(n_56834), .D(n_59968
		), .Z(n_208969101));
	notech_nand3 i_190455512(.A(n_56848), .B(n_187762157), .C(n_58494), .Z(n_209069102
		));
	notech_nor2 i_35255172(.A(n_58429), .B(n_28015), .Z(n_209269104));
	notech_or2 i_34755177(.A(n_57868), .B(\nbus_11365[30] ), .Z(n_209969111)
		);
	notech_nand2 i_37855146(.A(n_57481), .B(opa[9]), .Z(n_210469116));
	notech_or2 i_37555149(.A(n_57627), .B(n_29743), .Z(n_210769119));
	notech_or2 i_37255152(.A(n_57775), .B(n_60016), .Z(n_211069122));
	notech_nao3 i_32363(.A(n_32386), .B(n_32294), .C(n_56837), .Z(n_211169123
		));
	notech_ao4 i_79454773(.A(n_26649), .B(n_58106), .C(n_189962171), .D(n_171965248
		), .Z(n_211369125));
	notech_ao4 i_79254775(.A(n_291963186), .B(n_307991744), .C(n_308091743),
		 .D(n_28098), .Z(n_211569127));
	notech_and4 i_79654771(.A(n_211569127), .B(n_211369125), .C(n_210769119)
		, .D(n_211069122), .Z(n_211769129));
	notech_ao4 i_78954778(.A(n_57490), .B(\nbus_11358[9] ), .C(n_211169123),
		 .D(n_27992), .Z(n_211869130));
	notech_ao4 i_78854779(.A(n_27761), .B(n_58608), .C(n_29789), .D(n_307091753
		), .Z(n_212069132));
	notech_ao4 i_74954812(.A(n_154831963), .B(n_303091793), .C(n_151931934),
		 .D(n_30809), .Z(n_212269134));
	notech_ao4 i_74854813(.A(n_58084), .B(n_32252), .C(n_57875), .D(\nbus_11358[30] 
		), .Z(n_212469136));
	notech_nand3 i_75254810(.A(n_212269134), .B(n_212469136), .C(n_209969111
		), .Z(n_212569137));
	notech_ao4 i_74654815(.A(n_26929), .B(n_29591), .C(n_58147), .D(n_302991794
		), .Z(n_212669138));
	notech_or4 i_4953863(.A(n_32643), .B(n_2875), .C(n_2877), .D(n_60868), .Z
		(n_212969141));
	notech_nao3 i_5153861(.A(n_60153), .B(n_60338), .C(n_58740), .Z(n_213069142
		));
	notech_nand3 i_5253860(.A(n_60144), .B(n_60349), .C(n_326090758), .Z(n_213169143
		));
	notech_nao3 i_1453895(.A(n_346670477), .B(n_213069142), .C(n_349480995),
		 .Z(n_213369145));
	notech_nand2 i_5353859(.A(eval_flag), .B(n_213369145), .Z(n_213469146)
		);
	notech_nand3 i_49796(.A(n_221669228), .B(n_213469146), .C(n_213169143), 
		.Z(n_15683));
	notech_or2 i_51253439(.A(n_287827260), .B(n_3982), .Z(n_213569147));
	notech_or4 i_51153440(.A(n_56837), .B(n_56939), .C(n_56666), .D(n_28013)
		, .Z(n_214069152));
	notech_nand3 i_2920882(.A(n_222369235), .B(n_222269234), .C(n_213569147)
		, .Z(n_24250));
	notech_nor2 i_52953422(.A(n_287827260), .B(n_4016), .Z(n_214369155));
	notech_nao3 i_52353428(.A(n_62820), .B(opc_10[27]), .C(n_286827250), .Z(n_214469156
		));
	notech_or4 i_52853423(.A(n_56834), .B(n_56939), .C(n_56666), .D(n_28012)
		, .Z(n_214969161));
	notech_ao3 i_53053421(.A(opc[27]), .B(n_62824), .C(n_286927251), .Z(n_215069162
		));
	notech_or4 i_2820881(.A(n_222969241), .B(n_222669238), .C(n_215069162), 
		.D(n_214369155), .Z(n_24244));
	notech_or2 i_54453407(.A(n_287827260), .B(n_3983), .Z(n_215169163));
	notech_or4 i_54353408(.A(n_56834), .B(n_56939), .C(n_56666), .D(n_28011)
		, .Z(n_215669168));
	notech_nand3 i_2720880(.A(n_223769249), .B(n_223669248), .C(n_215169163)
		, .Z(n_24238));
	notech_or2 i_59453358(.A(n_4016), .B(n_306824332), .Z(n_215969171));
	notech_ao3 i_58853364(.A(n_62820), .B(opc_10[27]), .C(n_306624330), .Z(n_216069172
		));
	notech_or4 i_59353359(.A(n_56834), .B(n_56939), .C(n_56653), .D(n_28012)
		, .Z(n_216569177));
	notech_or4 i_59553357(.A(n_58805), .B(n_58494), .C(nbus_11295[27]), .D(n_60942
		), .Z(n_216669178));
	notech_nand3 i_2821009(.A(n_224469256), .B(n_216669178), .C(n_215969171)
		, .Z(n_23896));
	notech_or2 i_73153225(.A(n_305924323), .B(n_4016), .Z(n_216769179));
	notech_nor2 i_72453232(.A(n_154331958), .B(nbus_11295[27]), .Z(n_216869180
		));
	notech_or4 i_73253224(.A(n_58806), .B(n_58493), .C(nbus_11295[27]), .D(n_60942
		), .Z(n_217569187));
	notech_nand3 i_2821105(.A(n_225269264), .B(n_217569187), .C(n_216769179)
		, .Z(n_18991));
	notech_or2 i_78153175(.A(n_321538010), .B(n_3982), .Z(n_217669188));
	notech_or4 i_78053176(.A(n_56834), .B(n_56935), .C(n_56502), .D(n_28013)
		, .Z(n_218169193));
	notech_nand3 i_2921202(.A(n_225969271), .B(n_225869270), .C(n_217669188)
		, .Z(n_18648));
	notech_or2 i_80053158(.A(n_321538010), .B(n_4016), .Z(n_218469196));
	notech_ao3 i_79453164(.A(n_62820), .B(opc_10[27]), .C(n_319937994), .Z(n_218569197
		));
	notech_or4 i_79953159(.A(n_56832), .B(n_56935), .C(n_56502), .D(n_28012)
		, .Z(n_219069202));
	notech_or4 i_80153157(.A(n_58497), .B(n_58810), .C(nbus_11295[27]), .D(n_60942
		), .Z(n_219169203));
	notech_nand3 i_2821201(.A(n_226669278), .B(n_219169203), .C(n_218469196)
		, .Z(n_18642));
	notech_or2 i_81653143(.A(n_321538010), .B(n_3983), .Z(n_219269204));
	notech_or4 i_81553144(.A(n_56832), .B(n_56935), .C(n_56502), .D(n_28011)
		, .Z(n_219769209));
	notech_nand3 i_2721200(.A(n_227369285), .B(n_227269284), .C(n_219269204)
		, .Z(n_18636));
	notech_or2 i_128852682(.A(n_4016), .B(n_154831963), .Z(n_220069212));
	notech_ao3 i_128252688(.A(n_62818), .B(opc_10[27]), .C(n_151931934), .Z(n_220169213
		));
	notech_or4 i_128752683(.A(n_246891941), .B(n_2479), .C(n_56688), .D(n_28012
		), .Z(n_220669218));
	notech_or4 i_128952681(.A(n_58802), .B(n_58498), .C(nbus_11295[27]), .D(n_60942
		), .Z(n_220769219));
	notech_nand3 i_2821649(.A(n_228069292), .B(n_220769219), .C(n_220069212)
		, .Z(n_17942));
	notech_or2 i_145952516(.A(n_4016), .B(n_3837), .Z(n_220869220));
	notech_ao3 i_145352522(.A(n_62826), .B(opc_10[27]), .C(n_3843), .Z(n_220969221
		));
	notech_or4 i_145852517(.A(n_56832), .B(n_56935), .C(n_56605), .D(n_28012
		), .Z(n_221469226));
	notech_or4 i_146052515(.A(n_3845), .B(n_26767), .C(nbus_11295[27]), .D(n_60942
		), .Z(n_221569227));
	notech_nand3 i_2821873(.A(n_228769299), .B(n_221569227), .C(n_220869220)
		, .Z(n_20780));
	notech_nao3 i_185464477(.A(n_60144), .B(n_60349), .C(n_32446), .Z(n_221669228
		));
	notech_ao4 i_51653435(.A(n_26615), .B(n_29662), .C(n_130528582), .D(n_58139
		), .Z(n_221869230));
	notech_ao4 i_51553436(.A(n_57863), .B(\nbus_11358[28] ), .C(n_57861), .D
		(\nbus_11365[28] ), .Z(n_221969231));
	notech_and4 i_51953432(.A(n_221969231), .B(n_221869230), .C(n_242259503)
		, .D(n_214069152), .Z(n_222269234));
	notech_ao4 i_52053431(.A(n_286927251), .B(n_172792106), .C(n_286827250),
		 .D(n_174492092), .Z(n_222369235));
	notech_nao3 i_53453417(.A(n_214969161), .B(n_214469156), .C(n_1978), .Z(n_222669238
		));
	notech_ao4 i_53253419(.A(n_57863), .B(\nbus_11358[27] ), .C(n_57861), .D
		(\nbus_11365[27] ), .Z(n_222769239));
	notech_ao4 i_53353418(.A(n_26615), .B(n_29661), .C(n_131228589), .D(n_58139
		), .Z(n_222869240));
	notech_nand2 i_53553416(.A(n_222869240), .B(n_222769239), .Z(n_222969241
		));
	notech_ao4 i_54853403(.A(n_26615), .B(n_29660), .C(n_133728614), .D(n_58139
		), .Z(n_223269244));
	notech_ao4 i_54753404(.A(n_57863), .B(\nbus_11358[26] ), .C(n_57861), .D
		(\nbus_11365[26] ), .Z(n_223369245));
	notech_and4 i_55153400(.A(n_223369245), .B(n_223269244), .C(n_174892088)
		, .D(n_215669168), .Z(n_223669248));
	notech_ao4 i_55253399(.A(n_286927251), .B(n_174292094), .C(n_286827250),
		 .D(n_174992087), .Z(n_223769249));
	notech_nor2 i_59653356(.A(n_1978), .B(n_216069172), .Z(n_223969251));
	notech_ao4 i_59753355(.A(n_57864), .B(\nbus_11358[27] ), .C(n_314047718)
		, .D(\nbus_11365[27] ), .Z(n_224169253));
	notech_ao4 i_59853354(.A(n_307324337), .B(n_29661), .C(n_131228589), .D(n_58141
		), .Z(n_224269254));
	notech_and4 i_60153351(.A(n_224269254), .B(n_224169253), .C(n_216569177)
		, .D(n_223969251), .Z(n_224469256));
	notech_nor2 i_73353223(.A(n_1978), .B(n_216869180), .Z(n_224669258));
	notech_ao4 i_73453222(.A(n_57870), .B(\nbus_11365[27] ), .C(n_306124325)
		, .D(n_310091723), .Z(n_224769259));
	notech_ao4 i_73553221(.A(n_131228589), .B(n_58143), .C(n_57877), .D(\nbus_11358[27] 
		), .Z(n_224969261));
	notech_ao4 i_73653220(.A(n_58427), .B(n_28012), .C(n_29661), .D(n_26902)
		, .Z(n_225069262));
	notech_and4 i_73953217(.A(n_225069262), .B(n_224969261), .C(n_224769259)
		, .D(n_224669258), .Z(n_225269264));
	notech_ao4 i_78553171(.A(n_26918), .B(n_29662), .C(n_58145), .D(n_130528582
		), .Z(n_225469266));
	notech_ao4 i_78453172(.A(n_57873), .B(\nbus_11358[28] ), .C(n_57869), .D
		(\nbus_11365[28] ), .Z(n_225569267));
	notech_and4 i_78853168(.A(n_225569267), .B(n_225469266), .C(n_242259503)
		, .D(n_218169193), .Z(n_225869270));
	notech_ao4 i_78953167(.A(n_58082), .B(n_172792106), .C(n_319937994), .D(n_174492092
		), .Z(n_225969271));
	notech_nor2 i_80253156(.A(n_1978), .B(n_218569197), .Z(n_226169273));
	notech_ao4 i_80453155(.A(n_57873), .B(\nbus_11358[27] ), .C(n_57869), .D
		(\nbus_11365[27] ), .Z(n_226369275));
	notech_ao4 i_80553154(.A(n_29661), .B(n_26918), .C(n_131228589), .D(n_58145
		), .Z(n_226469276));
	notech_and4 i_80853151(.A(n_226469276), .B(n_226369275), .C(n_219069202)
		, .D(n_226169273), .Z(n_226669278));
	notech_ao4 i_82053139(.A(n_26918), .B(n_29660), .C(n_58145), .D(n_133728614
		), .Z(n_226869280));
	notech_ao4 i_81953140(.A(n_57873), .B(\nbus_11358[26] ), .C(n_57869), .D
		(\nbus_11365[26] ), .Z(n_226969281));
	notech_and4 i_82353136(.A(n_226969281), .B(n_226869280), .C(n_174892088)
		, .D(n_219769209), .Z(n_227269284));
	notech_ao4 i_82453135(.A(n_58082), .B(n_174292094), .C(n_319937994), .D(n_174992087
		), .Z(n_227369285));
	notech_nor2 i_129052680(.A(n_1978), .B(n_220169213), .Z(n_227569287));
	notech_ao4 i_129152679(.A(n_57875), .B(\nbus_11358[27] ), .C(n_57868), .D
		(\nbus_11365[27] ), .Z(n_227769289));
	notech_ao4 i_129252678(.A(n_29661), .B(n_26929), .C(n_131228589), .D(n_58147
		), .Z(n_227869290));
	notech_and4 i_129552675(.A(n_227869290), .B(n_227769289), .C(n_220669218
		), .D(n_227569287), .Z(n_228069292));
	notech_nor2 i_146152514(.A(n_1978), .B(n_220969221), .Z(n_228269294));
	notech_ao4 i_146252513(.A(n_3877), .B(\nbus_11358[27] ), .C(n_3878), .D(\nbus_11365[27] 
		), .Z(n_228469296));
	notech_ao4 i_146352512(.A(n_26642), .B(n_29661), .C(n_148228759), .D(n_131228589
		), .Z(n_228569297));
	notech_and4 i_146652509(.A(n_228569297), .B(n_228469296), .C(n_221469226
		), .D(n_228269294), .Z(n_228769299));
	notech_and2 i_5250614(.A(n_269569707), .B(n_58714), .Z(n_228969301));
	notech_and2 i_5350613(.A(n_58717), .B(n_269669708), .Z(n_229069302));
	notech_mux2 i_4450622(.S(n_32318), .A(n_285027232), .B(n_284927231), .Z(n_229169303
		));
	notech_and2 i_4550621(.A(n_265269664), .B(n_58714), .Z(n_229269304));
	notech_ao3 i_8950577(.A(tsc[22]), .B(n_27855), .C(n_24989), .Z(n_229769309
		));
	notech_or2 i_8850578(.A(n_151028787), .B(nbus_11295[22]), .Z(n_230069312
		));
	notech_or2 i_8550581(.A(n_60003), .B(n_151428791), .Z(n_230369315));
	notech_or2 i_8250584(.A(n_289227274), .B(n_151128788), .Z(n_230669318)
		);
	notech_ao3 i_9950567(.A(tsc[23]), .B(n_27855), .C(n_24989), .Z(n_230769319
		));
	notech_or2 i_9850568(.A(n_151028787), .B(nbus_11295[23]), .Z(n_231069322
		));
	notech_or2 i_9550571(.A(n_60002), .B(n_151428791), .Z(n_231369325));
	notech_or2 i_9250574(.A(n_289127273), .B(n_151128788), .Z(n_231669328)
		);
	notech_ao3 i_12050547(.A(tsc[25]), .B(n_27855), .C(n_24989), .Z(n_231769329
		));
	notech_or2 i_11950548(.A(n_151028787), .B(nbus_11295[25]), .Z(n_232069332
		));
	notech_or2 i_11650551(.A(n_151428791), .B(n_60000), .Z(n_232369335));
	notech_or2 i_11250554(.A(n_151128788), .B(n_288927271), .Z(n_232669338)
		);
	notech_or2 i_18050487(.A(n_150528782), .B(\nbus_11358[25] ), .Z(n_233169343
		));
	notech_or4 i_17750490(.A(n_61138), .B(n_60338), .C(n_19086), .D(n_28114)
		, .Z(n_233469346));
	notech_or2 i_17450493(.A(n_150228779), .B(n_288927271), .Z(n_233769349)
		);
	notech_or2 i_19150476(.A(n_57891), .B(n_57557), .Z(n_234269354));
	notech_or2 i_18850479(.A(n_59991), .B(n_311791706), .Z(n_234569357));
	notech_or4 i_18550482(.A(n_62842), .B(n_305970070), .C(n_60942), .D(n_57557
		), .Z(n_234869360));
	notech_or4 i_23250435(.A(n_56832), .B(n_56935), .C(n_26927), .D(n_28010)
		, .Z(n_235669368));
	notech_or2 i_22750440(.A(n_148728764), .B(n_288927271), .Z(n_236169373)
		);
	notech_or2 i_27250396(.A(n_3878), .B(\nbus_11365[24] ), .Z(n_236469376)
		);
	notech_or2 i_26750401(.A(n_289027272), .B(n_3837), .Z(n_236969381));
	notech_nor2 i_28050388(.A(n_3878), .B(\nbus_11365[25] ), .Z(n_237069382)
		);
	notech_or2 i_27550393(.A(n_3837), .B(n_288927271), .Z(n_237769389));
	notech_nor2 i_39750271(.A(n_57868), .B(\nbus_11365[25] ), .Z(n_237869390
		));
	notech_or2 i_39250276(.A(n_154831963), .B(n_288927271), .Z(n_238569397)
		);
	notech_nand2 i_40750264(.A(sav_esi[2]), .B(n_61138), .Z(n_239469406));
	notech_nand3 i_46650206(.A(n_1429), .B(n_7332), .C(\eflags[10] ), .Z(n_240369415
		));
	notech_or2 i_46350209(.A(n_144928726), .B(\nbus_11358[25] ), .Z(n_240669418
		));
	notech_nand3 i_46050212(.A(n_60144), .B(n_60241), .C(read_data[25]), .Z(n_240969421
		));
	notech_or2 i_45750215(.A(n_144428721), .B(n_288927271), .Z(n_241269424)
		);
	notech_or2 i_46950203(.A(n_289227274), .B(n_309891725), .Z(n_242169433)
		);
	notech_or2 i_47850194(.A(n_289127273), .B(n_309891725), .Z(n_243069442)
		);
	notech_or2 i_48750185(.A(n_289027272), .B(n_309891725), .Z(n_243969451)
		);
	notech_or2 i_49650176(.A(n_309891725), .B(n_288927271), .Z(n_244869460)
		);
	notech_nor2 i_62350056(.A(n_57869), .B(\nbus_11365[25] ), .Z(n_244969461
		));
	notech_or2 i_61850061(.A(n_321538010), .B(n_288927271), .Z(n_245669468)
		);
	notech_or2 i_65950020(.A(n_154331958), .B(nbus_11295[25]), .Z(n_245769469
		));
	notech_or2 i_65850021(.A(n_57870), .B(\nbus_11365[25] ), .Z(n_246069472)
		);
	notech_or2 i_65350026(.A(n_305924323), .B(n_288927271), .Z(n_246569477)
		);
	notech_nor2 i_75849928(.A(n_314047718), .B(\nbus_11365[25] ), .Z(n_246669478
		));
	notech_or2 i_75349933(.A(n_306824332), .B(n_288927271), .Z(n_247369485)
		);
	notech_ao3 i_82549862(.A(n_32304), .B(opd[25]), .C(n_56688), .Z(n_247469486
		));
	notech_nand2 i_82049867(.A(\regs_13_14[25] ), .B(n_287027252), .Z(n_248169493
		));
	notech_ao3 i_84749840(.A(n_60338), .B(opb[22]), .C(n_30822), .Z(n_248569497
		));
	notech_nor2 i_86049827(.A(n_304691777), .B(\nbus_11358[23] ), .Z(n_248969501
		));
	notech_ao3 i_87349814(.A(n_60338), .B(opb[24]), .C(n_30822), .Z(n_249369505
		));
	notech_or2 i_88549804(.A(n_57867), .B(\nbus_11365[25] ), .Z(n_249469506)
		);
	notech_or2 i_88449805(.A(n_57865), .B(\nbus_11358[25] ), .Z(n_249769509)
		);
	notech_or2 i_87949810(.A(n_305624320), .B(n_288927271), .Z(n_250269514)
		);
	notech_nor2 i_88849801(.A(n_304691777), .B(\nbus_11358[25] ), .Z(n_250669518
		));
	notech_or2 i_100249689(.A(n_308991734), .B(\nbus_11365[25] ), .Z(n_250969521
		));
	notech_or2 i_99949692(.A(n_122428501), .B(n_28151), .Z(n_251269524));
	notech_nao3 i_99649695(.A(n_19065), .B(read_data[25]), .C(n_59100), .Z(n_251569527
		));
	notech_nand2 i_99349698(.A(add_len_pc[25]), .B(n_26766), .Z(n_251869530)
		);
	notech_nand2 i_41050664(.A(opc[25]), .B(n_62824), .Z(n_253569547));
	notech_ao4 i_191148803(.A(n_56547), .B(n_28586), .C(n_26651), .D(n_28183
		), .Z(n_253669548));
	notech_ao4 i_191048804(.A(n_27036), .B(n_28553), .C(n_56557), .D(n_27887
		), .Z(n_253769549));
	notech_ao4 i_190848806(.A(n_56605), .B(n_28476), .C(n_56583), .D(n_28509
		), .Z(n_253969551));
	notech_ao4 i_190748807(.A(n_56630), .B(n_28444), .C(n_56619), .D(n_28412
		), .Z(n_254069552));
	notech_and4 i_191348801(.A(n_254069552), .B(n_253969551), .C(n_253769549
		), .D(n_253669548), .Z(n_254269554));
	notech_ao4 i_190448810(.A(n_26920), .B(n_28380), .C(n_56489), .D(n_28348
		), .Z(n_254369555));
	notech_ao4 i_190348811(.A(n_26927), .B(n_28315), .C(n_26649), .D(n_29887
		), .Z(n_254469556));
	notech_and2 i_190548809(.A(n_254469556), .B(n_254369555), .Z(n_254569557
		));
	notech_ao4 i_190148813(.A(n_56919), .B(n_29886), .C(n_56640), .D(n_28282
		), .Z(n_254669558));
	notech_ao4 i_190048814(.A(n_26924), .B(n_28250), .C(n_56653), .D(n_28215
		), .Z(n_254769559));
	notech_ao4 i_189748817(.A(n_124328520), .B(n_288927271), .C(n_309391730)
		, .D(n_253569547), .Z(n_255069562));
	notech_ao4 i_189548819(.A(n_121628493), .B(n_28010), .C(n_60144), .D(n_27267
		), .Z(n_255269564));
	notech_and4 i_189948815(.A(n_255269564), .B(n_255069562), .C(n_251869530
		), .D(n_251569527), .Z(n_255469566));
	notech_ao4 i_189248822(.A(n_26765), .B(n_29770), .C(n_309191732), .D(n_29885
		), .Z(n_255569567));
	notech_ao4 i_189048824(.A(n_309091733), .B(\nbus_11358[25] ), .C(n_122528502
		), .D(n_60000), .Z(n_255769569));
	notech_and4 i_189448820(.A(n_255769569), .B(n_255569567), .C(n_250969521
		), .D(n_251269524), .Z(n_255969571));
	notech_nand2 i_2550668(.A(opc_10[25]), .B(n_62824), .Z(n_256069572));
	notech_ao4 i_179548913(.A(n_58007), .B(n_256069572), .C(n_58008), .D(n_253569547
		), .Z(n_256169573));
	notech_ao4 i_179448914(.A(n_26937), .B(n_29770), .C(n_58423), .D(n_28010
		), .Z(n_256369575));
	notech_ao4 i_179148917(.A(n_58138), .B(n_60000), .C(n_57726), .D(n_28151
		), .Z(n_256569577));
	notech_ao4 i_179948909(.A(n_30803), .B(n_60000), .C(n_309591728), .D(n_29770
		), .Z(n_256769579));
	notech_ao4 i_179848910(.A(n_28114), .B(n_60338), .C(n_309491729), .D(\nbus_11365[25] 
		), .Z(n_256969581));
	notech_nao3 i_68150659(.A(n_256769579), .B(n_256969581), .C(n_250669518)
		, .Z(n_257069582));
	notech_and4 i_179348915(.A(n_256569577), .B(n_249469506), .C(n_249769509
		), .D(n_26575), .Z(n_257269584));
	notech_ao4 i_178848920(.A(n_60001), .B(n_30803), .C(n_309591728), .D(n_29769
		), .Z(n_257369585));
	notech_ao4 i_178748921(.A(n_28113), .B(n_60338), .C(n_309491729), .D(\nbus_11365[24] 
		), .Z(n_257569587));
	notech_nao3 i_68050660(.A(n_257369585), .B(n_257569587), .C(n_249369505)
		, .Z(n_257669588));
	notech_ao4 i_177748931(.A(n_60002), .B(n_30803), .C(n_309591728), .D(n_29765
		), .Z(n_257769589));
	notech_ao4 i_177648932(.A(n_28112), .B(n_60338), .C(n_309491729), .D(\nbus_11365[23] 
		), .Z(n_257969591));
	notech_nao3 i_67950661(.A(n_257769589), .B(n_257969591), .C(n_248969501)
		, .Z(n_258069592));
	notech_ao4 i_176548942(.A(n_60003), .B(n_30803), .C(n_309591728), .D(n_29708
		), .Z(n_258169593));
	notech_ao4 i_176448943(.A(n_28111), .B(n_60338), .C(n_309491729), .D(\nbus_11365[22] 
		), .Z(n_258369595));
	notech_nao3 i_67850662(.A(n_258169593), .B(n_258369595), .C(n_248569497)
		, .Z(n_258469596));
	notech_ao4 i_174448963(.A(n_253569547), .B(n_286927251), .C(n_256069572)
		, .D(n_286827250), .Z(n_258569597));
	notech_ao4 i_174348964(.A(n_57861), .B(\nbus_11365[25] ), .C(n_287827260
		), .D(n_288927271), .Z(n_258769599));
	notech_nand3 i_174648961(.A(n_258569597), .B(n_258769599), .C(n_248169493
		), .Z(n_258869600));
	notech_ao4 i_174148966(.A(n_58139), .B(n_60000), .C(n_57863), .D(\nbus_11358[25] 
		), .Z(n_258969601));
	notech_ao4 i_163249074(.A(n_306624330), .B(n_256069572), .C(n_307124335)
		, .D(n_253569547), .Z(n_259269604));
	notech_ao4 i_163149075(.A(n_307324337), .B(n_29770), .C(n_58425), .D(n_28010
		), .Z(n_259469606));
	notech_nand3 i_163449072(.A(n_259269604), .B(n_259469606), .C(n_247369485
		), .Z(n_259569607));
	notech_ao4 i_162949077(.A(n_57864), .B(\nbus_11358[25] ), .C(n_58141), .D
		(n_60000), .Z(n_259669608));
	notech_ao4 i_155649149(.A(n_306124325), .B(n_256069572), .C(n_58085), .D
		(n_253569547), .Z(n_259969611));
	notech_ao4 i_155549150(.A(n_26902), .B(n_29770), .C(n_58427), .D(n_28010
		), .Z(n_260169613));
	notech_ao4 i_155249153(.A(n_57877), .B(\nbus_11358[25] ), .C(n_58143), .D
		(n_60000), .Z(n_260369615));
	notech_and4 i_155449151(.A(n_260369615), .B(n_245769469), .C(n_26575), .D
		(n_246069472), .Z(n_260669618));
	notech_ao4 i_152349181(.A(n_256069572), .B(n_319937994), .C(n_58082), .D
		(n_253569547), .Z(n_260769619));
	notech_ao4 i_152249182(.A(n_26918), .B(n_29770), .C(n_321438009), .D(n_28010
		), .Z(n_260969621));
	notech_nand3 i_152549179(.A(n_260769619), .B(n_260969621), .C(n_245669468
		), .Z(n_261069622));
	notech_ao4 i_152049184(.A(n_57873), .B(\nbus_11358[25] ), .C(n_58145), .D
		(n_60000), .Z(n_261169623));
	notech_ao4 i_142849272(.A(n_295269964), .B(n_256069572), .C(n_253569547)
		, .D(n_26595), .Z(n_261469626));
	notech_ao4 i_142749273(.A(n_308091743), .B(n_28114), .C(n_4014), .D(n_28010
		), .Z(n_261669628));
	notech_and3 i_143049270(.A(n_261469626), .B(n_261669628), .C(n_244869460
		), .Z(n_261769629));
	notech_ao4 i_142449275(.A(n_143028707), .B(n_60000), .C(n_142928706), .D
		(n_29770), .Z(n_261869630));
	notech_ao4 i_142349276(.A(n_142728704), .B(\nbus_11365[25] ), .C(n_142828705
		), .D(\nbus_11358[25] ), .Z(n_261969631));
	notech_ao4 i_142049279(.A(n_225565784), .B(n_295269964), .C(n_221065739)
		, .D(n_26595), .Z(n_262169633));
	notech_ao4 i_141949280(.A(n_308091743), .B(n_28113), .C(n_4014), .D(n_28009
		), .Z(n_262369635));
	notech_and3 i_142249277(.A(n_262169633), .B(n_262369635), .C(n_243969451
		), .Z(n_262469636));
	notech_ao4 i_141749282(.A(n_60001), .B(n_143028707), .C(n_142928706), .D
		(n_29769), .Z(n_262569637));
	notech_ao4 i_141649283(.A(n_142728704), .B(\nbus_11365[24] ), .C(n_142828705
		), .D(\nbus_11358[24] ), .Z(n_262669638));
	notech_ao4 i_141349286(.A(n_225665785), .B(n_295269964), .C(n_222565754)
		, .D(n_26595), .Z(n_262869640));
	notech_ao4 i_141249287(.A(n_308091743), .B(n_28112), .C(n_4014), .D(n_28008
		), .Z(n_263069642));
	notech_and3 i_141549284(.A(n_262869640), .B(n_263069642), .C(n_243069442
		), .Z(n_263169643));
	notech_ao4 i_141049289(.A(n_60002), .B(n_143028707), .C(n_142928706), .D
		(n_29765), .Z(n_263269644));
	notech_ao4 i_140949290(.A(n_142728704), .B(\nbus_11365[23] ), .C(n_142828705
		), .D(\nbus_11358[23] ), .Z(n_263369645));
	notech_ao4 i_140649293(.A(n_225765786), .B(n_295269964), .C(n_224065769)
		, .D(n_26595), .Z(n_263569647));
	notech_ao4 i_140549294(.A(n_308091743), .B(n_28111), .C(n_4014), .D(n_28007
		), .Z(n_263769649));
	notech_and3 i_140849291(.A(n_263569647), .B(n_263769649), .C(n_242169433
		), .Z(n_263869650));
	notech_ao4 i_140349296(.A(n_60003), .B(n_143028707), .C(n_142928706), .D
		(n_29708), .Z(n_263969651));
	notech_ao4 i_140249297(.A(n_142728704), .B(\nbus_11365[22] ), .C(n_142828705
		), .D(\nbus_11358[22] ), .Z(n_264069652));
	notech_ao4 i_139949300(.A(n_27329), .B(n_256069572), .C(n_253569547), .D
		(n_26803), .Z(n_264269654));
	notech_ao4 i_139749302(.A(n_27319), .B(n_28010), .C(n_60148), .D(n_27214
		), .Z(n_264469656));
	notech_and4 i_140149298(.A(n_264469656), .B(n_264269654), .C(n_240969421
		), .D(n_241269424), .Z(n_264669658));
	notech_ao4 i_139449305(.A(n_145128728), .B(n_60000), .C(n_145028727), .D
		(n_29770), .Z(n_264769659));
	notech_ao4 i_139249307(.A(n_27335), .B(n_29884), .C(n_144828725), .D(\nbus_11365[25] 
		), .Z(n_264969661));
	notech_and4 i_139649303(.A(n_264969661), .B(n_264769659), .C(n_240369415
		), .D(n_240669418), .Z(n_265169663));
	notech_mux2 i_136149338(.S(n_32318), .A(n_312147737), .B(n_344466973), .Z
		(n_265269664));
	notech_ao4 i_135849341(.A(n_300891815), .B(n_229269304), .C(n_229169303)
		, .D(n_184068857), .Z(n_265369665));
	notech_ao4 i_135749342(.A(n_152472004), .B(n_185068867), .C(n_152572005)
		, .D(n_117968196), .Z(n_265469666));
	notech_ao4 i_135549344(.A(n_59991), .B(n_303691787), .C(n_58316), .D(n_297369985
		), .Z(n_265669668));
	notech_and4 i_136049339(.A(n_265669668), .B(n_265469666), .C(n_265369665
		), .D(n_239469406), .Z(n_265869670));
	notech_ao4 i_135249347(.A(n_297469986), .B(\nbus_11358[2] ), .C(n_58383)
		, .D(n_27984), .Z(n_265969671));
	notech_ao4 i_135149348(.A(n_344366972), .B(n_274369755), .C(n_297569987)
		, .D(n_57557), .Z(n_266069672));
	notech_ao4 i_134949350(.A(n_27334), .B(n_29883), .C(n_27335), .D(n_29882
		), .Z(n_266269674));
	notech_and3 i_135049349(.A(n_230865837), .B(n_266269674), .C(n_208365612
		), .Z(n_266369675));
	notech_ao4 i_134649353(.A(n_151931934), .B(n_256069572), .C(n_58084), .D
		(n_253569547), .Z(n_266569677));
	notech_ao4 i_134549354(.A(n_29770), .B(n_26929), .C(n_58429), .D(n_28010
		), .Z(n_266769679));
	notech_nand3 i_134849351(.A(n_266569677), .B(n_266769679), .C(n_238569397
		), .Z(n_266869680));
	notech_ao4 i_134349356(.A(n_57875), .B(\nbus_11358[25] ), .C(n_58147), .D
		(n_60000), .Z(n_266969681));
	notech_ao4 i_124849451(.A(n_3843), .B(n_256069572), .C(n_3858), .D(n_253569547
		), .Z(n_267269684));
	notech_ao4 i_124749452(.A(n_26642), .B(n_29770), .C(n_3857), .D(n_28010)
		, .Z(n_267469686));
	notech_nand3 i_125049449(.A(n_267269684), .B(n_267469686), .C(n_237769389
		), .Z(n_267569687));
	notech_ao4 i_124549454(.A(n_3877), .B(\nbus_11358[25] ), .C(n_148228759)
		, .D(n_60000), .Z(n_267669688));
	notech_ao4 i_124149458(.A(n_225565784), .B(n_3843), .C(n_221065739), .D(n_3858
		), .Z(n_267969691));
	notech_ao4 i_124049459(.A(n_29769), .B(n_26642), .C(n_3857), .D(n_28009)
		, .Z(n_268169693));
	notech_ao4 i_123749462(.A(n_3877), .B(\nbus_11358[24] ), .C(n_60001), .D
		(n_148228759), .Z(n_268369695));
	notech_and4 i_123949460(.A(n_125828535), .B(n_268369695), .C(n_236469376
		), .D(n_26619), .Z(n_268669698));
	notech_ao4 i_120749492(.A(n_310891715), .B(n_253569547), .C(n_310791716)
		, .D(n_256069572), .Z(n_268769699));
	notech_ao4 i_120649493(.A(n_149328770), .B(\nbus_11365[25] ), .C(n_149428771
		), .D(\nbus_11358[25] ), .Z(n_268969701));
	notech_and3 i_120949490(.A(n_268769699), .B(n_268969701), .C(n_236169373
		), .Z(n_269069702));
	notech_ao4 i_120349496(.A(n_149128768), .B(n_60000), .C(n_149228769), .D
		(n_29770), .Z(n_269169703));
	notech_ao4 i_120249497(.A(n_28114), .B(n_60338), .C(n_54643), .D(n_28979
		), .Z(n_269369705));
	notech_mux2 i_117349524(.S(n_32341), .A(n_312147737), .B(n_344466973), .Z
		(n_269569707));
	notech_mux2 i_117249525(.S(n_32341), .A(n_312347735), .B(n_312447734), .Z
		(n_269669708));
	notech_ao4 i_116949528(.A(n_306070071), .B(n_229069302), .C(n_24994), .D
		(n_228969301), .Z(n_269769709));
	notech_ao4 i_116749530(.A(n_26697), .B(n_58316), .C(n_152472004), .D(n_306170072
		), .Z(n_269969711));
	notech_and4 i_117149526(.A(n_269969711), .B(n_269769709), .C(n_234569357
		), .D(n_234869360), .Z(n_270169713));
	notech_ao4 i_116449533(.A(n_57882), .B(\nbus_11358[2] ), .C(n_27984), .D
		(n_58410), .Z(n_270269714));
	notech_ao4 i_116249535(.A(n_54643), .B(n_28964), .C(n_344366972), .D(n_306270073
		), .Z(n_270469716));
	notech_and3 i_116349534(.A(n_138971869), .B(n_143671916), .C(n_270469716
		), .Z(n_270569717));
	notech_ao4 i_115949538(.A(n_308791736), .B(n_256069572), .C(n_307891745)
		, .D(n_253569547), .Z(n_270769719));
	notech_ao4 i_115749540(.A(n_308591738), .B(n_28010), .C(n_60148), .D(n_27148
		), .Z(n_270969721));
	notech_and4 i_116149536(.A(n_270969721), .B(n_270769719), .C(n_233469346
		), .D(n_233769349), .Z(n_271169723));
	notech_ao4 i_115449543(.A(n_150728784), .B(n_60000), .C(n_150628783), .D
		(n_29770), .Z(n_271269724));
	notech_ao4 i_115349544(.A(n_29881), .B(n_26648), .C(n_150428781), .D(\nbus_11365[25] 
		), .Z(n_271469726));
	notech_ao4 i_110449591(.A(n_311391710), .B(n_256069572), .C(n_311491709)
		, .D(n_253569547), .Z(n_271669728));
	notech_ao4 i_110249593(.A(n_29770), .B(n_26696), .C(n_311291711), .D(n_28010
		), .Z(n_271869730));
	notech_and4 i_110649589(.A(n_271869730), .B(n_271669728), .C(n_232369335
		), .D(n_232669338), .Z(n_272069732));
	notech_ao4 i_109949596(.A(n_311091713), .B(n_57771), .C(n_311191712), .D
		(n_55965), .Z(n_272169733));
	notech_nand2 i_110049595(.A(n_272169733), .B(n_232069332), .Z(n_272269734
		));
	notech_ao4 i_108649609(.A(n_225665785), .B(n_311391710), .C(n_222565754)
		, .D(n_311491709), .Z(n_272569737));
	notech_ao4 i_108449611(.A(n_29765), .B(n_26696), .C(n_311291711), .D(n_28008
		), .Z(n_272769739));
	notech_and4 i_108849607(.A(n_272769739), .B(n_272569737), .C(n_231369325
		), .D(n_231669328), .Z(n_272969741));
	notech_ao4 i_108149614(.A(n_311091713), .B(\nbus_11365[23] ), .C(n_311191712
		), .D(\nbus_11358[23] ), .Z(n_273069742));
	notech_nand2 i_108249613(.A(n_273069742), .B(n_231069322), .Z(n_273169743
		));
	notech_ao4 i_107749618(.A(n_225765786), .B(n_311391710), .C(n_224065769)
		, .D(n_311491709), .Z(n_273469746));
	notech_ao4 i_107449620(.A(n_29708), .B(n_26696), .C(n_311291711), .D(n_28007
		), .Z(n_273669748));
	notech_and4 i_107949616(.A(n_273669748), .B(n_273469746), .C(n_230369315
		), .D(n_230669318), .Z(n_273869750));
	notech_ao4 i_107049623(.A(n_311091713), .B(\nbus_11365[22] ), .C(n_311191712
		), .D(\nbus_11358[22] ), .Z(n_273969751));
	notech_nand2 i_107149622(.A(n_273969751), .B(n_230069312), .Z(n_274069752
		));
	notech_or4 i_125358525(.A(n_300891815), .B(instrc[116]), .C(n_29658), .D
		(n_26770), .Z(n_274369755));
	notech_ao4 i_8347616(.A(n_60009), .B(n_26815), .C(n_29710), .D(n_313491689
		), .Z(n_274469756));
	notech_and3 i_8447615(.A(n_27348), .B(n_274369755), .C(n_276769779), .Z(n_274569757
		));
	notech_and2 i_8247617(.A(n_288869900), .B(n_275169763), .Z(n_275069762)
		);
	notech_or2 i_51847194(.A(n_313747721), .B(n_4011), .Z(n_275169763));
	notech_nand3 i_44947262(.A(n_60148), .B(n_60241), .C(read_data[16]), .Z(n_275969771
		));
	notech_or2 i_44647265(.A(n_313747721), .B(n_144428721), .Z(n_276269774)
		);
	notech_or4 i_45447257(.A(n_27346), .B(instrc[116]), .C(n_29658), .D(n_26770
		), .Z(n_276769779));
	notech_or4 i_51047201(.A(n_62858), .B(n_304991774), .C(n_62788), .D(\nbus_11365[16] 
		), .Z(n_277669788));
	notech_or2 i_52747186(.A(n_142828705), .B(\nbus_11358[17] ), .Z(n_278169793
		));
	notech_or4 i_52247191(.A(n_62858), .B(n_304991774), .C(n_62814), .D(\nbus_11365[17] 
		), .Z(n_278669798));
	notech_or2 i_53947176(.A(n_142828705), .B(\nbus_11358[18] ), .Z(n_279169803
		));
	notech_or4 i_53347181(.A(n_62858), .B(n_304991774), .C(n_62824), .D(\nbus_11365[18] 
		), .Z(n_279669808));
	notech_or2 i_54947166(.A(n_142828705), .B(\nbus_11358[19] ), .Z(n_280169813
		));
	notech_or4 i_54447171(.A(n_62858), .B(n_304991774), .C(n_62814), .D(\nbus_11365[19] 
		), .Z(n_280669818));
	notech_or4 i_55747161(.A(n_304991774), .B(nbus_11295[20]), .C(n_60940), 
		.D(n_26601), .Z(n_281569827));
	notech_or2 i_65847061(.A(n_138168398), .B(\nbus_11365[18] ), .Z(n_281669828
		));
	notech_or4 i_65747062(.A(n_58133), .B(n_58497), .C(n_56428), .D(\nbus_11358[18] 
		), .Z(n_281969831));
	notech_nao3 i_65247067(.A(n_62826), .B(opc_10[18]), .C(n_319937994), .Z(n_282469836
		));
	notech_or2 i_71947004(.A(n_154331958), .B(nbus_11295[19]), .Z(n_282569837
		));
	notech_or4 i_71847005(.A(n_56832), .B(n_56939), .C(n_56919), .D(n_28004)
		, .Z(n_282869840));
	notech_or2 i_71547008(.A(n_60006), .B(n_58143), .Z(n_283169843));
	notech_or2 i_71247011(.A(n_286869880), .B(\nbus_11365[19] ), .Z(n_283469846
		));
	notech_or2 i_72846995(.A(n_154331958), .B(nbus_11295[20]), .Z(n_283569847
		));
	notech_or4 i_72746996(.A(n_56832), .B(n_56939), .C(n_56919), .D(n_28005)
		, .Z(n_283869850));
	notech_or4 i_72247001(.A(n_58806), .B(n_58493), .C(nbus_11295[20]), .D(n_60938
		), .Z(n_284369855));
	notech_nor2 i_84346881(.A(n_57861), .B(\nbus_11365[17] ), .Z(n_284469856
		));
	notech_or2 i_83846886(.A(n_313647722), .B(n_287827260), .Z(n_285169863)
		);
	notech_nor2 i_92446808(.A(n_304691777), .B(\nbus_11358[17] ), .Z(n_285569867
		));
	notech_ao3 i_93746795(.A(n_60338), .B(opb[18]), .C(n_30822), .Z(n_285969871
		));
	notech_ao3 i_95046782(.A(n_60338), .B(opb[19]), .C(n_30822), .Z(n_286369875
		));
	notech_ao3 i_96446769(.A(n_60338), .B(opb[20]), .C(n_30822), .Z(n_286769879
		));
	notech_nand2 i_4947650(.A(n_26800), .B(n_26824), .Z(n_286869880));
	notech_ao4 i_216545618(.A(n_27761), .B(n_27746), .C(n_58319), .D(eval_flag
		), .Z(n_287069882));
	notech_ao4 i_199045792(.A(n_60005), .B(n_30803), .C(n_309591728), .D(n_29775
		), .Z(n_287269884));
	notech_ao4 i_198945793(.A(n_28109), .B(n_60340), .C(n_309491729), .D(\nbus_11365[20] 
		), .Z(n_287469886));
	notech_nao3 i_67647689(.A(n_287269884), .B(n_287469886), .C(n_286769879)
		, .Z(n_287569887));
	notech_ao4 i_197945803(.A(n_60006), .B(n_30803), .C(n_309591728), .D(n_29773
		), .Z(n_287669888));
	notech_ao4 i_197845804(.A(n_28108), .B(n_60331), .C(n_309491729), .D(\nbus_11365[19] 
		), .Z(n_287869890));
	notech_nao3 i_67547690(.A(n_287669888), .B(n_287869890), .C(n_286369875)
		, .Z(n_287969891));
	notech_ao4 i_196645814(.A(n_3864), .B(n_30803), .C(n_309591728), .D(n_29711
		), .Z(n_288069892));
	notech_ao4 i_196545815(.A(n_28107), .B(n_60331), .C(n_309491729), .D(\nbus_11365[18] 
		), .Z(n_288269894));
	notech_nao3 i_67447691(.A(n_288069892), .B(n_288269894), .C(n_285969871)
		, .Z(n_288369895));
	notech_ao4 i_195545825(.A(n_60008), .B(n_30803), .C(n_29772), .D(n_309591728
		), .Z(n_288469896));
	notech_ao4 i_195445826(.A(n_28106), .B(n_60331), .C(n_309491729), .D(\nbus_11365[17] 
		), .Z(n_288669898));
	notech_nao3 i_67347692(.A(n_288469896), .B(n_288669898), .C(n_285569867)
		, .Z(n_288769899));
	notech_ao4 i_4447655(.A(n_56688), .B(n_28001), .C(n_313747721), .D(n_32348
		), .Z(n_288869900));
	notech_ao4 i_183245931(.A(n_249672976), .B(n_286827250), .C(n_245572935)
		, .D(n_286927251), .Z(n_288969901));
	notech_ao4 i_183145932(.A(n_29772), .B(n_26615), .C(n_58424), .D(n_28002
		), .Z(n_289169903));
	notech_nand3 i_183445929(.A(n_285169863), .B(n_288969901), .C(n_289169903
		), .Z(n_289269904));
	notech_ao4 i_182945934(.A(n_57863), .B(\nbus_11358[17] ), .C(n_60008), .D
		(n_58139), .Z(n_289369905));
	notech_ao4 i_173046030(.A(n_247072950), .B(n_306124325), .C(n_313347725)
		, .D(n_305924323), .Z(n_289669908));
	notech_ao4 i_172946031(.A(n_29775), .B(n_26902), .C(n_60005), .D(n_58143
		), .Z(n_289869910));
	notech_ao4 i_172646034(.A(n_57877), .B(\nbus_11358[20] ), .C(n_57870), .D
		(\nbus_11365[20] ), .Z(n_290069912));
	notech_and4 i_172846032(.A(n_283869850), .B(n_290069912), .C(n_283569847
		), .D(n_26623), .Z(n_290369915));
	notech_ao4 i_172246038(.A(n_247972959), .B(n_306124325), .C(n_313447724)
		, .D(n_305924323), .Z(n_290469916));
	notech_ao4 i_172046040(.A(n_243072910), .B(n_58085), .C(n_253773017), .D
		(n_58493), .Z(n_290669918));
	notech_and4 i_172446036(.A(n_290669918), .B(n_290469916), .C(n_283169843
		), .D(n_283469846), .Z(n_290869920));
	notech_ao4 i_171746043(.A(n_57877), .B(\nbus_11358[19] ), .C(n_29773), .D
		(n_26902), .Z(n_290969921));
	notech_and4 i_171946041(.A(n_282869840), .B(n_290969921), .C(n_26622), .D
		(n_282569837), .Z(n_291269924));
	notech_ao4 i_166946089(.A(n_95222216), .B(n_58082), .C(n_60121865), .D(n_58497
		), .Z(n_291369925));
	notech_ao4 i_166846090(.A(n_321438009), .B(n_28003), .C(n_3861), .D(n_321538010
		), .Z(n_291569927));
	notech_ao4 i_166546093(.A(n_3864), .B(n_58145), .C(n_29711), .D(n_26918)
		, .Z(n_291769929));
	notech_and4 i_166746091(.A(n_291769929), .B(n_26621), .C(n_281669828), .D
		(n_281969831), .Z(n_292069932));
	notech_ao4 i_158746168(.A(n_247072950), .B(n_295269964), .C(n_313347725)
		, .D(n_309891725), .Z(n_292169933));
	notech_ao4 i_158646169(.A(n_60005), .B(n_143028707), .C(n_29775), .D(n_142928706
		), .Z(n_292369935));
	notech_and3 i_158946166(.A(n_292169933), .B(n_292369935), .C(n_281569827
		), .Z(n_292469936));
	notech_ao4 i_158446171(.A(n_142728704), .B(\nbus_11365[20] ), .C(n_142828705
		), .D(\nbus_11358[20] ), .Z(n_292569937));
	notech_ao4 i_158346172(.A(n_308091743), .B(n_28109), .C(n_4014), .D(n_28005
		), .Z(n_292669938));
	notech_ao4 i_158046175(.A(n_247972959), .B(n_295269964), .C(n_313447724)
		, .D(n_309891725), .Z(n_292869940));
	notech_ao4 i_157946176(.A(n_142928706), .B(n_29773), .C(n_243072910), .D
		(n_26595), .Z(n_293069942));
	notech_and3 i_158246173(.A(n_292869940), .B(n_293069942), .C(n_280669818
		), .Z(n_293169943));
	notech_ao4 i_157546179(.A(n_57935), .B(\nbus_11365[19] ), .C(n_60006), .D
		(n_143028707), .Z(n_293269944));
	notech_ao4 i_157446180(.A(n_308091743), .B(n_28108), .C(n_4014), .D(n_28004
		), .Z(n_293469946));
	notech_ao4 i_157146183(.A(n_77522039), .B(n_295269964), .C(n_3861), .D(n_309891725
		), .Z(n_293669948));
	notech_ao4 i_157046184(.A(n_142928706), .B(n_29711), .C(n_95222216), .D(n_26595
		), .Z(n_293869950));
	notech_and3 i_157346181(.A(n_293669948), .B(n_293869950), .C(n_279669808
		), .Z(n_293969951));
	notech_ao4 i_156746187(.A(n_57935), .B(\nbus_11365[18] ), .C(n_3864), .D
		(n_143028707), .Z(n_294069952));
	notech_ao4 i_156646188(.A(n_55726), .B(n_28107), .C(n_4014), .D(n_28003)
		, .Z(n_294269954));
	notech_ao4 i_156346191(.A(n_249672976), .B(n_295269964), .C(n_313647722)
		, .D(n_309891725), .Z(n_294469956));
	notech_ao4 i_156246192(.A(n_142928706), .B(n_29772), .C(n_245572935), .D
		(n_26595), .Z(n_294669958));
	notech_ao4 i_155946195(.A(n_57935), .B(\nbus_11365[17] ), .C(n_60008), .D
		(n_143028707), .Z(n_294869960));
	notech_ao4 i_155846196(.A(n_55726), .B(n_28106), .C(n_4014), .D(n_28002)
		, .Z(n_295069962));
	notech_and3 i_156146193(.A(n_294869960), .B(n_295069962), .C(n_278169793
		), .Z(n_295169963));
	notech_nao3 i_155746197(.A(n_246591944), .B(n_57068), .C(n_184792036), .Z
		(n_295269964));
	notech_ao4 i_155446200(.A(n_26649), .B(n_275069762), .C(n_254466073), .D
		(n_295269964), .Z(n_295369965));
	notech_ao4 i_155346201(.A(n_57935), .B(\nbus_11365[16] ), .C(n_252966058
		), .D(n_26595), .Z(n_295569967));
	notech_and3 i_155646198(.A(n_295369965), .B(n_295569967), .C(n_277669788
		), .Z(n_295669968));
	notech_ao4 i_155146203(.A(n_60009), .B(n_298469996), .C(n_29710), .D(n_142928706
		), .Z(n_295769969));
	notech_ao4 i_155046204(.A(n_55726), .B(n_28105), .C(n_142828705), .D(\nbus_11358[16] 
		), .Z(n_295869970));
	notech_ao4 i_150146251(.A(n_254466073), .B(n_274569757), .C(n_274469756)
		, .D(n_184892035), .Z(n_296169973));
	notech_ao4 i_150046252(.A(n_57160), .B(\nbus_11365[16] ), .C(n_144928726
		), .D(\nbus_11358[16] ), .Z(n_296269974));
	notech_ao4 i_149846254(.A(n_312324377), .B(n_303791786), .C(n_252966058)
		, .D(n_26803), .Z(n_296469976));
	notech_and4 i_150346249(.A(n_296469976), .B(n_296269974), .C(n_296169973
		), .D(n_276269774), .Z(n_296669978));
	notech_ao4 i_149546257(.A(n_27319), .B(n_28001), .C(n_60144), .D(n_27205
		), .Z(n_296769979));
	notech_ao4 i_6147638(.A(n_60009), .B(n_305691767), .C(n_29710), .D(n_305591768
		), .Z(n_296969981));
	notech_ao4 i_149346259(.A(n_27334), .B(n_29889), .C(n_27335), .D(n_29888
		), .Z(n_297069982));
	notech_and4 i_149746255(.A(n_296969981), .B(n_297069982), .C(n_296769979
		), .D(n_275969771), .Z(n_297269984));
	notech_and3 i_85258537(.A(n_303791786), .B(n_27346), .C(n_27349), .Z(n_297369985
		));
	notech_ao4 i_116161805(.A(n_61115), .B(n_27306), .C(n_26815), .D(n_118468201
		), .Z(n_297469986));
	notech_and2 i_116261804(.A(n_298991830), .B(n_118268199), .Z(n_297569987
		));
	notech_nand2 i_14544351(.A(n_27348), .B(n_298269994), .Z(n_297869990));
	notech_and2 i_14644350(.A(n_92619108), .B(n_309370104), .Z(n_297969991)
		);
	notech_nand3 i_52243983(.A(n_27163), .B(n_30946), .C(n_2026), .Z(n_298269994
		));
	notech_and2 i_13544361(.A(n_215576094), .B(n_298769998), .Z(n_298369995)
		);
	notech_and2 i_159647758(.A(n_306691757), .B(n_287069882), .Z(n_298469996
		));
	notech_or2 i_59343916(.A(n_314391680), .B(n_4011), .Z(n_298769998));
	notech_nand3 i_64643870(.A(n_60144), .B(n_60241), .C(read_data[6]), .Z(n_298869999
		));
	notech_nand3 i_124343319(.A(n_60331), .B(n_1901), .C(n_26627), .Z(n_298970000
		));
	notech_nand3 i_125843304(.A(n_57985), .B(n_27221), .C(n_122175165), .Z(n_299070001
		));
	notech_or4 i_125943303(.A(fsm[2]), .B(n_61165), .C(n_61154), .D(n_30470)
		, .Z(n_299170002));
	notech_nand3 i_49144011(.A(n_1429), .B(n_7288), .C(\eflags[10] ), .Z(n_299470005
		));
	notech_nand3 i_50743996(.A(n_1429), .B(n_7292), .C(\eflags[10] ), .Z(n_300970020
		));
	notech_nand3 i_51843986(.A(n_1429), .B(n_7294), .C(\eflags[10] ), .Z(n_302270033
		));
	notech_nand3 i_51743987(.A(n_1429), .B(n_7293), .C(n_29601), .Z(n_302570036
		));
	notech_or4 i_51443990(.A(n_62858), .B(n_184068857), .C(n_60938), .D(n_29723
		), .Z(n_302870039));
	notech_nand3 i_51043993(.A(n_62826), .B(opc[6]), .C(n_297869990), .Z(n_303170042
		));
	notech_nand2 i_9744397(.A(n_26939), .B(n_122175165), .Z(n_305970070));
	notech_nand2 i_35112(.A(n_26939), .B(n_26596), .Z(n_306070071));
	notech_or4 i_7644418(.A(n_57026), .B(n_26697), .C(instrc[119]), .D(n_27712
		), .Z(n_306170072));
	notech_or4 i_8044414(.A(n_57026), .B(instrc[119]), .C(n_27712), .D(n_24994
		), .Z(n_306270073));
	notech_or4 i_71044483(.A(n_60969), .B(n_60958), .C(n_62846), .D(\nbus_11307[3] 
		), .Z(n_306570076));
	notech_nao3 i_70944484(.A(n_62826), .B(opa[3]), .C(n_62846), .Z(n_306670077
		));
	notech_nand2 i_70644486(.A(opc[3]), .B(n_62788), .Z(n_306770078));
	notech_nand2 i_62044488(.A(opc_10[3]), .B(n_62810), .Z(n_306870079));
	notech_or4 i_61344491(.A(n_60970), .B(n_60959), .C(n_62846), .D(n_29728)
		, .Z(n_306970080));
	notech_ao4 i_204042550(.A(n_56547), .B(n_28563), .C(n_29893), .D(n_26649
		), .Z(n_307070081));
	notech_ao4 i_203942551(.A(n_27036), .B(n_28519), .C(n_56557), .D(n_27861
		), .Z(n_307170082));
	notech_ao4 i_203742553(.A(n_26651), .B(n_28161), .C(n_56583), .D(n_28486
		), .Z(n_307370084));
	notech_ao4 i_203642554(.A(n_56619), .B(n_28390), .C(n_56605), .D(n_28454
		), .Z(n_307470085));
	notech_and4 i_204242548(.A(n_307470085), .B(n_307370084), .C(n_307170082
		), .D(n_307070081), .Z(n_307670087));
	notech_ao4 i_203342557(.A(n_56489), .B(n_28325), .C(n_56630), .D(n_28422
		), .Z(n_307770088));
	notech_ao4 i_203242558(.A(n_26927), .B(n_28292), .C(n_26920), .D(n_28358
		), .Z(n_307870089));
	notech_and2 i_203442556(.A(n_307870089), .B(n_307770088), .Z(n_307970090
		));
	notech_ao4 i_203042560(.A(n_56919), .B(n_29892), .C(n_56640), .D(n_28260
		), .Z(n_308070091));
	notech_ao4 i_202942561(.A(n_26924), .B(n_28226), .C(n_56653), .D(n_28193
		), .Z(n_308170092));
	notech_and2 i_8444410(.A(n_306121225), .B(n_298869999), .Z(n_308470095)
		);
	notech_ao4 i_163242955(.A(n_26649), .B(n_298369995), .C(n_83019012), .D(n_295269964
		), .Z(n_308570096));
	notech_ao4 i_163142956(.A(n_142728704), .B(\nbus_11365[31] ), .C(n_96519147
		), .D(n_26595), .Z(n_308670097));
	notech_ao4 i_162942958(.A(n_142828705), .B(\nbus_11358[31] ), .C(n_314791676
		), .D(n_298469996), .Z(n_308870099));
	notech_ao4 i_162842959(.A(n_142928706), .B(n_29619), .C(n_55726), .D(n_28123
		), .Z(n_308970100));
	notech_ao4 i_157843007(.A(\nbus_11358[6] ), .B(n_112664655), .C(\nbus_11307[6] 
		), .D(n_26594), .Z(n_309170102));
	notech_ao4 i_158143004(.A(n_1393), .B(n_29723), .C(n_3874), .D(n_26815),
		 .Z(n_309370104));
	notech_ao4 i_157643009(.A(n_303221196), .B(n_56548), .C(n_300891815), .D
		(n_297969991), .Z(n_309470105));
	notech_and4 i_158043005(.A(n_302870039), .B(n_309470105), .C(n_309170102
		), .D(n_303170042), .Z(n_309670107));
	notech_ao4 i_157343012(.A(n_60144), .B(n_27195), .C(n_92019102), .D(n_274369755
		), .Z(n_309770108));
	notech_and4 i_157543010(.A(n_308470095), .B(n_302570036), .C(n_309770108
		), .D(n_302270033), .Z(n_310070111));
	notech_ao4 i_156943016(.A(n_281966348), .B(n_297369985), .C(n_281866347)
		, .D(n_117968196), .Z(n_310170112));
	notech_ao4 i_156843017(.A(n_282166350), .B(n_274369755), .C(n_282066349)
		, .D(n_185068867), .Z(n_310270113));
	notech_ao4 i_156643019(.A(n_308621250), .B(n_303691787), .C(n_282266351)
		, .D(n_300891815), .Z(n_310470115));
	notech_ao4 i_156543020(.A(n_59326), .B(n_28094), .C(n_60144), .D(n_27193
		), .Z(n_310570116));
	notech_and4 i_157143014(.A(n_310570116), .B(n_310470115), .C(n_310270113
		), .D(n_310170112), .Z(n_310770118));
	notech_ao4 i_156243023(.A(n_297469986), .B(\nbus_11358[5] ), .C(n_58383)
		, .D(n_27987), .Z(n_310870119));
	notech_ao4 i_156143024(.A(n_58001), .B(n_29651), .C(\nbus_11307[5] ), .D
		(n_297569987), .Z(n_310970120));
	notech_ao4 i_155943026(.A(n_27335), .B(n_29891), .C(n_60020), .D(n_58002
		), .Z(n_311170122));
	notech_and4 i_156443021(.A(n_311170122), .B(n_310970120), .C(n_310870119
		), .D(n_300970020), .Z(n_311370124));
	notech_ao4 i_155643029(.A(n_306670077), .B(n_117968196), .C(n_306570076)
		, .D(n_297369985), .Z(n_311470125));
	notech_ao4 i_155543030(.A(n_306870079), .B(n_274369755), .C(n_306770078)
		, .D(n_185068867), .Z(n_311570126));
	notech_ao4 i_155343032(.A(n_308721251), .B(n_303691787), .C(n_300891815)
		, .D(n_306970080), .Z(n_311770128));
	notech_ao4 i_155243033(.A(n_59326), .B(n_28092), .C(n_60144), .D(n_27190
		), .Z(n_311870129));
	notech_and4 i_155843027(.A(n_311870129), .B(n_311770128), .C(n_311570126
		), .D(n_311470125), .Z(n_312070131));
	notech_ao4 i_154943036(.A(n_297469986), .B(\nbus_11358[3] ), .C(n_58383)
		, .D(n_27985), .Z(n_312170132));
	notech_ao4 i_154843037(.A(n_58001), .B(n_29728), .C(n_297569987), .D(\nbus_11307[3] 
		), .Z(n_312270133));
	notech_ao4 i_154643039(.A(n_27335), .B(n_29890), .C(n_60022), .D(n_58002
		), .Z(n_312470135));
	notech_and4 i_155143034(.A(n_312470135), .B(n_312270133), .C(n_312170132
		), .D(n_299470005), .Z(n_312670137));
	notech_nand3 i_88141311(.A(n_39370), .B(n_32341), .C(n_27221), .Z(n_312770138
		));
	notech_nand2 i_167141297(.A(n_26880), .B(n_26938), .Z(n_312870139));
	notech_or4 i_126041264(.A(n_26062), .B(n_57087), .C(n_57068), .D(n_314070151
		), .Z(n_312970140));
	notech_or4 i_126641263(.A(n_57026), .B(instrc[119]), .C(n_27712), .D(n_314170152
		), .Z(n_313070141));
	notech_ao4 i_190941248(.A(n_59445), .B(n_26792), .C(n_209069102), .D(n_26805
		), .Z(n_313170142));
	notech_or2 i_196241247(.A(n_58805), .B(n_314270153), .Z(n_313270143));
	notech_and3 i_61041369(.A(n_311791706), .B(n_310691717), .C(n_321970230)
		, .Z(n_313370144));
	notech_ao4 i_95341370(.A(n_59445), .B(n_26880), .C(n_39370), .D(n_26596)
		, .Z(n_313470145));
	notech_and4 i_101941371(.A(n_59152), .B(n_315391670), .C(n_312770138), .D
		(n_50904), .Z(n_313570146));
	notech_and2 i_121841355(.A(n_52335319), .B(n_102135817), .Z(n_313670147)
		);
	notech_ao4 i_121941356(.A(n_61110), .B(n_30594), .C(n_299691827), .D(n_27349
		), .Z(n_313770148));
	notech_or4 i_115441350(.A(n_308391740), .B(n_306491759), .C(n_304791776)
		, .D(n_48163), .Z(n_313870149));
	notech_ao4 i_122341351(.A(n_32382), .B(n_306291761), .C(n_306891755), .D
		(n_27761), .Z(n_313970150));
	notech_and3 i_79040514(.A(n_23513), .B(n_23514), .C(n_316491659), .Z(n_314070151
		));
	notech_nor2 i_79140513(.A(n_39370), .B(n_26596), .Z(n_314170152));
	notech_nor2 i_79640508(.A(n_209069102), .B(n_26805), .Z(n_314270153));
	notech_or2 i_98240340(.A(n_4011), .B(n_56640), .Z(n_314570156));
	notech_nao3 i_98640336(.A(n_319191632), .B(n_319091633), .C(n_4011), .Z(n_314670157
		));
	notech_or2 i_43340841(.A(n_313570146), .B(\nbus_11358[8] ), .Z(n_314970160
		));
	notech_nand2 i_43240842(.A(opa[8]), .B(n_313470145), .Z(n_315270163));
	notech_nand3 i_42940845(.A(n_26880), .B(n_26938), .C(\opa_12[8] ), .Z(n_315570166
		));
	notech_nao3 i_42640848(.A(n_319091633), .B(n_246991940), .C(n_325270263)
		, .Z(n_315870169));
	notech_nand3 i_50940776(.A(n_1429), .B(n_7298), .C(\eflags[10] ), .Z(n_316170172
		));
	notech_nand2 i_50540779(.A(sav_esi[8]), .B(n_61138), .Z(n_316470175));
	notech_nand2 i_50140782(.A(opb[8]), .B(n_27289), .Z(n_316770178));
	notech_nand2 i_51840767(.A(opd[8]), .B(n_26640), .Z(n_317670187));
	notech_or2 i_51540770(.A(n_313970150), .B(n_29787), .Z(n_317970190));
	notech_or4 i_51240773(.A(n_27761), .B(n_28134), .C(n_60938), .D(n_26601)
		, .Z(n_318270193));
	notech_nao3 i_74740557(.A(n_11415), .B(n_32272), .C(n_2868), .Z(n_318570196
		));
	notech_nand2 i_74440560(.A(sav_epc[12]), .B(n_61138), .Z(n_318870199));
	notech_or4 i_74140563(.A(n_62858), .B(n_62766), .C(n_29679), .D(n_316891655
		), .Z(n_319170202));
	notech_or4 i_36378(.A(n_26062), .B(n_57087), .C(n_57068), .D(n_23512), .Z
		(n_319670207));
	notech_or4 i_35010(.A(n_57026), .B(instrc[119]), .C(n_27712), .D(n_25010
		), .Z(n_319770208));
	notech_or2 i_30197(.A(n_58805), .B(n_58478), .Z(n_319870209));
	notech_nand2 i_30194(.A(n_26792), .B(n_26884), .Z(n_319970210));
	notech_or4 i_28479(.A(n_60970), .B(n_60959), .C(n_62860), .D(n_29679), .Z
		(n_320070211));
	notech_nand2 i_28457(.A(opc_10[12]), .B(n_62782), .Z(n_320170212));
	notech_or4 i_101140321(.A(n_2938), .B(n_2937), .C(n_56832), .D(n_26927),
		 .Z(n_321970230));
	notech_or4 i_101440318(.A(n_2938), .B(n_2937), .C(n_56832), .D(n_56583),
		 .Z(n_322070231));
	notech_ao4 i_200939392(.A(n_59445), .B(n_26829), .C(n_26808), .D(n_26599
		), .Z(n_322670237));
	notech_ao4 i_191739482(.A(n_56557), .B(n_27870), .C(n_56548), .D(n_28573
		), .Z(n_322770238));
	notech_ao4 i_191639483(.A(n_28495), .B(n_56583), .C(n_27036), .D(n_28531
		), .Z(n_322870239));
	notech_ao4 i_191339485(.A(n_56605), .B(n_28463), .C(n_26651), .D(n_28170
		), .Z(n_323070241));
	notech_ao4 i_190839486(.A(n_28431), .B(n_56630), .C(n_56619), .D(n_28399
		), .Z(n_323170242));
	notech_and4 i_191939480(.A(n_323170242), .B(n_323070241), .C(n_322870239
		), .D(n_322770238), .Z(n_323370244));
	notech_ao4 i_190539489(.A(n_26920), .B(n_28367), .C(n_56489), .D(n_28335
		), .Z(n_323470245));
	notech_ao4 i_190439490(.A(n_28302), .B(n_26927), .C(n_26649), .D(n_29898
		), .Z(n_323570246));
	notech_and2 i_190639488(.A(n_323570246), .B(n_323470245), .Z(n_323670247
		));
	notech_ao4 i_190239492(.A(n_56919), .B(n_29896), .C(n_28269), .D(n_56640
		), .Z(n_323770248));
	notech_ao4 i_190139493(.A(n_28237), .B(n_26924), .C(n_28202), .D(n_26922
		), .Z(n_323870249));
	notech_ao4 i_177939610(.A(n_323680737), .B(n_320170212), .C(n_323580736)
		, .D(n_29679), .Z(n_324170252));
	notech_ao4 i_177839611(.A(n_290818107), .B(nbus_11295[12]), .C(n_290718106
		), .D(\nbus_11358[12] ), .Z(n_324270253));
	notech_ao4 i_177639613(.A(n_291718116), .B(n_27997), .C(n_26857), .D(\nbus_11307[12] 
		), .Z(n_324470255));
	notech_and4 i_178139608(.A(n_324470255), .B(n_324270253), .C(n_324170252
		), .D(n_319170202), .Z(n_324670257));
	notech_ao4 i_177339616(.A(n_315591668), .B(n_59965), .C(n_122628503), .D
		(n_29549), .Z(n_324770258));
	notech_ao4 i_177139618(.A(n_309291731), .B(n_28101), .C(n_316791656), .D
		(n_60013), .Z(n_324970260));
	notech_and4 i_177539614(.A(n_318570196), .B(n_324970260), .C(n_324770258
		), .D(n_318870199), .Z(n_325170262));
	notech_or4 i_65441275(.A(calc_sz[1]), .B(n_56834), .C(n_293018129), .D(n_246691943
		), .Z(n_325270263));
	notech_ao4 i_160039783(.A(n_308166610), .B(n_55735), .C(n_325270263), .D
		(n_26649), .Z(n_325370264));
	notech_ao4 i_159839785(.A(\nbus_11307[8] ), .B(n_26598), .C(n_309666625)
		, .D(n_4009), .Z(n_325570266));
	notech_and4 i_160239781(.A(n_325570266), .B(n_325370264), .C(n_317970190
		), .D(n_318270193), .Z(n_325770268));
	notech_ao4 i_159539788(.A(n_55726), .B(n_28097), .C(n_307091753), .D(n_29864
		), .Z(n_325870269));
	notech_ao4 i_159439789(.A(n_5933), .B(n_4007), .C(n_4008), .D(\nbus_11358[8] 
		), .Z(n_326070271));
	notech_ao4 i_159139792(.A(n_308166610), .B(n_27349), .C(n_309666625), .D
		(n_27157), .Z(n_326270273));
	notech_ao4 i_159039793(.A(n_293018129), .B(n_27142), .C(n_27348), .D(n_308066609
		), .Z(n_326370274));
	notech_ao4 i_158839795(.A(n_302691797), .B(\nbus_11307[8] ), .C(n_302591798
		), .D(n_27991), .Z(n_326570276));
	notech_and4 i_159339790(.A(n_326570276), .B(n_326370274), .C(n_326270273
		), .D(n_316770178), .Z(n_326770278));
	notech_ao4 i_158439798(.A(n_313770148), .B(n_29787), .C(n_5933), .D(n_313670147
		), .Z(n_326870279));
	notech_ao4 i_158139800(.A(n_27335), .B(n_29894), .C(n_32270), .D(n_28097
		), .Z(n_327070281));
	notech_and4 i_158739796(.A(n_327070281), .B(n_326870279), .C(n_316170172
		), .D(n_316470175), .Z(n_327270283));
	notech_ao4 i_138439978(.A(n_309666625), .B(n_313070141), .C(n_54643), .D
		(n_28968), .Z(n_327370284));
	notech_ao4 i_138239980(.A(n_308066609), .B(n_319770208), .C(n_308166610)
		, .D(n_25010), .Z(n_327570286));
	notech_and4 i_138639976(.A(n_327570286), .B(n_327370284), .C(n_315570166
		), .D(n_315870169), .Z(n_327770288));
	notech_ao4 i_137939983(.A(n_313370144), .B(n_27991), .C(n_5933), .D(n_312391700
		), .Z(n_327870289));
	notech_and4 i_138139981(.A(n_334480845), .B(n_327870289), .C(n_314970160
		), .D(n_315270163), .Z(n_328170292));
	notech_and2 i_61837648(.A(n_308815164), .B(n_306915145), .Z(n_328270293)
		);
	notech_or2 i_34637898(.A(n_55886), .B(\nbus_11358[28] ), .Z(n_328370294)
		);
	notech_nor2 i_34137903(.A(n_53512635), .B(n_27997), .Z(n_329070301));
	notech_or2 i_33237912(.A(n_3887), .B(n_29064), .Z(n_329970310));
	notech_or2 i_54237724(.A(n_53612636), .B(n_60000), .Z(n_330470315));
	notech_or2 i_53937727(.A(n_54212642), .B(n_57771), .Z(n_330770318));
	notech_ao4 i_205636252(.A(n_27094), .B(n_28422), .C(n_26950), .D(n_28563
		), .Z(n_336070371));
	notech_ao4 i_205536253(.A(n_56909), .B(n_29892), .C(n_56428), .D(n_28358
		), .Z(n_336170372));
	notech_ao4 i_205336255(.A(n_56448), .B(n_28226), .C(n_56437), .D(n_28193
		), .Z(n_336370374));
	notech_ao4 i_205236256(.A(n_56457), .B(n_28260), .C(n_27089), .D(n_28454
		), .Z(n_336470375));
	notech_and4 i_205836250(.A(n_336470375), .B(n_336370374), .C(n_336170372
		), .D(n_336070371), .Z(n_336670377));
	notech_ao4 i_204936259(.A(n_59349), .B(n_28519), .C(n_26664), .D(n_28325
		), .Z(n_336770378));
	notech_ao4 i_204836260(.A(n_56401), .B(n_28161), .C(n_28390), .D(n_56390
		), .Z(n_336870379));
	notech_and2 i_205036258(.A(n_336870379), .B(n_336770378), .Z(n_336970380
		));
	notech_ao4 i_204636262(.A(n_58014), .B(n_27861), .C(n_56468), .D(n_29893
		), .Z(n_337070381));
	notech_ao4 i_204536263(.A(n_28292), .B(n_57985), .C(n_60845), .D(n_28486
		), .Z(n_337170382));
	notech_ao4 i_193036378(.A(n_27094), .B(n_28431), .C(n_26950), .D(n_28573
		), .Z(n_337470385));
	notech_ao4 i_192936379(.A(n_56909), .B(n_29896), .C(n_56428), .D(n_28367
		), .Z(n_337570386));
	notech_ao4 i_192736381(.A(n_56448), .B(n_28237), .C(n_56437), .D(n_28202
		), .Z(n_337770388));
	notech_ao4 i_192636382(.A(n_56457), .B(n_28269), .C(n_27089), .D(n_28463
		), .Z(n_337870389));
	notech_and4 i_193236376(.A(n_337870389), .B(n_337770388), .C(n_337570386
		), .D(n_337470385), .Z(n_338070391));
	notech_ao4 i_192336385(.A(n_59349), .B(n_28531), .C(n_26664), .D(n_28335
		), .Z(n_338170392));
	notech_ao4 i_192236386(.A(n_56401), .B(n_28170), .C(n_56390), .D(n_28399
		), .Z(n_338270393));
	notech_and2 i_192436384(.A(n_338270393), .B(n_338170392), .Z(n_338370394
		));
	notech_ao4 i_192036388(.A(n_58014), .B(n_27870), .C(n_56468), .D(n_29898
		), .Z(n_338470395));
	notech_ao4 i_191936389(.A(n_28302), .B(n_57985), .C(n_27104), .D(n_28495
		), .Z(n_338570396));
	notech_ao4 i_177536532(.A(n_27094), .B(n_28444), .C(n_26950), .D(n_28586
		), .Z(n_338870399));
	notech_ao4 i_177336533(.A(n_56909), .B(n_29886), .C(n_56428), .D(n_28380
		), .Z(n_338970400));
	notech_ao4 i_177136535(.A(n_56448), .B(n_28250), .C(n_56437), .D(n_28215
		), .Z(n_339170402));
	notech_ao4 i_177036536(.A(n_56457), .B(n_28282), .C(n_27089), .D(n_28476
		), .Z(n_339270403));
	notech_and4 i_177736530(.A(n_339270403), .B(n_339170402), .C(n_338970400
		), .D(n_338870399), .Z(n_339470405));
	notech_ao4 i_176736539(.A(n_59349), .B(n_28553), .C(n_26664), .D(n_28348
		), .Z(n_339570406));
	notech_ao4 i_176636540(.A(n_56401), .B(n_28183), .C(n_28412), .D(n_56390
		), .Z(n_339670407));
	notech_and2 i_176836538(.A(n_339670407), .B(n_339570406), .Z(n_339770408
		));
	notech_ao4 i_176436542(.A(n_58014), .B(n_27887), .C(n_56468), .D(n_29887
		), .Z(n_339870409));
	notech_ao4 i_176336543(.A(n_28315), .B(n_57985), .C(n_27104), .D(n_28509
		), .Z(n_339970410));
	notech_ao4 i_163236674(.A(n_276383754), .B(n_29015), .C(n_3888), .D(n_28114
		), .Z(n_340270413));
	notech_ao4 i_163136675(.A(n_310315179), .B(n_55965), .C(n_3887), .D(n_29079
		), .Z(n_340370414));
	notech_ao4 i_162936677(.A(n_54012640), .B(n_29277), .C(n_388360286), .D(nbus_11295
		[25]), .Z(n_340570416));
	notech_and4 i_163436672(.A(n_340570416), .B(n_340370414), .C(n_340270413
		), .D(n_330770318), .Z(n_340770418));
	notech_ao4 i_162636680(.A(n_53412634), .B(n_29628), .C(n_53512635), .D(n_28010
		), .Z(n_340870419));
	notech_ao4 i_162436682(.A(n_3882), .B(n_29243), .C(n_52112621), .D(n_29208
		), .Z(n_341070421));
	notech_and4 i_162836678(.A(n_277183762), .B(n_341070421), .C(n_340870419
		), .D(n_330470315), .Z(n_341270423));
	notech_ao4 i_146336842(.A(n_276383754), .B(n_29014), .C(n_3888), .D(n_28101
		), .Z(n_341370424));
	notech_ao4 i_146236843(.A(n_33412434), .B(n_29190), .C(n_309615172), .D(\nbus_11358[12] 
		), .Z(n_341570426));
	notech_and3 i_146536840(.A(n_341370424), .B(n_341570426), .C(n_329970310
		), .Z(n_341670427));
	notech_ao4 i_146036845(.A(n_33512435), .B(n_28013), .C(n_33312433), .D(n_29013
		), .Z(n_341770428));
	notech_ao4 i_145936846(.A(n_388360286), .B(nbus_11295[12]), .C(n_33012430
		), .D(n_28999), .Z(n_341870429));
	notech_ao4 i_145536850(.A(n_54212642), .B(n_57644), .C(n_54012640), .D(n_29264
		), .Z(n_342170432));
	notech_ao4 i_145436851(.A(n_53612636), .B(n_60013), .C(n_53412634), .D(n_29647
		), .Z(n_342370434));
	notech_ao3 i_145736848(.A(n_342170432), .B(n_342370434), .C(n_329070301)
		, .Z(n_342470435));
	notech_ao4 i_145236853(.A(n_3892), .B(nbus_11295[4]), .C(n_3882), .D(n_29228
		), .Z(n_342570436));
	notech_and2 i_4038194(.A(n_309515171), .B(n_309115167), .Z(n_342670437)
		);
	notech_and4 i_145836847(.A(n_342670437), .B(n_342570436), .C(n_342470435
		), .D(n_328370294), .Z(n_342970440));
	notech_nand3 i_32507(.A(n_246591944), .B(n_57068), .C(n_27061), .Z(n_343270443
		));
	notech_ao4 i_32476(.A(n_27500), .B(n_308012096), .C(n_61110), .D(n_116468181
		), .Z(n_343370444));
	notech_ao4 i_53032297(.A(n_26602), .B(n_343870449), .C(n_2873), .D(n_2872
		), .Z(n_343570446));
	notech_and3 i_53132296(.A(n_27580), .B(n_3925), .C(n_27377), .Z(n_343770448
		));
	notech_and2 i_53232295(.A(n_27377), .B(n_343970450), .Z(n_343870449));
	notech_nand2 i_27332505(.A(n_27714), .B(n_32327), .Z(n_343970450));
	notech_ao3 i_41932382(.A(tsc[27]), .B(n_27855), .C(n_24989), .Z(n_344070451
		));
	notech_or2 i_41832383(.A(n_131228589), .B(n_151428791), .Z(n_344370454)
		);
	notech_or2 i_41532386(.A(n_151028787), .B(nbus_11295[27]), .Z(n_344670457
		));
	notech_or4 i_41232389(.A(nbus_11295[27]), .B(n_60938), .C(n_316491659), 
		.D(n_26942), .Z(n_344970460));
	notech_ao3 i_9732642(.A(n_60329), .B(opa[27]), .C(n_30821), .Z(n_345370464
		));
	notech_ao4 i_101831849(.A(n_60329), .B(n_28116), .C(n_304691777), .D(\nbus_11358[27] 
		), .Z(n_345470465));
	notech_ao4 i_101731850(.A(n_309591728), .B(n_29661), .C(n_131228589), .D
		(n_30803), .Z(n_345670467));
	notech_ao4 i_80932040(.A(n_311391710), .B(n_310091723), .C(n_311291711),
		 .D(n_28012), .Z(n_345770468));
	notech_ao4 i_80732042(.A(n_311091713), .B(\nbus_11365[27] ), .C(n_311191712
		), .D(\nbus_11358[27] ), .Z(n_345970470));
	notech_and4 i_81132038(.A(n_345970470), .B(n_345770468), .C(n_344670457)
		, .D(n_344970460), .Z(n_346170472));
	notech_ao4 i_80332045(.A(n_29661), .B(n_26696), .C(n_151128788), .D(n_4016
		), .Z(n_346270473));
	notech_nand2 i_80432044(.A(n_346270473), .B(n_344370454), .Z(n_346370474
		));
	notech_nand2 i_1318018(.A(n_113368150), .B(n_113268149), .Z(write_data_26
		[12]));
	notech_nand2 i_2618031(.A(n_113568152), .B(n_113468151), .Z(write_data_26
		[25]));
	notech_nand3 i_49004(.A(n_26992), .B(n_114668163), .C(n_115668173), .Z(\nbus_11306[0] 
		));
	notech_or4 i_79864511(.A(n_2985), .B(n_57818), .C(n_61138), .D(n_60234),
		 .Z(n_58219));
	notech_and3 i_123135130(.A(n_32382), .B(n_306391760), .C(n_27896), .Z(n_57818
		));
	notech_nand2 i_49765(.A(n_58219), .B(n_115568172), .Z(n_15649));
	notech_and4 i_56142(.A(n_114368160), .B(n_116968186), .C(n_116268179), .D
		(n_115568172), .Z(\nbus_11376[6] ));
	notech_nand3 i_56141(.A(n_116168178), .B(n_116968186), .C(n_114368160), 
		.Z(\nbus_11376[2] ));
	notech_and4 i_54156(.A(n_252840546), .B(n_117468191), .C(n_146461747), .D
		(n_116068177), .Z(\nbus_11356[8] ));
	notech_and4 i_54155(.A(n_146361746), .B(n_144961732), .C(n_248240500), .D
		(n_117468191), .Z(\nbus_11356[0] ));
	notech_nand3 i_114864492(.A(n_58815), .B(n_254240560), .C(n_62782), .Z(n_57901
		));
	notech_nand2 i_1164439(.A(n_58504), .B(n_58496), .Z(n_254240560));
	notech_or4 i_161264478(.A(n_245362720), .B(n_58480), .C(n_57087), .D(n_57055
		), .Z(n_57473));
	notech_or2 i_37947329(.A(n_310191722), .B(n_27461), .Z(n_239265921));
	notech_and2 i_104761818(.A(n_300791816), .B(n_2991), .Z(n_58002));
	notech_ao4 i_104861817(.A(n_61110), .B(n_30825), .C(n_300891815), .D(n_299691827
		), .Z(n_58001));
	notech_nand3 i_12288(.A(n_60144), .B(n_60234), .C(read_data[12]), .Z(n_47649
		));
	notech_nand2 i_1520772(.A(n_140368420), .B(n_139568412), .Z(n_24514));
	notech_nand2 i_1520868(.A(n_141368430), .B(n_140868425), .Z(n_24166));
	notech_nand2 i_1520996(.A(n_142268439), .B(n_141868435), .Z(n_23818));
	notech_nand2 i_1521092(.A(n_143268449), .B(n_142768444), .Z(n_18913));
	notech_nand2 i_1521188(.A(n_144168458), .B(n_143768454), .Z(n_18564));
	notech_nand3 i_3121396(.A(n_144768464), .B(n_144668463), .C(n_144568462)
		, .Z(n_25426));
	notech_and4 i_1521380(.A(n_145468471), .B(n_145668473), .C(n_145368470),
		 .D(n_130868325), .Z(n_25330));
	notech_and4 i_1421379(.A(n_146368480), .B(n_146568482), .C(n_146268479),
		 .D(n_129768314), .Z(n_25324));
	notech_and4 i_1421539(.A(n_147468491), .B(n_147368490), .C(n_147268489),
		 .D(n_147768494), .Z(n_18210));
	notech_nand2 i_1321538(.A(n_148968506), .B(n_148468501), .Z(n_18204));
	notech_nand2 i_521530(.A(n_150268519), .B(n_149668513), .Z(n_18156));
	notech_nand2 i_221527(.A(n_151568532), .B(n_150968526), .Z(n_18138));
	notech_nand2 i_1521636(.A(n_152468541), .B(n_152068537), .Z(n_17864));
	notech_and4 i_1521860(.A(n_153068547), .B(n_152968546), .C(n_122168238),
		 .D(n_153368550), .Z(n_20702));
	notech_and4 i_1521924(.A(n_154168558), .B(n_154068557), .C(n_121068227),
		 .D(n_154468561), .Z(n_17516));
	notech_and4 i_1421923(.A(n_155268569), .B(n_155168568), .C(n_119968216),
		 .D(n_155568572), .Z(n_17510));
	notech_and4 i_1517604(.A(n_156068577), .B(n_156668583), .C(n_119268209),
		 .D(n_155968576), .Z(n_16790));
	notech_ao4 i_95141375(.A(n_59445), .B(n_27179), .C(n_2414), .D(n_26707),
		 .Z(n_58098));
	notech_nand2 i_95241376(.A(n_311191712), .B(n_316291661), .Z(n_58097));
	notech_and3 i_60941374(.A(n_315691667), .B(n_311291711), .C(n_322070231)
		, .Z(n_58408));
	notech_or2 i_35847350(.A(n_3864), .B(n_147228749), .Z(n_238565914));
	notech_and2 i_191041337(.A(n_57084), .B(n_57731), .Z(n_57181));
	notech_and2 i_64341336(.A(n_58425), .B(n_314670157), .Z(n_58374));
	notech_and2 i_124041330(.A(n_57867), .B(n_26600), .Z(n_57809));
	notech_and3 i_124241332(.A(n_57865), .B(n_57470), .C(n_45139), .Z(n_57807
		));
	notech_and2 i_64141329(.A(n_58423), .B(n_314570156), .Z(n_58376));
	notech_or2 i_36547343(.A(n_310191722), .B(n_27459), .Z(n_237865907));
	notech_and2 i_63458550(.A(n_27319), .B(n_304391780), .Z(n_58383));
	notech_and2 i_64758548(.A(n_4014), .B(n_159168608), .Z(n_58370));
	notech_nand2 i_94758535(.A(n_23513), .B(n_316491659), .Z(n_58102));
	notech_ao4 i_97858532(.A(n_27746), .B(n_305191772), .C(n_58432), .D(eval_flag
		), .Z(n_58071));
	notech_ao4 i_122858526(.A(n_306291761), .B(n_26610), .C(n_306891755), .D
		(n_305191772), .Z(n_57821));
	notech_and2 i_133858521(.A(n_185268869), .B(n_27259), .Z(n_57711));
	notech_nao3 i_32465(.A(n_60144), .B(n_60329), .C(n_32378), .Z(n_280634762
		));
	notech_and4 i_1320770(.A(n_185768874), .B(n_185968876), .C(n_186968885),
		 .D(n_183168848), .Z(n_24502));
	notech_nand2 i_1320866(.A(n_188868903), .B(n_188468899), .Z(n_24154));
	notech_and4 i_1320994(.A(n_188968904), .B(n_189268906), .C(n_189768911),
		 .D(n_180268819), .Z(n_23806));
	notech_nand2 i_1321090(.A(n_190768920), .B(n_190268916), .Z(n_18901));
	notech_and4 i_1321186(.A(n_190868921), .B(n_191068923), .C(n_191568928),
		 .D(n_178368800), .Z(n_18552));
	notech_and4 i_1321378(.A(n_192168934), .B(n_192368936), .C(n_176968786),
		 .D(n_192068933), .Z(n_25318));
	notech_and4 i_1121376(.A(n_193068943), .B(n_193268945), .C(n_192968942),
		 .D(n_175868775), .Z(n_25306));
	notech_nand2 i_821373(.A(n_194668959), .B(n_194168954), .Z(n_25288));
	notech_nand2 i_521370(.A(n_195768970), .B(n_195268965), .Z(n_25270));
	notech_nand2 i_221367(.A(n_196968982), .B(n_196368976), .Z(n_25252));
	notech_and4 i_121366(.A(n_197668989), .B(n_198468996), .C(n_170868725), 
		.D(n_197568988), .Z(n_25246));
	notech_nand2 i_1121536(.A(n_199569007), .B(n_199069002), .Z(n_18192));
	notech_and4 i_121526(.A(n_200469016), .B(n_200769019), .C(n_200369015), 
		.D(n_167568692), .Z(n_18132));
	notech_and4 i_1321634(.A(n_200969021), .B(n_201169023), .C(n_201669028),
		 .D(n_167168688), .Z(n_17852));
	notech_and4 i_1321858(.A(n_201769029), .B(n_201969031), .C(n_202469036),
		 .D(n_166268679), .Z(n_20690));
	notech_or4 i_1621925(.A(n_164668663), .B(n_203469046), .C(n_26585), .D(n_26586
		), .Z(n_17522));
	notech_or4 i_1321922(.A(n_163468651), .B(n_186768883), .C(n_204269054), 
		.D(n_26582), .Z(n_17504));
	notech_and4 i_1221921(.A(n_205169063), .B(n_205069062), .C(n_162668643),
		 .D(n_205469066), .Z(n_17498));
	notech_and4 i_1121920(.A(n_161668633), .B(n_206169073), .C(n_206069072),
		 .D(n_206469076), .Z(n_17492));
	notech_or4 i_1021919(.A(n_160568622), .B(n_207769089), .C(n_26576), .D(n_26577
		), .Z(n_17486));
	notech_nand2 i_1317602(.A(n_208869100), .B(n_208369095), .Z(n_16778));
	notech_ao4 i_2758462(.A(n_27754), .B(n_27306), .C(n_27746), .D(n_56508),
		 .Z(n_57812));
	notech_and4 i_260758501(.A(n_56848), .B(n_55735), .C(n_304991774), .D(n_1441
		), .Z(n_56508));
	notech_or2 i_10558386(.A(n_32356), .B(n_303391790), .Z(n_269834654));
	notech_or2 i_34447364(.A(n_60008), .B(n_147228749), .Z(n_237165900));
	notech_or2 i_35147357(.A(n_310191722), .B(n_27457), .Z(n_236465893));
	notech_or4 i_33747371(.A(n_26613), .B(n_57087), .C(n_57068), .D(n_26770)
		, .Z(n_236165890));
	notech_nand2 i_167041296(.A(n_27179), .B(n_26941), .Z(n_57415));
	notech_or4 i_129847745(.A(n_26614), .B(n_57087), .C(n_57068), .D(n_26770
		), .Z(n_236065889));
	notech_or2 i_32947379(.A(n_60009), .B(n_147228749), .Z(n_235565884));
	notech_nand3 i_58555617(.A(n_60329), .B(n_1901), .C(n_32386), .Z(n_58432
		));
	notech_nao3 i_131855580(.A(n_209069102), .B(n_32331), .C(n_58099), .Z(n_57731
		));
	notech_or4 i_200855553(.A(n_32342), .B(n_32339), .C(n_58099), .D(n_58486
		), .Z(n_57084));
	notech_nor2 i_11774(.A(n_304891775), .B(n_306391760), .Z(n_48163));
	notech_and4 i_1021375(.A(n_211869130), .B(n_212069132), .C(n_211769129),
		 .D(n_210469116), .Z(n_25300));
	notech_or4 i_3121652(.A(n_117868195), .B(n_209269104), .C(n_212569137), 
		.D(n_26574), .Z(n_17960));
	notech_ao4 i_94355545(.A(n_58186), .B(n_27992), .C(n_59968), .D(n_32348)
		, .Z(n_58106));
	notech_or2 i_181353970(.A(n_1874), .B(n_3912), .Z(n_346670477));
	notech_or4 i_19598(.A(n_32643), .B(n_2875), .C(n_2839), .D(n_1864), .Z(n_346770478
		));
	notech_mux2 i_2611695(.S(n_60548), .A(regs_14[25]), .B(add_len_pc32[25])
		, .Z(add_len_pc[25]));
	notech_and4 i_144850673(.A(n_254769559), .B(n_254669558), .C(n_254269554
		), .D(n_254569557), .Z(n_288927271));
	notech_nand2 i_2620719(.A(n_255969571), .B(n_255469566), .Z(n_24906));
	notech_and4 i_2620783(.A(n_256169573), .B(n_256369575), .C(n_250269514),
		 .D(n_257269584), .Z(n_24580));
	notech_or4 i_2620879(.A(n_257069582), .B(n_247469486), .C(n_258869600), 
		.D(n_26578), .Z(n_24232));
	notech_or4 i_2621007(.A(n_257069582), .B(n_246669478), .C(n_259569607), 
		.D(n_26579), .Z(n_23884));
	notech_and4 i_2621103(.A(n_259969611), .B(n_260169613), .C(n_246569477),
		 .D(n_260669618), .Z(n_18979));
	notech_or4 i_2621199(.A(n_257069582), .B(n_244969461), .C(n_261069622), 
		.D(n_26581), .Z(n_18630));
	notech_nand3 i_2621391(.A(n_261969631), .B(n_261869630), .C(n_261769629)
		, .Z(n_25396));
	notech_nand3 i_2521390(.A(n_262669638), .B(n_262569637), .C(n_262469636)
		, .Z(n_25390));
	notech_nand3 i_2421389(.A(n_263369645), .B(n_263269644), .C(n_263169643)
		, .Z(n_25384));
	notech_nand3 i_2321388(.A(n_264069652), .B(n_263969651), .C(n_263869650)
		, .Z(n_25378));
	notech_nand2 i_2621551(.A(n_265169663), .B(n_264669658), .Z(n_18282));
	notech_and4 i_321528(.A(n_266069672), .B(n_265969671), .C(n_265869670), 
		.D(n_266369675), .Z(n_18144));
	notech_or4 i_2621647(.A(n_257069582), .B(n_237869390), .C(n_266869680), 
		.D(n_26583), .Z(n_17930));
	notech_or4 i_2621871(.A(n_257069582), .B(n_237069382), .C(n_267569687), 
		.D(n_26584), .Z(n_20768));
	notech_and4 i_2521870(.A(n_267969691), .B(n_268169693), .C(n_268669698),
		 .D(n_236969381), .Z(n_20762));
	notech_and4 i_2621935(.A(n_269169703), .B(n_269369705), .C(n_235669368),
		 .D(n_269069702), .Z(n_17582));
	notech_and4 i_321912(.A(n_270269714), .B(n_270169713), .C(n_234269354), 
		.D(n_270569717), .Z(n_17444));
	notech_and4 i_2617039(.A(n_271269724), .B(n_271469726), .C(n_271169723),
		 .D(n_233169343), .Z(n_17225));
	notech_or4 i_2617615(.A(n_231769329), .B(n_257069582), .C(n_272269734), 
		.D(n_26587), .Z(n_16856));
	notech_or4 i_2417613(.A(n_230769319), .B(n_258069592), .C(n_273169743), 
		.D(n_26588), .Z(n_16844));
	notech_or4 i_2317612(.A(n_258469596), .B(n_229769309), .C(n_274069752), 
		.D(n_26589), .Z(n_16838));
	notech_or2 i_33647372(.A(n_310191722), .B(n_27455), .Z(n_234865877));
	notech_or2 i_31647392(.A(n_3837), .B(n_59980), .Z(n_234565874));
	notech_or2 i_31947389(.A(n_148228759), .B(n_60004), .Z(n_234265871));
	notech_nao3 i_32247386(.A(opc_10[21]), .B(n_62782), .C(n_3843), .Z(n_233965868
		));
	notech_ao4 i_111447730(.A(n_304891775), .B(n_56939), .C(n_304991774), .D
		(n_306891755), .Z(n_57935));
	notech_ao4 i_193447727(.A(n_30821), .B(n_61110), .C(n_301091813), .D(n_300491819
		), .Z(n_233165860));
	notech_or4 i_1820871(.A(n_288769899), .B(n_284469856), .C(n_289269904), 
		.D(n_26590), .Z(n_24184));
	notech_and4 i_2121098(.A(n_289669908), .B(n_289869910), .C(n_290369915),
		 .D(n_284369855), .Z(n_18949));
	notech_nand2 i_2021097(.A(n_291269924), .B(n_290869920), .Z(n_18943));
	notech_and4 i_1921192(.A(n_291369925), .B(n_291569927), .C(n_292069932),
		 .D(n_282469836), .Z(n_18588));
	notech_nand3 i_2121386(.A(n_292669938), .B(n_292569937), .C(n_292469936)
		, .Z(n_25366));
	notech_and4 i_2021385(.A(n_293269944), .B(n_293469946), .C(n_280169813),
		 .D(n_293169943), .Z(n_25360));
	notech_and4 i_1921384(.A(n_294069952), .B(n_294269954), .C(n_279169803),
		 .D(n_293969951), .Z(n_25354));
	notech_and4 i_1821383(.A(n_294469956), .B(n_294669958), .C(n_278669798),
		 .D(n_295169963), .Z(n_25348));
	notech_nand3 i_1721382(.A(n_295869970), .B(n_295769969), .C(n_295669968)
		, .Z(n_25342));
	notech_nand2 i_1721542(.A(n_297269984), .B(n_296669978), .Z(n_18228));
	notech_nand3 i_57747141(.A(n_313991684), .B(n_60144), .C(n_60331), .Z(n_233065859
		));
	notech_or4 i_57647142(.A(n_61138), .B(n_60234), .C(n_26602), .D(n_32380)
		, .Z(n_232965858));
	notech_and2 i_69844525(.A(n_58432), .B(n_298970000), .Z(n_58319));
	notech_and2 i_8147618(.A(n_312324377), .B(n_259166120), .Z(n_232865857)
		);
	notech_nand2 i_8047619(.A(n_26700), .B(n_233065859), .Z(n_232765856));
	notech_and3 i_7947620(.A(n_301891805), .B(n_300391820), .C(n_232965858),
		 .Z(n_232665855));
	notech_ao4 i_193247739(.A(n_30821), .B(n_61110), .C(n_312191702), .D(n_319291631
		), .Z(n_232565854));
	notech_and3 i_8547614(.A(n_236065889), .B(n_344666975), .C(n_236165890),
		 .Z(n_232465853));
	notech_and4 i_130449395(.A(n_232165850), .B(n_231965848), .C(n_208865617
		), .D(n_209165620), .Z(n_232365852));
	notech_ao4 i_130049399(.A(n_146328740), .B(n_28618), .C(n_146228739), .D
		(n_29827), .Z(n_232165850));
	notech_and2 i_115844562(.A(n_58514), .B(n_299070001), .Z(n_57891));
	notech_and4 i_116744556(.A(n_312391700), .B(n_312770138), .C(n_58530), .D
		(n_151028787), .Z(n_57882));
	notech_and2 i_60744555(.A(n_310691717), .B(n_311691707), .Z(n_58410));
	notech_and2 i_50344519(.A(n_309491729), .B(n_299170002), .Z(n_58514));
	notech_ao4 i_130249397(.A(n_60000), .B(n_147228749), .C(n_147128748), .D
		(n_29770), .Z(n_231965848));
	notech_and4 i_131049389(.A(n_231665845), .B(n_231465843), .C(n_231365842
		), .D(n_209465623), .Z(n_231865847));
	notech_ao4 i_130549394(.A(n_310391720), .B(n_28010), .C(n_60148), .D(n_27183
		), .Z(n_231665845));
	notech_and4 i_3221397(.A(n_308970100), .B(n_308870099), .C(n_308670097),
		 .D(n_308570096), .Z(n_25432));
	notech_nand2 i_721532(.A(n_310070111), .B(n_309670107), .Z(n_18168));
	notech_nand2 i_621531(.A(n_311370124), .B(n_310770118), .Z(n_18162));
	notech_nand2 i_421529(.A(n_312670137), .B(n_312070131), .Z(n_18150));
	notech_and4 i_142644501(.A(n_308170092), .B(n_308070091), .C(n_307670087
		), .D(n_307970090), .Z(n_308721251));
	notech_ao4 i_130749392(.A(n_146928746), .B(n_57771), .C(n_288927271), .D
		(n_146428741), .Z(n_231465843));
	notech_ao4 i_130849391(.A(n_256069572), .B(n_301791806), .C(n_253569547)
		, .D(n_310491719), .Z(n_231365842));
	notech_and3 i_143249268(.A(n_230865837), .B(n_208365612), .C(n_231065839
		), .Z(n_231165840));
	notech_ao4 i_143149269(.A(n_28527), .B(n_29830), .C(n_28530), .D(n_29828
		), .Z(n_231065839));
	notech_ao4 i_114250652(.A(n_2992), .B(n_29733), .C(n_60023), .D(n_2991),
		 .Z(n_230865837));
	notech_ao4 i_143349267(.A(n_28236), .B(n_344366972), .C(n_268366212), .D
		(n_57557), .Z(n_230665835));
	notech_nand3 i_20583(.A(n_56848), .B(n_311991704), .C(n_2004), .Z(n_39370
		));
	notech_nand2 i_124141331(.A(n_57298), .B(n_57901), .Z(n_57808));
	notech_and4 i_143541317(.A(n_323870249), .B(n_323770248), .C(n_323370244
		), .D(n_323670247), .Z(n_59965));
	notech_mux2 i_1311682(.S(n_60548), .A(n_5172), .B(add_len_pc32[12]), .Z(add_len_pc
		[12]));
	notech_or4 i_9029(.A(n_32343), .B(n_32342), .C(n_314891675), .D(n_24994)
		, .Z(n_50904));
	notech_ao4 i_143449266(.A(n_268266211), .B(\nbus_11358[2] ), .C(n_303291791
		), .D(n_27984), .Z(n_230565834));
	notech_nand2 i_1320706(.A(n_325170262), .B(n_324670257), .Z(n_24828));
	notech_and4 i_921374(.A(n_325870269), .B(n_326070271), .C(n_325770268), 
		.D(n_317670187), .Z(n_25294));
	notech_nand2 i_921534(.A(n_327270283), .B(n_326770278), .Z(n_18180));
	notech_nand2 i_921918(.A(n_328170292), .B(n_327770288), .Z(n_17480));
	notech_and4 i_144249258(.A(n_230265831), .B(n_230065829), .C(n_229965828
		), .D(n_210765636), .Z(n_230465833));
	notech_ao4 i_143749263(.A(n_59991), .B(n_28502), .C(n_58316), .D(n_303891785
		), .Z(n_230265831));
	notech_and4 i_91438297(.A(n_337170382), .B(n_337070381), .C(n_336670377)
		, .D(n_336970380), .Z(n_60022));
	notech_and4 i_92338288(.A(n_338570396), .B(n_338470395), .C(n_338070391)
		, .D(n_338370394), .Z(n_60013));
	notech_and4 i_93638275(.A(n_339970410), .B(n_339870409), .C(n_339470405)
		, .D(n_339770408), .Z(n_60000));
	notech_nand2 i_2616239(.A(n_341270423), .B(n_340770418), .Z(n_19256));
	notech_and4 i_1316226(.A(n_341870429), .B(n_341770428), .C(n_342970440),
		 .D(n_341670427), .Z(n_19178));
	notech_or2 i_177438222(.A(n_54912649), .B(n_328270293), .Z(n_309115167)
		);
	notech_nand3 i_56143(.A(n_114368160), .B(n_343370444), .C(n_114568162), 
		.Z(\nbus_11376[8] ));
	notech_ao4 i_122635132(.A(calc_sz[1]), .B(n_246691943), .C(n_26782), .D(n_56941
		), .Z(n_57823));
	notech_or4 i_177735123(.A(n_2873), .B(n_2872), .C(n_27754), .D(n_26789),
		 .Z(n_57314));
	notech_and3 i_127735122(.A(n_26962), .B(n_56983), .C(n_27896), .Z(n_57772
		));
	notech_nao3 i_228871053(.A(calc_sz[0]), .B(calc_sz[1]), .C(n_2937), .Z(n_56809
		));
	notech_nand3 i_57335120(.A(n_27377), .B(n_60331), .C(n_2988), .Z(n_58444
		));
	notech_or4 i_98235094(.A(n_60938), .B(n_60909), .C(n_61138), .D(n_60234)
		, .Z(n_308012096));
	notech_ao4 i_143949261(.A(n_152472004), .B(n_28234), .C(n_152572005), .D
		(n_111664645), .Z(n_230065829));
	notech_or4 i_10935001(.A(n_32643), .B(n_2875), .C(n_2839), .D(n_60868), 
		.Z(n_2985));
	notech_ao4 i_144049260(.A(n_28544), .B(n_208065609), .C(n_207965608), .D
		(n_199965528), .Z(n_229965828));
	notech_nao3 i_29221(.A(n_345470465), .B(n_345670467), .C(n_345370464), .Z
		(n_1978));
	notech_or4 i_2817617(.A(n_344070451), .B(n_1978), .C(n_346370474), .D(n_26603
		), .Z(n_16868));
	notech_mux2 i_144349257(.S(n_32612), .A(n_312147737), .B(n_344466973), .Z
		(n_229865827));
	notech_and4 i_145249252(.A(n_229565824), .B(n_229365822), .C(n_211665645
		), .D(n_211965648), .Z(n_229765826));
	notech_ao4 i_144449256(.A(n_28530), .B(n_29831), .C(n_140128678), .D(\nbus_11365[22] 
		), .Z(n_229565824));
	notech_ao4 i_145049254(.A(n_140428681), .B(n_60003), .C(n_29708), .D(n_140328680
		), .Z(n_229365822));
	notech_and4 i_145749247(.A(n_229065819), .B(n_228865817), .C(n_212265651
		), .D(n_212565654), .Z(n_229265821));
	notech_ao4 i_145349251(.A(n_303591788), .B(n_28007), .C(n_60149), .D(n_27239
		), .Z(n_229065819));
	notech_ao4 i_145549249(.A(n_225765786), .B(n_309691727), .C(n_224065769)
		, .D(n_26678), .Z(n_228865817));
	notech_and4 i_146249242(.A(n_228565814), .B(n_228365812), .C(n_212865657
		), .D(n_213165660), .Z(n_228765816));
	notech_ao4 i_145849246(.A(n_28530), .B(n_29832), .C(n_140128678), .D(\nbus_11365[23] 
		), .Z(n_228565814));
	notech_ao4 i_146049244(.A(n_140428681), .B(n_60002), .C(n_140328680), .D
		(n_29765), .Z(n_228365812));
	notech_and4 i_146749237(.A(n_228065809), .B(n_227865807), .C(n_213465663
		), .D(n_213765666), .Z(n_228265811));
	notech_ao4 i_146349241(.A(n_303591788), .B(n_28008), .C(n_60148), .D(n_27240
		), .Z(n_228065809));
	notech_ao4 i_146549239(.A(n_225665785), .B(n_309691727), .C(n_222565754)
		, .D(n_26678), .Z(n_227865807));
	notech_and4 i_147249232(.A(n_227565804), .B(n_227365802), .C(n_214065669
		), .D(n_214365672), .Z(n_227765806));
	notech_ao4 i_146849236(.A(n_28530), .B(n_29833), .C(n_140128678), .D(\nbus_11365[24] 
		), .Z(n_227565804));
	notech_ao4 i_147049234(.A(n_140428681), .B(n_60001), .C(n_140328680), .D
		(n_29769), .Z(n_227365802));
	notech_and4 i_147749227(.A(n_227065799), .B(n_226865797), .C(n_214665675
		), .D(n_214965678), .Z(n_227265801));
	notech_ao4 i_147349231(.A(n_303591788), .B(n_28009), .C(n_60148), .D(n_27241
		), .Z(n_227065799));
	notech_ao4 i_147549229(.A(n_225565784), .B(n_309691727), .C(n_221065739)
		, .D(n_26678), .Z(n_226865797));
	notech_and4 i_148249222(.A(n_226565794), .B(n_226365792), .C(n_215265681
		), .D(n_215565684), .Z(n_226765796));
	notech_ao4 i_147849226(.A(n_28530), .B(n_29834), .C(n_140128678), .D(n_57771
		), .Z(n_226565794));
	notech_ao4 i_148049224(.A(n_60000), .B(n_140428681), .C(n_140328680), .D
		(n_29770), .Z(n_226365792));
	notech_and4 i_148749217(.A(n_226065789), .B(n_225865787), .C(n_215865687
		), .D(n_216165690), .Z(n_226265791));
	notech_ao4 i_148349221(.A(n_303591788), .B(n_28010), .C(n_60149), .D(n_27242
		), .Z(n_226065789));
	notech_ao4 i_148549219(.A(n_256069572), .B(n_309691727), .C(n_253569547)
		, .D(n_26678), .Z(n_225865787));
	notech_nand2 i_2250671(.A(opc_10[22]), .B(n_62808), .Z(n_225765786));
	notech_nand2 i_2350670(.A(opc_10[23]), .B(n_62822), .Z(n_225665785));
	notech_nand2 i_2450669(.A(opc_10[24]), .B(n_62822), .Z(n_225565784));
	notech_ao4 i_182248886(.A(n_26924), .B(n_28247), .C(n_26922), .D(n_28212
		), .Z(n_225265781));
	notech_ao4 i_182348885(.A(n_56921), .B(n_29835), .C(n_26969), .D(n_28279
		), .Z(n_225165780));
	notech_and2 i_182748881(.A(n_224965778), .B(n_224865777), .Z(n_225065779
		));
	notech_ao4 i_182548883(.A(n_26927), .B(n_28312), .C(n_26649), .D(n_29837
		), .Z(n_224965778));
	notech_ao4 i_182648882(.A(n_26920), .B(n_28377), .C(n_26933), .D(n_28345
		), .Z(n_224865777));
	notech_and4 i_183548873(.A(n_224565774), .B(n_224465773), .C(n_224265771
		), .D(n_224165770), .Z(n_224765776));
	notech_ao4 i_182948879(.A(n_56630), .B(n_28441), .C(n_56619), .D(n_28409
		), .Z(n_224565774));
	notech_ao4 i_183048878(.A(n_26928), .B(n_28473), .C(n_26651), .D(n_28180
		), .Z(n_224465773));
	notech_ao4 i_183248876(.A(n_26925), .B(n_28506), .C(n_27036), .D(n_28548
		), .Z(n_224265771));
	notech_ao4 i_183348875(.A(n_56557), .B(n_27883), .C(n_56548), .D(n_28583
		), .Z(n_224165770));
	notech_nand2 i_40250667(.A(opc[22]), .B(n_62822), .Z(n_224065769));
	notech_ao4 i_184748862(.A(n_26924), .B(n_28248), .C(n_26922), .D(n_28213
		), .Z(n_223765766));
	notech_ao4 i_184848861(.A(n_56921), .B(n_29838), .C(n_26969), .D(n_28280
		), .Z(n_223665765));
	notech_and2 i_185248857(.A(n_223465763), .B(n_223365762), .Z(n_223565764
		));
	notech_ao4 i_185048859(.A(n_26927), .B(n_28313), .C(n_26649), .D(n_29839
		), .Z(n_223465763));
	notech_ao4 i_185148858(.A(n_26920), .B(n_28378), .C(n_26933), .D(n_28346
		), .Z(n_223365762));
	notech_and4 i_186048849(.A(n_223065759), .B(n_222965758), .C(n_222765756
		), .D(n_222665755), .Z(n_223265761));
	notech_ao4 i_185448855(.A(n_56630), .B(n_28442), .C(n_56619), .D(n_28410
		), .Z(n_223065759));
	notech_ao4 i_185548854(.A(n_26928), .B(n_28474), .C(n_26651), .D(n_28181
		), .Z(n_222965758));
	notech_ao4 i_185748852(.A(n_26925), .B(n_28507), .C(n_27036), .D(n_28549
		), .Z(n_222765756));
	notech_ao4 i_185848851(.A(n_26721), .B(n_27884), .C(n_56548), .D(n_28584
		), .Z(n_222665755));
	notech_nand2 i_40350666(.A(opc[23]), .B(n_62794), .Z(n_222565754));
	notech_ao4 i_187148838(.A(n_26924), .B(n_28249), .C(n_26922), .D(n_28214
		), .Z(n_222265751));
	notech_ao4 i_187248837(.A(n_56921), .B(n_29840), .C(n_26969), .D(n_28281
		), .Z(n_222165750));
	notech_and2 i_187648833(.A(n_221965748), .B(n_221865747), .Z(n_222065749
		));
	notech_ao4 i_187448835(.A(n_26927), .B(n_28314), .C(n_26649), .D(n_29841
		), .Z(n_221965748));
	notech_ao4 i_187548834(.A(n_26920), .B(n_28379), .C(n_26933), .D(n_28347
		), .Z(n_221865747));
	notech_and4 i_188948825(.A(n_221565744), .B(n_221465743), .C(n_221265741
		), .D(n_221165740), .Z(n_221765746));
	notech_ao4 i_188248831(.A(n_56630), .B(n_28443), .C(n_56619), .D(n_28411
		), .Z(n_221565744));
	notech_ao4 i_188348830(.A(n_26928), .B(n_28475), .C(n_26651), .D(n_28182
		), .Z(n_221465743));
	notech_ao4 i_188648828(.A(n_26925), .B(n_28508), .C(n_27036), .D(n_28550
		), .Z(n_221265741));
	notech_ao4 i_188748827(.A(n_26721), .B(n_27886), .C(n_56548), .D(n_28585
		), .Z(n_221165740));
	notech_nand2 i_40550665(.A(opc[24]), .B(n_62804), .Z(n_221065739));
	notech_or2 i_56750111(.A(n_288927271), .B(n_139728674), .Z(n_216165690)
		);
	notech_nand3 i_57050108(.A(n_60149), .B(n_60234), .C(read_data[25]), .Z(n_215865687
		));
	notech_or2 i_57350105(.A(n_140228679), .B(n_55965), .Z(n_215565684));
	notech_nand3 i_57650102(.A(n_1430), .B(n_6399), .C(n_29601), .Z(n_215265681
		));
	notech_or2 i_55450123(.A(n_139728674), .B(n_289027272), .Z(n_214965678)
		);
	notech_nand3 i_55750120(.A(n_60149), .B(n_60241), .C(read_data[24]), .Z(n_214665675
		));
	notech_or2 i_56150117(.A(n_140228679), .B(\nbus_11358[24] ), .Z(n_214365672
		));
	notech_nand3 i_56450114(.A(n_1430), .B(n_6397), .C(n_29601), .Z(n_214065669
		));
	notech_or2 i_54150135(.A(n_139728674), .B(n_289127273), .Z(n_213765666)
		);
	notech_nand3 i_54450132(.A(n_60149), .B(n_60241), .C(read_data[23]), .Z(n_213465663
		));
	notech_or2 i_54750129(.A(n_140228679), .B(\nbus_11358[23] ), .Z(n_213165660
		));
	notech_nand3 i_55150126(.A(n_1430), .B(n_6395), .C(n_56163), .Z(n_212865657
		));
	notech_or2 i_52750147(.A(n_139728674), .B(n_289227274), .Z(n_212565654)
		);
	notech_nand3 i_53150144(.A(n_60148), .B(n_60241), .C(read_data[22]), .Z(n_212265651
		));
	notech_or2 i_53450141(.A(n_140228679), .B(\nbus_11358[22] ), .Z(n_211965648
		));
	notech_nand3 i_53750138(.A(n_1430), .B(n_6393), .C(n_56163), .Z(n_211665645
		));
	notech_nand2 i_50950163(.A(sav_edi[2]), .B(n_61138), .Z(n_210765636));
	notech_or4 i_34550323(.A(n_32555), .B(n_61138), .C(n_60331), .D(n_28114)
		, .Z(n_209465623));
	notech_or2 i_34850320(.A(n_147028747), .B(n_55965), .Z(n_209165620));
	notech_or2 i_35150317(.A(n_310191722), .B(n_27475), .Z(n_208865617));
	notech_nand3 i_52150152(.A(n_60148), .B(n_60234), .C(read_data[2]), .Z(n_208365612
		));
	notech_and2 i_4350623(.A(n_229865827), .B(n_58714), .Z(n_208065609));
	notech_mux2 i_4250624(.S(n_32612), .A(n_285027232), .B(n_284927231), .Z(n_207965608
		));
	notech_or4 i_45955066(.A(n_61175), .B(n_61165), .C(n_61154), .D(n_206965598
		), .Z(n_207465603));
	notech_or2 i_45855067(.A(n_58318), .B(eval_flag), .Z(n_207365602));
	notech_or2 i_29384(.A(n_32382), .B(n_26602), .Z(n_207265601));
	notech_ao4 i_7255445(.A(n_26702), .B(n_56983), .C(n_26962), .D(n_307791746
		), .Z(n_206965598));
	notech_ao4 i_135957182(.A(n_310191722), .B(n_27422), .C(n_146328740), .D
		(n_28593), .Z(n_206665595));
	notech_ao4 i_136057181(.A(n_310291721), .B(n_28089), .C(n_312991694), .D
		(\nbus_11358[0] ), .Z(n_206465593));
	notech_ao3 i_136657175(.A(n_206065589), .B(n_206265591), .C(n_26704), .Z
		(n_206365592));
	notech_ao4 i_136357178(.A(n_60148), .B(n_27153), .C(n_61110), .D(n_58689
		), .Z(n_206265591));
	notech_ao4 i_136457177(.A(n_191465443), .B(n_205265581), .C(n_191365442)
		, .D(n_205765586), .Z(n_206065589));
	notech_ao4 i_137057171(.A(\nbus_11358[0] ), .B(n_191765446), .C(n_26789)
		, .D(n_191665445), .Z(n_205965588));
	notech_or4 i_137157170(.A(n_32378), .B(n_61115), .C(n_32730), .D(n_56619
		), .Z(n_205765586));
	notech_ao4 i_136757174(.A(n_59434), .B(n_29742), .C(n_291163178), .D(n_54930
		), .Z(n_205665585));
	notech_ao4 i_136857173(.A(n_60025), .B(n_26611), .C(n_29742), .D(n_317191652
		), .Z(n_205465583));
	notech_or4 i_6758424(.A(n_32378), .B(n_205165580), .C(n_61142), .D(n_60234
		), .Z(n_205265581));
	notech_ao3 i_4458447(.A(n_246991940), .B(n_62892), .C(n_246891941), .Z(n_205165580
		));
	notech_and4 i_137757164(.A(n_204865577), .B(n_204665575), .C(n_204565574
		), .D(n_194765476), .Z(n_205065579));
	notech_ao4 i_137257169(.A(n_146328740), .B(n_28603), .C(n_146228739), .D
		(n_29820), .Z(n_204865577));
	notech_ao4 i_137457167(.A(n_3851), .B(n_313191692), .C(n_31433), .D(n_344666975
		), .Z(n_204665575));
	notech_ao4 i_137557166(.A(n_344866977), .B(n_27993), .C(n_31411), .D(n_26616
		), .Z(n_204565574));
	notech_and4 i_138357158(.A(n_204265571), .B(n_204065569), .C(n_203965568
		), .D(n_195465483), .Z(n_204465573));
	notech_ao4 i_137857163(.A(n_344966978), .B(\nbus_11307[10] ), .C(n_292266451
		), .D(n_29684), .Z(n_204265571));
	notech_ao4 i_138057161(.A(n_3850), .B(n_292366452), .C(n_310291721), .D(n_28099
		), .Z(n_204065569));
	notech_ao4 i_138157160(.A(n_60148), .B(n_27166), .C(n_346866997), .D(n_87532846
		), .Z(n_203965568));
	notech_and4 i_155956986(.A(n_185362136), .B(n_185262135), .C(n_158668603
		), .D(n_195965488), .Z(n_203765566));
	notech_ao4 i_156056985(.A(n_59993), .B(n_28502), .C(n_291163178), .D(n_28236
		), .Z(n_203465563));
	notech_and4 i_156856977(.A(n_203165560), .B(n_202965558), .C(n_202765556
		), .D(n_196565494), .Z(n_203365562));
	notech_ao4 i_156356982(.A(n_291363180), .B(n_199965528), .C(n_28527), .D
		(n_29821), .Z(n_203165560));
	notech_ao4 i_156556980(.A(n_28530), .B(n_29822), .C(n_303891785), .D(n_192565454
		), .Z(n_202965558));
	notech_ao4 i_156956976(.A(n_300591818), .B(\nbus_11307[0] ), .C(\nbus_11358[0] 
		), .D(n_26681), .Z(n_202865557));
	notech_ao4 i_156656979(.A(n_28544), .B(n_192465453), .C(n_175062033), .D
		(n_26705), .Z(n_202765556));
	notech_ao4 i_157056975(.A(n_29742), .B(n_300591818), .C(n_60025), .D(n_26681
		), .Z(n_202665555));
	notech_and4 i_164856899(.A(n_202365552), .B(n_202165550), .C(n_197665505
		), .D(n_197965508), .Z(n_202565554));
	notech_ao4 i_164456903(.A(n_31433), .B(n_297566504), .C(n_292466453), .D
		(n_27993), .Z(n_202365552));
	notech_ao4 i_164656901(.A(n_292566454), .B(\nbus_11307[10] ), .C(n_292866457
		), .D(n_29684), .Z(n_202165550));
	notech_and4 i_165556893(.A(n_201865547), .B(n_201665545), .C(n_201565544
		), .D(n_198265511), .Z(n_202065549));
	notech_ao4 i_164956898(.A(n_32270), .B(n_28099), .C(n_60148), .D(n_27226
		), .Z(n_201865547));
	notech_ao4 i_165156896(.A(n_31411), .B(n_28545), .C(n_87532846), .D(n_292166450
		), .Z(n_201665545));
	notech_ao4 i_165256895(.A(n_28527), .B(n_29824), .C(n_28530), .D(n_29823
		), .Z(n_201565544));
	notech_and4 i_166056888(.A(n_47649), .B(n_201265541), .C(n_201065539), .D
		(n_199165520), .Z(n_201465543));
	notech_ao4 i_165656892(.A(n_59965), .B(n_297466503), .C(n_297566504), .D
		(n_320170212), .Z(n_201265541));
	notech_ao4 i_165856890(.A(\nbus_11358[12] ), .B(n_26667), .C(n_292566454
		), .D(n_57644), .Z(n_201065539));
	notech_and4 i_166656882(.A(n_200765536), .B(n_200565534), .C(n_200465533
		), .D(n_199465523), .Z(n_200965538));
	notech_ao4 i_166156887(.A(n_292766456), .B(n_60013), .C(n_60148), .D(n_27228
		), .Z(n_200765536));
	notech_ao4 i_166356885(.A(n_320070211), .B(n_28545), .C(n_156768584), .D
		(n_292166450), .Z(n_200565534));
	notech_ao4 i_166456884(.A(n_28527), .B(n_29826), .C(n_54649), .D(n_29825
		), .Z(n_200465533));
	notech_ao4 i_29476(.A(\nbus_11307[9] ), .B(n_27305), .C(n_30594), .D(n_29743
		), .Z(n_200265531));
	notech_or4 i_14483(.A(calc_sz[1]), .B(n_246691943), .C(n_26602), .D(n_60016
		), .Z(n_200165530));
	notech_ao4 i_29478(.A(n_192865457), .B(n_192765456), .C(n_58318), .D(\nbus_11358[9] 
		), .Z(n_200065529));
	notech_nand2 i_31761(.A(n_26890), .B(n_26668), .Z(n_199965528));
	notech_or2 i_78157736(.A(n_292866457), .B(n_29679), .Z(n_199465523));
	notech_or2 i_78457733(.A(n_292466453), .B(n_27997), .Z(n_199165520));
	notech_or2 i_76857749(.A(n_3850), .B(n_292766456), .Z(n_198265511));
	notech_nand2 i_77157746(.A(opb[10]), .B(n_292666455), .Z(n_197965508));
	notech_or4 i_77457743(.A(n_32348), .B(n_27036), .C(n_3851), .D(n_61142),
		 .Z(n_197665505));
	notech_nao3 i_71757793(.A(opc[0]), .B(n_62804), .C(n_28234), .Z(n_196565494
		));
	notech_or2 i_72057790(.A(n_303291791), .B(n_27981), .Z(n_196265491));
	notech_nand2 i_72157789(.A(sav_edi[0]), .B(n_61142), .Z(n_195965488));
	notech_or2 i_51457980(.A(n_345066979), .B(\nbus_11358[10] ), .Z(n_195465483
		));
	notech_or2 i_52157973(.A(n_310191722), .B(n_27443), .Z(n_194765476));
	notech_and4 i_50557989(.A(n_60909), .B(n_62806), .C(\opa_12[0] ), .D(n_54930
		), .Z(n_194265471));
	notech_or4 i_48958005(.A(n_280634762), .B(n_191565444), .C(n_205165580),
		 .D(n_56983), .Z(n_193865467));
	notech_nand2 i_49458000(.A(n_7349), .B(n_26986), .Z(n_193365462));
	notech_and2 i_102557502(.A(n_60246), .B(n_28098), .Z(n_192865457));
	notech_and3 i_102457503(.A(n_60331), .B(n_200165530), .C(n_200265531), .Z
		(n_192765456));
	notech_and2 i_15458339(.A(n_58646), .B(n_202865557), .Z(n_192565454));
	notech_and2 i_15358340(.A(n_202665555), .B(n_58610), .Z(n_192465453));
	notech_ao4 i_15258341(.A(n_26770), .B(n_27119), .C(n_28332), .D(n_26683)
		, .Z(n_192365452));
	notech_or4 i_50257992(.A(calc_sz[3]), .B(n_2938), .C(n_26611), .D(calc_sz
		[2]), .Z(n_192165450));
	notech_nand3 i_50157993(.A(opc[0]), .B(n_62806), .C(n_17107), .Z(n_192065449
		));
	notech_or2 i_50057994(.A(n_317191652), .B(\nbus_11307[0] ), .Z(n_191965448
		));
	notech_or4 i_49957995(.A(n_59419), .B(\nbus_11307[0] ), .C(n_26789), .D(n_17107
		), .Z(n_191865447));
	notech_and2 i_12458368(.A(n_3814), .B(n_192165450), .Z(n_191765446));
	notech_and3 i_13158362(.A(n_58646), .B(n_192065449), .C(n_191965448), .Z
		(n_191665445));
	notech_ao3 i_16458329(.A(n_205465583), .B(n_205665585), .C(n_194265471),
		 .Z(n_191565444));
	notech_and2 i_16358330(.A(n_205965588), .B(n_191865447), .Z(n_191465443)
		);
	notech_ao4 i_12058371(.A(n_26789), .B(n_27981), .C(n_59993), .D(n_56983)
		, .Z(n_191365442));
	notech_nand2 i_164058508(.A(n_26890), .B(n_26683), .Z(n_191265441));
	notech_and4 i_127260523(.A(n_190565434), .B(n_190365432), .C(n_26754), .D
		(n_116964698), .Z(n_190765436));
	notech_ao4 i_126860527(.A(n_54643), .B(n_28957), .C(n_151028787), .D(nbus_11295
		[21]), .Z(n_190565434));
	notech_ao4 i_127060525(.A(n_311291711), .B(n_28006), .C(n_151128788), .D
		(n_59980), .Z(n_190365432));
	notech_and4 i_127860518(.A(n_190065429), .B(n_189865427), .C(n_117264701
		), .D(n_117564704), .Z(n_190265431));
	notech_ao4 i_127460522(.A(n_311191712), .B(\nbus_11358[21] ), .C(n_151428791
		), .D(n_60004), .Z(n_190065429));
	notech_ao4 i_127660520(.A(n_311391710), .B(n_110964638), .C(n_316491659)
		, .D(n_111164640), .Z(n_189865427));
	notech_and4 i_145660345(.A(n_125828535), .B(n_189565424), .C(n_189365422
		), .D(n_117964708), .Z(n_189765426));
	notech_ao4 i_145260349(.A(n_60331), .B(n_28110), .C(n_54643), .D(n_28977
		), .Z(n_189565424));
	notech_ao4 i_145460347(.A(n_310691717), .B(n_28006), .C(n_148728764), .D
		(n_59980), .Z(n_189365422));
	notech_and4 i_146160340(.A(n_189065419), .B(n_188865417), .C(n_118264711
		), .D(n_118564714), .Z(n_189265421));
	notech_ao4 i_145760344(.A(n_149428771), .B(\nbus_11358[21] ), .C(n_149128768
		), .D(n_60004), .Z(n_189065419));
	notech_ao4 i_145960342(.A(n_310791716), .B(n_110964638), .C(n_311991704)
		, .D(n_111164640), .Z(n_188865417));
	notech_and4 i_154660261(.A(n_188565414), .B(n_188365412), .C(n_188265411
		), .D(n_118864717), .Z(n_188765416));
	notech_ao4 i_154160266(.A(n_146328740), .B(n_28600), .C(n_146228739), .D
		(n_29794), .Z(n_188565414));
	notech_ao4 i_154360264(.A(n_31279), .B(n_26614), .C(n_310291721), .D(n_28096
		), .Z(n_188365412));
	notech_ao4 i_154460263(.A(n_31309), .B(n_236065889), .C(n_60148), .D(n_27162
		), .Z(n_188265411));
	notech_and4 i_155260255(.A(n_187965408), .B(n_187765406), .C(n_187665405
		), .D(n_119564724), .Z(n_188165410));
	notech_ao4 i_154760260(.A(n_303191792), .B(n_58000), .C(n_57999), .D(n_29614
		), .Z(n_187965408));
	notech_ao4 i_154960258(.A(n_31307), .B(n_111464643), .C(n_303391790), .D
		(n_111564644), .Z(n_187765406));
	notech_ao4 i_155060257(.A(n_111864647), .B(\nbus_11358[7] ), .C(n_111764646
		), .D(\nbus_11307[7] ), .Z(n_187665405));
	notech_and4 i_155960248(.A(n_187165400), .B(n_186965398), .C(n_120264731
		), .D(n_120564734), .Z(n_187365402));
	notech_ao4 i_155560252(.A(n_310191722), .B(n_27441), .C(n_146328740), .D
		(n_28602), .Z(n_187165400));
	notech_ao4 i_155760250(.A(n_291963186), .B(n_344666975), .C(n_310291721)
		, .D(n_28098), .Z(n_186965398));
	notech_and4 i_156760242(.A(n_120864737), .B(n_186665395), .C(n_186465393
		), .D(n_186365392), .Z(n_186865397));
	notech_ao4 i_156060247(.A(n_60148), .B(n_27165), .C(n_56619), .D(n_113864667
		), .Z(n_186665395));
	notech_ao4 i_156260245(.A(n_155165080), .B(n_29743), .C(n_26616), .D(n_112164650
		), .Z(n_186465393));
	notech_ao4 i_156360244(.A(\nbus_11358[9] ), .B(n_112064649), .C(\nbus_11307[9] 
		), .D(n_111964648), .Z(n_186365392));
	notech_and3 i_157160239(.A(n_65435450), .B(n_185965388), .C(n_121364742)
		, .Z(n_186165390));
	notech_ao4 i_156960240(.A(n_146328740), .B(n_28604), .C(n_146228739), .D
		(n_29795), .Z(n_185965388));
	notech_ao4 i_157260238(.A(n_31492), .B(n_346766996), .C(n_30088), .D(n_346866997
		), .Z(n_185765386));
	notech_ao4 i_157360237(.A(n_302891795), .B(n_313191692), .C(n_31476), .D
		(n_344666975), .Z(n_185665385));
	notech_and4 i_158260228(.A(n_185365382), .B(n_185265381), .C(n_185065379
		), .D(n_184965378), .Z(n_185565384));
	notech_ao4 i_157660234(.A(n_345066979), .B(\nbus_11358[11] ), .C(n_344966978
		), .D(\nbus_11307[11] ), .Z(n_185365382));
	notech_ao4 i_157760233(.A(n_344866977), .B(n_27996), .C(n_54874), .D(n_28100
		), .Z(n_185265381));
	notech_ao4 i_157960231(.A(n_29596), .B(n_346666995), .C(n_302491799), .D
		(n_267466203), .Z(n_185065379));
	notech_ao4 i_158060230(.A(n_26616), .B(n_31456), .C(n_60166), .D(n_27167
		), .Z(n_184965378));
	notech_and4 i_158860222(.A(n_184665375), .B(n_184465373), .C(n_184365372
		), .D(n_123064759), .Z(n_184865377));
	notech_ao4 i_158360227(.A(n_54883), .B(n_28605), .C(n_146228739), .D(n_29796
		), .Z(n_184665375));
	notech_ao4 i_158560225(.A(n_320170212), .B(n_344666975), .C(n_59965), .D
		(n_313191692), .Z(n_184465373));
	notech_ao4 i_158660224(.A(n_156768584), .B(n_346866997), .C(n_345066979)
		, .D(n_56221), .Z(n_184365372));
	notech_and4 i_159460216(.A(n_184065369), .B(n_183865367), .C(n_183765366
		), .D(n_123764766), .Z(n_184265371));
	notech_ao4 i_158960221(.A(n_344866977), .B(n_27997), .C(n_54874), .D(n_28101
		), .Z(n_184065369));
	notech_ao4 i_159160219(.A(n_26616), .B(n_320070211), .C(n_60166), .D(n_27168
		), .Z(n_183865367));
	notech_ao4 i_159260218(.A(n_60013), .B(n_292366452), .C(n_292266451), .D
		(n_29679), .Z(n_183765366));
	notech_and3 i_159760213(.A(n_164365172), .B(n_183365362), .C(n_124264771
		), .Z(n_183565364));
	notech_ao4 i_159660214(.A(n_54883), .B(n_28607), .C(n_146228739), .D(n_29797
		), .Z(n_183365362));
	notech_ao4 i_159860212(.A(n_59963), .B(n_313191692), .C(n_298366512), .D
		(n_346766996), .Z(n_183165360));
	notech_ao4 i_159960211(.A(n_298266511), .B(n_344666975), .C(n_344866977)
		, .D(n_27999), .Z(n_183065359));
	notech_and4 i_160860202(.A(n_182765356), .B(n_182665355), .C(n_182465353
		), .D(n_182365352), .Z(n_182965358));
	notech_ao4 i_160260208(.A(n_345066979), .B(\nbus_11358[14] ), .C(n_344966978
		), .D(\nbus_11307[14] ), .Z(n_182765356));
	notech_ao4 i_160360207(.A(n_60011), .B(n_267466203), .C(n_54874), .D(n_28103
		), .Z(n_182665355));
	notech_ao4 i_160560205(.A(n_346666995), .B(n_56257), .C(n_26616), .D(n_298166510
		), .Z(n_182465353));
	notech_ao4 i_160660204(.A(n_60166), .B(n_27169), .C(n_157165100), .D(n_346866997
		), .Z(n_182365352));
	notech_and4 i_161460197(.A(n_162665155), .B(n_182065349), .C(n_181865347
		), .D(n_126164790), .Z(n_182265351));
	notech_ao4 i_160960201(.A(n_310191722), .B(n_27453), .C(n_54883), .D(n_28608
		), .Z(n_182065349));
	notech_ao4 i_161160199(.A(n_298466513), .B(n_344666975), .C(n_54874), .D
		(n_28104), .Z(n_181865347));
	notech_and4 i_162060191(.A(n_181565344), .B(n_181365342), .C(n_181265341
		), .D(n_126464793), .Z(n_181765346));
	notech_ao4 i_161560196(.A(n_111064639), .B(n_346866997), .C(n_56619), .D
		(n_320137996), .Z(n_181565344));
	notech_ao4 i_161760194(.A(n_155165080), .B(n_29754), .C(n_26616), .D(n_112364652
		), .Z(n_181365342));
	notech_ao4 i_161860193(.A(\nbus_11307[15] ), .B(n_111964648), .C(n_112064649
		), .D(\nbus_11358[15] ), .Z(n_181265341));
	notech_and4 i_162660185(.A(n_180965338), .B(n_180765336), .C(n_180665335
		), .D(n_127164800), .Z(n_181165340));
	notech_ao4 i_162160190(.A(n_54883), .B(n_28614), .C(n_54865), .D(n_29798
		), .Z(n_180965338));
	notech_ao4 i_162360188(.A(n_54874), .B(n_28110), .C(n_249866027), .D(n_310491719
		), .Z(n_180765336));
	notech_ao4 i_162460187(.A(n_310391720), .B(n_28006), .C(n_146428741), .D
		(n_59980), .Z(n_180665335));
	notech_and4 i_163260179(.A(n_180365332), .B(n_180165330), .C(n_180065329
		), .D(n_127864807), .Z(n_180565334));
	notech_ao4 i_162760184(.A(n_147028747), .B(\nbus_11358[21] ), .C(n_147228749
		), .D(n_60004), .Z(n_180365332));
	notech_ao4 i_162960182(.A(n_232565854), .B(\nbus_11365[21] ), .C(n_60166
		), .D(n_27176), .Z(n_180165330));
	notech_ao4 i_163060181(.A(n_312191702), .B(n_111164640), .C(n_301791806)
		, .D(n_110964638), .Z(n_180065329));
	notech_and4 i_163760174(.A(n_179765326), .B(n_179565324), .C(n_128564814
		), .D(n_128864817), .Z(n_179965328));
	notech_ao4 i_163360178(.A(n_54883), .B(n_28623), .C(n_54865), .D(n_29799
		), .Z(n_179765326));
	notech_ao4 i_163560176(.A(n_32252), .B(n_310491719), .C(n_310391720), .D
		(n_28015), .Z(n_179565324));
	notech_and4 i_164360168(.A(n_179265321), .B(n_179065319), .C(n_178965318
		), .D(n_129164820), .Z(n_179465323));
	notech_ao4 i_163860173(.A(n_147128748), .B(n_29591), .C(n_147028747), .D
		(\nbus_11358[30] ), .Z(n_179265321));
	notech_ao4 i_164060171(.A(n_302991794), .B(n_147228749), .C(n_146928746)
		, .D(\nbus_11365[30] ), .Z(n_179065319));
	notech_ao4 i_164160170(.A(n_60166), .B(n_27187), .C(n_301791806), .D(n_30809
		), .Z(n_178965318));
	notech_and4 i_167360138(.A(n_129964828), .B(n_178565314), .C(n_129664825
		), .D(n_26754), .Z(n_178865317));
	notech_ao4 i_167160140(.A(n_154831963), .B(n_59980), .C(n_26929), .D(n_29681
		), .Z(n_178565314));
	notech_ao4 i_167460137(.A(n_57875), .B(\nbus_11358[21] ), .C(n_58147), .D
		(n_60004), .Z(n_178365312));
	notech_ao4 i_167560136(.A(n_151931934), .B(n_110964638), .C(n_58498), .D
		(n_111164640), .Z(n_178165310));
	notech_and3 i_170660106(.A(n_130692198), .B(n_62935425), .C(n_177865307)
		, .Z(n_177965308));
	notech_ao4 i_170560107(.A(n_27334), .B(n_29801), .C(n_27335), .D(n_29800
		), .Z(n_177865307));
	notech_ao4 i_170760105(.A(n_185068867), .B(n_31307), .C(n_300891815), .D
		(n_31279), .Z(n_177665305));
	notech_and4 i_171960097(.A(n_131264841), .B(n_177365302), .C(n_177165300
		), .D(n_177065299), .Z(n_177565304));
	notech_ao4 i_171060102(.A(n_58383), .B(n_27990), .C(n_60166), .D(n_27197
		), .Z(n_177365302));
	notech_ao4 i_171560100(.A(n_58002), .B(n_303191792), .C(n_58001), .D(n_29614
		), .Z(n_177165300));
	notech_ao4 i_171660099(.A(\nbus_11358[7] ), .B(n_112664655), .C(\nbus_11307[7] 
		), .D(n_26594), .Z(n_177065299));
	notech_and4 i_172360093(.A(n_168265211), .B(n_176665295), .C(n_131764846
		), .D(n_132064849), .Z(n_176965298));
	notech_ao4 i_172160095(.A(n_27348), .B(n_291963186), .C(n_27157), .D(n_189962171
		), .Z(n_176665295));
	notech_and4 i_172860088(.A(n_176365292), .B(n_176165290), .C(n_132364852
		), .D(n_132664855), .Z(n_176565294));
	notech_ao4 i_172460092(.A(n_56548), .B(n_113864667), .C(n_60016), .D(n_174165270
		), .Z(n_176365292));
	notech_ao4 i_172660090(.A(\nbus_11307[9] ), .B(n_26750), .C(n_27349), .D
		(n_112864657), .Z(n_176165290));
	notech_and3 i_177260051(.A(n_164365172), .B(n_175865287), .C(n_114764676
		), .Z(n_175965288));
	notech_ao4 i_177160052(.A(n_27334), .B(n_29803), .C(n_27335), .D(n_29802
		), .Z(n_175865287));
	notech_ao4 i_177360050(.A(n_27142), .B(n_59963), .C(n_27348), .D(n_298266511
		), .Z(n_175665285));
	notech_ao4 i_177460049(.A(n_302591798), .B(n_27999), .C(n_27349), .D(n_298166510
		), .Z(n_175565284));
	notech_and4 i_178260041(.A(n_175265281), .B(n_175065279), .C(n_174965278
		), .D(n_133564864), .Z(n_175465283));
	notech_ao4 i_177760046(.A(n_302691797), .B(\nbus_11307[14] ), .C(n_51735313
		), .D(n_298366512), .Z(n_175265281));
	notech_ao4 i_177960044(.A(n_60166), .B(n_27203), .C(n_27157), .D(n_157165100
		), .Z(n_175065279));
	notech_ao4 i_178060043(.A(n_52135317), .B(n_56257), .C(n_60011), .D(n_52335319
		), .Z(n_174965278));
	notech_and4 i_178960035(.A(n_162765156), .B(n_174565274), .C(n_134064869
		), .D(n_134364872), .Z(n_174865277));
	notech_ao4 i_178760037(.A(n_298466513), .B(n_27348), .C(n_60166), .D(n_27204
		), .Z(n_174565274));
	notech_and4 i_179460030(.A(n_174265271), .B(n_173965268), .C(n_134664875
		), .D(n_134964878), .Z(n_174465273));
	notech_ao4 i_179060034(.A(n_56548), .B(n_320137996), .C(n_60010), .D(n_174165270
		), .Z(n_174265271));
	notech_nand2 i_361720(.A(n_27344), .B(n_26591), .Z(n_174165270));
	notech_ao4 i_179260032(.A(\nbus_11358[15] ), .B(n_26751), .C(n_27349), .D
		(n_113264661), .Z(n_173965268));
	notech_and4 i_179960025(.A(n_173665265), .B(n_173465263), .C(n_135264881
		), .D(n_135564884), .Z(n_173865267));
	notech_ao4 i_179560029(.A(n_54658), .B(n_29804), .C(n_32270), .D(n_28110
		), .Z(n_173665265));
	notech_ao4 i_179760027(.A(n_27319), .B(n_28006), .C(n_144428721), .D(n_59980
		), .Z(n_173465263));
	notech_and4 i_180760019(.A(n_173165260), .B(n_172965258), .C(n_172865257
		), .D(n_135864887), .Z(n_173365262));
	notech_ao4 i_180060024(.A(n_144928726), .B(\nbus_11358[21] ), .C(n_145128728
		), .D(n_60004), .Z(n_173165260));
	notech_ao4 i_180460022(.A(n_57160), .B(\nbus_11365[21] ), .C(n_60162), .D
		(n_27210), .Z(n_172965258));
	notech_ao4 i_180560021(.A(n_27329), .B(n_110964638), .C(n_303791786), .D
		(n_111164640), .Z(n_172865257));
	notech_ao4 i_183759990(.A(n_307991744), .B(n_298466513), .C(n_55735), .D
		(n_58622), .Z(n_172665255));
	notech_ao4 i_183859989(.A(n_57490), .B(\nbus_11358[15] ), .C(n_184968866
		), .D(n_28104), .Z(n_172465253));
	notech_and3 i_184459983(.A(n_172065249), .B(n_172265251), .C(n_137264901
		), .Z(n_172365252));
	notech_ao4 i_184159986(.A(n_60010), .B(n_57775), .C(n_57627), .D(n_29754
		), .Z(n_172265251));
	notech_ao4 i_184259985(.A(n_26649), .B(n_58105), .C(n_111064639), .D(n_171965248
		), .Z(n_172065249));
	notech_nao3 i_184659982(.A(n_246591944), .B(n_57068), .C(n_57715), .Z(n_171965248
		));
	notech_ao4 i_184759981(.A(n_55726), .B(n_28110), .C(n_249866027), .D(n_26595
		), .Z(n_171765246));
	notech_ao4 i_184859980(.A(n_309891725), .B(n_59980), .C(n_142928706), .D
		(n_29681), .Z(n_171565244));
	notech_and3 i_185459974(.A(n_171165240), .B(n_171365242), .C(n_138264911
		), .Z(n_171465243));
	notech_ao4 i_185159977(.A(n_142828705), .B(\nbus_11358[21] ), .C(n_143028707
		), .D(n_60004), .Z(n_171365242));
	notech_ao4 i_185259976(.A(n_295269964), .B(n_110964638), .C(n_304991774)
		, .D(n_111164640), .Z(n_171165240));
	notech_and4 i_186859961(.A(n_170865237), .B(n_170665235), .C(n_170565234
		), .D(n_138564914), .Z(n_171065239));
	notech_ao4 i_186259966(.A(n_28236), .B(n_298066509), .C(n_28234), .D(n_297966508
		), .Z(n_170865237));
	notech_ao4 i_186459964(.A(n_59992), .B(n_28502), .C(n_303291791), .D(n_27983
		), .Z(n_170665235));
	notech_ao4 i_186559963(.A(n_297666505), .B(n_28544), .C(n_32270), .D(n_28090
		), .Z(n_170565234));
	notech_and4 i_187559954(.A(n_170265231), .B(n_170165230), .C(n_169965228
		), .D(n_169865227), .Z(n_170465233));
	notech_ao4 i_186959960(.A(n_28527), .B(n_29806), .C(n_54649), .D(n_29805
		), .Z(n_170265231));
	notech_ao4 i_187059959(.A(n_60162), .B(n_27218), .C(n_300091823), .D(n_60024
		), .Z(n_170165230));
	notech_ao4 i_187259957(.A(n_300291821), .B(n_29678), .C(n_268266211), .D
		(\nbus_11358[1] ), .Z(n_169965228));
	notech_ao4 i_187359956(.A(n_268366212), .B(\nbus_11307[1] ), .C(n_297866507
		), .D(n_111664645), .Z(n_169865227));
	notech_and4 i_188159948(.A(n_169565224), .B(n_169365222), .C(n_169265221
		), .D(n_140064929), .Z(n_169765226));
	notech_ao4 i_187659953(.A(n_291863185), .B(n_28236), .C(n_291763184), .D
		(n_28234), .Z(n_169565224));
	notech_ao4 i_187859951(.A(n_5723), .B(n_28502), .C(n_27986), .D(n_303291791
		), .Z(n_169365222));
	notech_ao4 i_187959950(.A(n_291463181), .B(n_28544), .C(n_32270), .D(n_28093
		), .Z(n_169265221));
	notech_and4 i_188859941(.A(n_168965218), .B(n_168865217), .C(n_168665215
		), .D(n_168565214), .Z(n_169165220));
	notech_ao4 i_188259947(.A(n_28527), .B(n_29808), .C(n_54649), .D(n_29807
		), .Z(n_168965218));
	notech_ao4 i_188359946(.A(n_60162), .B(n_27220), .C(n_300091823), .D(n_5743
		), .Z(n_168865217));
	notech_ao4 i_188559944(.A(n_300291821), .B(n_29725), .C(n_268266211), .D
		(\nbus_11358[4] ), .Z(n_168665215));
	notech_ao4 i_188659943(.A(n_268366212), .B(\nbus_11307[4] ), .C(n_291663183
		), .D(n_111664645), .Z(n_168565214));
	notech_and4 i_190759926(.A(n_141364942), .B(n_168265211), .C(n_141664945
		), .D(n_167965208), .Z(n_168465213));
	notech_and2 i_157061745(.A(n_120264731), .B(n_114064669), .Z(n_168265211
		));
	notech_ao4 i_190559928(.A(n_54649), .B(n_29809), .C(n_60166), .D(n_27225
		), .Z(n_167965208));
	notech_ao4 i_190859925(.A(n_60016), .B(n_301891805), .C(n_28545), .D(n_113764666
		), .Z(n_167665205));
	notech_and2 i_191159922(.A(n_167465203), .B(n_142264951), .Z(n_167565204
		));
	notech_ao4 i_191059923(.A(\nbus_11307[9] ), .B(n_26749), .C(n_113464663)
		, .D(n_167365202), .Z(n_167465203));
	notech_nao3 i_191459919(.A(n_30946), .B(n_28552), .C(n_189962171), .Z(n_167365202
		));
	notech_and3 i_191659917(.A(n_65435450), .B(n_167065199), .C(n_130992195)
		, .Z(n_167165200));
	notech_ao4 i_191559918(.A(n_30088), .B(n_292166450), .C(n_302891795), .D
		(n_297466503), .Z(n_167065199));
	notech_ao4 i_191759916(.A(\nbus_11358[11] ), .B(n_26667), .C(n_292566454
		), .D(\nbus_11307[11] ), .Z(n_166865197));
	notech_ao4 i_191859915(.A(n_292466453), .B(n_27996), .C(n_31456), .D(n_28545
		), .Z(n_166765196));
	notech_and4 i_192859907(.A(n_143164960), .B(n_166465193), .C(n_166265191
		), .D(n_166165190), .Z(n_166665195));
	notech_ao4 i_192259912(.A(n_28527), .B(n_29811), .C(n_54649), .D(n_29810
		), .Z(n_166465193));
	notech_ao4 i_192559910(.A(n_31492), .B(n_191265441), .C(n_60166), .D(n_27227
		), .Z(n_166265191));
	notech_ao4 i_192659909(.A(n_302491799), .B(n_163365162), .C(n_163165160)
		, .D(n_29596), .Z(n_166165190));
	notech_and3 i_193059905(.A(n_111364642), .B(n_114664675), .C(n_165865187
		), .Z(n_165965188));
	notech_ao4 i_192959906(.A(n_301691807), .B(n_297466503), .C(n_28527), .D
		(n_29812), .Z(n_165865187));
	notech_ao4 i_193159904(.A(n_54649), .B(n_29813), .C(n_31560), .D(n_297566504
		), .Z(n_165565184));
	notech_ao4 i_193259903(.A(n_27998), .B(n_292466453), .C(n_31540), .D(n_28545
		), .Z(n_165465183));
	notech_and4 i_194159895(.A(n_165165180), .B(n_164965178), .C(n_164865177
		), .D(n_144464973), .Z(n_165365182));
	notech_ao4 i_193659900(.A(n_292566454), .B(\nbus_11307[13] ), .C(n_31576
		), .D(n_191265441), .Z(n_165165180));
	notech_ao4 i_193859898(.A(n_60166), .B(n_27229), .C(n_30109), .D(n_292166450
		), .Z(n_164965178));
	notech_ao4 i_193959897(.A(n_302091803), .B(n_163365162), .C(n_163165160)
		, .D(n_29592), .Z(n_164865177));
	notech_and3 i_194359893(.A(n_164365172), .B(n_114764676), .C(n_164565174
		), .Z(n_164665175));
	notech_ao4 i_194259894(.A(n_59963), .B(n_297466503), .C(n_28527), .D(n_29814
		), .Z(n_164565174));
	notech_ao4 i_114561757(.A(n_102135817), .B(n_60011), .C(n_102035816), .D
		(n_56257), .Z(n_164365172));
	notech_ao4 i_194459892(.A(n_54649), .B(n_29815), .C(n_298266511), .D(n_297566504
		), .Z(n_164165170));
	notech_ao4 i_194559891(.A(n_292466453), .B(n_27999), .C(n_28545), .D(n_298166510
		), .Z(n_164065169));
	notech_and4 i_195359883(.A(n_163765166), .B(n_163565164), .C(n_163465163
		), .D(n_145764986), .Z(n_163965168));
	notech_ao4 i_194859888(.A(\nbus_11307[14] ), .B(n_292566454), .C(n_298366512
		), .D(n_191265441), .Z(n_163765166));
	notech_ao4 i_195059886(.A(n_60166), .B(n_27230), .C(n_292166450), .D(n_157165100
		), .Z(n_163565164));
	notech_ao4 i_195159885(.A(n_60011), .B(n_163365162), .C(n_56257), .D(n_163165160
		), .Z(n_163465163));
	notech_nao3 i_173761738(.A(n_32612), .B(n_26683), .C(n_304191782), .Z(n_163365162
		));
	notech_nao3 i_173961737(.A(n_59349), .B(n_26683), .C(n_304191782), .Z(n_163165160
		));
	notech_and4 i_195959877(.A(n_146264991), .B(n_162465153), .C(n_162765156
		), .D(n_146564994), .Z(n_162965158));
	notech_and2 i_170161744(.A(n_162665155), .B(n_115264681), .Z(n_162765156
		));
	notech_ao4 i_80461764(.A(n_299591828), .B(\nbus_11358[15] ), .C(n_61115)
		, .D(n_316137956), .Z(n_162665155));
	notech_ao4 i_195759879(.A(n_298466513), .B(n_297566504), .C(n_60166), .D
		(n_27231), .Z(n_162465153));
	notech_ao4 i_196059876(.A(n_60010), .B(n_301891805), .C(\nbus_11307[15] 
		), .D(n_26749), .Z(n_162165150));
	notech_ao3 i_196359873(.A(n_146964998), .B(n_147165000), .C(n_147064999)
		, .Z(n_162065149));
	notech_and4 i_197059866(.A(n_161565144), .B(n_161365142), .C(n_135064879
		), .D(n_147665005), .Z(n_161765146));
	notech_ao4 i_196659870(.A(n_28527), .B(n_29817), .C(n_54649), .D(n_29816
		), .Z(n_161565144));
	notech_ao4 i_196859868(.A(n_303591788), .B(n_28006), .C(n_139728674), .D
		(n_59980), .Z(n_161365142));
	notech_and4 i_197659860(.A(n_161065139), .B(n_160865137), .C(n_160765136
		), .D(n_147965008), .Z(n_161265141));
	notech_ao4 i_197159865(.A(n_140228679), .B(\nbus_11358[21] ), .C(n_140428681
		), .D(n_60004), .Z(n_161065139));
	notech_ao4 i_197359863(.A(n_233165860), .B(\nbus_11365[21] ), .C(n_60167
		), .D(n_27238), .Z(n_160865137));
	notech_ao4 i_197459862(.A(n_110964638), .B(n_309691727), .C(n_301091813)
		, .D(n_111164640), .Z(n_160765136));
	notech_and4 i_198159855(.A(n_160465133), .B(n_160265131), .C(n_148665015
		), .D(n_148965018), .Z(n_160665135));
	notech_ao4 i_197759859(.A(n_28527), .B(n_29819), .C(n_54649), .D(n_29818
		), .Z(n_160465133));
	notech_ao4 i_197959857(.A(n_32252), .B(n_26678), .C(n_303591788), .D(n_28015
		), .Z(n_160265131));
	notech_and4 i_198659850(.A(n_159965128), .B(n_159765126), .C(n_149265021
		), .D(n_149565024), .Z(n_160165130));
	notech_ao4 i_198259854(.A(n_140328680), .B(n_29591), .C(n_140228679), .D
		(\nbus_11358[30] ), .Z(n_159965128));
	notech_ao4 i_198459852(.A(n_140128678), .B(\nbus_11365[30] ), .C(n_60167
		), .D(n_27244), .Z(n_159765126));
	notech_and4 i_201659820(.A(n_159365122), .B(n_149665025), .C(n_26754), .D
		(n_149965028), .Z(n_159665125));
	notech_ao4 i_201459822(.A(n_57873), .B(\nbus_11358[21] ), .C(n_58145), .D
		(n_60004), .Z(n_159365122));
	notech_ao4 i_201759819(.A(n_138168398), .B(\nbus_11365[21] ), .C(n_58497
		), .D(n_111164640), .Z(n_159165120));
	notech_ao4 i_201859818(.A(n_321438009), .B(n_28006), .C(n_110964638), .D
		(n_319937994), .Z(n_158965118));
	notech_nand2 i_206159777(.A(n_158565114), .B(n_150865037), .Z(n_158665115
		));
	notech_ao4 i_206059778(.A(n_58427), .B(n_28006), .C(n_305924323), .D(n_59980
		), .Z(n_158565114));
	notech_and4 i_206759771(.A(n_158265111), .B(n_158065109), .C(n_151165040
		), .D(n_151465043), .Z(n_158465113));
	notech_ao4 i_206359775(.A(n_57877), .B(\nbus_11358[21] ), .C(n_58143), .D
		(n_60004), .Z(n_158265111));
	notech_ao4 i_206559773(.A(n_306124325), .B(n_110964638), .C(n_58493), .D
		(n_111164640), .Z(n_158065109));
	notech_and4 i_213859700(.A(n_151865047), .B(n_157665105), .C(n_151565044
		), .D(n_26754), .Z(n_157965108));
	notech_ao4 i_213659702(.A(n_306824332), .B(n_59980), .C(n_307324337), .D
		(n_29681), .Z(n_157665105));
	notech_ao4 i_213959699(.A(n_57864), .B(\nbus_11358[21] ), .C(n_58141), .D
		(n_60004), .Z(n_157465103));
	notech_ao4 i_214059698(.A(n_306624330), .B(n_110964638), .C(n_58494), .D
		(n_111164640), .Z(n_157265101));
	notech_nand2 i_4061778(.A(opc[14]), .B(n_62806), .Z(n_157165100));
	notech_ao4 i_218059658(.A(n_58424), .B(n_28006), .C(n_287827260), .D(n_59980
		), .Z(n_156865097));
	notech_nand3 i_218559653(.A(n_156465093), .B(n_156665095), .C(n_153165060
		), .Z(n_156765096));
	notech_ao4 i_218259656(.A(n_26615), .B(n_29681), .C(n_57863), .D(\nbus_11358[21] 
		), .Z(n_156665095));
	notech_ao4 i_218359655(.A(n_57861), .B(\nbus_11365[21] ), .C(n_286827250
		), .D(n_110964638), .Z(n_156465093));
	notech_and4 i_222059618(.A(n_156065089), .B(n_153265061), .C(n_26754), .D
		(n_153565064), .Z(n_156365092));
	notech_ao4 i_221859620(.A(n_57865), .B(n_56329), .C(n_57867), .D(\nbus_11365[21] 
		), .Z(n_156065089));
	notech_ao4 i_222159617(.A(n_58008), .B(n_249866027), .C(n_58138), .D(n_60004
		), .Z(n_155865087));
	notech_ao4 i_222259616(.A(n_305624320), .B(n_59980), .C(n_58007), .D(n_110964638
		), .Z(n_155665085));
	notech_ao4 i_224259596(.A(n_30594), .B(n_29754), .C(n_27305), .D(\nbus_11307[15] 
		), .Z(n_155565084));
	notech_ao4 i_224359595(.A(n_60331), .B(n_28110), .C(n_309591728), .D(n_29681
		), .Z(n_155465083));
	notech_ao4 i_224459594(.A(n_30803), .B(n_60004), .C(n_309491729), .D(\nbus_11365[21] 
		), .Z(n_155265081));
	notech_or2 i_161722(.A(n_26616), .B(n_319291631), .Z(n_155165080));
	notech_or4 i_123160562(.A(n_56834), .B(n_26962), .C(n_61142), .D(n_56619
		), .Z(n_154865077));
	notech_nor2 i_120360588(.A(n_304691777), .B(n_56329), .Z(n_154765076));
	notech_or4 i_116860623(.A(n_56834), .B(n_56939), .C(n_26969), .D(n_28006
		), .Z(n_154065069));
	notech_or2 i_117360618(.A(n_57726), .B(n_28147), .Z(n_153565064));
	notech_nand2 i_117460617(.A(n_57569), .B(\regs_13_14[21] ), .Z(n_153265061
		));
	notech_or2 i_111460669(.A(n_58139), .B(n_60004), .Z(n_153165060));
	notech_ao3 i_111960664(.A(opc[21]), .B(n_62806), .C(n_286927251), .Z(n_152465053
		));
	notech_nao3 i_105560718(.A(n_26792), .B(opa[21]), .C(n_58494), .Z(n_152365052
		));
	notech_or4 i_106260713(.A(n_56832), .B(n_56939), .C(n_26922), .D(n_28006
		), .Z(n_151865047));
	notech_or4 i_106360712(.A(n_58805), .B(n_58494), .C(nbus_11295[21]), .D(n_60938
		), .Z(n_151565044));
	notech_or2 i_95860803(.A(n_286869880), .B(\nbus_11365[21] ), .Z(n_151465043
		));
	notech_nand2 i_96160800(.A(n_58144), .B(\regs_13_14[21] ), .Z(n_151165040
		));
	notech_or4 i_96460797(.A(n_58806), .B(n_58493), .C(nbus_11295[21]), .D(n_60938
		), .Z(n_150865037));
	notech_nor2 i_96560796(.A(n_154331958), .B(nbus_11295[21]), .Z(n_150565034
		));
	notech_or2 i_90660852(.A(n_321538010), .B(n_59980), .Z(n_150465033));
	notech_nand2 i_91360847(.A(n_58146), .B(\regs_13_14[21] ), .Z(n_149965028
		));
	notech_or4 i_91460846(.A(n_58497), .B(n_58810), .C(nbus_11295[21]), .D(n_60938
		), .Z(n_149665025));
	notech_or2 i_86460893(.A(n_140428681), .B(n_302991794), .Z(n_149565024)
		);
	notech_or2 i_86760890(.A(n_139728674), .B(n_303091793), .Z(n_149265021)
		);
	notech_nao3 i_87060887(.A(n_62798), .B(opc_10[30]), .C(n_309691727), .Z(n_148965018
		));
	notech_nand3 i_87360884(.A(n_60167), .B(n_60246), .C(read_data[30]), .Z(n_148665015
		));
	notech_or2 i_85560902(.A(n_140328680), .B(n_29681), .Z(n_147965008));
	notech_nand3 i_85860899(.A(opc[21]), .B(n_62822), .C(n_309791726), .Z(n_147665005
		));
	notech_nand2 i_83460922(.A(n_113664665), .B(opb[15]), .Z(n_147165000));
	notech_ao4 i_83360923(.A(n_234791985), .B(n_1427), .C(n_26646), .D(n_115164680
		), .Z(n_147064999));
	notech_or4 i_83260924(.A(n_26890), .B(n_113464663), .C(nbus_11295[15]), 
		.D(n_60938), .Z(n_146964998));
	notech_or2 i_83760919(.A(n_27036), .B(n_320137996), .Z(n_146864997));
	notech_nand3 i_84060916(.A(n_1430), .B(n_6380), .C(\eflags[10] ), .Z(n_146564994
		));
	notech_nand3 i_84160915(.A(n_1430), .B(n_6379), .C(n_56163), .Z(n_146264991
		));
	notech_nand2 i_82260934(.A(n_292666455), .B(opb[14]), .Z(n_145764986));
	notech_nand2 i_80760948(.A(opb[13]), .B(n_292666455), .Z(n_144464973));
	notech_or4 i_79060964(.A(n_26890), .B(n_60938), .C(n_28137), .D(n_28545)
		, .Z(n_143164960));
	notech_nand2 i_77160983(.A(opb[9]), .B(n_113664665), .Z(n_142264951));
	notech_or2 i_77460980(.A(n_113864667), .B(n_27036), .Z(n_141964948));
	notech_nand3 i_77760977(.A(n_1430), .B(n_6367), .C(n_56163), .Z(n_141664945
		));
	notech_or4 i_77860976(.A(n_26890), .B(n_28135), .C(n_60938), .D(n_28545)
		, .Z(n_141364942));
	notech_or4 i_75061002(.A(n_62858), .B(n_303891785), .C(n_62822), .D(\nbus_11307[4] 
		), .Z(n_140064929));
	notech_or4 i_73561017(.A(n_62858), .B(n_303891785), .C(n_62822), .D(\nbus_11307[1] 
		), .Z(n_138564914));
	notech_or2 i_70461048(.A(n_57935), .B(\nbus_11365[21] ), .Z(n_138264911)
		);
	notech_or4 i_70961043(.A(n_56832), .B(n_56939), .C(n_26649), .D(n_28006)
		, .Z(n_137764906));
	notech_nand2 i_69461058(.A(n_57481), .B(opa[15]), .Z(n_137264901));
	notech_or4 i_69961053(.A(n_56832), .B(n_56983), .C(n_26649), .D(n_28000)
		, .Z(n_136764896));
	notech_or2 i_64361102(.A(n_145028727), .B(n_29681), .Z(n_135864887));
	notech_nand3 i_64661099(.A(opc[21]), .B(n_62806), .C(n_27340), .Z(n_135564884
		));
	notech_nand3 i_64961096(.A(n_1429), .B(n_7324), .C(\eflags[10] ), .Z(n_135264881
		));
	notech_nand3 i_64761098(.A(n_60167), .B(n_60246), .C(read_data[21]), .Z(n_135064879
		));
	notech_nand2 i_62461117(.A(opa[15]), .B(n_112964658), .Z(n_134964878));
	notech_nao3 i_62761114(.A(opc[15]), .B(n_62806), .C(n_27157), .Z(n_134664875
		));
	notech_nand3 i_63261111(.A(n_1429), .B(n_7311), .C(n_56163), .Z(n_134364872
		));
	notech_nand3 i_63361110(.A(n_1429), .B(n_7312), .C(\eflags[10] ), .Z(n_134064869
		));
	notech_nand2 i_61561126(.A(n_27289), .B(opb[14]), .Z(n_133564864));
	notech_nand2 i_55261179(.A(opb[9]), .B(n_113064659), .Z(n_132664855));
	notech_nand2 i_55561176(.A(sav_esi[9]), .B(n_61142), .Z(n_132364852));
	notech_nand3 i_55961173(.A(n_1429), .B(n_7299), .C(n_56163), .Z(n_132064849
		));
	notech_nand3 i_56061172(.A(n_1429), .B(n_7300), .C(\eflags[10] ), .Z(n_131764846
		));
	notech_or4 i_54361188(.A(n_32356), .B(n_56548), .C(n_303391790), .D(n_61138
		), .Z(n_131264841));
	notech_or4 i_54661185(.A(n_300891815), .B(n_31309), .C(n_26770), .D(n_27712
		), .Z(n_130964838));
	notech_or2 i_50061231(.A(n_241372893), .B(\nbus_11365[21] ), .Z(n_130464833
		));
	notech_or4 i_50561226(.A(n_246891941), .B(n_2479), .C(n_56688), .D(n_28006
		), .Z(n_129964828));
	notech_or4 i_50661225(.A(n_58802), .B(n_58498), .C(nbus_11295[21]), .D(n_60938
		), .Z(n_129664825));
	notech_or2 i_46061269(.A(n_303091793), .B(n_146428741), .Z(n_129164820)
		);
	notech_or4 i_46361266(.A(n_32555), .B(n_61138), .C(n_60331), .D(n_28121)
		, .Z(n_128864817));
	notech_or2 i_46661263(.A(n_310191722), .B(n_27485), .Z(n_128564814));
	notech_or2 i_44661283(.A(n_147128748), .B(n_29681), .Z(n_127864807));
	notech_or2 i_45361276(.A(n_54894), .B(n_27465), .Z(n_127164800));
	notech_nand2 i_43361296(.A(sav_esp[15]), .B(n_61138), .Z(n_126464793));
	notech_nand2 i_43661293(.A(n_7364), .B(n_26986), .Z(n_126164790));
	notech_ao4 i_133468528(.A(n_326990767), .B(n_60023), .C(n_56390), .D(n_27426
		), .Z(n_110271582));
	notech_ao4 i_133368529(.A(n_326790765), .B(n_27730), .C(n_326890766), .D
		(n_27768), .Z(n_110371583));
	notech_ao4 i_130468558(.A(n_326990767), .B(n_60008), .C(n_56390), .D(n_27457
		), .Z(n_110471584));
	notech_ao4 i_130368559(.A(n_326790765), .B(n_27747), .C(n_326890766), .D
		(n_27788), .Z(n_110571585));
	notech_ao4 i_130268560(.A(n_326990767), .B(n_60006), .C(n_56391), .D(n_27461
		), .Z(n_110671586));
	notech_ao4 i_130168561(.A(n_326790765), .B(n_27749), .C(n_326890766), .D
		(n_27790), .Z(n_110771587));
	notech_ao4 i_130068562(.A(n_326990767), .B(n_60005), .C(n_56391), .D(n_27463
		), .Z(n_110871588));
	notech_ao4 i_129968563(.A(n_326790765), .B(n_27750), .C(n_326890766), .D
		(n_27791), .Z(n_110971589));
	notech_nand2 i_40467023(.A(n_329263509), .B(imm[4]), .Z(n_111071590));
	notech_or4 i_40367024(.A(opz[0]), .B(opz[1]), .C(n_28051), .D(n_26651), 
		.Z(n_111171591));
	notech_and2 i_40767020(.A(n_329263509), .B(imm[5]), .Z(n_111271592));
	notech_ao4 i_615643(.A(n_62041235), .B(n_28094), .C(n_317887452), .D(n_28392
		), .Z(n_22745));
	notech_or2 i_158967433(.A(n_111271592), .B(n_83341448), .Z(\nbus_11317[5] 
		));
	notech_nor2 i_112366305(.A(n_112271602), .B(n_27987), .Z(n_112171601));
	notech_and2 i_7267329(.A(n_115671636), .B(n_115771637), .Z(n_112271602)
		);
	notech_ao4 i_7167330(.A(n_25140866), .B(n_115871638), .C(n_330063517), .D
		(opd[4]), .Z(n_112371603));
	notech_nao3 i_111966309(.A(n_9241), .B(n_60331), .C(n_60051), .Z(n_113071610
		));
	notech_ao4 i_112066308(.A(n_111271592), .B(n_83341448), .C(n_121261495),
		 .D(n_26781), .Z(n_113171611));
	notech_nand2 i_112266306(.A(add_src[5]), .B(n_26723), .Z(n_113271612));
	notech_nor2 i_112166307(.A(n_24540860), .B(n_28094), .Z(n_113371613));
	notech_nor2 i_112466304(.A(n_112371603), .B(opd[5]), .Z(n_113471614));
	notech_or4 i_612923(.A(n_116671646), .B(n_113471614), .C(n_112171601), .D
		(n_113371613), .Z(n_25973));
	notech_or2 i_114766281(.A(n_115671636), .B(n_27986), .Z(n_113671616));
	notech_ao4 i_7367328(.A(n_25140866), .B(n_27985), .C(n_330963526), .D(n_25540870
		), .Z(n_113771617));
	notech_nao3 i_114366285(.A(n_9236), .B(n_60331), .C(n_60051), .Z(n_114471624
		));
	notech_or2 i_114466284(.A(n_29904), .B(n_329363510), .Z(n_114571625));
	notech_nand2 i_114666282(.A(add_src[4]), .B(n_26723), .Z(n_114671626));
	notech_or2 i_114566283(.A(n_24540860), .B(n_28093), .Z(n_114771627));
	notech_or2 i_114866280(.A(n_113771617), .B(opd[4]), .Z(n_114871628));
	notech_nand3 i_512922(.A(n_117771657), .B(n_114871628), .C(n_113671616),
		 .Z(n_25968));
	notech_nand2 i_149965930(.A(write_data_33[5]), .B(n_60246), .Z(n_115371633
		));
	notech_nand3 i_618811(.A(n_118071660), .B(n_117971659), .C(n_115371633),
		 .Z(n_25729));
	notech_mux2 i_1767383(.S(opd[3]), .A(n_55508), .B(n_27040885), .Z(n_115571635
		));
	notech_and2 i_3467367(.A(n_115571635), .B(n_26785), .Z(n_115671636));
	notech_mux2 i_110966319(.S(opd[4]), .A(n_55508), .B(n_27040885), .Z(n_115771637
		));
	notech_nand2 i_111266316(.A(opd[4]), .B(opd[3]), .Z(n_115871638));
	notech_ao4 i_112566303(.A(n_40241017), .B(n_29091), .C(n_39041005), .D(n_28931
		), .Z(n_115971639));
	notech_ao4 i_112666302(.A(n_53841153), .B(n_29900), .C(n_54141156), .D(n_29899
		), .Z(n_116171641));
	notech_ao4 i_112766301(.A(n_53341148), .B(nbus_11295[5]), .C(n_53641151)
		, .D(\nbus_11307[5] ), .Z(n_116271642));
	notech_and4 i_113066298(.A(n_116271642), .B(n_116171641), .C(n_115971639
		), .D(n_113071610), .Z(n_116471644));
	notech_nao3 i_113266296(.A(n_116471644), .B(n_113271612), .C(n_113171611
		), .Z(n_116671646));
	notech_ao4 i_114966279(.A(n_40241017), .B(n_29090), .C(n_39041005), .D(n_28930
		), .Z(n_116971649));
	notech_ao4 i_115066278(.A(n_53841153), .B(n_29903), .C(n_54141156), .D(n_29901
		), .Z(n_117171651));
	notech_ao4 i_115166277(.A(n_53341148), .B(nbus_11295[4]), .C(n_53641151)
		, .D(\nbus_11307[4] ), .Z(n_117271652));
	notech_and4 i_115466274(.A(n_117271652), .B(n_117171651), .C(n_116971649
		), .D(n_114471624), .Z(n_117471654));
	notech_and4 i_115766271(.A(n_117471654), .B(n_114571625), .C(n_114671626
		), .D(n_114771627), .Z(n_117771657));
	notech_ao4 i_150165928(.A(n_318291641), .B(\nbus_11358[5] ), .C(n_318391640
		), .D(nbus_11295[5]), .Z(n_117971659));
	notech_ao4 i_150065929(.A(n_315391670), .B(n_27863), .C(n_59152), .D(n_28456
		), .Z(n_118071660));
	notech_ao4 i_16264292(.A(\nbus_11307[7] ), .B(n_26895), .C(\nbus_11358[7] 
		), .D(n_57758), .Z(n_118271662));
	notech_and3 i_16364291(.A(n_322373703), .B(n_58084), .C(n_120171681), .Z
		(n_118371663));
	notech_nand2 i_16064294(.A(n_58717), .B(n_125371733), .Z(n_118671666));
	notech_ao4 i_15364301(.A(n_59434), .B(\nbus_11307[7] ), .C(n_58573), .D(\nbus_11358[7] 
		), .Z(n_118871668));
	notech_and3 i_15464300(.A(n_58008), .B(n_58007), .C(n_57473), .Z(n_118971669
		));
	notech_or4 i_85963617(.A(n_101413114), .B(n_58100), .C(n_57229), .D(instrc
		[121]), .Z(n_119171671));
	notech_ao3 i_58263888(.A(n_26811), .B(\opa_12[7] ), .C(n_26812), .Z(n_119371673
		));
	notech_or4 i_57763893(.A(n_246891941), .B(n_2479), .C(n_56688), .D(n_27990
		), .Z(n_120071680));
	notech_or4 i_58563885(.A(n_57087), .B(n_29652), .C(n_26770), .D(n_58506)
		, .Z(n_120171681));
	notech_nao3 i_59663876(.A(opc[9]), .B(n_62806), .C(n_128571765), .Z(n_120271682
		));
	notech_or2 i_59463877(.A(n_60016), .B(n_57329), .Z(n_120571685));
	notech_or2 i_58863882(.A(n_58106), .B(n_26933), .Z(n_121071690));
	notech_or4 i_64863824(.A(n_62858), .B(n_58162), .C(n_62806), .D(n_57557)
		, .Z(n_121571695));
	notech_nao3 i_64563827(.A(opd[2]), .B(n_58078), .C(n_56921), .Z(n_121871698
		));
	notech_nao3 i_64063832(.A(n_58806), .B(n_118671666), .C(n_26804), .Z(n_121971699
		));
	notech_ao4 i_64163831(.A(n_305291771), .B(n_189362166), .C(n_26647), .D(n_125471734
		), .Z(n_122071700));
	notech_ao3 i_64263830(.A(n_62798), .B(opc[2]), .C(n_153279036), .Z(n_122171701
		));
	notech_and3 i_82763647(.A(n_59445), .B(\opa_12[7] ), .C(n_26808), .Z(n_122671706
		));
	notech_or4 i_82663648(.A(n_56832), .B(n_56939), .C(n_26969), .D(n_27990)
		, .Z(n_122971709));
	notech_or4 i_82363651(.A(n_30854), .B(n_245362720), .C(n_31309), .D(n_58488
		), .Z(n_123271712));
	notech_or4 i_82063654(.A(n_62858), .B(n_124171721), .C(n_60938), .D(\nbus_11307[7] 
		), .Z(n_123571715));
	notech_nao3 i_11864336(.A(n_56448), .B(n_56482), .C(n_58100), .Z(n_123671716
		));
	notech_nao3 i_29533(.A(n_319191632), .B(n_58078), .C(n_246891941), .Z(n_123771717
		));
	notech_nao3 i_7564378(.A(n_56457), .B(n_26731), .C(n_56529), .Z(n_123871718
		));
	notech_or4 i_12564329(.A(n_245362720), .B(n_56529), .C(n_57082), .D(n_29652
		), .Z(n_123971719));
	notech_or2 i_29516(.A(n_58815), .B(n_58488), .Z(n_124071720));
	notech_or2 i_8564368(.A(n_56529), .B(n_58815), .Z(n_124171721));
	notech_nao3 i_12264332(.A(n_32386), .B(n_32298), .C(n_56839), .Z(n_124271722
		));
	notech_ao4 i_154562952(.A(n_31307), .B(n_118971669), .C(n_56529), .D(n_118871668
		), .Z(n_124471724));
	notech_ao4 i_154362954(.A(n_123871718), .B(\nbus_11307[7] ), .C(n_154079044
		), .D(n_29614), .Z(n_124671726));
	notech_and4 i_154762950(.A(n_124671726), .B(n_123571715), .C(n_124471724
		), .D(n_123271712), .Z(n_124871728));
	notech_ao4 i_154062957(.A(n_57947), .B(n_26969), .C(n_303191792), .D(n_57470
		), .Z(n_124971729));
	notech_nand2 i_154162956(.A(n_124971729), .B(n_122971709), .Z(n_125071730
		));
	notech_mux2 i_139763095(.S(n_32325), .A(n_312347735), .B(n_312447734), .Z
		(n_125371733));
	notech_mux2 i_139663096(.S(n_32325), .A(n_26645), .B(n_26644), .Z(n_125471734
		));
	notech_ao3 i_139463098(.A(n_121971699), .B(n_26629), .C(n_122171701), .Z
		(n_125671736));
	notech_ao4 i_139163101(.A(n_153379037), .B(n_152572005), .C(n_153479038)
		, .D(n_57557), .Z(n_125771737));
	notech_ao4 i_138863104(.A(n_58047), .B(\nbus_11358[2] ), .C(n_59991), .D
		(n_153779041), .Z(n_126071740));
	notech_ao4 i_138663106(.A(n_257980080), .B(n_344366972), .C(n_154331958)
		, .D(nbus_11295[2]), .Z(n_126271742));
	notech_and4 i_139063102(.A(n_126271742), .B(n_126071740), .C(n_26672), .D
		(n_121571695), .Z(n_126471744));
	notech_ao4 i_133563156(.A(n_303673516), .B(n_27992), .C(n_58608), .D(n_58482
		), .Z(n_126571745));
	notech_ao4 i_133463157(.A(n_58054), .B(\nbus_11358[9] ), .C(\nbus_11307[9] 
		), .D(n_26679), .Z(n_126771747));
	notech_ao4 i_133163160(.A(n_325273732), .B(n_29743), .C(n_291963186), .D
		(n_322373703), .Z(n_126971749));
	notech_and4 i_133363158(.A(n_200065529), .B(n_126971749), .C(n_120271682
		), .D(n_120571685), .Z(n_127271752));
	notech_ao4 i_132663165(.A(n_31307), .B(n_118371663), .C(n_26852), .D(n_118271662
		), .Z(n_127471754));
	notech_ao4 i_132563166(.A(n_57947), .B(n_26933), .C(n_31279), .D(n_26812
		), .Z(n_127671756));
	notech_nand3 i_132863163(.A(n_127471754), .B(n_127671756), .C(n_120071680
		), .Z(n_127771757));
	notech_ao4 i_132363168(.A(n_303191792), .B(n_284880349), .C(n_31309), .D
		(n_57915), .Z(n_127871758));
	notech_and2 i_76661765(.A(n_128671766), .B(n_134171821), .Z(n_128171761)
		);
	notech_nand2 i_176061733(.A(n_58802), .B(n_26662), .Z(n_128371763));
	notech_nao3 i_181061729(.A(n_26664), .B(n_26662), .C(n_58184), .Z(n_128471764
		));
	notech_and2 i_150961785(.A(n_57915), .B(n_128771767), .Z(n_128571765));
	notech_or2 i_119760594(.A(n_58318), .B(\nbus_11358[15] ), .Z(n_128671766
		));
	notech_nao3 i_121160580(.A(n_57730), .B(n_30946), .C(n_30854), .Z(n_128771767
		));
	notech_or4 i_47661253(.A(n_58802), .B(n_60940), .C(n_28139), .D(n_58482)
		, .Z(n_132071800));
	notech_nand2 i_47561254(.A(opd[13]), .B(n_58378), .Z(n_132371803));
	notech_nand2 i_47261257(.A(opa[13]), .B(n_58055), .Z(n_132671806));
	notech_or4 i_46961260(.A(n_58184), .B(n_58482), .C(n_302091803), .D(n_26664
		), .Z(n_132971809));
	notech_or4 i_49661234(.A(n_58802), .B(n_28141), .C(n_60940), .D(n_58482)
		, .Z(n_133071810));
	notech_or4 i_49561235(.A(n_62858), .B(n_62806), .C(n_29754), .D(n_58482)
		, .Z(n_133371813));
	notech_nand2 i_49061240(.A(opa[15]), .B(n_58055), .Z(n_133871818));
	notech_mux2 i_224159597(.S(n_60329), .A(n_28104), .B(n_316137956), .Z(n_134171821
		));
	notech_ao4 i_166760144(.A(n_58105), .B(n_26933), .C(n_111064639), .D(n_128571765
		), .Z(n_134471824));
	notech_ao4 i_166660145(.A(n_60010), .B(n_57329), .C(n_29754), .D(n_325273732
		), .Z(n_134671826));
	notech_ao4 i_166360148(.A(n_303673516), .B(n_28000), .C(\nbus_11358[15] 
		), .D(n_58054), .Z(n_134871828));
	notech_and4 i_166560146(.A(n_128171761), .B(n_133071810), .C(n_134871828
		), .D(n_133371813), .Z(n_135171831));
	notech_ao4 i_165060161(.A(n_31576), .B(n_128371763), .C(n_128471764), .D
		(n_29592), .Z(n_135271832));
	notech_ao4 i_164860163(.A(n_30109), .B(n_58040), .C(n_94935745), .D(n_26933
		), .Z(n_135471834));
	notech_and4 i_165260159(.A(n_135471834), .B(n_135271832), .C(n_132671806
		), .D(n_132971809), .Z(n_135671836));
	notech_ao4 i_164560166(.A(n_58482), .B(n_31540), .C(n_58054), .D(\nbus_11358[13] 
		), .Z(n_135771837));
	notech_and4 i_164760164(.A(n_93835734), .B(n_135771837), .C(n_132071800)
		, .D(n_132371803), .Z(n_136071840));
	notech_ao4 i_153860269(.A(n_291763184), .B(n_111464643), .C(n_5723), .D(n_111564644
		), .Z(n_136171841));
	notech_ao4 i_153760270(.A(n_57999), .B(n_29725), .C(n_291563182), .D(n_56512
		), .Z(n_136271842));
	notech_ao4 i_153560272(.A(n_58367), .B(n_27986), .C(n_5743), .D(n_58000)
		, .Z(n_136471844));
	notech_ao4 i_153460273(.A(n_291863185), .B(n_236065889), .C(n_60167), .D
		(n_27159), .Z(n_136571845));
	notech_and4 i_154060267(.A(n_136571845), .B(n_136471844), .C(n_136271842
		), .D(n_136171841), .Z(n_136771847));
	notech_ao4 i_153160276(.A(n_57885), .B(\nbus_11358[4] ), .C(n_291463181)
		, .D(n_26614), .Z(n_136871848));
	notech_ao4 i_153060277(.A(n_291663183), .B(n_281566344), .C(n_57886), .D
		(\nbus_11307[4] ), .Z(n_136971849));
	notech_ao4 i_152860279(.A(n_54865), .B(n_29908), .C(n_54874), .D(n_28093
		), .Z(n_137171851));
	notech_ao4 i_152760280(.A(n_54894), .B(n_27430), .C(n_54883), .D(n_28597
		), .Z(n_137271852));
	notech_and4 i_153360274(.A(n_137271852), .B(n_137171851), .C(n_136971849
		), .D(n_136871848), .Z(n_137471854));
	notech_ao4 i_152460283(.A(n_111464643), .B(n_297966508), .C(n_111564644)
		, .D(n_59992), .Z(n_137571855));
	notech_ao4 i_152260284(.A(n_57999), .B(n_29678), .C(n_56512), .D(n_297766506
		), .Z(n_137671856));
	notech_ao4 i_152060286(.A(n_58367), .B(n_27983), .C(n_58000), .D(n_60024
		), .Z(n_137871858));
	notech_ao4 i_151860287(.A(n_236065889), .B(n_298066509), .C(n_60167), .D
		(n_27154), .Z(n_137971859));
	notech_and4 i_152660281(.A(n_137971859), .B(n_137871858), .C(n_137671856
		), .D(n_137571855), .Z(n_138171861));
	notech_ao4 i_151560290(.A(n_57885), .B(\nbus_11358[1] ), .C(n_297666505)
		, .D(n_26614), .Z(n_138271862));
	notech_ao4 i_151460291(.A(n_297866507), .B(n_281566344), .C(n_57886), .D
		(\nbus_11307[1] ), .Z(n_138371863));
	notech_ao4 i_151260293(.A(n_54865), .B(n_29906), .C(n_54874), .D(n_28090
		), .Z(n_138571865));
	notech_ao4 i_151060294(.A(n_54894), .B(n_27424), .C(n_54883), .D(n_28594
		), .Z(n_138671866));
	notech_and4 i_151760288(.A(n_138671866), .B(n_138571865), .C(n_138371863
		), .D(n_138271862), .Z(n_138871868));
	notech_or2 i_10458387(.A(n_58432), .B(n_60023), .Z(n_138971869));
	notech_and2 i_7158420(.A(n_26054), .B(n_57729), .Z(n_139071870));
	notech_and2 i_17358320(.A(n_145471934), .B(n_58714), .Z(n_139171871));
	notech_and2 i_17458319(.A(n_58717), .B(n_145571935), .Z(n_139271872));
	notech_or2 i_21858275(.A(n_151028787), .B(nbus_11295[2]), .Z(n_139371873
		));
	notech_or4 i_21358280(.A(n_62858), .B(n_56516), .C(n_62808), .D(n_57557)
		, .Z(n_140071880));
	notech_or4 i_54257952(.A(n_58802), .B(n_60940), .C(n_28136), .D(n_58482)
		, .Z(n_140971889));
	notech_nand2 i_54157953(.A(opd[10]), .B(n_58378), .Z(n_141271892));
	notech_or2 i_53657958(.A(n_3850), .B(n_57329), .Z(n_141771897));
	notech_nao3 i_55257942(.A(n_62798), .B(opc[11]), .C(n_58040), .Z(n_141871898
		));
	notech_or4 i_55157943(.A(n_62858), .B(n_128371763), .C(n_60940), .D(n_29596
		), .Z(n_142171901));
	notech_nand2 i_54857946(.A(n_58378), .B(opd[11]), .Z(n_142471904));
	notech_nand2 i_54557949(.A(opa[11]), .B(n_58055), .Z(n_142771907));
	notech_or2 i_9658395(.A(n_23514), .B(n_23510), .Z(n_142871908));
	notech_or2 i_13458359(.A(n_3844), .B(n_139071870), .Z(n_142971909));
	notech_nand2 i_29937(.A(n_58817), .B(n_58487), .Z(n_143071910));
	notech_or4 i_29947(.A(n_59387), .B(n_246891941), .C(n_29178), .D(n_26810
		), .Z(n_143471914));
	notech_or4 i_29721(.A(n_59387), .B(n_246891941), .C(n_32356), .D(n_29178
		), .Z(n_143571915));
	notech_ao4 i_189556655(.A(n_58391), .B(n_29733), .C(n_60329), .D(n_28091
		), .Z(n_143671916));
	notech_ao4 i_140757134(.A(n_29596), .B(n_128471764), .C(n_302491799), .D
		(n_57329), .Z(n_143771917));
	notech_ao4 i_140557136(.A(n_31456), .B(n_58482), .C(n_58054), .D(\nbus_11358[11] 
		), .Z(n_143971919));
	notech_and4 i_140957132(.A(n_143971919), .B(n_143771917), .C(n_142471904
		), .D(n_142771907), .Z(n_144171921));
	notech_ao4 i_140257139(.A(n_31476), .B(n_322373703), .C(n_30528), .D(n_26933
		), .Z(n_144271922));
	notech_and4 i_140457137(.A(n_187368889), .B(n_144271922), .C(n_141871898
		), .D(n_142171901), .Z(n_144571925));
	notech_ao4 i_139857143(.A(n_87532846), .B(n_58040), .C(n_187568890), .D(n_26933
		), .Z(n_144671926));
	notech_ao4 i_139757144(.A(\nbus_11307[10] ), .B(n_26679), .C(n_325273732
		), .D(n_29684), .Z(n_144871928));
	notech_ao4 i_139457147(.A(n_31411), .B(n_58482), .C(n_58054), .D(\nbus_11358[10] 
		), .Z(n_145071930));
	notech_and4 i_139657145(.A(n_187968894), .B(n_140971889), .C(n_145071930
		), .D(n_141271892), .Z(n_145371933));
	notech_mux2 i_110357425(.S(n_32323), .A(n_312147737), .B(n_344466973), .Z
		(n_145471934));
	notech_mux2 i_110157426(.S(n_32323), .A(n_312347735), .B(n_312447734), .Z
		(n_145571935));
	notech_ao4 i_109857429(.A(n_139271872), .B(n_142871908), .C(n_23514), .D
		(n_139171871), .Z(n_145671936));
	notech_ao4 i_109757430(.A(n_137375317), .B(n_152572005), .C(n_57892), .D
		(n_57557), .Z(n_145771937));
	notech_ao4 i_109557432(.A(n_137575319), .B(n_344366972), .C(n_137475318)
		, .D(n_152472004), .Z(n_145971939));
	notech_and4 i_110057427(.A(n_145971939), .B(n_145771937), .C(n_145671936
		), .D(n_140071880), .Z(n_146171941));
	notech_ao4 i_109257435(.A(n_58411), .B(n_27984), .C(n_57893), .D(\nbus_11358[2] 
		), .Z(n_146271942));
	notech_ao4 i_109157436(.A(n_54643), .B(n_28945), .C(n_315691667), .D(n_59991
		), .Z(n_146371943));
	notech_and4 i_109057437(.A(n_138971869), .B(n_143671916), .C(n_3849), .D
		(n_139371873), .Z(n_146671946));
	notech_or2 i_47155054(.A(n_26060), .B(n_57729), .Z(n_146871948));
	notech_nand2 i_34145(.A(n_26767), .B(n_27023), .Z(n_146971949));
	notech_or4 i_29528(.A(n_61175), .B(n_61165), .C(n_61154), .D(n_3852), .Z
		(n_147071950));
	notech_nand3 i_30289(.A(n_319191632), .B(n_319091633), .C(n_58078), .Z(n_147171951
		));
	notech_nao3 i_30070(.A(n_319191632), .B(n_319091633), .C(n_32356), .Z(n_147271952
		));
	notech_or2 i_30287(.A(n_151731932), .B(n_280073280), .Z(n_147371953));
	notech_nand2 i_31002(.A(n_58806), .B(n_58485), .Z(n_147471954));
	notech_nao3 i_34149(.A(n_319091633), .B(n_58078), .C(n_2479), .Z(n_147571955
		));
	notech_or4 i_33924(.A(n_2479), .B(n_56839), .C(n_27192), .D(n_56983), .Z
		(n_147671956));
	notech_or4 i_34146(.A(n_26062), .B(n_29652), .C(n_29658), .D(n_58163), .Z
		(n_147771957));
	notech_nand2 i_34154(.A(n_26767), .B(n_26698), .Z(n_147871958));
	notech_or2 i_57653375(.A(n_306824332), .B(n_3982), .Z(n_147971959));
	notech_or4 i_57553376(.A(n_56839), .B(n_56939), .C(n_26922), .D(n_28013)
		, .Z(n_148471964));
	notech_nand3 i_2921010(.A(n_150871988), .B(n_150771987), .C(n_147971959)
		, .Z(n_23902));
	notech_or2 i_126952699(.A(n_154831963), .B(n_3982), .Z(n_148771967));
	notech_or4 i_126852700(.A(n_246891941), .B(n_2479), .C(n_56689), .D(n_28013
		), .Z(n_149271972));
	notech_nand3 i_2921650(.A(n_151571995), .B(n_151471994), .C(n_148771967)
		, .Z(n_17948));
	notech_or2 i_130352667(.A(n_154831963), .B(n_3983), .Z(n_149571975));
	notech_or4 i_130252668(.A(n_246891941), .B(n_2479), .C(n_56689), .D(n_28011
		), .Z(n_150071980));
	notech_nand3 i_2721648(.A(n_152272002), .B(n_152172001), .C(n_149571975)
		, .Z(n_17936));
	notech_ao4 i_58153371(.A(n_307324337), .B(n_29662), .C(n_130528582), .D(n_58141
		), .Z(n_150371983));
	notech_ao4 i_58053372(.A(n_57864), .B(\nbus_11358[28] ), .C(n_314047718)
		, .D(\nbus_11365[28] ), .Z(n_150471984));
	notech_and4 i_58453368(.A(n_148471964), .B(n_150471984), .C(n_150371983)
		, .D(n_242259503), .Z(n_150771987));
	notech_ao4 i_58553367(.A(n_307124335), .B(n_172792106), .C(n_306624330),
		 .D(n_174492092), .Z(n_150871988));
	notech_ao4 i_127352695(.A(n_26929), .B(n_29662), .C(n_58147), .D(n_130528582
		), .Z(n_151071990));
	notech_ao4 i_127252696(.A(n_57875), .B(\nbus_11358[28] ), .C(n_57868), .D
		(\nbus_11365[28] ), .Z(n_151171991));
	notech_and4 i_127652692(.A(n_149271972), .B(n_151171991), .C(n_151071990
		), .D(n_242259503), .Z(n_151471994));
	notech_ao4 i_127752691(.A(n_58084), .B(n_172792106), .C(n_151931934), .D
		(n_174492092), .Z(n_151571995));
	notech_ao4 i_130752663(.A(n_29660), .B(n_26929), .C(n_133728614), .D(n_58147
		), .Z(n_151771997));
	notech_ao4 i_130652664(.A(n_57875), .B(\nbus_11358[26] ), .C(n_57868), .D
		(\nbus_11365[26] ), .Z(n_151871998));
	notech_and4 i_131052660(.A(n_150071980), .B(n_151871998), .C(n_151771997
		), .D(n_174892088), .Z(n_152172001));
	notech_ao4 i_131152659(.A(n_58084), .B(n_174292094), .C(n_151931934), .D
		(n_174992087), .Z(n_152272002));
	notech_nand2 i_70450658(.A(n_62798), .B(opc[2]), .Z(n_152472004));
	notech_nao3 i_71250657(.A(n_62798), .B(opa[2]), .C(n_62860), .Z(n_152572005
		));
	notech_nand3 i_77150656(.A(n_143671916), .B(n_181672296), .C(n_138971869
		), .Z(n_152672006));
	notech_mux2 i_5050616(.S(n_32335), .A(n_285027232), .B(n_284927231), .Z(n_152772007
		));
	notech_and2 i_5150615(.A(n_195572435), .B(n_58714), .Z(n_152872008));
	notech_and3 i_4850618(.A(n_162972109), .B(n_194072420), .C(n_58714), .Z(n_153172011
		));
	notech_and2 i_4950617(.A(n_58717), .B(n_193972419), .Z(n_153272012));
	notech_mux2 i_4650620(.S(n_32344), .A(n_285027232), .B(n_284927231), .Z(n_153372013
		));
	notech_mux2 i_4050626(.S(n_32322), .A(n_285027232), .B(n_284927231), .Z(n_153772017
		));
	notech_and2 i_4150625(.A(n_185672336), .B(n_58714), .Z(n_153872018));
	notech_mux2 i_3550631(.S(n_32331), .A(n_285027232), .B(n_284927231), .Z(n_154172021
		));
	notech_and2 i_3650630(.A(n_184872328), .B(n_58714), .Z(n_154272022));
	notech_nand2 i_3250634(.A(n_58717), .B(n_183872318), .Z(n_154672026));
	notech_ao4 i_3150635(.A(n_32309), .B(n_28126), .C(n_315891665), .D(n_29733
		), .Z(n_154972029));
	notech_or2 i_15850509(.A(n_150528782), .B(\nbus_11358[23] ), .Z(n_155872038
		));
	notech_or4 i_15550512(.A(n_61138), .B(n_60329), .C(n_19086), .D(n_28112)
		, .Z(n_156172041));
	notech_or2 i_15250515(.A(n_289127273), .B(n_150228779), .Z(n_156472044)
		);
	notech_or2 i_16950498(.A(n_150528782), .B(\nbus_11358[24] ), .Z(n_156972049
		));
	notech_or4 i_16650501(.A(n_61143), .B(n_60329), .C(n_19086), .D(n_28113)
		, .Z(n_157272052));
	notech_or2 i_16350504(.A(n_289027272), .B(n_150228779), .Z(n_157572055)
		);
	notech_nao3 i_20650461(.A(tsc[54]), .B(n_27855), .C(n_24989), .Z(n_157872058
		));
	notech_or2 i_20350464(.A(n_149228769), .B(n_29708), .Z(n_158172061));
	notech_or2 i_20050467(.A(n_289227274), .B(n_148728764), .Z(n_158472064)
		);
	notech_or4 i_21450453(.A(n_56839), .B(n_56939), .C(n_26927), .D(n_28008)
		, .Z(n_158872068));
	notech_or2 i_20950458(.A(n_148728764), .B(n_289127273), .Z(n_159372073)
		);
	notech_nao3 i_22450443(.A(tsc[56]), .B(n_27855), .C(n_24989), .Z(n_159672076
		));
	notech_or2 i_22150446(.A(n_149228769), .B(n_29769), .Z(n_159972079));
	notech_or2 i_21850449(.A(n_148728764), .B(n_289027272), .Z(n_160272082)
		);
	notech_or4 i_24450424(.A(n_26767), .B(n_3853), .C(n_28126), .D(n_60940),
		 .Z(n_160372083));
	notech_or4 i_24250425(.A(n_3854), .B(n_139071870), .C(n_32335), .D(n_57557
		), .Z(n_160672086));
	notech_or2 i_23950428(.A(n_59991), .B(n_147671956), .Z(n_160972089));
	notech_or4 i_23650431(.A(n_62842), .B(n_147871958), .C(n_60940), .D(n_57557
		), .Z(n_161272092));
	notech_nand2 i_29750371(.A(n_26644), .B(n_32334), .Z(n_162972109));
	notech_or2 i_31250356(.A(n_54894), .B(n_27469), .Z(n_163672116));
	notech_or2 i_30950359(.A(n_147028747), .B(\nbus_11358[22] ), .Z(n_163972119
		));
	notech_or4 i_30650362(.A(n_32555), .B(n_61145), .C(n_60340), .D(n_28111)
		, .Z(n_164272122));
	notech_or2 i_32550343(.A(n_54894), .B(n_27471), .Z(n_164972129));
	notech_or2 i_32250346(.A(n_147028747), .B(\nbus_11358[23] ), .Z(n_165272132
		));
	notech_or4 i_31950349(.A(n_32555), .B(n_61145), .C(n_60340), .D(n_28112)
		, .Z(n_165572135));
	notech_or2 i_33850330(.A(n_54894), .B(n_27473), .Z(n_166272142));
	notech_or2 i_33550333(.A(n_147028747), .B(\nbus_11358[24] ), .Z(n_166572145
		));
	notech_or4 i_33250336(.A(n_32555), .B(n_61145), .C(n_60329), .D(n_28113)
		, .Z(n_166872148));
	notech_or4 i_36150307(.A(n_26812), .B(n_58802), .C(n_28126), .D(n_60940)
		, .Z(n_167372153));
	notech_or4 i_36050308(.A(n_58184), .B(n_26852), .C(n_32344), .D(n_57557)
		, .Z(n_167672156));
	notech_or4 i_35750311(.A(n_246891941), .B(n_2479), .C(n_32356), .D(n_59991
		), .Z(n_167972159));
	notech_nao3 i_35250316(.A(n_58802), .B(n_26631), .C(n_26812), .Z(n_168072160
		));
	notech_ao4 i_35350315(.A(n_305291771), .B(n_189662168), .C(n_26647), .D(n_189672376
		), .Z(n_168172161));
	notech_or4 i_35450314(.A(n_62858), .B(n_284480345), .C(n_60938), .D(n_57557
		), .Z(n_168272162));
	notech_nand3 i_43050242(.A(n_54834), .B(n_7326), .C(\eflags[10] ), .Z(n_168772167
		));
	notech_or2 i_42750245(.A(n_144928726), .B(\nbus_11358[22] ), .Z(n_169072170
		));
	notech_nand3 i_42450248(.A(n_60167), .B(n_60246), .C(read_data[22]), .Z(n_169372173
		));
	notech_or2 i_42150251(.A(n_144428721), .B(n_289227274), .Z(n_169672176)
		);
	notech_nand3 i_44250230(.A(n_54834), .B(n_7328), .C(\eflags[10] ), .Z(n_169972179
		));
	notech_or2 i_43950233(.A(n_144928726), .B(\nbus_11358[23] ), .Z(n_170272182
		));
	notech_nand3 i_43650236(.A(n_60167), .B(n_60246), .C(read_data[23]), .Z(n_170572185
		));
	notech_or2 i_43350239(.A(n_144428721), .B(n_289127273), .Z(n_170872188)
		);
	notech_nand3 i_45450218(.A(n_54834), .B(n_7330), .C(\eflags[10] ), .Z(n_171172191
		));
	notech_or2 i_45150221(.A(n_144928726), .B(\nbus_11358[24] ), .Z(n_171472194
		));
	notech_nand3 i_44850224(.A(n_60167), .B(n_60246), .C(read_data[24]), .Z(n_171772197
		));
	notech_or2 i_44550227(.A(n_144428721), .B(n_289027272), .Z(n_172072200)
		);
	notech_or4 i_58650092(.A(n_58489), .B(n_58810), .C(n_28126), .D(n_60938)
		, .Z(n_172172201));
	notech_or4 i_58550093(.A(n_58133), .B(n_26906), .C(n_32322), .D(n_57557)
		, .Z(n_172472204));
	notech_or2 i_58250096(.A(n_304273522), .B(n_59991), .Z(n_172772207));
	notech_or4 i_57950099(.A(n_62854), .B(n_303873518), .C(n_60938), .D(n_57557
		), .Z(n_173072210));
	notech_ao3 i_72049966(.A(opc_10[2]), .B(n_62806), .C(n_57141), .Z(n_173372213
		));
	notech_ao4 i_71549971(.A(n_209069102), .B(n_26884), .C(n_26671), .D(n_26636
		), .Z(n_174072220));
	notech_ao3 i_76649920(.A(opc_10[2]), .B(n_62814), .C(n_57139), .Z(n_174572225
		));
	notech_and3 i_75949927(.A(n_58487), .B(n_58817), .C(n_154672026), .Z(n_175072230
		));
	notech_ao4 i_76049926(.A(n_305291771), .B(n_240762674), .C(n_26647), .D(n_183972319
		), .Z(n_175172231));
	notech_ao4 i_76149925(.A(n_281173291), .B(n_26828), .C(n_26671), .D(n_26632
		), .Z(n_175272232));
	notech_or2 i_83549852(.A(n_60023), .B(n_57470), .Z(n_175972239));
	notech_or4 i_83449853(.A(n_58087), .B(n_56529), .C(n_32338), .D(n_57557)
		, .Z(n_176272242));
	notech_nand3 i_83149856(.A(n_58632), .B(n_26808), .C(\opa_12[2] ), .Z(n_176572245
		));
	notech_or4 i_82849859(.A(n_62840), .B(n_56529), .C(n_62814), .D(n_57557)
		, .Z(n_176872248));
	notech_or4 i_90249787(.A(n_317391650), .B(n_317091653), .C(n_60023), .D(n_56401
		), .Z(n_177172251));
	notech_or2 i_89949790(.A(n_58406), .B(n_27984), .Z(n_177472254));
	notech_nand2 i_89649793(.A(sav_epc[2]), .B(n_61145), .Z(n_177772257));
	notech_nand2 i_30281(.A(n_58805), .B(n_26805), .Z(n_178472264));
	notech_nand2 i_33261(.A(n_58802), .B(n_58490), .Z(n_178572265));
	notech_ao4 i_194748769(.A(n_26721), .B(n_27860), .C(n_56548), .D(n_28562
		), .Z(n_180272282));
	notech_ao4 i_194648770(.A(n_26925), .B(n_28485), .C(n_27036), .D(n_28518
		), .Z(n_180372283));
	notech_ao4 i_194448772(.A(n_26928), .B(n_28453), .C(n_26651), .D(n_28160
		), .Z(n_180572285));
	notech_ao4 i_194348773(.A(n_56630), .B(n_28421), .C(n_56619), .D(n_28389
		), .Z(n_180672286));
	notech_and4 i_194948767(.A(n_180672286), .B(n_180572285), .C(n_180372283
		), .D(n_180272282), .Z(n_180872288));
	notech_ao4 i_194048776(.A(n_26920), .B(n_28357), .C(n_26933), .D(n_28324
		), .Z(n_180972289));
	notech_ao4 i_193948777(.A(n_26927), .B(n_28291), .C(n_56513), .D(n_29931
		), .Z(n_181072290));
	notech_and2 i_194148775(.A(n_181072290), .B(n_180972289), .Z(n_181172291
		));
	notech_ao4 i_193748779(.A(n_56921), .B(n_29930), .C(n_26969), .D(n_28259
		), .Z(n_181272292));
	notech_ao4 i_193648780(.A(n_26924), .B(n_28225), .C(n_26922), .D(n_28192
		), .Z(n_181372293));
	notech_ao4 i_191448800(.A(n_147071950), .B(n_57557), .C(n_58530), .D(\nbus_11358[2] 
		), .Z(n_181672296));
	notech_ao4 i_180948899(.A(n_285963126), .B(n_152572005), .C(n_317091653)
		, .D(n_154972029), .Z(n_181772297));
	notech_ao4 i_180848900(.A(n_122628503), .B(n_29540), .C(n_286063127), .D
		(n_152472004), .Z(n_181872298));
	notech_ao4 i_180648902(.A(n_317991644), .B(n_59991), .C(n_56533), .D(n_58316
		), .Z(n_182072300));
	notech_and4 i_181148897(.A(n_182072300), .B(n_181872298), .C(n_181772297
		), .D(n_177772257), .Z(n_182272302));
	notech_ao4 i_180348905(.A(n_309191732), .B(n_29929), .C(n_309291731), .D
		(n_28091), .Z(n_182372303));
	notech_ao4 i_180148907(.A(n_285663123), .B(n_57557), .C(n_58081), .D(\nbus_11358[2] 
		), .Z(n_182572305));
	notech_and4 i_180548903(.A(n_177172251), .B(n_182572305), .C(n_182372303
		), .D(n_177472254), .Z(n_182772307));
	notech_ao4 i_175348954(.A(n_152472004), .B(n_123971719), .C(n_152572005)
		, .D(n_124171721), .Z(n_182872308));
	notech_ao4 i_175148956(.A(n_57298), .B(n_28126), .C(n_59991), .D(n_124271722
		), .Z(n_183072310));
	notech_and4 i_175548952(.A(n_183072310), .B(n_182872308), .C(n_176572245
		), .D(n_176872248), .Z(n_183272312));
	notech_ao4 i_174848959(.A(\nbus_11358[2] ), .B(n_58044), .C(n_27984), .D
		(n_123771717), .Z(n_183372313));
	notech_and4 i_175048957(.A(n_175972239), .B(n_183372313), .C(n_26672), .D
		(n_176272242), .Z(n_183672316));
	notech_mux2 i_164249064(.S(n_58817), .A(n_152472004), .B(n_152572005), .Z
		(n_183772317));
	notech_mux2 i_164449062(.S(n_32332), .A(n_312347735), .B(n_312447734), .Z
		(n_183872318));
	notech_mux2 i_164349063(.S(n_32332), .A(n_26645), .B(n_26644), .Z(n_183972319
		));
	notech_ao4 i_163849068(.A(n_143471914), .B(n_27984), .C(n_59991), .D(n_143571915
		), .Z(n_184272322));
	notech_or4 i_164149065(.A(n_175172231), .B(n_175272232), .C(n_175072230)
		, .D(n_26633), .Z(n_184372323));
	notech_ao4 i_163649070(.A(n_123671716), .B(n_57557), .C(n_57573), .D(\nbus_11358[2] 
		), .Z(n_184472324));
	notech_mux2 i_160549101(.S(n_58805), .A(n_152472004), .B(n_152572005), .Z
		(n_184772327));
	notech_mux2 i_160649100(.S(n_32331), .A(n_312147737), .B(n_344466973), .Z
		(n_184872328));
	notech_ao4 i_160249104(.A(n_58486), .B(n_154272022), .C(n_178472264), .D
		(n_154172021), .Z(n_184972329));
	notech_ao4 i_160149105(.A(n_27984), .B(n_147171951), .C(n_59991), .D(n_147271952
		), .Z(n_185172331));
	notech_nao3 i_160449102(.A(n_184972329), .B(n_185172331), .C(n_174072220
		), .Z(n_185272332));
	notech_ao4 i_159949107(.A(n_147371953), .B(n_57557), .C(n_57154), .D(\nbus_11358[2] 
		), .Z(n_185372333));
	notech_mux2 i_149749207(.S(n_32322), .A(n_312147737), .B(n_344466973), .Z
		(n_185672336));
	notech_ao4 i_149449210(.A(n_58489), .B(n_153872018), .C(n_304073520), .D
		(n_153772017), .Z(n_185772337));
	notech_ao4 i_149249212(.A(n_26906), .B(n_58316), .C(n_303773517), .D(n_152472004
		), .Z(n_185972339));
	notech_and4 i_149649208(.A(n_185972339), .B(n_185772337), .C(n_172772207
		), .D(n_173072210), .Z(n_186172341));
	notech_ao4 i_148949215(.A(n_304173521), .B(\nbus_11358[2] ), .C(n_27984)
		, .D(n_303973519), .Z(n_186272342));
	notech_and4 i_149149213(.A(n_172172201), .B(n_186272342), .C(n_26672), .D
		(n_172472204), .Z(n_186572345));
	notech_ao4 i_138949310(.A(n_27329), .B(n_225565784), .C(n_221065739), .D
		(n_26803), .Z(n_186672346));
	notech_ao4 i_138749312(.A(n_27319), .B(n_28009), .C(n_60167), .D(n_27213
		), .Z(n_186872348));
	notech_and4 i_139149308(.A(n_186872348), .B(n_186672346), .C(n_171772197
		), .D(n_172072200), .Z(n_187072350));
	notech_ao4 i_138449315(.A(n_145128728), .B(n_60001), .C(n_145028727), .D
		(n_29769), .Z(n_187172351));
	notech_ao4 i_138249317(.A(n_54658), .B(n_29928), .C(n_144828725), .D(\nbus_11365[24] 
		), .Z(n_187372353));
	notech_and4 i_138649313(.A(n_187372353), .B(n_187172351), .C(n_171172191
		), .D(n_171472194), .Z(n_187572355));
	notech_ao4 i_137949320(.A(n_225665785), .B(n_27329), .C(n_222565754), .D
		(n_26803), .Z(n_187672356));
	notech_ao4 i_137749322(.A(n_27319), .B(n_28008), .C(n_60166), .D(n_27212
		), .Z(n_187872358));
	notech_and4 i_138149318(.A(n_187872358), .B(n_187672356), .C(n_170572185
		), .D(n_170872188), .Z(n_188072360));
	notech_ao4 i_137449325(.A(n_145128728), .B(n_60002), .C(n_145028727), .D
		(n_29765), .Z(n_188172361));
	notech_ao4 i_137249327(.A(n_54658), .B(n_29927), .C(n_144828725), .D(\nbus_11365[23] 
		), .Z(n_188372363));
	notech_and4 i_137649323(.A(n_188372363), .B(n_188172361), .C(n_169972179
		), .D(n_170272182), .Z(n_188572365));
	notech_ao4 i_136949330(.A(n_27329), .B(n_225765786), .C(n_224065769), .D
		(n_26803), .Z(n_188672366));
	notech_ao4 i_136749332(.A(n_27319), .B(n_28007), .C(n_60167), .D(n_27211
		), .Z(n_188872368));
	notech_and4 i_137149328(.A(n_188872368), .B(n_188672366), .C(n_169372173
		), .D(n_169672176), .Z(n_189072370));
	notech_ao4 i_136449335(.A(n_145128728), .B(n_60003), .C(n_145028727), .D
		(n_29708), .Z(n_189172371));
	notech_ao4 i_136249337(.A(n_54658), .B(n_29926), .C(n_144828725), .D(\nbus_11365[22] 
		), .Z(n_189372373));
	notech_and4 i_136649333(.A(n_189372373), .B(n_189172371), .C(n_168772167
		), .D(n_169072170), .Z(n_189572375));
	notech_mux2 i_132049379(.S(n_32344), .A(n_26645), .B(n_26644), .Z(n_189672376
		));
	notech_ao3 i_131849381(.A(n_168072160), .B(n_168272162), .C(n_168172161)
		, .Z(n_189872378));
	notech_ao4 i_131549384(.A(n_26852), .B(n_58316), .C(n_284680347), .D(n_152472004
		), .Z(n_189972379));
	notech_ao4 i_131249387(.A(n_57982), .B(\nbus_11358[2] ), .C(n_284580346)
		, .D(n_27984), .Z(n_190272382));
	notech_and4 i_131449385(.A(n_167372153), .B(n_190272382), .C(n_26672), .D
		(n_167672156), .Z(n_190572385));
	notech_ao4 i_129749402(.A(n_301791806), .B(n_225565784), .C(n_310491719)
		, .D(n_221065739), .Z(n_190672386));
	notech_ao4 i_129649403(.A(n_146928746), .B(\nbus_11365[24] ), .C(n_146428741
		), .D(n_289027272), .Z(n_190772387));
	notech_ao4 i_129449405(.A(n_310391720), .B(n_28009), .C(n_60167), .D(n_27182
		), .Z(n_190972389));
	notech_and4 i_129949400(.A(n_190972389), .B(n_190772387), .C(n_190672386
		), .D(n_166872148), .Z(n_191172391));
	notech_ao4 i_129149408(.A(n_147228749), .B(n_60001), .C(n_147128748), .D
		(n_29769), .Z(n_191272392));
	notech_ao4 i_128949410(.A(n_54883), .B(n_28617), .C(n_54865), .D(n_29918
		), .Z(n_191472394));
	notech_and4 i_129349406(.A(n_191472394), .B(n_191272392), .C(n_166272142
		), .D(n_166572145), .Z(n_191672396));
	notech_ao4 i_128649413(.A(n_301791806), .B(n_225665785), .C(n_310491719)
		, .D(n_222565754), .Z(n_191772397));
	notech_ao4 i_128549414(.A(n_146928746), .B(\nbus_11365[23] ), .C(n_146428741
		), .D(n_289127273), .Z(n_191872398));
	notech_ao4 i_128349416(.A(n_310391720), .B(n_28008), .C(n_60167), .D(n_27181
		), .Z(n_192072400));
	notech_and4 i_128849411(.A(n_192072400), .B(n_191872398), .C(n_191772397
		), .D(n_165572135), .Z(n_192272402));
	notech_ao4 i_128049419(.A(n_147228749), .B(n_60002), .C(n_147128748), .D
		(n_29765), .Z(n_192372403));
	notech_ao4 i_127849421(.A(n_54883), .B(n_28616), .C(n_54865), .D(n_29916
		), .Z(n_192572405));
	notech_and4 i_128249417(.A(n_192572405), .B(n_192372403), .C(n_164972129
		), .D(n_165272132), .Z(n_192772407));
	notech_ao4 i_127549424(.A(n_301791806), .B(n_225765786), .C(n_310491719)
		, .D(n_224065769), .Z(n_192872408));
	notech_ao4 i_127449425(.A(n_146928746), .B(\nbus_11365[22] ), .C(n_146428741
		), .D(n_289227274), .Z(n_192972409));
	notech_ao4 i_127249427(.A(n_310391720), .B(n_28007), .C(n_60167), .D(n_27178
		), .Z(n_193172411));
	notech_and4 i_127749422(.A(n_193172411), .B(n_192972409), .C(n_192872408
		), .D(n_164272122), .Z(n_193372413));
	notech_ao4 i_126949430(.A(n_147228749), .B(n_60003), .C(n_147128748), .D
		(n_29708), .Z(n_193472414));
	notech_ao4 i_126749432(.A(n_54883), .B(n_28615), .C(n_54865), .D(n_29914
		), .Z(n_193672416));
	notech_and4 i_127149428(.A(n_193672416), .B(n_193472414), .C(n_163672116
		), .D(n_163972119), .Z(n_193872418));
	notech_mux2 i_126649433(.S(n_32334), .A(n_312347735), .B(n_312447734), .Z
		(n_193972419));
	notech_ao4 i_126549434(.A(n_312147737), .B(n_32334), .C(n_153272012), .D
		(n_17107), .Z(n_194072420));
	notech_ao4 i_126149438(.A(n_281566344), .B(n_152572005), .C(n_26614), .D
		(n_153172011), .Z(n_194272422));
	notech_ao4 i_126049439(.A(n_56512), .B(n_58316), .C(n_111464643), .D(n_152472004
		), .Z(n_194372423));
	notech_ao4 i_125849441(.A(n_60158), .B(n_27156), .C(n_111564644), .D(n_59991
		), .Z(n_194572425));
	notech_ao4 i_125749442(.A(n_58367), .B(n_27984), .C(n_54874), .D(n_28091
		), .Z(n_194672426));
	notech_and4 i_126349436(.A(n_194672426), .B(n_194572425), .C(n_194372423
		), .D(n_194272422), .Z(n_194872428));
	notech_ao4 i_125449445(.A(n_57886), .B(n_57552), .C(n_57885), .D(\nbus_11358[2] 
		), .Z(n_194972429));
	notech_ao4 i_125349446(.A(n_54865), .B(n_29913), .C(n_236065889), .D(n_344366972
		), .Z(n_195072430));
	notech_ao4 i_125149448(.A(n_54894), .B(n_27426), .C(n_54883), .D(n_28595
		), .Z(n_195272432));
	notech_and4 i_125649443(.A(n_230865837), .B(n_195272432), .C(n_195072430
		), .D(n_194972429), .Z(n_195472434));
	notech_mux2 i_122049479(.S(n_32335), .A(n_312147737), .B(n_344466973), .Z
		(n_195572435));
	notech_ao4 i_121749482(.A(n_3853), .B(n_152872008), .C(n_146971949), .D(n_152772007
		), .Z(n_195672436));
	notech_ao4 i_121549484(.A(n_58163), .B(n_58316), .C(n_152472004), .D(n_147771957
		), .Z(n_195872438));
	notech_and4 i_121949480(.A(n_195872438), .B(n_195672436), .C(n_160972089
		), .D(n_161272092), .Z(n_196072440));
	notech_ao4 i_121249487(.A(\nbus_11358[2] ), .B(n_57980), .C(n_147571955)
		, .D(n_27984), .Z(n_196172441));
	notech_ao3 i_121149488(.A(n_160372083), .B(n_125828535), .C(n_152672006)
		, .Z(n_196472444));
	notech_ao4 i_119949500(.A(n_221065739), .B(n_310891715), .C(n_225565784)
		, .D(n_310791716), .Z(n_196672446));
	notech_ao4 i_119749502(.A(n_149328770), .B(\nbus_11365[24] ), .C(n_149428771
		), .D(\nbus_11358[24] ), .Z(n_196872448));
	notech_and4 i_120149498(.A(n_196872448), .B(n_196672446), .C(n_159972079
		), .D(n_160272082), .Z(n_197072450));
	notech_ao4 i_119449505(.A(n_310691717), .B(n_28009), .C(n_149128768), .D
		(n_60001), .Z(n_197172451));
	notech_ao4 i_119349506(.A(n_3867), .B(n_27025), .C(n_28113), .D(n_60340)
		, .Z(n_197372453));
	notech_ao4 i_119049509(.A(n_222565754), .B(n_310891715), .C(n_225665785)
		, .D(n_310791716), .Z(n_197572455));
	notech_ao4 i_118949510(.A(n_149328770), .B(\nbus_11365[23] ), .C(n_149428771
		), .D(\nbus_11358[23] ), .Z(n_197772457));
	notech_and3 i_119249507(.A(n_197572455), .B(n_197772457), .C(n_159372073
		), .Z(n_197872458));
	notech_ao4 i_118449513(.A(n_149128768), .B(n_60002), .C(n_149228769), .D
		(n_29765), .Z(n_197972459));
	notech_ao4 i_118349514(.A(n_28112), .B(n_60329), .C(n_54643), .D(n_28978
		), .Z(n_198172461));
	notech_ao4 i_118049517(.A(n_224065769), .B(n_310891715), .C(n_225765786)
		, .D(n_310791716), .Z(n_198372463));
	notech_ao4 i_117849519(.A(n_149328770), .B(\nbus_11365[22] ), .C(n_149428771
		), .D(\nbus_11358[22] ), .Z(n_198572465));
	notech_and4 i_118249515(.A(n_198572465), .B(n_198372463), .C(n_158172061
		), .D(n_158472064), .Z(n_198772467));
	notech_ao4 i_117549522(.A(n_310691717), .B(n_28007), .C(n_149128768), .D
		(n_60003), .Z(n_198872468));
	notech_ao4 i_117449523(.A(n_28111), .B(n_60329), .C(n_3867), .D(n_27025)
		, .Z(n_199072470));
	notech_ao4 i_115049547(.A(n_225565784), .B(n_308791736), .C(n_221065739)
		, .D(n_307891745), .Z(n_199272472));
	notech_ao4 i_114849549(.A(n_308591738), .B(n_28009), .C(n_60158), .D(n_27147
		), .Z(n_199472474));
	notech_and4 i_115249545(.A(n_199472474), .B(n_199272472), .C(n_157272052
		), .D(n_157572055), .Z(n_199672476));
	notech_ao4 i_114549552(.A(n_60001), .B(n_150728784), .C(n_150628783), .D
		(n_29769), .Z(n_199772477));
	notech_ao4 i_114449553(.A(n_26648), .B(n_29911), .C(n_150428781), .D(\nbus_11365[24] 
		), .Z(n_199972479));
	notech_ao4 i_114049556(.A(n_225665785), .B(n_308791736), .C(n_222565754)
		, .D(n_307891745), .Z(n_200172481));
	notech_ao4 i_113849558(.A(n_308591738), .B(n_28008), .C(n_60158), .D(n_27146
		), .Z(n_200372483));
	notech_and4 i_114349554(.A(n_200372483), .B(n_200172481), .C(n_156172041
		), .D(n_156472044), .Z(n_200572485));
	notech_ao4 i_113549561(.A(n_60002), .B(n_150728784), .C(n_150628783), .D
		(n_29765), .Z(n_200672486));
	notech_ao4 i_113449562(.A(n_26648), .B(n_29910), .C(n_150428781), .D(\nbus_11365[23] 
		), .Z(n_200872488));
	notech_or4 i_11347586(.A(n_317591648), .B(n_27104), .C(n_316491659), .D(\nbus_11358[17] 
		), .Z(n_201772497));
	notech_nand2 i_11047589(.A(n_151328790), .B(\regs_13_14[17] ), .Z(n_202072500
		));
	notech_or4 i_10747592(.A(n_316491659), .B(n_26942), .C(nbus_11295[17]), 
		.D(n_60940), .Z(n_202372503));
	notech_or4 i_13647564(.A(n_317591648), .B(n_27104), .C(n_316491659), .D(\nbus_11358[19] 
		), .Z(n_202872508));
	notech_nand2 i_13347567(.A(\regs_13_14[19] ), .B(n_151328790), .Z(n_203172511
		));
	notech_or4 i_13047570(.A(n_316491659), .B(n_26942), .C(nbus_11295[19]), 
		.D(n_60940), .Z(n_203472514));
	notech_ao3 i_14847552(.A(tsc[20]), .B(n_27855), .C(n_24989), .Z(n_203572515
		));
	notech_or2 i_14747553(.A(n_151028787), .B(nbus_11295[20]), .Z(n_203872518
		));
	notech_or4 i_14447556(.A(n_56839), .B(n_56935), .C(n_26925), .D(n_28005)
		, .Z(n_204172521));
	notech_or2 i_14147559(.A(n_151128788), .B(n_313347725), .Z(n_204472524)
		);
	notech_nao3 i_17747523(.A(\regs_1_0[17] ), .B(n_19086), .C(n_32270), .Z(n_204772527
		));
	notech_or2 i_17447526(.A(n_60008), .B(n_150728784), .Z(n_205072530));
	notech_or4 i_17147529(.A(n_56689), .B(n_26721), .C(n_61145), .D(n_28002)
		, .Z(n_205372533));
	notech_nao3 i_16847532(.A(opc_10[17]), .B(n_62786), .C(n_308791736), .Z(n_205672536
		));
	notech_nao3 i_20147499(.A(\regs_1_0[19] ), .B(n_19086), .C(n_32270), .Z(n_205972539
		));
	notech_or2 i_19847502(.A(n_150728784), .B(n_60006), .Z(n_206272542));
	notech_or4 i_19547505(.A(n_56689), .B(n_26721), .C(n_61145), .D(n_28004)
		, .Z(n_206572545));
	notech_nao3 i_19247508(.A(opc_10[19]), .B(n_62808), .C(n_308791736), .Z(n_206872548
		));
	notech_or2 i_21047490(.A(n_150528782), .B(\nbus_11358[20] ), .Z(n_207372553
		));
	notech_or4 i_20747493(.A(n_61145), .B(n_60329), .C(n_19086), .D(n_28109)
		, .Z(n_207672556));
	notech_or2 i_20447496(.A(n_150228779), .B(n_313347725), .Z(n_207972559)
		);
	notech_or2 i_23147469(.A(n_149428771), .B(\nbus_11358[17] ), .Z(n_208372563
		));
	notech_or4 i_22847472(.A(n_56839), .B(n_56935), .C(n_26927), .D(n_28002)
		, .Z(n_208672566));
	notech_or4 i_22547475(.A(n_311891705), .B(n_26939), .C(n_28143), .D(n_60940
		), .Z(n_208972569));
	notech_or2 i_24147459(.A(n_149428771), .B(\nbus_11358[18] ), .Z(n_209372573
		));
	notech_or4 i_23847462(.A(n_56839), .B(n_56944), .C(n_26927), .D(n_28003)
		, .Z(n_209672576));
	notech_or4 i_23547465(.A(n_311891705), .B(n_26939), .C(n_60949), .D(n_28144
		), .Z(n_209972579));
	notech_or2 i_25147449(.A(n_149428771), .B(\nbus_11358[19] ), .Z(n_210372583
		));
	notech_or4 i_24847452(.A(n_56839), .B(n_56935), .C(n_56527), .D(n_28004)
		, .Z(n_210672586));
	notech_or4 i_24547455(.A(n_311891705), .B(n_26939), .C(n_28145), .D(n_60949
		), .Z(n_210972589));
	notech_or2 i_26047440(.A(n_149328770), .B(\nbus_11365[20] ), .Z(n_211372593
		));
	notech_or2 i_25547445(.A(n_148728764), .B(n_313347725), .Z(n_211872598)
		);
	notech_or4 i_27947421(.A(n_3854), .B(n_3845), .C(n_27089), .D(\nbus_11358[17] 
		), .Z(n_212172601));
	notech_or4 i_27647424(.A(n_56839), .B(n_56935), .C(n_26928), .D(n_28002)
		, .Z(n_212472604));
	notech_or4 i_27347427(.A(n_3845), .B(n_26767), .C(nbus_11295[17]), .D(n_60947
		), .Z(n_212772607));
	notech_or4 i_30147403(.A(n_3854), .B(n_3845), .C(n_27089), .D(\nbus_11358[19] 
		), .Z(n_213072610));
	notech_or4 i_29847406(.A(n_56839), .B(n_56935), .C(n_26928), .D(n_28004)
		, .Z(n_213372613));
	notech_or4 i_29547409(.A(n_3845), .B(n_26767), .C(nbus_11295[19]), .D(n_60949
		), .Z(n_213672616));
	notech_nor2 i_31347395(.A(n_3878), .B(\nbus_11365[20] ), .Z(n_213772617)
		);
	notech_or2 i_30447400(.A(n_3837), .B(n_313347725), .Z(n_214472624));
	notech_or4 i_41147298(.A(n_58184), .B(n_58498), .C(n_26664), .D(\nbus_11358[17] 
		), .Z(n_214572625));
	notech_or2 i_41047299(.A(n_58147), .B(n_60008), .Z(n_214872628));
	notech_or4 i_40547304(.A(n_58802), .B(n_58498), .C(nbus_11295[17]), .D(n_60949
		), .Z(n_215372633));
	notech_or4 i_42147289(.A(n_58184), .B(n_58498), .C(n_26664), .D(\nbus_11358[18] 
		), .Z(n_215472634));
	notech_or2 i_42047290(.A(n_58147), .B(n_3864), .Z(n_215772637));
	notech_or4 i_41447295(.A(n_58802), .B(n_58498), .C(n_60949), .D(nbus_11295
		[18]), .Z(n_216272642));
	notech_or4 i_43047280(.A(n_58184), .B(n_58498), .C(n_26664), .D(\nbus_11358[19] 
		), .Z(n_216372643));
	notech_or2 i_42947281(.A(n_58147), .B(n_60006), .Z(n_216672646));
	notech_or4 i_42447286(.A(n_58802), .B(n_58498), .C(nbus_11295[19]), .D(n_60947
		), .Z(n_217172651));
	notech_nor2 i_43847272(.A(n_57868), .B(\nbus_11365[20] ), .Z(n_217272652
		));
	notech_or2 i_43347277(.A(n_154831963), .B(n_313347725), .Z(n_217972659)
		);
	notech_nand3 i_46947242(.A(n_54834), .B(n_7316), .C(n_56172), .Z(n_218272662
		));
	notech_or4 i_46647245(.A(n_56689), .B(n_56548), .C(n_61145), .D(n_28002)
		, .Z(n_218572665));
	notech_or2 i_46347248(.A(n_145028727), .B(n_29772), .Z(n_218872668));
	notech_nand3 i_48247229(.A(n_54834), .B(n_7318), .C(n_56172), .Z(n_219572675
		));
	notech_or4 i_47947232(.A(n_56689), .B(n_56548), .C(n_61145), .D(n_28003)
		, .Z(n_219872678));
	notech_or2 i_47647235(.A(n_145028727), .B(n_29711), .Z(n_220172681));
	notech_nand3 i_49547216(.A(n_54834), .B(n_7320), .C(n_56172), .Z(n_220872688
		));
	notech_or4 i_49247219(.A(n_56689), .B(n_56548), .C(n_61145), .D(n_28004)
		, .Z(n_221172691));
	notech_or2 i_48947222(.A(n_145028727), .B(n_29773), .Z(n_221472694));
	notech_nand3 i_50747204(.A(n_54834), .B(n_7322), .C(n_56172), .Z(n_222172701
		));
	notech_or4 i_50447207(.A(n_56689), .B(n_56542), .C(n_61145), .D(n_28005)
		, .Z(n_222472704));
	notech_or2 i_50147210(.A(n_145028727), .B(n_29775), .Z(n_222772707));
	notech_nand3 i_49847213(.A(opc[20]), .B(n_62806), .C(n_27340), .Z(n_223072710
		));
	notech_or2 i_64947070(.A(n_138168398), .B(\nbus_11365[17] ), .Z(n_223172711
		));
	notech_or4 i_64847071(.A(n_58133), .B(n_58497), .C(n_56428), .D(\nbus_11358[17] 
		), .Z(n_223472714));
	notech_nao3 i_64347076(.A(opc_10[17]), .B(n_62788), .C(n_319937994), .Z(n_223972719
		));
	notech_or2 i_66747052(.A(n_138168398), .B(\nbus_11365[19] ), .Z(n_224072720
		));
	notech_or4 i_66647053(.A(n_58133), .B(n_58497), .C(n_56428), .D(\nbus_11358[19] 
		), .Z(n_224372723));
	notech_nao3 i_66147058(.A(opc_10[19]), .B(n_62806), .C(n_319937994), .Z(n_224872728
		));
	notech_nor2 i_67947044(.A(n_57869), .B(\nbus_11365[20] ), .Z(n_224972729
		));
	notech_or2 i_67047049(.A(n_321538010), .B(n_313347725), .Z(n_225672736)
		);
	notech_nor2 i_69947024(.A(n_154331958), .B(nbus_11295[17]), .Z(n_225772737
		));
	notech_or4 i_69847025(.A(n_56839), .B(n_56944), .C(n_56921), .D(n_28002)
		, .Z(n_226072740));
	notech_or2 i_69547028(.A(n_58143), .B(n_60008), .Z(n_226372743));
	notech_or2 i_69247031(.A(n_286869880), .B(\nbus_11365[17] ), .Z(n_226672746
		));
	notech_or4 i_80146923(.A(n_56839), .B(n_56944), .C(n_26922), .D(n_28002)
		, .Z(n_226772747));
	notech_or4 i_80046924(.A(n_58099), .B(n_58494), .C(n_56437), .D(\nbus_11358[17] 
		), .Z(n_227072750));
	notech_or2 i_79546929(.A(n_313647722), .B(n_306824332), .Z(n_227572755)
		);
	notech_or4 i_81946905(.A(n_56839), .B(n_56944), .C(n_26922), .D(n_28004)
		, .Z(n_227672756));
	notech_or4 i_81846906(.A(n_58099), .B(n_58494), .C(n_56437), .D(\nbus_11358[19] 
		), .Z(n_227972759));
	notech_or2 i_81346911(.A(n_306824332), .B(n_313447724), .Z(n_228472764)
		);
	notech_or4 i_82746897(.A(n_56839), .B(n_56944), .C(n_26922), .D(n_28005)
		, .Z(n_228572765));
	notech_or4 i_82246902(.A(n_58805), .B(n_58494), .C(nbus_11295[20]), .D(n_60947
		), .Z(n_229272772));
	notech_nor2 i_85146873(.A(n_57861), .B(\nbus_11365[18] ), .Z(n_229372773
		));
	notech_or2 i_84646878(.A(n_287827260), .B(n_3861), .Z(n_230072780));
	notech_nor2 i_85946865(.A(n_57861), .B(\nbus_11365[19] ), .Z(n_230172781
		));
	notech_or2 i_85446870(.A(n_287827260), .B(n_313447724), .Z(n_230872788)
		);
	notech_nor2 i_86746857(.A(n_57861), .B(\nbus_11365[20] ), .Z(n_230972789
		));
	notech_or2 i_86246862(.A(n_287827260), .B(n_313347725), .Z(n_231672796)
		);
	notech_or4 i_92146811(.A(n_56839), .B(n_56944), .C(n_26969), .D(n_28002)
		, .Z(n_231772797));
	notech_or2 i_92046812(.A(n_58138), .B(n_60008), .Z(n_232072800));
	notech_nao3 i_91546817(.A(opc_10[17]), .B(n_62806), .C(n_58007), .Z(n_232572805
		));
	notech_or4 i_93446798(.A(n_56837), .B(n_56935), .C(n_26969), .D(n_28003)
		, .Z(n_232672806));
	notech_or2 i_93346799(.A(n_58138), .B(n_3864), .Z(n_232972809));
	notech_nao3 i_92846804(.A(n_62798), .B(opc_10[18]), .C(n_58007), .Z(n_233472814
		));
	notech_or4 i_94746785(.A(n_56837), .B(n_56935), .C(n_26969), .D(n_28004)
		, .Z(n_233572815));
	notech_or2 i_94646786(.A(n_58138), .B(n_60006), .Z(n_233872818));
	notech_nao3 i_94146791(.A(opc_10[19]), .B(n_62806), .C(n_58007), .Z(n_234372823
		));
	notech_or4 i_96046772(.A(n_56837), .B(n_56935), .C(n_26969), .D(n_28005)
		, .Z(n_234472824));
	notech_or2 i_95946773(.A(n_58138), .B(n_60005), .Z(n_234772827));
	notech_nao3 i_95446778(.A(opc_10[20]), .B(n_62788), .C(n_58007), .Z(n_235272832
		));
	notech_or2 i_103346700(.A(n_308991734), .B(\nbus_11365[18] ), .Z(n_237172851
		));
	notech_or2 i_103046703(.A(n_122428501), .B(n_28144), .Z(n_237472854));
	notech_nao3 i_102746706(.A(n_19065), .B(read_data[18]), .C(n_59100), .Z(n_237772857
		));
	notech_nand2 i_102446709(.A(add_len_pc[18]), .B(n_26766), .Z(n_238072860
		));
	notech_nand2 i_5147648(.A(n_26916), .B(n_26811), .Z(n_241372893));
	notech_or2 i_4847651(.A(n_58494), .B(n_57926), .Z(n_241472894));
	notech_nand2 i_41747693(.A(opc[20]), .B(n_62788), .Z(n_241572895));
	notech_ao4 i_211045673(.A(n_56542), .B(n_28581), .C(n_27036), .D(n_28541
		), .Z(n_241672896));
	notech_ao4 i_210945674(.A(n_28504), .B(n_26925), .C(n_26721), .D(n_27881
		), .Z(n_241772897));
	notech_ao4 i_210745676(.A(n_26928), .B(n_28471), .C(n_26651), .D(n_28178
		), .Z(n_241972899));
	notech_ao4 i_210645677(.A(n_56632), .B(n_28439), .C(n_56614), .D(n_28407
		), .Z(n_242072900));
	notech_and4 i_211245671(.A(n_242072900), .B(n_241972899), .C(n_241772897
		), .D(n_241672896), .Z(n_242272902));
	notech_ao4 i_210345680(.A(n_26920), .B(n_28375), .C(n_26933), .D(n_28343
		), .Z(n_242372903));
	notech_ao4 i_210245681(.A(n_56527), .B(n_28310), .C(n_56513), .D(n_29944
		), .Z(n_242472904));
	notech_and2 i_210445679(.A(n_242472904), .B(n_242372903), .Z(n_242572905
		));
	notech_ao4 i_210045683(.A(n_56921), .B(n_29943), .C(n_26969), .D(n_28277
		), .Z(n_242672906));
	notech_ao4 i_209945684(.A(n_26924), .B(n_28245), .C(n_26922), .D(n_28210
		), .Z(n_242772907));
	notech_nand2 i_28947701(.A(opc[19]), .B(n_62806), .Z(n_243072910));
	notech_ao4 i_208645697(.A(n_56542), .B(n_28580), .C(n_56566), .D(n_28540
		), .Z(n_243172911));
	notech_ao4 i_208545698(.A(n_28503), .B(n_26925), .C(n_26721), .D(n_27878
		), .Z(n_243272912));
	notech_ao4 i_208345700(.A(n_26928), .B(n_28470), .C(n_26651), .D(n_28177
		), .Z(n_243472914));
	notech_ao4 i_208245701(.A(n_56632), .B(n_28438), .C(n_56614), .D(n_28406
		), .Z(n_243572915));
	notech_and4 i_208845695(.A(n_243572915), .B(n_243472914), .C(n_243272912
		), .D(n_243172911), .Z(n_243772917));
	notech_ao4 i_207945704(.A(n_26920), .B(n_28374), .C(n_26933), .D(n_28342
		), .Z(n_243872918));
	notech_ao4 i_207845705(.A(n_56527), .B(n_28309), .C(n_56513), .D(n_29942
		), .Z(n_243972919));
	notech_and2 i_208045703(.A(n_243972919), .B(n_243872918), .Z(n_244072920
		));
	notech_ao4 i_207645707(.A(n_56921), .B(n_29941), .C(n_26969), .D(n_28276
		), .Z(n_244172921));
	notech_ao4 i_207545708(.A(n_26924), .B(n_28244), .C(n_26922), .D(n_28209
		), .Z(n_244272922));
	notech_ao4 i_204845735(.A(n_124328520), .B(n_3861), .C(n_309391730), .D(n_95222216
		), .Z(n_244572925));
	notech_ao4 i_204645737(.A(n_121628493), .B(n_28003), .C(n_60158), .D(n_27260
		), .Z(n_244772927));
	notech_and4 i_205045733(.A(n_244772927), .B(n_244572925), .C(n_238072860
		), .D(n_237772857), .Z(n_244972929));
	notech_ao4 i_204345740(.A(n_26765), .B(n_29711), .C(n_309191732), .D(n_29940
		), .Z(n_245072930));
	notech_ao4 i_204145742(.A(n_309091733), .B(\nbus_11358[18] ), .C(n_122528502
		), .D(n_3864), .Z(n_245272932));
	notech_and4 i_204545738(.A(n_245272932), .B(n_245072930), .C(n_237172851
		), .D(n_237472854), .Z(n_245472934));
	notech_nand2 i_29347698(.A(opc[17]), .B(n_62788), .Z(n_245572935));
	notech_ao4 i_203845745(.A(n_56547), .B(n_28578), .C(n_56566), .D(n_28538
		), .Z(n_245672936));
	notech_ao4 i_203745746(.A(n_28500), .B(n_26925), .C(n_26721), .D(n_27875
		), .Z(n_245772937));
	notech_ao4 i_203545748(.A(n_26928), .B(n_28468), .C(n_26651), .D(n_28175
		), .Z(n_245972939));
	notech_ao4 i_203445749(.A(n_56632), .B(n_28436), .C(n_56614), .D(n_28404
		), .Z(n_246072940));
	notech_and4 i_204045743(.A(n_246072940), .B(n_245972939), .C(n_245772937
		), .D(n_245672936), .Z(n_246272942));
	notech_ao4 i_203145752(.A(n_26920), .B(n_28372), .C(n_26933), .D(n_28340
		), .Z(n_246372943));
	notech_ao4 i_203045753(.A(n_56527), .B(n_28307), .C(n_56513), .D(n_29939
		), .Z(n_246472944));
	notech_and2 i_203245751(.A(n_246472944), .B(n_246372943), .Z(n_246572945
		));
	notech_ao4 i_202845755(.A(n_56921), .B(n_29938), .C(n_26969), .D(n_28274
		), .Z(n_246672946));
	notech_ao4 i_202745756(.A(n_26924), .B(n_28242), .C(n_26922), .D(n_28207
		), .Z(n_246772947));
	notech_nand2 i_2047702(.A(opc_10[20]), .B(n_62806), .Z(n_247072950));
	notech_ao4 i_198645796(.A(n_58008), .B(n_241572895), .C(n_305624320), .D
		(n_313347725), .Z(n_247172951));
	notech_ao4 i_198545797(.A(n_57726), .B(n_28146), .C(n_26937), .D(n_29775
		), .Z(n_247372953));
	notech_ao4 i_198245800(.A(n_57867), .B(\nbus_11365[20] ), .C(n_57865), .D
		(\nbus_11358[20] ), .Z(n_247572955));
	notech_and4 i_198445798(.A(n_234472824), .B(n_247572955), .C(n_26623), .D
		(n_234772827), .Z(n_247872958));
	notech_nand2 i_1947703(.A(opc_10[19]), .B(n_62788), .Z(n_247972959));
	notech_ao4 i_197345807(.A(n_58008), .B(n_243072910), .C(n_305624320), .D
		(n_313447724), .Z(n_248072960));
	notech_ao4 i_197245808(.A(n_57726), .B(n_28145), .C(n_26937), .D(n_29773
		), .Z(n_248272962));
	notech_ao4 i_196945811(.A(n_57867), .B(\nbus_11365[19] ), .C(n_57865), .D
		(\nbus_11358[19] ), .Z(n_248472964));
	notech_and4 i_197145809(.A(n_233572815), .B(n_248472964), .C(n_26622), .D
		(n_233872818), .Z(n_248772967));
	notech_ao4 i_196245818(.A(n_58008), .B(n_95222216), .C(n_3861), .D(n_305624320
		), .Z(n_248872968));
	notech_ao4 i_196145819(.A(n_57726), .B(n_28144), .C(n_26937), .D(n_29711
		), .Z(n_249072970));
	notech_ao4 i_195845822(.A(n_57867), .B(\nbus_11365[18] ), .C(n_57865), .D
		(\nbus_11358[18] ), .Z(n_249272972));
	notech_and4 i_196045820(.A(n_232672806), .B(n_249272972), .C(n_26621), .D
		(n_232972809), .Z(n_249572975));
	notech_nand2 i_1747705(.A(opc_10[17]), .B(n_62822), .Z(n_249672976));
	notech_ao4 i_195145829(.A(n_58008), .B(n_245572935), .C(n_313647722), .D
		(n_305624320), .Z(n_249772977));
	notech_ao4 i_195045830(.A(n_57726), .B(n_28143), .C(n_26937), .D(n_29772
		), .Z(n_249972979));
	notech_ao4 i_194745833(.A(n_57867), .B(\nbus_11365[17] ), .C(n_57865), .D
		(\nbus_11358[17] ), .Z(n_250172981));
	notech_and4 i_194945831(.A(n_231772797), .B(n_250172981), .C(n_26624), .D
		(n_232072800), .Z(n_250472984));
	notech_ao4 i_185445910(.A(n_286827250), .B(n_247072950), .C(n_286927251)
		, .D(n_241572895), .Z(n_250572985));
	notech_ao4 i_185345911(.A(n_26615), .B(n_29775), .C(n_58424), .D(n_28005
		), .Z(n_250772987));
	notech_nand3 i_185645908(.A(n_250572985), .B(n_250772987), .C(n_231672796
		), .Z(n_250872988));
	notech_ao4 i_185145913(.A(n_57863), .B(\nbus_11358[20] ), .C(n_58139), .D
		(n_60005), .Z(n_250972989));
	notech_ao4 i_184745917(.A(n_286827250), .B(n_247972959), .C(n_286927251)
		, .D(n_243072910), .Z(n_251272992));
	notech_ao4 i_184645918(.A(n_26615), .B(n_29773), .C(n_58424), .D(n_28004
		), .Z(n_251472994));
	notech_nand3 i_184945915(.A(n_251272992), .B(n_251472994), .C(n_230872788
		), .Z(n_251572995));
	notech_ao4 i_184445920(.A(n_57863), .B(\nbus_11358[19] ), .C(n_58139), .D
		(n_60006), .Z(n_251672996));
	notech_ao4 i_184045924(.A(n_286827250), .B(n_77522039), .C(n_286927251),
		 .D(n_95222216), .Z(n_251972999));
	notech_ao4 i_183945925(.A(n_26615), .B(n_29711), .C(n_58424), .D(n_28003
		), .Z(n_252173001));
	notech_nand3 i_184245922(.A(n_251972999), .B(n_252173001), .C(n_230072780
		), .Z(n_252273002));
	notech_ao4 i_183745927(.A(n_57863), .B(\nbus_11358[18] ), .C(n_58139), .D
		(n_3864), .Z(n_252373003));
	notech_ao4 i_181845945(.A(n_306824332), .B(n_313347725), .C(n_247072950)
		, .D(n_306624330), .Z(n_252673006));
	notech_ao4 i_181745946(.A(n_314047718), .B(\nbus_11365[20] ), .C(n_29775
		), .D(n_307324337), .Z(n_252873008));
	notech_ao4 i_181545948(.A(\nbus_11358[20] ), .B(n_57864), .C(n_58141), .D
		(n_60005), .Z(n_253073010));
	notech_and3 i_181645947(.A(n_228572765), .B(n_253073010), .C(n_26623), .Z
		(n_253273012));
	notech_ao4 i_181145952(.A(n_247972959), .B(n_306624330), .C(\nbus_11365[19] 
		), .D(n_241472894), .Z(n_253373013));
	notech_ao4 i_181045953(.A(n_29773), .B(n_307324337), .C(n_243072910), .D
		(n_307124335), .Z(n_253573015));
	notech_or4 i_30847696(.A(n_60970), .B(n_60959), .C(n_62860), .D(\nbus_11365[19] 
		), .Z(n_253773017));
	notech_ao4 i_180745956(.A(n_58141), .B(n_60006), .C(n_58494), .D(n_253773017
		), .Z(n_253873018));
	notech_and4 i_180945954(.A(n_227672756), .B(n_253873018), .C(n_26622), .D
		(n_227972759), .Z(n_254173021));
	notech_ao4 i_179445968(.A(n_249672976), .B(n_306624330), .C(n_241472894)
		, .D(\nbus_11365[17] ), .Z(n_254273022));
	notech_ao4 i_179145969(.A(n_29772), .B(n_307324337), .C(n_245572935), .D
		(n_307124335), .Z(n_254473024));
	notech_or4 i_31147694(.A(n_60970), .B(n_60959), .C(n_62860), .D(\nbus_11365[17] 
		), .Z(n_254673026));
	notech_ao4 i_178845972(.A(n_58141), .B(n_60008), .C(n_58494), .D(n_254673026
		), .Z(n_254773027));
	notech_and4 i_179045970(.A(n_226772747), .B(n_254773027), .C(n_26624), .D
		(n_227072750), .Z(n_255073030));
	notech_ao4 i_170446056(.A(n_306124325), .B(n_249672976), .C(n_313647722)
		, .D(n_305924323), .Z(n_255173031));
	notech_ao4 i_170146058(.A(n_58085), .B(n_245572935), .C(n_58493), .D(n_254673026
		), .Z(n_255373033));
	notech_and4 i_170646054(.A(n_255373033), .B(n_255173031), .C(n_226372743
		), .D(n_226672746), .Z(n_255573035));
	notech_ao4 i_169746061(.A(n_57877), .B(\nbus_11358[17] ), .C(n_26902), .D
		(n_29772), .Z(n_255673036));
	notech_nand2 i_169846060(.A(n_255673036), .B(n_226072740), .Z(n_255773037
		));
	notech_ao4 i_168446074(.A(n_319937994), .B(n_247072950), .C(n_58082), .D
		(n_241572895), .Z(n_256073040));
	notech_ao4 i_168346075(.A(n_26918), .B(n_29775), .C(n_321438009), .D(n_28005
		), .Z(n_256273042));
	notech_nand3 i_168646072(.A(n_256073040), .B(n_256273042), .C(n_225672736
		), .Z(n_256373043));
	notech_ao4 i_168146077(.A(n_57873), .B(\nbus_11358[20] ), .C(n_58145), .D
		(n_60005), .Z(n_256473044));
	notech_ao4 i_167746081(.A(n_58082), .B(n_243072910), .C(n_58497), .D(n_253773017
		), .Z(n_256773047));
	notech_ao4 i_167646082(.A(n_321438009), .B(n_28004), .C(n_321538010), .D
		(n_313447724), .Z(n_256973049));
	notech_ao4 i_167346085(.A(n_58145), .B(n_60006), .C(n_26918), .D(n_29773
		), .Z(n_257173051));
	notech_and4 i_167546083(.A(n_257173051), .B(n_26622), .C(n_224072720), .D
		(n_224372723), .Z(n_257473054));
	notech_ao4 i_166146097(.A(n_58082), .B(n_245572935), .C(n_58497), .D(n_254673026
		), .Z(n_257573055));
	notech_ao4 i_166046098(.A(n_321438009), .B(n_28002), .C(n_313647722), .D
		(n_321538010), .Z(n_257773057));
	notech_ao4 i_165746101(.A(n_58145), .B(n_60008), .C(n_26918), .D(n_29772
		), .Z(n_257973059));
	notech_and4 i_165946099(.A(n_257973059), .B(n_26624), .C(n_223172711), .D
		(n_223472714), .Z(n_258273062));
	notech_ao4 i_154746207(.A(n_27329), .B(n_247072950), .C(n_144928726), .D
		(\nbus_11358[20] ), .Z(n_258373063));
	notech_ao4 i_154546209(.A(n_144828725), .B(\nbus_11365[20] ), .C(n_144428721
		), .D(n_313347725), .Z(n_258573065));
	notech_and4 i_154946205(.A(n_258573065), .B(n_258373063), .C(n_222772707
		), .D(n_223072710), .Z(n_258773067));
	notech_ao4 i_154246212(.A(n_60158), .B(n_27209), .C(n_145128728), .D(n_60005
		), .Z(n_258873068));
	notech_ao4 i_154046214(.A(n_54658), .B(n_29937), .C(n_32270), .D(n_28109
		), .Z(n_259073070));
	notech_and4 i_154446210(.A(n_259073070), .B(n_258873068), .C(n_222172701
		), .D(n_222472704), .Z(n_259273072));
	notech_ao4 i_153746217(.A(n_57160), .B(\nbus_11365[19] ), .C(n_144928726
		), .D(n_56311), .Z(n_259373073));
	notech_ao4 i_153646218(.A(n_243072910), .B(n_26803), .C(n_27329), .D(n_247972959
		), .Z(n_259473074));
	notech_ao4 i_153446220(.A(n_144428721), .B(n_313447724), .C(n_303791786)
		, .D(n_253773017), .Z(n_259673076));
	notech_and4 i_153946215(.A(n_259673076), .B(n_259473074), .C(n_259373073
		), .D(n_221472694), .Z(n_259873078));
	notech_ao4 i_153146223(.A(n_60158), .B(n_27208), .C(n_145128728), .D(n_60006
		), .Z(n_259973079));
	notech_ao4 i_152946225(.A(n_54658), .B(n_29936), .C(n_32270), .D(n_28108
		), .Z(n_260173081));
	notech_and4 i_153346221(.A(n_260173081), .B(n_259973079), .C(n_220872688
		), .D(n_221172691), .Z(n_260373083));
	notech_ao4 i_152646228(.A(n_57160), .B(\nbus_11365[18] ), .C(n_144928726
		), .D(\nbus_11358[18] ), .Z(n_260473084));
	notech_ao4 i_152546229(.A(n_95222216), .B(n_26803), .C(n_77522039), .D(n_27329
		), .Z(n_260573085));
	notech_ao4 i_152346231(.A(n_3861), .B(n_144428721), .C(n_303791786), .D(n_60121865
		), .Z(n_260773087));
	notech_and4 i_152846226(.A(n_260773087), .B(n_260573085), .C(n_260473084
		), .D(n_220172681), .Z(n_260973089));
	notech_ao4 i_152046234(.A(n_60158), .B(n_27207), .C(n_3864), .D(n_145128728
		), .Z(n_261073090));
	notech_ao4 i_151846236(.A(n_54658), .B(n_29935), .C(n_32270), .D(n_28107
		), .Z(n_261273092));
	notech_and4 i_152246232(.A(n_261273092), .B(n_261073090), .C(n_219572675
		), .D(n_219872678), .Z(n_261473094));
	notech_ao4 i_151546239(.A(n_57160), .B(\nbus_11365[17] ), .C(n_144928726
		), .D(n_56293), .Z(n_261573095));
	notech_ao4 i_151446240(.A(n_245572935), .B(n_26803), .C(n_27329), .D(n_249672976
		), .Z(n_261673096));
	notech_ao4 i_151146242(.A(n_144428721), .B(n_313647722), .C(n_303791786)
		, .D(n_254673026), .Z(n_261873098));
	notech_and4 i_151746237(.A(n_261873098), .B(n_261673096), .C(n_261573095
		), .D(n_218872668), .Z(n_262073100));
	notech_ao4 i_150846245(.A(n_60158), .B(n_27206), .C(n_60008), .D(n_145128728
		), .Z(n_262173101));
	notech_ao4 i_150646247(.A(n_54658), .B(n_29933), .C(n_32270), .D(n_28106
		), .Z(n_262373103));
	notech_and4 i_151046243(.A(n_262373103), .B(n_262173101), .C(n_218272662
		), .D(n_218572665), .Z(n_262573105));
	notech_ao4 i_149046262(.A(n_247072950), .B(n_151931934), .C(n_241572895)
		, .D(n_58084), .Z(n_262673106));
	notech_ao4 i_148946263(.A(n_26929), .B(n_29775), .C(n_58429), .D(n_28005
		), .Z(n_262873108));
	notech_nand3 i_149246260(.A(n_262673106), .B(n_262873108), .C(n_217972659
		), .Z(n_262973109));
	notech_ao4 i_148746265(.A(n_57875), .B(\nbus_11358[20] ), .C(n_58147), .D
		(n_60005), .Z(n_263073110));
	notech_ao4 i_148346269(.A(n_58498), .B(n_253773017), .C(n_241372893), .D
		(\nbus_11365[19] ), .Z(n_263373113));
	notech_ao4 i_148246270(.A(n_154831963), .B(n_313447724), .C(n_151931934)
		, .D(n_247972959), .Z(n_263573115));
	notech_ao4 i_147946273(.A(n_26929), .B(n_29773), .C(n_58429), .D(n_28004
		), .Z(n_263773117));
	notech_and4 i_148146271(.A(n_263773117), .B(n_26622), .C(n_216372643), .D
		(n_216672646), .Z(n_264073120));
	notech_ao4 i_147346277(.A(n_60121865), .B(n_58498), .C(n_241372893), .D(\nbus_11365[18] 
		), .Z(n_264173121));
	notech_ao4 i_147246278(.A(n_3861), .B(n_154831963), .C(n_77522039), .D(n_151931934
		), .Z(n_264373123));
	notech_ao4 i_146946281(.A(n_26929), .B(n_29711), .C(n_58429), .D(n_28003
		), .Z(n_264573125));
	notech_and4 i_147146279(.A(n_264573125), .B(n_26621), .C(n_215472634), .D
		(n_215772637), .Z(n_264873128));
	notech_ao4 i_146546285(.A(n_58498), .B(n_254673026), .C(n_241372893), .D
		(\nbus_11365[17] ), .Z(n_264973129));
	notech_ao4 i_146446286(.A(n_313647722), .B(n_154831963), .C(n_249672976)
		, .D(n_151931934), .Z(n_265173131));
	notech_ao4 i_146146289(.A(n_26929), .B(n_29772), .C(n_58429), .D(n_28002
		), .Z(n_265373133));
	notech_and4 i_146346287(.A(n_265373133), .B(n_26624), .C(n_214572625), .D
		(n_214872628), .Z(n_265673136));
	notech_ao4 i_137446370(.A(n_247072950), .B(n_3843), .C(n_3858), .D(n_241572895
		), .Z(n_265773137));
	notech_ao4 i_137346371(.A(n_26642), .B(n_29775), .C(n_3857), .D(n_28005)
		, .Z(n_265973139));
	notech_nand3 i_137646368(.A(n_265773137), .B(n_265973139), .C(n_214472624
		), .Z(n_266073140));
	notech_ao4 i_137146373(.A(n_3877), .B(\nbus_11358[20] ), .C(n_148228759)
		, .D(n_60005), .Z(n_266173141));
	notech_ao4 i_136746377(.A(n_3845), .B(n_253773017), .C(n_263180132), .D(\nbus_11365[19] 
		), .Z(n_266473144));
	notech_ao4 i_136546379(.A(n_3837), .B(n_313447724), .C(n_247972959), .D(n_3843
		), .Z(n_266673146));
	notech_and4 i_136946375(.A(n_213372613), .B(n_266673146), .C(n_266473144
		), .D(n_213672616), .Z(n_266873148));
	notech_ao4 i_136246382(.A(n_148228759), .B(n_60006), .C(n_26642), .D(n_29773
		), .Z(n_266973149));
	notech_and4 i_136446380(.A(n_125828535), .B(n_266973149), .C(n_26622), .D
		(n_213072610), .Z(n_267273152));
	notech_ao4 i_134946395(.A(n_3845), .B(n_254673026), .C(n_263180132), .D(\nbus_11365[17] 
		), .Z(n_267373153));
	notech_ao4 i_134746397(.A(n_313647722), .B(n_3837), .C(n_249672976), .D(n_3843
		), .Z(n_267573155));
	notech_and4 i_135146393(.A(n_212472604), .B(n_267573155), .C(n_267373153
		), .D(n_212772607), .Z(n_267773157));
	notech_ao4 i_134446400(.A(n_148228759), .B(n_60008), .C(n_26642), .D(n_29772
		), .Z(n_267873158));
	notech_and4 i_134646398(.A(n_125828535), .B(n_267873158), .C(n_26624), .D
		(n_212172601), .Z(n_268173161));
	notech_ao4 i_133146412(.A(n_247072950), .B(n_310791716), .C(n_241572895)
		, .D(n_310891715), .Z(n_268273162));
	notech_ao4 i_133046413(.A(n_149228769), .B(n_29775), .C(n_310691717), .D
		(n_28005), .Z(n_268473164));
	notech_and3 i_133346410(.A(n_268273162), .B(n_268473164), .C(n_211872598
		), .Z(n_268573165));
	notech_ao4 i_132746416(.A(n_56320), .B(n_149428771), .C(n_149128768), .D
		(n_60005), .Z(n_268673166));
	notech_ao4 i_132646417(.A(n_28109), .B(n_60329), .C(n_54643), .D(n_28976
		), .Z(n_268873168));
	notech_ao4 i_132246420(.A(n_243072910), .B(n_310891715), .C(n_311991704)
		, .D(n_253773017), .Z(n_269073170));
	notech_ao4 i_132046422(.A(n_57173), .B(n_57707), .C(n_148728764), .D(n_313447724
		), .Z(n_269273172));
	notech_and4 i_132546418(.A(n_210672586), .B(n_269273172), .C(n_269073170
		), .D(n_210972589), .Z(n_269473174));
	notech_ao4 i_131746425(.A(n_149128768), .B(n_60006), .C(n_149228769), .D
		(n_29773), .Z(n_269573175));
	notech_ao4 i_131646426(.A(n_28108), .B(n_60329), .C(n_54643), .D(n_28974
		), .Z(n_269773177));
	notech_ao4 i_131346429(.A(n_95222216), .B(n_310891715), .C(n_60121865), 
		.D(n_311991704), .Z(n_269973179));
	notech_ao4 i_131146431(.A(n_57173), .B(\nbus_11365[18] ), .C(n_3861), .D
		(n_148728764), .Z(n_270173181));
	notech_and4 i_131546427(.A(n_209672576), .B(n_270173181), .C(n_269973179
		), .D(n_209972579), .Z(n_270373183));
	notech_ao4 i_130846434(.A(n_3864), .B(n_149128768), .C(n_149228769), .D(n_29711
		), .Z(n_270473184));
	notech_ao4 i_130646436(.A(n_28107), .B(n_60329), .C(n_54643), .D(n_28972
		), .Z(n_270673186));
	notech_and4 i_131046432(.A(n_125828535), .B(n_270673186), .C(n_270473184
		), .D(n_209372573), .Z(n_270873188));
	notech_ao4 i_130346439(.A(n_245572935), .B(n_310891715), .C(n_311991704)
		, .D(n_254673026), .Z(n_270973189));
	notech_ao4 i_130146441(.A(n_57173), .B(n_57689), .C(n_148728764), .D(n_313647722
		), .Z(n_271173191));
	notech_and4 i_130546437(.A(n_208672566), .B(n_271173191), .C(n_270973189
		), .D(n_208972569), .Z(n_271373193));
	notech_ao4 i_129746444(.A(n_149128768), .B(n_60008), .C(n_149228769), .D
		(n_29772), .Z(n_271473194));
	notech_ao4 i_129646445(.A(n_28106), .B(n_60329), .C(n_54643), .D(n_28971
		), .Z(n_271673196));
	notech_ao4 i_128346458(.A(n_308791736), .B(n_247072950), .C(n_307891745)
		, .D(n_241572895), .Z(n_271873198));
	notech_ao4 i_128146460(.A(n_308591738), .B(n_28005), .C(n_60157), .D(n_27140
		), .Z(n_272073200));
	notech_and4 i_128546456(.A(n_272073200), .B(n_271873198), .C(n_207672556
		), .D(n_207972559), .Z(n_272273202));
	notech_ao4 i_127846463(.A(n_150728784), .B(n_60005), .C(n_150628783), .D
		(n_29775), .Z(n_272373203));
	notech_ao4 i_127746464(.A(n_26648), .B(n_29932), .C(n_150428781), .D(n_57720
		), .Z(n_272573205));
	notech_ao4 i_127446467(.A(n_307891745), .B(n_243072910), .C(n_306791756)
		, .D(n_253773017), .Z(n_272773207));
	notech_ao4 i_127246469(.A(n_60157), .B(n_27139), .C(n_150228779), .D(n_313447724
		), .Z(n_272973209));
	notech_and4 i_127646465(.A(n_272973209), .B(n_272773207), .C(n_206572545
		), .D(n_206872548), .Z(n_273173211));
	notech_ao4 i_126946472(.A(n_150628783), .B(n_29773), .C(n_59100), .D(n_28108
		), .Z(n_273273212));
	notech_ao4 i_126746474(.A(n_3836), .B(n_57707), .C(n_150528782), .D(n_56311
		), .Z(n_273473214));
	notech_and4 i_127146470(.A(n_273473214), .B(n_273273212), .C(n_206272542
		), .D(n_205972539), .Z(n_273673216));
	notech_ao4 i_125346488(.A(n_307891745), .B(n_245572935), .C(n_306791756)
		, .D(n_254673026), .Z(n_273773217));
	notech_ao4 i_125146490(.A(n_60157), .B(n_27137), .C(n_150228779), .D(n_313647722
		), .Z(n_273973219));
	notech_and4 i_125546486(.A(n_273973219), .B(n_273773217), .C(n_205372533
		), .D(n_205672536), .Z(n_274173221));
	notech_ao4 i_124746493(.A(n_150628783), .B(n_29772), .C(n_59100), .D(n_28106
		), .Z(n_274273222));
	notech_ao4 i_124546495(.A(n_3836), .B(n_57689), .C(n_150528782), .D(n_56293
		), .Z(n_274473224));
	notech_and4 i_124946491(.A(n_274473224), .B(n_274273222), .C(n_205072530
		), .D(n_204772527), .Z(n_274673226));
	notech_ao4 i_122846512(.A(n_311391710), .B(n_247072950), .C(n_311491709)
		, .D(n_241572895), .Z(n_274773227));
	notech_ao4 i_122646514(.A(n_151428791), .B(n_60005), .C(n_29775), .D(n_26696
		), .Z(n_274973229));
	notech_and4 i_123046510(.A(n_274973229), .B(n_274773227), .C(n_204172521
		), .D(n_204472524), .Z(n_275173231));
	notech_ao4 i_122346517(.A(n_311091713), .B(n_57720), .C(n_311191712), .D
		(n_56320), .Z(n_275273232));
	notech_nand2 i_122446516(.A(n_275273232), .B(n_203872518), .Z(n_275373233
		));
	notech_ao4 i_121946521(.A(n_253773017), .B(n_316491659), .C(n_57707), .D
		(n_306024324), .Z(n_275673236));
	notech_ao4 i_121746523(.A(n_151128788), .B(n_313447724), .C(n_311391710)
		, .D(n_247972959), .Z(n_275873238));
	notech_and4 i_122146519(.A(n_275873238), .B(n_275673236), .C(n_203172511
		), .D(n_203472514), .Z(n_276073240));
	notech_ao4 i_121446526(.A(n_311291711), .B(n_28004), .C(n_151428791), .D
		(n_60006), .Z(n_276173241));
	notech_ao4 i_121246528(.A(n_54643), .B(n_28956), .C(n_151028787), .D(nbus_11295
		[19]), .Z(n_276373243));
	notech_and4 i_121646524(.A(n_276373243), .B(n_202872508), .C(n_276173241
		), .D(n_26622), .Z(n_276573245));
	notech_ao4 i_119846541(.A(n_254673026), .B(n_316491659), .C(n_306024324)
		, .D(n_57689), .Z(n_276673246));
	notech_ao4 i_119646543(.A(n_151128788), .B(n_313647722), .C(n_311391710)
		, .D(n_249672976), .Z(n_276873248));
	notech_and4 i_120046539(.A(n_276873248), .B(n_276673246), .C(n_202072500
		), .D(n_202372503), .Z(n_277073250));
	notech_ao4 i_119346546(.A(n_28002), .B(n_311291711), .C(n_60008), .D(n_151428791
		), .Z(n_277173251));
	notech_ao4 i_119146548(.A(n_54643), .B(n_28954), .C(n_151028787), .D(nbus_11295
		[17]), .Z(n_277373253));
	notech_and4 i_119546544(.A(n_277373253), .B(n_201772497), .C(n_277173251
		), .D(n_26624), .Z(n_277573255));
	notech_or4 i_17044326(.A(n_60970), .B(n_60959), .C(n_60909), .D(n_29723)
		, .Z(n_277673256));
	notech_mux2 i_13044366(.S(n_32322), .A(n_305721221), .B(n_305621220), .Z
		(n_277873258));
	notech_and2 i_13144365(.A(n_92519107), .B(n_318173661), .Z(n_277973259)
		);
	notech_and3 i_12944367(.A(n_58082), .B(n_57765), .C(n_289073370), .Z(n_278273262
		));
	notech_ao4 i_5844436(.A(n_58505), .B(n_57500), .C(n_58421), .D(n_304573525
		), .Z(n_278373263));
	notech_mux2 i_12744369(.S(n_32325), .A(n_305721221), .B(n_305621220), .Z
		(n_278673266));
	notech_and2 i_12844368(.A(n_92519107), .B(n_316073640), .Z(n_278773267)
		);
	notech_and2 i_12544371(.A(n_58085), .B(n_279373273), .Z(n_279073270));
	notech_and4 i_5244442(.A(n_56848), .B(n_125961542), .C(n_58477), .D(n_58493
		), .Z(n_279173271));
	notech_ao4 i_12644370(.A(n_59435), .B(\nbus_11307[7] ), .C(n_304373523),
		 .D(n_26784), .Z(n_279273272));
	notech_or4 i_81243718(.A(n_57026), .B(n_30854), .C(n_57827), .D(n_29653)
		, .Z(n_279373273));
	notech_mux2 i_11944376(.S(n_32331), .A(n_305721221), .B(n_305621220), .Z
		(n_279573275));
	notech_and2 i_12044375(.A(n_92519107), .B(n_314273622), .Z(n_279673276)
		);
	notech_nor2 i_263255552(.A(n_209069102), .B(n_26884), .Z(n_280073280));
	notech_and4 i_11844377(.A(n_58285), .B(n_293473414), .C(n_293773417), .D
		(n_313273612), .Z(n_280173281));
	notech_mux2 i_11544380(.S(n_32332), .A(n_305721221), .B(n_305621220), .Z
		(n_280273282));
	notech_and2 i_11644379(.A(n_92519107), .B(n_312473604), .Z(n_280373283)
		);
	notech_and2 i_11344382(.A(n_228579786), .B(n_281073290), .Z(n_280773287)
		);
	notech_nor2 i_102250712(.A(n_281173291), .B(n_26828), .Z(n_280873288));
	notech_and3 i_11444381(.A(n_58285), .B(n_295873438), .C(n_311473594), .Z
		(n_280973289));
	notech_nao3 i_98143564(.A(n_281173291), .B(n_32332), .C(n_58100), .Z(n_281073290
		));
	notech_nand2 i_101850713(.A(n_58503), .B(n_58495), .Z(n_281173291));
	notech_mux2 i_11144384(.S(n_32338), .A(n_305721221), .B(n_305621220), .Z
		(n_281273292));
	notech_and2 i_11244383(.A(n_92519107), .B(n_310173581), .Z(n_281373293)
		);
	notech_and2 i_11044385(.A(n_305973539), .B(n_92619108), .Z(n_281673296)
		);
	notech_ao4 i_8844406(.A(n_59419), .B(n_29723), .C(n_60893), .D(n_281973299
		), .Z(n_281773297));
	notech_mux2 i_4344451(.S(n_32365), .A(n_29723), .B(n_3874), .Z(n_281973299
		));
	notech_or2 i_55243955(.A(n_58071), .B(n_60022), .Z(n_284873328));
	notech_or2 i_54943958(.A(n_57812), .B(\nbus_11358[3] ), .Z(n_285173331)
		);
	notech_or2 i_54643961(.A(n_211169123), .B(n_308721251), .Z(n_285473334)
		);
	notech_or4 i_54343964(.A(n_56508), .B(n_26601), .C(nbus_11295[3]), .D(n_60947
		), .Z(n_285773337));
	notech_or2 i_56443943(.A(n_60020), .B(n_58071), .Z(n_286073340));
	notech_or2 i_56143946(.A(n_57812), .B(\nbus_11358[5] ), .Z(n_286373343)
		);
	notech_or4 i_55843949(.A(n_56837), .B(n_26610), .C(n_308621250), .D(n_56513
		), .Z(n_286673346));
	notech_or4 i_55543952(.A(n_56508), .B(nbus_11295[5]), .C(n_60947), .D(n_26601
		), .Z(n_286973349));
	notech_or4 i_72843796(.A(n_58489), .B(n_58810), .C(n_60947), .D(n_28131)
		, .Z(n_287073350));
	notech_or4 i_72343801(.A(n_58810), .B(n_26906), .C(n_60947), .D(nbus_11295
		[6]), .Z(n_287773357));
	notech_nor2 i_74543780(.A(n_321438009), .B(n_27990), .Z(n_288073360));
	notech_nao3 i_74443781(.A(n_318891635), .B(n_318791636), .C(n_57947), .Z
		(n_288373363));
	notech_or2 i_74143784(.A(n_278373263), .B(\nbus_11307[7] ), .Z(n_288673366
		));
	notech_or2 i_73843787(.A(n_285080351), .B(n_303191792), .Z(n_288973369)
		);
	notech_nao3 i_74643779(.A(n_30945), .B(n_190062172), .C(n_58505), .Z(n_289073370
		));
	notech_or2 i_79343736(.A(n_58047), .B(\nbus_11358[6] ), .Z(n_289573375)
		);
	notech_or4 i_79043739(.A(n_58806), .B(n_58162), .C(n_60947), .D(nbus_11295
		[6]), .Z(n_289873378));
	notech_nao3 i_78743742(.A(n_58806), .B(n_26676), .C(n_58162), .Z(n_290173381
		));
	notech_nao3 i_80943721(.A(n_26824), .B(\opa_12[7] ), .C(n_26804), .Z(n_290873388
		));
	notech_nao3 i_80543724(.A(n_318791636), .B(n_319191632), .C(n_57947), .Z
		(n_291173391));
	notech_or4 i_80243727(.A(n_26804), .B(n_58806), .C(n_60949), .D(n_28133)
		, .Z(n_291473394));
	notech_or4 i_90743634(.A(n_58099), .B(n_280073280), .C(n_32331), .D(\nbus_11307[6] 
		), .Z(n_291573395));
	notech_ao4 i_90143639(.A(n_209069102), .B(n_26884), .C(n_26677), .D(n_314173621
		), .Z(n_292273402));
	notech_or2 i_92043621(.A(n_57084), .B(n_303191792), .Z(n_292773407));
	notech_nao3 i_92443617(.A(n_56437), .B(opa[7]), .C(n_58099), .Z(n_293473414
		));
	notech_or2 i_92343618(.A(n_57322), .B(\nbus_11358[7] ), .Z(n_293773417)
		);
	notech_or4 i_96343579(.A(n_58100), .B(n_26807), .C(n_32332), .D(\nbus_11307[6] 
		), .Z(n_293873418));
	notech_ao4 i_95743584(.A(n_281173291), .B(n_26828), .C(n_26677), .D(n_312373603
		), .Z(n_294573425));
	notech_ao3 i_98043565(.A(n_26737), .B(n_58487), .C(n_303191792), .Z(n_295073430
		));
	notech_ao3 i_97543570(.A(n_62798), .B(opc_10[7]), .C(n_57139), .Z(n_295773437
		));
	notech_nao3 i_98443561(.A(n_56448), .B(opa[7]), .C(n_58100), .Z(n_295873438
		));
	notech_or4 i_103343513(.A(n_58087), .B(n_56529), .C(n_32338), .D(\nbus_11307[6] 
		), .Z(n_296173441));
	notech_or2 i_103243514(.A(n_58044), .B(\nbus_11358[6] ), .Z(n_296473444)
		);
	notech_nao3 i_102943517(.A(n_62798), .B(opc[6]), .C(n_123971719), .Z(n_296773447
		));
	notech_or4 i_102643520(.A(n_62864), .B(n_124171721), .C(n_60949), .D(\nbus_11307[6] 
		), .Z(n_297073450));
	notech_nao3 i_104143506(.A(n_60329), .B(opa[6]), .C(n_3852), .Z(n_297173451
		));
	notech_or4 i_107843471(.A(n_317391650), .B(n_317091653), .C(n_60022), .D
		(n_56401), .Z(n_297873458));
	notech_or4 i_110943440(.A(n_317391650), .B(n_317091653), .C(n_60020), .D
		(n_56401), .Z(n_299373473));
	notech_or4 i_114143411(.A(n_317391650), .B(n_56533), .C(n_32365), .D(\nbus_11307[6] 
		), .Z(n_300873488));
	notech_nao3 i_113843414(.A(n_19065), .B(read_data[6]), .C(n_59100), .Z(n_301173491
		));
	notech_nand2 i_113543417(.A(add_len_pc[6]), .B(n_26766), .Z(n_301473494)
		);
	notech_or4 i_118643375(.A(n_317391650), .B(n_317091653), .C(n_303191792)
		, .D(n_56401), .Z(n_302373503));
	notech_or4 i_33058(.A(n_246891941), .B(n_2479), .C(n_56837), .D(n_26610)
		, .Z(n_303673516));
	notech_or2 i_10144393(.A(n_58810), .B(n_26906), .Z(n_303773517));
	notech_nand2 i_9844396(.A(n_58810), .B(n_58167), .Z(n_303873518));
	notech_or4 i_31339(.A(n_59387), .B(n_29178), .C(n_27198), .D(n_26810), .Z
		(n_303973519));
	notech_nand2 i_31329(.A(n_58810), .B(n_26908), .Z(n_304073520));
	notech_or4 i_6644428(.A(n_32326), .B(n_58133), .C(n_26906), .D(n_26735),
		 .Z(n_304173521));
	notech_or4 i_31124(.A(n_59387), .B(n_32356), .C(n_29178), .D(n_27198), .Z
		(n_304273522));
	notech_nao3 i_6544429(.A(n_62798), .B(opa[7]), .C(n_62848), .Z(n_304373523
		));
	notech_or2 i_106344540(.A(n_295921141), .B(n_26906), .Z(n_304473524));
	notech_and2 i_2744466(.A(n_58481), .B(n_58497), .Z(n_304573525));
	notech_ao4 i_210642484(.A(n_286163128), .B(n_31309), .C(n_285963126), .D
		(n_304373523), .Z(n_304673526));
	notech_ao4 i_210542485(.A(n_317091653), .B(n_31279), .C(n_286063127), .D
		(n_31307), .Z(n_304773527));
	notech_ao4 i_210342487(.A(n_122628503), .B(n_29544), .C(n_56533), .D(n_58285
		), .Z(n_304973529));
	notech_ao4 i_210242488(.A(n_60157), .B(n_27252), .C(n_317991644), .D(n_303391790
		), .Z(n_305073530));
	notech_and4 i_210842482(.A(n_305073530), .B(n_304973529), .C(n_304773527
		), .D(n_304673526), .Z(n_305273532));
	notech_ao4 i_209942491(.A(n_309191732), .B(n_29949), .C(n_309291731), .D
		(n_28096), .Z(n_305373533));
	notech_ao4 i_209842492(.A(n_58081), .B(\nbus_11358[7] ), .C(n_58406), .D
		(n_27990), .Z(n_305473534));
	notech_ao4 i_209642494(.A(n_286363130), .B(n_29614), .C(n_285663123), .D
		(\nbus_11307[7] ), .Z(n_305673536));
	notech_and4 i_210142489(.A(n_305673536), .B(n_305473534), .C(n_305373533
		), .D(n_302373503), .Z(n_305873538));
	notech_ao4 i_209542495(.A(n_60868), .B(n_281973299), .C(n_32393), .D(n_281773297
		), .Z(n_305973539));
	notech_nao3 i_5944435(.A(n_62826), .B(opa[6]), .C(n_62848), .Z(n_306073540
		));
	notech_ao4 i_207842512(.A(n_285963126), .B(n_306073540), .C(n_317091653)
		, .D(n_281673296), .Z(n_306173541));
	notech_or4 i_5044444(.A(n_60970), .B(n_60959), .C(n_62848), .D(\nbus_11307[6] 
		), .Z(n_306273542));
	notech_ao4 i_207742513(.A(n_286163128), .B(n_92019102), .C(n_56533), .D(n_306273542
		), .Z(n_306373543));
	notech_ao4 i_207542515(.A(n_3868), .B(n_317991644), .C(n_26802), .D(n_286063127
		), .Z(n_306573545));
	notech_and4 i_208042510(.A(n_306573545), .B(n_306373543), .C(n_306173541
		), .D(n_301473494), .Z(n_306773547));
	notech_ao4 i_207242518(.A(n_58406), .B(n_27989), .C(n_60158), .D(n_27251
		), .Z(n_306873548));
	notech_ao4 i_207042520(.A(n_58081), .B(\nbus_11358[6] ), .C(n_309191732)
		, .D(n_29948), .Z(n_307073550));
	notech_and4 i_207442516(.A(n_307073550), .B(n_306873548), .C(n_300873488
		), .D(n_301173491), .Z(n_307273552));
	notech_ao4 i_205342537(.A(n_281966348), .B(n_56533), .C(n_281866347), .D
		(n_285963126), .Z(n_307373553));
	notech_ao4 i_205242538(.A(n_282166350), .B(n_286163128), .C(n_282066349)
		, .D(n_286063127), .Z(n_307473554));
	notech_ao4 i_205042540(.A(n_308621250), .B(n_317991644), .C(n_282266351)
		, .D(n_317091653), .Z(n_307673556));
	notech_ao4 i_204942541(.A(n_60157), .B(n_27250), .C(n_122628503), .D(n_29543
		), .Z(n_307773557));
	notech_and4 i_205542535(.A(n_307773557), .B(n_307673556), .C(n_307473554
		), .D(n_307373553), .Z(n_307973559));
	notech_ao4 i_204642544(.A(n_309191732), .B(n_29947), .C(n_309291731), .D
		(n_28094), .Z(n_308073560));
	notech_ao4 i_204542545(.A(n_58081), .B(\nbus_11358[5] ), .C(n_58406), .D
		(n_27987), .Z(n_308173561));
	notech_ao4 i_204342547(.A(n_286363130), .B(n_29651), .C(n_285663123), .D
		(\nbus_11307[5] ), .Z(n_308373563));
	notech_and4 i_204842542(.A(n_308373563), .B(n_308173561), .C(n_308073560
		), .D(n_299373473), .Z(n_308573565));
	notech_ao4 i_202642564(.A(n_306670077), .B(n_285963126), .C(n_306570076)
		, .D(n_56533), .Z(n_308673566));
	notech_ao4 i_202542565(.A(n_286163128), .B(n_306870079), .C(n_306770078)
		, .D(n_286063127), .Z(n_308773567));
	notech_ao4 i_202342567(.A(n_308721251), .B(n_317991644), .C(n_306970080)
		, .D(n_317091653), .Z(n_308973569));
	notech_ao4 i_202242568(.A(n_60157), .B(n_27248), .C(n_122628503), .D(n_29541
		), .Z(n_309073570));
	notech_and4 i_202842562(.A(n_309073570), .B(n_308973569), .C(n_308773567
		), .D(n_308673566), .Z(n_309273572));
	notech_ao4 i_201942571(.A(n_309191732), .B(n_29946), .C(n_309291731), .D
		(n_28092), .Z(n_309373573));
	notech_ao4 i_201842572(.A(n_58081), .B(\nbus_11358[3] ), .C(n_58406), .D
		(n_27985), .Z(n_309473574));
	notech_ao4 i_201642574(.A(n_286363130), .B(n_29728), .C(n_285663123), .D
		(\nbus_11307[3] ), .Z(n_309673576));
	notech_and4 i_202142569(.A(n_297873458), .B(n_309673576), .C(n_309473574
		), .D(n_309373573), .Z(n_309873578));
	notech_nand3 i_4944445(.A(n_62826), .B(n_62848), .C(\opa_12[6] ), .Z(n_309973579
		));
	notech_nao3 i_4844446(.A(n_62864), .B(n_62822), .C(n_3874), .Z(n_310073580
		));
	notech_mux2 i_200542585(.S(n_32338), .A(n_309973579), .B(n_310073580), .Z
		(n_310173581));
	notech_ao4 i_199942590(.A(n_124071720), .B(n_281373293), .C(n_58488), .D
		(n_281273292), .Z(n_310273582));
	notech_ao4 i_199742592(.A(n_92019102), .B(n_153979043), .C(n_56529), .D(n_306273542
		), .Z(n_310473584));
	notech_and4 i_200242588(.A(n_310473584), .B(n_297073450), .C(n_310273582
		), .D(n_296773447), .Z(n_310673586));
	notech_ao4 i_199442595(.A(n_123771717), .B(n_27989), .C(n_3868), .D(n_124271722
		), .Z(n_310773587));
	notech_ao4 i_200442586(.A(n_60329), .B(n_28095), .C(n_58391), .D(n_29723
		), .Z(n_310973589));
	notech_and3 i_76944480(.A(n_3873), .B(n_310973589), .C(n_297173451), .Z(n_311173591
		));
	notech_and4 i_199642593(.A(n_311173591), .B(n_310773587), .C(n_296173441
		), .D(n_296473444), .Z(n_311373593));
	notech_mux2 i_195942630(.S(n_58817), .A(n_31307), .B(n_304373523), .Z(n_311473594
		));
	notech_ao4 i_195542634(.A(n_280973289), .B(n_280873288), .C(\nbus_11358[7] 
		), .D(n_280773287), .Z(n_311673596));
	notech_ao4 i_195442635(.A(n_57947), .B(n_26924), .C(n_31279), .D(n_26816
		), .Z(n_311873598));
	notech_nao3 i_195742632(.A(n_311673596), .B(n_311873598), .C(n_295773437
		), .Z(n_311973599));
	notech_ao4 i_195242637(.A(n_153879042), .B(n_29614), .C(n_58424), .D(n_27990
		), .Z(n_312073600));
	notech_mux2 i_194942640(.S(n_58817), .A(n_91719099), .B(n_26676), .Z(n_312373603
		));
	notech_mux2 i_195042639(.S(n_32332), .A(n_309973579), .B(n_310073580), .Z
		(n_312473604));
	notech_ao4 i_194642643(.A(n_143071910), .B(n_280373283), .C(n_280273282)
		, .D(n_26816), .Z(n_312573605));
	notech_ao4 i_194542644(.A(n_3868), .B(n_143571915), .C(n_92019102), .D(n_57139
		), .Z(n_312773607));
	notech_ao3 i_194842641(.A(n_312573605), .B(n_312773607), .C(n_294573425)
		, .Z(n_312873608));
	notech_ao4 i_194342646(.A(n_57573), .B(\nbus_11358[6] ), .C(n_143471914)
		, .D(n_27989), .Z(n_312973609));
	notech_mux2 i_191342676(.S(n_58805), .A(n_31307), .B(n_304373523), .Z(n_313273612
		));
	notech_ao4 i_191042679(.A(n_31309), .B(n_57141), .C(n_280173281), .D(n_280073280
		), .Z(n_313573615));
	notech_ao4 i_190942680(.A(n_58425), .B(n_27990), .C(n_58486), .D(n_31279
		), .Z(n_313673616));
	notech_ao4 i_190742682(.A(n_247679977), .B(n_29614), .C(n_57947), .D(n_56653
		), .Z(n_313873618));
	notech_and3 i_190842681(.A(n_313873618), .B(n_26708), .C(n_292773407), .Z
		(n_314073620));
	notech_mux2 i_190442685(.S(n_58805), .A(n_91719099), .B(n_26676), .Z(n_314173621
		));
	notech_mux2 i_190542684(.S(n_32331), .A(n_309973579), .B(n_310073580), .Z
		(n_314273622));
	notech_ao4 i_190142688(.A(n_178472264), .B(n_279673276), .C(n_58486), .D
		(n_279573275), .Z(n_314373623));
	notech_ao4 i_190042689(.A(n_3868), .B(n_147271952), .C(n_92019102), .D(n_57141
		), .Z(n_314573625));
	notech_ao3 i_190342686(.A(n_314373623), .B(n_314573625), .C(n_292273402)
		, .Z(n_314673626));
	notech_ao4 i_189842691(.A(n_57154), .B(\nbus_11358[6] ), .C(n_147171951)
		, .D(n_27989), .Z(n_314773627));
	notech_ao4 i_182842761(.A(n_279273272), .B(n_279173271), .C(n_31307), .D
		(n_279073270), .Z(n_315073630));
	notech_ao4 i_182642763(.A(n_58427), .B(n_27990), .C(n_26804), .D(n_31279
		), .Z(n_315273632));
	notech_and4 i_183042759(.A(n_315273632), .B(n_315073630), .C(n_291173391
		), .D(n_291473394), .Z(n_315473634));
	notech_ao4 i_182342766(.A(n_153479038), .B(\nbus_11307[7] ), .C(n_58047)
		, .D(\nbus_11358[7] ), .Z(n_315573635));
	notech_ao4 i_182142768(.A(n_154331958), .B(nbus_11295[7]), .C(n_153579039
		), .D(n_303191792), .Z(n_315773637));
	notech_and4 i_182542764(.A(n_315773637), .B(n_315573635), .C(n_290873388
		), .D(n_26708), .Z(n_315973639));
	notech_mux2 i_182042769(.S(n_32325), .A(n_309973579), .B(n_310073580), .Z
		(n_316073640));
	notech_ao4 i_181742772(.A(n_278773267), .B(n_147471954), .C(n_26804), .D
		(n_278673266), .Z(n_316173641));
	notech_ao4 i_181542774(.A(n_92019102), .B(n_257980080), .C(n_58162), .D(n_306273542
		), .Z(n_316373643));
	notech_and4 i_181942770(.A(n_316373643), .B(n_290173381), .C(n_316173641
		), .D(n_289873378), .Z(n_316573645));
	notech_ao4 i_181242777(.A(n_27989), .B(n_153179035), .C(n_3868), .D(n_153779041
		), .Z(n_316673646));
	notech_ao4 i_181042779(.A(n_154331958), .B(nbus_11295[6]), .C(n_153479038
		), .D(\nbus_11307[6] ), .Z(n_316873648));
	notech_and4 i_181442775(.A(n_311173591), .B(n_316873648), .C(n_316673646
		), .D(n_289573375), .Z(n_317073650));
	notech_ao4 i_177742811(.A(n_284980350), .B(n_29614), .C(n_31307), .D(n_278273262
		), .Z(n_317273652));
	notech_ao4 i_177542813(.A(n_31309), .B(n_57923), .C(n_304173521), .D(\nbus_11358[7] 
		), .Z(n_317473654));
	notech_and4 i_177942809(.A(n_317473654), .B(n_317273652), .C(n_288673366
		), .D(n_288973369), .Z(n_317673656));
	notech_ao4 i_177242816(.A(n_58489), .B(n_31279), .C(n_304573525), .D(n_58285
		), .Z(n_317773657));
	notech_nand2 i_177342815(.A(n_317773657), .B(n_288373363), .Z(n_317873658
		));
	notech_mux2 i_177042818(.S(n_32322), .A(n_309973579), .B(n_310073580), .Z
		(n_318173661));
	notech_ao4 i_176742821(.A(n_304073520), .B(n_277973259), .C(n_58489), .D
		(n_277873258), .Z(n_318273662));
	notech_ao4 i_176642822(.A(n_278373263), .B(\nbus_11307[6] ), .C(n_304173521
		), .D(\nbus_11358[6] ), .Z(n_318473664));
	notech_and3 i_176942819(.A(n_318273662), .B(n_318473664), .C(n_287773357
		), .Z(n_318573665));
	notech_ao4 i_176442824(.A(n_304573525), .B(n_306273542), .C(n_302621190)
		, .D(n_26920), .Z(n_318673666));
	notech_ao4 i_161142976(.A(n_281966348), .B(n_56508), .C(n_281866347), .D
		(n_184168858), .Z(n_318973669));
	notech_ao4 i_160942978(.A(n_282266351), .B(n_305191772), .C(n_282166350)
		, .D(n_343270443), .Z(n_319173671));
	notech_and4 i_161342974(.A(n_319173671), .B(n_318973669), .C(n_286673346
		), .D(n_286973349), .Z(n_319373673));
	notech_ao4 i_160642981(.A(n_58370), .B(n_27987), .C(n_184968866), .D(n_28094
		), .Z(n_319473674));
	notech_ao4 i_160442983(.A(n_57821), .B(n_29651), .C(n_57711), .D(\nbus_11307[5] 
		), .Z(n_319673676));
	notech_and4 i_160842979(.A(n_319673676), .B(n_319473674), .C(n_286073340
		), .D(n_286373343), .Z(n_319873678));
	notech_ao4 i_160142986(.A(n_184168858), .B(n_306670077), .C(n_56508), .D
		(n_306570076), .Z(n_319973679));
	notech_ao4 i_159942988(.A(n_306970080), .B(n_305191772), .C(n_343270443)
		, .D(n_306870079), .Z(n_320173681));
	notech_and4 i_160342984(.A(n_320173681), .B(n_319973679), .C(n_285473334
		), .D(n_285773337), .Z(n_320373683));
	notech_ao4 i_159642991(.A(n_58370), .B(n_27985), .C(n_184968866), .D(n_28092
		), .Z(n_320473684));
	notech_ao4 i_159442993(.A(n_57821), .B(n_29728), .C(n_57711), .D(\nbus_11307[3] 
		), .Z(n_320673686));
	notech_and4 i_159842989(.A(n_320673686), .B(n_320473684), .C(n_284873328
		), .D(n_285173331), .Z(n_320873688));
	notech_ao4 i_146543110(.A(n_306570076), .B(n_56512), .C(n_306670077), .D
		(n_281566344), .Z(n_320973689));
	notech_ao4 i_146443111(.A(n_306870079), .B(n_236065889), .C(n_306770078)
		, .D(n_111464643), .Z(n_321073690));
	notech_ao4 i_146043113(.A(n_308721251), .B(n_111564644), .C(n_306970080)
		, .D(n_26614), .Z(n_321273692));
	notech_ao4 i_145943114(.A(n_57885), .B(\nbus_11358[3] ), .C(n_57886), .D
		(\nbus_11307[3] ), .Z(n_321373693));
	notech_and4 i_146743108(.A(n_321373693), .B(n_321273692), .C(n_321073690
		), .D(n_320973689), .Z(n_321573695));
	notech_ao4 i_145643117(.A(n_28092), .B(n_54874), .C(n_60158), .D(n_27158
		), .Z(n_321673696));
	notech_ao4 i_145343118(.A(n_57999), .B(n_29728), .C(n_58367), .D(n_27985
		), .Z(n_321773697));
	notech_ao4 i_145143120(.A(n_54865), .B(n_29945), .C(n_60022), .D(n_58000
		), .Z(n_321973699));
	notech_ao4 i_145043121(.A(n_54894), .B(n_27428), .C(n_54883), .D(n_28596
		), .Z(n_322073700));
	notech_and4 i_145843115(.A(n_322073700), .B(n_321973699), .C(n_321773697
		), .D(n_321673696), .Z(n_322273702));
	notech_or4 i_128364486(.A(n_57082), .B(n_57055), .C(n_26770), .D(n_58482
		), .Z(n_322373703));
	notech_or2 i_100240326(.A(n_4011), .B(n_56489), .Z(n_322673706));
	notech_nao3 i_100340325(.A(n_58173), .B(n_30946), .C(n_30854), .Z(n_322773707
		));
	notech_or2 i_49240789(.A(n_5933), .B(n_57329), .Z(n_322873708));
	notech_or2 i_49040790(.A(n_58054), .B(\nbus_11358[8] ), .Z(n_323173711)
		);
	notech_or4 i_48440795(.A(n_58802), .B(n_28134), .C(n_60949), .D(n_58482)
		, .Z(n_323673716));
	notech_nao3 i_63840654(.A(n_11404), .B(n_32272), .C(n_2868), .Z(n_323973719
		));
	notech_nand2 i_33176(.A(n_26811), .B(n_26662), .Z(n_325273732));
	notech_ao4 i_169439693(.A(n_286163128), .B(n_298066509), .C(n_286363130)
		, .D(n_29678), .Z(n_325373733));
	notech_ao4 i_169339694(.A(n_285963126), .B(n_297866507), .C(n_286063127)
		, .D(n_297966508), .Z(n_325473734));
	notech_ao4 i_169139696(.A(n_317091653), .B(n_297666505), .C(n_285663123)
		, .D(\nbus_11307[1] ), .Z(n_325673736));
	notech_ao4 i_169039697(.A(n_58406), .B(n_27983), .C(n_56533), .D(n_297766506
		), .Z(n_325773737));
	notech_and4 i_169639691(.A(n_325773737), .B(n_325673736), .C(n_325473734
		), .D(n_325373733), .Z(n_325973739));
	notech_ao4 i_168739700(.A(n_122628503), .B(n_29539), .C(n_58081), .D(\nbus_11358[1] 
		), .Z(n_326073740));
	notech_ao4 i_168639701(.A(n_27247), .B(n_60162), .C(n_317991644), .D(n_59992
		), .Z(n_326173741));
	notech_ao4 i_168439703(.A(n_309291731), .B(n_28090), .C(n_316991654), .D
		(n_60024), .Z(n_326373743));
	notech_and4 i_168939698(.A(n_323973719), .B(n_326373743), .C(n_326173741
		), .D(n_326073740), .Z(n_326573745));
	notech_ao4 i_157839803(.A(n_308166610), .B(n_58482), .C(n_325270263), .D
		(n_56485), .Z(n_326673746));
	notech_ao4 i_157739804(.A(n_325273732), .B(n_29787), .C(n_309666625), .D
		(n_58040), .Z(n_326873748));
	notech_ao4 i_157439807(.A(\nbus_11307[8] ), .B(n_26679), .C(n_27991), .D
		(n_26680), .Z(n_327073750));
	notech_and4 i_157639805(.A(n_334480845), .B(n_322873708), .C(n_327073750
		), .D(n_323173711), .Z(n_327373753));
	notech_or2 i_44037820(.A(n_53612636), .B(n_60008), .Z(n_327873758));
	notech_or2 i_43737823(.A(n_54212642), .B(n_57689), .Z(n_328173761));
	notech_or2 i_47037796(.A(n_53612636), .B(n_60006), .Z(n_329073770));
	notech_or2 i_46737799(.A(n_54212642), .B(n_57707), .Z(n_329373773));
	notech_or2 i_48237784(.A(n_53612636), .B(n_60005), .Z(n_330273782));
	notech_or2 i_47937787(.A(n_54212642), .B(n_57720), .Z(n_330573785));
	notech_ao4 i_214036168(.A(n_27094), .B(n_28421), .C(n_26950), .D(n_28562
		), .Z(n_337473854));
	notech_ao4 i_213936169(.A(n_56909), .B(n_29930), .C(n_56428), .D(n_28357
		), .Z(n_337573855));
	notech_ao4 i_213736171(.A(n_56448), .B(n_28225), .C(n_56437), .D(n_28192
		), .Z(n_337773857));
	notech_ao4 i_213636172(.A(n_56457), .B(n_28259), .C(n_28453), .D(n_27089
		), .Z(n_337873858));
	notech_and4 i_214236166(.A(n_337873858), .B(n_337773857), .C(n_337573855
		), .D(n_337473854), .Z(n_338073860));
	notech_ao4 i_213336175(.A(n_59349), .B(n_28518), .C(n_28324), .D(n_26664
		), .Z(n_338173861));
	notech_ao4 i_213236176(.A(n_56401), .B(n_28160), .C(n_28389), .D(n_56391
		), .Z(n_338273862));
	notech_and2 i_213436174(.A(n_338273862), .B(n_338173861), .Z(n_338373863
		));
	notech_ao4 i_213036178(.A(n_58014), .B(n_27860), .C(n_56468), .D(n_29931
		), .Z(n_338473864));
	notech_ao4 i_212936179(.A(n_57985), .B(n_28291), .C(n_28485), .D(n_27104
		), .Z(n_338573865));
	notech_ao4 i_187436434(.A(n_27094), .B(n_28436), .C(n_26950), .D(n_28578
		), .Z(n_338873868));
	notech_ao4 i_187336435(.A(n_56909), .B(n_29938), .C(n_56428), .D(n_28372
		), .Z(n_338973869));
	notech_ao4 i_187136437(.A(n_56448), .B(n_28242), .C(n_56437), .D(n_28207
		), .Z(n_339173871));
	notech_ao4 i_187036438(.A(n_56457), .B(n_28274), .C(n_28468), .D(n_27089
		), .Z(n_339273872));
	notech_and4 i_187636432(.A(n_339273872), .B(n_339173871), .C(n_338973869
		), .D(n_338873868), .Z(n_339473874));
	notech_ao4 i_186736441(.A(n_59349), .B(n_28538), .C(n_28340), .D(n_26664
		), .Z(n_339573875));
	notech_ao4 i_186636442(.A(n_56401), .B(n_28175), .C(n_28404), .D(n_56391
		), .Z(n_339673876));
	notech_and2 i_186836440(.A(n_339673876), .B(n_339573875), .Z(n_339773877
		));
	notech_ao4 i_186436444(.A(n_58014), .B(n_27875), .C(n_56468), .D(n_29939
		), .Z(n_339873878));
	notech_ao4 i_186336445(.A(n_57985), .B(n_28307), .C(n_28500), .D(n_27104
		), .Z(n_339973879));
	notech_ao4 i_186036448(.A(n_27094), .B(n_28438), .C(n_26950), .D(n_28580
		), .Z(n_340273882));
	notech_ao4 i_185936449(.A(n_56909), .B(n_29941), .C(n_56428), .D(n_28374
		), .Z(n_340373883));
	notech_ao4 i_185736451(.A(n_56448), .B(n_28244), .C(n_56437), .D(n_28209
		), .Z(n_340573885));
	notech_ao4 i_185636452(.A(n_56457), .B(n_28276), .C(n_28470), .D(n_27089
		), .Z(n_340673886));
	notech_and4 i_186236446(.A(n_340673886), .B(n_340573885), .C(n_340373883
		), .D(n_340273882), .Z(n_340873888));
	notech_ao4 i_185336455(.A(n_59349), .B(n_28540), .C(n_28342), .D(n_26664
		), .Z(n_340973889));
	notech_ao4 i_185236456(.A(n_56401), .B(n_28177), .C(n_28406), .D(n_56391
		), .Z(n_341073890));
	notech_and2 i_185436454(.A(n_341073890), .B(n_340973889), .Z(n_341173891
		));
	notech_ao4 i_185036458(.A(n_58014), .B(n_27878), .C(n_56468), .D(n_29942
		), .Z(n_341273892));
	notech_ao4 i_184936459(.A(n_57985), .B(n_28309), .C(n_28503), .D(n_27104
		), .Z(n_341373893));
	notech_ao4 i_184636462(.A(n_27094), .B(n_28439), .C(n_26950), .D(n_28581
		), .Z(n_341673896));
	notech_ao4 i_184536463(.A(n_56909), .B(n_29943), .C(n_56428), .D(n_28375
		), .Z(n_341773897));
	notech_ao4 i_184336465(.A(n_56448), .B(n_28245), .C(n_56437), .D(n_28210
		), .Z(n_341973899));
	notech_ao4 i_184236466(.A(n_56457), .B(n_28277), .C(n_28471), .D(n_27089
		), .Z(n_342073900));
	notech_and4 i_184836460(.A(n_342073900), .B(n_341973899), .C(n_341773897
		), .D(n_341673896), .Z(n_342273902));
	notech_ao4 i_183936469(.A(n_59344), .B(n_28541), .C(n_28343), .D(n_56371
		), .Z(n_342373903));
	notech_ao4 i_183836470(.A(n_56400), .B(n_28178), .C(n_28407), .D(n_56391
		), .Z(n_342473904));
	notech_and2 i_184036468(.A(n_342473904), .B(n_342373903), .Z(n_342573905
		));
	notech_ao4 i_183636472(.A(n_58014), .B(n_27881), .C(n_56468), .D(n_29944
		), .Z(n_342673906));
	notech_ao4 i_183536473(.A(n_57985), .B(n_28310), .C(n_28504), .D(n_27104
		), .Z(n_342773907));
	notech_ao4 i_157636729(.A(n_276383754), .B(n_29020), .C(n_3888), .D(n_28109
		), .Z(n_343073910));
	notech_ao4 i_157536730(.A(n_310315179), .B(n_56320), .C(n_3887), .D(n_29074
		), .Z(n_343173911));
	notech_ao4 i_157336732(.A(n_54012640), .B(n_29272), .C(n_388360286), .D(nbus_11295
		[20]), .Z(n_343373913));
	notech_and4 i_157836727(.A(n_343373913), .B(n_343173911), .C(n_343073910
		), .D(n_330573785), .Z(n_343573915));
	notech_ao4 i_157036735(.A(n_53412634), .B(n_29634), .C(n_53512635), .D(n_28005
		), .Z(n_343673916));
	notech_ao4 i_156836737(.A(n_3882), .B(n_29237), .C(n_52112621), .D(n_29200
		), .Z(n_343873918));
	notech_and4 i_157236733(.A(n_293087204), .B(n_343873918), .C(n_343673916
		), .D(n_330273782), .Z(n_344073920));
	notech_ao4 i_156536740(.A(n_276383754), .B(n_29019), .C(n_3888), .D(n_28108
		), .Z(n_344173921));
	notech_ao4 i_156436741(.A(n_310315179), .B(n_56311), .C(n_3887), .D(n_29073
		), .Z(n_344273922));
	notech_ao4 i_156236743(.A(n_54012640), .B(n_29271), .C(n_388360286), .D(nbus_11295
		[19]), .Z(n_344473924));
	notech_and4 i_156736738(.A(n_344473924), .B(n_344273922), .C(n_344173921
		), .D(n_329373773), .Z(n_344673926));
	notech_ao4 i_155936746(.A(n_53412634), .B(n_29640), .C(n_53512635), .D(n_28004
		), .Z(n_344773927));
	notech_ao4 i_155736748(.A(n_3882), .B(n_29236), .C(n_52112621), .D(n_29199
		), .Z(n_344973929));
	notech_and4 i_156136744(.A(n_293087204), .B(n_344973929), .C(n_344773927
		), .D(n_329073770), .Z(n_345173931));
	notech_ao4 i_154336762(.A(n_276383754), .B(n_29018), .C(n_3888), .D(n_28106
		), .Z(n_345273932));
	notech_ao4 i_154236763(.A(n_310315179), .B(n_56293), .C(n_3887), .D(n_29070
		), .Z(n_345373933));
	notech_ao4 i_154036765(.A(n_54012640), .B(n_29269), .C(n_388360286), .D(nbus_11295
		[17]), .Z(n_345573935));
	notech_and4 i_154536760(.A(n_345573935), .B(n_345373933), .C(n_345273932
		), .D(n_328173761), .Z(n_345773937));
	notech_ao4 i_153736768(.A(n_53412634), .B(n_29631), .C(n_53512635), .D(n_28002
		), .Z(n_345873938));
	notech_ao4 i_153536770(.A(n_3882), .B(n_29234), .C(n_52112621), .D(n_29197
		), .Z(n_346073940));
	notech_and4 i_153936766(.A(n_346073940), .B(n_345873938), .C(n_277183762
		), .D(n_327873758), .Z(n_346273942));
	notech_nand2 i_318008(.A(n_110371583), .B(n_110271582), .Z(write_data_26
		[2]));
	notech_nand2 i_1818023(.A(n_110571585), .B(n_110471584), .Z(write_data_26
		[17]));
	notech_nand2 i_2018025(.A(n_110771587), .B(n_110671586), .Z(write_data_26
		[19]));
	notech_nand2 i_2118026(.A(n_110971589), .B(n_110871588), .Z(write_data_26
		[20]));
	notech_nao3 i_172467434(.A(n_111171591), .B(n_111071590), .C(n_83341448)
		, .Z(n_346373943));
	notech_and2 i_100564495(.A(n_57299), .B(n_132978833), .Z(n_58044));
	notech_and2 i_150864481(.A(n_57863), .B(n_119171671), .Z(n_57573));
	notech_ao3 i_258164472(.A(n_305391770), .B(n_253162798), .C(n_254240560)
		, .Z(n_56529));
	notech_or4 i_820765(.A(n_121375157), .B(n_122671706), .C(n_125071730), .D
		(n_26628), .Z(n_24472));
	notech_and4 i_321080(.A(n_125771737), .B(n_126471744), .C(n_121871698), 
		.D(n_125671736), .Z(n_18841));
	notech_and4 i_1021631(.A(n_126571745), .B(n_126771747), .C(n_127271752),
		 .D(n_121071690), .Z(n_17834));
	notech_or4 i_821629(.A(n_121375157), .B(n_119371673), .C(n_127771757), .D
		(n_26630), .Z(n_17822));
	notech_or2 i_42661303(.A(n_54894), .B(n_27451), .Z(n_124264771));
	notech_nand3 i_263358500(.A(n_58503), .B(n_58479), .C(n_58495), .Z(n_56482
		));
	notech_or2 i_40461325(.A(n_344966978), .B(n_57644), .Z(n_123764766));
	notech_and2 i_186258511(.A(n_58503), .B(n_58479), .Z(n_57229));
	notech_nand3 i_128461798(.A(n_30945), .B(n_190062172), .C(n_26821), .Z(n_57765
		));
	notech_or4 i_113444509(.A(n_26812), .B(n_57082), .C(n_57055), .D(n_54916
		), .Z(n_57915));
	notech_or2 i_41161318(.A(n_54894), .B(n_27447), .Z(n_123064759));
	notech_and4 i_1621637(.A(n_134471824), .B(n_134671826), .C(n_135171831),
		 .D(n_133871818), .Z(n_17870));
	notech_nand2 i_1421635(.A(n_136071840), .B(n_135671836), .Z(n_17858));
	notech_nand2 i_521786(.A(n_137471854), .B(n_136771847), .Z(n_21008));
	notech_nand2 i_221783(.A(n_138871868), .B(n_138171861), .Z(n_20990));
	notech_nand3 i_131944508(.A(n_56848), .B(n_188562161), .C(n_58498), .Z(n_57730
		));
	notech_or4 i_195358510(.A(n_245362720), .B(n_57087), .C(instrc[116]), .D
		(n_26816), .Z(n_57139));
	notech_nao3 i_62644577(.A(n_32386), .B(n_60349), .C(n_308891735), .Z(n_58391
		));
	notech_nand2 i_1221633(.A(n_144571925), .B(n_144171921), .Z(n_17846));
	notech_and4 i_1121632(.A(n_144671926), .B(n_144871928), .C(n_145371933),
		 .D(n_141771897), .Z(n_17840));
	notech_and4 i_317592(.A(n_146371943), .B(n_146271942), .C(n_146671946), 
		.D(n_146171941), .Z(n_16718));
	notech_and3 i_132055551(.A(n_211359194), .B(n_56848), .C(n_3845), .Z(n_57729
		));
	notech_and2 i_83155600(.A(n_32352), .B(n_56689), .Z(n_58186));
	notech_and3 i_84055599(.A(n_211359194), .B(n_56848), .C(n_26054), .Z(n_58177
		));
	notech_and4 i_85455597(.A(n_56848), .B(n_26054), .C(n_211359194), .D(n_3845
		), .Z(n_58163));
	notech_and2 i_106955590(.A(n_25875), .B(n_146871948), .Z(n_57980));
	notech_or4 i_112755587(.A(n_26062), .B(n_57055), .C(n_29658), .D(n_3853)
		, .Z(n_57922));
	notech_and2 i_193755556(.A(n_57025), .B(n_57731), .Z(n_57154));
	notech_or2 i_195155554(.A(n_58805), .B(n_58486), .Z(n_57141));
	notech_or2 i_39761332(.A(n_54894), .B(n_27445), .Z(n_121364742));
	notech_nao3 i_37661353(.A(opc[9]), .B(n_62822), .C(n_346866997), .Z(n_120864737
		));
	notech_and4 i_142550724(.A(n_181372293), .B(n_181272292), .C(n_180872288
		), .D(n_181172291), .Z(n_59991));
	notech_or4 i_70150717(.A(n_60970), .B(n_60959), .C(n_62848), .D(n_57552)
		, .Z(n_58316));
	notech_nand2 i_37961350(.A(n_7358), .B(n_26986), .Z(n_120564734));
	notech_mux2 i_311672(.S(n_60548), .A(n_5162), .B(add_len_pc32[2]), .Z(add_len_pc
		[2]));
	notech_nand2 i_320696(.A(n_182772307), .B(n_182272302), .Z(n_24768));
	notech_nand2 i_320760(.A(n_183672316), .B(n_183272312), .Z(n_24442));
	notech_or4 i_320856(.A(n_174572225), .B(n_184372323), .C(n_152672006), .D
		(n_26635), .Z(n_24094));
	notech_or4 i_320984(.A(n_152672006), .B(n_173372213), .C(n_185272332), .D
		(n_26637), .Z(n_23746));
	notech_nand2 i_321176(.A(n_186572345), .B(n_186172341), .Z(n_18492));
	notech_nand2 i_2521550(.A(n_187572355), .B(n_187072350), .Z(n_18276));
	notech_nand2 i_2421549(.A(n_188572365), .B(n_188072360), .Z(n_18270));
	notech_nand2 i_2321548(.A(n_189572375), .B(n_189072370), .Z(n_18264));
	notech_and4 i_321624(.A(n_167972159), .B(n_189972379), .C(n_190572385), 
		.D(n_189872378), .Z(n_17792));
	notech_nand2 i_2521806(.A(n_191672396), .B(n_191172391), .Z(n_21128));
	notech_nand2 i_2421805(.A(n_192772407), .B(n_192272402), .Z(n_21122));
	notech_nand2 i_2321804(.A(n_193872418), .B(n_193372413), .Z(n_21116));
	notech_nand2 i_321784(.A(n_195472434), .B(n_194872428), .Z(n_20996));
	notech_and4 i_321848(.A(n_196172441), .B(n_196072440), .C(n_160672086), 
		.D(n_196472444), .Z(n_20630));
	notech_and4 i_2521934(.A(n_197172451), .B(n_197372453), .C(n_197072450),
		 .D(n_159672076), .Z(n_17576));
	notech_and4 i_2421933(.A(n_197972459), .B(n_198172461), .C(n_158872068),
		 .D(n_197872458), .Z(n_17570));
	notech_and4 i_2321932(.A(n_198872468), .B(n_199072470), .C(n_198772467),
		 .D(n_157872058), .Z(n_17564));
	notech_and4 i_2517038(.A(n_199772477), .B(n_199972479), .C(n_199672476),
		 .D(n_156972049), .Z(n_17219));
	notech_and4 i_2417037(.A(n_200672486), .B(n_200872488), .C(n_200572485),
		 .D(n_155872038), .Z(n_17213));
	notech_nand3 i_12255(.A(n_60358), .B(n_60162), .C(n_114164670), .Z(n_120264731
		));
	notech_nand3 i_4744447(.A(n_58481), .B(n_58505), .C(n_58497), .Z(n_58167
		));
	notech_or2 i_36261367(.A(n_58367), .B(n_27990), .Z(n_119564724));
	notech_mux2 i_1911688(.S(n_60548), .A(regs_14[18]), .B(add_len_pc32[18])
		, .Z(add_len_pc[18]));
	notech_and4 i_144047710(.A(n_246772947), .B(n_246672946), .C(n_246272942
		), .D(n_246572945), .Z(n_313647722));
	notech_and4 i_144247708(.A(n_244272922), .B(n_244172921), .C(n_243772917
		), .D(n_244072920), .Z(n_313447724));
	notech_and4 i_144347707(.A(n_242772907), .B(n_242672906), .C(n_242272902
		), .D(n_242572905), .Z(n_313347725));
	notech_nand2 i_1920712(.A(n_245472934), .B(n_244972929), .Z(n_24864));
	notech_and4 i_2120778(.A(n_247172951), .B(n_247372953), .C(n_247872958),
		 .D(n_235272832), .Z(n_24550));
	notech_and4 i_2020777(.A(n_248072960), .B(n_248272962), .C(n_248772967),
		 .D(n_234372823), .Z(n_24544));
	notech_and4 i_1920776(.A(n_248872968), .B(n_249072970), .C(n_249572975),
		 .D(n_233472814), .Z(n_24538));
	notech_and4 i_1820775(.A(n_249772977), .B(n_249972979), .C(n_250472984),
		 .D(n_232572805), .Z(n_24532));
	notech_or4 i_2120874(.A(n_287569887), .B(n_230972789), .C(n_250872988), 
		.D(n_26652), .Z(n_24202));
	notech_or4 i_2020873(.A(n_287969891), .B(n_230172781), .C(n_251572995), 
		.D(n_26653), .Z(n_24196));
	notech_or4 i_1920872(.A(n_288369895), .B(n_229372773), .C(n_252273002), 
		.D(n_26654), .Z(n_24190));
	notech_and4 i_2121002(.A(n_252673006), .B(n_252873008), .C(n_229272772),
		 .D(n_253273012), .Z(n_23854));
	notech_and4 i_2021001(.A(n_253373013), .B(n_253573015), .C(n_254173021),
		 .D(n_228472764), .Z(n_23848));
	notech_and4 i_1820999(.A(n_227572755), .B(n_254273022), .C(n_254473024),
		 .D(n_255073030), .Z(n_23836));
	notech_or4 i_1821095(.A(n_288769899), .B(n_225772737), .C(n_255773037), 
		.D(n_26655), .Z(n_18931));
	notech_or4 i_2121194(.A(n_287569887), .B(n_224972729), .C(n_256373043), 
		.D(n_26656), .Z(n_18600));
	notech_and4 i_2021193(.A(n_256773047), .B(n_256973049), .C(n_224872728),
		 .D(n_257473054), .Z(n_18594));
	notech_and4 i_1821191(.A(n_257573055), .B(n_257773057), .C(n_223972719),
		 .D(n_258273062), .Z(n_18582));
	notech_nand2 i_2121546(.A(n_259273072), .B(n_258773067), .Z(n_18252));
	notech_nand2 i_2021545(.A(n_260373083), .B(n_259873078), .Z(n_18246));
	notech_nand2 i_1921544(.A(n_261473094), .B(n_260973089), .Z(n_18240));
	notech_nand2 i_1821543(.A(n_262573105), .B(n_262073100), .Z(n_18234));
	notech_or4 i_2121642(.A(n_287569887), .B(n_217272652), .C(n_262973109), 
		.D(n_26657), .Z(n_17900));
	notech_and4 i_2021641(.A(n_263373113), .B(n_263573115), .C(n_217172651),
		 .D(n_264073120), .Z(n_17894));
	notech_and4 i_1921640(.A(n_264173121), .B(n_264373123), .C(n_216272642),
		 .D(n_264873128), .Z(n_17888));
	notech_and4 i_1821639(.A(n_264973129), .B(n_265173131), .C(n_215372633),
		 .D(n_265673136), .Z(n_17882));
	notech_or4 i_2121866(.A(n_287569887), .B(n_213772617), .C(n_266073140), 
		.D(n_26658), .Z(n_20738));
	notech_nand2 i_2021865(.A(n_267273152), .B(n_266873148), .Z(n_20732));
	notech_nand2 i_1821863(.A(n_268173161), .B(n_267773157), .Z(n_20720));
	notech_and4 i_2121930(.A(n_268673166), .B(n_268873168), .C(n_211372593),
		 .D(n_268573165), .Z(n_17552));
	notech_and4 i_2021929(.A(n_269573175), .B(n_269773177), .C(n_269473174),
		 .D(n_210372583), .Z(n_17546));
	notech_nand2 i_1921928(.A(n_270873188), .B(n_270373183), .Z(n_17540));
	notech_and4 i_1821927(.A(n_271473194), .B(n_271673196), .C(n_271373193),
		 .D(n_208372563), .Z(n_17534));
	notech_and4 i_2117034(.A(n_272373203), .B(n_272573205), .C(n_272273202),
		 .D(n_207372553), .Z(n_17195));
	notech_nand2 i_2017033(.A(n_273673216), .B(n_273173211), .Z(n_17189));
	notech_nand2 i_1817031(.A(n_274673226), .B(n_274173221), .Z(n_17177));
	notech_or4 i_2117610(.A(n_203572515), .B(n_287569887), .C(n_275373233), 
		.D(n_26659), .Z(n_16826));
	notech_nand2 i_2017609(.A(n_276573245), .B(n_276073240), .Z(n_16820));
	notech_nand2 i_1817607(.A(n_277573255), .B(n_277073250), .Z(n_16808));
	notech_nand2 i_5347646(.A(n_26707), .B(n_27179), .Z(n_306024324));
	notech_ao4 i_191847740(.A(n_30821), .B(n_60246), .C(n_311991704), .D(n_315191672
		), .Z(n_57173));
	notech_nao3 i_36961360(.A(n_319391630), .B(temp_sp[7]), .C(n_27552), .Z(n_118864717
		));
	notech_or2 i_26961459(.A(n_57173), .B(\nbus_11365[21] ), .Z(n_118564714)
		);
	notech_or2 i_27261456(.A(n_149228769), .B(n_29681), .Z(n_118264711));
	notech_or4 i_27561453(.A(n_311991704), .B(n_26939), .C(nbus_11295[21]), 
		.D(n_60949), .Z(n_117964708));
	notech_nao3 i_7761651(.A(opa[21]), .B(n_26707), .C(n_319891625), .Z(n_117564704
		));
	notech_nand2 i_8061648(.A(\regs_13_14[21] ), .B(n_151328790), .Z(n_117264701
		));
	notech_or4 i_8361645(.A(n_316491659), .B(n_26942), .C(nbus_11295[21]), .D
		(n_60949), .Z(n_116964698));
	notech_nand2 i_97144544(.A(n_32348), .B(n_58186), .Z(n_58078));
	notech_mux2 i_411673(.S(n_60548), .A(n_5163), .B(add_len_pc32[3]), .Z(add_len_pc
		[3]));
	notech_mux2 i_611675(.S(n_60548), .A(n_5165), .B(add_len_pc32[5]), .Z(add_len_pc
		[5]));
	notech_mux2 i_711676(.S(n_60548), .A(n_5166), .B(add_len_pc32[6]), .Z(add_len_pc
		[6]));
	notech_mux2 i_811677(.S(n_60548), .A(n_5167), .B(add_len_pc32[7]), .Z(add_len_pc
		[7]));
	notech_or4 i_73244522(.A(n_60970), .B(n_60959), .C(n_62860), .D(\nbus_11307[7] 
		), .Z(n_58285));
	notech_or2 i_121560576(.A(n_268666215), .B(n_300591818), .Z(n_116264691)
		);
	notech_or4 i_48744518(.A(fsm[2]), .B(n_61165), .C(n_61154), .D(n_27306),
		 .Z(n_58530));
	notech_nao3 i_121460577(.A(n_281666345), .B(n_32334), .C(n_2351), .Z(n_116164690
		));
	notech_nao3 i_112644513(.A(n_30945), .B(n_190062172), .C(n_58489), .Z(n_57923
		));
	notech_nand2 i_820701(.A(n_305873538), .B(n_305273532), .Z(n_24798));
	notech_nand2 i_720700(.A(n_307273552), .B(n_306773547), .Z(n_24792));
	notech_nand2 i_620699(.A(n_308573565), .B(n_307973559), .Z(n_24786));
	notech_nand2 i_420697(.A(n_309873578), .B(n_309273572), .Z(n_24774));
	notech_nand2 i_720764(.A(n_311373593), .B(n_310673586), .Z(n_24466));
	notech_or4 i_820861(.A(n_121375157), .B(n_295073430), .C(n_311973599), .D
		(n_26660), .Z(n_24124));
	notech_and4 i_720860(.A(n_311173591), .B(n_312973609), .C(n_293873418), 
		.D(n_312873608), .Z(n_24118));
	notech_nand3 i_820989(.A(n_313673616), .B(n_313573615), .C(n_314073620),
		 .Z(n_23776));
	notech_and4 i_720988(.A(n_311173591), .B(n_314773627), .C(n_291573395), 
		.D(n_314673626), .Z(n_23770));
	notech_nand2 i_821085(.A(n_315973639), .B(n_315473634), .Z(n_18871));
	notech_nand2 i_721084(.A(n_317073650), .B(n_316573645), .Z(n_18865));
	notech_or4 i_821181(.A(n_121375157), .B(n_288073360), .C(n_317873658), .D
		(n_26661), .Z(n_18522));
	notech_and4 i_721180(.A(n_311173591), .B(n_318673666), .C(n_287073350), 
		.D(n_318573665), .Z(n_18516));
	notech_nand2 i_621371(.A(n_319873678), .B(n_319373673), .Z(n_25276));
	notech_nand2 i_421369(.A(n_320873688), .B(n_320373683), .Z(n_25264));
	notech_nand2 i_421785(.A(n_322273702), .B(n_321573695), .Z(n_21002));
	notech_and2 i_344474(.A(n_92619108), .B(n_277673256), .Z(n_305721221));
	notech_ao4 i_2044473(.A(n_59435), .B(n_29723), .C(n_60868), .D(n_3874), 
		.Z(n_305621220));
	notech_or4 i_120060591(.A(calc_sz[1]), .B(n_246691943), .C(n_26602), .D(n_60010
		), .Z(n_115964688));
	notech_and2 i_100941360(.A(n_58084), .B(n_322773707), .Z(n_58040));
	notech_and2 i_99541359(.A(n_57875), .B(n_58194), .Z(n_58054));
	notech_ao4 i_99441358(.A(n_59445), .B(n_26811), .C(n_58173), .D(n_26916)
		, .Z(n_58055));
	notech_nand2 i_63941357(.A(n_58429), .B(n_322673706), .Z(n_58378));
	notech_mux2 i_211671(.S(n_60548), .A(n_5161), .B(add_len_pc32[1]), .Z(add_len_pc
		[1]));
	notech_nand2 i_220695(.A(n_326573745), .B(n_325973739), .Z(n_24762));
	notech_and4 i_921630(.A(n_323673716), .B(n_326673746), .C(n_326873748), 
		.D(n_327373753), .Z(n_17828));
	notech_nand3 i_84360913(.A(n_60162), .B(n_60246), .C(read_data[15]), .Z(n_115264681
		));
	notech_and4 i_91338309(.A(n_338573865), .B(n_338473864), .C(n_338073860)
		, .D(n_338373863), .Z(n_60023));
	notech_and4 i_92838283(.A(n_339973879), .B(n_339873878), .C(n_339473874)
		, .D(n_339773877), .Z(n_60008));
	notech_and4 i_93038281(.A(n_341373893), .B(n_341273892), .C(n_340873888)
		, .D(n_341173891), .Z(n_60006));
	notech_and4 i_93138280(.A(n_342773907), .B(n_342673906), .C(n_342273902)
		, .D(n_342573905), .Z(n_60005));
	notech_nand2 i_2116234(.A(n_344073920), .B(n_343573915), .Z(n_19226));
	notech_nand2 i_2016233(.A(n_345173931), .B(n_344673926), .Z(n_19220));
	notech_nand2 i_1816231(.A(n_346273942), .B(n_345773937), .Z(n_19208));
	notech_and2 i_84260914(.A(n_27302), .B(\opa_12[15] ), .Z(n_115164680));
	notech_nand3 i_82960927(.A(n_60162), .B(n_60246), .C(read_data[14]), .Z(n_114764676
		));
	notech_nand3 i_81460941(.A(n_60162), .B(n_60246), .C(read_data[13]), .Z(n_114664675
		));
	notech_and3 i_4261686(.A(n_32355), .B(n_32370), .C(n_32351), .Z(n_114464673
		));
	notech_nand2 i_4361685(.A(n_1476), .B(opb[9]), .Z(n_114264671));
	notech_nand3 i_78160973(.A(n_200165530), .B(n_200265531), .C(n_114264671
		), .Z(n_114164670));
	notech_nand3 i_78060974(.A(n_60162), .B(n_60241), .C(read_data[9]), .Z(n_114064669
		));
	notech_nand2 i_77960975(.A(n_27302), .B(\opa_12[9] ), .Z(n_113964668));
	notech_ao4 i_115261756(.A(n_59968), .B(n_32347), .C(n_27992), .D(n_114464673
		), .Z(n_113864667));
	notech_and2 i_1361711(.A(n_58608), .B(n_113964668), .Z(n_113764666));
	notech_nand2 i_1161712(.A(n_300991814), .B(n_300391820), .Z(n_113664665)
		);
	notech_ao4 i_1061713(.A(n_59445), .B(n_27302), .C(n_28542), .D(n_26748),
		 .Z(n_113564664));
	notech_and3 i_1461710(.A(n_28544), .B(n_28543), .C(n_301091813), .Z(n_113464663
		));
	notech_nand2 i_63461109(.A(n_27304), .B(\opa_12[15] ), .Z(n_113364662)
		);
	notech_and2 i_1761707(.A(n_58622), .B(n_113364662), .Z(n_113264661));
	notech_nand2 i_56161171(.A(n_27304), .B(\opa_12[9] ), .Z(n_113164660));
	notech_nand2 i_2361702(.A(n_300791816), .B(n_313791686), .Z(n_113064659)
		);
	notech_nand2 i_2261703(.A(n_313891685), .B(n_315091673), .Z(n_112964658)
		);
	notech_and2 i_2061704(.A(n_58608), .B(n_113164660), .Z(n_112864657));
	notech_and2 i_2561700(.A(n_313791686), .B(n_174165270), .Z(n_112664655)
		);
	notech_ao4 i_2461701(.A(n_59445), .B(n_27304), .C(n_27163), .D(n_26591),
		 .Z(n_112564654));
	notech_ao4 i_2861697(.A(n_59434), .B(n_29754), .C(n_26611), .D(n_60010),
		 .Z(n_112364652));
	notech_ao4 i_3161694(.A(n_26611), .B(n_60016), .C(n_59434), .D(n_29743),
		 .Z(n_112164650));
	notech_and3 i_3061695(.A(n_312991694), .B(n_116164690), .C(n_347066999),
		 .Z(n_112064649));
	notech_and2 i_2961696(.A(n_346966998), .B(n_344566974), .Z(n_111964648)
		);
	notech_and4 i_3361692(.A(n_312991694), .B(n_28222), .C(n_116164690), .D(n_312791696
		), .Z(n_111864647));
	notech_and3 i_3261693(.A(n_298991830), .B(n_344566974), .C(n_312891695),
		 .Z(n_111764646));
	notech_nand2 i_151961749(.A(n_26890), .B(n_27280), .Z(n_111664645));
	notech_or4 i_140761750(.A(n_59387), .B(n_246891941), .C(n_32355), .D(instrc
		[115]), .Z(n_111564644));
	notech_or4 i_135961751(.A(n_56512), .B(n_57087), .C(instrc[116]), .D(n_54916
		), .Z(n_111464643));
	notech_ao4 i_114461758(.A(n_102135817), .B(n_302091803), .C(n_102035816)
		, .D(n_29592), .Z(n_111364642));
	notech_nao3 i_67761768(.A(n_155265081), .B(n_155465083), .C(n_154765076)
		, .Z(n_111264641));
	notech_or4 i_31061777(.A(n_60970), .B(n_60959), .C(n_62848), .D(n_57733)
		, .Z(n_111164640));
	notech_nand2 i_3961779(.A(opc[15]), .B(n_62794), .Z(n_111064639));
	notech_nand2 i_2161781(.A(opc_10[21]), .B(n_62822), .Z(n_110964638));
	notech_ao4 i_155062947(.A(n_323180732), .B(n_29743), .C(n_57473), .D(n_291963186
		), .Z(n_110664635));
	notech_and3 i_155562942(.A(n_110264631), .B(n_110464633), .C(n_110164630
		), .Z(n_110564634));
	notech_ao4 i_155262945(.A(n_26823), .B(nbus_11295[9]), .C(n_58480), .D(n_58608
		), .Z(n_110464633));
	notech_ao4 i_155362944(.A(n_250240520), .B(\nbus_11358[9] ), .C(n_26846)
		, .D(\nbus_11307[9] ), .Z(n_110264631));
	notech_or2 i_83263643(.A(n_56636), .B(n_252740545), .Z(n_110164630));
	notech_or2 i_83763638(.A(n_57299), .B(n_60016), .Z(n_109464623));
	notech_or2 i_83863637(.A(n_32356), .B(n_27992), .Z(n_109364622));
	notech_ao4 i_129768565(.A(n_326790765), .B(n_27751), .C(n_326890766), .D
		(n_27792), .Z(n_109264621));
	notech_ao4 i_129868564(.A(n_326990767), .B(n_60004), .C(n_56391), .D(n_27465
		), .Z(n_109164620));
	notech_and4 i_34083472(.A(n_327063487), .B(n_328163498), .C(n_22995), .D
		(n_22035), .Z(n_331163528));
	notech_nand3 i_35731(.A(n_59259), .B(n_27983), .C(n_27985), .Z(n_330963526
		));
	notech_nand2 i_35730(.A(n_59259), .B(n_27983), .Z(n_330863525));
	notech_nand2 i_12083471(.A(over_seg[5]), .B(n_60548), .Z(n_58812));
	notech_or4 i_34246(.A(fsm[2]), .B(n_61165), .C(n_61154), .D(n_60893), .Z
		(n_330763524));
	notech_nao3 i_25283469(.A(over_seg[5]), .B(n_60548), .C(n_326591251), .Z
		(n_330563522));
	notech_or4 i_3423(.A(n_27925), .B(n_60868), .C(n_32747), .D(\opcode[3] )
		, .Z(n_330463521));
	notech_nao3 i_14832593(.A(fsm[2]), .B(n_32562), .C(n_61165), .Z(n_17189930
		));
	notech_nand2 i_12632615(.A(n_27378), .B(n_314863415), .Z(n_17409952));
	notech_or4 i_11332628(.A(n_32270), .B(n_26900), .C(n_60373), .D(n_1862),
		 .Z(n_17539965));
	notech_or4 i_8732652(.A(n_61115), .B(n_315291671), .C(n_62848), .D(n_62822
		), .Z(n_17779989));
	notech_and4 i_226951(.A(n_324891268), .B(n_324791269), .C(n_325791259), 
		.D(n_325191265), .Z(n_19653));
	notech_nand2 i_9850(.A(n_314963416), .B(n_61110), .Z(n_14843));
	notech_nand3 i_9840(.A(n_317963446), .B(n_61110), .C(n_317863445), .Z(n_21585
		));
	notech_or4 i_35332738(.A(n_32566), .B(n_26580), .C(n_32403), .D(n_19036)
		, .Z(n_58664));
	notech_or2 i_180632739(.A(n_320063467), .B(n_26761), .Z(n_57285));
	notech_and2 i_23132740(.A(n_324263481), .B(n_23006), .Z(n_58786));
	notech_or4 i_9832641(.A(n_61145), .B(n_60358), .C(n_26900), .D(n_60373),
		 .Z(n_17669978));
	notech_or4 i_32119(.A(n_60970), .B(n_60959), .C(n_62848), .D(n_60241), .Z
		(n_190710119));
	notech_or4 i_3434(.A(n_4958709), .B(n_32695), .C(n_32747), .D(n_2838), .Z
		(n_60054));
	notech_nand2 i_5949(.A(sema_rw), .B(n_320391620), .Z(n_53739));
	notech_or4 i_35532862(.A(n_32580), .B(n_61145), .C(n_29655), .D(n_27065)
		, .Z(n_58662));
	notech_or2 i_5962(.A(n_266891921), .B(n_32476), .Z(n_53731));
	notech_or4 i_3068(.A(n_60970), .B(n_60959), .C(n_319691627), .D(n_62848)
		, .Z(n_60074));
	notech_nao3 i_52253(.A(n_60162), .B(n_60358), .C(n_60054), .Z(n_60136)
		);
	notech_or2 i_8160(.A(n_315963426), .B(n_29793), .Z(n_51771));
	notech_nand2 i_56532(.A(n_51771), .B(n_60129), .Z(\nbus_11380[0] ));
	notech_nand2 i_56533(.A(n_61560), .B(n_316263429), .Z(n_60129));
	notech_or4 i_5735053(.A(n_60970), .B(n_60959), .C(n_60909), .D(n_60241),
		 .Z(n_303747815));
	notech_or4 i_3485(.A(n_62868), .B(n_62892), .C(n_27573), .D(n_59434), .Z
		(n_60051));
	notech_nand2 i_3138203(.A(n_28049), .B(n_28050), .Z(n_307215148));
	notech_and4 i_91538296(.A(n_312763394), .B(n_312663393), .C(n_312263389)
		, .D(n_312563392), .Z(n_5743));
	notech_nand3 i_9271(.A(n_28049), .B(n_28050), .C(opz[2]), .Z(n_50662));
	notech_or4 i_98041270(.A(opc[3]), .B(opc[2]), .C(opc[1]), .D(opc[0]), .Z
		(n_291118110));
	notech_nand2 i_97641271(.A(opc[1]), .B(opc[0]), .Z(n_291218111));
	notech_nand2 i_90341273(.A(nbus_11295[1]), .B(nbus_11295[0]), .Z(n_291418113
		));
	notech_nand2 i_917022(.A(n_305163318), .B(n_304663313), .Z(n_17123));
	notech_and4 i_921022(.A(n_289363160), .B(n_303363300), .C(n_303563302), 
		.D(n_304063307), .Z(n_14022));
	notech_nand2 i_520698(.A(n_303263299), .B(n_302663293), .Z(n_24780));
	notech_nand3 i_108441265(.A(opc[1]), .B(opc[0]), .C(opc[2]), .Z(n_290618105
		));
	notech_or4 i_40941308(.A(n_60969), .B(n_60958), .C(n_62848), .D(n_29743)
		, .Z(n_58608));
	notech_mux2 i_511674(.S(n_60548), .A(n_5164), .B(add_len_pc32[4]), .Z(add_len_pc
		[4]));
	notech_and3 i_61141321(.A(n_315591668), .B(n_318691637), .C(n_121628493)
		, .Z(n_58406));
	notech_and4 i_142741322(.A(n_300263269), .B(n_300163268), .C(n_299763264
		), .D(n_300063267), .Z(n_5723));
	notech_and3 i_257741323(.A(n_316591658), .B(n_32350), .C(n_316891655), .Z
		(n_56533));
	notech_and3 i_96841324(.A(n_309091733), .B(n_316791656), .C(n_318191642)
		, .Z(n_58081));
	notech_nand2 i_167941387(.A(rep_en2), .B(n_27378), .Z(n_57406));
	notech_or4 i_115341393(.A(n_291418113), .B(opc[3]), .C(opc[2]), .D(opc[4
		]), .Z(n_57896));
	notech_or4 i_34241402(.A(rep_en1), .B(rep_en3), .C(rep_en2), .D(rep_en4)
		, .Z(n_58675));
	notech_or4 i_32041403(.A(rep_en1), .B(rep_en3), .C(rep_en2), .D(n_27380)
		, .Z(n_58697));
	notech_or2 i_10244392(.A(n_58133), .B(n_32322), .Z(n_295921141));
	notech_ao4 i_4044454(.A(n_58133), .B(n_32322), .C(n_59419), .D(n_26753),
		 .Z(n_58421));
	notech_nand2 i_421017(.A(n_285263119), .B(n_284763114), .Z(n_13992));
	notech_nand2 i_621019(.A(n_284263109), .B(n_283763104), .Z(n_14004));
	notech_nand2 i_721020(.A(n_283263099), .B(n_282863095), .Z(n_14010));
	notech_or4 i_3221045(.A(n_215876097), .B(n_280463071), .C(n_281963086), 
		.D(n_26842), .Z(n_14160));
	notech_ao4 i_51244512(.A(n_56859), .B(n_26962), .C(n_32352), .D(n_32292)
		, .Z(n_58505));
	notech_ao4 i_52844514(.A(n_56858), .B(n_26610), .C(n_32356), .D(n_32292)
		, .Z(n_58489));
	notech_or4 i_69244516(.A(instrc[122]), .B(n_58133), .C(instrc[121]), .D(n_26735
		), .Z(n_58325));
	notech_or4 i_12244517(.A(n_57026), .B(n_57087), .C(instrc[116]), .D(n_29653
		), .Z(n_58810));
	notech_nand2 i_30402(.A(n_26763), .B(n_26945), .Z(n_309721261));
	notech_and3 i_115944563(.A(n_28222), .B(n_274663013), .C(n_188857101), .Z
		(n_57890));
	notech_and2 i_116044564(.A(n_298991830), .B(n_276363030), .Z(n_57889));
	notech_ao4 i_88444569(.A(n_60893), .B(n_26753), .C(n_62822), .D(n_60909)
		, .Z(n_58133));
	notech_ao4 i_52044579(.A(n_56859), .B(n_56935), .C(n_56689), .D(n_32292)
		, .Z(n_58497));
	notech_nao3 i_82544585(.A(n_58172), .B(n_32322), .C(n_58133), .Z(n_58192
		));
	notech_and2 i_158344535(.A(n_59434), .B(n_58421), .Z(n_57500));
	notech_ao4 i_53644590(.A(n_56859), .B(n_32382), .C(n_32348), .D(n_32292)
		, .Z(n_58481));
	notech_nand3 i_84641340(.A(n_56848), .B(n_125961542), .C(n_26804), .Z(n_58171
		));
	notech_nand2 i_158241388(.A(n_59434), .B(n_58422), .Z(n_57501));
	notech_and4 i_1721030(.A(n_273963006), .B(n_274163008), .C(n_274563012),
		 .D(n_254362810), .Z(n_14070));
	notech_and4 i_1821031(.A(n_273563002), .B(n_273763004), .C(n_254762814),
		 .D(n_273463001), .Z(n_14076));
	notech_and4 i_1921032(.A(n_272762994), .B(n_272962996), .C(n_255662823),
		 .D(n_272662993), .Z(n_14082));
	notech_and4 i_2021033(.A(n_271962986), .B(n_272162988), .C(n_256562832),
		 .D(n_271862985), .Z(n_14088));
	notech_nand3 i_2121034(.A(n_271362980), .B(n_271262979), .C(n_271162978)
		, .Z(n_14094));
	notech_and4 i_2221035(.A(n_258262849), .B(n_270462971), .C(n_270662973),
		 .D(n_270362970), .Z(n_14100));
	notech_nand2 i_1720710(.A(n_269962966), .B(n_269462961), .Z(n_24852));
	notech_nand2 i_1820711(.A(n_268962956), .B(n_268462951), .Z(n_24858));
	notech_nand2 i_2020713(.A(n_267962946), .B(n_267462941), .Z(n_24870));
	notech_nand2 i_2120714(.A(n_266962936), .B(n_266462931), .Z(n_24876));
	notech_nand2 i_2220715(.A(n_265962926), .B(n_265462921), .Z(n_24882));
	notech_or4 i_125047719(.A(n_26062), .B(n_57087), .C(n_57055), .D(n_24589
		), .Z(n_57799));
	notech_mux2 i_2211691(.S(n_60548), .A(regs_14[21]), .B(add_len_pc32[21])
		, .Z(add_len_pc[21]));
	notech_mux2 i_2111690(.S(n_60548), .A(regs_14[20]), .B(add_len_pc32[20])
		, .Z(add_len_pc[20]));
	notech_mux2 i_2011689(.S(n_60548), .A(regs_14[19]), .B(add_len_pc32[19])
		, .Z(add_len_pc[19]));
	notech_mux2 i_1811687(.S(n_60548), .A(regs_14[17]), .B(add_len_pc32[17])
		, .Z(add_len_pc[17]));
	notech_mux2 i_1711686(.S(n_60548), .A(regs_14[16]), .B(add_len_pc32[16])
		, .Z(add_len_pc[16]));
	notech_and2 i_199241380(.A(n_59434), .B(n_57926), .Z(n_57100));
	notech_or4 i_120847744(.A(n_26062), .B(n_24583), .C(n_57087), .D(n_57055
		), .Z(n_57841));
	notech_or4 i_201647746(.A(n_245362720), .B(n_57088), .C(n_57055), .D(n_60949
		), .Z(n_57076));
	notech_nao3 i_179247754(.A(n_32338), .B(n_26731), .C(n_58480), .Z(n_57299
		));
	notech_ao4 i_157647759(.A(n_32338), .B(n_58087), .C(n_59419), .D(n_58815
		), .Z(n_57505));
	notech_or4 i_179347767(.A(n_30854), .B(n_245362720), .C(n_60949), .D(n_58488
		), .Z(n_57298));
	notech_ao4 i_52147769(.A(n_56859), .B(n_56935), .C(n_56688), .D(n_32298)
		, .Z(n_58496));
	notech_nand3 i_14798(.A(n_32338), .B(n_26731), .C(n_26599), .Z(n_45139)
		);
	notech_nand3 i_161547774(.A(n_32338), .B(n_26731), .C(n_26808), .Z(n_57470
		));
	notech_nand3 i_82741395(.A(n_58171), .B(n_32325), .C(n_26790), .Z(n_58190
		));
	notech_ao4 i_53747779(.A(n_56858), .B(n_32382), .C(n_32348), .D(n_32298)
		, .Z(n_58480));
	notech_ao4 i_52947780(.A(n_56858), .B(n_26610), .C(n_32356), .D(n_32298)
		, .Z(n_58488));
	notech_ao4 i_51347781(.A(n_56858), .B(n_26962), .C(n_32352), .D(n_32298)
		, .Z(n_58504));
	notech_ao4 i_96247753(.A(n_60893), .B(n_58815), .C(n_62792), .D(n_60909)
		, .Z(n_58087));
	notech_nand2 i_44447782(.A(n_32338), .B(n_26731), .Z(n_58573));
	notech_nand2 i_38547783(.A(n_59434), .B(n_57505), .Z(n_58632));
	notech_nand2 i_321016(.A(n_250462771), .B(n_250062767), .Z(n_13986));
	notech_nand3 i_2321036(.A(n_249362760), .B(n_249262759), .C(n_249162758)
		, .Z(n_14106));
	notech_nand3 i_2421037(.A(n_248662753), .B(n_248562752), .C(n_248462751)
		, .Z(n_14112));
	notech_nand3 i_2521038(.A(n_247962746), .B(n_247862745), .C(n_247762744)
		, .Z(n_14118));
	notech_nand3 i_2621039(.A(n_247262739), .B(n_247162738), .C(n_247062737)
		, .Z(n_14124));
	notech_ao4 i_51450681(.A(n_56858), .B(n_26962), .C(n_32352), .D(n_32304)
		, .Z(n_58503));
	notech_or4 i_25905(.A(n_246362730), .B(n_245962726), .C(n_245662723), .D
		(n_246562732), .Z(n_288827270));
	notech_or2 i_184250682(.A(n_58100), .B(n_56448), .Z(n_57249));
	notech_or2 i_155050707(.A(n_288827270), .B(n_27052), .Z(n_5380));
	notech_nao3 i_264450692(.A(n_58503), .B(n_27024), .C(n_240762674), .Z(n_56471
		));
	notech_ao4 i_94950704(.A(n_60893), .B(n_26769), .C(n_62822), .D(n_60909)
		, .Z(n_58100));
	notech_ao4 i_156750706(.A(n_246791942), .B(n_2479), .C(n_59344), .D(n_29734
		), .Z(n_57514));
	notech_nand2 i_209850709(.A(n_59434), .B(n_57927), .Z(n_56994));
	notech_or2 i_177550705(.A(n_58100), .B(n_32332), .Z(n_57316));
	notech_ao4 i_112250711(.A(n_58100), .B(n_32332), .C(n_59419), .D(n_26769
		), .Z(n_57927));
	notech_ao4 i_53850720(.A(n_56858), .B(n_32382), .C(n_32348), .D(n_32304)
		, .Z(n_58479));
	notech_or2 i_53050721(.A(n_240762674), .B(n_305291771), .Z(n_58487));
	notech_ao4 i_52250722(.A(n_56859), .B(n_56935), .C(n_56684), .D(n_32304)
		, .Z(n_58495));
	notech_nand2 i_206371079(.A(n_60241), .B(read_data[27]), .Z(n_57029));
	notech_and3 i_87947773(.A(n_57299), .B(n_57470), .C(n_45139), .Z(n_58138
		));
	notech_and2 i_132347766(.A(n_57298), .B(n_252762794), .Z(n_57726));
	notech_ao4 i_151247760(.A(n_59445), .B(n_26829), .C(n_26808), .D(n_252662793
		), .Z(n_57569));
	notech_and2 i_87850715(.A(n_228579786), .B(n_240362670), .Z(n_58139));
	notech_and2 i_87647775(.A(n_57025), .B(n_252962796), .Z(n_58141));
	notech_ao4 i_87347777(.A(n_59445), .B(n_26824), .C(n_58171), .D(n_26825)
		, .Z(n_58144));
	notech_and2 i_87447776(.A(n_58190), .B(n_228479785), .Z(n_58143));
	notech_ao4 i_87144536(.A(n_59445), .B(n_26813), .C(n_58172), .D(n_26821)
		, .Z(n_58146));
	notech_and2 i_87244537(.A(n_181779321), .B(n_58192), .Z(n_58145));
	notech_and3 i_11938270(.A(n_28049), .B(n_28050), .C(n_28051), .Z(n_58813
		));
	notech_or2 i_96744510(.A(n_58810), .B(n_58497), .Z(n_58082));
	notech_or4 i_117644515(.A(n_32326), .B(n_58133), .C(n_26735), .D(n_58497
		), .Z(n_57873));
	notech_or2 i_118044511(.A(n_57500), .B(n_58497), .Z(n_57869));
	notech_or4 i_96444581(.A(n_57026), .B(n_30854), .C(n_29653), .D(n_58493)
		, .Z(n_58085));
	notech_or4 i_5247647(.A(n_57026), .B(n_30854), .C(n_29653), .D(n_250662773
		), .Z(n_306124325));
	notech_nand3 i_5447645(.A(n_319191632), .B(n_318791636), .C(n_57988), .Z
		(n_305924323));
	notech_nao3 i_59044589(.A(n_319191632), .B(n_318791636), .C(n_56684), .Z
		(n_58427));
	notech_nand2 i_117941391(.A(n_57501), .B(n_26800), .Z(n_57870));
	notech_or2 i_4247657(.A(n_58805), .B(n_58494), .Z(n_307124335));
	notech_or2 i_4747652(.A(n_58805), .B(n_250562772), .Z(n_306624330));
	notech_nand3 i_4547654(.A(n_319191632), .B(n_57988), .C(n_319091633), .Z
		(n_306824332));
	notech_nao3 i_59244588(.A(n_319191632), .B(n_319091633), .C(n_56684), .Z
		(n_58425));
	notech_or2 i_4047659(.A(n_57100), .B(n_250562772), .Z(n_307324337));
	notech_or2 i_30060(.A(n_58494), .B(n_57100), .Z(n_314047718));
	notech_or4 i_107350654(.A(n_245362720), .B(n_57088), .C(instrc[116]), .D
		(n_58495), .Z(n_286927251));
	notech_or4 i_107650653(.A(n_245362720), .B(n_57088), .C(instrc[116]), .D
		(n_240162668), .Z(n_286827250));
	notech_nao3 i_55850663(.A(n_318891635), .B(n_57988), .C(n_246891941), .Z
		(n_287827260));
	notech_or4 i_59350718(.A(n_59387), .B(n_246891941), .C(n_56684), .D(n_29178
		), .Z(n_58424));
	notech_ao4 i_87750655(.A(n_59445), .B(n_26827), .C(n_56471), .D(n_26828)
		, .Z(n_287027252));
	notech_or4 i_118650710(.A(n_101413114), .B(n_58100), .C(instrc[121]), .D
		(n_58495), .Z(n_57863));
	notech_nand2 i_118850708(.A(n_56994), .B(n_26826), .Z(n_57861));
	notech_or4 i_104147716(.A(n_245362720), .B(n_58496), .C(n_57088), .D(n_57055
		), .Z(n_58008));
	notech_or4 i_104247717(.A(n_245362720), .B(n_57088), .C(n_29652), .D(n_58504
		), .Z(n_58007));
	notech_nao3 i_5747642(.A(n_319191632), .B(n_313391690), .C(n_246891941),
		 .Z(n_305624320));
	notech_nao3 i_59447778(.A(n_32380), .B(n_32298), .C(n_56837), .Z(n_58423
		));
	notech_nao3 i_118447768(.A(n_32338), .B(n_26731), .C(n_58496), .Z(n_57865
		));
	notech_nand2 i_118247770(.A(n_58632), .B(n_26641), .Z(n_57867));
	notech_and3 i_18056(.A(n_26964), .B(n_60241), .C(n_26985), .Z(n_330363520
		));
	notech_or4 i_4435066(.A(n_2839), .B(n_25617), .C(n_2864), .D(n_27123), .Z
		(n_305047803));
	notech_or4 i_24453985(.A(n_27917), .B(n_62848), .C(n_60949), .D(n_60246)
		, .Z(n_58773));
	notech_or4 i_107855517(.A(n_57088), .B(n_29652), .C(n_54916), .D(n_187662156
		), .Z(n_151931934));
	notech_ao4 i_51155533(.A(n_56859), .B(n_26962), .C(n_32352), .D(n_32291)
		, .Z(n_58506));
	notech_ao4 i_51555536(.A(n_56859), .B(n_26962), .C(n_32352), .D(n_32301)
		, .Z(n_58502));
	notech_or4 i_30771(.A(n_61175), .B(n_61165), .C(n_61154), .D(n_32257), .Z
		(n_154331958));
	notech_nand2 i_33068(.A(n_57988), .B(n_32291), .Z(n_154831963));
	notech_or4 i_176955537(.A(instrc[122]), .B(n_32339), .C(n_58099), .D(n_29179
		), .Z(n_57322));
	notech_or4 i_206755557(.A(n_32342), .B(n_32339), .C(n_58099), .D(n_58478
		), .Z(n_57025));
	notech_ao4 i_95055566(.A(n_60894), .B(n_26791), .C(n_62822), .D(n_60909)
		, .Z(n_58099));
	notech_or2 i_129155534(.A(n_58184), .B(n_56367), .Z(n_57758));
	notech_ao4 i_83355577(.A(n_60893), .B(n_26809), .C(n_62822), .D(n_60909)
		, .Z(n_58184));
	notech_or2 i_118155584(.A(n_26895), .B(n_58498), .Z(n_57868));
	notech_nao3 i_117455585(.A(n_32344), .B(n_26916), .C(n_58184), .Z(n_57875
		));
	notech_or2 i_181455515(.A(n_58099), .B(n_32331), .Z(n_151731932));
	notech_ao4 i_112355588(.A(n_58099), .B(n_32331), .C(n_59419), .D(n_26791
		), .Z(n_57926));
	notech_or4 i_96555592(.A(n_57088), .B(n_29652), .C(n_54916), .D(n_58498)
		, .Z(n_58084));
	notech_nao3 i_176255568(.A(n_32344), .B(n_26662), .C(n_58184), .Z(n_57329
		));
	notech_and2 i_87055595(.A(n_57329), .B(n_58194), .Z(n_58147));
	notech_ao4 i_86955596(.A(n_59445), .B(n_26811), .C(n_58173), .D(n_26662)
		, .Z(n_58148));
	notech_nao3 i_82355601(.A(n_58173), .B(n_32344), .C(n_58184), .Z(n_58194
		));
	notech_nand2 i_147955579(.A(n_59434), .B(n_58419), .Z(n_57602));
	notech_nand3 i_84455598(.A(n_56848), .B(n_188562161), .C(n_26812), .Z(n_58173
		));
	notech_ao4 i_59855615(.A(n_58184), .B(n_32344), .C(n_59418), .D(n_26809)
		, .Z(n_58419));
	notech_or4 i_58855616(.A(n_246891941), .B(n_2479), .C(n_56837), .D(n_56935
		), .Z(n_58429));
	notech_ao4 i_53955623(.A(n_56859), .B(n_32382), .C(n_32348), .D(n_32301)
		, .Z(n_58478));
	notech_ao4 i_53555624(.A(n_56859), .B(n_32382), .C(n_32348), .D(n_32291)
		, .Z(n_58482));
	notech_or2 i_53255626(.A(n_189362166), .B(n_305291771), .Z(n_58485));
	notech_ao4 i_53155627(.A(n_56859), .B(n_26610), .C(n_32356), .D(n_32301)
		, .Z(n_58486));
	notech_or2 i_52755628(.A(n_189662168), .B(n_305291771), .Z(n_58490));
	notech_ao4 i_51955631(.A(n_56859), .B(n_56935), .C(n_56684), .D(n_32291)
		, .Z(n_58498));
	notech_nao3 i_19155641(.A(n_57026), .B(n_29653), .C(n_30854), .Z(n_58802
		));
	notech_or4 i_14155643(.A(n_57026), .B(n_29653), .C(n_29658), .D(n_29652)
		, .Z(n_58805));
	notech_nand2 i_4158450(.A(n_60246), .B(read_data[4]), .Z(n_276134717));
	notech_and4 i_142341327(.A(n_298663253), .B(n_298563252), .C(n_298163248
		), .D(n_298463251), .Z(n_59993));
	notech_and4 i_117014(.A(n_186462146), .B(n_186362145), .C(n_186162144), 
		.D(n_186762149), .Z(n_17075));
	notech_and4 i_1121024(.A(n_184462127), .B(n_184662129), .C(n_185162134),
		 .D(n_179162074), .Z(n_14034));
	notech_nand2 i_1221025(.A(n_184362126), .B(n_183962122), .Z(n_14040));
	notech_and4 i_1321026(.A(n_182762110), .B(n_182962112), .C(n_183462117),
		 .D(n_181062093), .Z(n_14046));
	notech_nand2 i_24300(.A(n_56809), .B(opd[0]), .Z(n_35658));
	notech_ao4 i_52355630(.A(n_56859), .B(n_56935), .C(n_56684), .D(n_32301)
		, .Z(n_58494));
	notech_or2 i_118558528(.A(n_57322), .B(n_58494), .Z(n_57864));
	notech_and2 i_32858556(.A(n_182262105), .B(n_176362046), .Z(n_58689));
	notech_nand2 i_84544587(.A(n_58505), .B(n_58489), .Z(n_58172));
	notech_and4 i_143241320(.A(n_301763284), .B(n_301663283), .C(n_301263279
		), .D(n_301563282), .Z(n_59968));
	notech_nand2 i_192161727(.A(n_152961812), .B(n_26945), .Z(n_316537960)
		);
	notech_or2 i_108161760(.A(n_58810), .B(n_152861811), .Z(n_319937994));
	notech_or4 i_58961775(.A(n_59387), .B(n_56684), .C(n_29178), .D(n_27198)
		, .Z(n_321438009));
	notech_nand3 i_55661776(.A(n_318891635), .B(n_57988), .C(n_318791636), .Z
		(n_321538010));
	notech_nand2 i_517018(.A(n_174862031), .B(n_174262025), .Z(n_17099));
	notech_nand2 i_817021(.A(n_173562018), .B(n_172962012), .Z(n_17117));
	notech_nand2 i_1017023(.A(n_172362006), .B(n_171862001), .Z(n_17129));
	notech_nand2 i_1217025(.A(n_171261995), .B(n_170661989), .Z(n_17141));
	notech_or4 i_1617029(.A(n_159861881), .B(n_168761970), .C(n_26952), .D(n_26951
		), .Z(n_17165));
	notech_nand2 i_1421027(.A(n_168261965), .B(n_167861961), .Z(n_14052));
	notech_nand2 i_1521028(.A(n_167361956), .B(n_166961952), .Z(n_14058));
	notech_and4 i_1621029(.A(n_165761940), .B(n_165961942), .C(n_166461947),
		 .D(n_163461917), .Z(n_14064));
	notech_nand3 i_3121044(.A(n_165561938), .B(n_165461937), .C(n_165361936)
		, .Z(n_14154));
	notech_nand3 i_30428(.A(n_318891635), .B(n_57988), .C(n_319091633), .Z(n_322438019
		));
	notech_and2 i_146661796(.A(n_188857101), .B(n_274663013), .Z(n_57615));
	notech_ao4 i_146561797(.A(n_59445), .B(n_27079), .C(n_175762040), .D(n_26775
		), .Z(n_57616));
	notech_ao4 i_111361806(.A(n_61117), .B(n_30594), .C(n_305891765), .D(n_24589
		), .Z(n_57936));
	notech_and2 i_111261807(.A(n_102135817), .B(n_188857101), .Z(n_57937));
	notech_and3 i_106661808(.A(n_299591828), .B(n_274663013), .C(n_153561818
		), .Z(n_57983));
	notech_ao4 i_106561809(.A(n_61117), .B(n_27305), .C(n_307391750), .D(n_152761810
		), .Z(n_57984));
	notech_nand3 i_106161810(.A(n_32352), .B(n_32356), .C(n_56813), .Z(n_57988
		));
	notech_ao4 i_104661819(.A(n_61117), .B(n_30825), .C(n_24583), .D(n_305891765
		), .Z(n_58003));
	notech_and2 i_104561820(.A(n_2991), .B(n_153561818), .Z(n_58004));
	notech_or2 i_84861827(.A(n_175762040), .B(n_26775), .Z(n_58169));
	notech_and3 i_63661831(.A(n_308591738), .B(n_308491739), .C(n_306091763)
		, .Z(n_58381));
	notech_and3 i_60861832(.A(n_308591738), .B(n_308491739), .C(n_305791766)
		, .Z(n_58409));
	notech_or4 i_37141378(.A(n_60964), .B(n_60953), .C(n_62850), .D(\nbus_11307[0] 
		), .Z(n_58646));
	notech_or4 i_13355644(.A(n_57026), .B(n_57088), .C(n_29652), .D(n_29653)
		, .Z(n_58806));
	notech_and4 i_92038291(.A(n_314163408), .B(n_314063407), .C(n_313663403)
		, .D(n_313963406), .Z(n_60016));
	notech_ao4 i_127655543(.A(n_59993), .B(n_32356), .C(n_56837), .D(n_35658
		), .Z(n_57773));
	notech_and4 i_91138301(.A(n_311363380), .B(n_311263379), .C(n_310863375)
		, .D(n_311163378), .Z(n_60025));
	notech_or4 i_40741377(.A(n_60964), .B(n_60953), .C(n_62848), .D(n_29742)
		, .Z(n_58610));
	notech_ao4 i_7464379(.A(n_27907), .B(n_125461537), .C(n_61117), .D(n_127961562
		), .Z(n_248240500));
	notech_ao4 i_88555542(.A(n_60893), .B(n_26784), .C(n_62822), .D(n_60909)
		, .Z(n_58132));
	notech_ao4 i_4164412(.A(n_26975), .B(n_143561718), .C(n_27377), .D(n_26983
		), .Z(n_251540533));
	notech_nao3 i_11550723(.A(n_29658), .B(n_29652), .C(n_245362720), .Z(n_58817
		));
	notech_and4 i_11747718(.A(n_57026), .B(n_29658), .C(instrc[116]), .D(instrc
		[119]), .Z(n_58815));
	notech_or4 i_2864425(.A(n_60868), .B(n_27907), .C(n_61145), .D(n_60246),
		 .Z(n_252840546));
	notech_ao4 i_1964434(.A(n_32356), .B(n_5723), .C(n_26810), .D(n_27986), 
		.Z(n_253740555));
	notech_and4 i_121014(.A(n_186962151), .B(n_151361796), .C(n_151261795), 
		.D(n_130861591), .Z(n_13974));
	notech_nand2 i_221015(.A(n_150461787), .B(n_150061783), .Z(n_13980));
	notech_nand2 i_521018(.A(n_149561778), .B(n_149161774), .Z(n_13998));
	notech_or4 i_821021(.A(n_121375157), .B(n_133961622), .C(n_148461767), .D
		(n_26966), .Z(n_14016));
	notech_and4 i_1021023(.A(n_147061753), .B(n_147261755), .C(n_135861641),
		 .D(n_147661759), .Z(n_14028));
	notech_nand2 i_3564418(.A(pipe_mul[1]), .B(n_27376), .Z(n_252140539));
	notech_or4 i_13307(.A(n_32259), .B(n_32643), .C(n_61117), .D(n_59434), .Z
		(n_46630));
	notech_or4 i_2596(.A(n_319063457), .B(n_319263459), .C(n_319163458), .D(n_319363460
		), .Z(n_60094));
	notech_and4 i_121064489(.A(n_60094), .B(n_32605), .C(n_3792), .D(n_32562
		), .Z(n_57839));
	notech_or4 i_117264490(.A(n_32326), .B(n_32339), .C(n_58132), .D(n_58493
		), .Z(n_57877));
	notech_ao4 i_59564502(.A(n_32325), .B(n_58132), .C(n_59418), .D(n_26784)
		, .Z(n_58422));
	notech_nao3 i_59164503(.A(n_32380), .B(n_32287), .C(n_56837), .Z(n_58426
		));
	notech_ao4 i_54064505(.A(n_56859), .B(n_32382), .C(n_56813), .D(n_32299)
		, .Z(n_58477));
	notech_ao4 i_52464508(.A(n_56859), .B(n_56935), .C(n_56684), .D(n_32299)
		, .Z(n_58493));
	notech_and4 i_54157(.A(n_146361746), .B(n_144961732), .C(n_136961652), .D
		(n_144161724), .Z(\nbus_11356[16] ));
	notech_ao4 i_56145(.A(n_3598), .B(n_61145), .C(n_251540533), .D(n_32476)
		, .Z(\nbus_11376[10] ));
	notech_nand2 i_56146(.A(n_27570), .B(n_129161574), .Z(\nbus_11376[12] )
		);
	notech_or4 i_48701(.A(n_141261695), .B(n_138061663), .C(n_26994), .D(n_26976
		), .Z(\nbus_11302[0] ));
	notech_ao4 i_146853910(.A(n_28533), .B(n_330763524), .C(n_32656), .D(n_60241
		), .Z(n_330263519));
	notech_or4 i_37773(.A(n_59418), .B(n_27917), .C(n_60246), .D(n_26782), .Z
		(n_39041005));
	notech_or4 i_37778(.A(n_59418), .B(n_27917), .C(n_60229), .D(n_27896), .Z
		(n_40241017));
	notech_or4 i_25353984(.A(n_2875), .B(n_28081), .C(n_32443), .D(n_303747815
		), .Z(n_53341148));
	notech_or4 i_25453983(.A(n_305047803), .B(n_62834), .C(n_62822), .D(n_60229
		), .Z(n_53641151));
	notech_or4 i_25553982(.A(n_2875), .B(n_25617), .C(n_2877), .D(n_27105), 
		.Z(n_53841153));
	notech_or4 i_26453924(.A(n_27907), .B(n_62848), .C(n_60949), .D(n_60229)
		, .Z(n_54141156));
	notech_nand2 i_256938310(.A(n_50662), .B(n_305263319), .Z(n_60095));
	notech_or4 i_24935152(.A(n_61175), .B(n_61165), .C(n_61154), .D(n_60051)
		, .Z(n_58768));
	notech_or4 i_5067351(.A(n_55524), .B(n_330963526), .C(n_60373), .D(opd[0
		]), .Z(n_330063517));
	notech_nand2 i_4767354(.A(n_329663513), .B(n_123561518), .Z(n_329963516)
		);
	notech_nand2 i_4167360(.A(n_56542), .B(n_56632), .Z(n_329863515));
	notech_nor2 i_5885(.A(n_58813), .B(n_26721), .Z(n_329763514));
	notech_or2 i_35653(.A(n_19109), .B(n_60358), .Z(n_188810100));
	notech_nao3 i_1867382(.A(n_19101), .B(n_27981), .C(n_55524), .Z(n_25540870
		));
	notech_mux2 i_1367387(.S(opd[1]), .A(n_55508), .B(n_27040885), .Z(n_329663513
		));
	notech_nand3 i_134267397(.A(n_329663513), .B(n_123561518), .C(n_123661519
		), .Z(n_329563512));
	notech_ao4 i_98367398(.A(n_55524), .B(n_124061523), .C(n_329363510), .D(n_56566
		), .Z(n_329463511));
	notech_nor2 i_25967404(.A(n_121261495), .B(n_26781), .Z(n_329363510));
	notech_nand2 i_10267406(.A(n_19109), .B(n_60229), .Z(n_67341288));
	notech_nand3 i_3267407(.A(n_56542), .B(n_56632), .C(n_26920), .Z(n_329263509
		));
	notech_ao4 i_37759(.A(n_27907), .B(n_59418), .C(n_60893), .D(n_28533), .Z
		(n_329163508));
	notech_nao3 i_172367435(.A(n_121161494), .B(n_121061493), .C(n_83341448)
		, .Z(n_328963506));
	notech_nand2 i_318136(.A(n_120861491), .B(n_120761490), .Z(write_data_27
		[2]));
	notech_mux2 i_3212309(.S(n_60548), .A(n_6084), .B(regs_14[31]), .Z(pc_out
		[31]));
	notech_mux2 i_2612303(.S(n_60548), .A(n_6078), .B(regs_14[25]), .Z(pc_out
		[25]));
	notech_mux2 i_2512302(.S(n_60550), .A(n_6077), .B(regs_14[24]), .Z(pc_out
		[24]));
	notech_mux2 i_2412301(.S(n_60550), .A(n_6076), .B(regs_14[23]), .Z(pc_out
		[23]));
	notech_mux2 i_2312300(.S(n_60550), .A(n_6075), .B(regs_14[22]), .Z(pc_out
		[22]));
	notech_mux2 i_2112298(.S(n_60550), .A(n_6073), .B(regs_14[20]), .Z(pc_out
		[20]));
	notech_ao4 i_113383448(.A(n_32579), .B(n_327363490), .C(n_1878), .D(n_27069
		), .Z(n_328763504));
	notech_and2 i_37495(.A(n_22024), .B(n_330463521), .Z(n_328463501));
	notech_and3 i_33183443(.A(n_326963486), .B(n_326891248), .C(n_326791249)
		, .Z(n_328163498));
	notech_nand3 i_426953(.A(n_328763504), .B(n_327863495), .C(n_327563492),
		 .Z(n_19665));
	notech_nao3 i_113183440(.A(n_60162), .B(n_60358), .C(n_327463491), .Z(n_327863495
		));
	notech_nand3 i_112983438(.A(n_327263489), .B(n_330563522), .C(n_22015), 
		.Z(n_327663493));
	notech_nand2 i_113283437(.A(n_60158), .B(n_327663493), .Z(n_327563492)
		);
	notech_and2 i_112883436(.A(n_331163528), .B(n_328463501), .Z(n_327463491
		));
	notech_ao4 i_112383435(.A(n_29655), .B(n_26755), .C(n_3790), .D(n_26758)
		, .Z(n_327363490));
	notech_or4 i_112683434(.A(n_5221), .B(n_330963526), .C(n_2946), .D(n_60373
		), .Z(n_327263489));
	notech_or4 i_57883432(.A(n_2839), .B(n_2888), .C(n_60949), .D(n_60909), 
		.Z(n_327063487));
	notech_or4 i_57583431(.A(n_59418), .B(n_27501), .C(n_32747), .D(n_62892)
		, .Z(n_326963486));
	notech_or4 i_57383430(.A(n_27501), .B(n_1868), .C(n_60949), .D(n_60909),
		 .Z(n_326891248));
	notech_or4 i_57483429(.A(n_27501), .B(\opcode[0] ), .C(n_32730), .D(n_59435
		), .Z(n_326791249));
	notech_ao4 i_45383427(.A(n_27907), .B(n_330763524), .C(n_60229), .D(n_326491252
		), .Z(n_326591251));
	notech_and3 i_45283426(.A(n_1897), .B(n_1898), .C(n_1881), .Z(n_326491252
		));
	notech_nand3 i_76232085(.A(n_19137), .B(n_26964), .C(n_60229), .Z(n_325891258
		));
	notech_and4 i_78532062(.A(n_58662), .B(n_53731), .C(n_325491262), .D(n_60136
		), .Z(n_325791259));
	notech_and4 i_78432063(.A(n_320163468), .B(n_17779989), .C(n_53739), .D(n_317163438
		), .Z(n_325491262));
	notech_and3 i_78732060(.A(n_324463483), .B(n_17539965), .C(n_5968810), .Z
		(n_325191265));
	notech_ao4 i_78832059(.A(n_18998), .B(n_27069), .C(write_ack), .D(n_57285
		), .Z(n_324891268));
	notech_ao4 i_78932058(.A(n_319391630), .B(n_58664), .C(n_61117), .D(n_315663423
		), .Z(n_324791269));
	notech_ao4 i_21832552(.A(n_17669978), .B(n_29656), .C(n_32579), .D(n_324363482
		), .Z(n_324463483));
	notech_nand2 i_80032047(.A(n_19022), .B(n_29655), .Z(n_324363482));
	notech_ao4 i_99631871(.A(n_60868), .B(n_27904), .C(n_27063), .D(n_1881),
		 .Z(n_324263481));
	notech_ao4 i_107731792(.A(n_61117), .B(n_316963436), .C(n_317063437), .D
		(n_61145), .Z(n_324091270));
	notech_and3 i_108131788(.A(n_53341148), .B(n_53641151), .C(n_53841153), 
		.Z(n_323791273));
	notech_or4 i_24332531(.A(n_32565), .B(n_3812), .C(n_314463411), .D(n_19043
		), .Z(n_323563479));
	notech_or4 i_111931754(.A(opc[30]), .B(opc[31]), .C(opc[27]), .D(n_322991279
		), .Z(n_323291277));
	notech_nao3 i_111831755(.A(nbus_11295[29]), .B(nbus_11295[26]), .C(opc[
		28]), .Z(n_322991279));
	notech_or4 i_112431749(.A(opc[23]), .B(opc[24]), .C(opc[25]), .D(n_322491283
		), .Z(n_322791280));
	notech_nand3 i_112331750(.A(nbus_11295[20]), .B(nbus_11295[21]), .C(nbus_11295
		[22]), .Z(n_322491283));
	notech_or4 i_113131743(.A(opc[17]), .B(opc[18]), .C(opc[19]), .D(n_321891287
		), .Z(n_322163476));
	notech_nand3 i_112931744(.A(nbus_11295[14]), .B(nbus_11295[15]), .C(nbus_11295
		[16]), .Z(n_321891287));
	notech_or4 i_113931738(.A(opc[11]), .B(opc[12]), .C(opc[13]), .D(n_321391291
		), .Z(n_321663474));
	notech_nand3 i_113831739(.A(nbus_11295[8]), .B(nbus_11295[9]), .C(nbus_11295
		[10]), .Z(n_321391291));
	notech_xor2 i_114231735(.A(opc[3]), .B(n_60095), .Z(n_320991294));
	notech_and2 i_141332701(.A(n_320163468), .B(n_317163438), .Z(n_320263469
		));
	notech_or2 i_30032483(.A(n_5018715), .B(n_320063467), .Z(n_320163468));
	notech_nand3 i_16132581(.A(n_19137), .B(n_60158), .C(n_60229), .Z(n_320063467
		));
	notech_or4 i_35946(.A(n_61175), .B(n_61165), .C(n_27037), .D(n_19101), .Z
		(n_319963466));
	notech_nor2 i_65432181(.A(n_50662), .B(opc[4]), .Z(n_319763464));
	notech_and2 i_65532180(.A(opc[4]), .B(n_50662), .Z(n_319463461));
	notech_and2 i_64832187(.A(n_317463441), .B(n_17409952), .Z(n_319363460)
		);
	notech_ao4 i_64732188(.A(n_291118110), .B(opc[4]), .C(n_27054), .D(n_317763444
		), .Z(n_319263459));
	notech_and2 i_65032185(.A(n_317663443), .B(n_26759), .Z(n_319163458));
	notech_and3 i_64932186(.A(\nbus_11307[0] ), .B(n_27050), .C(n_317563442)
		, .Z(n_319063457));
	notech_and3 i_37523(.A(n_32434), .B(n_2419), .C(n_58786), .Z(n_318563452
		));
	notech_ao4 i_22532545(.A(n_319391630), .B(n_19029), .C(n_29282), .D(n_315463421
		), .Z(n_318063447));
	notech_or2 i_38332417(.A(n_320063467), .B(n_26964), .Z(n_317963446));
	notech_or4 i_38232418(.A(n_318063447), .B(n_61145), .C(n_19050), .D(n_325891258
		), .Z(n_317863445));
	notech_ao3 i_65132184(.A(rep_en5), .B(\nbus_11365[31] ), .C(n_58675), .Z
		(n_317763444));
	notech_or4 i_34732447(.A(n_323291277), .B(n_322791280), .C(n_322163476),
		 .D(n_321663474), .Z(n_317663443));
	notech_or4 i_34632448(.A(n_290618105), .B(n_319463461), .C(n_319763464),
		 .D(n_320991294), .Z(n_317563442));
	notech_or4 i_34532449(.A(opc[6]), .B(opc[7]), .C(n_57896), .D(opc[5]), .Z
		(n_317463441));
	notech_nand2 i_36932431(.A(n_1880), .B(n_60074), .Z(n_317263439));
	notech_nand3 i_64132194(.A(n_60158), .B(n_60356), .C(n_317263439), .Z(n_317163438
		));
	notech_and4 i_62432210(.A(n_58773), .B(n_1887), .C(n_58768), .D(n_323791273
		), .Z(n_317063437));
	notech_and4 i_62332211(.A(n_313784128), .B(n_32656), .C(n_329163508), .D
		(n_60074), .Z(n_316963436));
	notech_ao4 i_62232212(.A(n_319791626), .B(n_26964), .C(n_25397), .D(n_56566
		), .Z(n_316763434));
	notech_ao4 i_62132213(.A(n_323563479), .B(n_325684247), .C(n_316763434),
		 .D(n_32581), .Z(n_316463431));
	notech_or4 i_29932484(.A(n_316463431), .B(n_61145), .C(n_60358), .D(n_26900
		), .Z(n_316363430));
	notech_nand2 i_62032214(.A(n_324091270), .B(n_316363430), .Z(n_316263429
		));
	notech_ao4 i_61932215(.A(n_320163468), .B(n_29657), .C(n_5221), .D(n_17539965
		), .Z(n_315963426));
	notech_and4 i_36132438(.A(n_319591628), .B(n_318563452), .C(n_328463501)
		, .D(n_328163498), .Z(n_315663423));
	notech_ao3 i_20032570(.A(n_27065), .B(n_320291621), .C(n_18981), .Z(n_315463421
		));
	notech_mux2 i_27632503(.S(n_19043), .A(n_19036), .B(n_3848598), .Z(n_315063417
		));
	notech_or4 i_37932421(.A(n_19127), .B(n_315063417), .C(n_61143), .D(n_60358
		), .Z(n_314963416));
	notech_nao3 i_26841404(.A(rep_en3), .B(n_27378), .C(rep_en2), .Z(n_314863415
		));
	notech_nand3 i_26932715(.A(n_60158), .B(n_60229), .C(n_32586), .Z(n_314663413
		));
	notech_or4 i_35817(.A(n_2875), .B(n_28081), .C(n_2877), .D(n_1864), .Z(n_314563412
		));
	notech_nand3 i_28996(.A(n_19093), .B(n_60373), .C(n_26964), .Z(n_314463411
		));
	notech_ao4 i_196136347(.A(n_57985), .B(n_28298), .C(n_28492), .D(n_27104
		), .Z(n_314163408));
	notech_ao4 i_196236346(.A(n_27867), .B(n_58014), .C(n_56468), .D(n_29789
		), .Z(n_314063407));
	notech_and2 i_196636342(.A(n_313863405), .B(n_313763404), .Z(n_313963406
		));
	notech_ao4 i_196436344(.A(n_56396), .B(n_28167), .C(n_56391), .D(n_28396
		), .Z(n_313863405));
	notech_ao4 i_196536343(.A(n_28526), .B(n_59344), .C(n_56367), .D(n_28331
		), .Z(n_313763404));
	notech_and4 i_197436334(.A(n_313463401), .B(n_313363400), .C(n_313163398
		), .D(n_313063397), .Z(n_313663403));
	notech_ao4 i_196836340(.A(n_56452), .B(n_28266), .C(n_27089), .D(n_28460
		), .Z(n_313463401));
	notech_ao4 i_196936339(.A(n_56447), .B(n_28232), .C(n_56432), .D(n_28199
		), .Z(n_313363400));
	notech_ao4 i_197136337(.A(n_56909), .B(n_29788), .C(n_28364), .D(n_56427
		), .Z(n_313163398));
	notech_ao4 i_197236336(.A(n_27094), .B(n_28428), .C(n_26950), .D(n_28570
		), .Z(n_313063397));
	notech_ao4 i_203136277(.A(n_57976), .B(n_28293), .C(n_28487), .D(n_27104
		), .Z(n_312763394));
	notech_ao4 i_203236276(.A(n_27862), .B(n_58014), .C(n_56468), .D(n_29791
		), .Z(n_312663393));
	notech_and2 i_203636272(.A(n_312463391), .B(n_312363390), .Z(n_312563392
		));
	notech_ao4 i_203436274(.A(n_56396), .B(n_28162), .C(n_56391), .D(n_28391
		), .Z(n_312463391));
	notech_ao4 i_203536273(.A(n_28520), .B(n_59344), .C(n_56367), .D(n_28326
		), .Z(n_312363390));
	notech_and4 i_204436264(.A(n_312063387), .B(n_311963386), .C(n_311763384
		), .D(n_311663383), .Z(n_312263389));
	notech_ao4 i_203836270(.A(n_56452), .B(n_28261), .C(n_27089), .D(n_28455
		), .Z(n_312063387));
	notech_ao4 i_203936269(.A(n_56443), .B(n_28227), .C(n_56432), .D(n_28194
		), .Z(n_311963386));
	notech_ao4 i_204136267(.A(n_56909), .B(n_29790), .C(n_28359), .D(n_56423
		), .Z(n_311763384));
	notech_ao4 i_204236266(.A(n_56414), .B(n_28423), .C(n_56405), .D(n_28564
		), .Z(n_311663383));
	notech_ao4 i_207336235(.A(n_57976), .B(n_28289), .C(n_28483), .D(n_27104
		), .Z(n_311363380));
	notech_ao4 i_207436234(.A(n_27858), .B(n_58014), .C(n_56463), .D(n_29792
		), .Z(n_311263379));
	notech_and2 i_207836230(.A(n_311063377), .B(n_310963376), .Z(n_311163378
		));
	notech_ao4 i_207636232(.A(n_56396), .B(n_28158), .C(n_56391), .D(n_28387
		), .Z(n_311063377));
	notech_ao4 i_207736231(.A(n_59344), .B(n_28516), .C(n_28322), .D(n_56371
		), .Z(n_310963376));
	notech_and4 i_208636222(.A(n_310663373), .B(n_310563372), .C(n_310363370
		), .D(n_310263369), .Z(n_310863375));
	notech_ao4 i_208036228(.A(n_28257), .B(n_56452), .C(n_58020), .D(n_28451
		), .Z(n_310663373));
	notech_ao4 i_208136227(.A(n_56443), .B(n_28223), .C(n_56432), .D(n_28190
		), .Z(n_310563372));
	notech_ao4 i_208336225(.A(n_56909), .B(n_27849), .C(n_28355), .D(n_56423
		), .Z(n_310363370));
	notech_ao4 i_208436224(.A(n_56414), .B(n_28419), .C(n_56405), .D(n_28560
		), .Z(n_310263369));
	notech_nand3 i_116837134(.A(opz[1]), .B(n_28051), .C(n_28049), .Z(n_305263319
		));
	notech_and4 i_137139991(.A(n_304963316), .B(n_304763314), .C(n_287463141
		), .D(n_287763144), .Z(n_305163318));
	notech_ao4 i_136739995(.A(n_151761800), .B(n_29786), .C(n_5933), .D(n_57937
		), .Z(n_304963316));
	notech_ao4 i_136939993(.A(n_57983), .B(\nbus_11358[8] ), .C(n_58381), .D
		(n_27991), .Z(n_304763314));
	notech_and4 i_137739985(.A(n_304463311), .B(n_304263309), .C(n_304163308
		), .D(n_288063147), .Z(n_304663313));
	notech_ao4 i_137239990(.A(n_57984), .B(\nbus_11307[8] ), .C(n_60162), .D
		(n_27127), .Z(n_304463311));
	notech_ao4 i_137439988(.A(n_293018129), .B(n_305791766), .C(n_309666625)
		, .D(n_152061803), .Z(n_304263309));
	notech_ao4 i_137539987(.A(n_308066609), .B(n_57799), .C(n_308166610), .D
		(n_24589), .Z(n_304163308));
	notech_and4 i_163639748(.A(n_334480845), .B(n_303763304), .C(n_288563152
		), .D(n_288863155), .Z(n_304063307));
	notech_ao4 i_163439750(.A(n_5933), .B(n_285563122), .C(n_29787), .D(n_291063177
		), .Z(n_303763304));
	notech_ao4 i_163739747(.A(n_308066609), .B(n_290963176), .C(n_308166610)
		, .D(n_286463131), .Z(n_303563302));
	notech_ao4 i_163839746(.A(\nbus_11307[8] ), .B(n_285763124), .C(n_309666625
		), .D(n_286263129), .Z(n_303363300));
	notech_and4 i_170239685(.A(n_289663163), .B(n_303063297), .C(n_302863295
		), .D(n_302763294), .Z(n_303263299));
	notech_ao4 i_169739690(.A(n_28093), .B(n_309291731), .C(n_5743), .D(n_316991654
		), .Z(n_303063297));
	notech_ao4 i_169939688(.A(n_60162), .B(n_27249), .C(n_58081), .D(\nbus_11358[4] 
		), .Z(n_302863295));
	notech_ao4 i_170039687(.A(n_317991644), .B(n_5723), .C(n_58406), .D(n_27986
		), .Z(n_302763294));
	notech_and4 i_170939678(.A(n_302463291), .B(n_302363290), .C(n_302163288
		), .D(n_302063287), .Z(n_302663293));
	notech_ao4 i_170339684(.A(n_122628503), .B(n_29542), .C(n_291563182), .D
		(n_56533), .Z(n_302463291));
	notech_ao4 i_170439683(.A(n_317091653), .B(n_291463181), .C(n_285663123)
		, .D(\nbus_11307[4] ), .Z(n_302363290));
	notech_ao4 i_170639681(.A(n_291663183), .B(n_285963126), .C(n_291763184)
		, .D(n_286063127), .Z(n_302163288));
	notech_ao4 i_170739680(.A(n_291863185), .B(n_286163128), .C(n_286363130)
		, .D(n_29725), .Z(n_302063287));
	notech_ao4 i_194839451(.A(n_28232), .B(n_26924), .C(n_28199), .D(n_56649
		), .Z(n_301763284));
	notech_ao4 i_194939450(.A(n_56921), .B(n_29788), .C(n_28266), .D(n_56636
		), .Z(n_301663283));
	notech_and2 i_195339446(.A(n_301463281), .B(n_301363280), .Z(n_301563282
		));
	notech_ao4 i_195139448(.A(n_56527), .B(n_28298), .C(n_56513), .D(n_29789
		), .Z(n_301463281));
	notech_ao4 i_195239447(.A(n_26920), .B(n_28364), .C(n_56485), .D(n_28331
		), .Z(n_301363280));
	notech_and4 i_196139438(.A(n_301063277), .B(n_300963276), .C(n_300763274
		), .D(n_300663273), .Z(n_301263279));
	notech_ao4 i_195539444(.A(n_28428), .B(n_56632), .C(n_56614), .D(n_28396
		), .Z(n_301063277));
	notech_ao4 i_195639443(.A(n_26928), .B(n_28460), .C(n_56592), .D(n_28167
		), .Z(n_300963276));
	notech_ao4 i_195839441(.A(n_26925), .B(n_28492), .C(n_56566), .D(n_28526
		), .Z(n_300763274));
	notech_ao4 i_195939440(.A(n_26721), .B(n_27867), .C(n_56542), .D(n_28570
		), .Z(n_300663273));
	notech_ao4 i_196439436(.A(n_28227), .B(n_26924), .C(n_28194), .D(n_56649
		), .Z(n_300263269));
	notech_ao4 i_196539435(.A(n_56921), .B(n_29790), .C(n_28261), .D(n_56636
		), .Z(n_300163268));
	notech_and2 i_196939431(.A(n_299963266), .B(n_299863265), .Z(n_300063267
		));
	notech_ao4 i_196739433(.A(n_28293), .B(n_56527), .C(n_56513), .D(n_29791
		), .Z(n_299963266));
	notech_ao4 i_196839432(.A(n_56502), .B(n_28359), .C(n_56485), .D(n_28326
		), .Z(n_299863265));
	notech_and4 i_197739423(.A(n_299563262), .B(n_299463261), .C(n_299263259
		), .D(n_299163258), .Z(n_299763264));
	notech_ao4 i_197139429(.A(n_28423), .B(n_56632), .C(n_56614), .D(n_28391
		), .Z(n_299563262));
	notech_ao4 i_197239428(.A(n_26928), .B(n_28455), .C(n_56592), .D(n_28162
		), .Z(n_299463261));
	notech_ao4 i_197439426(.A(n_28487), .B(n_26925), .C(n_56566), .D(n_28520
		), .Z(n_299263259));
	notech_ao4 i_197539425(.A(n_26721), .B(n_27862), .C(n_56542), .D(n_28564
		), .Z(n_299163258));
	notech_ao4 i_199539406(.A(n_28223), .B(n_56662), .C(n_28190), .D(n_56649
		), .Z(n_298663253));
	notech_ao4 i_199639405(.A(n_56921), .B(n_27849), .C(n_56636), .D(n_28257
		), .Z(n_298563252));
	notech_and2 i_200039401(.A(n_298363250), .B(n_298263249), .Z(n_298463251
		));
	notech_ao4 i_199839403(.A(n_28289), .B(n_56527), .C(n_56513), .D(n_29792
		), .Z(n_298363250));
	notech_ao4 i_199939402(.A(n_56498), .B(n_28355), .C(n_56485), .D(n_28322
		), .Z(n_298263249));
	notech_and4 i_200839393(.A(n_297963246), .B(n_297863245), .C(n_297663243
		), .D(n_297563242), .Z(n_298163248));
	notech_ao4 i_200239399(.A(n_56632), .B(n_28419), .C(n_56614), .D(n_28387
		), .Z(n_297963246));
	notech_ao4 i_200339398(.A(n_26928), .B(n_28451), .C(n_56592), .D(n_28158
		), .Z(n_297863245));
	notech_ao4 i_200539396(.A(n_28483), .B(n_26925), .C(n_56566), .D(n_28516
		), .Z(n_297663243));
	notech_ao4 i_200639395(.A(n_27858), .B(n_56553), .C(n_28560), .D(n_56542
		), .Z(n_297563242));
	notech_ao4 i_105864494(.A(n_175162034), .B(n_32319), .C(n_59419), .D(n_26945
		), .Z(n_297363240));
	notech_or2 i_98840334(.A(n_125561538), .B(n_287163138), .Z(n_296963236)
		);
	notech_or4 i_160564479(.A(n_32342), .B(n_175162034), .C(n_285463121), .D
		(n_26735), .Z(n_296863235));
	notech_nand2 i_28583(.A(opc_10[9]), .B(n_62806), .Z(n_291963186));
	notech_nand2 i_28817(.A(opc_10[4]), .B(n_62806), .Z(n_291863185));
	notech_nand2 i_28818(.A(opc[4]), .B(n_62778), .Z(n_291763184));
	notech_nao3 i_28821(.A(n_62826), .B(opa[4]), .C(n_62860), .Z(n_291663183
		));
	notech_or4 i_28823(.A(n_60964), .B(n_60953), .C(n_62846), .D(\nbus_11307[4] 
		), .Z(n_291563182));
	notech_or4 i_28841(.A(n_60964), .B(n_60953), .C(n_62860), .D(n_29725), .Z
		(n_291463181));
	notech_nand3 i_29092(.A(n_60909), .B(n_62808), .C(\opa_12[0] ), .Z(n_291363180
		));
	notech_nand2 i_29096(.A(opc[0]), .B(n_62808), .Z(n_291263179));
	notech_nand2 i_29097(.A(opc_10[0]), .B(n_62816), .Z(n_291163178));
	notech_or2 i_30533(.A(n_286463131), .B(n_297363240), .Z(n_291063177));
	notech_or2 i_30539(.A(n_286463131), .B(n_174962032), .Z(n_290963176));
	notech_nao3 i_66440639(.A(n_11407), .B(n_32272), .C(n_2868), .Z(n_289663163
		));
	notech_nao3 i_55740728(.A(n_318891635), .B(n_319091633), .C(n_325270263)
		, .Z(n_289363160));
	notech_or2 i_56240723(.A(n_286563132), .B(n_27991), .Z(n_288863155));
	notech_nand2 i_56340722(.A(opb[8]), .B(n_286663133), .Z(n_288563152));
	notech_or4 i_41740857(.A(n_61143), .B(n_60358), .C(n_19086), .D(n_28097)
		, .Z(n_288063147));
	notech_or2 i_42040854(.A(n_57936), .B(n_29787), .Z(n_287763144));
	notech_nand3 i_42340851(.A(n_310991714), .B(\regs_1[8] ), .C(n_28680), .Z
		(n_287463141));
	notech_and3 i_90864498(.A(n_56848), .B(n_127161554), .C(n_281263079), .Z
		(n_287163138));
	notech_or4 i_98740335(.A(n_59387), .B(n_4011), .C(n_29178), .D(n_27192),
		 .Z(n_287063137));
	notech_nand2 i_79440510(.A(n_287163138), .B(n_285463121), .Z(n_286763134
		));
	notech_nand3 i_109841339(.A(n_296863235), .B(n_285363120), .C(n_296963236
		), .Z(n_286663133));
	notech_and2 i_64641338(.A(n_58426), .B(n_287063137), .Z(n_286563132));
	notech_ao4 i_54164504(.A(n_56858), .B(n_32382), .C(n_56813), .D(n_32287)
		, .Z(n_286463131));
	notech_or2 i_154641252(.A(n_317091653), .B(n_318991634), .Z(n_286363130)
		);
	notech_nand2 i_139641257(.A(n_286763134), .B(n_26945), .Z(n_286263129)
		);
	notech_nao3 i_139141258(.A(n_246591944), .B(n_29652), .C(n_317091653), .Z
		(n_286163128));
	notech_nao3 i_130641260(.A(n_29652), .B(n_246591944), .C(n_56533), .Z(n_286063127
		));
	notech_or2 i_128641262(.A(n_32393), .B(n_56533), .Z(n_285963126));
	notech_nand2 i_38441394(.A(n_59435), .B(n_297363240), .Z(n_285863125));
	notech_nand2 i_100641269(.A(n_286763134), .B(n_285863125), .Z(n_285763124
		));
	notech_nao3 i_96941272(.A(n_56396), .B(n_27194), .C(n_56533), .Z(n_285663123
		));
	notech_or4 i_176841305(.A(n_32342), .B(n_175162034), .C(n_286463131), .D
		(n_26735), .Z(n_285563122));
	notech_ao4 i_53364506(.A(n_56854), .B(n_26610), .C(n_32356), .D(n_32287)
		, .Z(n_285463121));
	notech_or4 i_68864501(.A(n_32643), .B(n_32259), .C(n_60229), .D(n_59435)
		, .Z(n_285363120));
	notech_and4 i_184342746(.A(n_216676105), .B(n_285063117), .C(n_284863115
		), .D(n_277463041), .Z(n_285263119));
	notech_ao4 i_183942750(.A(n_60022), .B(n_296863235), .C(n_29728), .D(n_136461647
		), .Z(n_285063117));
	notech_ao4 i_184142748(.A(n_275463021), .B(\nbus_11358[3] ), .C(n_135961642
		), .D(n_27985), .Z(n_284863115));
	notech_and4 i_184842741(.A(n_277763044), .B(n_284563112), .C(n_284363110
		), .D(n_278063047), .Z(n_284763114));
	notech_ao4 i_184442745(.A(n_306970080), .B(n_285463121), .C(n_306870079)
		, .D(n_274763014), .Z(n_284563112));
	notech_ao4 i_184642743(.A(n_306670077), .B(n_136361646), .C(n_306570076)
		, .D(n_275363020), .Z(n_284363110));
	notech_and4 i_185342736(.A(n_216276101), .B(n_284063107), .C(n_283863105
		), .D(n_278563052), .Z(n_284263109));
	notech_ao4 i_184942740(.A(n_60020), .B(n_296863235), .C(n_136461647), .D
		(n_29651), .Z(n_284063107));
	notech_ao4 i_185142738(.A(n_275463021), .B(\nbus_11358[5] ), .C(n_135961642
		), .D(n_27987), .Z(n_283863105));
	notech_and4 i_185842731(.A(n_278863055), .B(n_283563102), .C(n_283363100
		), .D(n_279163058), .Z(n_283763104));
	notech_ao4 i_185442735(.A(n_282266351), .B(n_285463121), .C(n_282166350)
		, .D(n_274763014), .Z(n_283563102));
	notech_ao4 i_185642733(.A(n_281966348), .B(n_275363020), .C(n_281866347)
		, .D(n_136361646), .Z(n_283363100));
	notech_and4 i_186242727(.A(n_311173591), .B(n_282963096), .C(n_279263059
		), .D(n_279563062), .Z(n_283263099));
	notech_ao4 i_186042729(.A(n_135961642), .B(n_27989), .C(n_3868), .D(n_136561648
		), .Z(n_282963096));
	notech_and4 i_186742722(.A(n_282663093), .B(n_280163068), .C(n_282463091
		), .D(n_279863065), .Z(n_282863095));
	notech_ao4 i_186342726(.A(n_92019102), .B(n_274763014), .C(n_275363020),
		 .D(n_306273542), .Z(n_282663093));
	notech_ao4 i_186542724(.A(n_136161644), .B(n_275263019), .C(n_285463121)
		, .D(n_275163018), .Z(n_282463091));
	notech_mux2 i_186842721(.S(n_32319), .A(n_309973579), .B(n_310073580), .Z
		(n_282363090));
	notech_ao4 i_187042719(.A(n_314791676), .B(n_164761930), .C(n_29619), .D
		(n_275863025), .Z(n_282063087));
	notech_nand3 i_187542714(.A(n_281663083), .B(n_281863085), .C(n_281163078
		), .Z(n_281963086));
	notech_ao4 i_187242717(.A(n_314391680), .B(n_136561648), .C(n_83019012),
		 .D(n_275763024), .Z(n_281863085));
	notech_ao4 i_187342716(.A(n_306221226), .B(n_56632), .C(\nbus_11365[31] 
		), .D(n_151661799), .Z(n_281663083));
	notech_nand2 i_35552(.A(n_26718), .B(n_26960), .Z(n_281463081));
	notech_nand2 i_9644398(.A(n_26718), .B(n_58169), .Z(n_281363080));
	notech_ao4 i_52564507(.A(n_56854), .B(n_56946), .C(n_56684), .D(n_32287)
		, .Z(n_281263079));
	notech_or4 i_86543669(.A(n_281263079), .B(n_174962032), .C(n_60949), .D(nbus_11295
		[31]), .Z(n_281163078));
	notech_nor2 i_87443664(.A(n_275963026), .B(\nbus_11358[31] ), .Z(n_280463071
		));
	notech_or4 i_85043683(.A(n_62856), .B(n_136361646), .C(n_60949), .D(\nbus_11307[6] 
		), .Z(n_280163068));
	notech_or4 i_85443680(.A(n_275363020), .B(n_60947), .C(nbus_11295[6]), .D
		(n_174962032), .Z(n_279863065));
	notech_or2 i_85743677(.A(n_275463021), .B(\nbus_11358[6] ), .Z(n_279563062
		));
	notech_nao3 i_85843676(.A(n_126061543), .B(opa[6]), .C(n_140661689), .Z(n_279263059
		));
	notech_nao3 i_83843694(.A(opc[5]), .B(n_62808), .C(n_136261645), .Z(n_279163058
		));
	notech_or4 i_84143691(.A(n_56837), .B(n_26610), .C(n_56632), .D(n_308621250
		), .Z(n_278863055));
	notech_nao3 i_84443688(.A(n_126061543), .B(opa[5]), .C(n_140661689), .Z(n_278563052
		));
	notech_or4 i_82743705(.A(n_275363020), .B(nbus_11295[3]), .C(n_60945), .D
		(n_174962032), .Z(n_278063047));
	notech_or4 i_83043702(.A(n_56839), .B(n_26610), .C(n_56632), .D(n_308721251
		), .Z(n_277763044));
	notech_nao3 i_83343699(.A(n_126061543), .B(opa[3]), .C(n_140661689), .Z(n_277463041
		));
	notech_or2 i_126043302(.A(n_305991764), .B(n_26774), .Z(n_276363030));
	notech_nand3 i_131764485(.A(n_56848), .B(n_127161554), .C(n_286463131), 
		.Z(n_276163028));
	notech_nand2 i_124543317(.A(n_276163028), .B(n_26945), .Z(n_276063027)
		);
	notech_and2 i_98764497(.A(n_285363120), .B(n_164361926), .Z(n_275963026)
		);
	notech_and2 i_147344530(.A(n_274963016), .B(n_275063017), .Z(n_275863025
		));
	notech_and2 i_150544532(.A(n_274763014), .B(n_276063027), .Z(n_275763024
		));
	notech_and2 i_109764493(.A(n_275963026), .B(n_127061553), .Z(n_275463021
		));
	notech_and2 i_123364487(.A(n_287163138), .B(n_286463131), .Z(n_275363020
		));
	notech_and2 i_12444372(.A(n_92519107), .B(n_282363090), .Z(n_275263019)
		);
	notech_mux2 i_12344373(.S(n_32319), .A(n_305721221), .B(n_305621220), .Z
		(n_275163018));
	notech_nand2 i_13623(.A(n_285863125), .B(n_26834), .Z(n_275063017));
	notech_nand2 i_186864476(.A(n_285863125), .B(n_164961932), .Z(n_274963016
		));
	notech_nao3 i_186964475(.A(n_164961932), .B(n_32319), .C(n_175162034), .Z
		(n_274863015));
	notech_or2 i_116864491(.A(n_285463121), .B(n_174962032), .Z(n_274763014)
		);
	notech_nao3 i_88761826(.A(n_175762040), .B(n_32316), .C(n_307691747), .Z
		(n_274663013));
	notech_and3 i_173546025(.A(n_194675885), .B(n_274363010), .C(n_253662803
		), .Z(n_274563012));
	notech_ao4 i_173446026(.A(n_60009), .B(n_164761930), .C(n_29710), .D(n_275863025
		), .Z(n_274363010));
	notech_ao4 i_173646024(.A(n_313747721), .B(n_136561648), .C(n_254466073)
		, .D(n_275763024), .Z(n_274163008));
	notech_ao4 i_173746023(.A(n_311224366), .B(n_56632), .C(n_281263079), .D
		(n_250762774), .Z(n_273963006));
	notech_ao4 i_174046020(.A(n_28106), .B(n_60358), .C(n_251362780), .D(n_56293
		), .Z(n_273763004));
	notech_ao4 i_174146019(.A(n_251162778), .B(n_29772), .C(n_58426), .D(n_28002
		), .Z(n_273563002));
	notech_and3 i_174746013(.A(n_273162998), .B(n_273363000), .C(n_255262819
		), .Z(n_273463001));
	notech_ao4 i_174446016(.A(n_313647722), .B(n_322438019), .C(n_249672976)
		, .D(n_316537960), .Z(n_273363000));
	notech_ao4 i_174546015(.A(n_254673026), .B(n_281263079), .C(n_251062777)
		, .D(n_57689), .Z(n_273162998));
	notech_ao4 i_174846012(.A(n_28107), .B(n_60358), .C(n_251362780), .D(\nbus_11358[18] 
		), .Z(n_272962996));
	notech_ao4 i_174946011(.A(n_251162778), .B(n_29711), .C(n_58426), .D(n_28003
		), .Z(n_272762994));
	notech_and3 i_175546005(.A(n_272362990), .B(n_272562992), .C(n_256162828
		), .Z(n_272662993));
	notech_ao4 i_175246008(.A(n_3861), .B(n_322438019), .C(n_77522039), .D(n_316537960
		), .Z(n_272562992));
	notech_ao4 i_175346007(.A(n_60121865), .B(n_281263079), .C(n_251062777),
		 .D(\nbus_11365[18] ), .Z(n_272362990));
	notech_ao4 i_175646004(.A(n_28108), .B(n_60358), .C(n_251362780), .D(n_56311
		), .Z(n_272162988));
	notech_ao4 i_175746003(.A(n_251162778), .B(n_29773), .C(n_58426), .D(n_28004
		), .Z(n_271962986));
	notech_and3 i_176345997(.A(n_271562982), .B(n_271762984), .C(n_257062837
		), .Z(n_271862985));
	notech_ao4 i_176046000(.A(n_313447724), .B(n_322438019), .C(n_247972959)
		, .D(n_316537960), .Z(n_271762984));
	notech_ao4 i_176145999(.A(n_253773017), .B(n_281263079), .C(n_251062777)
		, .D(n_57707), .Z(n_271562982));
	notech_ao4 i_176445996(.A(n_28109), .B(n_60358), .C(n_250962776), .D(n_57720
		), .Z(n_271362980));
	notech_ao4 i_176545995(.A(n_56320), .B(n_251362780), .C(n_60005), .D(n_251262779
		), .Z(n_271262979));
	notech_and3 i_177045990(.A(n_270862975), .B(n_271062977), .C(n_257862845
		), .Z(n_271162978));
	notech_ao4 i_176745993(.A(n_251162778), .B(n_29775), .C(n_58426), .D(n_28005
		), .Z(n_271062977));
	notech_ao4 i_176845992(.A(n_247072950), .B(n_316537960), .C(n_241572895)
		, .D(n_309721261), .Z(n_270862975));
	notech_ao4 i_177145989(.A(n_60358), .B(n_28110), .C(n_110964638), .D(n_316537960
		), .Z(n_270662973));
	notech_ao4 i_177245988(.A(n_251362780), .B(n_56329), .C(n_60004), .D(n_251262779
		), .Z(n_270462971));
	notech_and3 i_177845982(.A(n_270062967), .B(n_270262969), .C(n_258762854
		), .Z(n_270362970));
	notech_ao4 i_177545985(.A(n_251162778), .B(n_29681), .C(n_58426), .D(n_28006
		), .Z(n_270262969));
	notech_ao4 i_177645984(.A(n_251062777), .B(n_57733), .C(n_249866027), .D
		(n_309721261), .Z(n_270062967));
	notech_and4 i_199645786(.A(n_269762964), .B(n_269562962), .C(n_259062857
		), .D(n_259362860), .Z(n_269962966));
	notech_ao4 i_199245790(.A(\nbus_11358[16] ), .B(n_309091733), .C(n_60009
		), .D(n_122528502), .Z(n_269762964));
	notech_ao4 i_199445788(.A(n_29710), .B(n_26765), .C(n_309191732), .D(n_29776
		), .Z(n_269562962));
	notech_and4 i_200145781(.A(n_269262959), .B(n_269062957), .C(n_259962866
		), .D(n_259662863), .Z(n_269462961));
	notech_ao4 i_199745785(.A(n_121628493), .B(n_28001), .C(n_60162), .D(n_27256
		), .Z(n_269262959));
	notech_ao4 i_199945783(.A(n_313747721), .B(n_124328520), .C(n_252966058)
		, .D(n_309391730), .Z(n_269062957));
	notech_and4 i_202145762(.A(n_268762954), .B(n_268562952), .C(n_260262869
		), .D(n_260562872), .Z(n_268962956));
	notech_ao4 i_201745766(.A(n_309091733), .B(n_56293), .C(n_60008), .D(n_122528502
		), .Z(n_268762954));
	notech_ao4 i_201945764(.A(n_29772), .B(n_26765), .C(n_309191732), .D(n_29779
		), .Z(n_268562952));
	notech_and4 i_202645757(.A(n_268262949), .B(n_268062947), .C(n_261162878
		), .D(n_260862875), .Z(n_268462951));
	notech_ao4 i_202245761(.A(n_121628493), .B(n_28002), .C(n_60122), .D(n_27258
		), .Z(n_268262949));
	notech_ao4 i_202445759(.A(n_313647722), .B(n_124328520), .C(n_245572935)
		, .D(n_309391730), .Z(n_268062947));
	notech_and4 i_206945714(.A(n_267762944), .B(n_267562942), .C(n_261462881
		), .D(n_261762884), .Z(n_267962946));
	notech_ao4 i_206545718(.A(n_309091733), .B(n_56311), .C(n_60006), .D(n_122528502
		), .Z(n_267762944));
	notech_ao4 i_206745716(.A(n_29773), .B(n_26765), .C(n_309191732), .D(n_29780
		), .Z(n_267562942));
	notech_and4 i_207445709(.A(n_267262939), .B(n_267062937), .C(n_262362890
		), .D(n_262062887), .Z(n_267462941));
	notech_ao4 i_207045713(.A(n_121628493), .B(n_28004), .C(n_60122), .D(n_27261
		), .Z(n_267262939));
	notech_ao4 i_207245711(.A(n_313447724), .B(n_124328520), .C(n_243072910)
		, .D(n_309391730), .Z(n_267062937));
	notech_and4 i_209345690(.A(n_266762934), .B(n_266562932), .C(n_262662893
		), .D(n_262962896), .Z(n_266962936));
	notech_ao4 i_208945694(.A(n_309091733), .B(n_56320), .C(n_60005), .D(n_122528502
		), .Z(n_266762934));
	notech_ao4 i_209145692(.A(n_29775), .B(n_26765), .C(n_309191732), .D(n_29784
		), .Z(n_266562932));
	notech_and4 i_209845685(.A(n_266262929), .B(n_266062927), .C(n_263562902
		), .D(n_263262899), .Z(n_266462931));
	notech_ao4 i_209445689(.A(n_121628493), .B(n_28005), .C(n_60122), .D(n_27262
		), .Z(n_266262929));
	notech_ao4 i_209645687(.A(n_313347725), .B(n_124328520), .C(n_241572895)
		, .D(n_309391730), .Z(n_266062927));
	notech_and4 i_211745666(.A(n_265762924), .B(n_265562922), .C(n_263862905
		), .D(n_264162908), .Z(n_265962926));
	notech_ao4 i_211345670(.A(n_309091733), .B(n_56329), .C(n_60004), .D(n_122528502
		), .Z(n_265762924));
	notech_ao4 i_211545668(.A(n_29681), .B(n_26765), .C(n_56091), .D(n_29785
		), .Z(n_265562922));
	notech_and4 i_212245661(.A(n_265262919), .B(n_265062917), .C(n_264762914
		), .D(n_264462911), .Z(n_265462921));
	notech_ao4 i_211845665(.A(n_121628493), .B(n_28006), .C(n_60122), .D(n_27263
		), .Z(n_265262919));
	notech_ao4 i_212045663(.A(n_122628503), .B(n_29553), .C(n_249866027), .D
		(n_309391730), .Z(n_265062917));
	notech_and3 i_7047629(.A(n_56848), .B(n_187762157), .C(n_58486), .Z(n_264862915
		));
	notech_or2 i_111146625(.A(n_59980), .B(n_124328520), .Z(n_264762914));
	notech_nao3 i_111546622(.A(n_19065), .B(read_data[21]), .C(n_59100), .Z(n_264462911
		));
	notech_or2 i_111846619(.A(n_122428501), .B(n_28147), .Z(n_264162908));
	notech_or2 i_112146616(.A(n_308991734), .B(n_57733), .Z(n_263862905));
	notech_nand2 i_108246653(.A(add_len_pc[20]), .B(n_26766), .Z(n_263562902
		));
	notech_nao3 i_108546650(.A(n_19065), .B(read_data[20]), .C(n_59100), .Z(n_263262899
		));
	notech_or2 i_108846647(.A(n_122428501), .B(n_28146), .Z(n_262962896));
	notech_or2 i_109146644(.A(n_308991734), .B(n_57720), .Z(n_262662893));
	notech_nand2 i_105446681(.A(add_len_pc[19]), .B(n_26766), .Z(n_262362890
		));
	notech_nao3 i_105746678(.A(n_19065), .B(read_data[19]), .C(n_59100), .Z(n_262062887
		));
	notech_or2 i_106046675(.A(n_122428501), .B(n_28145), .Z(n_261762884));
	notech_or2 i_106346672(.A(n_308991734), .B(n_57707), .Z(n_261462881));
	notech_nand2 i_99646737(.A(add_len_pc[17]), .B(n_26766), .Z(n_261162878)
		);
	notech_nao3 i_99946734(.A(n_19065), .B(read_data[17]), .C(n_59100), .Z(n_260862875
		));
	notech_or2 i_100246731(.A(n_122428501), .B(n_28143), .Z(n_260562872));
	notech_or2 i_100546728(.A(n_308991734), .B(n_57689), .Z(n_260262869));
	notech_nand2 i_96846765(.A(add_len_pc[16]), .B(n_26766), .Z(n_259962866)
		);
	notech_nao3 i_97146762(.A(n_19065), .B(read_data[16]), .C(n_59100), .Z(n_259662863
		));
	notech_or2 i_97446759(.A(n_122428501), .B(n_28142), .Z(n_259362860));
	notech_or2 i_97746756(.A(n_308991734), .B(\nbus_11365[16] ), .Z(n_259062857
		));
	notech_or2 i_77646948(.A(n_59980), .B(n_322438019), .Z(n_258762854));
	notech_or4 i_78146943(.A(n_62856), .B(n_281263079), .C(n_62808), .D(n_57733
		), .Z(n_258262849));
	notech_or2 i_76746956(.A(n_313347725), .B(n_322438019), .Z(n_257862845)
		);
	notech_or4 i_75846965(.A(n_281263079), .B(nbus_11295[19]), .C(n_60945), 
		.D(n_174962032), .Z(n_257062837));
	notech_or2 i_76346960(.A(n_60006), .B(n_251262779), .Z(n_256562832));
	notech_or4 i_74946974(.A(n_281263079), .B(n_60945), .C(nbus_11295[18]), 
		.D(n_174962032), .Z(n_256162828));
	notech_or2 i_75446969(.A(n_3864), .B(n_251262779), .Z(n_255662823));
	notech_or4 i_74046983(.A(n_281263079), .B(nbus_11295[17]), .C(n_60945), 
		.D(n_174962032), .Z(n_255262819));
	notech_or2 i_74546978(.A(n_60008), .B(n_251262779), .Z(n_254762814));
	notech_or4 i_73146992(.A(n_281263079), .B(nbus_11295[16]), .C(n_60945), 
		.D(n_174962032), .Z(n_254362810));
	notech_or2 i_73646987(.A(n_275963026), .B(\nbus_11358[16] ), .Z(n_253662803
		));
	notech_or4 i_117446563(.A(calc_sz[1]), .B(n_246691943), .C(n_56837), .D(n_32298
		), .Z(n_253162798));
	notech_or4 i_117246565(.A(n_32342), .B(n_32339), .C(n_54756), .D(n_264862915
		), .Z(n_252962796));
	notech_or4 i_116946568(.A(n_30854), .B(n_54727), .C(n_58480), .D(n_60945
		), .Z(n_252762794));
	notech_nand3 i_7647623(.A(n_305391770), .B(n_253162798), .C(n_58504), .Z
		(n_252662793));
	notech_ao4 i_156561747(.A(n_60358), .B(n_28104), .C(n_30565), .D(n_60010
		), .Z(n_115075094));
	notech_ao4 i_156661746(.A(n_30569), .B(\nbus_11358[15] ), .C(n_30568), .D
		(\nbus_11307[15] ), .Z(n_115175095));
	notech_and4 i_3461691(.A(n_59152), .B(n_315391670), .C(n_312391700), .D(n_312770138
		), .Z(n_115275096));
	notech_and2 i_3561690(.A(n_31279), .B(n_119475138), .Z(n_115375097));
	notech_ao3 i_7461654(.A(tsc[15]), .B(n_27855), .C(n_59469), .Z(n_115875102
		));
	notech_or2 i_7361655(.A(n_151028787), .B(nbus_11295[15]), .Z(n_116175105
		));
	notech_nand2 i_7061658(.A(opb[15]), .B(n_58097), .Z(n_116475108));
	notech_nao3 i_24261486(.A(n_319091633), .B(n_246991940), .C(n_269834654)
		, .Z(n_116975113));
	notech_nand2 i_23761491(.A(n_200075939), .B(opa[7]), .Z(n_117675120));
	notech_ao3 i_92260838(.A(n_62826), .B(opc[30]), .C(n_58082), .Z(n_117975123
		));
	notech_or2 i_91760843(.A(n_321538010), .B(n_303091793), .Z(n_118675130)
		);
	notech_ao4 i_202559811(.A(n_321438009), .B(n_28015), .C(n_319937994), .D
		(n_30809), .Z(n_118775131));
	notech_ao4 i_202459812(.A(n_302991794), .B(n_58145), .C(\nbus_11365[30] 
		), .D(n_57869), .Z(n_118975133));
	notech_nand3 i_202759809(.A(n_118775131), .B(n_118975133), .C(n_118675130
		), .Z(n_119075134));
	notech_ao4 i_202259814(.A(n_29591), .B(n_26918), .C(n_57873), .D(\nbus_11358[30] 
		), .Z(n_119175135));
	notech_ao4 i_142960372(.A(n_29614), .B(n_315191672), .C(n_303191792), .D
		(n_24996), .Z(n_119475138));
	notech_ao4 i_142660375(.A(n_24994), .B(n_115375097), .C(\nbus_11358[7] )
		, .D(n_115275096), .Z(n_119575139));
	notech_ao4 i_142560376(.A(n_31307), .B(n_306170072), .C(n_58410), .D(n_27990
		), .Z(n_119775141));
	notech_ao4 i_142360378(.A(n_54643), .B(n_28967), .C(n_31309), .D(n_306270073
		), .Z(n_119975143));
	notech_and3 i_142460377(.A(n_116975113), .B(n_119975143), .C(n_26708), .Z
		(n_120175145));
	notech_ao4 i_126560530(.A(n_111064639), .B(n_312970140), .C(n_26925), .D
		(n_320538000), .Z(n_120275146));
	notech_ao4 i_126460531(.A(\nbus_11307[15] ), .B(n_26819), .C(n_23512), .D
		(n_58622), .Z(n_120375147));
	notech_ao4 i_126260533(.A(n_60010), .B(n_316691657), .C(n_121675160), .D
		(n_29754), .Z(n_120575149));
	notech_and4 i_126760528(.A(n_120575149), .B(n_120375147), .C(n_120275146
		), .D(n_116475108), .Z(n_120775151));
	notech_ao4 i_125960536(.A(n_298466513), .B(n_319670207), .C(n_28000), .D
		(n_58408), .Z(n_120875152));
	notech_ao3 i_125860537(.A(n_115175095), .B(n_115075094), .C(n_115875102)
		, .Z(n_121175155));
	notech_nand3 i_65858480(.A(n_138375327), .B(n_138575329), .C(n_138175325
		), .Z(n_121375157));
	notech_and4 i_17558318(.A(n_58530), .B(n_316691657), .C(n_311191712), .D
		(n_124675190), .Z(n_121475158));
	notech_and2 i_17258321(.A(n_31279), .B(n_147275416), .Z(n_121575159));
	notech_ao4 i_141458499(.A(n_30594), .B(n_60229), .C(n_319891625), .D(n_23512
		), .Z(n_121675160));
	notech_and2 i_17158322(.A(n_31456), .B(n_144075384), .Z(n_121775161));
	notech_mux2 i_12358369(.S(n_32323), .A(n_29596), .B(n_302491799), .Z(n_121875162
		));
	notech_or2 i_12258370(.A(n_39370), .B(n_26938), .Z(n_122175165));
	notech_nand2 i_16758326(.A(n_58514), .B(n_122375167), .Z(n_122275166));
	notech_nao3 i_33758157(.A(n_57976), .B(n_27221), .C(n_26697), .Z(n_122375167
		));
	notech_ao4 i_16558328(.A(n_183858934), .B(\nbus_11307[7] ), .C(n_26060),
		 .D(\nbus_11358[7] ), .Z(n_122475168));
	notech_and3 i_16658327(.A(n_3858), .B(n_25884), .C(n_137275316), .Z(n_122575169
		));
	notech_nao3 i_104057487(.A(n_60845), .B(n_27177), .C(n_56516), .Z(n_122975173
		));
	notech_or4 i_19358300(.A(n_32326), .B(n_32343), .C(n_23513), .D(n_317591648
		), .Z(n_124675190));
	notech_or2 i_23558258(.A(n_151028787), .B(nbus_11295[4]), .Z(n_126075204
		));
	notech_or2 i_24458249(.A(n_151028787), .B(nbus_11295[7]), .Z(n_127375217
		));
	notech_nao3 i_24358250(.A(tsc[7]), .B(n_27855), .C(n_59469), .Z(n_127675220
		));
	notech_or4 i_23858255(.A(n_56516), .B(n_60945), .C(nbus_11295[7]), .D(n_26942
		), .Z(n_128175225));
	notech_or2 i_25358240(.A(n_58408), .B(n_27992), .Z(n_129075234));
	notech_ao3 i_26858225(.A(tsc[10]), .B(n_55820), .C(n_59469), .Z(n_129575239
		));
	notech_or4 i_26758226(.A(n_60945), .B(n_28136), .C(n_26942), .D(n_23512)
		, .Z(n_129875242));
	notech_or4 i_26458229(.A(n_62856), .B(n_62808), .C(n_29684), .D(n_23512)
		, .Z(n_130175245));
	notech_nao3 i_27758216(.A(tsc[11]), .B(n_55820), .C(n_59469), .Z(n_130675250
		));
	notech_nao3 i_27658217(.A(n_62826), .B(opc[11]), .C(n_312970140), .Z(n_130975253
		));
	notech_nand2 i_27158222(.A(opb[11]), .B(n_58097), .Z(n_131475258));
	notech_nao3 i_32358170(.A(n_26939), .B(n_122175165), .C(n_175062033), .Z
		(n_132875272));
	notech_nand2 i_32458169(.A(opa[0]), .B(n_122275166), .Z(n_132975273));
	notech_or4 i_34758147(.A(n_56837), .B(n_26610), .C(n_59992), .D(n_56527)
		, .Z(n_133475278));
	notech_or4 i_34458150(.A(n_62856), .B(n_26697), .C(n_62808), .D(\nbus_11307[1] 
		), .Z(n_133775281));
	notech_or4 i_42758067(.A(n_62864), .B(n_147871958), .C(n_60945), .D(\nbus_11307[1] 
		), .Z(n_134275286));
	notech_or4 i_42658068(.A(n_56837), .B(n_26610), .C(n_26928), .D(n_59992)
		, .Z(n_134575289));
	notech_or4 i_42358071(.A(n_62854), .B(n_58163), .C(n_62780), .D(\nbus_11307[1] 
		), .Z(n_134875292));
	notech_or4 i_43658058(.A(n_26767), .B(n_3853), .C(n_28128), .D(n_60945),
		 .Z(n_135775301));
	notech_nao3 i_43358061(.A(n_58078), .B(opd[4]), .C(n_56601), .Z(n_136075304
		));
	notech_or2 i_43058064(.A(n_57980), .B(\nbus_11358[4] ), .Z(n_136375307)
		);
	notech_or4 i_44658048(.A(n_26767), .B(n_3853), .C(n_60945), .D(n_28133),
		 .Z(n_136475308));
	notech_nao3 i_44158053(.A(n_27029), .B(\opa_12[7] ), .C(n_3853), .Z(n_137175315
		));
	notech_or4 i_44958045(.A(n_26062), .B(n_29652), .C(n_29658), .D(n_26055)
		, .Z(n_137275316));
	notech_or2 i_9458397(.A(n_56516), .B(n_23510), .Z(n_137375317));
	notech_or4 i_8858403(.A(n_26062), .B(n_56516), .C(n_57088), .D(instrc[
		116]), .Z(n_137475318));
	notech_or4 i_8758404(.A(n_26062), .B(n_23514), .C(n_57088), .D(instrc[
		116]), .Z(n_137575319));
	notech_nand2 i_11358378(.A(n_27029), .B(n_27023), .Z(n_137675320));
	notech_nand2 i_102857499(.A(read_data[7]), .B(n_60229), .Z(n_138175325)
		);
	notech_ao4 i_190756643(.A(n_58391), .B(n_29614), .C(n_58432), .D(n_303191792
		), .Z(n_138375327));
	notech_ao4 i_190656644(.A(n_58514), .B(\nbus_11307[7] ), .C(n_58530), .D
		(\nbus_11358[7] ), .Z(n_138575329));
	notech_ao4 i_131957220(.A(n_31307), .B(n_122575169), .C(n_58163), .D(n_122475168
		), .Z(n_138775331));
	notech_ao4 i_131857221(.A(n_3857), .B(n_56100), .C(n_56601), .D(n_57947)
		, .Z(n_138975333));
	notech_ao4 i_131657223(.A(n_31279), .B(n_3853), .C(n_303191792), .D(n_154175485
		), .Z(n_139175335));
	notech_and3 i_131757222(.A(n_136475308), .B(n_139175335), .C(n_26708), .Z
		(n_139375337));
	notech_ao4 i_131257227(.A(n_137675320), .B(n_29725), .C(n_142971909), .D
		(\nbus_11307[4] ), .Z(n_139475338));
	notech_ao4 i_130957229(.A(n_3853), .B(n_291463181), .C(n_5743), .D(n_154175485
		), .Z(n_139675340));
	notech_and4 i_131457225(.A(n_139675340), .B(n_139475338), .C(n_136075304
		), .D(n_136375307), .Z(n_139875342));
	notech_ao4 i_130657232(.A(n_291763184), .B(n_147771957), .C(n_58163), .D
		(n_291563182), .Z(n_139975343));
	notech_ao4 i_130457234(.A(n_291663183), .B(n_147871958), .C(n_147671956)
		, .D(n_5723), .Z(n_140175345));
	notech_and4 i_130857230(.A(n_181462097), .B(n_140175345), .C(n_135775301
		), .D(n_139975343), .Z(n_140375347));
	notech_ao4 i_130157237(.A(n_137675320), .B(n_29678), .C(n_142971909), .D
		(\nbus_11307[1] ), .Z(n_140475348));
	notech_ao4 i_130057238(.A(n_60024), .B(n_154175485), .C(n_57980), .D(\nbus_11358[1] 
		), .Z(n_140575349));
	notech_ao4 i_129857240(.A(n_147571955), .B(n_27983), .C(n_297666505), .D
		(n_3853), .Z(n_140775351));
	notech_and4 i_130357235(.A(n_140775351), .B(n_140575349), .C(n_140475348
		), .D(n_134875292), .Z(n_140975353));
	notech_ao4 i_129557243(.A(n_298066509), .B(n_57922), .C(n_147771957), .D
		(n_297966508), .Z(n_141075354));
	notech_and4 i_129257244(.A(n_229779798), .B(n_134275286), .C(n_125828535
		), .D(n_229679797), .Z(n_141375357));
	notech_ao4 i_122257312(.A(n_60024), .B(n_57619), .C(n_57882), .D(\nbus_11358[1] 
		), .Z(n_141575359));
	notech_ao4 i_122157313(.A(n_57891), .B(\nbus_11307[1] ), .C(n_57938), .D
		(n_29678), .Z(n_141675360));
	notech_ao4 i_121957315(.A(n_58410), .B(n_27983), .C(n_297666505), .D(n_24994
		), .Z(n_141875362));
	notech_and4 i_122457310(.A(n_141875362), .B(n_141675360), .C(n_141575359
		), .D(n_133775281), .Z(n_142075364));
	notech_ao4 i_121557318(.A(n_298066509), .B(n_306270073), .C(n_297966508)
		, .D(n_306170072), .Z(n_142175365));
	notech_ao4 i_121357320(.A(n_54643), .B(n_28962), .C(n_305970070), .D(n_297866507
		), .Z(n_142375367));
	notech_and4 i_121857316(.A(n_276234718), .B(n_142375367), .C(n_142175365
		), .D(n_133475278), .Z(n_142575369));
	notech_ao4 i_120857325(.A(n_58410), .B(n_27981), .C(n_24994), .D(n_58610
		), .Z(n_142875372));
	notech_and3 i_121057323(.A(n_142875372), .B(n_132975273), .C(n_132875272
		), .Z(n_142975373));
	notech_ao4 i_120657327(.A(n_60025), .B(n_57619), .C(n_199975938), .D(n_29742
		), .Z(n_143075374));
	notech_ao4 i_120557328(.A(n_291363180), .B(n_306070071), .C(n_311791706)
		, .D(n_59993), .Z(n_143175375));
	notech_ao4 i_120257331(.A(n_291263179), .B(n_306170072), .C(n_291163178)
		, .D(n_306270073), .Z(n_143475378));
	notech_ao4 i_120157332(.A(n_54643), .B(n_28961), .C(n_57882), .D(\nbus_11358[0] 
		), .Z(n_143575379));
	notech_ao4 i_119857334(.A(n_60358), .B(n_28089), .C(n_26697), .D(n_58646
		), .Z(n_143775381));
	notech_and4 i_120457329(.A(n_125828535), .B(n_143775381), .C(n_143575379
		), .D(n_143475378), .Z(n_143975383));
	notech_ao4 i_115957371(.A(n_31492), .B(n_23510), .C(n_317591648), .D(n_121875162
		), .Z(n_144075384));
	notech_ao4 i_115557374(.A(n_26819), .B(\nbus_11307[11] ), .C(n_23512), .D
		(n_121775161), .Z(n_144175385));
	notech_ao4 i_115457375(.A(n_30528), .B(n_26925), .C(n_58408), .D(n_27996
		), .Z(n_144375387));
	notech_ao4 i_115157378(.A(n_31476), .B(n_319670207), .C(n_151028787), .D
		(nbus_11295[11]), .Z(n_144575389));
	notech_and4 i_115357376(.A(n_187368889), .B(n_144575389), .C(n_130675250
		), .D(n_130975253), .Z(n_144875392));
	notech_ao4 i_114757382(.A(n_87532846), .B(n_312970140), .C(n_187568890),
		 .D(n_56579), .Z(n_144975393));
	notech_ao4 i_114657383(.A(n_29684), .B(n_57415), .C(n_3850), .D(n_316691657
		), .Z(n_145075394));
	notech_ao4 i_114457385(.A(\nbus_11358[10] ), .B(n_26820), .C(\nbus_11307[10] 
		), .D(n_26819), .Z(n_145275396));
	notech_and4 i_114957380(.A(n_145275396), .B(n_145075394), .C(n_144975393
		), .D(n_130175245), .Z(n_145475398));
	notech_ao4 i_114157388(.A(n_151028787), .B(nbus_11295[10]), .C(n_58408),
		 .D(n_27993), .Z(n_145575399));
	notech_ao3 i_114057389(.A(n_3849), .B(n_187968894), .C(n_129575239), .Z(n_145875402
		));
	notech_ao4 i_113657393(.A(n_208969101), .B(n_56579), .C(n_121675160), .D
		(n_29743), .Z(n_146075404));
	notech_ao4 i_113557394(.A(n_60016), .B(n_316691657), .C(\nbus_11307[9] )
		, .D(n_26819), .Z(n_146175405));
	notech_ao4 i_113357396(.A(n_58608), .B(n_23512), .C(\nbus_11358[9] ), .D
		(n_26820), .Z(n_146375407));
	notech_and4 i_113857391(.A(n_146375407), .B(n_146175405), .C(n_146075404
		), .D(n_129075234), .Z(n_146575409));
	notech_ao4 i_113057399(.A(n_189962171), .B(n_312970140), .C(n_291963186)
		, .D(n_319670207), .Z(n_146675410));
	notech_ao4 i_112957400(.A(n_59124), .B(nbus_11295[9]), .C(n_54643), .D(n_28951
		), .Z(n_146775411));
	notech_and3 i_112857401(.A(n_207569087), .B(n_207469086), .C(n_3849), .Z
		(n_147075414));
	notech_ao4 i_112657403(.A(n_319891625), .B(n_29614), .C(n_23507), .D(n_303191792
		), .Z(n_147275416));
	notech_ao4 i_112357406(.A(n_56579), .B(n_269834654), .C(n_23514), .D(n_121575159
		), .Z(n_147375417));
	notech_ao4 i_112257407(.A(n_58411), .B(n_56100), .C(n_31309), .D(n_137575319
		), .Z(n_147575419));
	notech_ao4 i_111957410(.A(\nbus_11307[7] ), .B(n_26699), .C(\nbus_11358[7] 
		), .D(n_215476093), .Z(n_147775421));
	notech_and4 i_112157408(.A(n_147775421), .B(n_26708), .C(n_127375217), .D
		(n_127675220), .Z(n_148075424));
	notech_ao4 i_111557414(.A(n_291663183), .B(n_137375317), .C(n_57892), .D
		(\nbus_11307[4] ), .Z(n_148175425));
	notech_ao4 i_111457415(.A(n_291863185), .B(n_137575319), .C(n_291763184)
		, .D(n_137475318), .Z(n_148275426));
	notech_ao4 i_111257417(.A(n_5743), .B(n_199875937), .C(n_56516), .D(n_291563182
		), .Z(n_148475428));
	notech_ao4 i_111157418(.A(n_199575934), .B(n_29725), .C(n_57893), .D(\nbus_11358[4] 
		), .Z(n_148575429));
	notech_and4 i_111757412(.A(n_148575429), .B(n_148475428), .C(n_148275426
		), .D(n_148175425), .Z(n_148775431));
	notech_ao4 i_110757421(.A(n_5723), .B(n_315691667), .C(n_58411), .D(n_27986
		), .Z(n_148875432));
	notech_ao4 i_110657422(.A(n_54643), .B(n_28947), .C(n_291463181), .D(n_23514
		), .Z(n_148975433));
	notech_and3 i_110557423(.A(n_3849), .B(n_276134717), .C(n_126075204), .Z
		(n_149275436));
	notech_ao4 i_108657441(.A(n_297866507), .B(n_137375317), .C(n_57892), .D
		(\nbus_11307[1] ), .Z(n_149475438));
	notech_ao4 i_108557442(.A(n_298066509), .B(n_137575319), .C(n_297966508)
		, .D(n_137475318), .Z(n_149575439));
	notech_ao4 i_108357444(.A(n_60024), .B(n_199875937), .C(n_297766506), .D
		(n_56516), .Z(n_149775441));
	notech_ao4 i_108257445(.A(n_199575934), .B(n_29678), .C(n_57893), .D(\nbus_11358[1] 
		), .Z(n_149875442));
	notech_and4 i_108857439(.A(n_149875442), .B(n_149775441), .C(n_149575439
		), .D(n_149475438), .Z(n_150075444));
	notech_ao4 i_107957448(.A(n_59992), .B(n_315691667), .C(n_58411), .D(n_27983
		), .Z(n_150175445));
	notech_ao4 i_107857449(.A(n_54638), .B(n_28944), .C(n_297666505), .D(n_23514
		), .Z(n_150275446));
	notech_ao4 i_107657451(.A(n_3867), .B(n_3596), .C(n_59124), .D(nbus_11295
		[1]), .Z(n_150475448));
	notech_and4 i_108157446(.A(n_150475448), .B(n_150275446), .C(n_150175445
		), .D(n_276234718), .Z(n_150675450));
	notech_ao4 i_107257455(.A(\nbus_11307[0] ), .B(n_57892), .C(n_121475158)
		, .D(\nbus_11358[0] ), .Z(n_150875452));
	notech_ao4 i_107157456(.A(n_175062033), .B(n_137375317), .C(n_142871908)
		, .D(n_291363180), .Z(n_150975453));
	notech_ao4 i_106957458(.A(n_291163178), .B(n_137575319), .C(n_291263179)
		, .D(n_137475318), .Z(n_151175455));
	notech_ao4 i_106857459(.A(n_60025), .B(n_199875937), .C(n_56516), .D(n_58646
		), .Z(n_151275456));
	notech_and4 i_107457453(.A(n_151275456), .B(n_151175455), .C(n_150975453
		), .D(n_150875452), .Z(n_151475458));
	notech_ao4 i_106557462(.A(n_59993), .B(n_315691667), .C(n_27981), .D(n_58411
		), .Z(n_151575459));
	notech_ao4 i_106457463(.A(n_199775936), .B(n_29742), .C(n_23514), .D(n_58610
		), .Z(n_151675460));
	notech_ao4 i_106257465(.A(n_59124), .B(nbus_11295[0]), .C(n_54638), .D(n_28943
		), .Z(n_151875462));
	notech_and3 i_106357464(.A(n_3867), .B(n_151875462), .C(n_57548), .Z(n_152075464
		));
	notech_ao3 i_78755519(.A(n_154275486), .B(n_154475488), .C(n_154075484),
		 .Z(n_152275466));
	notech_ao4 i_10555412(.A(n_3853), .B(n_29742), .C(n_58163), .D(\nbus_11307[0] 
		), .Z(n_152375467));
	notech_or4 i_32755197(.A(n_62864), .B(n_62808), .C(n_29742), .D(n_3853),
		 .Z(n_152675470));
	notech_ao3 i_32655198(.A(n_59445), .B(opa[0]), .C(n_58163), .Z(n_152975473
		));
	notech_or4 i_32355201(.A(n_3854), .B(n_3853), .C(n_60025), .D(n_58020), 
		.Z(n_153275476));
	notech_nor2 i_45155074(.A(n_60025), .B(n_58432), .Z(n_154075484));
	notech_or4 i_34137(.A(n_32614), .B(n_32342), .C(n_3854), .D(n_3853), .Z(n_154175485
		));
	notech_ao4 i_94654639(.A(n_58530), .B(\nbus_11358[0] ), .C(n_147071950),
		 .D(\nbus_11307[0] ), .Z(n_154275486));
	notech_ao4 i_94554640(.A(n_60358), .B(n_28089), .C(n_58391), .D(n_29742)
		, .Z(n_154475488));
	notech_ao4 i_71554846(.A(n_146971949), .B(n_291363180), .C(n_152375467),
		 .D(n_3844), .Z(n_154575489));
	notech_ao4 i_71454847(.A(n_147671956), .B(n_59993), .C(n_147571955), .D(n_27981
		), .Z(n_154675490));
	notech_ao4 i_71254849(.A(n_147871958), .B(n_175062033), .C(n_147771957),
		 .D(n_291263179), .Z(n_154875492));
	notech_and4 i_71754844(.A(n_153275476), .B(n_154875492), .C(n_154675490)
		, .D(n_154575489), .Z(n_155075494));
	notech_ao4 i_70954852(.A(n_57980), .B(\nbus_11358[0] ), .C(n_291163178),
		 .D(n_57922), .Z(n_155175495));
	notech_nand3 i_70854853(.A(n_152275466), .B(n_125828535), .C(n_152675470
		), .Z(n_155475498));
	notech_or2 i_25650412(.A(n_3878), .B(\nbus_11365[22] ), .Z(n_156475508)
		);
	notech_or2 i_25150417(.A(n_289227274), .B(n_3837), .Z(n_156975513));
	notech_nor2 i_26450404(.A(n_3878), .B(\nbus_11365[23] ), .Z(n_157075514)
		);
	notech_or2 i_25950409(.A(n_289127273), .B(n_3837), .Z(n_157775521));
	notech_nor2 i_38150287(.A(n_57868), .B(\nbus_11365[23] ), .Z(n_157875522
		));
	notech_or2 i_37650292(.A(n_154831963), .B(n_289127273), .Z(n_158575529)
		);
	notech_nor2 i_38950279(.A(n_57868), .B(\nbus_11365[24] ), .Z(n_158675530
		));
	notech_or2 i_38450284(.A(n_289027272), .B(n_154831963), .Z(n_159375537)
		);
	notech_nor2 i_59950080(.A(n_57869), .B(\nbus_11365[22] ), .Z(n_159475538
		));
	notech_or2 i_59450085(.A(n_289227274), .B(n_321538010), .Z(n_160175545)
		);
	notech_nor2 i_60750072(.A(n_57869), .B(\nbus_11365[23] ), .Z(n_160275546
		));
	notech_or2 i_60250077(.A(n_289127273), .B(n_321538010), .Z(n_160975553)
		);
	notech_nor2 i_61550064(.A(n_57869), .B(\nbus_11365[24] ), .Z(n_161075554
		));
	notech_or2 i_61050069(.A(n_289027272), .B(n_321538010), .Z(n_161775561)
		);
	notech_or2 i_63250047(.A(n_154331958), .B(nbus_11295[22]), .Z(n_161875562
		));
	notech_or2 i_63150048(.A(n_57870), .B(\nbus_11365[22] ), .Z(n_162175565)
		);
	notech_or2 i_62650053(.A(n_305924323), .B(n_289227274), .Z(n_162675570)
		);
	notech_or2 i_64150038(.A(n_154331958), .B(nbus_11295[23]), .Z(n_162775571
		));
	notech_or2 i_64050039(.A(n_57870), .B(\nbus_11365[23] ), .Z(n_163075574)
		);
	notech_or2 i_63550044(.A(n_305924323), .B(n_289127273), .Z(n_163575579)
		);
	notech_or2 i_65050029(.A(n_154331958), .B(nbus_11295[24]), .Z(n_163675580
		));
	notech_or2 i_64950030(.A(n_57870), .B(\nbus_11365[24] ), .Z(n_163975583)
		);
	notech_or2 i_64450035(.A(n_305924323), .B(n_289027272), .Z(n_164475588)
		);
	notech_nor2 i_73449952(.A(n_314047718), .B(\nbus_11365[22] ), .Z(n_164575589
		));
	notech_or2 i_72949957(.A(n_306824332), .B(n_289227274), .Z(n_165275596)
		);
	notech_nor2 i_74249944(.A(n_314047718), .B(\nbus_11365[23] ), .Z(n_165375597
		));
	notech_or2 i_73749949(.A(n_306824332), .B(n_289127273), .Z(n_166075604)
		);
	notech_nor2 i_75049936(.A(n_314047718), .B(\nbus_11365[24] ), .Z(n_166175605
		));
	notech_or2 i_74549941(.A(n_306824332), .B(n_289027272), .Z(n_166875612)
		);
	notech_ao3 i_80949878(.A(n_32304), .B(opd[23]), .C(n_56684), .Z(n_166975613
		));
	notech_nand2 i_80449883(.A(n_287027252), .B(\regs_13_14[23] ), .Z(n_167675620
		));
	notech_or2 i_84449843(.A(n_57867), .B(\nbus_11365[22] ), .Z(n_167775621)
		);
	notech_or2 i_84349844(.A(n_57865), .B(\nbus_11358[22] ), .Z(n_168075624)
		);
	notech_or2 i_83849849(.A(n_305624320), .B(n_289227274), .Z(n_168575629)
		);
	notech_or2 i_87049817(.A(n_57867), .B(\nbus_11365[24] ), .Z(n_168675630)
		);
	notech_or2 i_86949818(.A(n_57865), .B(\nbus_11358[24] ), .Z(n_168975633)
		);
	notech_or2 i_86449823(.A(n_305624320), .B(n_289027272), .Z(n_169475638)
		);
	notech_or2 i_91649773(.A(n_308991734), .B(\nbus_11365[22] ), .Z(n_169775641
		));
	notech_or2 i_91349776(.A(n_122428501), .B(n_28148), .Z(n_170075644));
	notech_nao3 i_91049779(.A(n_19065), .B(read_data[22]), .C(n_59100), .Z(n_170375647
		));
	notech_nand2 i_90749782(.A(add_len_pc[22]), .B(n_26766), .Z(n_170675650)
		);
	notech_or2 i_94449745(.A(n_308991734), .B(n_57751), .Z(n_170975653));
	notech_or2 i_94149748(.A(n_122428501), .B(n_28149), .Z(n_171275656));
	notech_nao3 i_93849751(.A(n_19065), .B(read_data[23]), .C(n_59100), .Z(n_171575659
		));
	notech_nand2 i_93549754(.A(add_len_pc[23]), .B(n_26766), .Z(n_171875662)
		);
	notech_or2 i_97349717(.A(n_308991734), .B(n_57761), .Z(n_172175665));
	notech_or2 i_97049720(.A(n_122428501), .B(n_28150), .Z(n_172475668));
	notech_nao3 i_96749723(.A(n_19065), .B(read_data[24]), .C(n_59100), .Z(n_172775671
		));
	notech_nand2 i_96449726(.A(add_len_pc[24]), .B(n_26766), .Z(n_173075674)
		);
	notech_ao4 i_186848841(.A(n_124328520), .B(n_289027272), .C(n_309391730)
		, .D(n_221065739), .Z(n_173175675));
	notech_ao4 i_186648843(.A(n_121628493), .B(n_28009), .C(n_60122), .D(n_27266
		), .Z(n_173375677));
	notech_and4 i_187048839(.A(n_173375677), .B(n_173175675), .C(n_173075674
		), .D(n_172775671), .Z(n_173575679));
	notech_ao4 i_186348846(.A(n_26765), .B(n_29769), .C(n_56091), .D(n_29952
		), .Z(n_173675680));
	notech_ao4 i_186148848(.A(n_309091733), .B(\nbus_11358[24] ), .C(n_122528502
		), .D(n_60001), .Z(n_173875682));
	notech_and4 i_186548844(.A(n_173875682), .B(n_173675680), .C(n_172175665
		), .D(n_172475668), .Z(n_174075684));
	notech_ao4 i_184448865(.A(n_124328520), .B(n_289127273), .C(n_309391730)
		, .D(n_222565754), .Z(n_174175685));
	notech_ao4 i_184148867(.A(n_121628493), .B(n_28008), .C(n_60122), .D(n_27265
		), .Z(n_174375687));
	notech_and4 i_184648863(.A(n_174375687), .B(n_174175685), .C(n_171875662
		), .D(n_171575659), .Z(n_174575689));
	notech_ao4 i_183848870(.A(n_26765), .B(n_29765), .C(n_56091), .D(n_29951
		), .Z(n_174675690));
	notech_ao4 i_183648872(.A(n_309091733), .B(\nbus_11358[23] ), .C(n_122528502
		), .D(n_60002), .Z(n_174875692));
	notech_and4 i_184048868(.A(n_174875692), .B(n_174675690), .C(n_170975653
		), .D(n_171275656), .Z(n_175075694));
	notech_ao4 i_181948889(.A(n_124328520), .B(n_289227274), .C(n_309391730)
		, .D(n_224065769), .Z(n_175175695));
	notech_ao4 i_181748891(.A(n_121628493), .B(n_28007), .C(n_60122), .D(n_27264
		), .Z(n_175375697));
	notech_and4 i_182148887(.A(n_175375697), .B(n_175175695), .C(n_170675650
		), .D(n_170375647), .Z(n_175575699));
	notech_ao4 i_181448894(.A(n_26765), .B(n_29708), .C(n_56091), .D(n_29950
		), .Z(n_175675700));
	notech_ao4 i_181248896(.A(n_309091733), .B(\nbus_11358[22] ), .C(n_122528502
		), .D(n_60003), .Z(n_175875702));
	notech_and4 i_181648892(.A(n_175875702), .B(n_175675700), .C(n_169775641
		), .D(n_170075644), .Z(n_176075704));
	notech_ao4 i_178448924(.A(n_58007), .B(n_225565784), .C(n_58008), .D(n_221065739
		), .Z(n_176175705));
	notech_ao4 i_178348925(.A(n_26937), .B(n_29769), .C(n_58423), .D(n_28009
		), .Z(n_176375707));
	notech_ao4 i_178048928(.A(n_58138), .B(n_60001), .C(n_57726), .D(n_28150
		), .Z(n_176575709));
	notech_and4 i_178248926(.A(n_176575709), .B(n_26619), .C(n_168675630), .D
		(n_168975633), .Z(n_176875712));
	notech_ao4 i_176148946(.A(n_58007), .B(n_225765786), .C(n_58008), .D(n_224065769
		), .Z(n_176975713));
	notech_ao4 i_176048947(.A(n_26937), .B(n_29708), .C(n_58423), .D(n_28007
		), .Z(n_177175715));
	notech_ao4 i_175748950(.A(n_58138), .B(n_60003), .C(n_57726), .D(n_28148
		), .Z(n_177375717));
	notech_and4 i_175948948(.A(n_177375717), .B(n_167775621), .C(n_168075624
		), .D(n_26617), .Z(n_177675720));
	notech_ao4 i_173048977(.A(n_286927251), .B(n_222565754), .C(n_286827250)
		, .D(n_225665785), .Z(n_177775721));
	notech_ao4 i_172948978(.A(n_57861), .B(n_57751), .C(n_287827260), .D(n_289127273
		), .Z(n_177975723));
	notech_nand3 i_173248975(.A(n_177775721), .B(n_177975723), .C(n_167675620
		), .Z(n_178075724));
	notech_ao4 i_172748980(.A(n_58139), .B(n_60002), .C(n_57863), .D(\nbus_11358[23] 
		), .Z(n_178175725));
	notech_ao4 i_162549081(.A(n_306624330), .B(n_225565784), .C(n_307124335)
		, .D(n_221065739), .Z(n_178475728));
	notech_ao4 i_162449082(.A(n_307324337), .B(n_29769), .C(n_58425), .D(n_28009
		), .Z(n_178675730));
	notech_nand3 i_162749079(.A(n_178475728), .B(n_178675730), .C(n_166875612
		), .Z(n_178775731));
	notech_ao4 i_162249084(.A(n_57864), .B(\nbus_11358[24] ), .C(n_58141), .D
		(n_60001), .Z(n_178875732));
	notech_ao4 i_161849088(.A(n_306624330), .B(n_225665785), .C(n_307124335)
		, .D(n_222565754), .Z(n_179175735));
	notech_ao4 i_161749089(.A(n_307324337), .B(n_29765), .C(n_58425), .D(n_28008
		), .Z(n_179375737));
	notech_nand3 i_162049086(.A(n_179175735), .B(n_179375737), .C(n_166075604
		), .Z(n_179475738));
	notech_ao4 i_161549091(.A(n_57864), .B(\nbus_11358[23] ), .C(n_58141), .D
		(n_60002), .Z(n_179575739));
	notech_ao4 i_161149095(.A(n_306624330), .B(n_225765786), .C(n_307124335)
		, .D(n_224065769), .Z(n_179875742));
	notech_ao4 i_161049096(.A(n_307324337), .B(n_29708), .C(n_58425), .D(n_28007
		), .Z(n_180075744));
	notech_nand3 i_161349093(.A(n_179875742), .B(n_180075744), .C(n_165275596
		), .Z(n_180175745));
	notech_ao4 i_160849098(.A(n_57864), .B(\nbus_11358[22] ), .C(n_58141), .D
		(n_60003), .Z(n_180275746));
	notech_ao4 i_154749157(.A(n_306124325), .B(n_225565784), .C(n_58085), .D
		(n_221065739), .Z(n_180575749));
	notech_ao4 i_154649158(.A(n_26902), .B(n_29769), .C(n_58427), .D(n_28009
		), .Z(n_180775751));
	notech_ao4 i_154349161(.A(n_57877), .B(\nbus_11358[24] ), .C(n_58143), .D
		(n_60001), .Z(n_180975753));
	notech_and4 i_154549159(.A(n_180975753), .B(n_26619), .C(n_163675580), .D
		(n_163975583), .Z(n_181275756));
	notech_ao4 i_153949165(.A(n_306124325), .B(n_225665785), .C(n_58085), .D
		(n_222565754), .Z(n_181375757));
	notech_ao4 i_153849166(.A(n_26902), .B(n_29765), .C(n_58427), .D(n_28008
		), .Z(n_181575759));
	notech_ao4 i_153549169(.A(n_57877), .B(\nbus_11358[23] ), .C(n_58143), .D
		(n_60002), .Z(n_181775761));
	notech_and4 i_153749167(.A(n_181775761), .B(n_26618), .C(n_162775571), .D
		(n_163075574), .Z(n_182075764));
	notech_ao4 i_153149173(.A(n_306124325), .B(n_225765786), .C(n_58085), .D
		(n_224065769), .Z(n_182175765));
	notech_ao4 i_153049174(.A(n_26902), .B(n_29708), .C(n_58427), .D(n_28007
		), .Z(n_182375767));
	notech_ao4 i_152749177(.A(n_57877), .B(\nbus_11358[22] ), .C(n_58143), .D
		(n_60003), .Z(n_182575769));
	notech_and4 i_152949175(.A(n_182575769), .B(n_26617), .C(n_161875562), .D
		(n_162175565), .Z(n_182875772));
	notech_ao4 i_151649188(.A(n_225565784), .B(n_319937994), .C(n_221065739)
		, .D(n_58082), .Z(n_182975773));
	notech_ao4 i_151549189(.A(n_29769), .B(n_26918), .C(n_321438009), .D(n_28009
		), .Z(n_183175775));
	notech_nand3 i_151849186(.A(n_182975773), .B(n_183175775), .C(n_161775561
		), .Z(n_183275776));
	notech_ao4 i_151349191(.A(n_57873), .B(\nbus_11358[24] ), .C(n_60001), .D
		(n_58145), .Z(n_183375777));
	notech_ao4 i_150949195(.A(n_225665785), .B(n_319937994), .C(n_222565754)
		, .D(n_58082), .Z(n_183675780));
	notech_ao4 i_150849196(.A(n_29765), .B(n_26918), .C(n_321438009), .D(n_28008
		), .Z(n_183875782));
	notech_nand3 i_151149193(.A(n_183675780), .B(n_183875782), .C(n_160975553
		), .Z(n_183975783));
	notech_ao4 i_150649198(.A(n_57873), .B(\nbus_11358[23] ), .C(n_60002), .D
		(n_58145), .Z(n_184075784));
	notech_ao4 i_150249202(.A(n_225765786), .B(n_319937994), .C(n_224065769)
		, .D(n_58082), .Z(n_184375787));
	notech_ao4 i_150149203(.A(n_29708), .B(n_26918), .C(n_321438009), .D(n_28007
		), .Z(n_184575789));
	notech_nand3 i_150449200(.A(n_184375787), .B(n_184575789), .C(n_160175545
		), .Z(n_184675790));
	notech_ao4 i_149949205(.A(n_57873), .B(\nbus_11358[22] ), .C(n_60003), .D
		(n_58145), .Z(n_184775791));
	notech_ao4 i_133949360(.A(n_225565784), .B(n_151931934), .C(n_221065739)
		, .D(n_58084), .Z(n_185075794));
	notech_ao4 i_133849361(.A(n_29769), .B(n_26929), .C(n_58429), .D(n_28009
		), .Z(n_185275796));
	notech_nand3 i_134149358(.A(n_185075794), .B(n_185275796), .C(n_159375537
		), .Z(n_185375797));
	notech_ao4 i_133649363(.A(n_57875), .B(\nbus_11358[24] ), .C(n_60001), .D
		(n_58147), .Z(n_185475798));
	notech_ao4 i_133249367(.A(n_151931934), .B(n_225665785), .C(n_58084), .D
		(n_222565754), .Z(n_185775801));
	notech_ao4 i_133149368(.A(n_26929), .B(n_29765), .C(n_58429), .D(n_28008
		), .Z(n_185975803));
	notech_nand3 i_133449365(.A(n_185775801), .B(n_185975803), .C(n_158575529
		), .Z(n_186075804));
	notech_ao4 i_132949370(.A(n_57875), .B(n_56347), .C(n_58147), .D(n_60002
		), .Z(n_186175805));
	notech_ao4 i_123349466(.A(n_225665785), .B(n_3843), .C(n_222565754), .D(n_3858
		), .Z(n_186475808));
	notech_ao4 i_123249467(.A(n_29765), .B(n_26642), .C(n_3857), .D(n_28008)
		, .Z(n_186675810));
	notech_nand3 i_123549464(.A(n_186475808), .B(n_186675810), .C(n_157775521
		), .Z(n_186775811));
	notech_ao4 i_123049469(.A(n_3877), .B(n_56347), .C(n_60002), .D(n_148228759
		), .Z(n_186875812));
	notech_ao4 i_122649473(.A(n_225765786), .B(n_3843), .C(n_224065769), .D(n_3858
		), .Z(n_187175815));
	notech_ao4 i_122549474(.A(n_29708), .B(n_26642), .C(n_3857), .D(n_28007)
		, .Z(n_187375817));
	notech_ao4 i_122249477(.A(n_3877), .B(\nbus_11358[22] ), .C(n_60003), .D
		(n_148228759), .Z(n_187575819));
	notech_and4 i_122449475(.A(n_54667), .B(n_187575819), .C(n_26617), .D(n_156475508
		), .Z(n_188075822));
	notech_ao4 i_9047609(.A(n_316491659), .B(n_319891625), .C(n_30821), .D(n_60223
		), .Z(n_188175823));
	notech_ao4 i_9147608(.A(n_30822), .B(n_60223), .C(n_23507), .D(n_54974),
		 .Z(n_188275824));
	notech_and3 i_9247607(.A(n_316691657), .B(n_316291661), .C(n_30803), .Z(n_188375825
		));
	notech_and2 i_9347606(.A(n_309591728), .B(n_26696), .Z(n_188575826));
	notech_or4 i_88146847(.A(n_56837), .B(n_313747721), .C(n_2938), .D(n_2937
		), .Z(n_188675827));
	notech_or4 i_116146576(.A(n_54727), .B(n_57087), .C(instrc[116]), .D(n_57229
		), .Z(n_188775828));
	notech_or4 i_10247597(.A(n_56832), .B(n_56944), .C(n_56579), .D(n_28001)
		, .Z(n_189275833));
	notech_or4 i_9947600(.A(nbus_11295[16]), .B(n_60945), .C(n_54974), .D(n_26942
		), .Z(n_189575836));
	notech_or2 i_9647603(.A(n_60009), .B(n_188375825), .Z(n_189875839));
	notech_or4 i_12547575(.A(n_317591648), .B(n_60841), .C(n_54974), .D(\nbus_11358[18] 
		), .Z(n_190375844));
	notech_nand2 i_12247578(.A(n_151328790), .B(\regs_13_14[18] ), .Z(n_190875847
		));
	notech_or4 i_11947581(.A(n_60945), .B(nbus_11295[18]), .C(n_54974), .D(n_26942
		), .Z(n_191175850));
	notech_or2 i_22147479(.A(n_149428771), .B(\nbus_11358[16] ), .Z(n_191575854
		));
	notech_or4 i_21847482(.A(n_56824), .B(n_56946), .C(n_56527), .D(n_28001)
		, .Z(n_191875857));
	notech_or4 i_21547485(.A(n_26062), .B(n_311891705), .C(n_254466073), .D(n_27712
		), .Z(n_192175860));
	notech_or4 i_27047430(.A(n_3854), .B(n_3845), .C(n_58020), .D(\nbus_11358[16] 
		), .Z(n_192275861));
	notech_or2 i_26947431(.A(n_60009), .B(n_148228759), .Z(n_192575864));
	notech_or4 i_26447436(.A(n_62864), .B(n_3845), .C(n_62808), .D(\nbus_11365[16] 
		), .Z(n_193075869));
	notech_or4 i_81046914(.A(n_56824), .B(n_56946), .C(n_56649), .D(n_28003)
		, .Z(n_193175870));
	notech_or4 i_80946915(.A(n_54756), .B(n_58494), .C(n_56432), .D(n_56302)
		, .Z(n_193475873));
	notech_or2 i_80446920(.A(n_3861), .B(n_306824332), .Z(n_193975878));
	notech_nand2 i_7547624(.A(n_60223), .B(read_data[16]), .Z(n_194075879)
		);
	notech_nor2 i_88646842(.A(n_60009), .B(n_58319), .Z(n_194175880));
	notech_ao4 i_186845898(.A(n_29710), .B(n_201175950), .C(n_307624340), .D
		(n_60223), .Z(n_194475883));
	notech_ao3 i_76847688(.A(n_194075879), .B(n_194475883), .C(n_194175880),
		 .Z(n_194675885));
	notech_ao4 i_180345960(.A(n_77522039), .B(n_306624330), .C(n_241472894),
		 .D(\nbus_11365[18] ), .Z(n_194775886));
	notech_ao4 i_180245961(.A(n_29711), .B(n_307324337), .C(n_95222216), .D(n_307124335
		), .Z(n_194975888));
	notech_ao4 i_179945964(.A(n_3864), .B(n_58141), .C(n_58494), .D(n_60121865
		), .Z(n_195175890));
	notech_and4 i_180145962(.A(n_193175870), .B(n_195175890), .C(n_26621), .D
		(n_193475873), .Z(n_195475893));
	notech_ao4 i_134046404(.A(n_56601), .B(n_311224366), .C(n_263180132), .D
		(\nbus_11365[16] ), .Z(n_195575894));
	notech_ao4 i_133946405(.A(n_254466073), .B(n_57595), .C(n_252966058), .D
		(n_3858), .Z(n_195775896));
	notech_ao4 i_133646408(.A(n_29710), .B(n_26642), .C(n_313747721), .D(n_147671956
		), .Z(n_195975898));
	notech_and4 i_133846406(.A(n_194675885), .B(n_195975898), .C(n_192275861
		), .D(n_192575864), .Z(n_196275901));
	notech_ao4 i_129346448(.A(n_310891715), .B(n_252966058), .C(n_311991704)
		, .D(n_312324377), .Z(n_196375902));
	notech_ao4 i_129146450(.A(n_57173), .B(\nbus_11365[16] ), .C(n_313747721
		), .D(n_148728764), .Z(n_196575904));
	notech_and4 i_129546446(.A(n_191875857), .B(n_196575904), .C(n_192175860
		), .D(n_196375902), .Z(n_196775906));
	notech_ao4 i_128846453(.A(n_60009), .B(n_149128768), .C(n_149228769), .D
		(n_29710), .Z(n_196875907));
	notech_ao4 i_128646455(.A(n_60356), .B(n_28105), .C(n_54638), .D(n_28970
		), .Z(n_197075909));
	notech_and4 i_129046451(.A(n_54667), .B(n_197075909), .C(n_196875907), .D
		(n_191575854), .Z(n_197275911));
	notech_ao4 i_120946531(.A(n_60121865), .B(n_54974), .C(n_306024324), .D(n_57698
		), .Z(n_197375912));
	notech_ao4 i_120646533(.A(n_3861), .B(n_151128788), .C(n_77522039), .D(n_311391710
		), .Z(n_197575914));
	notech_and4 i_121146529(.A(n_197575914), .B(n_197375912), .C(n_190875847
		), .D(n_191175850), .Z(n_197775916));
	notech_ao4 i_120346536(.A(n_311291711), .B(n_28003), .C(n_151428791), .D
		(n_3864), .Z(n_197875917));
	notech_ao4 i_120146538(.A(n_54638), .B(n_28955), .C(n_59124), .D(nbus_11295
		[18]), .Z(n_198075919));
	notech_and4 i_120546534(.A(n_198075919), .B(n_190375844), .C(n_197875917
		), .D(n_26621), .Z(n_198275921));
	notech_ao4 i_118846551(.A(\nbus_11358[16] ), .B(n_188275824), .C(\nbus_11365[16] 
		), .D(n_188175823), .Z(n_198375922));
	notech_ao4 i_118646553(.A(n_312324377), .B(n_54974), .C(n_29710), .D(n_188575826
		), .Z(n_198575924));
	notech_and4 i_119046549(.A(n_189575836), .B(n_198575924), .C(n_198375922
		), .D(n_189875839), .Z(n_198775926));
	notech_ao4 i_118146556(.A(n_313747721), .B(n_151128788), .C(n_254466073)
		, .D(n_311391710), .Z(n_198875927));
	notech_ao4 i_117946558(.A(n_54638), .B(n_28953), .C(n_59124), .D(nbus_11295
		[16]), .Z(n_199075929));
	notech_and4 i_118546554(.A(n_199075929), .B(n_189275833), .C(n_198875927
		), .D(n_194075879), .Z(n_199275931));
	notech_nand3 i_131158522(.A(n_58102), .B(n_27177), .C(n_32323), .Z(n_199375932
		));
	notech_ao4 i_111058530(.A(n_30825), .B(n_60223), .C(n_23514), .D(n_319891625
		), .Z(n_199575934));
	notech_and2 i_16844328(.A(n_58530), .B(n_215476093), .Z(n_199675935));
	notech_ao4 i_132744566(.A(n_30825), .B(n_60223), .C(n_23514), .D(n_317691647
		), .Z(n_199775936));
	notech_ao4 i_146158519(.A(n_26610), .B(n_30818), .C(n_23514), .D(n_23507
		), .Z(n_199875937));
	notech_ao4 i_132844557(.A(n_30825), .B(n_60229), .C(n_314991674), .D(n_24994
		), .Z(n_199975938));
	notech_ao4 i_146344559(.A(n_59445), .B(n_26880), .C(n_39370), .D(n_26938
		), .Z(n_200075939));
	notech_and2 i_15744339(.A(n_92619108), .B(n_200575944), .Z(n_200375942)
		);
	notech_ao4 i_15844338(.A(n_26060), .B(\nbus_11358[6] ), .C(n_183858934),
		 .D(\nbus_11307[6] ), .Z(n_200475943));
	notech_nao3 i_35844138(.A(n_58024), .B(\opa_12[6] ), .C(n_3854), .Z(n_200575944
		));
	notech_or4 i_105343494(.A(n_2938), .B(n_2937), .C(n_56824), .D(n_314391680
		), .Z(n_200875947));
	notech_and2 i_145544526(.A(n_58391), .B(n_201275951), .Z(n_201175950));
	notech_nao3 i_124443318(.A(n_26627), .B(n_60356), .C(n_308891735), .Z(n_201275951
		));
	notech_or2 i_124743315(.A(n_54814), .B(n_201475953), .Z(n_201375952));
	notech_and2 i_10744388(.A(n_58505), .B(n_58481), .Z(n_201475953));
	notech_or4 i_125443308(.A(n_26062), .B(n_29652), .C(n_29658), .D(n_58177
		), .Z(n_201575954));
	notech_or2 i_17844318(.A(n_59124), .B(nbus_11295[3]), .Z(n_202875967));
	notech_or2 i_19144305(.A(n_59124), .B(nbus_11295[5]), .Z(n_204175980));
	notech_or2 i_20744289(.A(n_58411), .B(n_27989), .Z(n_205075989));
	notech_nand2 i_20444292(.A(opa[6]), .B(n_215276091), .Z(n_205375992));
	notech_or2 i_28544211(.A(n_58410), .B(n_27985), .Z(n_206576004));
	notech_or2 i_29744199(.A(n_58410), .B(n_27987), .Z(n_207776016));
	notech_nao3 i_31344183(.A(tsc[38]), .B(n_55820), .C(n_59469), .Z(n_208276021
		));
	notech_nand2 i_31244184(.A(n_200075939), .B(opa[6]), .Z(n_208576024));
	notech_or2 i_30944187(.A(n_57882), .B(\nbus_11358[6] ), .Z(n_208876027)
		);
	notech_or4 i_33644160(.A(n_3854), .B(n_139071870), .C(n_32335), .D(\nbus_11307[3] 
		), .Z(n_209776036));
	notech_or2 i_33344163(.A(n_308721251), .B(n_147671956), .Z(n_210076039)
		);
	notech_or4 i_33044166(.A(n_26767), .B(n_58163), .C(nbus_11295[3]), .D(n_60947
		), .Z(n_210376042));
	notech_or4 i_34744149(.A(n_3854), .B(n_139071870), .C(n_32335), .D(\nbus_11307[5] 
		), .Z(n_210876047));
	notech_or2 i_34444152(.A(n_308621250), .B(n_147671956), .Z(n_211176050)
		);
	notech_or4 i_34144155(.A(n_26767), .B(n_58163), .C(nbus_11295[5]), .D(n_60947
		), .Z(n_211476053));
	notech_nao3 i_35744139(.A(n_58078), .B(opd[6]), .C(n_56601), .Z(n_211776056
		));
	notech_or4 i_35244144(.A(n_62864), .B(n_146971949), .C(n_60947), .D(n_29723
		), .Z(n_212276061));
	notech_or2 i_75543770(.A(n_314791676), .B(n_58145), .Z(n_212376062));
	notech_and2 i_99243553(.A(\regs_13_14[31] ), .B(n_287027252), .Z(n_213076069
		));
	notech_nand3 i_98743558(.A(n_57115), .B(n_62808), .C(opc_10[31]), .Z(n_213776076
		));
	notech_nand2 i_9244402(.A(read_data[3]), .B(n_60223), .Z(n_213876077));
	notech_ao3 i_100643539(.A(n_60356), .B(\opa_12[3] ), .C(n_30825), .Z(n_214276081
		));
	notech_nand2 i_9544399(.A(read_data[5]), .B(n_60223), .Z(n_214376082));
	notech_ao3 i_102243524(.A(n_60356), .B(\opa_12[5] ), .C(n_30825), .Z(n_214776086
		));
	notech_ao4 i_36463(.A(n_59445), .B(n_27179), .C(n_58102), .D(n_26941), .Z
		(n_215276091));
	notech_and2 i_150344506(.A(n_199375932), .B(n_316691657), .Z(n_215476093
		));
	notech_ao4 i_6344431(.A(n_56688), .B(n_28016), .C(n_56813), .D(n_314391680
		), .Z(n_215576094));
	notech_ao4 i_201542575(.A(n_314791676), .B(n_58319), .C(n_314691677), .D
		(n_60223), .Z(n_215676095));
	notech_ao4 i_201442576(.A(n_28123), .B(n_60356), .C(n_201175950), .D(n_29619
		), .Z(n_215776096));
	notech_nand2 i_75944481(.A(n_215776096), .B(n_215676095), .Z(n_215876097
		));
	notech_ao4 i_199142598(.A(\nbus_11307[5] ), .B(n_147071950), .C(\nbus_11358[5] 
		), .D(n_58530), .Z(n_215976098));
	notech_ao4 i_199042599(.A(n_60020), .B(n_58432), .C(n_60356), .D(n_28094
		), .Z(n_216176100));
	notech_ao3 i_77444478(.A(n_215976098), .B(n_216176100), .C(n_214776086),
		 .Z(n_216276101));
	notech_ao4 i_197842611(.A(n_147071950), .B(\nbus_11307[3] ), .C(n_58530)
		, .D(\nbus_11358[3] ), .Z(n_216376102));
	notech_ao4 i_197742612(.A(n_60022), .B(n_58432), .C(n_60356), .D(n_28092
		), .Z(n_216576104));
	notech_ao3 i_77244479(.A(n_216376102), .B(n_216576104), .C(n_214276081),
		 .Z(n_216676105));
	notech_ao4 i_196442625(.A(n_96519147), .B(n_286927251), .C(n_56662), .D(n_306221226
		), .Z(n_216776106));
	notech_ao4 i_196342626(.A(n_57861), .B(\nbus_11365[31] ), .C(n_314391680
		), .D(n_143571915), .Z(n_216976108));
	notech_nand3 i_196642623(.A(n_216776106), .B(n_216976108), .C(n_213776076
		), .Z(n_217076109));
	notech_ao4 i_196142628(.A(n_57863), .B(\nbus_11358[31] ), .C(n_314791676
		), .D(n_58139), .Z(n_217176110));
	notech_ao4 i_178542803(.A(n_96519147), .B(n_58082), .C(n_303721201), .D(n_56498
		), .Z(n_217476113));
	notech_ao4 i_178442804(.A(n_57869), .B(\nbus_11365[31] ), .C(n_83019012)
		, .D(n_57596), .Z(n_217576114));
	notech_ao4 i_178242806(.A(n_29619), .B(n_26918), .C(n_57873), .D(\nbus_11358[31] 
		), .Z(n_217776116));
	notech_ao3 i_178342805(.A(n_217776116), .B(n_212376062), .C(n_215876097)
		, .Z(n_217976118));
	notech_ao4 i_144043131(.A(n_58163), .B(n_200475943), .C(n_3853), .D(n_200375942
		), .Z(n_218076119));
	notech_ao4 i_143943132(.A(n_26802), .B(n_147771957), .C(n_92019102), .D(n_57922
		), .Z(n_218276121));
	notech_ao4 i_143643135(.A(n_3874), .B(n_154175485), .C(n_3868), .D(n_147671956
		), .Z(n_218476123));
	notech_and4 i_143843133(.A(n_54667), .B(n_218476123), .C(n_311173591), .D
		(n_211776056), .Z(n_218776126));
	notech_ao4 i_143243139(.A(n_281966348), .B(n_58163), .C(n_281866347), .D
		(n_147871958), .Z(n_218876127));
	notech_ao4 i_142743141(.A(n_282266351), .B(n_3853), .C(n_282166350), .D(n_57922
		), .Z(n_219076129));
	notech_and4 i_143443137(.A(n_219076129), .B(n_218876127), .C(n_211176050
		), .D(n_211476053), .Z(n_219276131));
	notech_ao4 i_142343144(.A(n_57980), .B(\nbus_11358[5] ), .C(n_147571955)
		, .D(n_27987), .Z(n_219376132));
	notech_ao4 i_142143146(.A(n_60020), .B(n_154175485), .C(n_137675320), .D
		(n_29651), .Z(n_219576134));
	notech_and4 i_142543142(.A(n_216276101), .B(n_219576134), .C(n_219376132
		), .D(n_210876047), .Z(n_219776136));
	notech_ao4 i_141843149(.A(n_306670077), .B(n_147871958), .C(n_306570076)
		, .D(n_58163), .Z(n_219876137));
	notech_ao4 i_141643151(.A(n_306970080), .B(n_3853), .C(n_306870079), .D(n_57922
		), .Z(n_220076139));
	notech_and4 i_142043147(.A(n_220076139), .B(n_219876137), .C(n_210076039
		), .D(n_210376042), .Z(n_220276141));
	notech_ao4 i_141343154(.A(n_57980), .B(\nbus_11358[3] ), .C(n_147571955)
		, .D(n_27985), .Z(n_220376142));
	notech_ao4 i_141143156(.A(n_60022), .B(n_154175485), .C(n_29728), .D(n_137675320
		), .Z(n_220576144));
	notech_and4 i_141543152(.A(n_216676105), .B(n_220576144), .C(n_220376142
		), .D(n_209776036), .Z(n_220776146));
	notech_ao4 i_140043167(.A(n_26802), .B(n_306170072), .C(n_92019102), .D(n_306270073
		), .Z(n_220876147));
	notech_ao4 i_139943168(.A(n_92619108), .B(n_24994), .C(n_92519107), .D(n_306070071
		), .Z(n_220976148));
	notech_ao4 i_139743170(.A(n_58410), .B(n_27989), .C(n_3868), .D(n_311791706
		), .Z(n_221176150));
	notech_and4 i_140243165(.A(n_221176150), .B(n_220976148), .C(n_220876147
		), .D(n_208876027), .Z(n_221376152));
	notech_ao4 i_139443173(.A(n_3874), .B(n_57619), .C(n_199975938), .D(n_29723
		), .Z(n_221476153));
	notech_ao4 i_6744427(.A(n_28095), .B(n_60356), .C(n_58514), .D(\nbus_11307[6] 
		), .Z(n_221676155));
	notech_and3 i_139343174(.A(n_221676155), .B(n_54667), .C(n_208276021), .Z
		(n_221876157));
	notech_ao4 i_138943178(.A(n_282166350), .B(n_306270073), .C(n_281866347)
		, .D(n_305970070), .Z(n_222076159));
	notech_ao4 i_138843179(.A(n_281966348), .B(n_26697), .C(n_282066349), .D
		(n_306170072), .Z(n_222176160));
	notech_ao4 i_138643181(.A(n_308621250), .B(n_311791706), .C(n_282266351)
		, .D(n_24994), .Z(n_222376162));
	notech_and4 i_139143176(.A(n_222376162), .B(n_222176160), .C(n_222076159
		), .D(n_207776016), .Z(n_222576164));
	notech_ao4 i_138343184(.A(n_60020), .B(n_57619), .C(n_57882), .D(\nbus_11358[5] 
		), .Z(n_222676165));
	notech_ao4 i_138243185(.A(\nbus_11307[5] ), .B(n_57891), .C(n_57938), .D
		(n_29651), .Z(n_222776166));
	notech_ao4 i_138043187(.A(n_28094), .B(n_60356), .C(n_54638), .D(n_28966
		), .Z(n_222976168));
	notech_and4 i_138543182(.A(n_54667), .B(n_222976168), .C(n_222776166), .D
		(n_222676165), .Z(n_223176170));
	notech_ao4 i_137743190(.A(n_306270073), .B(n_306870079), .C(n_306670077)
		, .D(n_305970070), .Z(n_223276171));
	notech_ao4 i_137643191(.A(n_306570076), .B(n_26697), .C(n_306770078), .D
		(n_306170072), .Z(n_223376172));
	notech_ao4 i_137443193(.A(n_308721251), .B(n_311791706), .C(n_306970080)
		, .D(n_24994), .Z(n_223576174));
	notech_and4 i_137943188(.A(n_223576174), .B(n_223376172), .C(n_223276171
		), .D(n_206576004), .Z(n_223776176));
	notech_ao4 i_137143196(.A(n_60022), .B(n_57619), .C(n_57882), .D(\nbus_11358[3] 
		), .Z(n_223876177));
	notech_ao4 i_137043197(.A(n_57891), .B(\nbus_11307[3] ), .C(n_57938), .D
		(n_29728), .Z(n_223976178));
	notech_ao4 i_136843199(.A(n_28092), .B(n_60356), .C(n_54638), .D(n_28965
		), .Z(n_224176180));
	notech_and4 i_137343194(.A(n_54667), .B(n_224176180), .C(n_223976178), .D
		(n_223876177), .Z(n_224376182));
	notech_ao4 i_130343260(.A(n_142871908), .B(n_92519107), .C(\nbus_11358[6] 
		), .D(n_199675935), .Z(n_224476183));
	notech_ao4 i_130143261(.A(n_92619108), .B(n_23514), .C(n_92019102), .D(n_137575319
		), .Z(n_224576184));
	notech_ao4 i_129943263(.A(n_315691667), .B(n_3868), .C(n_26802), .D(n_137475318
		), .Z(n_224776186));
	notech_and4 i_130543258(.A(n_224776186), .B(n_224576184), .C(n_224476183
		), .D(n_205375992), .Z(n_224976188));
	notech_ao4 i_129643266(.A(n_3874), .B(n_199875937), .C(n_199775936), .D(n_29723
		), .Z(n_225076189));
	notech_ao4 i_129443268(.A(n_54638), .B(n_28949), .C(n_59124), .D(nbus_11295
		[6]), .Z(n_225276191));
	notech_and4 i_129843264(.A(n_225276191), .B(n_221676155), .C(n_225076189
		), .D(n_205075989), .Z(n_225476193));
	notech_ao4 i_129143271(.A(n_281966348), .B(n_56516), .C(n_281866347), .D
		(n_137375317), .Z(n_225576194));
	notech_ao4 i_129043272(.A(n_282166350), .B(n_137575319), .C(n_282066349)
		, .D(n_137475318), .Z(n_225676195));
	notech_ao4 i_128843274(.A(n_308621250), .B(n_315691667), .C(n_282266351)
		, .D(n_23514), .Z(n_225876197));
	notech_and4 i_129343269(.A(n_225876197), .B(n_225676195), .C(n_225576194
		), .D(n_204175980), .Z(n_226076199));
	notech_ao4 i_128543277(.A(n_57893), .B(\nbus_11358[5] ), .C(n_58411), .D
		(n_27987), .Z(n_226176200));
	notech_ao4 i_128443278(.A(n_199575934), .B(n_29651), .C(n_57892), .D(\nbus_11307[5] 
		), .Z(n_226276201));
	notech_ao4 i_128243280(.A(n_54638), .B(n_28948), .C(n_60020), .D(n_199875937
		), .Z(n_226476203));
	notech_and4 i_128743275(.A(n_226476203), .B(n_226276201), .C(n_226176200
		), .D(n_214376082), .Z(n_226676205));
	notech_ao4 i_127943283(.A(n_306670077), .B(n_137375317), .C(n_306570076)
		, .D(n_56516), .Z(n_226776206));
	notech_ao4 i_127843284(.A(n_306870079), .B(n_137575319), .C(n_306770078)
		, .D(n_137475318), .Z(n_226876207));
	notech_ao4 i_127643286(.A(n_308721251), .B(n_315691667), .C(n_306970080)
		, .D(n_23514), .Z(n_227076209));
	notech_and4 i_128143281(.A(n_227076209), .B(n_226876207), .C(n_226776206
		), .D(n_202875967), .Z(n_227276211));
	notech_ao4 i_127343289(.A(n_57893), .B(\nbus_11358[3] ), .C(n_58411), .D
		(n_27985), .Z(n_227376212));
	notech_ao4 i_127243290(.A(n_199575934), .B(n_29728), .C(n_57892), .D(\nbus_11307[3] 
		), .Z(n_227476213));
	notech_ao4 i_127043292(.A(n_54638), .B(n_28946), .C(n_60022), .D(n_199875937
		), .Z(n_227676215));
	notech_and4 i_127543287(.A(n_227676215), .B(n_227476213), .C(n_227376212
		), .D(n_213876077), .Z(n_227876217));
	notech_or4 i_28035102(.A(n_2888), .B(n_2877), .C(n_1864), .D(n_60234), .Z
		(n_227976218));
	notech_and3 i_15334958(.A(n_22322), .B(n_1884), .C(n_236276301), .Z(n_228176220
		));
	notech_ao4 i_15234959(.A(n_2653), .B(n_60234), .C(n_23045), .D(nbus_11310
		[1]), .Z(n_228276221));
	notech_ao4 i_14634965(.A(n_23045), .B(nbus_11310[8]), .C(n_230076239), .D
		(n_60234), .Z(n_228476223));
	notech_ao4 i_14534966(.A(n_23045), .B(nbus_11310[9]), .C(n_230076239), .D
		(n_60234), .Z(n_228676225));
	notech_ao4 i_14434967(.A(n_23045), .B(nbus_11310[10]), .C(n_230076239), 
		.D(n_60234), .Z(n_228876227));
	notech_ao4 i_14334968(.A(n_23045), .B(nbus_11310[11]), .C(n_230076239), 
		.D(n_60234), .Z(n_229076229));
	notech_ao4 i_14234969(.A(n_23045), .B(nbus_11310[12]), .C(n_230076239), 
		.D(n_60234), .Z(n_229276231));
	notech_ao4 i_14134970(.A(n_23045), .B(nbus_11310[13]), .C(n_230076239), 
		.D(n_60234), .Z(n_229476233));
	notech_ao4 i_14034971(.A(n_23045), .B(nbus_11310[14]), .C(n_230076239), 
		.D(n_60234), .Z(n_229676235));
	notech_ao4 i_13934972(.A(n_23045), .B(nbus_11310[15]), .C(n_60234), .D(n_230076239
		), .Z(n_229876237));
	notech_and3 i_66634466(.A(n_25385), .B(n_2678), .C(n_2654), .Z(n_230076239
		));
	notech_and4 i_13834973(.A(n_23052), .B(n_23049), .C(n_81910939), .D(n_230276241
		), .Z(n_230176240));
	notech_or2 i_68834444(.A(n_23045), .B(nbus_11310[16]), .Z(n_230276241)
		);
	notech_and4 i_13734974(.A(n_23052), .B(n_23049), .C(n_81910939), .D(n_230476243
		), .Z(n_230376242));
	notech_or2 i_71034422(.A(n_23045), .B(nbus_11310[17]), .Z(n_230476243)
		);
	notech_and4 i_13634975(.A(n_23052), .B(n_23049), .C(n_81910939), .D(n_230676245
		), .Z(n_230576244));
	notech_or2 i_73334400(.A(n_23045), .B(nbus_11310[18]), .Z(n_230676245)
		);
	notech_and4 i_13534976(.A(n_23052), .B(n_23049), .C(n_81910939), .D(n_230876247
		), .Z(n_230776246));
	notech_or2 i_75534378(.A(n_23045), .B(nbus_11310[19]), .Z(n_230876247)
		);
	notech_and4 i_13434977(.A(n_23052), .B(n_23049), .C(n_81910939), .D(n_231076249
		), .Z(n_230976248));
	notech_or2 i_77734356(.A(n_23045), .B(nbus_11310[20]), .Z(n_231076249)
		);
	notech_and4 i_13334978(.A(n_23052), .B(n_23049), .C(n_81910939), .D(n_231276251
		), .Z(n_231176250));
	notech_or2 i_80034334(.A(n_23045), .B(nbus_11310[21]), .Z(n_231276251)
		);
	notech_and4 i_13134979(.A(n_23052), .B(n_23049), .C(n_81910939), .D(n_231476253
		), .Z(n_231376252));
	notech_or2 i_82234312(.A(n_23045), .B(nbus_11310[22]), .Z(n_231476253)
		);
	notech_and4 i_13034980(.A(n_23052), .B(n_23049), .C(n_81910939), .D(n_231676255
		), .Z(n_231576254));
	notech_or2 i_84434290(.A(n_57143), .B(nbus_11310[23]), .Z(n_231676255)
		);
	notech_and4 i_12934981(.A(n_23052), .B(n_23049), .C(n_81910939), .D(n_231876257
		), .Z(n_231776256));
	notech_or2 i_86634268(.A(n_57143), .B(nbus_11310[24]), .Z(n_231876257)
		);
	notech_and4 i_12834982(.A(n_23052), .B(n_23049), .C(n_81910939), .D(n_232076259
		), .Z(n_231976258));
	notech_or2 i_88834246(.A(n_57143), .B(nbus_11310[25]), .Z(n_232076259)
		);
	notech_and4 i_12734983(.A(n_23052), .B(n_23049), .C(n_81910939), .D(n_232276261
		), .Z(n_232176260));
	notech_or2 i_91034224(.A(n_57143), .B(nbus_11310[26]), .Z(n_232276261)
		);
	notech_and4 i_12634984(.A(n_23052), .B(n_23049), .C(n_81910939), .D(n_232476263
		), .Z(n_232376262));
	notech_or2 i_93234202(.A(n_57143), .B(nbus_11310[27]), .Z(n_232476263)
		);
	notech_and4 i_12534985(.A(n_23052), .B(n_57155), .C(n_81910939), .D(n_232676265
		), .Z(n_232576264));
	notech_or2 i_95434180(.A(n_57143), .B(nbus_11310[28]), .Z(n_232676265)
		);
	notech_and4 i_12434986(.A(n_23052), .B(n_57155), .C(n_81910939), .D(n_232876267
		), .Z(n_232776266));
	notech_or2 i_97634158(.A(n_57143), .B(nbus_11310[29]), .Z(n_232876267)
		);
	notech_and4 i_12334987(.A(n_23052), .B(n_57155), .C(n_81910939), .D(n_233076269
		), .Z(n_232976268));
	notech_or2 i_99934136(.A(n_57143), .B(nbus_11310[30]), .Z(n_233076269)
		);
	notech_and4 i_12234988(.A(n_23052), .B(n_57155), .C(n_81910939), .D(n_233276271
		), .Z(n_233176270));
	notech_or2 i_102134114(.A(n_57143), .B(nbus_11310[31]), .Z(n_233276271)
		);
	notech_nand3 i_21834893(.A(n_27784), .B(n_2944), .C(nbus_158[0]), .Z(n_233676275
		));
	notech_nao3 i_21134900(.A(n_295591839), .B(nbus_163[0]), .C(n_27907), .Z
		(n_234376282));
	notech_nao3 i_20434907(.A(n_2947), .B(n_10901), .C(n_19093), .Z(n_235076289
		));
	notech_nand2 i_19734914(.A(readio_data[0]), .B(n_26711), .Z(n_235776296)
		);
	notech_or2 i_21934892(.A(n_57143), .B(nbus_11310[0]), .Z(n_236276301));
	notech_nand3 i_25234863(.A(nbus_158[1]), .B(n_27784), .C(n_2944), .Z(n_236576304
		));
	notech_nao3 i_24434870(.A(nbus_163[1]), .B(n_295591839), .C(n_27907), .Z
		(n_237276311));
	notech_nao3 i_23734877(.A(n_2947), .B(n_10902), .C(n_19093), .Z(n_237976318
		));
	notech_nao3 i_43934692(.A(nbus_14521[8]), .B(n_32316), .C(n_2949), .Z(n_240876347
		));
	notech_nao3 i_46934662(.A(nbus_14521[9]), .B(n_32316), .C(n_2949), .Z(n_243776376
		));
	notech_nao3 i_49934632(.A(nbus_14521[10]), .B(n_32316), .C(n_2949), .Z(n_246676405
		));
	notech_nao3 i_52934602(.A(nbus_14521[11]), .B(n_32316), .C(n_2949), .Z(n_249576434
		));
	notech_nao3 i_55934572(.A(nbus_14521[12]), .B(n_32316), .C(n_2949), .Z(n_252476463
		));
	notech_nao3 i_59034542(.A(n_32316), .B(nbus_14521[13]), .C(n_2949), .Z(n_255376492
		));
	notech_nao3 i_62034512(.A(nbus_14521[14]), .B(n_32316), .C(n_2949), .Z(n_258276521
		));
	notech_nao3 i_65034482(.A(resa_arithbox[15]), .B(n_60356), .C(n_2941), .Z
		(n_261176550));
	notech_nao3 i_68734445(.A(resa_shift4box[16]), .B(n_27877), .C(n_293591841
		), .Z(n_262476563));
	notech_or2 i_68634446(.A(n_57537), .B(nbus_11295[16]), .Z(n_262776566)
		);
	notech_nao3 i_68334449(.A(cr2_reg[16]), .B(n_32341), .C(n_2949), .Z(n_263076569
		));
	notech_nao3 i_68034452(.A(resa_arithbox[16]), .B(n_60356), .C(n_2941), .Z
		(n_263376572));
	notech_or2 i_67534457(.A(n_1876), .B(n_29710), .Z(n_263876577));
	notech_nao3 i_67234460(.A(n_60356), .B(opc[0]), .C(n_25385), .Z(n_264176580
		));
	notech_nand2 i_66934463(.A(nbus_164[16]), .B(n_296076899), .Z(n_264476583
		));
	notech_nao3 i_70934423(.A(resa_shift4box[17]), .B(n_27877), .C(n_293591841
		), .Z(n_264576584));
	notech_or2 i_70834424(.A(n_57537), .B(nbus_11295[17]), .Z(n_264876587)
		);
	notech_nao3 i_70534427(.A(cr2_reg[17]), .B(n_32341), .C(n_2949), .Z(n_265176590
		));
	notech_nao3 i_70234430(.A(resa_arithbox[17]), .B(n_60356), .C(n_2941), .Z
		(n_265476593));
	notech_or2 i_69734435(.A(n_1876), .B(n_29772), .Z(n_265976598));
	notech_nao3 i_69434438(.A(n_60356), .B(opc[1]), .C(n_25385), .Z(n_266276601
		));
	notech_nand2 i_69134441(.A(nbus_164[17]), .B(n_296076899), .Z(n_266576604
		));
	notech_nao3 i_73234401(.A(resa_shift4box[18]), .B(n_27877), .C(n_293591841
		), .Z(n_266676605));
	notech_or2 i_73134402(.A(n_57538), .B(nbus_11295[18]), .Z(n_266976608)
		);
	notech_nao3 i_72834405(.A(cr2_reg[18]), .B(n_32341), .C(n_2949), .Z(n_267276611
		));
	notech_nao3 i_72534408(.A(resa_arithbox[18]), .B(n_60356), .C(n_2941), .Z
		(n_267576614));
	notech_or2 i_72034413(.A(n_1876), .B(n_29711), .Z(n_268076619));
	notech_nao3 i_71734416(.A(n_60356), .B(opc[2]), .C(n_25385), .Z(n_268376622
		));
	notech_nand2 i_71334419(.A(nbus_164[18]), .B(n_296076899), .Z(n_268676625
		));
	notech_nao3 i_75434379(.A(resa_shift4box[19]), .B(n_27877), .C(n_293591841
		), .Z(n_268776626));
	notech_or2 i_75334380(.A(n_57538), .B(nbus_11295[19]), .Z(n_269076629)
		);
	notech_nao3 i_75034383(.A(cr2_reg[19]), .B(n_32341), .C(n_2949), .Z(n_269376632
		));
	notech_nao3 i_74734386(.A(resa_arithbox[19]), .B(n_60358), .C(n_2941), .Z
		(n_269676635));
	notech_or2 i_74234391(.A(n_1876), .B(n_29773), .Z(n_270176640));
	notech_nao3 i_73934394(.A(n_60349), .B(opc[3]), .C(n_25385), .Z(n_270476643
		));
	notech_nand2 i_73634397(.A(nbus_164[19]), .B(n_296076899), .Z(n_270776646
		));
	notech_nao3 i_77634357(.A(resa_shift4box[20]), .B(n_27877), .C(n_293591841
		), .Z(n_270876647));
	notech_or2 i_77534358(.A(n_57538), .B(nbus_11295[20]), .Z(n_271176650)
		);
	notech_nao3 i_77234361(.A(cr2_reg[20]), .B(n_32341), .C(n_2949), .Z(n_271476653
		));
	notech_nao3 i_76934364(.A(resa_arithbox[20]), .B(n_60349), .C(n_2941), .Z
		(n_271776656));
	notech_or2 i_76434369(.A(n_1876), .B(n_29775), .Z(n_272276661));
	notech_nao3 i_76134372(.A(n_60349), .B(opc[4]), .C(n_25385), .Z(n_272576664
		));
	notech_nand2 i_75834375(.A(nbus_164[20]), .B(n_296076899), .Z(n_272876667
		));
	notech_nao3 i_79934335(.A(resa_shift4box[21]), .B(n_27877), .C(n_293591841
		), .Z(n_272976668));
	notech_or2 i_79834336(.A(n_57537), .B(nbus_11295[21]), .Z(n_273276671)
		);
	notech_nao3 i_79434339(.A(cr2_reg[21]), .B(n_32341), .C(n_2949), .Z(n_273576674
		));
	notech_nao3 i_79134342(.A(resa_arithbox[21]), .B(n_60349), .C(n_2941), .Z
		(n_273876677));
	notech_or2 i_78634347(.A(n_1876), .B(n_29681), .Z(n_274376682));
	notech_nao3 i_78334350(.A(n_60347), .B(opc[5]), .C(n_25385), .Z(n_274676685
		));
	notech_nand2 i_78034353(.A(nbus_164[21]), .B(n_296076899), .Z(n_274976688
		));
	notech_nao3 i_82134313(.A(resa_shift4box[22]), .B(n_27877), .C(n_293591841
		), .Z(n_275076689));
	notech_or2 i_82034314(.A(n_57537), .B(nbus_11295[22]), .Z(n_275376692)
		);
	notech_nao3 i_81734317(.A(cr2_reg[22]), .B(n_32341), .C(n_2949), .Z(n_275676695
		));
	notech_nao3 i_81434320(.A(resa_arithbox[22]), .B(n_60347), .C(n_2941), .Z
		(n_275976698));
	notech_or2 i_80934325(.A(n_1876), .B(n_29708), .Z(n_276476703));
	notech_nao3 i_80634328(.A(n_60349), .B(opc[6]), .C(n_25385), .Z(n_276776706
		));
	notech_nand2 i_80334331(.A(nbus_164[22]), .B(n_296076899), .Z(n_277076709
		));
	notech_nao3 i_84334291(.A(resa_shift4box[23]), .B(n_27877), .C(n_293591841
		), .Z(n_277176710));
	notech_or2 i_84234292(.A(n_57537), .B(nbus_11295[23]), .Z(n_277476713)
		);
	notech_nao3 i_83934295(.A(cr2_reg[23]), .B(n_32341), .C(n_2949), .Z(n_277776716
		));
	notech_nao3 i_83634298(.A(resa_arithbox[23]), .B(n_60349), .C(n_2941), .Z
		(n_278076719));
	notech_or2 i_83134303(.A(n_1876), .B(n_29765), .Z(n_278576724));
	notech_nao3 i_82834306(.A(n_60349), .B(opc[7]), .C(n_25385), .Z(n_278876727
		));
	notech_nand2 i_82534309(.A(nbus_164[23]), .B(n_296076899), .Z(n_279176730
		));
	notech_nao3 i_86534269(.A(resa_shift4box[24]), .B(n_27877), .C(n_293591841
		), .Z(n_279276731));
	notech_or2 i_86434270(.A(n_57537), .B(nbus_11295[24]), .Z(n_279576734)
		);
	notech_nao3 i_86134273(.A(cr2_reg[24]), .B(n_32341), .C(n_2949), .Z(n_279876737
		));
	notech_nao3 i_85834276(.A(resa_arithbox[24]), .B(n_60349), .C(n_2941), .Z
		(n_280176740));
	notech_or2 i_85334281(.A(n_1876), .B(n_29769), .Z(n_280676745));
	notech_nao3 i_85034284(.A(n_60349), .B(opc[8]), .C(n_25385), .Z(n_280976748
		));
	notech_nand2 i_84734287(.A(nbus_164[24]), .B(n_296076899), .Z(n_281276751
		));
	notech_nao3 i_88734247(.A(resa_shift4box[25]), .B(n_27877), .C(n_293591841
		), .Z(n_281376752));
	notech_or2 i_88634248(.A(n_57537), .B(nbus_11295[25]), .Z(n_281676755)
		);
	notech_nao3 i_88334251(.A(cr2_reg[25]), .B(n_57992), .C(n_57933), .Z(n_281976758
		));
	notech_nao3 i_88034254(.A(resa_arithbox[25]), .B(n_60349), .C(n_2941), .Z
		(n_282276761));
	notech_or2 i_87534259(.A(n_1876), .B(n_29770), .Z(n_282776766));
	notech_nao3 i_87234262(.A(n_60349), .B(opc[9]), .C(n_25385), .Z(n_283076769
		));
	notech_nand2 i_86934265(.A(nbus_164[25]), .B(n_296076899), .Z(n_283376772
		));
	notech_nao3 i_90934225(.A(resa_shift4box[26]), .B(n_27877), .C(n_293591841
		), .Z(n_283476773));
	notech_or2 i_90834226(.A(n_57538), .B(nbus_11295[26]), .Z(n_283776776)
		);
	notech_nao3 i_90534229(.A(cr2_reg[26]), .B(n_57992), .C(n_57933), .Z(n_284076779
		));
	notech_nao3 i_90234232(.A(resa_arithbox[26]), .B(n_60349), .C(n_58072), 
		.Z(n_284376782));
	notech_or2 i_89734237(.A(n_1876), .B(n_29660), .Z(n_284876787));
	notech_nao3 i_89434240(.A(n_60349), .B(opc[10]), .C(n_58046), .Z(n_285176790
		));
	notech_nand2 i_89134243(.A(nbus_164[26]), .B(n_296076899), .Z(n_285476793
		));
	notech_nao3 i_93134203(.A(resa_shift4box[27]), .B(n_27877), .C(n_293591841
		), .Z(n_285576794));
	notech_or2 i_93034204(.A(n_57538), .B(nbus_11295[27]), .Z(n_285876797)
		);
	notech_nao3 i_92734207(.A(cr2_reg[27]), .B(n_57992), .C(n_57933), .Z(n_286176800
		));
	notech_nao3 i_92434210(.A(resa_arithbox[27]), .B(n_60349), .C(n_58072), 
		.Z(n_286476803));
	notech_or2 i_91934215(.A(n_1876), .B(n_29661), .Z(n_286976808));
	notech_nao3 i_91634218(.A(n_60349), .B(opc[11]), .C(n_58046), .Z(n_287276811
		));
	notech_nand2 i_91334221(.A(nbus_164[27]), .B(n_296076899), .Z(n_287576814
		));
	notech_nao3 i_95334181(.A(resa_shift4box[28]), .B(n_27877), .C(n_293591841
		), .Z(n_287676815));
	notech_or2 i_95234182(.A(n_57538), .B(nbus_11295[28]), .Z(n_287976818)
		);
	notech_nao3 i_94934185(.A(cr2_reg[28]), .B(n_57992), .C(n_57933), .Z(n_288276821
		));
	notech_nao3 i_94634188(.A(resa_arithbox[28]), .B(n_60347), .C(n_58072), 
		.Z(n_288576824));
	notech_or2 i_94134193(.A(n_1876), .B(n_29662), .Z(n_289076829));
	notech_nao3 i_93834196(.A(n_60347), .B(opc[12]), .C(n_58046), .Z(n_289376832
		));
	notech_nand2 i_93534199(.A(nbus_164[28]), .B(n_296076899), .Z(n_289676835
		));
	notech_nao3 i_97534159(.A(resa_shift4box[29]), .B(n_57899), .C(n_293591841
		), .Z(n_289776836));
	notech_or2 i_97434160(.A(n_57538), .B(nbus_11295[29]), .Z(n_290076839)
		);
	notech_nao3 i_97134163(.A(cr2_reg[29]), .B(n_57992), .C(n_57933), .Z(n_290376842
		));
	notech_nao3 i_96834166(.A(resa_arithbox[29]), .B(n_60347), .C(n_58072), 
		.Z(n_290676845));
	notech_or2 i_96334171(.A(n_1876), .B(n_29659), .Z(n_291176850));
	notech_nao3 i_96034174(.A(n_60347), .B(opc[13]), .C(n_58046), .Z(n_291476853
		));
	notech_nand2 i_95734177(.A(nbus_164[29]), .B(n_296076899), .Z(n_291776856
		));
	notech_nao3 i_99834137(.A(resa_shift4box[30]), .B(n_57899), .C(n_293591841
		), .Z(n_291876857));
	notech_or2 i_99734138(.A(n_57538), .B(nbus_11295[30]), .Z(n_292176860)
		);
	notech_nao3 i_99434141(.A(cr2_reg[30]), .B(n_57992), .C(n_57933), .Z(n_292476863
		));
	notech_nao3 i_99134144(.A(resa_arithbox[30]), .B(n_60347), .C(n_58072), 
		.Z(n_292776866));
	notech_or2 i_98634149(.A(n_1876), .B(n_29591), .Z(n_293276871));
	notech_nao3 i_98334152(.A(n_60358), .B(opc[14]), .C(n_58046), .Z(n_293576874
		));
	notech_nand2 i_97934155(.A(nbus_164[30]), .B(n_296076899), .Z(n_293876877
		));
	notech_nao3 i_102034115(.A(resa_shift4box[31]), .B(n_57899), .C(n_293591841
		), .Z(n_293976878));
	notech_nao3 i_101934116(.A(n_10932), .B(n_2947), .C(n_19093), .Z(n_294276881
		));
	notech_nao3 i_101634119(.A(nbus_14521[31]), .B(n_32316), .C(n_57933), .Z
		(n_294576884));
	notech_nand3 i_101334122(.A(nbus_157[31]), .B(n_27906), .C(n_60347), .Z(n_294876887
		));
	notech_nand2 i_100834127(.A(resa_shiftbox[31]), .B(n_26712), .Z(n_295376892
		));
	notech_nao3 i_100534130(.A(n_60347), .B(opc[15]), .C(n_58046), .Z(n_295676895
		));
	notech_nand2 i_100234133(.A(nbus_164[31]), .B(n_296076899), .Z(n_295976898
		));
	notech_nor2 i_42035098(.A(n_27917), .B(n_303747815), .Z(n_296076899));
	notech_or4 i_42735096(.A(n_25625), .B(n_28081), .C(n_59435), .D(n_60234)
		, .Z(n_296376902));
	notech_ao4 i_193433219(.A(n_296376902), .B(n_28016), .C(n_233176270), .D
		(\nbus_11365[31] ), .Z(n_296476903));
	notech_ao4 i_193233221(.A(n_227976218), .B(n_30017), .C(n_308547770), .D
		(n_28908), .Z(n_296676905));
	notech_and4 i_193633217(.A(n_296676905), .B(n_296476903), .C(n_295676895
		), .D(n_295976898), .Z(n_296876907));
	notech_ao4 i_192933224(.A(n_57538), .B(nbus_11295[31]), .C(n_23059), .D(n_27941
		), .Z(n_296976908));
	notech_ao4 i_192833225(.A(n_1877), .B(n_28832), .C(n_1876), .D(n_29619),
		 .Z(n_297176910));
	notech_and4 i_193733216(.A(n_296976908), .B(n_297176910), .C(n_296876907
		), .D(n_295376892), .Z(n_297376912));
	notech_ao4 i_192433229(.A(n_23003), .B(\nbus_11358[31] ), .C(n_27879), .D
		(n_28769), .Z(n_297476913));
	notech_ao4 i_192233231(.A(n_23019), .B(n_27847), .C(n_27781), .D(n_28737
		), .Z(n_297676915));
	notech_and4 i_192633227(.A(n_297676915), .B(n_297476913), .C(n_294576884
		), .D(n_294876887), .Z(n_297876917));
	notech_ao4 i_191933234(.A(n_23029), .B(n_28717), .C(n_23031), .D(n_27691
		), .Z(n_297976918));
	notech_and4 i_192133232(.A(n_3901), .B(n_297976918), .C(n_293976878), .D
		(n_294276881), .Z(n_298276921));
	notech_ao4 i_191433239(.A(n_296376902), .B(n_28015), .C(n_232976268), .D
		(\nbus_11365[30] ), .Z(n_298476923));
	notech_ao4 i_191233241(.A(n_57379), .B(n_30016), .C(n_308547770), .D(n_28907
		), .Z(n_298676925));
	notech_and4 i_191633237(.A(n_298676925), .B(n_298476923), .C(n_293576874
		), .D(n_293876877), .Z(n_298876927));
	notech_ao4 i_190933244(.A(n_18756873), .B(n_28877), .C(n_23059), .D(n_27940
		), .Z(n_298976928));
	notech_ao4 i_190833245(.A(n_27879), .B(n_28768), .C(n_1877), .D(n_28831)
		, .Z(n_299176930));
	notech_and4 i_191733236(.A(n_298976928), .B(n_299176930), .C(n_298876927
		), .D(n_293276871), .Z(n_299376932));
	notech_ao4 i_190433249(.A(n_23009), .B(n_28801), .C(n_23003), .D(\nbus_11358[30] 
		), .Z(n_299476933));
	notech_ao4 i_190233251(.A(n_23023), .B(n_27675), .C(n_23019), .D(n_27539
		), .Z(n_299676935));
	notech_and4 i_190633247(.A(n_299676935), .B(n_299476933), .C(n_292476863
		), .D(n_292776866), .Z(n_299876937));
	notech_ao4 i_189933254(.A(n_23940), .B(n_30015), .C(n_23029), .D(n_28716
		), .Z(n_299976938));
	notech_and4 i_190133252(.A(n_3901), .B(n_299976938), .C(n_291876857), .D
		(n_292176860), .Z(n_300276941));
	notech_ao4 i_189433259(.A(n_296376902), .B(n_28014), .C(n_232776266), .D
		(\nbus_11365[29] ), .Z(n_300476943));
	notech_ao4 i_189233261(.A(n_227976218), .B(n_30014), .C(n_308547770), .D
		(n_28906), .Z(n_300676945));
	notech_and4 i_189633257(.A(n_300676945), .B(n_300476943), .C(n_291476853
		), .D(n_291776856), .Z(n_300876947));
	notech_ao4 i_188933264(.A(n_18756873), .B(n_28876), .C(n_23059), .D(n_27939
		), .Z(n_300976948));
	notech_ao4 i_188833265(.A(n_27879), .B(n_28767), .C(n_1877), .D(n_28830)
		, .Z(n_301176950));
	notech_and4 i_189733256(.A(n_300976948), .B(n_301176950), .C(n_300876947
		), .D(n_291176850), .Z(n_301376952));
	notech_ao4 i_188433269(.A(n_23009), .B(n_28800), .C(n_23003), .D(\nbus_11358[29] 
		), .Z(n_301476953));
	notech_ao4 i_188233271(.A(n_23023), .B(n_27674), .C(n_23019), .D(n_27538
		), .Z(n_301676955));
	notech_and4 i_188633267(.A(n_301676955), .B(n_301476953), .C(n_290376842
		), .D(n_290676845), .Z(n_301876957));
	notech_ao4 i_187933274(.A(n_30013), .B(n_23940), .C(n_23029), .D(n_28715
		), .Z(n_301976958));
	notech_and4 i_188133272(.A(n_3901), .B(n_301976958), .C(n_289776836), .D
		(n_290076839), .Z(n_302276961));
	notech_ao4 i_187433279(.A(n_296376902), .B(n_28013), .C(n_232576264), .D
		(\nbus_11365[28] ), .Z(n_302476963));
	notech_ao4 i_187233281(.A(n_227976218), .B(n_30012), .C(n_308547770), .D
		(n_28905), .Z(n_302676965));
	notech_and4 i_187633277(.A(n_302676965), .B(n_302476963), .C(n_289376832
		), .D(n_289676835), .Z(n_302876967));
	notech_ao4 i_186933284(.A(n_18756873), .B(n_28875), .C(n_23059), .D(n_27938
		), .Z(n_302976968));
	notech_ao4 i_186833285(.A(n_27879), .B(n_28766), .C(n_1877), .D(n_28829)
		, .Z(n_303176970));
	notech_and4 i_187733276(.A(n_302976968), .B(n_303176970), .C(n_302876967
		), .D(n_289076829), .Z(n_303376972));
	notech_ao4 i_186433289(.A(n_23009), .B(n_28799), .C(n_23003), .D(\nbus_11358[28] 
		), .Z(n_303476973));
	notech_ao4 i_186233291(.A(n_23023), .B(n_27673), .C(n_23019), .D(n_27537
		), .Z(n_303676975));
	notech_and4 i_186633287(.A(n_303676975), .B(n_303476973), .C(n_288276821
		), .D(n_288576824), .Z(n_303876977));
	notech_ao4 i_185933294(.A(n_23940), .B(n_30011), .C(n_23029), .D(n_28714
		), .Z(n_303976978));
	notech_and4 i_186133292(.A(n_3901), .B(n_303976978), .C(n_287676815), .D
		(n_287976818), .Z(n_304276981));
	notech_ao4 i_185433299(.A(n_296376902), .B(n_28012), .C(n_232376262), .D
		(\nbus_11365[27] ), .Z(n_304476983));
	notech_ao4 i_185233301(.A(n_227976218), .B(n_30010), .C(n_308547770), .D
		(n_28904), .Z(n_304676985));
	notech_and4 i_185633297(.A(n_304676985), .B(n_304476983), .C(n_287276811
		), .D(n_287576814), .Z(n_304876987));
	notech_ao4 i_184833304(.A(n_18756873), .B(n_28874), .C(n_23059), .D(n_27937
		), .Z(n_304976988));
	notech_ao4 i_184733305(.A(n_27879), .B(n_28765), .C(n_1877), .D(n_28828)
		, .Z(n_305176990));
	notech_and4 i_185733296(.A(n_304976988), .B(n_305176990), .C(n_304876987
		), .D(n_286976808), .Z(n_305376992));
	notech_ao4 i_184333309(.A(n_23009), .B(n_28798), .C(n_23003), .D(\nbus_11358[27] 
		), .Z(n_305476993));
	notech_ao4 i_184133311(.A(n_23023), .B(n_27672), .C(n_23019), .D(n_27536
		), .Z(n_305676995));
	notech_and4 i_184533307(.A(n_305676995), .B(n_305476993), .C(n_286176800
		), .D(n_286476803), .Z(n_305876997));
	notech_ao4 i_183833314(.A(n_23940), .B(n_30009), .C(n_23029), .D(n_28713
		), .Z(n_305976998));
	notech_and4 i_184033312(.A(n_3901), .B(n_305976998), .C(n_285576794), .D
		(n_285876797), .Z(n_306277001));
	notech_ao4 i_183333319(.A(n_296376902), .B(n_28011), .C(n_232176260), .D
		(\nbus_11365[26] ), .Z(n_306477003));
	notech_ao4 i_183133321(.A(n_57379), .B(n_30008), .C(n_308547770), .D(n_28903
		), .Z(n_306677005));
	notech_and4 i_183533317(.A(n_306677005), .B(n_306477003), .C(n_285176790
		), .D(n_285476793), .Z(n_306877007));
	notech_ao4 i_182833324(.A(n_18756873), .B(n_28873), .C(n_23059), .D(n_27936
		), .Z(n_306977008));
	notech_ao4 i_182733325(.A(n_27879), .B(n_28764), .C(n_1877), .D(n_28827)
		, .Z(n_307177010));
	notech_and4 i_183633316(.A(n_306977008), .B(n_307177010), .C(n_306877007
		), .D(n_284876787), .Z(n_307377012));
	notech_ao4 i_182333329(.A(n_23009), .B(n_28797), .C(n_23003), .D(\nbus_11358[26] 
		), .Z(n_307477013));
	notech_ao4 i_182133331(.A(n_23023), .B(n_27671), .C(n_23019), .D(n_27534
		), .Z(n_307677015));
	notech_and4 i_182533327(.A(n_307677015), .B(n_307477013), .C(n_284076779
		), .D(n_284376782), .Z(n_307877017));
	notech_ao4 i_181833334(.A(n_23940), .B(n_30007), .C(n_23029), .D(n_28712
		), .Z(n_307977018));
	notech_and4 i_182033332(.A(n_3901), .B(n_307977018), .C(n_283476773), .D
		(n_283776776), .Z(n_308277021));
	notech_ao4 i_181333339(.A(n_296376902), .B(n_28010), .C(n_231976258), .D
		(n_57771), .Z(n_308477023));
	notech_ao4 i_181133341(.A(n_57379), .B(n_30006), .C(n_308547770), .D(n_28902
		), .Z(n_308677025));
	notech_and4 i_181533337(.A(n_308677025), .B(n_308477023), .C(n_283076769
		), .D(n_283376772), .Z(n_308877027));
	notech_ao4 i_180833344(.A(n_18756873), .B(n_28872), .C(n_23059), .D(n_27935
		), .Z(n_308977028));
	notech_ao4 i_180733345(.A(n_27879), .B(n_28763), .C(n_1877), .D(n_28826)
		, .Z(n_309177030));
	notech_and4 i_181633336(.A(n_308977028), .B(n_309177030), .C(n_308877027
		), .D(n_282776766), .Z(n_309377032));
	notech_ao4 i_180333349(.A(n_23009), .B(n_28796), .C(n_23003), .D(n_55965
		), .Z(n_309477033));
	notech_ao4 i_180133351(.A(n_23023), .B(n_27670), .C(n_23019), .D(n_27533
		), .Z(n_309677035));
	notech_and4 i_180533347(.A(n_309677035), .B(n_309477033), .C(n_281976758
		), .D(n_282276761), .Z(n_309877037));
	notech_ao4 i_179833354(.A(n_23940), .B(n_30005), .C(n_23029), .D(n_28711
		), .Z(n_309977038));
	notech_and4 i_180033352(.A(n_3901), .B(n_309977038), .C(n_281376752), .D
		(n_281676755), .Z(n_310277041));
	notech_ao4 i_179333359(.A(n_296376902), .B(n_28009), .C(n_231776256), .D
		(n_57761), .Z(n_310477043));
	notech_ao4 i_179133361(.A(n_57379), .B(n_30004), .C(n_308547770), .D(n_28901
		), .Z(n_310677045));
	notech_and4 i_179533357(.A(n_310677045), .B(n_310477043), .C(n_280976748
		), .D(n_281276751), .Z(n_310877047));
	notech_ao4 i_178833364(.A(n_18756873), .B(n_28867), .C(n_23059), .D(n_27934
		), .Z(n_310977048));
	notech_ao4 i_178733365(.A(n_27879), .B(n_28762), .C(n_1877), .D(n_28825)
		, .Z(n_311177050));
	notech_and4 i_179633356(.A(n_310977048), .B(n_311177050), .C(n_310877047
		), .D(n_280676745), .Z(n_311377052));
	notech_ao4 i_178333369(.A(n_23009), .B(n_28795), .C(n_23003), .D(n_56475
		), .Z(n_311477053));
	notech_ao4 i_178133371(.A(n_23023), .B(n_27669), .C(n_23019), .D(n_27532
		), .Z(n_311677055));
	notech_and4 i_178533367(.A(n_311677055), .B(n_311477053), .C(n_279876737
		), .D(n_280176740), .Z(n_311877057));
	notech_ao4 i_177833374(.A(n_23940), .B(n_30003), .C(n_23029), .D(n_28710
		), .Z(n_311977058));
	notech_and4 i_178033372(.A(n_3901), .B(n_311977058), .C(n_279276731), .D
		(n_279576734), .Z(n_312277061));
	notech_ao4 i_177233379(.A(n_296376902), .B(n_28008), .C(n_231576254), .D
		(n_57751), .Z(n_312477063));
	notech_ao4 i_177033381(.A(n_57379), .B(n_30002), .C(n_308547770), .D(n_28900
		), .Z(n_312677065));
	notech_and4 i_177433377(.A(n_312677065), .B(n_312477063), .C(n_278876727
		), .D(n_279176730), .Z(n_312877067));
	notech_ao4 i_176733384(.A(n_18756873), .B(n_28863), .C(n_23059), .D(n_27933
		), .Z(n_312977068));
	notech_ao4 i_176633385(.A(n_27879), .B(n_28761), .C(n_1877), .D(n_28824)
		, .Z(n_313177070));
	notech_and4 i_177533376(.A(n_312977068), .B(n_313177070), .C(n_312877067
		), .D(n_278576724), .Z(n_313377072));
	notech_ao4 i_176233389(.A(n_23009), .B(n_28794), .C(n_23003), .D(n_56347
		), .Z(n_313477073));
	notech_ao4 i_176033391(.A(n_23023), .B(n_27668), .C(n_23019), .D(n_27531
		), .Z(n_313677075));
	notech_and4 i_176433387(.A(n_313677075), .B(n_313477073), .C(n_277776716
		), .D(n_278076719), .Z(n_313877077));
	notech_ao4 i_175733394(.A(n_23940), .B(n_30001), .C(n_23029), .D(n_28709
		), .Z(n_313977078));
	notech_and4 i_175933392(.A(n_3901), .B(n_313977078), .C(n_277176710), .D
		(n_277476713), .Z(n_314277081));
	notech_ao4 i_175233399(.A(n_296376902), .B(n_28007), .C(n_231376252), .D
		(n_57742), .Z(n_314477083));
	notech_ao4 i_175033401(.A(n_57379), .B(n_30000), .C(n_308547770), .D(n_28899
		), .Z(n_314677085));
	notech_and4 i_175433397(.A(n_314677085), .B(n_314477083), .C(n_276776706
		), .D(n_277076709), .Z(n_314877087));
	notech_ao4 i_174733404(.A(n_18756873), .B(n_28861), .C(n_23059), .D(n_27932
		), .Z(n_314977088));
	notech_ao4 i_174633405(.A(n_27879), .B(n_28760), .C(n_1877), .D(n_28823)
		, .Z(n_315177090));
	notech_and4 i_175533396(.A(n_314977088), .B(n_315177090), .C(n_314877087
		), .D(n_276476703), .Z(n_315377092));
	notech_ao4 i_174233409(.A(n_23009), .B(n_28793), .C(n_23003), .D(n_56338
		), .Z(n_315477093));
	notech_ao4 i_174033411(.A(n_23023), .B(n_27667), .C(n_23019), .D(n_27530
		), .Z(n_315677095));
	notech_and4 i_174433407(.A(n_315677095), .B(n_315477093), .C(n_275676695
		), .D(n_275976698), .Z(n_315877097));
	notech_ao4 i_173733414(.A(n_23940), .B(n_29999), .C(n_23029), .D(n_28708
		), .Z(n_315977098));
	notech_and4 i_173933412(.A(n_3901), .B(n_315977098), .C(n_275076689), .D
		(n_275376692), .Z(n_316277101));
	notech_ao4 i_173233419(.A(n_296376902), .B(n_28006), .C(n_231176250), .D
		(n_57733), .Z(n_316477103));
	notech_ao4 i_173033421(.A(n_57379), .B(n_29998), .C(n_308547770), .D(n_28898
		), .Z(n_316677105));
	notech_and4 i_173433417(.A(n_316677105), .B(n_316477103), .C(n_274676685
		), .D(n_274976688), .Z(n_316877107));
	notech_ao4 i_172733424(.A(n_18756873), .B(n_28859), .C(n_23059), .D(n_27931
		), .Z(n_316977108));
	notech_ao4 i_172633425(.A(n_27879), .B(n_28759), .C(n_1877), .D(n_28822)
		, .Z(n_317177110));
	notech_and4 i_173533416(.A(n_316977108), .B(n_317177110), .C(n_316877107
		), .D(n_274376682), .Z(n_317377112));
	notech_ao4 i_172233429(.A(n_23009), .B(n_28792), .C(n_23003), .D(n_56329
		), .Z(n_317477113));
	notech_ao4 i_172033431(.A(n_23023), .B(n_27666), .C(n_23019), .D(n_27529
		), .Z(n_317677115));
	notech_and4 i_172433427(.A(n_317677115), .B(n_317477113), .C(n_273576674
		), .D(n_273876677), .Z(n_317877117));
	notech_ao4 i_171633434(.A(n_23940), .B(n_29997), .C(n_23029), .D(n_28707
		), .Z(n_317977118));
	notech_and4 i_171833432(.A(n_3901), .B(n_317977118), .C(n_272976668), .D
		(n_273276671), .Z(n_318277121));
	notech_ao4 i_171133439(.A(n_296376902), .B(n_28005), .C(n_230976248), .D
		(n_57720), .Z(n_318477123));
	notech_ao4 i_170933441(.A(n_227976218), .B(n_29996), .C(n_308547770), .D
		(n_28897), .Z(n_318677125));
	notech_and4 i_171333437(.A(n_318677125), .B(n_318477123), .C(n_272576664
		), .D(n_272876667), .Z(n_318877127));
	notech_ao4 i_170633444(.A(n_18756873), .B(n_28858), .C(n_23059), .D(n_27930
		), .Z(n_318977128));
	notech_ao4 i_170533445(.A(n_27879), .B(n_28758), .C(n_1877), .D(n_28821)
		, .Z(n_319177130));
	notech_and4 i_171433436(.A(n_318977128), .B(n_319177130), .C(n_318877127
		), .D(n_272276661), .Z(n_319377132));
	notech_ao4 i_170133449(.A(n_23009), .B(n_28791), .C(n_23003), .D(n_56320
		), .Z(n_319477133));
	notech_ao4 i_169933451(.A(n_23023), .B(n_27665), .C(n_23019), .D(n_27528
		), .Z(n_319677135));
	notech_and4 i_170333447(.A(n_319677135), .B(n_319477133), .C(n_271476653
		), .D(n_271776656), .Z(n_319877137));
	notech_ao4 i_169633454(.A(n_23940), .B(n_29995), .C(n_23029), .D(n_28706
		), .Z(n_319977138));
	notech_and4 i_169833452(.A(n_3901), .B(n_319977138), .C(n_270876647), .D
		(n_271176650), .Z(n_320277141));
	notech_ao4 i_169033459(.A(n_57177), .B(n_28004), .C(n_230776246), .D(n_57707
		), .Z(n_320477143));
	notech_ao4 i_168833461(.A(n_227976218), .B(n_29994), .C(n_308547770), .D
		(n_28896), .Z(n_320677145));
	notech_and4 i_169333457(.A(n_320677145), .B(n_320477143), .C(n_270476643
		), .D(n_270776646), .Z(n_320877147));
	notech_ao4 i_168533464(.A(n_18756873), .B(n_28856), .C(n_23059), .D(n_27929
		), .Z(n_320977148));
	notech_ao4 i_168433465(.A(n_27879), .B(n_28757), .C(n_1877), .D(n_28820)
		, .Z(n_321177150));
	notech_and4 i_169433456(.A(n_320977148), .B(n_321177150), .C(n_320877147
		), .D(n_270176640), .Z(n_321377152));
	notech_ao4 i_168033469(.A(n_23009), .B(n_28790), .C(n_23003), .D(n_56311
		), .Z(n_321477153));
	notech_ao4 i_167833471(.A(n_23023), .B(n_27664), .C(n_23019), .D(n_27527
		), .Z(n_321677155));
	notech_and4 i_168233467(.A(n_321677155), .B(n_321477153), .C(n_269376632
		), .D(n_269676635), .Z(n_321877157));
	notech_ao4 i_167533474(.A(n_23940), .B(n_29991), .C(n_23029), .D(n_28705
		), .Z(n_321977158));
	notech_and4 i_167733472(.A(n_3901), .B(n_321977158), .C(n_268776626), .D
		(n_269076629), .Z(n_322277161));
	notech_ao4 i_167033479(.A(n_57177), .B(n_28003), .C(n_230576244), .D(n_57698
		), .Z(n_322477163));
	notech_ao4 i_166833481(.A(n_227976218), .B(n_29988), .C(n_308547770), .D
		(n_28895), .Z(n_322677165));
	notech_and4 i_167233477(.A(n_322677165), .B(n_322477163), .C(n_268376622
		), .D(n_268676625), .Z(n_322877167));
	notech_ao4 i_166533484(.A(n_18756873), .B(n_28855), .C(n_23059), .D(n_27928
		), .Z(n_322977168));
	notech_ao4 i_166433485(.A(n_27879), .B(n_28756), .C(n_1877), .D(n_28819)
		, .Z(n_323177170));
	notech_and4 i_167333476(.A(n_322977168), .B(n_323177170), .C(n_322877167
		), .D(n_268076619), .Z(n_323377172));
	notech_ao4 i_166033489(.A(n_23009), .B(n_28789), .C(n_23003), .D(n_56302
		), .Z(n_323477173));
	notech_ao4 i_165833491(.A(n_55764), .B(n_27663), .C(n_23019), .D(n_27526
		), .Z(n_323677175));
	notech_and4 i_166233487(.A(n_323677175), .B(n_323477173), .C(n_267276611
		), .D(n_267576614), .Z(n_323877177));
	notech_ao4 i_165533494(.A(n_23940), .B(n_29987), .C(n_23029), .D(n_28704
		), .Z(n_323977178));
	notech_and4 i_165733492(.A(n_57948), .B(n_323977178), .C(n_266676605), .D
		(n_266976608), .Z(n_324277181));
	notech_ao4 i_164933499(.A(n_57177), .B(n_28002), .C(n_230376242), .D(n_57689
		), .Z(n_324477183));
	notech_ao4 i_164733501(.A(n_227976218), .B(n_29986), .C(n_308547770), .D
		(n_28894), .Z(n_324677185));
	notech_and4 i_165233497(.A(n_324677185), .B(n_324477183), .C(n_266276601
		), .D(n_266576604), .Z(n_324877187));
	notech_ao4 i_164333504(.A(n_18756873), .B(n_28854), .C(n_23059), .D(n_27927
		), .Z(n_324977188));
	notech_ao4 i_164233505(.A(n_27879), .B(n_28755), .C(n_1877), .D(n_28818)
		, .Z(n_325177190));
	notech_and4 i_165333496(.A(n_324977188), .B(n_325177190), .C(n_324877187
		), .D(n_265976598), .Z(n_325377192));
	notech_ao4 i_163833509(.A(n_23009), .B(n_28788), .C(n_23003), .D(n_56293
		), .Z(n_325477193));
	notech_ao4 i_163633511(.A(n_55764), .B(n_27662), .C(n_23019), .D(n_27525
		), .Z(n_325677195));
	notech_and4 i_164033507(.A(n_325677195), .B(n_325477193), .C(n_265176590
		), .D(n_265476593), .Z(n_325877197));
	notech_ao4 i_163333514(.A(n_23940), .B(n_29985), .C(n_57920), .D(n_28703
		), .Z(n_325977198));
	notech_and4 i_163533512(.A(n_57948), .B(n_325977198), .C(n_264576584), .D
		(n_264876587), .Z(n_326277201));
	notech_ao4 i_162833519(.A(n_57177), .B(n_28001), .C(n_230176240), .D(\nbus_11365[16] 
		), .Z(n_326477203));
	notech_ao4 i_162633521(.A(n_227976218), .B(n_29983), .C(n_308547770), .D
		(n_28893), .Z(n_326677205));
	notech_and4 i_163033517(.A(n_326677205), .B(n_326477203), .C(n_264176580
		), .D(n_264476583), .Z(n_326877207));
	notech_ao4 i_162333524(.A(n_18756873), .B(n_28852), .C(n_23059), .D(n_27926
		), .Z(n_326977208));
	notech_ao4 i_162233525(.A(n_27879), .B(n_28754), .C(n_1877), .D(n_28817)
		, .Z(n_327177210));
	notech_and4 i_163133516(.A(n_326977208), .B(n_327177210), .C(n_326877207
		), .D(n_263876577), .Z(n_327377212));
	notech_ao4 i_161833529(.A(n_23009), .B(n_28787), .C(n_23003), .D(\nbus_11358[16] 
		), .Z(n_327477213));
	notech_ao4 i_161633531(.A(n_55764), .B(n_27661), .C(n_23019), .D(n_28682
		), .Z(n_327677215));
	notech_and4 i_162033527(.A(n_327677215), .B(n_327477213), .C(n_263076569
		), .D(n_263376572), .Z(n_327877217));
	notech_ao4 i_161333534(.A(n_23940), .B(n_29982), .C(n_57920), .D(n_28702
		), .Z(n_327977218));
	notech_and4 i_161533532(.A(n_57948), .B(n_327977218), .C(n_262476563), .D
		(n_262776566), .Z(n_328277221));
	notech_or4 i_4835062(.A(n_32729), .B(n_25625), .C(n_59435), .D(n_60229),
		 .Z(n_328577224));
	notech_ao4 i_160733540(.A(n_328577224), .B(\nbus_11365[31] ), .C(n_229876237
		), .D(\nbus_11307[15] ), .Z(n_328677225));
	notech_or4 i_4735063(.A(n_27907), .B(n_59435), .C(n_26782), .D(n_60229),
		 .Z(n_328777226));
	notech_ao4 i_160633541(.A(n_3903), .B(n_56100), .C(n_328777226), .D(n_28678
		), .Z(n_328877227));
	notech_ao4 i_160433543(.A(n_57177), .B(n_28000), .C(n_3902), .D(\nbus_11358[7] 
		), .Z(n_329077229));
	notech_ao4 i_160333544(.A(n_57538), .B(nbus_11295[15]), .C(n_57524), .D(n_27923
		), .Z(n_329177230));
	notech_and4 i_160933538(.A(n_329177230), .B(n_329077229), .C(n_328877227
		), .D(n_328677225), .Z(n_329377232));
	notech_ao4 i_160033547(.A(n_57848), .B(\nbus_11358[15] ), .C(n_57165), .D
		(\nbus_11307[7] ), .Z(n_329477233));
	notech_ao4 i_159933548(.A(n_57498), .B(n_29754), .C(n_18756873), .D(n_28850
		), .Z(n_329577234));
	notech_ao4 i_159733550(.A(n_22571), .B(\nbus_11358[31] ), .C(n_57512), .D
		(n_28816), .Z(n_329777236));
	notech_and4 i_160233545(.A(n_329777236), .B(n_329577234), .C(n_329477233
		), .D(n_261176550), .Z(n_329977238));
	notech_ao4 i_159333554(.A(n_55764), .B(n_27660), .C(n_57859), .D(n_27524
		), .Z(n_330177240));
	notech_ao4 i_159233555(.A(n_57920), .B(n_28701), .C(n_23031), .D(n_27690
		), .Z(n_330277241));
	notech_ao4 i_159033557(.A(n_23040), .B(n_28697), .C(n_55773), .D(n_29981
		), .Z(n_330477243));
	notech_ao4 i_158933558(.A(n_22585), .B(n_28924), .C(n_22572), .D(n_28667
		), .Z(n_330577244));
	notech_and4 i_159533552(.A(n_330577244), .B(n_330477243), .C(n_330277241
		), .D(n_330177240), .Z(n_330777246));
	notech_ao4 i_158633561(.A(n_22582), .B(n_28648), .C(n_22579), .D(n_28892
		), .Z(n_330877247));
	notech_ao4 i_158533562(.A(n_22591), .B(n_28753), .C(n_22590), .D(n_29980
		), .Z(n_330977248));
	notech_ao4 i_158333564(.A(n_28076), .B(n_29979), .C(n_22594), .D(n_28786
		), .Z(n_331177250));
	notech_and4 i_158833559(.A(n_57948), .B(n_331177250), .C(n_330977248), .D
		(n_330877247), .Z(n_331377252));
	notech_ao4 i_157933568(.A(n_328577224), .B(\nbus_11365[30] ), .C(n_229676235
		), .D(n_57662), .Z(n_331577254));
	notech_ao4 i_157833569(.A(n_3903), .B(n_27989), .C(n_328777226), .D(n_28677
		), .Z(n_331677255));
	notech_ao4 i_157533571(.A(n_57177), .B(n_27999), .C(n_3902), .D(n_56082)
		, .Z(n_331877257));
	notech_ao4 i_157433572(.A(n_57165), .B(n_57592), .C(n_57524), .D(n_27918
		), .Z(n_331977258));
	notech_and4 i_158133566(.A(n_331977258), .B(n_331877257), .C(n_331677255
		), .D(n_331577254), .Z(n_332177260));
	notech_ao4 i_157133575(.A(n_57498), .B(n_56257), .C(n_57121), .D(n_28849
		), .Z(n_332277261));
	notech_ao4 i_157033576(.A(n_57848), .B(\nbus_11358[14] ), .C(n_57512), .D
		(n_28815), .Z(n_332377262));
	notech_ao4 i_156833578(.A(n_57859), .B(n_27523), .C(n_27781), .D(n_28736
		), .Z(n_332577264));
	notech_and4 i_157333573(.A(n_332577264), .B(n_332377262), .C(n_332277261
		), .D(n_258276521), .Z(n_332777266));
	notech_ao4 i_156433582(.A(n_57920), .B(n_28700), .C(n_23031), .D(n_27689
		), .Z(n_332977268));
	notech_ao4 i_156333583(.A(n_57538), .B(nbus_11295[14]), .C(n_55773), .D(n_29978
		), .Z(n_333077269));
	notech_ao4 i_156133585(.A(n_22571), .B(\nbus_11358[30] ), .C(n_23040), .D
		(n_28696), .Z(n_333277271));
	notech_ao4 i_156033586(.A(n_22585), .B(n_28923), .C(n_22572), .D(n_28666
		), .Z(n_333377272));
	notech_and4 i_156633580(.A(n_333377272), .B(n_333277271), .C(n_333077269
		), .D(n_332977268), .Z(n_333577274));
	notech_ao4 i_155733589(.A(n_22582), .B(n_28647), .C(n_22579), .D(n_28891
		), .Z(n_333677275));
	notech_ao4 i_155633590(.A(n_22591), .B(n_28752), .C(n_22590), .D(n_29977
		), .Z(n_333777276));
	notech_ao4 i_155433592(.A(n_28076), .B(n_29976), .C(n_22594), .D(n_28785
		), .Z(n_333977278));
	notech_and4 i_155933587(.A(n_57948), .B(n_333977278), .C(n_333777276), .D
		(n_333677275), .Z(n_334177280));
	notech_ao4 i_155033596(.A(n_328577224), .B(\nbus_11365[29] ), .C(n_229476233
		), .D(\nbus_11307[13] ), .Z(n_334377282));
	notech_ao4 i_154933597(.A(n_3903), .B(n_27987), .C(n_328777226), .D(n_28676
		), .Z(n_334477283));
	notech_ao4 i_154733599(.A(n_57177), .B(n_27998), .C(n_3902), .D(\nbus_11358[5] 
		), .Z(n_334677285));
	notech_ao4 i_154633600(.A(n_57165), .B(\nbus_11307[5] ), .C(n_57524), .D
		(n_27916), .Z(n_334777286));
	notech_and4 i_155233594(.A(n_334777286), .B(n_334677285), .C(n_334477283
		), .D(n_334377282), .Z(n_334977288));
	notech_ao4 i_154333603(.A(n_57498), .B(n_29592), .C(n_57121), .D(n_28847
		), .Z(n_335077289));
	notech_ao4 i_154233604(.A(n_57848), .B(\nbus_11358[13] ), .C(n_57512), .D
		(n_28814), .Z(n_335177290));
	notech_ao4 i_154033606(.A(n_57859), .B(n_27522), .C(n_27781), .D(n_28735
		), .Z(n_335377292));
	notech_and4 i_154533601(.A(n_335377292), .B(n_335177290), .C(n_335077289
		), .D(n_255376492), .Z(n_335577294));
	notech_ao4 i_153633610(.A(n_57920), .B(n_28699), .C(n_23031), .D(n_27688
		), .Z(n_335777296));
	notech_ao4 i_153533611(.A(nbus_11295[13]), .B(n_57538), .C(n_55773), .D(n_29975
		), .Z(n_335877297));
	notech_ao4 i_153333613(.A(n_22571), .B(\nbus_11358[29] ), .C(n_23040), .D
		(n_28695), .Z(n_336077299));
	notech_ao4 i_153233614(.A(n_22585), .B(n_28922), .C(n_22572), .D(n_28665
		), .Z(n_336177300));
	notech_and4 i_153833608(.A(n_336177300), .B(n_336077299), .C(n_335877297
		), .D(n_335777296), .Z(n_336377302));
	notech_ao4 i_152933617(.A(n_22582), .B(n_28645), .C(n_22579), .D(n_28890
		), .Z(n_336477303));
	notech_ao4 i_152833618(.A(n_22591), .B(n_28751), .C(n_22590), .D(n_29974
		), .Z(n_336577304));
	notech_ao4 i_152633620(.A(n_28076), .B(n_29973), .C(n_22594), .D(n_28784
		), .Z(n_336777306));
	notech_and4 i_153133615(.A(n_57948), .B(n_336777306), .C(n_336577304), .D
		(n_336477303), .Z(n_336977308));
	notech_ao4 i_152233624(.A(n_328577224), .B(\nbus_11365[28] ), .C(n_229276231
		), .D(n_57644), .Z(n_337177310));
	notech_ao4 i_152133625(.A(n_3903), .B(n_27986), .C(n_328777226), .D(n_28675
		), .Z(n_337277311));
	notech_ao4 i_151933627(.A(n_57177), .B(n_27997), .C(n_3902), .D(\nbus_11358[4] 
		), .Z(n_337477313));
	notech_ao4 i_151833628(.A(n_57165), .B(\nbus_11307[4] ), .C(n_57524), .D
		(n_27915), .Z(n_337577314));
	notech_and4 i_152433622(.A(n_337577314), .B(n_337477313), .C(n_337277311
		), .D(n_337177310), .Z(n_337777316));
	notech_ao4 i_151433631(.A(n_57498), .B(n_29679), .C(n_57121), .D(n_28846
		), .Z(n_337877317));
	notech_ao4 i_151233632(.A(n_57848), .B(n_56221), .C(n_57512), .D(n_28813
		), .Z(n_337977318));
	notech_ao4 i_151033634(.A(n_57859), .B(n_27521), .C(n_27781), .D(n_28733
		), .Z(n_338177320));
	notech_and4 i_151733629(.A(n_338177320), .B(n_337977318), .C(n_337877317
		), .D(n_252476463), .Z(n_338377322));
	notech_ao4 i_150633638(.A(n_57920), .B(n_28698), .C(n_23031), .D(n_27687
		), .Z(n_338577324));
	notech_ao4 i_150533639(.A(n_57538), .B(nbus_11295[12]), .C(n_55773), .D(n_29972
		), .Z(n_338677325));
	notech_ao4 i_150333641(.A(n_22571), .B(\nbus_11358[28] ), .C(n_23040), .D
		(n_28694), .Z(n_338877327));
	notech_ao4 i_150233642(.A(n_22585), .B(n_28921), .C(n_22572), .D(n_28664
		), .Z(n_338977328));
	notech_and4 i_150833636(.A(n_338977328), .B(n_338877327), .C(n_338677325
		), .D(n_338577324), .Z(n_339177330));
	notech_ao4 i_149933645(.A(n_22582), .B(n_28644), .C(n_22579), .D(n_28889
		), .Z(n_339277331));
	notech_ao4 i_149833646(.A(n_22591), .B(n_28750), .C(n_22590), .D(n_29971
		), .Z(n_339377332));
	notech_ao4 i_149633648(.A(n_28076), .B(n_29970), .C(n_22594), .D(n_28783
		), .Z(n_339577334));
	notech_and4 i_150133643(.A(n_57948), .B(n_339577334), .C(n_339377332), .D
		(n_339277331), .Z(n_339777336));
	notech_ao4 i_149233652(.A(n_328577224), .B(\nbus_11365[27] ), .C(n_229076229
		), .D(\nbus_11307[11] ), .Z(n_339977338));
	notech_ao4 i_149133653(.A(n_3903), .B(n_59223), .C(n_328777226), .D(n_28674
		), .Z(n_340077339));
	notech_ao4 i_148933655(.A(n_57177), .B(n_27996), .C(n_3902), .D(\nbus_11358[3] 
		), .Z(n_340277341));
	notech_ao4 i_148833656(.A(n_57165), .B(\nbus_11307[3] ), .C(n_57524), .D
		(n_27914), .Z(n_340377342));
	notech_and4 i_149433650(.A(n_340377342), .B(n_340277341), .C(n_340077339
		), .D(n_339977338), .Z(n_340577344));
	notech_ao4 i_148533659(.A(n_57498), .B(n_29596), .C(n_57121), .D(n_28845
		), .Z(n_340677345));
	notech_ao4 i_148433660(.A(n_57848), .B(\nbus_11358[11] ), .C(n_57512), .D
		(n_28812), .Z(n_340777346));
	notech_ao4 i_148233662(.A(n_57859), .B(n_27520), .C(n_27781), .D(n_28732
		), .Z(n_340977348));
	notech_and4 i_148733657(.A(n_340977348), .B(n_340777346), .C(n_340677345
		), .D(n_249576434), .Z(n_341177350));
	notech_ao4 i_147833666(.A(n_57920), .B(n_27699), .C(n_23031), .D(n_27686
		), .Z(n_341377352));
	notech_ao4 i_147733667(.A(n_57538), .B(nbus_11295[11]), .C(n_55773), .D(n_29969
		), .Z(n_341477353));
	notech_ao4 i_147533669(.A(n_22571), .B(\nbus_11358[27] ), .C(n_23040), .D
		(n_28693), .Z(n_341677355));
	notech_ao4 i_147433670(.A(n_22585), .B(n_28920), .C(n_22572), .D(n_28663
		), .Z(n_341777356));
	notech_and4 i_148033664(.A(n_341777356), .B(n_341677355), .C(n_341477353
		), .D(n_341377352), .Z(n_341977358));
	notech_ao4 i_147133673(.A(n_22582), .B(n_28643), .C(n_22579), .D(n_28888
		), .Z(n_342077359));
	notech_ao4 i_147033674(.A(n_22591), .B(n_28749), .C(n_22590), .D(n_29968
		), .Z(n_342177360));
	notech_ao4 i_146833676(.A(n_28076), .B(n_29966), .C(n_22594), .D(n_28781
		), .Z(n_342377362));
	notech_and4 i_147333671(.A(n_57948), .B(n_342377362), .C(n_342177360), .D
		(n_342077359), .Z(n_342577364));
	notech_ao4 i_146433680(.A(n_328577224), .B(\nbus_11365[26] ), .C(n_228876227
		), .D(\nbus_11307[10] ), .Z(n_342777366));
	notech_ao4 i_146333681(.A(n_3903), .B(n_59259), .C(n_328777226), .D(n_28673
		), .Z(n_342877367));
	notech_ao4 i_146133683(.A(n_57177), .B(n_27993), .C(n_3902), .D(n_55992)
		, .Z(n_343077369));
	notech_ao4 i_146033684(.A(n_57165), .B(n_57552), .C(n_57524), .D(n_27913
		), .Z(n_343177370));
	notech_and4 i_146633678(.A(n_343177370), .B(n_343077369), .C(n_342877367
		), .D(n_342777366), .Z(n_343377372));
	notech_ao4 i_145733687(.A(n_57498), .B(n_29684), .C(n_57121), .D(n_28844
		), .Z(n_343477373));
	notech_ao4 i_145633688(.A(n_57848), .B(\nbus_11358[10] ), .C(n_57512), .D
		(n_28811), .Z(n_343577374));
	notech_ao4 i_145433690(.A(n_57859), .B(n_27519), .C(n_27781), .D(n_28730
		), .Z(n_343777376));
	notech_and4 i_145933685(.A(n_343777376), .B(n_343577374), .C(n_343477373
		), .D(n_246676405), .Z(n_343977378));
	notech_ao4 i_145033694(.A(n_57920), .B(n_27698), .C(n_23031), .D(n_27685
		), .Z(n_344177380));
	notech_ao4 i_144933695(.A(n_57533), .B(nbus_11295[10]), .C(n_55773), .D(n_29965
		), .Z(n_344277381));
	notech_ao4 i_144733697(.A(n_22571), .B(\nbus_11358[26] ), .C(n_23040), .D
		(n_28692), .Z(n_344477383));
	notech_ao4 i_144633698(.A(n_22585), .B(n_28919), .C(n_22572), .D(n_28662
		), .Z(n_344577384));
	notech_and4 i_145233692(.A(n_344577384), .B(n_344477383), .C(n_344277381
		), .D(n_344177380), .Z(n_344777386));
	notech_ao4 i_144333701(.A(n_22582), .B(n_28642), .C(n_22579), .D(n_28887
		), .Z(n_344877387));
	notech_ao4 i_144233702(.A(n_22591), .B(n_28748), .C(n_22590), .D(n_29964
		), .Z(n_344977388));
	notech_ao4 i_144033704(.A(n_28076), .B(n_29963), .C(n_22594), .D(n_28780
		), .Z(n_345177390));
	notech_and4 i_144533699(.A(n_57948), .B(n_345177390), .C(n_344977388), .D
		(n_344877387), .Z(n_345377392));
	notech_ao4 i_143633708(.A(n_328577224), .B(n_57771), .C(n_228676225), .D
		(\nbus_11307[9] ), .Z(n_345577394));
	notech_ao4 i_143533709(.A(n_3903), .B(n_27983), .C(n_328777226), .D(n_28672
		), .Z(n_345677395));
	notech_ao4 i_143333711(.A(n_57177), .B(n_27992), .C(n_3902), .D(\nbus_11358[1] 
		), .Z(n_345877397));
	notech_ao4 i_143233712(.A(n_57165), .B(\nbus_11307[1] ), .C(n_57524), .D
		(n_27912), .Z(n_345977398));
	notech_and4 i_143833706(.A(n_345977398), .B(n_345877397), .C(n_345677395
		), .D(n_345577394), .Z(n_346177400));
	notech_ao4 i_142933715(.A(n_57498), .B(n_29743), .C(n_57121), .D(n_28842
		), .Z(n_346277401));
	notech_ao4 i_142833716(.A(n_57848), .B(\nbus_11358[9] ), .C(n_57512), .D
		(n_28810), .Z(n_346377402));
	notech_ao4 i_142633718(.A(n_57859), .B(n_27518), .C(n_27781), .D(n_28729
		), .Z(n_346577404));
	notech_and4 i_143133713(.A(n_346577404), .B(n_346377402), .C(n_346277401
		), .D(n_243776376), .Z(n_346777406));
	notech_ao4 i_142233722(.A(n_57920), .B(n_27697), .C(n_23031), .D(n_27684
		), .Z(n_346977408));
	notech_ao4 i_142133723(.A(n_57533), .B(nbus_11295[9]), .C(n_55773), .D(n_29962
		), .Z(n_347077409));
	notech_ao4 i_141933725(.A(n_22571), .B(n_55965), .C(n_23040), .D(n_28691
		), .Z(n_347277411));
	notech_ao4 i_141833726(.A(n_22585), .B(n_28918), .C(n_22572), .D(n_28661
		), .Z(n_347377412));
	notech_and4 i_142433720(.A(n_347377412), .B(n_347277411), .C(n_347077409
		), .D(n_346977408), .Z(n_347577414));
	notech_ao4 i_141533729(.A(n_22582), .B(n_28641), .C(n_22579), .D(n_28886
		), .Z(n_347677415));
	notech_ao4 i_141433730(.A(n_22591), .B(n_28747), .C(n_22590), .D(n_29961
		), .Z(n_347777416));
	notech_ao4 i_141233732(.A(n_28076), .B(n_29960), .C(n_22594), .D(n_28779
		), .Z(n_347977418));
	notech_and4 i_141733727(.A(n_3901), .B(n_347977418), .C(n_347777416), .D
		(n_347677415), .Z(n_348177420));
	notech_ao4 i_140833736(.A(n_328577224), .B(n_57761), .C(n_228476223), .D
		(\nbus_11307[8] ), .Z(n_348377422));
	notech_ao4 i_140733737(.A(n_3903), .B(n_27981), .C(n_328777226), .D(n_28671
		), .Z(n_348477423));
	notech_ao4 i_140533739(.A(n_57177), .B(n_27991), .C(n_3902), .D(\nbus_11358[0] 
		), .Z(n_348677425));
	notech_ao4 i_140433740(.A(n_57165), .B(\nbus_11307[0] ), .C(n_57524), .D
		(n_27911), .Z(n_348777426));
	notech_and4 i_141033734(.A(n_348777426), .B(n_348677425), .C(n_348477423
		), .D(n_348377422), .Z(n_348977428));
	notech_ao4 i_140133743(.A(n_57498), .B(n_29787), .C(n_57121), .D(n_28840
		), .Z(n_349077429));
	notech_ao4 i_140033744(.A(n_57848), .B(\nbus_11358[8] ), .C(n_57512), .D
		(n_28809), .Z(n_349177430));
	notech_ao4 i_139833746(.A(n_57859), .B(n_27517), .C(n_27781), .D(n_28728
		), .Z(n_349377432));
	notech_and4 i_140333741(.A(n_349377432), .B(n_349177430), .C(n_349077429
		), .D(n_240876347), .Z(n_349577434));
	notech_ao4 i_139433750(.A(n_23029), .B(n_27696), .C(n_23031), .D(n_27683
		), .Z(n_349777436));
	notech_ao4 i_139333751(.A(n_57533), .B(nbus_11295[8]), .C(n_55773), .D(n_29959
		), .Z(n_349877437));
	notech_ao4 i_139133753(.A(n_22571), .B(n_56475), .C(n_23040), .D(n_28690
		), .Z(n_350077439));
	notech_ao4 i_139033754(.A(n_22585), .B(n_28917), .C(n_22572), .D(n_28660
		), .Z(n_350177440));
	notech_and4 i_139633748(.A(n_350177440), .B(n_350077439), .C(n_349877437
		), .D(n_349777436), .Z(n_350377442));
	notech_ao4 i_138733757(.A(n_22582), .B(n_28640), .C(n_22579), .D(n_28885
		), .Z(n_350477443));
	notech_ao4 i_138633758(.A(n_22591), .B(n_28746), .C(n_22590), .D(n_29958
		), .Z(n_350577444));
	notech_ao4 i_138433760(.A(n_28076), .B(n_29956), .C(n_22594), .D(n_28778
		), .Z(n_350777446));
	notech_and4 i_138933755(.A(n_57948), .B(n_350777446), .C(n_350577444), .D
		(n_350477443), .Z(n_350977448));
	notech_ao4 i_122733912(.A(n_22322), .B(n_307947775), .C(n_228276221), .D
		(\nbus_11307[1] ), .Z(n_351177450));
	notech_ao4 i_122533913(.A(n_57165), .B(\nbus_11307[9] ), .C(n_57524), .D
		(n_27898), .Z(n_351277451));
	notech_ao4 i_122333915(.A(n_57121), .B(n_28834), .C(n_57155), .D(\nbus_11358[9] 
		), .Z(n_351477453));
	notech_ao4 i_122233916(.A(n_57512), .B(n_28803), .C(n_57498), .D(n_29678
		), .Z(n_351577454));
	notech_and4 i_122933910(.A(n_351577454), .B(n_351477453), .C(n_351277451
		), .D(n_351177450), .Z(n_351777456));
	notech_ao4 i_121933919(.A(n_27781), .B(n_28719), .C(n_57848), .D(\nbus_11358[1] 
		), .Z(n_351877457));
	notech_ao4 i_121833920(.A(n_55764), .B(n_27654), .C(n_27512), .D(n_57859
		), .Z(n_351977458));
	notech_ao4 i_121633922(.A(n_57920), .B(n_27693), .C(n_23031), .D(n_27677
		), .Z(n_352177460));
	notech_and4 i_122133917(.A(n_352177460), .B(n_351977458), .C(n_351877457
		), .D(n_237976318), .Z(n_352377462));
	notech_ao4 i_121233926(.A(n_23040), .B(n_28684), .C(n_57533), .D(nbus_11295
		[1]), .Z(n_352577464));
	notech_ao4 i_121133927(.A(n_22572), .B(n_28650), .C(n_22571), .D(n_56293
		), .Z(n_352677465));
	notech_ao4 i_120933929(.A(n_22579), .B(n_28879), .C(n_22585), .D(n_28910
		), .Z(n_352877467));
	notech_and4 i_121433924(.A(n_352877467), .B(n_352677465), .C(n_352577464
		), .D(n_237276311), .Z(n_353077469));
	notech_ao4 i_120633932(.A(n_22591), .B(n_28739), .C(n_22590), .D(n_29955
		), .Z(n_353177470));
	notech_ao4 i_120533933(.A(n_28076), .B(n_29004), .C(n_22594), .D(n_28771
		), .Z(n_353277471));
	notech_ao4 i_120333935(.A(n_22309), .B(n_28626), .C(n_22313), .D(n_59241
		), .Z(n_353477473));
	notech_and4 i_120833930(.A(n_353477473), .B(n_353277471), .C(n_353177470
		), .D(n_236576304), .Z(n_353677475));
	notech_ao4 i_119833940(.A(n_57524), .B(n_27897), .C(\nbus_11307[0] ), .D
		(n_228176220), .Z(n_353977478));
	notech_ao4 i_119733941(.A(n_57155), .B(\nbus_11358[8] ), .C(n_57165), .D
		(\nbus_11307[8] ), .Z(n_354077479));
	notech_ao4 i_119533943(.A(n_57498), .B(n_56037), .C(n_57121), .D(n_28833
		), .Z(n_354277481));
	notech_and4 i_120033938(.A(n_354277481), .B(n_354077479), .C(n_353977478
		), .D(n_235776296), .Z(n_354477483));
	notech_ao4 i_119233946(.A(n_27781), .B(n_28718), .C(n_57848), .D(\nbus_11358[0] 
		), .Z(n_354577484));
	notech_ao4 i_119133947(.A(n_55764), .B(n_27653), .C(n_57859), .D(n_28680
		), .Z(n_354677485));
	notech_ao4 i_118733949(.A(n_57920), .B(n_27692), .C(n_23031), .D(n_27676
		), .Z(n_354877487));
	notech_and4 i_119433944(.A(n_354877487), .B(n_354677485), .C(n_354577484
		), .D(n_235076289), .Z(n_355077489));
	notech_ao4 i_118333953(.A(n_23040), .B(n_28683), .C(n_57533), .D(nbus_11295
		[0]), .Z(n_355277491));
	notech_ao4 i_118233954(.A(n_22572), .B(n_28649), .C(n_22571), .D(\nbus_11358[16] 
		), .Z(n_355377492));
	notech_ao4 i_118033956(.A(n_22579), .B(n_28878), .C(n_22585), .D(n_28909
		), .Z(n_355577494));
	notech_and4 i_118533951(.A(n_355577494), .B(n_355377492), .C(n_355277491
		), .D(n_234376282), .Z(n_355777496));
	notech_ao4 i_117733959(.A(n_22591), .B(n_28738), .C(n_22590), .D(n_29953
		), .Z(n_355877497));
	notech_ao4 i_117633960(.A(n_28076), .B(n_29003), .C(n_22594), .D(n_28770
		), .Z(n_355977498));
	notech_ao4 i_117433962(.A(n_22309), .B(n_28625), .C(n_22313), .D(n_27981
		), .Z(n_356177500));
	notech_and4 i_117933957(.A(n_356177500), .B(n_355977498), .C(n_355877497
		), .D(n_233676275), .Z(n_356377502));
	notech_or4 i_3121204(.A(n_117868195), .B(n_117975123), .C(n_119075134), 
		.D(n_26682), .Z(n_18660));
	notech_and4 i_821917(.A(n_119575139), .B(n_119775141), .C(n_117675120), 
		.D(n_120175145), .Z(n_17474));
	notech_and4 i_1617605(.A(n_120875152), .B(n_120775151), .C(n_116175105),
		 .D(n_121175155), .Z(n_16796));
	notech_and2 i_60658551(.A(n_311291711), .B(n_317891645), .Z(n_58411));
	notech_ao4 i_110258531(.A(n_32356), .B(n_303391790), .C(n_304291781), .D
		(n_56100), .Z(n_57947));
	notech_and3 i_115658529(.A(n_58530), .B(n_316691657), .C(n_199375932), .Z
		(n_57893));
	notech_nand2 i_153358518(.A(n_60229), .B(read_data[0]), .Z(n_57548));
	notech_and3 i_259958503(.A(n_23513), .B(n_23512), .C(n_54974), .Z(n_56516
		));
	notech_and4 i_821853(.A(n_138775331), .B(n_138975333), .C(n_137175315), 
		.D(n_139375337), .Z(n_20660));
	notech_nand2 i_521850(.A(n_140375347), .B(n_139875342), .Z(n_20642));
	notech_and4 i_221847(.A(n_141075354), .B(n_140975353), .C(n_134575289), 
		.D(n_141375357), .Z(n_20624));
	notech_nand2 i_221911(.A(n_142575369), .B(n_142075364), .Z(n_17438));
	notech_and4 i_121910(.A(n_143175375), .B(n_143075374), .C(n_143975383), 
		.D(n_142975373), .Z(n_17432));
	notech_and4 i_1217601(.A(n_144175385), .B(n_144375387), .C(n_144875392),
		 .D(n_131475258), .Z(n_16772));
	notech_and4 i_1117600(.A(n_129875242), .B(n_145575399), .C(n_145475398),
		 .D(n_145875402), .Z(n_16766));
	notech_and4 i_1017599(.A(n_146775411), .B(n_146675410), .C(n_146575409),
		 .D(n_147075414), .Z(n_16760));
	notech_and4 i_817597(.A(n_147375417), .B(n_147575419), .C(n_128175225), 
		.D(n_148075424), .Z(n_16748));
	notech_and4 i_517594(.A(n_148975433), .B(n_148875432), .C(n_148775431), 
		.D(n_149275436), .Z(n_16730));
	notech_nand2 i_217591(.A(n_150675450), .B(n_150075444), .Z(n_16712));
	notech_and4 i_117590(.A(n_151675460), .B(n_151575459), .C(n_151475458), 
		.D(n_152075464), .Z(n_16706));
	notech_nand2 i_4058451(.A(read_data[1]), .B(n_60229), .Z(n_276234718));
	notech_and2 i_9858393(.A(n_58514), .B(n_122975173), .Z(n_57892));
	notech_and3 i_189161792(.A(n_304691777), .B(n_285363120), .C(n_164361926
		), .Z(n_251362780));
	notech_or4 i_121846(.A(n_152975473), .B(n_155475498), .C(n_26685), .D(n_26684
		), .Z(n_20618));
	notech_mux2 i_2311692(.S(n_60550), .A(regs_14[22]), .B(add_len_pc32[22])
		, .Z(add_len_pc[22]));
	notech_mux2 i_2411693(.S(n_60550), .A(regs_14[23]), .B(add_len_pc32[23])
		, .Z(add_len_pc[23]));
	notech_mux2 i_2511694(.S(n_60550), .A(regs_14[24]), .B(add_len_pc32[24])
		, .Z(add_len_pc[24]));
	notech_nand2 i_2520718(.A(n_174075684), .B(n_173575679), .Z(n_24900));
	notech_nand2 i_2420717(.A(n_175075694), .B(n_174575689), .Z(n_24894));
	notech_nand2 i_2320716(.A(n_176075704), .B(n_175575699), .Z(n_24888));
	notech_and4 i_2520782(.A(n_176175705), .B(n_176375707), .C(n_169475638),
		 .D(n_176875712), .Z(n_24574));
	notech_and4 i_2320780(.A(n_176975713), .B(n_177175715), .C(n_168575629),
		 .D(n_177675720), .Z(n_24562));
	notech_or4 i_2420877(.A(n_258069592), .B(n_166975613), .C(n_178075724), 
		.D(n_26686), .Z(n_24220));
	notech_or4 i_2521006(.A(n_257669588), .B(n_166175605), .C(n_178775731), 
		.D(n_26687), .Z(n_23878));
	notech_or4 i_2421005(.A(n_258069592), .B(n_165375597), .C(n_179475738), 
		.D(n_26688), .Z(n_23872));
	notech_or4 i_2321004(.A(n_258469596), .B(n_164575589), .C(n_180175745), 
		.D(n_26689), .Z(n_23866));
	notech_and4 i_2521102(.A(n_180575749), .B(n_180775751), .C(n_164475588),
		 .D(n_181275756), .Z(n_18973));
	notech_and4 i_2421101(.A(n_181375757), .B(n_181575759), .C(n_163575579),
		 .D(n_182075764), .Z(n_18967));
	notech_and4 i_2321100(.A(n_182175765), .B(n_182375767), .C(n_162675570),
		 .D(n_182875772), .Z(n_18961));
	notech_or4 i_2521198(.A(n_257669588), .B(n_161075554), .C(n_183275776), 
		.D(n_26690), .Z(n_18624));
	notech_or4 i_2421197(.A(n_258069592), .B(n_160275546), .C(n_183975783), 
		.D(n_26691), .Z(n_18618));
	notech_or4 i_2321196(.A(n_258469596), .B(n_159475538), .C(n_184675790), 
		.D(n_26692), .Z(n_18612));
	notech_or4 i_2521646(.A(n_257669588), .B(n_158675530), .C(n_185375797), 
		.D(n_26693), .Z(n_17924));
	notech_or4 i_2421645(.A(n_258069592), .B(n_157875522), .C(n_186075804), 
		.D(n_26694), .Z(n_17918));
	notech_or4 i_2421869(.A(n_258069592), .B(n_157075514), .C(n_186775811), 
		.D(n_26695), .Z(n_20756));
	notech_and4 i_2321868(.A(n_187175815), .B(n_187375817), .C(n_188075822),
		 .D(n_156975513), .Z(n_20750));
	notech_nand2 i_197747747(.A(n_57139), .B(n_188775828), .Z(n_57115));
	notech_and4 i_1921000(.A(n_194775886), .B(n_194975888), .C(n_195475893),
		 .D(n_193975878), .Z(n_23842));
	notech_and4 i_1721862(.A(n_195575894), .B(n_195775896), .C(n_196275901),
		 .D(n_193075869), .Z(n_20714));
	notech_nand2 i_1721926(.A(n_197275911), .B(n_196775906), .Z(n_17528));
	notech_nand2 i_1917608(.A(n_198275921), .B(n_197775916), .Z(n_16814));
	notech_nand2 i_1717606(.A(n_199275931), .B(n_198775926), .Z(n_16802));
	notech_and2 i_110147686(.A(n_288869900), .B(n_188675827), .Z(n_311224366
		));
	notech_and2 i_148644553(.A(n_57922), .B(n_201575954), .Z(n_57595));
	notech_and3 i_190161791(.A(n_285563122), .B(n_274863015), .C(n_30803), .Z
		(n_251262779));
	notech_ao4 i_111144561(.A(n_30825), .B(n_60229), .C(n_315191672), .D(n_24994
		), .Z(n_57938));
	notech_and2 i_146244558(.A(n_50904), .B(n_58432), .Z(n_57619));
	notech_and2 i_148544538(.A(n_57923), .B(n_201375952), .Z(n_57596));
	notech_ao3 i_190261790(.A(n_309591728), .B(n_274963016), .C(n_26845), .Z
		(n_251162778));
	notech_ao4 i_3447665(.A(n_30821), .B(n_60234), .C(n_281263079), .D(n_297363240
		), .Z(n_251062777));
	notech_or4 i_3220885(.A(n_215876097), .B(n_213076069), .C(n_217076109), 
		.D(n_26701), .Z(n_24268));
	notech_nand3 i_3221205(.A(n_217576114), .B(n_217476113), .C(n_217976118)
		, .Z(n_18666));
	notech_and4 i_721852(.A(n_212276061), .B(n_218076119), .C(n_218276121), 
		.D(n_218776126), .Z(n_20654));
	notech_nand2 i_621851(.A(n_219776136), .B(n_219276131), .Z(n_20648));
	notech_nand2 i_421849(.A(n_220776146), .B(n_220276141), .Z(n_20636));
	notech_and4 i_721916(.A(n_221476153), .B(n_221376152), .C(n_208576024), 
		.D(n_221876157), .Z(n_17468));
	notech_nand2 i_621915(.A(n_223176170), .B(n_222576164), .Z(n_17462));
	notech_nand2 i_421913(.A(n_224376182), .B(n_223776176), .Z(n_17450));
	notech_nand2 i_717596(.A(n_225476193), .B(n_224976188), .Z(n_16742));
	notech_nand2 i_617595(.A(n_226676205), .B(n_226076199), .Z(n_16736));
	notech_nand2 i_417593(.A(n_227876217), .B(n_227276211), .Z(n_16724));
	notech_and2 i_102144476(.A(n_215576094), .B(n_200875947), .Z(n_306221226
		));
	notech_and2 i_189061793(.A(n_309491729), .B(n_151661799), .Z(n_250962776
		));
	notech_nand2 i_73746986(.A(opa[16]), .B(n_26833), .Z(n_250862775));
	notech_and2 i_7847621(.A(n_312324377), .B(n_250862775), .Z(n_250762774)
		);
	notech_and4 i_3147668(.A(n_56848), .B(n_125961542), .C(n_26804), .D(n_58477
		), .Z(n_250662773));
	notech_and4 i_259147687(.A(n_56848), .B(n_187762157), .C(n_58486), .D(n_58478
		), .Z(n_250562772));
	notech_and4 i_156249143(.A(n_240962676), .B(n_250162768), .C(n_241262679
		), .D(n_26672), .Z(n_250462771));
	notech_nand3 i_3217781(.A(n_298276921), .B(n_297876917), .C(n_297376912)
		, .Z(n_22401));
	notech_nand3 i_3117780(.A(n_300276941), .B(n_299876937), .C(n_299376932)
		, .Z(n_22395));
	notech_nand3 i_3017779(.A(n_302276961), .B(n_301876957), .C(n_301376952)
		, .Z(n_22389));
	notech_nand3 i_2917778(.A(n_304276981), .B(n_303876977), .C(n_303376972)
		, .Z(n_22383));
	notech_nand3 i_2817777(.A(n_306277001), .B(n_305876997), .C(n_305376992)
		, .Z(n_22377));
	notech_nand3 i_2717776(.A(n_308277021), .B(n_307877017), .C(n_307377012)
		, .Z(n_22371));
	notech_nand3 i_2617775(.A(n_310277041), .B(n_309877037), .C(n_309377032)
		, .Z(n_22365));
	notech_nand3 i_2517774(.A(n_312277061), .B(n_311877057), .C(n_311377052)
		, .Z(n_22359));
	notech_nand3 i_2417773(.A(n_314277081), .B(n_313877077), .C(n_313377072)
		, .Z(n_22353));
	notech_nand3 i_2317772(.A(n_316277101), .B(n_315877097), .C(n_315377092)
		, .Z(n_22347));
	notech_nand3 i_2217771(.A(n_318277121), .B(n_317877117), .C(n_317377112)
		, .Z(n_22341));
	notech_nand3 i_2117770(.A(n_320277141), .B(n_319877137), .C(n_319377132)
		, .Z(n_22335));
	notech_nand3 i_2017769(.A(n_322277161), .B(n_321877157), .C(n_321377152)
		, .Z(n_22329));
	notech_nand3 i_1917768(.A(n_324277181), .B(n_323877177), .C(n_323377172)
		, .Z(n_22323));
	notech_nand3 i_1817767(.A(n_326277201), .B(n_325877197), .C(n_325377192)
		, .Z(n_22317));
	notech_nand3 i_1717766(.A(n_328277221), .B(n_327877217), .C(n_327377212)
		, .Z(n_22311));
	notech_and4 i_1617765(.A(n_331377252), .B(n_330777246), .C(n_329977238),
		 .D(n_329377232), .Z(n_22305));
	notech_and4 i_1517764(.A(n_334177280), .B(n_333577274), .C(n_332777266),
		 .D(n_332177260), .Z(n_22299));
	notech_and4 i_1417763(.A(n_336977308), .B(n_336377302), .C(n_335577294),
		 .D(n_334977288), .Z(n_22293));
	notech_and4 i_1317762(.A(n_339777336), .B(n_339177330), .C(n_338377322),
		 .D(n_337777316), .Z(n_22287));
	notech_and4 i_1217761(.A(n_342577364), .B(n_341977358), .C(n_341177350),
		 .D(n_340577344), .Z(n_22281));
	notech_and4 i_1117760(.A(n_345377392), .B(n_344777386), .C(n_343977378),
		 .D(n_343377372), .Z(n_22275));
	notech_and4 i_1017759(.A(n_348177420), .B(n_347577414), .C(n_346777406),
		 .D(n_346177400), .Z(n_22269));
	notech_and4 i_917758(.A(n_350977448), .B(n_350377442), .C(n_349577434), 
		.D(n_348977428), .Z(n_22263));
	notech_and4 i_217751(.A(n_353677475), .B(n_353077469), .C(n_352377462), 
		.D(n_351777456), .Z(n_22221));
	notech_and4 i_117750(.A(n_356377502), .B(n_355777496), .C(n_355077489), 
		.D(n_354477483), .Z(n_22215));
	notech_or4 i_40035099(.A(n_27907), .B(n_62808), .C(n_60910), .D(n_60234)
		, .Z(n_308547770));
	notech_xor2 i_113835093(.A(\nbus_11307[0] ), .B(opa[1]), .Z(n_307947775)
		);
	notech_ao4 i_156049145(.A(n_55992), .B(n_275463021), .C(n_59259), .D(n_135961642
		), .Z(n_250162768));
	notech_and4 i_156849138(.A(n_241562682), .B(n_249862765), .C(n_249662763
		), .D(n_241862685), .Z(n_250062767));
	notech_ao4 i_156349142(.A(n_275363020), .B(n_58316), .C(n_152472004), .D
		(n_136261645), .Z(n_249862765));
	notech_ao4 i_156549140(.A(n_285463121), .B(n_239862665), .C(n_136161644)
		, .D(n_239762664), .Z(n_249662763));
	notech_mux2 i_156949137(.S(n_32319), .A(n_312147737), .B(n_344466973), .Z
		(n_249562762));
	notech_ao4 i_157049136(.A(n_28111), .B(n_60347), .C(n_250962776), .D(n_57742
		), .Z(n_249362760));
	notech_ao4 i_157149135(.A(n_251362780), .B(n_56338), .C(n_60003), .D(n_251262779
		), .Z(n_249262759));
	notech_and3 i_157649130(.A(n_248862755), .B(n_249062757), .C(n_242862695
		), .Z(n_249162758));
	notech_ao4 i_157349133(.A(n_251162778), .B(n_29708), .C(n_58426), .D(n_28007
		), .Z(n_249062757));
	notech_ao4 i_157449132(.A(n_225765786), .B(n_316537960), .C(n_224065769)
		, .D(n_309721261), .Z(n_248862755));
	notech_ao4 i_157749129(.A(n_28112), .B(n_60347), .C(n_250962776), .D(n_57751
		), .Z(n_248662753));
	notech_ao4 i_157849128(.A(n_251362780), .B(n_56347), .C(n_60002), .D(n_251262779
		), .Z(n_248562752));
	notech_and3 i_158349123(.A(n_248162748), .B(n_248362750), .C(n_243662703
		), .Z(n_248462751));
	notech_ao4 i_158049126(.A(n_251162778), .B(n_29765), .C(n_28008), .D(n_58426
		), .Z(n_248362750));
	notech_ao4 i_158149125(.A(n_225665785), .B(n_316537960), .C(n_222565754)
		, .D(n_309721261), .Z(n_248162748));
	notech_ao4 i_158449122(.A(n_28113), .B(n_60347), .C(n_250962776), .D(n_57761
		), .Z(n_247962746));
	notech_ao4 i_158549121(.A(n_251362780), .B(n_56475), .C(n_60001), .D(n_251262779
		), .Z(n_247862745));
	notech_and3 i_159049116(.A(n_247462741), .B(n_247662743), .C(n_244462711
		), .Z(n_247762744));
	notech_ao4 i_158749119(.A(n_251162778), .B(n_29769), .C(n_58426), .D(n_28009
		), .Z(n_247662743));
	notech_ao4 i_158849118(.A(n_225565784), .B(n_316537960), .C(n_221065739)
		, .D(n_309721261), .Z(n_247462741));
	notech_ao4 i_159149115(.A(n_28114), .B(n_60347), .C(n_250962776), .D(n_57771
		), .Z(n_247262739));
	notech_ao4 i_159249114(.A(n_251362780), .B(n_55965), .C(n_60000), .D(n_251262779
		), .Z(n_247162738));
	notech_and3 i_159749109(.A(n_246762734), .B(n_246962736), .C(n_245262719
		), .Z(n_247062737));
	notech_ao4 i_159449112(.A(n_251162778), .B(n_29770), .C(n_58426), .D(n_28010
		), .Z(n_246962736));
	notech_ao4 i_159549111(.A(n_316537960), .B(n_256069572), .C(n_253569547)
		, .D(n_309721261), .Z(n_246762734));
	notech_nao3 i_192348793(.A(n_57514), .B(n_27112), .C(fsmf[2]), .Z(n_246562732
		));
	notech_or4 i_192648790(.A(fsmf[3]), .B(fsmf[0]), .C(fsmf[1]), .D(instrc[
		6]), .Z(n_246362730));
	notech_or4 i_193048786(.A(instrc[4]), .B(instrc[7]), .C(instrc[5]), .D(instrc
		[3]), .Z(n_245962726));
	notech_or4 i_193348783(.A(instrc[2]), .B(instrc[1]), .C(n_29771), .D(n_29117
		), .Z(n_245662723));
	notech_nand2 i_29122(.A(n_57026), .B(instrc[119]), .Z(n_245362720));
	notech_or2 i_70649979(.A(n_288927271), .B(n_322438019), .Z(n_245262719)
		);
	notech_or2 i_69649987(.A(n_289027272), .B(n_322438019), .Z(n_244462711)
		);
	notech_or2 i_68849995(.A(n_289127273), .B(n_322438019), .Z(n_243662703)
		);
	notech_or2 i_67650003(.A(n_289227274), .B(n_322438019), .Z(n_242862695)
		);
	notech_or4 i_66250017(.A(n_62864), .B(n_136361646), .C(n_60947), .D(n_57552
		), .Z(n_241862685));
	notech_or4 i_66550014(.A(n_56824), .B(n_26610), .C(n_59991), .D(n_56632)
		, .Z(n_241562682));
	notech_nao3 i_66850011(.A(n_126061543), .B(opa[2]), .C(n_140661689), .Z(n_241262679
		));
	notech_or4 i_66950010(.A(n_285463121), .B(n_28126), .C(n_60947), .D(n_174962032
		), .Z(n_240962676));
	notech_ao3 i_104549648(.A(n_32386), .B(n_56662), .C(n_56824), .Z(n_240762674
		));
	notech_nao3 i_104149652(.A(n_56471), .B(n_32332), .C(n_58100), .Z(n_240362670
		));
	notech_and3 i_103349660(.A(n_58503), .B(n_26816), .C(n_58479), .Z(n_240162668
		));
	notech_and2 i_3950627(.A(n_249562762), .B(n_58714), .Z(n_239862665));
	notech_mux2 i_3850628(.S(n_32319), .A(n_285027232), .B(n_284927231), .Z(n_239762664
		));
	notech_and4 i_190852070(.A(n_239462661), .B(n_239362660), .C(n_239162658
		), .D(n_239062657), .Z(n_239662663));
	notech_ao4 i_190252076(.A(n_58789), .B(n_28620), .C(n_58791), .D(n_29373
		), .Z(n_239462661));
	notech_ao4 i_190152077(.A(n_59152), .B(n_29311), .C(n_27065), .D(n_29342
		), .Z(n_239362660));
	notech_ao4 i_190052078(.A(n_1887), .B(n_29764), .C(n_330563522), .D(n_27830
		), .Z(n_239162658));
	notech_ao4 i_189952079(.A(n_310247754), .B(n_29763), .C(n_310447752), .D
		(n_29762), .Z(n_239062657));
	notech_ao4 i_190452074(.A(n_58788), .B(n_28414), .C(n_58750), .D(n_28012
		), .Z(n_238862655));
	notech_ao4 i_190352075(.A(n_58751), .B(\nbus_11358[27] ), .C(n_310347753
		), .D(nbus_11295[27]), .Z(n_238762654));
	notech_ao4 i_166452312(.A(n_311491709), .B(n_170292129), .C(n_311391710)
		, .D(n_174392093), .Z(n_238562652));
	notech_and4 i_166252314(.A(n_238162648), .B(n_238062647), .C(n_237862645
		), .D(n_215762424), .Z(n_238362650));
	notech_ao4 i_165952317(.A(n_26696), .B(n_29659), .C(n_151428791), .D(n_128228559
		), .Z(n_238162648));
	notech_ao4 i_165852318(.A(n_311191712), .B(\nbus_11358[29] ), .C(n_311091713
		), .D(\nbus_11365[29] ), .Z(n_238062647));
	notech_ao4 i_165752319(.A(n_59124), .B(nbus_11295[29]), .C(n_54638), .D(n_28960
		), .Z(n_237862645));
	notech_and4 i_153952437(.A(n_237262639), .B(n_237062637), .C(n_236962636
		), .D(n_237462641), .Z(n_237662643));
	notech_and3 i_153652440(.A(n_54667), .B(n_57029), .C(n_214862415), .Z(n_237462641
		));
	notech_ao4 i_153552441(.A(n_149228769), .B(n_29661), .C(n_149128768), .D
		(n_131228589), .Z(n_237262639));
	notech_ao4 i_153452442(.A(n_149428771), .B(\nbus_11358[27] ), .C(n_149328770
		), .D(\nbus_11365[27] ), .Z(n_237062637));
	notech_ao4 i_153352443(.A(n_310791716), .B(n_310091723), .C(n_54643), .D
		(n_28982), .Z(n_236962636));
	notech_ao4 i_148452492(.A(n_3858), .B(n_174292094), .C(n_3843), .D(n_174992087
		), .Z(n_236762634));
	notech_and4 i_148252494(.A(n_54667), .B(n_236362630), .C(n_236162628), .D
		(n_213462401), .Z(n_236562632));
	notech_ao4 i_147952497(.A(n_148228759), .B(n_133728614), .C(n_3877), .D(\nbus_11358[26] 
		), .Z(n_236362630));
	notech_ao4 i_148052496(.A(n_3857), .B(n_28011), .C(n_26642), .D(n_29660)
		, .Z(n_236162628));
	notech_ao4 i_142952542(.A(n_170292129), .B(n_3858), .C(n_174392093), .D(n_3843
		), .Z(n_235962626));
	notech_and4 i_142752544(.A(n_54667), .B(n_235562622), .C(n_235362620), .D
		(n_212662393), .Z(n_235762624));
	notech_ao4 i_142452547(.A(n_128228559), .B(n_148228759), .C(n_3877), .D(\nbus_11358[29] 
		), .Z(n_235562622));
	notech_ao4 i_142552546(.A(n_28014), .B(n_3857), .C(n_29659), .D(n_26642)
		, .Z(n_235362620));
	notech_and3 i_138652584(.A(n_234362610), .B(n_234262609), .C(n_235062617
		), .Z(n_235162618));
	notech_and4 i_138552585(.A(n_234862615), .B(n_234762614), .C(n_234562612
		), .D(n_212362390), .Z(n_235062617));
	notech_ao4 i_137952591(.A(n_147028747), .B(\nbus_11358[27] ), .C(n_146928746
		), .D(\nbus_11365[27] ), .Z(n_234862615));
	notech_ao4 i_137852592(.A(n_301791806), .B(n_310091723), .C(n_146228739)
		, .D(n_29761), .Z(n_234762614));
	notech_ao4 i_137752593(.A(n_54883), .B(n_28620), .C(n_54894), .D(n_27479
		), .Z(n_234562612));
	notech_ao4 i_138152589(.A(n_310391720), .B(n_28012), .C(n_310291721), .D
		(n_28116), .Z(n_234362610));
	notech_ao4 i_138052590(.A(n_147128748), .B(n_29661), .C(n_131228589), .D
		(n_147228749), .Z(n_234262609));
	notech_ao4 i_126152707(.A(n_170292129), .B(n_58084), .C(n_174392093), .D
		(n_151931934), .Z(n_234062607));
	notech_and4 i_126052708(.A(n_210962376), .B(n_233662603), .C(n_233562602
		), .D(n_220562472), .Z(n_233962606));
	notech_ao4 i_125652712(.A(n_57875), .B(\nbus_11358[29] ), .C(\nbus_11365[29] 
		), .D(n_57868), .Z(n_233662603));
	notech_ao4 i_125752711(.A(n_26929), .B(n_29659), .C(n_58147), .D(n_128228559
		), .Z(n_233562602));
	notech_nand3 i_110752860(.A(n_233062597), .B(n_232962596), .C(n_232862595
		), .Z(n_233262599));
	notech_ao4 i_110452863(.A(n_142928706), .B(n_29660), .C(n_133728614), .D
		(n_143028707), .Z(n_233062597));
	notech_ao4 i_110352864(.A(n_142828705), .B(\nbus_11358[26] ), .C(n_142728704
		), .D(\nbus_11365[26] ), .Z(n_232962596));
	notech_ao4 i_110552862(.A(n_4014), .B(n_28011), .C(n_55726), .D(n_28115)
		, .Z(n_232862595));
	notech_and4 i_109052876(.A(n_232462591), .B(n_232362590), .C(n_209362360
		), .D(n_232162588), .Z(n_232662593));
	notech_ao4 i_108752879(.A(n_55726), .B(n_28116), .C(n_142928706), .D(n_29661
		), .Z(n_232462591));
	notech_ao4 i_108652880(.A(n_131228589), .B(n_143028707), .C(n_142828705)
		, .D(n_55938), .Z(n_232362590));
	notech_ao4 i_108552881(.A(n_142728704), .B(\nbus_11365[27] ), .C(n_310091723
		), .D(n_295269964), .Z(n_232162588));
	notech_nand3 i_107252894(.A(n_231662583), .B(n_231562582), .C(n_231462581
		), .Z(n_231862585));
	notech_ao4 i_106952897(.A(n_142928706), .B(n_29662), .C(n_143028707), .D
		(n_130528582), .Z(n_231662583));
	notech_ao4 i_106852898(.A(n_142828705), .B(\nbus_11358[28] ), .C(n_142728704
		), .D(\nbus_11365[28] ), .Z(n_231562582));
	notech_ao4 i_107052896(.A(n_4014), .B(n_28013), .C(n_55726), .D(n_28117)
		, .Z(n_231462581));
	notech_nand3 i_89553067(.A(n_230962576), .B(n_230862575), .C(n_230762574
		), .Z(n_231162578));
	notech_ao4 i_88853073(.A(n_140128678), .B(\nbus_11365[27] ), .C(n_310091723
		), .D(n_309691727), .Z(n_230962576));
	notech_ao4 i_88753074(.A(n_54649), .B(n_29760), .C(n_28527), .D(n_29759)
		, .Z(n_230862575));
	notech_ao4 i_89153070(.A(n_60122), .B(n_27243), .C(n_303591788), .D(n_28012
		), .Z(n_230762574));
	notech_nand2 i_89453068(.A(n_230562572), .B(n_230462571), .Z(n_230662573
		));
	notech_ao4 i_89053071(.A(n_32270), .B(n_28116), .C(n_140328680), .D(n_29661
		), .Z(n_230562572));
	notech_ao4 i_88953072(.A(n_131228589), .B(n_140428681), .C(n_140228679),
		 .D(n_55938), .Z(n_230462571));
	notech_ao4 i_77353183(.A(n_170292129), .B(n_58082), .C(n_174392093), .D(n_319937994
		), .Z(n_230262569));
	notech_and4 i_77253184(.A(n_229862565), .B(n_229762564), .C(n_220562472)
		, .D(n_206262329), .Z(n_230162568));
	notech_ao4 i_76853188(.A(n_57873), .B(\nbus_11358[29] ), .C(n_57869), .D
		(\nbus_11365[29] ), .Z(n_229862565));
	notech_ao4 i_76953187(.A(n_26918), .B(n_29659), .C(n_58145), .D(n_128228559
		), .Z(n_229762564));
	notech_ao4 i_75753199(.A(n_174292094), .B(n_58085), .C(n_174992087), .D(n_306124325
		), .Z(n_229562562));
	notech_and4 i_75653200(.A(n_229162558), .B(n_229062557), .C(n_228962556)
		, .D(n_174892088), .Z(n_229462561));
	notech_ao4 i_75253204(.A(n_58143), .B(n_133728614), .C(n_57877), .D(\nbus_11358[26] 
		), .Z(n_229162558));
	notech_ao4 i_75153205(.A(n_57870), .B(\nbus_11365[26] ), .C(n_154331958)
		, .D(nbus_11295[26]), .Z(n_229062557));
	notech_ao4 i_75353203(.A(n_58427), .B(n_28011), .C(n_26902), .D(n_29660)
		, .Z(n_228962556));
	notech_ao4 i_72153235(.A(n_172792106), .B(n_58085), .C(n_174492092), .D(n_306124325
		), .Z(n_228762554));
	notech_and4 i_72053236(.A(n_228362550), .B(n_228262549), .C(n_228162548)
		, .D(n_242259503), .Z(n_228662553));
	notech_ao4 i_71653240(.A(n_58143), .B(n_130528582), .C(n_57877), .D(\nbus_11358[28] 
		), .Z(n_228362550));
	notech_ao4 i_71553241(.A(n_57870), .B(\nbus_11365[28] ), .C(n_154331958)
		, .D(nbus_11295[28]), .Z(n_228262549));
	notech_ao4 i_71753239(.A(n_58427), .B(n_28013), .C(n_26902), .D(n_29662)
		, .Z(n_228162548));
	notech_ao4 i_70353253(.A(n_170292129), .B(n_58085), .C(n_174392093), .D(n_306124325
		), .Z(n_227962546));
	notech_and4 i_70253254(.A(n_227562542), .B(n_227462541), .C(n_227362540)
		, .D(n_220562472), .Z(n_227862545));
	notech_ao4 i_69853258(.A(n_58143), .B(n_128228559), .C(n_57877), .D(\nbus_11358[29] 
		), .Z(n_227562542));
	notech_ao4 i_69753259(.A(n_57870), .B(\nbus_11365[29] ), .C(n_56356), .D
		(nbus_11295[29]), .Z(n_227462541));
	notech_ao4 i_69953257(.A(n_58427), .B(n_28014), .C(n_26902), .D(n_29659)
		, .Z(n_227362540));
	notech_and4 i_66653287(.A(n_226962536), .B(n_226862535), .C(n_202862295)
		, .D(n_226662533), .Z(n_227162538));
	notech_ao4 i_66353290(.A(n_251162778), .B(n_29661), .C(n_251262779), .D(n_131228589
		), .Z(n_226962536));
	notech_ao4 i_66253291(.A(n_251362780), .B(n_55938), .C(n_250962776), .D(n_57792
		), .Z(n_226862535));
	notech_ao4 i_66153292(.A(n_60347), .B(n_28116), .C(n_316537960), .D(n_310091723
		), .Z(n_226662533));
	notech_and4 i_63253320(.A(n_201962286), .B(n_226062527), .C(n_225962526)
		, .D(n_3883), .Z(n_226362530));
	notech_ao4 i_62853324(.A(n_251362780), .B(\nbus_11358[29] ), .C(n_250962776
		), .D(\nbus_11365[29] ), .Z(n_226062527));
	notech_ao4 i_62953323(.A(n_251162778), .B(n_29659), .C(n_251262779), .D(n_128228559
		), .Z(n_225962526));
	notech_ao4 i_61753335(.A(n_174292094), .B(n_307124335), .C(n_174992087),
		 .D(n_306624330), .Z(n_225762524));
	notech_and4 i_61653336(.A(n_201162278), .B(n_225362520), .C(n_225262519)
		, .D(n_174892088), .Z(n_225662523));
	notech_ao4 i_61253340(.A(n_57864), .B(\nbus_11358[26] ), .C(n_314047718)
		, .D(\nbus_11365[26] ), .Z(n_225362520));
	notech_ao4 i_61353339(.A(n_307324337), .B(n_29660), .C(n_58141), .D(n_133728614
		), .Z(n_225262519));
	notech_ao4 i_56853383(.A(n_170292129), .B(n_307124335), .C(n_174392093),
		 .D(n_306624330), .Z(n_225062517));
	notech_and4 i_56753384(.A(n_200362270), .B(n_224662513), .C(n_224562512)
		, .D(n_220562472), .Z(n_224962516));
	notech_ao4 i_56353388(.A(n_57864), .B(\nbus_11358[29] ), .C(n_314047718)
		, .D(\nbus_11365[29] ), .Z(n_224662513));
	notech_ao4 i_56453387(.A(n_307324337), .B(n_29659), .C(n_58141), .D(n_128228559
		), .Z(n_224562512));
	notech_ao4 i_50453447(.A(n_170292129), .B(n_286927251), .C(n_174392093),
		 .D(n_286827250), .Z(n_224362510));
	notech_and4 i_50353448(.A(n_223962506), .B(n_223862505), .C(n_220562472)
		, .D(n_199562262), .Z(n_224262509));
	notech_ao4 i_49953452(.A(n_57863), .B(\nbus_11358[29] ), .C(n_57861), .D
		(\nbus_11365[29] ), .Z(n_223962506));
	notech_ao4 i_50053451(.A(n_26615), .B(n_29659), .C(n_58139), .D(n_128228559
		), .Z(n_223862505));
	notech_ao4 i_48853463(.A(n_174292094), .B(n_58008), .C(n_174992087), .D(n_58007
		), .Z(n_223662503));
	notech_and4 i_48753464(.A(n_223262499), .B(n_223162498), .C(n_223062497)
		, .D(n_174892088), .Z(n_223562502));
	notech_ao4 i_48353468(.A(n_57726), .B(n_28152), .C(n_58138), .D(n_133728614
		), .Z(n_223262499));
	notech_ao4 i_48253469(.A(n_57865), .B(\nbus_11358[26] ), .C(n_57867), .D
		(\nbus_11365[26] ), .Z(n_223162498));
	notech_ao4 i_48453467(.A(n_58423), .B(n_28011), .C(n_26937), .D(n_29660)
		, .Z(n_223062497));
	notech_and4 i_46253488(.A(n_222662493), .B(n_222562492), .C(n_222362490)
		, .D(n_222262489), .Z(n_222862495));
	notech_ao4 i_45953491(.A(n_58423), .B(n_28012), .C(n_26937), .D(n_29661)
		, .Z(n_222662493));
	notech_ao4 i_45853492(.A(n_57726), .B(n_28153), .C(n_58138), .D(n_131228589
		), .Z(n_222562492));
	notech_ao4 i_45753493(.A(n_57865), .B(n_55938), .C(n_57867), .D(n_57792)
		, .Z(n_222362490));
	notech_nor2 i_45653494(.A(n_1978), .B(n_196962240), .Z(n_222262489));
	notech_ao4 i_44453506(.A(n_172792106), .B(n_58008), .C(n_174492092), .D(n_58007
		), .Z(n_222062487));
	notech_and4 i_44353507(.A(n_221662483), .B(n_221562482), .C(n_221462481)
		, .D(n_242259503), .Z(n_221962486));
	notech_ao4 i_43953511(.A(n_57726), .B(n_28154), .C(n_58138), .D(n_130528582
		), .Z(n_221662483));
	notech_ao4 i_43853512(.A(n_57865), .B(\nbus_11358[28] ), .C(n_57867), .D
		(\nbus_11365[28] ), .Z(n_221562482));
	notech_ao4 i_44053510(.A(n_58423), .B(n_28013), .C(n_26937), .D(n_29662)
		, .Z(n_221462481));
	notech_ao4 i_41753531(.A(n_170292129), .B(n_58008), .C(n_174392093), .D(n_58007
		), .Z(n_221262479));
	notech_and4 i_41653532(.A(n_220862475), .B(n_220762474), .C(n_220662473)
		, .D(n_220562472), .Z(n_221162478));
	notech_ao4 i_41253536(.A(n_57726), .B(n_28155), .C(n_58138), .D(n_128228559
		), .Z(n_220862475));
	notech_ao4 i_41153537(.A(n_57865), .B(\nbus_11358[29] ), .C(n_57867), .D
		(\nbus_11365[29] ), .Z(n_220762474));
	notech_ao4 i_41353535(.A(n_28014), .B(n_58423), .C(n_26937), .D(n_29659)
		, .Z(n_220662473));
	notech_and3 i_68553916(.A(n_220362470), .B(n_220262469), .C(n_3883), .Z(n_220562472
		));
	notech_ao4 i_39953548(.A(n_309591728), .B(n_29659), .C(n_30803), .D(n_128228559
		), .Z(n_220362470));
	notech_ao4 i_39853549(.A(n_304691777), .B(\nbus_11358[29] ), .C(n_309491729
		), .D(\nbus_11365[29] ), .Z(n_220262469));
	notech_nand3 i_38953557(.A(n_219362460), .B(n_219262459), .C(n_219862465
		), .Z(n_219962466));
	notech_and3 i_38853558(.A(n_219662463), .B(n_219562462), .C(n_194262214)
		, .Z(n_219862465));
	notech_ao4 i_38253564(.A(n_309091733), .B(\nbus_11358[26] ), .C(n_308991734
		), .D(\nbus_11365[26] ), .Z(n_219662463));
	notech_ao4 i_38553561(.A(n_121628493), .B(n_28011), .C(n_309291731), .D(n_28115
		), .Z(n_219562462));
	notech_ao4 i_38453562(.A(n_56091), .B(n_29758), .C(n_26765), .D(n_29660)
		, .Z(n_219362460));
	notech_ao4 i_38353563(.A(n_122428501), .B(n_28152), .C(n_122528502), .D(n_133728614
		), .Z(n_219262459));
	notech_nand3 i_33653610(.A(n_218362450), .B(n_218262449), .C(n_218862455
		), .Z(n_218962456));
	notech_and3 i_33553611(.A(n_218662453), .B(n_218562452), .C(n_193062202)
		, .Z(n_218862455));
	notech_ao4 i_32953617(.A(n_309091733), .B(n_55938), .C(n_308991734), .D(n_57792
		), .Z(n_218662453));
	notech_ao4 i_33253614(.A(n_121628493), .B(n_28012), .C(n_309291731), .D(n_28116
		), .Z(n_218562452));
	notech_ao4 i_33153615(.A(n_56091), .B(n_29757), .C(n_26765), .D(n_29661)
		, .Z(n_218362450));
	notech_ao4 i_33053616(.A(n_122428501), .B(n_28153), .C(n_122528502), .D(n_131228589
		), .Z(n_218262449));
	notech_nand3 i_31353633(.A(n_217362440), .B(n_217262439), .C(n_217862445
		), .Z(n_217962446));
	notech_and3 i_31253634(.A(n_217662443), .B(n_217562442), .C(n_191862190)
		, .Z(n_217862445));
	notech_ao4 i_30653640(.A(n_309091733), .B(\nbus_11358[28] ), .C(n_308991734
		), .D(\nbus_11365[28] ), .Z(n_217662443));
	notech_ao4 i_30953637(.A(n_121628493), .B(n_28013), .C(n_309291731), .D(n_28117
		), .Z(n_217562442));
	notech_ao4 i_30853638(.A(n_309191732), .B(n_29756), .C(n_26765), .D(n_29662
		), .Z(n_217362440));
	notech_ao4 i_30753639(.A(n_122428501), .B(n_28154), .C(n_122528502), .D(n_130528582
		), .Z(n_217262439));
	notech_nand3 i_2818993(.A(n_238862655), .B(n_238762654), .C(n_239662663)
		, .Z(n_25650));
	notech_and4 i_3017619(.A(n_238362650), .B(n_238562652), .C(n_220562472),
		 .D(n_215062417), .Z(n_16880));
	notech_or2 i_165352323(.A(n_311291711), .B(n_28014), .Z(n_215762424));
	notech_or2 i_165452322(.A(n_151128788), .B(n_3981), .Z(n_215062417));
	notech_nand3 i_2821937(.A(n_214962416), .B(n_237662643), .C(n_214162408)
		, .Z(n_17594));
	notech_or4 i_153152445(.A(n_311991704), .B(n_26939), .C(nbus_11295[27]),
		 .D(n_60947), .Z(n_214962416));
	notech_or4 i_152952447(.A(n_56824), .B(n_56946), .C(n_56527), .D(n_28012
		), .Z(n_214862415));
	notech_or2 i_153052446(.A(n_148728764), .B(n_4016), .Z(n_214162408));
	notech_and4 i_2721872(.A(n_236562632), .B(n_236762634), .C(n_174892088),
		 .D(n_213362400), .Z(n_20774));
	notech_or2 i_147052506(.A(n_3878), .B(\nbus_11365[26] ), .Z(n_213462401)
		);
	notech_or2 i_147552501(.A(n_3837), .B(n_3983), .Z(n_213362400));
	notech_and4 i_3021875(.A(n_220562472), .B(n_235762624), .C(n_235962626),
		 .D(n_212562392), .Z(n_20792));
	notech_or2 i_141552556(.A(n_3878), .B(\nbus_11365[29] ), .Z(n_212662393)
		);
	notech_or2 i_142052551(.A(n_3981), .B(n_3837), .Z(n_212562392));
	notech_nand3 i_2821809(.A(n_212462391), .B(n_235162618), .C(n_211262379)
		, .Z(n_21146));
	notech_or4 i_137652594(.A(n_312191702), .B(nbus_11295[27]), .C(n_60947),
		 .D(n_54930), .Z(n_212462391));
	notech_nand2 i_137452596(.A(sav_esp[27]), .B(n_61143), .Z(n_212362390)
		);
	notech_or2 i_137552595(.A(n_4016), .B(n_146428741), .Z(n_211262379));
	notech_nand3 i_3021651(.A(n_234062607), .B(n_233962606), .C(n_210462371)
		, .Z(n_17954));
	notech_or4 i_125252716(.A(n_59275), .B(n_2479), .C(n_56688), .D(n_28014)
		, .Z(n_210962376));
	notech_or2 i_125352715(.A(n_3981), .B(n_154831963), .Z(n_210462371));
	notech_or4 i_2721392(.A(n_210262369), .B(n_233262599), .C(n_210362370), 
		.D(n_209562362), .Z(n_25402));
	notech_and3 i_110252865(.A(opc[26]), .B(n_62808), .C(n_4010), .Z(n_210362370
		));
	notech_ao3 i_110152866(.A(opc_10[26]), .B(n_62808), .C(n_295269964), .Z(n_210262369
		));
	notech_nor2 i_110052867(.A(n_3983), .B(n_309891725), .Z(n_209562362));
	notech_nand3 i_2821393(.A(n_232662593), .B(n_209462361), .C(n_208662353)
		, .Z(n_25408));
	notech_or4 i_108452882(.A(n_304991774), .B(n_57881), .C(n_60945), .D(n_26601
		), .Z(n_209462361));
	notech_or4 i_108252884(.A(n_56824), .B(n_56944), .C(n_56513), .D(n_28012
		), .Z(n_209362360));
	notech_or2 i_108352883(.A(n_4016), .B(n_309891725), .Z(n_208662353));
	notech_or4 i_2921394(.A(n_208462351), .B(n_231862585), .C(n_208562352), 
		.D(n_207762344), .Z(n_25414));
	notech_and3 i_106752899(.A(opc[28]), .B(n_62808), .C(n_4010), .Z(n_208562352
		));
	notech_ao3 i_106652900(.A(opc_10[28]), .B(n_62808), .C(n_295269964), .Z(n_208462351
		));
	notech_nor2 i_106552901(.A(n_309891725), .B(n_3982), .Z(n_207762344));
	notech_or4 i_2821361(.A(n_231162578), .B(n_230662573), .C(n_207662343), 
		.D(n_206562332), .Z(n_21498));
	notech_and3 i_88653075(.A(opc[27]), .B(n_62808), .C(n_309791726), .Z(n_207662343
		));
	notech_nor2 i_88553076(.A(n_4016), .B(n_139728674), .Z(n_206562332));
	notech_nand3 i_3021203(.A(n_230262569), .B(n_230162568), .C(n_205762324)
		, .Z(n_18654));
	notech_or2 i_76453192(.A(n_321438009), .B(n_28014), .Z(n_206262329));
	notech_or2 i_76553191(.A(n_3981), .B(n_321538010), .Z(n_205762324));
	notech_nand3 i_2721104(.A(n_229562562), .B(n_229462561), .C(n_204862315)
		, .Z(n_18985));
	notech_or2 i_74853208(.A(n_3983), .B(n_305924323), .Z(n_204862315));
	notech_nand3 i_2921106(.A(n_228762554), .B(n_228662553), .C(n_203962306)
		, .Z(n_18997));
	notech_or2 i_71253244(.A(n_3982), .B(n_305924323), .Z(n_203962306));
	notech_nand3 i_3021107(.A(n_227962546), .B(n_227862545), .C(n_203062297)
		, .Z(n_19003));
	notech_or2 i_69453262(.A(n_3981), .B(n_305924323), .Z(n_203062297));
	notech_nand3 i_2821041(.A(n_227162538), .B(n_202962296), .C(n_202262289)
		, .Z(n_14136));
	notech_or4 i_66053293(.A(n_281263079), .B(n_174962032), .C(n_57881), .D(n_60945
		), .Z(n_202962296));
	notech_or4 i_65853295(.A(n_56824), .B(n_56944), .C(n_56632), .D(n_28012)
		, .Z(n_202862295));
	notech_or2 i_65953294(.A(n_322438019), .B(n_4016), .Z(n_202262289));
	notech_or4 i_3021043(.A(n_202062287), .B(n_202162288), .C(n_201462281), 
		.D(n_26911), .Z(n_14148));
	notech_and3 i_62753325(.A(opc[29]), .B(n_62780), .C(n_26762), .Z(n_202162288
		));
	notech_ao3 i_62653326(.A(opc_10[29]), .B(n_62808), .C(n_316537960), .Z(n_202062287
		));
	notech_or4 i_62453328(.A(n_56824), .B(n_56625), .C(n_56944), .D(n_28014)
		, .Z(n_201962286));
	notech_nor2 i_62553327(.A(n_322438019), .B(n_3981), .Z(n_201462281));
	notech_nand3 i_2721008(.A(n_225762524), .B(n_225662523), .C(n_200662273)
		, .Z(n_23890));
	notech_or4 i_60853344(.A(n_56827), .B(n_56944), .C(n_56649), .D(n_28011)
		, .Z(n_201162278));
	notech_or2 i_60953343(.A(n_3983), .B(n_306824332), .Z(n_200662273));
	notech_nand3 i_3021011(.A(n_225062517), .B(n_224962516), .C(n_199862265)
		, .Z(n_23908));
	notech_or4 i_55953392(.A(n_56827), .B(n_56944), .C(n_56649), .D(n_28014)
		, .Z(n_200362270));
	notech_or2 i_56053391(.A(n_3981), .B(n_306824332), .Z(n_199862265));
	notech_nand3 i_3020883(.A(n_224362510), .B(n_224262509), .C(n_199062257)
		, .Z(n_24256));
	notech_or4 i_49553456(.A(n_56824), .B(n_56946), .C(n_56662), .D(n_28014)
		, .Z(n_199562262));
	notech_or2 i_49653455(.A(n_3981), .B(n_287827260), .Z(n_199062257));
	notech_nand3 i_2720784(.A(n_223662503), .B(n_223562502), .C(n_197762248)
		, .Z(n_24586));
	notech_or2 i_47953472(.A(n_3983), .B(n_305624320), .Z(n_197762248));
	notech_nand3 i_2820785(.A(n_222862495), .B(n_197662247), .C(n_196862239)
		, .Z(n_24592));
	notech_nao3 i_45553495(.A(opc[27]), .B(n_62782), .C(n_58008), .Z(n_197662247
		));
	notech_and4 i_44753503(.A(n_58815), .B(n_62782), .C(opc_10[27]), .D(n_26599
		), .Z(n_196962240));
	notech_or2 i_45453496(.A(n_4016), .B(n_305624320), .Z(n_196862239));
	notech_nand3 i_2920786(.A(n_222062487), .B(n_221962486), .C(n_195962230)
		, .Z(n_24598));
	notech_or2 i_43553515(.A(n_3982), .B(n_305624320), .Z(n_195962230));
	notech_nand3 i_3020787(.A(n_221262479), .B(n_221162478), .C(n_194962221)
		, .Z(n_24604));
	notech_or2 i_40853540(.A(n_3981), .B(n_305624320), .Z(n_194962221));
	notech_or4 i_2720720(.A(n_194362215), .B(n_219962466), .C(n_194462216), 
		.D(n_193362205), .Z(n_24912));
	notech_ao3 i_38153565(.A(opc[26]), .B(n_62792), .C(n_309391730), .Z(n_194462216
		));
	notech_and2 i_37953567(.A(add_len_pc[26]), .B(n_26766), .Z(n_194362215)
		);
	notech_nand2 i_37853568(.A(sav_epc[26]), .B(n_61143), .Z(n_194262214));
	notech_nor2 i_38053566(.A(n_124328520), .B(n_3983), .Z(n_193362205));
	notech_mux2 i_2711696(.S(n_60550), .A(regs_14[26]), .B(add_len_pc32[26])
		, .Z(add_len_pc[26]));
	notech_or4 i_2820721(.A(n_193162203), .B(n_218962456), .C(n_193262204), 
		.D(n_192162193), .Z(n_24918));
	notech_ao3 i_32853618(.A(opc[27]), .B(n_62782), .C(n_309391730), .Z(n_193262204
		));
	notech_and2 i_32753619(.A(add_len_pc[27]), .B(n_26766), .Z(n_193162203)
		);
	notech_nand2 i_32553621(.A(sav_epc[27]), .B(n_61143), .Z(n_193062202));
	notech_mux2 i_2811697(.S(n_60550), .A(regs_14[27]), .B(add_len_pc32[27])
		, .Z(add_len_pc[27]));
	notech_nor2 i_32653620(.A(n_124328520), .B(n_4016), .Z(n_192162193));
	notech_or4 i_2920722(.A(n_191962191), .B(n_217962446), .C(n_192062192), 
		.D(n_190962181), .Z(n_24924));
	notech_ao3 i_30553641(.A(opc[28]), .B(n_62782), .C(n_309391730), .Z(n_192062192
		));
	notech_and2 i_30353643(.A(add_len_pc[28]), .B(n_26766), .Z(n_191962191)
		);
	notech_nand2 i_30253644(.A(sav_epc[28]), .B(n_61143), .Z(n_191862190));
	notech_nor2 i_30453642(.A(n_124328520), .B(n_3982), .Z(n_190962181));
	notech_mux2 i_2911698(.S(n_60550), .A(regs_14[28]), .B(add_len_pc32[28])
		, .Z(add_len_pc[28]));
	notech_nand3 i_16853767(.A(n_319191632), .B(n_318791636), .C(n_57369), .Z
		(n_190262174));
	notech_nor2 i_30749(.A(n_57026), .B(n_29653), .Z(n_190062172));
	notech_nand2 i_29906(.A(opc[9]), .B(n_62782), .Z(n_189962171));
	notech_ao3 i_49255035(.A(n_32386), .B(n_56485), .C(n_56824), .Z(n_189662168
		));
	notech_ao3 i_49055037(.A(n_32386), .B(n_56921), .C(n_56824), .Z(n_189362166
		));
	notech_or4 i_47655049(.A(n_2938), .B(n_2937), .C(n_56824), .D(n_32291), 
		.Z(n_188562161));
	notech_or4 i_46655059(.A(n_2938), .B(n_2937), .C(n_56822), .D(n_32301), 
		.Z(n_187762157));
	notech_and4 i_46255063(.A(n_56848), .B(n_188562161), .C(n_26812), .D(n_58482
		), .Z(n_187662156));
	notech_mux2 i_170555509(.S(n_60347), .A(n_28089), .B(n_58689), .Z(n_186962151
		));
	notech_and3 i_117157359(.A(n_185262135), .B(n_185362136), .C(n_176762050
		), .Z(n_186762149));
	notech_ao4 i_117257358(.A(n_151761800), .B(n_29755), .C(n_59100), .D(n_28089
		), .Z(n_186462146));
	notech_ao4 i_117357357(.A(n_151961802), .B(n_291263179), .C(n_57841), .D
		(n_291163178), .Z(n_186362145));
	notech_and4 i_118257349(.A(n_185962142), .B(n_185762140), .C(n_185562138
		), .D(n_177462057), .Z(n_186162144));
	notech_ao4 i_117657354(.A(n_59993), .B(n_306091763), .C(n_58409), .D(n_27981
		), .Z(n_185962142));
	notech_ao4 i_117957352(.A(n_60117), .B(n_27116), .C(n_26774), .D(n_175562038
		), .Z(n_185762140));
	notech_ao4 i_118357348(.A(n_24590), .B(\nbus_11358[0] ), .C(n_305991764)
		, .D(\nbus_11307[0] ), .Z(n_185662139));
	notech_ao4 i_118057351(.A(n_24583), .B(n_175462037), .C(n_175062033), .D
		(n_26947), .Z(n_185562138));
	notech_ao4 i_118457347(.A(n_24590), .B(n_60025), .C(n_56037), .D(n_305991764
		), .Z(n_185462137));
	notech_ao4 i_7658415(.A(n_28222), .B(\nbus_11358[0] ), .C(n_298991830), 
		.D(\nbus_11307[0] ), .Z(n_185362136));
	notech_ao4 i_7758414(.A(n_2991), .B(n_60025), .C(n_56037), .D(n_2992), .Z
		(n_185262135));
	notech_and4 i_173356815(.A(n_187968894), .B(n_178362066), .C(n_184862131
		), .D(n_178662069), .Z(n_185162134));
	notech_ao4 i_173156817(.A(n_31411), .B(n_286463131), .C(\nbus_11358[10] 
		), .D(n_26835), .Z(n_184862131));
	notech_ao4 i_173456814(.A(\nbus_11307[10] ), .B(n_285763124), .C(n_291063177
		), .D(n_29684), .Z(n_184662129));
	notech_ao4 i_173556813(.A(n_87532846), .B(n_286263129), .C(n_187568890),
		 .D(n_56625), .Z(n_184462127));
	notech_and4 i_174156807(.A(n_187368889), .B(n_179562078), .C(n_184062123
		), .D(n_179262075), .Z(n_184362126));
	notech_ao4 i_173956809(.A(n_30528), .B(n_56625), .C(n_27996), .D(n_286563132
		), .Z(n_184062123));
	notech_and4 i_174656802(.A(n_183762120), .B(n_180162084), .C(n_183562118
		), .D(n_179862081), .Z(n_183962122));
	notech_ao4 i_174256806(.A(\nbus_11358[11] ), .B(n_26835), .C(\nbus_11307[11] 
		), .D(n_285763124), .Z(n_183762120));
	notech_ao4 i_174456804(.A(n_31492), .B(n_181262095), .C(n_302491799), .D
		(n_181162094), .Z(n_183562118));
	notech_and4 i_175056798(.A(n_180262085), .B(n_183162114), .C(n_26609), .D
		(n_180562088), .Z(n_183462117));
	notech_ao4 i_174856800(.A(n_320070211), .B(n_286463131), .C(n_56221), .D
		(n_26835), .Z(n_183162114));
	notech_ao4 i_175156797(.A(n_57644), .B(n_285763124), .C(n_291063177), .D
		(n_29679), .Z(n_182962112));
	notech_ao4 i_175256796(.A(n_286263129), .B(n_156768584), .C(n_185668873)
		, .D(n_56625), .Z(n_182762110));
	notech_ao4 i_189756653(.A(n_58432), .B(n_5743), .C(n_58391), .D(n_29725)
		, .Z(n_182562108));
	notech_ao4 i_189856652(.A(n_60347), .B(n_28093), .C(n_147071950), .D(\nbus_11307[4] 
		), .Z(n_182362106));
	notech_ao4 i_193156619(.A(n_3852), .B(n_59742), .C(n_26610), .D(n_176262045
		), .Z(n_182262105));
	notech_nand3 i_5858433(.A(n_2988), .B(n_60347), .C(opb[4]), .Z(n_181862101
		));
	notech_and3 i_29560(.A(n_182362106), .B(n_182562108), .C(n_181862101), .Z
		(n_181462097));
	notech_nand2 i_30546(.A(n_26834), .B(n_174962032), .Z(n_181262095));
	notech_or4 i_30547(.A(n_286463131), .B(n_175162034), .C(n_32342), .D(n_26735
		), .Z(n_181162094));
	notech_or2 i_88557637(.A(n_60013), .B(n_285563122), .Z(n_181062093));
	notech_or2 i_89057632(.A(n_286563132), .B(n_27997), .Z(n_180562088));
	notech_or4 i_89157631(.A(n_286463131), .B(n_28138), .C(n_60945), .D(n_54794
		), .Z(n_180262085));
	notech_or4 i_87557647(.A(n_286463131), .B(n_175162034), .C(n_32319), .D(n_29596
		), .Z(n_180162084));
	notech_or4 i_87857644(.A(n_62864), .B(n_62782), .C(n_29596), .D(n_286463131
		), .Z(n_179862081));
	notech_or4 i_88157641(.A(n_286463131), .B(n_60947), .C(n_28137), .D(n_54794
		), .Z(n_179562078));
	notech_nao3 i_88257640(.A(n_62826), .B(opc[11]), .C(n_286263129), .Z(n_179262075
		));
	notech_or2 i_86657656(.A(n_3850), .B(n_285563122), .Z(n_179162074));
	notech_or2 i_87157651(.A(n_286563132), .B(n_27993), .Z(n_178662069));
	notech_or4 i_87257650(.A(n_54774), .B(n_60947), .C(n_28136), .D(n_54794)
		, .Z(n_178362066));
	notech_or4 i_29958194(.A(n_62864), .B(n_281463081), .C(n_60945), .D(n_56037
		), .Z(n_177462057));
	notech_nand3 i_30458189(.A(n_310991714), .B(\regs_1[0] ), .C(n_28680), .Z
		(n_176762050));
	notech_and3 i_11758374(.A(n_26702), .B(n_26643), .C(n_26634), .Z(n_176562048
		));
	notech_nand2 i_105857469(.A(n_2988), .B(opb[0]), .Z(n_176362046));
	notech_ao4 i_13758356(.A(n_60025), .B(n_26602), .C(n_56037), .D(n_176562048
		), .Z(n_176262045));
	notech_nand2 i_81761828(.A(n_24582), .B(n_306791756), .Z(n_175762040));
	notech_and2 i_17058323(.A(n_58646), .B(n_185662139), .Z(n_175562038));
	notech_and2 i_16958324(.A(n_185462137), .B(n_58610), .Z(n_175462037));
	notech_ao4 i_16858325(.A(n_30854), .B(n_26062), .C(n_175762040), .D(n_26775
		), .Z(n_175362036));
	notech_nand2 i_161361795(.A(n_26718), .B(n_26775), .Z(n_175262035));
	notech_ao4 i_82964500(.A(n_60893), .B(n_26945), .C(n_62782), .D(n_60910)
		, .Z(n_175162034));
	notech_nao3 i_117758476(.A(n_62826), .B(opa[0]), .C(n_62848), .Z(n_175062033
		));
	notech_or4 i_11664510(.A(n_57026), .B(n_29653), .C(n_29658), .D(instrc[
		116]), .Z(n_174962032));
	notech_and4 i_130960489(.A(n_174662029), .B(n_174462027), .C(n_174362026
		), .D(n_153861821), .Z(n_174862031));
	notech_ao4 i_130360494(.A(n_291663183), .B(n_281363080), .C(n_57889), .D
		(\nbus_11307[4] ), .Z(n_174662029));
	notech_ao4 i_130560492(.A(n_57890), .B(\nbus_11358[4] ), .C(n_24583), .D
		(n_291463181), .Z(n_174462027));
	notech_ao4 i_130660491(.A(n_5723), .B(n_306091763), .C(n_57841), .D(n_291863185
		), .Z(n_174362026));
	notech_and4 i_131660482(.A(n_174062023), .B(n_173962022), .C(n_173762020
		), .D(n_173662019), .Z(n_174262025));
	notech_ao4 i_131060488(.A(n_60117), .B(n_27121), .C(n_58409), .D(n_27986
		), .Z(n_174062023));
	notech_ao4 i_131160487(.A(n_291563182), .B(n_26774), .C(n_5743), .D(n_58004
		), .Z(n_173962022));
	notech_ao4 i_131360485(.A(n_58003), .B(n_29725), .C(n_151761800), .D(n_29745
		), .Z(n_173762020));
	notech_ao4 i_131460484(.A(n_151861801), .B(n_29746), .C(n_291763184), .D
		(n_151961802), .Z(n_173662019));
	notech_and4 i_132260476(.A(n_62935425), .B(n_173362016), .C(n_173162014)
		, .D(n_173062013), .Z(n_173562018));
	notech_ao4 i_131760481(.A(n_24583), .B(n_31279), .C(n_59100), .D(n_28096
		), .Z(n_173362016));
	notech_ao4 i_131960479(.A(n_303391790), .B(n_306091763), .C(n_31309), .D
		(n_57841), .Z(n_173162014));
	notech_ao4 i_132060478(.A(n_60117), .B(n_27126), .C(n_58409), .D(n_56100
		), .Z(n_173062013));
	notech_and4 i_132860470(.A(n_172762010), .B(n_172562008), .C(n_172462007
		), .D(n_155961842), .Z(n_172962012));
	notech_ao4 i_132360475(.A(n_58003), .B(n_29614), .C(\nbus_11307[7] ), .D
		(n_26773), .Z(n_172762010));
	notech_ao4 i_132560473(.A(\nbus_11358[7] ), .B(n_57615), .C(n_151761800)
		, .D(n_29747), .Z(n_172562008));
	notech_ao4 i_132660472(.A(n_151861801), .B(n_29748), .C(n_31307), .D(n_151961802
		), .Z(n_172462007));
	notech_and4 i_133460465(.A(n_172162004), .B(n_156961852), .C(n_171962002
		), .D(n_156661849), .Z(n_172362006));
	notech_ao4 i_133060469(.A(n_59100), .B(n_28098), .C(n_59968), .D(n_305791766
		), .Z(n_172162004));
	notech_ao4 i_133260467(.A(n_60117), .B(n_27129), .C(n_58381), .D(n_27992
		), .Z(n_171962002));
	notech_and4 i_134060459(.A(n_171661999), .B(n_171461997), .C(n_171361996
		), .D(n_157261855), .Z(n_171862001));
	notech_ao4 i_133560464(.A(\nbus_11358[9] ), .B(n_57983), .C(n_57937), .D
		(n_60016), .Z(n_171661999));
	notech_ao4 i_133760462(.A(n_57936), .B(n_29743), .C(n_151761800), .D(n_29749
		), .Z(n_171461997));
	notech_ao4 i_133860461(.A(n_151861801), .B(n_29750), .C(n_152061803), .D
		(n_189962171), .Z(n_171361996));
	notech_and4 i_134660453(.A(n_65435450), .B(n_171061993), .C(n_170861991)
		, .D(n_170761990), .Z(n_171261995));
	notech_ao4 i_134160458(.A(n_31456), .B(n_24589), .C(n_59100), .D(n_28100
		), .Z(n_171061993));
	notech_ao4 i_134360456(.A(n_302891795), .B(n_305791766), .C(n_31476), .D
		(n_57799), .Z(n_170861991));
	notech_ao4 i_134460455(.A(n_60117), .B(n_27131), .C(n_58381), .D(n_27996
		), .Z(n_170761990));
	notech_and4 i_135360446(.A(n_170461987), .B(n_170361986), .C(n_170161984
		), .D(n_170061983), .Z(n_170661989));
	notech_ao4 i_134760452(.A(n_57984), .B(\nbus_11307[11] ), .C(n_57983), .D
		(\nbus_11358[11] ), .Z(n_170461987));
	notech_ao4 i_134860451(.A(n_31492), .B(n_175262035), .C(n_151761800), .D
		(n_29751), .Z(n_170361986));
	notech_ao4 i_135060449(.A(n_151861801), .B(n_29752), .C(n_30088), .D(n_152061803
		), .Z(n_170161984));
	notech_ao4 i_135160448(.A(n_302491799), .B(n_188857101), .C(n_169761980)
		, .D(n_29596), .Z(n_170061983));
	notech_nao3 i_174161736(.A(n_58009), .B(n_26775), .C(n_307691747), .Z(n_169761980
		));
	notech_and4 i_140160399(.A(n_162665155), .B(n_169361976), .C(n_169161974
		), .D(n_159561878), .Z(n_169561978));
	notech_ao4 i_139760403(.A(\nbus_11358[15] ), .B(n_307591748), .C(n_59100
		), .D(n_28104), .Z(n_169361976));
	notech_ao4 i_139960401(.A(n_298466513), .B(n_57799), .C(n_60117), .D(n_27136
		), .Z(n_169161974));
	notech_ao4 i_140260398(.A(n_151861801), .B(n_29753), .C(n_320137996), .D
		(n_56553), .Z(n_168861971));
	notech_nao3 i_140560395(.A(n_159961882), .B(n_26953), .C(n_160161884), .Z
		(n_168761970));
	notech_ao4 i_140960392(.A(n_60010), .B(n_24590), .C(n_305891765), .D(n_29754
		), .Z(n_168561968));
	notech_ao4 i_140860393(.A(n_307391750), .B(\nbus_11307[15] ), .C(n_111064639
		), .D(n_26718), .Z(n_168361966));
	notech_and4 i_207959759(.A(n_93835734), .B(n_160961892), .C(n_167961962)
		, .D(n_160661889), .Z(n_168261965));
	notech_ao4 i_207759761(.A(n_286563132), .B(n_27998), .C(n_31540), .D(n_54774
		), .Z(n_167961962));
	notech_and4 i_208459754(.A(n_167661959), .B(n_161561898), .C(n_167461957
		), .D(n_161261895), .Z(n_167861961));
	notech_ao4 i_208059758(.A(\nbus_11307[13] ), .B(n_285763124), .C(n_302091803
		), .D(n_181162094), .Z(n_167661959));
	notech_ao4 i_208259756(.A(n_30109), .B(n_286263129), .C(n_94935745), .D(n_56625
		), .Z(n_167461957));
	notech_and4 i_208859750(.A(n_140168418), .B(n_161961902), .C(n_167061953
		), .D(n_161661899), .Z(n_167361956));
	notech_ao4 i_208659752(.A(n_286563132), .B(n_27999), .C(n_298166510), .D
		(n_54774), .Z(n_167061953));
	notech_and4 i_209359745(.A(n_166761950), .B(n_166561948), .C(n_162261905
		), .D(n_162561908), .Z(n_166961952));
	notech_ao4 i_208959749(.A(n_57662), .B(n_285763124), .C(n_60011), .D(n_181162094
		), .Z(n_166761950));
	notech_ao4 i_209159747(.A(n_157165100), .B(n_286263129), .C(n_139068407)
		, .D(n_56625), .Z(n_166561948));
	notech_and4 i_209759741(.A(n_128171761), .B(n_162661909), .C(n_166161944
		), .D(n_162961912), .Z(n_166461947));
	notech_ao4 i_209559743(.A(n_136561648), .B(n_28000), .C(n_152661809), .D
		(\nbus_11358[15] ), .Z(n_166161944));
	notech_ao4 i_209859740(.A(n_60010), .B(n_285563122), .C(n_291063177), .D
		(n_29754), .Z(n_165961942));
	notech_ao4 i_209959739(.A(n_58105), .B(n_56625), .C(n_111064639), .D(n_152461807
		), .Z(n_165761940));
	notech_ao4 i_210259736(.A(n_60347), .B(n_28121), .C(n_32252), .D(n_309721261
		), .Z(n_165561938));
	notech_ao4 i_210359735(.A(n_58426), .B(n_28015), .C(n_250962776), .D(\nbus_11365[30] 
		), .Z(n_165461937));
	notech_and3 i_210859730(.A(n_165061933), .B(n_165261935), .C(n_164261925
		), .Z(n_165361936));
	notech_ao4 i_210559733(.A(n_251362780), .B(\nbus_11358[30] ), .C(n_302991794
		), .D(n_251262779), .Z(n_165261935));
	notech_ao4 i_210659732(.A(n_303091793), .B(n_322438019), .C(n_30809), .D
		(n_316537960), .Z(n_165061933));
	notech_nand3 i_187364474(.A(n_56848), .B(n_127161554), .C(n_285463121), 
		.Z(n_164961932));
	notech_and2 i_225159587(.A(n_285563122), .B(n_274863015), .Z(n_164761930
		));
	notech_nao3 i_13627(.A(n_32319), .B(n_26763), .C(n_175162034), .Z(n_164361926
		));
	notech_or2 i_100860755(.A(n_251162778), .B(n_29591), .Z(n_164261925));
	notech_nand2 i_99960764(.A(opa[15]), .B(n_152561808), .Z(n_163461917));
	notech_or4 i_100460759(.A(n_62864), .B(n_62782), .C(n_56266), .D(n_54774
		), .Z(n_162961912));
	notech_or4 i_100560758(.A(n_54774), .B(n_28141), .C(n_60938), .D(n_54794
		), .Z(n_162661909));
	notech_or4 i_98760774(.A(n_54774), .B(n_175162034), .C(n_32319), .D(n_56257
		), .Z(n_162561908));
	notech_nand2 i_99060771(.A(n_286663133), .B(opb[14]), .Z(n_162261905));
	notech_or4 i_99360768(.A(n_54774), .B(n_28140), .C(n_60928), .D(n_54794)
		, .Z(n_161961902));
	notech_or4 i_99460767(.A(n_62864), .B(n_181262095), .C(n_60928), .D(n_29680
		), .Z(n_161661899));
	notech_or4 i_97760784(.A(n_54774), .B(n_175162034), .C(n_32319), .D(n_29592
		), .Z(n_161561898));
	notech_nand2 i_98060781(.A(opb[13]), .B(n_286663133), .Z(n_161261895));
	notech_or4 i_98360778(.A(n_54774), .B(n_60928), .C(n_28139), .D(n_54794)
		, .Z(n_160961892));
	notech_or4 i_98460777(.A(n_62864), .B(n_181262095), .C(n_60928), .D(n_29592
		), .Z(n_160661889));
	notech_ao4 i_20961519(.A(n_2349), .B(n_1440), .C(n_152361806), .D(n_26955
		), .Z(n_160161884));
	notech_ao4 i_20861520(.A(n_234791985), .B(n_1442), .C(n_26646), .D(n_26954
		), .Z(n_160061883));
	notech_or4 i_20761521(.A(n_26718), .B(nbus_11295[15]), .C(n_60928), .D(n_307491749
		), .Z(n_159961882));
	notech_and3 i_21261516(.A(n_8129), .B(n_60550), .C(n_310991714), .Z(n_159861881
		));
	notech_nao3 i_21561513(.A(opa[15]), .B(n_27274), .C(n_307391750), .Z(n_159561878
		));
	notech_or2 i_14561583(.A(n_57984), .B(\nbus_11307[9] ), .Z(n_157261855)
		);
	notech_or4 i_14861580(.A(n_56863), .B(n_26062), .C(n_291963186), .D(n_24589
		), .Z(n_156961852));
	notech_or4 i_15161577(.A(n_62830), .B(n_62782), .C(n_56127), .D(n_24589)
		, .Z(n_156661849));
	notech_or2 i_13261596(.A(n_303191792), .B(n_58004), .Z(n_155961842));
	notech_or4 i_12561603(.A(n_61143), .B(n_60292), .C(n_19086), .D(n_28093)
		, .Z(n_153861821));
	notech_or4 i_122960564(.A(n_32326), .B(n_32614), .C(n_307691747), .D(n_24583
		), .Z(n_153561818));
	notech_nand3 i_119460597(.A(n_146961752), .B(n_285463121), .C(n_286463131
		), .Z(n_152961812));
	notech_and3 i_119360598(.A(n_58505), .B(n_58489), .C(n_58481), .Z(n_152861811
		));
	notech_and3 i_118460607(.A(n_24582), .B(n_306791756), .C(n_24583), .Z(n_152761810
		));
	notech_and2 i_160164480(.A(n_275963026), .B(n_274863015), .Z(n_152661809
		));
	notech_ao4 i_147264484(.A(n_59445), .B(n_26833), .C(n_164961932), .D(n_26763
		), .Z(n_152561808));
	notech_and2 i_149564483(.A(n_274763014), .B(n_126961552), .Z(n_152461807
		));
	notech_nor2 i_22261506(.A(n_24590), .B(\nbus_11358[15] ), .Z(n_152361806
		));
	notech_or4 i_130861753(.A(n_26062), .B(n_57088), .C(n_29652), .D(n_152761810
		), .Z(n_152061803));
	notech_or4 i_124561755(.A(n_55581), .B(n_57088), .C(n_29652), .D(n_26774
		), .Z(n_151961802));
	notech_or4 i_63061773(.A(n_61143), .B(n_60292), .C(n_26983), .D(n_60550)
		, .Z(n_151861801));
	notech_or4 i_62961774(.A(n_61143), .B(n_60303), .C(n_26983), .D(n_28680)
		, .Z(n_151761800));
	notech_nand2 i_13613(.A(n_285863125), .B(n_26763), .Z(n_151661799));
	notech_ao4 i_141763075(.A(n_285363120), .B(\nbus_11358[0] ), .C(n_291163178
		), .D(n_274763014), .Z(n_151361796));
	notech_and4 i_142363070(.A(n_131361596), .B(n_151161794), .C(n_131561598
		), .D(n_26961), .Z(n_151261795));
	notech_ao4 i_142063073(.A(n_56046), .B(n_296863235), .C(n_291363180), .D
		(n_136161644), .Z(n_151161794));
	notech_ao4 i_142563068(.A(n_125561538), .B(n_56028), .C(n_140661689), .D
		(n_59742), .Z(n_150661789));
	notech_and4 i_143063063(.A(n_228879789), .B(n_150161784), .C(n_131961602
		), .D(n_132261605), .Z(n_150461787));
	notech_ao4 i_142863065(.A(n_298066509), .B(n_274763014), .C(n_297766506)
		, .D(n_275363020), .Z(n_150161784));
	notech_and4 i_143563058(.A(n_149861781), .B(n_132861611), .C(n_149661779
		), .D(n_132561608), .Z(n_150061783));
	notech_ao4 i_143163062(.A(n_253640554), .B(n_56625), .C(n_297966508), .D
		(n_136261645), .Z(n_149861781));
	notech_ao4 i_143363060(.A(n_136461647), .B(n_29678), .C(n_136061643), .D
		(\nbus_11307[1] ), .Z(n_149661779));
	notech_and4 i_143963054(.A(n_181462097), .B(n_149261775), .C(n_132961612
		), .D(n_133261615), .Z(n_149561778));
	notech_ao4 i_143763056(.A(n_291863185), .B(n_274763014), .C(n_291563182)
		, .D(n_275363020), .Z(n_149261775));
	notech_and4 i_144463049(.A(n_148961772), .B(n_148761770), .C(n_133561618
		), .D(n_133861621), .Z(n_149161774));
	notech_ao4 i_144063053(.A(n_56625), .B(n_253740555), .C(n_136261645), .D
		(n_291763184), .Z(n_148961772));
	notech_ao4 i_144263051(.A(n_136461647), .B(n_29725), .C(\nbus_11307[4] )
		, .D(n_136061643), .Z(n_148761770));
	notech_nand2 i_144763046(.A(n_148361766), .B(n_134261625), .Z(n_148461767
		));
	notech_ao4 i_144663047(.A(n_58426), .B(n_56100), .C(n_56109), .D(n_285363120
		), .Z(n_148361766));
	notech_and4 i_145363040(.A(n_134561628), .B(n_148061763), .C(n_147861761
		), .D(n_134861631), .Z(n_148261765));
	notech_ao4 i_144963044(.A(n_296863235), .B(n_303191792), .C(n_31307), .D
		(n_136261645), .Z(n_148061763));
	notech_ao4 i_145163042(.A(n_136461647), .B(n_29614), .C(n_275363020), .D
		(n_126661549), .Z(n_147861761));
	notech_ao4 i_145463039(.A(n_125561538), .B(n_56109), .C(n_57957), .D(n_140661689
		), .Z(n_147761760));
	notech_and3 i_145763036(.A(n_200065529), .B(n_147461757), .C(n_135161634
		), .Z(n_147661759));
	notech_ao4 i_145663037(.A(n_291063177), .B(n_56127), .C(n_291963186), .D
		(n_290963176), .Z(n_147461757));
	notech_ao4 i_145863035(.A(n_58608), .B(n_54774), .C(\nbus_11307[9] ), .D
		(n_26958), .Z(n_147261755));
	notech_ao4 i_145963034(.A(\nbus_11358[9] ), .B(n_152661809), .C(n_252740545
		), .D(n_56625), .Z(n_147061753));
	notech_ao4 i_5064403(.A(n_56854), .B(n_26962), .C(n_32352), .D(n_32287),
		 .Z(n_146961752));
	notech_and2 i_141864451(.A(n_146361746), .B(n_144961732), .Z(n_146461747
		));
	notech_ao4 i_162662875(.A(n_61117), .B(n_128261565), .C(n_128161564), .D
		(n_27084), .Z(n_146361746));
	notech_ao4 i_162862873(.A(n_60868), .B(n_319691627), .C(n_60893), .D(n_2884
		), .Z(n_146061743));
	notech_and3 i_163162870(.A(n_1870), .B(n_1871), .C(n_2678), .Z(n_145961742
		));
	notech_and4 i_163862863(.A(n_23007), .B(n_2684), .C(n_2677), .D(n_145461737
		), .Z(n_145761740));
	notech_and4 i_163762864(.A(n_58072), .B(n_145361736), .C(n_32652), .D(n_137661659
		), .Z(n_145461737));
	notech_and4 i_163562866(.A(n_1906), .B(n_1907), .C(n_2895), .D(n_137861661
		), .Z(n_145361736));
	notech_ao4 i_162762874(.A(n_59322), .B(n_128061563), .C(n_144261725), .D
		(n_144361726), .Z(n_144961732));
	notech_ao4 i_5164402(.A(n_26900), .B(n_319963466), .C(n_5380), .D(n_125361536
		), .Z(n_144861731));
	notech_or4 i_164262859(.A(n_32596), .B(n_32555), .C(n_19006), .D(n_19057
		), .Z(n_144761730));
	notech_or4 i_164662856(.A(n_32581), .B(n_59322), .C(n_26900), .D(n_29744
		), .Z(n_144361726));
	notech_or4 i_164762855(.A(n_27037), .B(n_26757), .C(n_19086), .D(n_19079
		), .Z(n_144261725));
	notech_ao4 i_162562876(.A(n_248240500), .B(n_27896), .C(n_144061723), .D
		(n_252140539), .Z(n_144161724));
	notech_or4 i_164862854(.A(n_1864), .B(n_28079), .C(n_61143), .D(n_60229)
		, .Z(n_144061723));
	notech_and4 i_172162781(.A(n_19065), .B(n_19072), .C(n_137961662), .D(n_26985
		), .Z(n_143861721));
	notech_or4 i_172662777(.A(n_19022), .B(n_19036), .C(n_32555), .D(n_143261715
		), .Z(n_143561718));
	notech_or4 i_172462779(.A(n_27037), .B(n_3790), .C(n_3923), .D(n_19086),
		 .Z(n_143261715));
	notech_ao4 i_177862725(.A(n_26981), .B(n_252940547), .C(n_125561538), .D
		(n_129461577), .Z(n_142761710));
	notech_ao4 i_178762716(.A(n_30294), .B(n_142361706), .C(n_142261705), .D
		(n_26735), .Z(n_142461707));
	notech_nao3 i_12164333(.A(instrc[125]), .B(n_26849), .C(instrc[126]), .Z
		(n_142361706));
	notech_ao4 i_92170128(.A(n_154379047), .B(n_27766), .C(n_27107), .D(n_27422
		), .Z(n_113978643));
	notech_ao4 i_92070129(.A(n_154179045), .B(n_56037), .C(n_27728), .D(n_154279046
		), .Z(n_114078644));
	notech_and2 i_1567385(.A(n_30303), .B(n_131578819), .Z(n_114178645));
	notech_nao3 i_2367377(.A(n_126178765), .B(instrc[107]), .C(n_30933), .Z(n_114278646
		));
	notech_nand2 i_1267388(.A(n_27198), .B(n_27192), .Z(n_114378647));
	notech_or4 i_21767201(.A(n_32326), .B(n_32614), .C(n_32334), .D(n_3730),
		 .Z(n_114578649));
	notech_or4 i_21967200(.A(n_30344), .B(n_57026), .C(n_56863), .D(instrc[
		119]), .Z(n_114678650));
	notech_nand3 i_22067199(.A(n_26858), .B(n_28130), .C(n_29667), .Z(n_114778651
		));
	notech_or4 i_22167198(.A(n_29633), .B(n_57462), .C(instrc[103]), .D(n_26724
		), .Z(n_114878652));
	notech_or4 i_22267197(.A(n_190010112), .B(n_29642), .C(instrc[90]), .D(n_26727
		), .Z(n_114978653));
	notech_or4 i_22367196(.A(instrc[105]), .B(n_57369), .C(n_26728), .D(n_26892
		), .Z(n_115078654));
	notech_nand3 i_22467195(.A(n_125078754), .B(n_29638), .C(n_29636), .Z(n_115178655
		));
	notech_ao4 i_2467376(.A(n_59445), .B(n_27079), .C(n_32380), .D(n_56939),
		 .Z(n_115978663));
	notech_ao4 i_4667355(.A(n_116378667), .B(n_24590), .C(n_56822), .D(n_56553
		), .Z(n_116178665));
	notech_ao4 i_467391(.A(n_56822), .B(n_32280), .C(n_2480), .D(n_62892), .Z
		(n_116378667));
	notech_ao4 i_4867353(.A(n_123978743), .B(n_26719), .C(n_26718), .D(n_60928
		), .Z(n_116478668));
	notech_or4 i_25367167(.A(instrc[122]), .B(n_32614), .C(n_30312), .D(instrc
		[121]), .Z(n_116578669));
	notech_and4 i_7667325(.A(n_115078654), .B(n_124778751), .C(n_114978653),
		 .D(n_115178655), .Z(n_116678670));
	notech_nao3 i_25567165(.A(n_60117), .B(n_27714), .C(n_116878672), .Z(n_116778671
		));
	notech_ao4 i_7567326(.A(n_116478668), .B(n_116378667), .C(n_116178665), 
		.D(1'b0), .Z(n_116878672));
	notech_nand2 i_7467327(.A(n_3835), .B(n_116578669), .Z(n_116978673));
	notech_ao4 i_4567356(.A(n_7298943), .B(n_3593), .C(n_252940547), .D(n_30294
		), .Z(n_117078674));
	notech_nand3 i_25667164(.A(n_60122), .B(n_60292), .C(n_116978673), .Z(n_117178675
		));
	notech_or4 i_25767163(.A(instrc[127]), .B(n_340380904), .C(n_117078674),
		 .D(n_29632), .Z(n_117278676));
	notech_or2 i_25467166(.A(n_116678670), .B(n_252940547), .Z(n_117378677)
		);
	notech_nao3 i_50691(.A(n_116778671), .B(n_126078764), .C(n_349480995), .Z
		(\nbus_11330[0] ));
	notech_nand3 i_36967057(.A(n_3914), .B(n_11064), .C(n_114278646), .Z(n_117678680
		));
	notech_nor2 i_36867058(.A(n_349880999), .B(n_27769), .Z(n_117978683));
	notech_nao3 i_418265(.A(n_126578769), .B(n_117678680), .C(n_117978683), 
		.Z(write_data_28[3]));
	notech_and2 i_37367053(.A(imm[0]), .B(n_329263509), .Z(n_118078684));
	notech_nand2 i_6867333(.A(n_56579), .B(n_56557), .Z(n_118178685));
	notech_and2 i_37667051(.A(opz[0]), .B(n_118178685), .Z(n_118278686));
	notech_and4 i_37567052(.A(n_59387), .B(n_114378647), .C(instrc[115]), .D
		(instrc[104]), .Z(n_118378687));
	notech_nand2 i_38367044(.A(imm[1]), .B(n_329263509), .Z(n_118478688));
	notech_nand3 i_38467043(.A(n_114378647), .B(n_56925), .C(instrc[105]), .Z
		(n_118778691));
	notech_nand2 i_39267035(.A(imm[2]), .B(n_329263509), .Z(n_118878692));
	notech_ao3 i_5267349(.A(instrc[115]), .B(n_59397), .C(n_59387), .Z(n_119078694
		));
	notech_nand3 i_39367034(.A(n_56925), .B(n_114378647), .C(n_57369), .Z(n_119278696
		));
	notech_ao4 i_315640(.A(n_62041235), .B(n_28091), .C(n_317887452), .D(n_28389
		), .Z(n_22730));
	notech_and4 i_172967436(.A(n_127678780), .B(n_127578779), .C(n_119278696
		), .D(n_118878692), .Z(nbus_11317_2100235));
	notech_nand2 i_119966229(.A(opd[2]), .B(n_329963516), .Z(n_119578699));
	notech_or4 i_119866230(.A(n_55508), .B(n_59241), .C(n_27981), .D(opd[2])
		, .Z(n_120478708));
	notech_or2 i_119466234(.A(nbus_11317_2100235), .B(n_329363510), .Z(n_120578709
		));
	notech_or2 i_119666232(.A(n_329463511), .B(n_29054), .Z(n_120678710));
	notech_nand3 i_312920(.A(n_128978793), .B(n_128878792), .C(n_119578699),
		 .Z(n_25958));
	notech_or2 i_122366205(.A(n_329663513), .B(n_27981), .Z(n_120978713));
	notech_or4 i_121966209(.A(n_25625), .B(n_25617), .C(n_190710119), .D(\nbus_11307[1] 
		), .Z(n_121678720));
	notech_nao3 i_122566203(.A(opd[1]), .B(n_59187), .C(n_55508), .Z(n_121778721
		));
	notech_or2 i_122066208(.A(n_349680997100234), .B(n_329363510), .Z(n_121878722
		));
	notech_or2 i_122266206(.A(n_329463511), .B(n_29053), .Z(n_121978723));
	notech_and4 i_212919(.A(n_129878802), .B(n_130078804), .C(n_121978723), 
		.D(n_120978713), .Z(n_25953));
	notech_ao4 i_124666182(.A(n_118078684), .B(n_127078774), .C(n_121261495)
		, .D(n_26781), .Z(n_123078734));
	notech_nor2 i_124866180(.A(n_329463511), .B(n_29052), .Z(n_123178735));
	notech_or4 i_112918(.A(n_123078734), .B(n_123178735), .C(n_26729), .D(n_26730
		), .Z(n_25948));
	notech_nand2 i_152665903(.A(write_data_33[2]), .B(n_60229), .Z(n_123778741
		));
	notech_nand3 i_318808(.A(n_131378817), .B(n_131278816), .C(n_123778741),
		 .Z(n_25714));
	notech_or4 i_25067170(.A(n_340380904), .B(n_32747), .C(instrc[127]), .D(n_29632
		), .Z(n_123978743));
	notech_and4 i_24167179(.A(n_114678650), .B(n_114578649), .C(n_114878652)
		, .D(n_114778651), .Z(n_124778751));
	notech_and3 i_23667183(.A(n_29666), .B(instrc[92]), .C(n_30366), .Z(n_125078754
		));
	notech_and4 i_26267159(.A(n_3821), .B(n_117278676), .C(n_117378677), .D(n_117178675
		), .Z(n_126078764));
	notech_ao4 i_1667384(.A(n_57369), .B(instrc[105]), .C(n_30939), .D(n_29735
		), .Z(n_126178765));
	notech_ao4 i_37067056(.A(n_349780998), .B(n_27731), .C(n_3914), .D(n_27428
		), .Z(n_126578769));
	notech_or4 i_37967048(.A(n_32284), .B(n_119078694), .C(n_118278686), .D(n_118378687
		), .Z(n_127078774));
	notech_ao4 i_38567042(.A(n_28050), .B(n_56579), .C(n_59275), .D(n_27577)
		, .Z(n_127178775));
	notech_ao4 i_38667041(.A(n_29177), .B(n_26720), .C(n_57940), .D(n_56557)
		, .Z(n_127278776));
	notech_ao4 i_39467033(.A(n_59275), .B(n_59355), .C(n_28051), .D(n_56579)
		, .Z(n_127578779));
	notech_ao4 i_39567032(.A(n_57710), .B(n_56553), .C(n_29177), .D(n_26720)
		, .Z(n_127678780));
	notech_ao4 i_120066228(.A(n_40241017), .B(n_29088), .C(n_39041005), .D(n_28928
		), .Z(n_127978783));
	notech_ao4 i_120166227(.A(n_53841153), .B(n_30020), .C(n_54141156), .D(n_30019
		), .Z(n_128078784));
	notech_ao4 i_120266226(.A(n_53341148), .B(nbus_11295[2]), .C(n_53641151)
		, .D(n_57552), .Z(n_128278786));
	notech_ao4 i_120366225(.A(n_1894), .B(n_60229), .C(n_58768), .D(n_30021)
		, .Z(n_128378787));
	notech_and4 i_120666222(.A(n_128378787), .B(n_128278786), .C(n_128078784
		), .D(n_127978783), .Z(n_128578789));
	notech_and4 i_120966219(.A(n_120478708), .B(n_128578789), .C(n_120578709
		), .D(n_120678710), .Z(n_128878792));
	notech_ao4 i_121066218(.A(n_25540870), .B(n_330863525), .C(n_24540860), 
		.D(n_28091), .Z(n_128978793));
	notech_ao4 i_122766201(.A(n_53841153), .B(n_30023), .C(n_54141156), .D(n_30022
		), .Z(n_129178795));
	notech_ao4 i_122866200(.A(n_58768), .B(n_30024), .C(n_53341148), .D(nbus_11295
		[1]), .Z(n_129278796));
	notech_ao4 i_122666202(.A(n_40241017), .B(n_29087), .C(n_39041005), .D(n_28927
		), .Z(n_129478798));
	notech_and3 i_123166197(.A(n_129478798), .B(n_121678720), .C(n_121778721
		), .Z(n_129678800));
	notech_and4 i_123366195(.A(n_129278796), .B(n_129178795), .C(n_129678800
		), .D(n_121878722), .Z(n_129878802));
	notech_ao4 i_123566193(.A(n_25540870), .B(opd[1]), .C(n_24540860), .D(n_28090
		), .Z(n_130078804));
	notech_ao4 i_124966179(.A(n_40241017), .B(n_29086), .C(n_39041005), .D(n_28926
		), .Z(n_130278806));
	notech_ao4 i_125066178(.A(n_53841153), .B(n_30027), .C(n_54141156), .D(n_30026
		), .Z(n_130378807));
	notech_ao4 i_125166177(.A(n_53341148), .B(nbus_11295[0]), .C(n_53641151)
		, .D(n_59742), .Z(n_130578809));
	notech_ao4 i_125266176(.A(n_55508), .B(opd[0]), .C(n_58768), .D(n_30029)
		, .Z(n_130678810));
	notech_and4 i_125566173(.A(n_130678810), .B(n_130578809), .C(n_130378807
		), .D(n_130278806), .Z(n_130878812));
	notech_ao4 i_125866170(.A(n_27040885), .B(opd[0]), .C(n_24540860), .D(n_28089
		), .Z(n_131178815));
	notech_ao4 i_152865901(.A(n_318291641), .B(n_55992), .C(n_318391640), .D
		(nbus_11295[2]), .Z(n_131278816));
	notech_ao4 i_152765902(.A(n_315391670), .B(n_27860), .C(n_59152), .D(n_28453
		), .Z(n_131378817));
	notech_nand2 i_138464463(.A(n_29735), .B(instrc[107]), .Z(n_131578819)
		);
	notech_nand2 i_3864415(.A(n_26973), .B(n_160079104), .Z(n_131678820));
	notech_and4 i_5664397(.A(n_340380904), .B(instrc[127]), .C(n_26891), .D(n_133378837
		), .Z(n_131778821));
	notech_nao3 i_10364350(.A(n_305391770), .B(n_253162798), .C(n_254240560)
		, .Z(n_131878822));
	notech_nand2 i_15564299(.A(n_57901), .B(n_132178825), .Z(n_131978823));
	notech_ao4 i_15664298(.A(n_59435), .B(n_56037), .C(n_58087), .D(n_132378827
		), .Z(n_132078824));
	notech_or4 i_78963684(.A(n_56863), .B(n_54727), .C(n_58480), .D(n_60928)
		, .Z(n_132178825));
	notech_mux2 i_9964354(.S(n_32338), .A(n_56037), .B(n_56046), .Z(n_132378827
		));
	notech_nand3 i_84963626(.A(n_254240560), .B(n_32338), .C(n_26731), .Z(n_132978833
		));
	notech_or4 i_86063616(.A(n_57026), .B(n_56863), .C(n_29653), .D(n_133178835
		), .Z(n_133078834));
	notech_and3 i_14964305(.A(n_56848), .B(n_125961542), .C(n_58493), .Z(n_133178835
		));
	notech_or4 i_86463612(.A(n_32326), .B(n_32339), .C(n_57827), .D(n_58132)
		, .Z(n_133278836));
	notech_nand2 i_88563591(.A(instrc[124]), .B(n_26968), .Z(n_133378837));
	notech_ao3 i_13564319(.A(n_184658942), .B(n_133878842), .C(n_3823), .Z(n_133478838
		));
	notech_ao4 i_13664318(.A(instrc[124]), .B(n_343180932), .C(n_3908), .D(n_160079104
		), .Z(n_133578839));
	notech_nand2 i_101963461(.A(n_56498), .B(n_27033), .Z(n_133878842));
	notech_and2 i_102263458(.A(n_56498), .B(n_26836), .Z(n_134178845));
	notech_ao3 i_102363457(.A(n_345280953), .B(n_26849), .C(n_57500), .Z(n_134278846
		));
	notech_ao3 i_13364321(.A(n_184658942), .B(n_27034), .C(n_134678850), .Z(n_134378847
		));
	notech_ao4 i_3264421(.A(n_56909), .B(n_58132), .C(n_164179145), .D(n_26973
		), .Z(n_134478848));
	notech_and4 i_13464320(.A(n_30905), .B(n_3828), .C(n_27035), .D(n_134778851
		), .Z(n_134578849));
	notech_and2 i_103563445(.A(n_341380914), .B(n_56921), .Z(n_134678850));
	notech_nand2 i_103663444(.A(n_56914), .B(n_26836), .Z(n_134778851));
	notech_ao4 i_10464349(.A(n_59445), .B(n_26792), .C(n_135578859), .D(n_26734
		), .Z(n_134978853));
	notech_ao4 i_12964325(.A(n_3824), .B(n_54765), .C(n_3829), .D(n_57322), 
		.Z(n_135078854));
	notech_nand3 i_7064383(.A(n_27035), .B(n_30905), .C(n_135878862), .Z(n_135578859
		));
	notech_ao4 i_6264391(.A(n_56946), .B(n_3695), .C(n_30910), .D(n_32301), 
		.Z(n_135778861));
	notech_nand2 i_108163400(.A(n_3825), .B(n_56649), .Z(n_135878862));
	notech_ao4 i_12664328(.A(n_3594), .B(n_60926), .C(n_3833), .D(n_32304), 
		.Z(n_136078864));
	notech_and2 i_110063382(.A(n_56662), .B(n_26837), .Z(n_136578869));
	notech_and4 i_110263380(.A(n_62868), .B(n_56994), .C(n_30931), .D(n_26849
		), .Z(n_136678870));
	notech_or4 i_56163909(.A(n_62864), .B(n_284480345), .C(n_60926), .D(\nbus_11307[1] 
		), .Z(n_137178875));
	notech_or2 i_55863912(.A(n_57982), .B(\nbus_11358[1] ), .Z(n_137478878)
		);
	notech_or4 i_55563915(.A(n_59275), .B(n_59355), .C(n_32356), .D(n_59992)
		, .Z(n_137778881));
	notech_or4 i_57263898(.A(n_62864), .B(n_284480345), .C(n_60926), .D(\nbus_11307[4] 
		), .Z(n_138278886));
	notech_or2 i_56963901(.A(n_57982), .B(\nbus_11358[4] ), .Z(n_138578889)
		);
	notech_or4 i_56663904(.A(n_59275), .B(n_59355), .C(n_32356), .D(n_5723),
		 .Z(n_138878892));
	notech_or4 i_60663866(.A(n_62830), .B(n_303873518), .C(n_60926), .D(n_57542
		), .Z(n_139378897));
	notech_or4 i_60363869(.A(n_58133), .B(n_26906), .C(n_56423), .D(\nbus_11358[1] 
		), .Z(n_139678900));
	notech_or4 i_60063872(.A(n_56822), .B(n_56983), .C(n_56498), .D(n_59992)
		, .Z(n_139978903));
	notech_or4 i_61763855(.A(n_62864), .B(n_303873518), .C(n_60926), .D(\nbus_11307[4] 
		), .Z(n_140478908));
	notech_or4 i_61463858(.A(n_58133), .B(n_26906), .C(n_56423), .D(\nbus_11358[4] 
		), .Z(n_140778911));
	notech_or2 i_61163861(.A(n_304273522), .B(n_5723), .Z(n_141078914));
	notech_nao3 i_62863844(.A(opc[9]), .B(n_62782), .C(n_181879322), .Z(n_141178915
		));
	notech_or2 i_62763845(.A(n_60016), .B(n_181779321), .Z(n_141478918));
	notech_nao3 i_62263850(.A(n_318891635), .B(n_318791636), .C(n_58106), .Z
		(n_141978923));
	notech_or4 i_63763835(.A(n_62864), .B(n_26804), .C(n_62782), .D(n_56019)
		, .Z(n_142478928));
	notech_nao3 i_63463838(.A(n_318791636), .B(n_56925), .C(n_253640554), .Z
		(n_142778931));
	notech_or4 i_63163841(.A(n_58806), .B(n_58162), .C(nbus_11295[1]), .D(n_60926
		), .Z(n_143078934));
	notech_or4 i_66363809(.A(n_62860), .B(n_26804), .C(n_62782), .D(n_56055)
		, .Z(n_143578939));
	notech_or2 i_66063812(.A(n_253740555), .B(n_56914), .Z(n_143878942));
	notech_or4 i_65763815(.A(n_58806), .B(n_58162), .C(nbus_11295[4]), .D(n_60928
		), .Z(n_144178945));
	notech_or4 i_67463798(.A(n_58132), .B(n_58477), .C(n_60016), .D(n_56909)
		, .Z(n_144278946));
	notech_nand3 i_67363799(.A(n_26825), .B(n_26824), .C(\opa_12[9] ), .Z(n_144578949
		));
	notech_or4 i_66863804(.A(n_62854), .B(n_62782), .C(n_56127), .D(n_58477)
		, .Z(n_145078954));
	notech_or4 i_73763736(.A(n_62854), .B(n_247579976), .C(n_60928), .D(\nbus_11307[4] 
		), .Z(n_145578959));
	notech_or2 i_73463739(.A(n_57154), .B(\nbus_11358[4] ), .Z(n_145878962)
		);
	notech_or2 i_73163742(.A(n_147271952), .B(n_5723), .Z(n_146178965));
	notech_or4 i_75763716(.A(n_58817), .B(n_26816), .C(n_28125), .D(n_60928)
		, .Z(n_146678970));
	notech_nand3 i_75463719(.A(n_32304), .B(n_58078), .C(opd[1]), .Z(n_146978973
		));
	notech_or4 i_75163722(.A(n_54709), .B(n_60024), .C(n_56443), .D(n_26816)
		, .Z(n_147278976));
	notech_or4 i_76863705(.A(n_58817), .B(n_26816), .C(n_28128), .D(n_60931)
		, .Z(n_147778981));
	notech_nand3 i_76563708(.A(n_32304), .B(n_58078), .C(opd[4]), .Z(n_148078984
		));
	notech_or2 i_76263711(.A(n_5743), .B(n_301180512), .Z(n_148378987));
	notech_nao3 i_78063693(.A(opc[9]), .B(n_62782), .C(n_323080731), .Z(n_148478988
		));
	notech_or2 i_77963694(.A(n_60016), .B(n_228579786), .Z(n_148778991));
	notech_nand2 i_77663697(.A(opb[9]), .B(n_57179), .Z(n_149078994));
	notech_or2 i_77363700(.A(n_56662), .B(n_58106), .Z(n_149378997));
	notech_or2 i_78863685(.A(n_58044), .B(n_56028), .Z(n_149478998));
	notech_nand3 i_78163692(.A(n_58632), .B(opa[0]), .C(n_131878822), .Z(n_149979003
		));
	notech_nand2 i_78263691(.A(opc[0]), .B(n_131978823), .Z(n_150079004));
	notech_or2 i_78363690(.A(n_58488), .B(n_132078824), .Z(n_150179005));
	notech_or4 i_80363671(.A(n_62860), .B(n_62782), .C(n_56019), .D(n_58488)
		, .Z(n_150279006));
	notech_or4 i_80263672(.A(n_58087), .B(n_58488), .C(n_60024), .D(n_56452)
		, .Z(n_150579009));
	notech_or2 i_79963675(.A(n_253640554), .B(n_56636), .Z(n_150879012));
	notech_nand3 i_79563678(.A(n_26829), .B(n_26808), .C(\opa_12[1] ), .Z(n_151179015
		));
	notech_or4 i_81563659(.A(n_62840), .B(n_62782), .C(n_56055), .D(n_58488)
		, .Z(n_151279016));
	notech_or2 i_81463660(.A(n_5743), .B(n_57470), .Z(n_151579019));
	notech_or2 i_81163663(.A(n_253740555), .B(n_56636), .Z(n_151879022));
	notech_nand3 i_80863666(.A(n_26829), .B(n_26808), .C(\opa_12[4] ), .Z(n_152179025
		));
	notech_or4 i_84763628(.A(n_58087), .B(n_54678), .C(n_60010), .D(n_56452)
		, .Z(n_152279026));
	notech_nao3 i_84663629(.A(n_26829), .B(\opa_12[15] ), .C(n_54678), .Z(n_152579029
		));
	notech_or2 i_84163634(.A(n_250240520), .B(\nbus_11358[15] ), .Z(n_153079034
		));
	notech_nand3 i_31012(.A(n_56925), .B(n_318791636), .C(n_58078), .Z(n_153179035
		));
	notech_or4 i_9264361(.A(n_57026), .B(n_56863), .C(n_29653), .D(n_58162),
		 .Z(n_153279036));
	notech_nand2 i_8864365(.A(n_58806), .B(n_26843), .Z(n_153379037));
	notech_nao3 i_8964364(.A(n_56903), .B(n_26790), .C(n_58162), .Z(n_153479038
		));
	notech_or4 i_12364331(.A(n_32326), .B(n_32339), .C(n_26804), .D(n_58132)
		, .Z(n_153579039));
	notech_or2 i_11164342(.A(n_26804), .B(n_58422), .Z(n_153679040));
	notech_nao3 i_30766(.A(n_32386), .B(n_32299), .C(n_56822), .Z(n_153779041
		));
	notech_nand2 i_11364340(.A(n_26827), .B(n_58487), .Z(n_153879042));
	notech_or4 i_6164392(.A(n_54727), .B(n_57088), .C(n_29652), .D(n_58488),
		 .Z(n_153979043));
	notech_nand2 i_7964374(.A(n_26829), .B(n_26808), .Z(n_154079044));
	notech_or2 i_38869(.A(n_131778821), .B(n_3922), .Z(n_154179045));
	notech_or4 i_38871(.A(instrc[124]), .B(n_29663), .C(n_26885), .D(n_3922)
		, .Z(n_154279046));
	notech_nand3 i_38874(.A(n_30931), .B(n_26898), .C(n_131678820), .Z(n_154379047
		));
	notech_ao4 i_101463466(.A(n_26883), .B(n_134178845), .C(n_134278846), .D
		(n_26733), .Z(n_154679050));
	notech_or2 i_101563465(.A(n_131578819), .B(n_344880949), .Z(n_154779051)
		);
	notech_or2 i_101663464(.A(n_26735), .B(n_344580946), .Z(n_154879052));
	notech_or2 i_101363467(.A(n_133578839), .B(n_340380904), .Z(n_155179055)
		);
	notech_or4 i_100863472(.A(instrc[116]), .B(n_57088), .C(n_345480955), .D
		(n_29653), .Z(n_155279056));
	notech_or4 i_100963471(.A(n_345880959), .B(instrc[98]), .C(n_314663413),
		 .D(instrc[96]), .Z(n_155379057));
	notech_and4 i_101063470(.A(n_29635), .B(n_29665), .C(instrc[103]), .D(n_29967
		), .Z(n_155479058));
	notech_or2 i_103263448(.A(n_345680957), .B(n_340380904), .Z(n_155979063)
		);
	notech_ao3 i_102963451(.A(n_29631), .B(instrc[91]), .C(n_75738777), .Z(n_156279066
		));
	notech_and4 i_102463456(.A(n_30350), .B(n_29635), .C(n_29665), .D(instrc
		[103]), .Z(n_156379067));
	notech_or4 i_102563455(.A(n_57078), .B(n_57051), .C(n_29653), .D(n_345480955
		), .Z(n_156479068));
	notech_or4 i_102663454(.A(instrc[93]), .B(n_346280963), .C(instrc[94]), 
		.D(n_26972), .Z(n_156579069));
	notech_nand3 i_107663405(.A(n_319091633), .B(n_56925), .C(n_26836), .Z(n_156879072
		));
	notech_or2 i_107363408(.A(n_251040528), .B(n_54765), .Z(n_157179075));
	notech_ao3 i_107063411(.A(instrc[89]), .B(instrc[91]), .C(n_75738777), .Z
		(n_157479078));
	notech_and4 i_106663415(.A(n_30357), .B(n_29666), .C(instrc[93]), .D(n_26847
		), .Z(n_157579079));
	notech_and4 i_106763414(.A(instrc[119]), .B(n_57078), .C(instrc[116]), .D
		(n_26859), .Z(n_157679080));
	notech_ao3 i_106463417(.A(instrc[96]), .B(instrc[99]), .C(n_77438794), .Z
		(n_157779081));
	notech_and4 i_106563416(.A(n_62868), .B(n_76638786), .C(n_134978853), .D
		(n_30322), .Z(n_157879082));
	notech_ao3 i_109863384(.A(n_318891635), .B(n_26836), .C(n_59275), .Z(n_158179085
		));
	notech_or2 i_109263389(.A(n_58817), .B(n_136078864), .Z(n_158279086));
	notech_ao4 i_109363388(.A(n_136578869), .B(n_26840), .C(n_323480735), .D
		(n_161179115), .Z(n_158379087));
	notech_ao4 i_109463387(.A(n_136678870), .B(n_26737), .C(n_3822), .D(n_26738
		), .Z(n_158479088));
	notech_or4 i_108963392(.A(n_29954), .B(instrc[93]), .C(n_29666), .D(n_346280963
		), .Z(n_158579089));
	notech_or4 i_109063391(.A(n_29667), .B(n_314663413), .C(n_345880959), .D
		(instrc[96]), .Z(n_158679090));
	notech_or4 i_109163390(.A(n_346080961), .B(n_30306), .C(instrc[88]), .D(n_314663413
		), .Z(n_158779091));
	notech_or4 i_108763394(.A(instrc[116]), .B(n_29653), .C(n_57078), .D(n_26971
		), .Z(n_158879092));
	notech_or4 i_108863393(.A(n_26968), .B(n_3908), .C(instrc[124]), .D(n_29663
		), .Z(n_158979093));
	notech_or4 i_108563396(.A(n_29665), .B(n_29637), .C(instrc[101]), .D(n_26899
		), .Z(n_159079094));
	notech_or4 i_108663395(.A(instrc[125]), .B(n_26838), .C(instrc[124]), .D
		(n_340480905), .Z(n_159179095));
	notech_and2 i_7664377(.A(n_57051), .B(instrc[119]), .Z(n_159379097));
	notech_nand2 i_205264448(.A(n_29632), .B(instrc[127]), .Z(n_160079104)
		);
	notech_and4 i_184262661(.A(n_158979093), .B(n_159179095), .C(n_158879092
		), .D(n_159079094), .Z(n_160379107));
	notech_and4 i_184362660(.A(n_158579089), .B(n_158779091), .C(n_160379107
		), .D(n_158679090), .Z(n_160979113));
	notech_or2 i_864442(.A(n_136678870), .B(n_26737), .Z(n_161179115));
	notech_ao4 i_184462659(.A(n_56946), .B(n_3695), .C(n_32304), .D(n_3915),
		 .Z(n_161279116));
	notech_nao3 i_183662667(.A(n_158279086), .B(n_26739), .C(n_158479088), .Z
		(n_161479118));
	notech_ao4 i_183362670(.A(n_345980960), .B(n_26735), .C(n_131578819), .D
		(n_346180962), .Z(n_161579119));
	notech_or4 i_6064393(.A(n_61143), .B(n_60292), .C(n_26900), .D(instrc[98
		]), .Z(n_161879122));
	notech_or4 i_182462679(.A(n_157679080), .B(n_157579079), .C(n_157879082)
		, .D(n_157779081), .Z(n_162579129));
	notech_nand3 i_182762676(.A(instrc[101]), .B(instrc[103]), .C(n_30350), 
		.Z(n_162679130));
	notech_ao4 i_182062683(.A(n_135078854), .B(n_32301), .C(instrc[102]), .D
		(n_162679130), .Z(n_162779131));
	notech_ao4 i_181762686(.A(n_74738767), .B(n_32339), .C(n_74838768), .D(n_30303
		), .Z(n_163079134));
	notech_ao4 i_181562688(.A(n_345680957), .B(n_26885), .C(n_57322), .D(n_74438764
		), .Z(n_163279136));
	notech_and4 i_181962684(.A(n_163279136), .B(n_163079134), .C(n_156879072
		), .D(n_157179075), .Z(n_163479138));
	notech_or4 i_177462729(.A(n_314663413), .B(n_29638), .C(instrc[93]), .D(instrc
		[94]), .Z(n_163679140));
	notech_nao3 i_177162732(.A(n_156479068), .B(n_156579069), .C(n_156379067
		), .Z(n_164079144));
	notech_nao3 i_177362730(.A(n_62868), .B(n_57501), .C(n_340380904), .Z(n_164179145
		));
	notech_ao4 i_176862735(.A(n_134578849), .B(n_134478848), .C(n_58806), .D
		(n_134378847), .Z(n_164279146));
	notech_ao4 i_176562738(.A(n_56914), .B(n_3829), .C(n_161879122), .D(n_345780958
		), .Z(n_164579149));
	notech_ao4 i_176362740(.A(n_32339), .B(n_344580946), .C(n_344880949), .D
		(n_30303), .Z(n_164779151));
	notech_and4 i_176762736(.A(n_318091643), .B(n_164779151), .C(n_155979063
		), .D(n_164579149), .Z(n_164979153));
	notech_ao3 i_175662747(.A(n_155279056), .B(n_155379057), .C(n_155479058)
		, .Z(n_165479158));
	notech_ao4 i_175362750(.A(n_54814), .B(n_133478838), .C(n_163679140), .D
		(n_29954), .Z(n_165579159));
	notech_ao4 i_174962754(.A(n_344680947), .B(n_346080961), .C(n_56498), .D
		(n_3829), .Z(n_166179165));
	notech_and4 i_175262751(.A(n_154779051), .B(n_166179165), .C(n_154879052
		), .D(n_26745), .Z(n_166279166));
	notech_ao4 i_156162936(.A(\nbus_11307[15] ), .B(n_26846), .C(n_124271722
		), .D(n_28000), .Z(n_166679170));
	notech_ao4 i_156062937(.A(n_58105), .B(n_56636), .C(n_54678), .D(n_58622
		), .Z(n_166879172));
	notech_ao4 i_155762940(.A(n_298466513), .B(n_57473), .C(nbus_11295[15]),
		 .D(n_26823), .Z(n_167079174));
	notech_and4 i_155962938(.A(n_128171761), .B(n_167079174), .C(n_152279026
		), .D(n_152579029), .Z(n_167379177));
	notech_ao4 i_153662961(.A(n_124171721), .B(n_291663183), .C(n_291763184)
		, .D(n_123971719), .Z(n_167479178));
	notech_ao4 i_153462963(.A(n_291863185), .B(n_153979043), .C(n_123871718)
		, .D(n_57574), .Z(n_167679180));
	notech_and4 i_153862959(.A(n_167679180), .B(n_167479178), .C(n_151879022
		), .D(n_152179025), .Z(n_167879182));
	notech_ao4 i_153162966(.A(n_58044), .B(\nbus_11358[4] ), .C(n_56529), .D
		(n_291563182), .Z(n_167979183));
	notech_and4 i_153362964(.A(n_181462097), .B(n_167979183), .C(n_151279016
		), .D(n_151579019), .Z(n_168279186));
	notech_ao4 i_152762970(.A(n_124171721), .B(n_297866507), .C(n_123971719)
		, .D(n_297966508), .Z(n_168379187));
	notech_ao4 i_152562972(.A(n_298066509), .B(n_153979043), .C(n_123871718)
		, .D(n_57542), .Z(n_168579189));
	notech_and4 i_152962968(.A(n_168579189), .B(n_168379187), .C(n_150879012
		), .D(n_151179015), .Z(n_168779191));
	notech_ao4 i_152262975(.A(n_58044), .B(\nbus_11358[1] ), .C(n_56529), .D
		(n_297766506), .Z(n_168879192));
	notech_and4 i_152462973(.A(n_228879789), .B(n_168879192), .C(n_150279006
		), .D(n_150579009), .Z(n_169179195));
	notech_ao4 i_151662981(.A(n_291163178), .B(n_153979043), .C(n_124271722)
		, .D(n_59993), .Z(n_169579199));
	notech_and4 i_151962978(.A(n_169579199), .B(n_150079004), .C(n_149979003
		), .D(n_150179005), .Z(n_169679200));
	notech_ao4 i_151462983(.A(n_291363180), .B(n_124071720), .C(n_123771717)
		, .D(n_59187), .Z(n_169779201));
	notech_ao4 i_151062987(.A(n_143571915), .B(n_27992), .C(n_58479), .D(n_58608
		), .Z(n_170079204));
	notech_ao4 i_150762989(.A(n_57613), .B(n_26856), .C(n_322880729), .D(nbus_11295
		[9]), .Z(n_170279206));
	notech_and4 i_151262985(.A(n_170279206), .B(n_170079204), .C(n_149078994
		), .D(n_149378997), .Z(n_170479208));
	notech_ao4 i_150462992(.A(n_322980730), .B(n_56127), .C(n_291963186), .D
		(n_322780728), .Z(n_170579209));
	notech_and4 i_150662990(.A(n_200065529), .B(n_170579209), .C(n_148778991
		), .D(n_148478988), .Z(n_170879212));
	notech_ao4 i_150062996(.A(n_153879042), .B(n_56055), .C(n_123671716), .D
		(n_57574), .Z(n_170979213));
	notech_ao4 i_149862998(.A(n_291463181), .B(n_26816), .C(n_57573), .D(n_56064
		), .Z(n_171179215));
	notech_and4 i_150262994(.A(n_171179215), .B(n_170979213), .C(n_148078984
		), .D(n_148378987), .Z(n_171379217));
	notech_ao4 i_149363001(.A(n_291563182), .B(n_26807), .C(n_143571915), .D
		(n_5723), .Z(n_171479218));
	notech_ao4 i_149163003(.A(n_291663183), .B(n_229479795), .C(n_291763184)
		, .D(n_229379794), .Z(n_171679220));
	notech_and4 i_149762999(.A(n_181462097), .B(n_171679220), .C(n_171479218
		), .D(n_147778981), .Z(n_171879222));
	notech_ao4 i_148863006(.A(n_153879042), .B(n_56019), .C(n_123671716), .D
		(n_57542), .Z(n_171979223));
	notech_ao4 i_148663008(.A(n_297666505), .B(n_26816), .C(n_57573), .D(n_56010
		), .Z(n_172179225));
	notech_and4 i_149063004(.A(n_172179225), .B(n_171979223), .C(n_146978973
		), .D(n_147278976), .Z(n_172379227));
	notech_ao4 i_148363011(.A(n_26807), .B(n_297766506), .C(n_143571915), .D
		(n_59992), .Z(n_172479228));
	notech_ao4 i_148163013(.A(n_297866507), .B(n_229479795), .C(n_297966508)
		, .D(n_229379794), .Z(n_172679230));
	notech_and4 i_148563009(.A(n_228879789), .B(n_172679230), .C(n_146678970
		), .D(n_172479228), .Z(n_172879232));
	notech_ao4 i_146963024(.A(n_147171951), .B(n_27986), .C(n_58486), .D(n_291463181
		), .Z(n_172979233));
	notech_ao4 i_146763026(.A(n_147371953), .B(n_57574), .C(n_291563182), .D
		(n_266380164), .Z(n_173179235));
	notech_and4 i_147163022(.A(n_173179235), .B(n_172979233), .C(n_145878962
		), .D(n_146178965), .Z(n_173379237));
	notech_ao4 i_146463029(.A(n_291763184), .B(n_247479975), .C(n_57141), .D
		(n_291863185), .Z(n_173479238));
	notech_ao4 i_146263031(.A(n_247679977), .B(n_56055), .C(n_5743), .D(n_57084
		), .Z(n_173679240));
	notech_and4 i_146663027(.A(n_181462097), .B(n_173679240), .C(n_173479238
		), .D(n_145578959), .Z(n_173879242));
	notech_ao4 i_141363079(.A(n_189962171), .B(n_181979323), .C(n_56914), .D
		(n_252740545), .Z(n_173979243));
	notech_ao4 i_141263080(.A(n_57613), .B(n_26854), .C(n_56356), .D(nbus_11295
		[9]), .Z(n_174179245));
	notech_ao4 i_140963083(.A(n_291963186), .B(n_322580726), .C(\nbus_11358[9] 
		), .D(n_26853), .Z(n_174379247));
	notech_and4 i_141163081(.A(n_200065529), .B(n_144278946), .C(n_174379247
		), .D(n_144578949), .Z(n_174679250));
	notech_ao4 i_140563087(.A(n_56055), .B(n_153679040), .C(n_5743), .D(n_153579039
		), .Z(n_174779251));
	notech_ao4 i_140363089(.A(n_291663183), .B(n_153379037), .C(n_153479038)
		, .D(n_57574), .Z(n_174979253));
	notech_and4 i_140763085(.A(n_174979253), .B(n_174779251), .C(n_143878942
		), .D(n_144178945), .Z(n_175179255));
	notech_ao4 i_140063092(.A(n_291563182), .B(n_58162), .C(n_58047), .D(n_56064
		), .Z(n_175279256));
	notech_ao4 i_139863094(.A(n_56356), .B(nbus_11295[4]), .C(n_291863185), 
		.D(n_257980080), .Z(n_175479258));
	notech_and4 i_140263090(.A(n_181462097), .B(n_175479258), .C(n_175279256
		), .D(n_143578939), .Z(n_175679260));
	notech_ao4 i_138263109(.A(n_153679040), .B(n_56019), .C(n_60024), .D(n_153579039
		), .Z(n_175779261));
	notech_ao4 i_138063111(.A(n_297866507), .B(n_153379037), .C(n_153479038)
		, .D(n_57542), .Z(n_175979263));
	notech_and4 i_138563107(.A(n_175979263), .B(n_175779261), .C(n_142778931
		), .D(n_143078934), .Z(n_176179265));
	notech_ao4 i_137763114(.A(n_297766506), .B(n_58162), .C(n_58047), .D(n_56010
		), .Z(n_176279266));
	notech_ao4 i_137563116(.A(n_56356), .B(nbus_11295[1]), .C(n_298066509), 
		.D(n_257980080), .Z(n_176479268));
	notech_and4 i_137963112(.A(n_228879789), .B(n_176479268), .C(n_176279266
		), .D(n_142478928), .Z(n_176679270));
	notech_ao4 i_137263119(.A(n_304273522), .B(n_27992), .C(n_58608), .D(n_58481
		), .Z(n_176779271));
	notech_ao4 i_137163120(.A(n_58052), .B(n_56136), .C(n_57613), .D(n_26851
		), .Z(n_176979273));
	notech_ao4 i_136863123(.A(n_197279473), .B(n_56127), .C(n_291963186), .D
		(n_57765), .Z(n_177179275));
	notech_and4 i_137063121(.A(n_200065529), .B(n_177179275), .C(n_141178915
		), .D(n_141478918), .Z(n_177479278));
	notech_ao4 i_136463127(.A(n_303973519), .B(n_27986), .C(n_58489), .D(n_291463181
		), .Z(n_177579279));
	notech_ao4 i_136263129(.A(n_304473524), .B(n_57574), .C(n_26906), .D(n_291563182
		), .Z(n_177779281));
	notech_and4 i_136663125(.A(n_177779281), .B(n_177579279), .C(n_140778911
		), .D(n_141078914), .Z(n_177979283));
	notech_ao4 i_135963132(.A(n_303773517), .B(n_291763184), .C(n_57923), .D
		(n_291863185), .Z(n_178079284));
	notech_ao4 i_135763134(.A(n_56055), .B(n_284980350), .C(n_5743), .D(n_285080351
		), .Z(n_178279286));
	notech_and4 i_136163130(.A(n_181462097), .B(n_178279286), .C(n_178079284
		), .D(n_140478908), .Z(n_178479288));
	notech_ao4 i_135463137(.A(n_303973519), .B(n_59241), .C(n_58489), .D(n_297666505
		), .Z(n_178579289));
	notech_ao4 i_135263139(.A(n_304473524), .B(n_57542), .C(n_26906), .D(n_297766506
		), .Z(n_178779291));
	notech_and4 i_135663135(.A(n_178779291), .B(n_178579289), .C(n_139678900
		), .D(n_139978903), .Z(n_178979293));
	notech_ao4 i_134963142(.A(n_303773517), .B(n_297966508), .C(n_57923), .D
		(n_298066509), .Z(n_179079294));
	notech_ao4 i_134763144(.A(n_284980350), .B(n_56019), .C(n_60024), .D(n_285080351
		), .Z(n_179279296));
	notech_and4 i_135163140(.A(n_228879789), .B(n_179279296), .C(n_139378897
		), .D(n_179079294), .Z(n_179479298));
	notech_ao4 i_131963172(.A(n_284580346), .B(n_27986), .C(n_291463181), .D
		(n_26812), .Z(n_179579299));
	notech_ao4 i_131663174(.A(n_284380344), .B(n_57574), .C(n_291563182), .D
		(n_26852), .Z(n_179779301));
	notech_and4 i_132163170(.A(n_179779301), .B(n_138878892), .C(n_179579299
		), .D(n_138578889), .Z(n_179979303));
	notech_ao4 i_131363177(.A(n_291763184), .B(n_284680347), .C(n_291863185)
		, .D(n_57915), .Z(n_180079304));
	notech_ao4 i_131163179(.A(n_56055), .B(n_284780348), .C(n_5743), .D(n_284880349
		), .Z(n_180279306));
	notech_and4 i_131563175(.A(n_180279306), .B(n_180079304), .C(n_181462097
		), .D(n_138278886), .Z(n_180479308));
	notech_ao4 i_130863182(.A(n_284580346), .B(n_59241), .C(n_297666505), .D
		(n_26812), .Z(n_180579309));
	notech_ao4 i_130663184(.A(n_284380344), .B(n_57542), .C(n_297766506), .D
		(n_26852), .Z(n_180779311));
	notech_and4 i_131063180(.A(n_180779311), .B(n_180579309), .C(n_137478878
		), .D(n_137778881), .Z(n_180979313));
	notech_ao4 i_130363187(.A(n_297966508), .B(n_284680347), .C(n_298066509)
		, .D(n_57915), .Z(n_181079314));
	notech_ao4 i_130163189(.A(n_284780348), .B(n_56019), .C(n_60024), .D(n_284880349
		), .Z(n_181279316));
	notech_and4 i_130563185(.A(n_181279316), .B(n_137178875), .C(n_181079314
		), .D(n_228879789), .Z(n_181479318));
	notech_nao3 i_180261731(.A(n_56423), .B(n_26821), .C(n_58133), .Z(n_181679320
		));
	notech_or4 i_180361730(.A(n_32326), .B(n_58133), .C(n_26735), .D(n_58481
		), .Z(n_181779321));
	notech_and2 i_151161784(.A(n_57923), .B(n_182079324), .Z(n_181879322));
	notech_and2 i_149664482(.A(n_257980080), .B(n_133078834), .Z(n_181979323
		));
	notech_or2 i_121060581(.A(n_54814), .B(n_182179325), .Z(n_182079324));
	notech_and2 i_561718(.A(n_58505), .B(n_58497), .Z(n_182179325));
	notech_nand3 i_123060563(.A(n_58172), .B(n_30945), .C(n_190062172), .Z(n_182279326
		));
	notech_or4 i_123260561(.A(n_59387), .B(n_4011), .C(n_29178), .D(n_27198)
		, .Z(n_182379327));
	notech_nao3 i_5361675(.A(tsc[13]), .B(n_55820), .C(n_59469), .Z(n_182479328
		));
	notech_or4 i_5261676(.A(n_60931), .B(n_28139), .C(n_26942), .D(n_23512),
		 .Z(n_182779331));
	notech_nand2 i_4961679(.A(opb[13]), .B(n_58097), .Z(n_183079334));
	notech_nao3 i_4661682(.A(n_62826), .B(opc[13]), .C(n_312970140), .Z(n_183379337
		));
	notech_ao3 i_9561633(.A(tsc[30]), .B(n_55820), .C(n_59469), .Z(n_183479338
		));
	notech_or2 i_9461634(.A(n_59124), .B(nbus_11295[30]), .Z(n_183779341));
	notech_or4 i_9161637(.A(n_56822), .B(n_56946), .C(n_56579), .D(n_28015),
		 .Z(n_184079344));
	notech_or4 i_8861640(.A(n_317591648), .B(n_60841), .C(n_54974), .D(\nbus_11358[30] 
		), .Z(n_184379347));
	notech_nao3 i_28561443(.A(tsc[62]), .B(n_55820), .C(n_59469), .Z(n_184679350
		));
	notech_or4 i_28261446(.A(n_56822), .B(n_56946), .C(n_56527), .D(n_28015)
		, .Z(n_184979353));
	notech_or2 i_27961449(.A(n_149428771), .B(\nbus_11358[30] ), .Z(n_185279356
		));
	notech_or4 i_31561414(.A(n_55581), .B(n_298466513), .C(n_27119), .D(n_26054
		), .Z(n_185379357));
	notech_or4 i_31461415(.A(n_62856), .B(n_62806), .C(n_56266), .D(n_26054)
		, .Z(n_185679360));
	notech_nand2 i_30861420(.A(n_302191802), .B(opa[15]), .Z(n_186179365));
	notech_or4 i_32361406(.A(n_3845), .B(n_26767), .C(n_60928), .D(nbus_11295
		[30]), .Z(n_186479368));
	notech_or2 i_31861411(.A(n_3878), .B(\nbus_11365[30] ), .Z(n_186979373)
		);
	notech_or4 i_88360874(.A(n_62856), .B(\opcode[2] ), .C(n_29592), .D(n_58481
		), .Z(n_187079374));
	notech_nand2 i_88260875(.A(opd[13]), .B(n_58377), .Z(n_187379377));
	notech_or4 i_87960878(.A(n_54814), .B(n_60928), .C(n_28139), .D(n_58481)
		, .Z(n_187679380));
	notech_nao3 i_87660881(.A(n_54814), .B(n_26821), .C(n_31576), .Z(n_187979383
		));
	notech_or4 i_90360855(.A(n_62858), .B(n_62788), .C(n_56266), .D(n_58481)
		, .Z(n_188079384));
	notech_or4 i_90260856(.A(n_56822), .B(n_56979), .C(n_56498), .D(n_28000)
		, .Z(n_188379387));
	notech_nand3 i_89760861(.A(n_26813), .B(n_26821), .C(\opa_12[15] ), .Z(n_188879392
		));
	notech_or2 i_93160829(.A(n_56356), .B(nbus_11295[13]), .Z(n_189379397)
		);
	notech_nand2 i_92860832(.A(opb[13]), .B(n_58050), .Z(n_189779400));
	notech_or4 i_92560835(.A(n_58477), .B(n_58132), .C(n_32325), .D(n_29592)
		, .Z(n_190079403));
	notech_or2 i_95560806(.A(n_56356), .B(nbus_11295[15]), .Z(n_190179404)
		);
	notech_or4 i_95460807(.A(n_58806), .B(n_28141), .C(n_60928), .D(n_58477)
		, .Z(n_190479407));
	notech_nand2 i_95160810(.A(opb[15]), .B(n_58050), .Z(n_190779410));
	notech_nand2 i_94860813(.A(opa[15]), .B(n_58051), .Z(n_191079413));
	notech_nao3 i_102460740(.A(n_54765), .B(n_26884), .C(n_31576), .Z(n_191179414
		));
	notech_or4 i_102360741(.A(n_54765), .B(n_58478), .C(n_60928), .D(n_28139
		), .Z(n_191479417));
	notech_or2 i_102060744(.A(n_57181), .B(\nbus_11358[13] ), .Z(n_191779420
		));
	notech_or4 i_101760747(.A(n_54756), .B(n_58478), .C(n_32331), .D(n_56239
		), .Z(n_192079423));
	notech_or4 i_104360721(.A(n_54765), .B(n_58478), .C(n_28141), .D(n_60928
		), .Z(n_192179424));
	notech_or4 i_104260722(.A(n_62860), .B(n_62788), .C(n_56266), .D(n_58478
		), .Z(n_192479427));
	notech_nand2 i_103760727(.A(n_313170142), .B(opa[15]), .Z(n_192979432)
		);
	notech_or4 i_108560695(.A(n_58817), .B(n_58495), .C(n_60928), .D(nbus_11295
		[13]), .Z(n_193479437));
	notech_nand2 i_108260698(.A(opb[13]), .B(n_57179), .Z(n_193779440));
	notech_or4 i_107760701(.A(n_54709), .B(n_58479), .C(n_32332), .D(n_56239
		), .Z(n_194079443));
	notech_or4 i_110960672(.A(n_58817), .B(n_58495), .C(n_60928), .D(nbus_11295
		[15]), .Z(n_194179444));
	notech_or4 i_110860673(.A(n_54718), .B(n_28141), .C(n_60928), .D(n_58479
		), .Z(n_194479447));
	notech_nand2 i_110560676(.A(opb[15]), .B(n_57179), .Z(n_194779450));
	notech_nand2 i_110260679(.A(opa[15]), .B(n_57180), .Z(n_195079453));
	notech_or4 i_113760646(.A(n_54678), .B(n_58815), .C(n_59419), .D(n_56239
		), .Z(n_195179454));
	notech_or4 i_113660647(.A(n_58087), .B(n_54678), .C(n_302091803), .D(n_56452
		), .Z(n_195479457));
	notech_nand2 i_113360650(.A(opc[13]), .B(n_57808), .Z(n_195779460));
	notech_or4 i_113060653(.A(n_62856), .B(n_54678), .C(n_62788), .D(n_56239
		), .Z(n_196079463));
	notech_or2 i_118360608(.A(n_57726), .B(n_28156), .Z(n_196179464));
	notech_or4 i_118260609(.A(n_56863), .B(n_54727), .C(n_30809), .D(n_58504
		), .Z(n_196579467));
	notech_or2 i_117760614(.A(n_57865), .B(\nbus_11358[30] ), .Z(n_197179472
		));
	notech_nand2 i_31241(.A(n_26813), .B(n_26821), .Z(n_197279473));
	notech_ao4 i_223059608(.A(n_58138), .B(n_302991794), .C(n_57867), .D(\nbus_11365[30] 
		), .Z(n_197579476));
	notech_ao4 i_222959609(.A(n_305624320), .B(n_303091793), .C(n_26937), .D
		(n_29591), .Z(n_197779478));
	notech_ao4 i_222659612(.A(n_58008), .B(n_32252), .C(n_58423), .D(n_28015
		), .Z(n_197979480));
	notech_and4 i_222859610(.A(n_197979480), .B(n_26604), .C(n_196179464), .D
		(n_196579467), .Z(n_198279483));
	notech_ao4 i_219959639(.A(n_184868865), .B(n_56239), .C(n_94935745), .D(n_56636
		), .Z(n_198379484));
	notech_ao4 i_219759641(.A(n_57809), .B(\nbus_11307[13] ), .C(n_58376), .D
		(n_27998), .Z(n_198579486));
	notech_and4 i_220159637(.A(n_198579486), .B(n_198379484), .C(n_195779460
		), .D(n_196079463), .Z(n_198779488));
	notech_ao4 i_219459644(.A(n_31560), .B(n_57473), .C(n_57807), .D(\nbus_11358[13] 
		), .Z(n_198879489));
	notech_and4 i_219659642(.A(n_93835734), .B(n_198879489), .C(n_195179454)
		, .D(n_195479457), .Z(n_199179492));
	notech_ao4 i_217659662(.A(n_58105), .B(n_56662), .C(n_323080731), .D(n_111064639
		), .Z(n_199279493));
	notech_ao4 i_217459664(.A(n_60010), .B(n_228579786), .C(n_56266), .D(n_322980730
		), .Z(n_199479495));
	notech_and4 i_217859660(.A(n_199479495), .B(n_199279493), .C(n_194779450
		), .D(n_195079453), .Z(n_199679497));
	notech_ao4 i_217159667(.A(n_58479), .B(n_58622), .C(n_143571915), .D(n_28000
		), .Z(n_199779498));
	notech_and4 i_217359665(.A(n_128171761), .B(n_194479447), .C(n_199779498
		), .D(n_194179444), .Z(n_200079501));
	notech_ao4 i_215759681(.A(n_30109), .B(n_323080731), .C(n_94935745), .D(n_56662
		), .Z(n_200179502));
	notech_ao4 i_215559683(.A(\nbus_11307[13] ), .B(n_26856), .C(n_302091803
		), .D(n_228579786), .Z(n_200379504));
	notech_and4 i_215959679(.A(n_200379504), .B(n_200179502), .C(n_193779440
		), .D(n_194079443), .Z(n_200579506));
	notech_ao4 i_215259686(.A(n_58375), .B(n_27998), .C(n_31540), .D(n_58479
		), .Z(n_200679507));
	notech_ao4 i_215059688(.A(n_31576), .B(n_228779788), .C(n_31560), .D(n_322780728
		), .Z(n_200879509));
	notech_and4 i_215459684(.A(n_93835734), .B(n_200879509), .C(n_200679507)
		, .D(n_193479437), .Z(n_201079511));
	notech_ao4 i_213259706(.A(n_56649), .B(n_58105), .C(n_313270143), .D(n_111064639
		), .Z(n_201179512));
	notech_ao4 i_213159707(.A(n_57025), .B(n_60010), .C(n_319970210), .D(n_56266
		), .Z(n_201379514));
	notech_ao4 i_212859710(.A(n_147271952), .B(n_28000), .C(n_57181), .D(\nbus_11358[15] 
		), .Z(n_201579516));
	notech_and4 i_213059708(.A(n_128171761), .B(n_201579516), .C(n_192179424
		), .D(n_192479427), .Z(n_201879519));
	notech_ao4 i_211559723(.A(n_313270143), .B(n_30109), .C(n_94935745), .D(n_56649
		), .Z(n_201979520));
	notech_ao4 i_211359725(.A(n_26607), .B(\nbus_11307[13] ), .C(n_184368860
		), .D(n_302091803), .Z(n_202179522));
	notech_and4 i_211759721(.A(n_202179522), .B(n_192079423), .C(n_201979520
		), .D(n_191779420), .Z(n_202379524));
	notech_ao4 i_211059728(.A(n_58374), .B(n_27998), .C(n_54736), .D(n_31540
		), .Z(n_202479525));
	notech_and4 i_211259726(.A(n_93835734), .B(n_191479417), .C(n_202479525)
		, .D(n_191179414), .Z(n_202779528));
	notech_ao4 i_205659782(.A(n_58105), .B(n_56914), .C(n_111064639), .D(n_181979323
		), .Z(n_202879529));
	notech_ao4 i_205459784(.A(n_60010), .B(n_228479785), .C(n_56266), .D(n_322680727
		), .Z(n_203079531));
	notech_and4 i_205859780(.A(n_203079531), .B(n_202879529), .C(n_190779410
		), .D(n_191079413), .Z(n_203279533));
	notech_ao4 i_205159787(.A(n_58477), .B(n_58622), .C(n_153779041), .D(n_28000
		), .Z(n_203379534));
	notech_and4 i_205359785(.A(n_128171761), .B(n_190479407), .C(n_203379534
		), .D(n_190179404), .Z(n_203679537));
	notech_ao4 i_203559801(.A(n_30109), .B(n_58041), .C(n_94935745), .D(n_56914
		), .Z(n_203779538));
	notech_ao4 i_203359803(.A(\nbus_11307[13] ), .B(n_26854), .C(n_302091803
		), .D(n_228479785), .Z(n_203979540));
	notech_and4 i_203759799(.A(n_203979540), .B(n_190079403), .C(n_203779538
		), .D(n_189779400), .Z(n_204179542));
	notech_ao4 i_203059806(.A(n_58372), .B(n_27998), .C(n_31540), .D(n_58477
		), .Z(n_204279543));
	notech_ao4 i_202859808(.A(n_31576), .B(n_228379784), .C(n_31560), .D(n_322580726
		), .Z(n_204479545));
	notech_and4 i_203259804(.A(n_93835734), .B(n_204479545), .C(n_204279543)
		, .D(n_189379397), .Z(n_204679547));
	notech_ao4 i_201059826(.A(n_58105), .B(n_56498), .C(n_111064639), .D(n_181879322
		), .Z(n_204779548));
	notech_ao4 i_200959827(.A(n_58052), .B(n_56275), .C(n_298466513), .D(n_57765
		), .Z(n_204979550));
	notech_ao4 i_200659830(.A(n_60010), .B(n_181779321), .C(\nbus_11307[15] 
		), .D(n_26851), .Z(n_205179552));
	notech_and4 i_200859828(.A(n_128171761), .B(n_205179552), .C(n_188079384
		), .D(n_188379387), .Z(n_205479555));
	notech_ao4 i_199359843(.A(n_181679320), .B(n_56239), .C(n_302091803), .D
		(n_181779321), .Z(n_205579556));
	notech_ao4 i_199159845(.A(n_30109), .B(n_58038), .C(n_94935745), .D(n_56498
		), .Z(n_205779558));
	notech_and4 i_199559841(.A(n_205779558), .B(n_205579556), .C(n_187679380
		), .D(n_187979383), .Z(n_205979560));
	notech_ao4 i_198859848(.A(n_26851), .B(\nbus_11307[13] ), .C(\nbus_11358[13] 
		), .D(n_58052), .Z(n_206079561));
	notech_and4 i_199059846(.A(n_93835734), .B(n_206079561), .C(n_187079374)
		, .D(n_187379377), .Z(n_206379564));
	notech_ao4 i_150660297(.A(n_3837), .B(n_303091793), .C(n_3843), .D(n_30809
		), .Z(n_206479565));
	notech_ao4 i_150560298(.A(n_3877), .B(\nbus_11358[30] ), .C(n_148228759)
		, .D(n_302991794), .Z(n_206679567));
	notech_ao4 i_150260301(.A(n_3857), .B(n_28015), .C(n_26642), .D(n_29591)
		, .Z(n_206879569));
	notech_and4 i_150460299(.A(n_54667), .B(n_206879569), .C(n_26604), .D(n_186479368
		), .Z(n_207179572));
	notech_ao4 i_149860305(.A(n_56601), .B(n_58105), .C(n_111064639), .D(n_210879609
		), .Z(n_207279573));
	notech_ao4 i_149760306(.A(n_60010), .B(n_25875), .C(n_56266), .D(n_322480725
		), .Z(n_207479575));
	notech_ao4 i_149460309(.A(n_147671956), .B(n_28000), .C(n_302291801), .D
		(n_56275), .Z(n_207679577));
	notech_and4 i_149660307(.A(n_207679577), .B(n_128171761), .C(n_185379357
		), .D(n_185679360), .Z(n_207979580));
	notech_ao4 i_147060333(.A(n_149128768), .B(n_302991794), .C(n_149328770)
		, .D(\nbus_11365[30] ), .Z(n_208079581));
	notech_ao4 i_146860335(.A(n_148728764), .B(n_303091793), .C(n_149228769)
		, .D(n_29591), .Z(n_208279583));
	notech_and4 i_147260331(.A(n_208279583), .B(n_208079581), .C(n_184979353
		), .D(n_185279356), .Z(n_208479585));
	notech_ao4 i_146360338(.A(n_310791716), .B(n_30809), .C(n_310891715), .D
		(n_32252), .Z(n_208579586));
	notech_ao4 i_146260339(.A(n_60292), .B(n_28121), .C(n_3867), .D(n_27025)
		, .Z(n_208779588));
	notech_ao4 i_128660511(.A(n_302991794), .B(n_151428791), .C(\nbus_11365[30] 
		), .D(n_311091713), .Z(n_208979590));
	notech_ao4 i_128360513(.A(n_303091793), .B(n_151128788), .C(n_29591), .D
		(n_26696), .Z(n_209179592));
	notech_and4 i_128860509(.A(n_209179592), .B(n_208979590), .C(n_184079344
		), .D(n_184379347), .Z(n_209379594));
	notech_ao4 i_128060516(.A(n_30809), .B(n_311391710), .C(n_32252), .D(n_311491709
		), .Z(n_209479595));
	notech_nand2 i_128160515(.A(n_209479595), .B(n_183779341), .Z(n_209579596
		));
	notech_or2 i_124660549(.A(n_316191662), .B(n_56239), .Z(n_209879599));
	notech_ao4 i_124260552(.A(n_94935745), .B(n_56579), .C(n_23512), .D(n_209879599
		), .Z(n_209979600));
	notech_ao4 i_124060554(.A(n_26819), .B(\nbus_11307[13] ), .C(n_302091803
		), .D(n_316691657), .Z(n_210179602));
	notech_and4 i_124460550(.A(n_210179602), .B(n_209979600), .C(n_183079334
		), .D(n_183379337), .Z(n_210379604));
	notech_ao4 i_123660557(.A(n_151028787), .B(nbus_11295[13]), .C(n_58408),
		 .D(n_27998), .Z(n_210479605));
	notech_and4 i_123860555(.A(n_210479605), .B(n_93835734), .C(n_182479328)
		, .D(n_182779331), .Z(n_210779608));
	notech_and2 i_151058498(.A(n_57922), .B(n_212179622), .Z(n_210879609));
	notech_ao3 i_53257962(.A(n_56367), .B(opa[0]), .C(n_58184), .Z(n_211179612
		));
	notech_ao3 i_53357961(.A(n_56367), .B(\opa_12[0] ), .C(n_58184), .Z(n_211279613
		));
	notech_and2 i_14658347(.A(n_58646), .B(n_211679617), .Z(n_211379614));
	notech_and2 i_14758346(.A(n_236479865), .B(n_58610), .Z(n_211479615));
	notech_nand3 i_14858345(.A(n_57864), .B(n_57025), .C(n_220979710), .Z(n_211579616
		));
	notech_nao3 i_90157621(.A(n_56432), .B(opa[0]), .C(n_54756), .Z(n_211679617
		));
	notech_and2 i_14358350(.A(n_58646), .B(n_212079621), .Z(n_211779618));
	notech_and3 i_14458349(.A(n_228579786), .B(n_57863), .C(n_323280733), .Z
		(n_211879619));
	notech_nao3 i_94357580(.A(n_56443), .B(opa[0]), .C(n_54709), .Z(n_212079621
		));
	notech_or4 i_103157496(.A(n_55581), .B(n_57051), .C(n_29658), .D(n_57729
		), .Z(n_212179622));
	notech_or4 i_45858036(.A(n_56822), .B(n_56979), .C(n_56601), .D(n_27992)
		, .Z(n_212279623));
	notech_or4 i_45758037(.A(n_62856), .B(n_62788), .C(n_56127), .D(n_26054)
		, .Z(n_212579626));
	notech_nand3 i_45258042(.A(n_27029), .B(n_26669), .C(\opa_12[9] ), .Z(n_213079631
		));
	notech_or4 i_46758027(.A(n_26767), .B(n_60926), .C(n_28136), .D(n_26054)
		, .Z(n_213379634));
	notech_or2 i_46458030(.A(n_302291801), .B(\nbus_11358[10] ), .Z(n_213679637
		));
	notech_or4 i_46158033(.A(n_3854), .B(n_26054), .C(n_3850), .D(n_58024), 
		.Z(n_213979640));
	notech_nao3 i_47758017(.A(n_62826), .B(opc[11]), .C(n_301991804), .Z(n_214079641
		));
	notech_or4 i_47658018(.A(n_26767), .B(n_60924), .C(n_28137), .D(n_54934)
		, .Z(n_214379644));
	notech_or4 i_47358021(.A(n_62856), .B(n_62788), .C(n_29596), .D(n_54934)
		, .Z(n_214679647));
	notech_or4 i_47058024(.A(n_54954), .B(n_54934), .C(n_32335), .D(n_29596)
		, .Z(n_214979650));
	notech_or2 i_53157963(.A(n_57982), .B(n_56028), .Z(n_215079651));
	notech_or4 i_53057964(.A(n_58802), .B(n_26852), .C(nbus_11295[0]), .D(n_60924
		), .Z(n_215379654));
	notech_or4 i_52757967(.A(n_56675), .B(n_59993), .C(n_59275), .D(n_59355)
		, .Z(n_215679657));
	notech_ao4 i_52257972(.A(n_57730), .B(n_26662), .C(n_26904), .D(n_211179612
		), .Z(n_215779658));
	notech_ao4 i_52357971(.A(n_189662168), .B(n_305291771), .C(n_26905), .D(n_211279613
		), .Z(n_215879659));
	notech_or4 i_52457970(.A(n_62856), .B(n_284480345), .C(n_60924), .D(n_59742
		), .Z(n_215979660));
	notech_or4 i_80857709(.A(n_54814), .B(n_60924), .C(n_28136), .D(n_58481)
		, .Z(n_216079661));
	notech_nand2 i_80757710(.A(opd[10]), .B(n_58377), .Z(n_216379664));
	notech_or2 i_80257715(.A(n_3850), .B(n_181779321), .Z(n_216879669));
	notech_nao3 i_81857699(.A(n_62798), .B(opc[11]), .C(n_58038), .Z(n_216979670
		));
	notech_nao3 i_81757700(.A(n_54814), .B(n_26821), .C(n_31492), .Z(n_217279673
		));
	notech_nand2 i_81457703(.A(n_58377), .B(opd[11]), .Z(n_217579676));
	notech_nand2 i_81157706(.A(opa[11]), .B(n_58053), .Z(n_217879679));
	notech_or4 i_83957680(.A(n_58806), .B(n_60924), .C(n_28136), .D(n_56803)
		, .Z(n_217979680));
	notech_or2 i_83757681(.A(n_56356), .B(nbus_11295[10]), .Z(n_218279683)
		);
	notech_nand2 i_83457684(.A(opb[10]), .B(n_58050), .Z(n_218579686));
	notech_or4 i_83157687(.A(n_58132), .B(n_56803), .C(n_3850), .D(n_56903),
		 .Z(n_218879689));
	notech_or2 i_84957671(.A(n_56356), .B(nbus_11295[11]), .Z(n_219379694)
		);
	notech_or4 i_84557674(.A(n_62860), .B(n_62788), .C(n_29596), .D(n_56803)
		, .Z(n_219679697));
	notech_or4 i_84257677(.A(n_58132), .B(n_56803), .C(n_302491799), .D(n_56903
		), .Z(n_219979700));
	notech_or4 i_90057622(.A(n_54765), .B(n_266380164), .C(nbus_11295[0]), .D
		(n_60924), .Z(n_220079701));
	notech_or4 i_89957623(.A(n_54765), .B(n_28124), .C(n_60924), .D(n_58486)
		, .Z(n_220379704));
	notech_nand2 i_89457628(.A(opb[0]), .B(n_211579616), .Z(n_220879709));
	notech_or4 i_90457618(.A(n_32342), .B(n_32339), .C(n_54756), .D(n_58502)
		, .Z(n_220979710));
	notech_or4 i_91457609(.A(n_54765), .B(n_60924), .C(n_28136), .D(n_54736)
		, .Z(n_221279713));
	notech_or2 i_91357610(.A(n_58374), .B(n_27993), .Z(n_221579716));
	notech_or2 i_90857615(.A(n_3850), .B(n_57025), .Z(n_222079721));
	notech_nao3 i_92457599(.A(n_62798), .B(opc[11]), .C(n_313270143), .Z(n_222179722
		));
	notech_or4 i_92357600(.A(n_54765), .B(n_60924), .C(n_28137), .D(n_54736)
		, .Z(n_222479725));
	notech_or4 i_92057603(.A(n_62856), .B(n_62788), .C(n_56190), .D(n_54736)
		, .Z(n_222779728));
	notech_or4 i_91757606(.A(n_54756), .B(n_54736), .C(n_32331), .D(n_56190)
		, .Z(n_223079731));
	notech_or4 i_94257581(.A(n_54718), .B(n_28124), .C(n_60924), .D(n_26816)
		, .Z(n_223179732));
	notech_or4 i_94157582(.A(n_54718), .B(n_26807), .C(nbus_11295[0]), .D(n_60924
		), .Z(n_223479735));
	notech_ao4 i_93657587(.A(n_305291771), .B(n_240762674), .C(n_26905), .D(n_26771
		), .Z(n_223979740));
	notech_or4 i_95757568(.A(n_54718), .B(n_60924), .C(n_28136), .D(n_58479)
		, .Z(n_224279743));
	notech_or4 i_95657569(.A(n_54718), .B(n_58495), .C(n_60924), .D(nbus_11295
		[10]), .Z(n_224579746));
	notech_nand2 i_95257572(.A(opb[10]), .B(n_57179), .Z(n_224879749));
	notech_or2 i_94957575(.A(n_3850), .B(n_228579786), .Z(n_225179752));
	notech_or4 i_96757559(.A(n_54718), .B(n_58495), .C(n_60926), .D(nbus_11295
		[11]), .Z(n_225679757));
	notech_or4 i_96357562(.A(n_62858), .B(n_62810), .C(n_56190), .D(n_58479)
		, .Z(n_225979760));
	notech_or4 i_96057565(.A(n_62856), .B(n_228779788), .C(n_60926), .D(n_56190
		), .Z(n_226279763));
	notech_or2 i_98957538(.A(n_3850), .B(n_57299), .Z(n_226379764));
	notech_nao3 i_98857539(.A(n_26829), .B(\opa_12[10] ), .C(n_54678), .Z(n_226679767
		));
	notech_or2 i_98357544(.A(n_58376), .B(n_27993), .Z(n_227179772));
	notech_nao3 i_100457523(.A(n_62798), .B(opc_10[11]), .C(n_57473), .Z(n_227279773
		));
	notech_or2 i_100357524(.A(n_57807), .B(\nbus_11358[11] ), .Z(n_227579776
		));
	notech_or2 i_100057527(.A(n_30528), .B(n_56636), .Z(n_227879779));
	notech_or4 i_99757530(.A(n_54678), .B(n_58087), .C(n_32338), .D(n_56190)
		, .Z(n_228179782));
	notech_nand3 i_30918(.A(n_26790), .B(n_26825), .C(n_56903), .Z(n_228279783
		));
	notech_nand2 i_30917(.A(n_58806), .B(n_26825), .Z(n_228379784));
	notech_or4 i_30916(.A(n_32326), .B(n_32339), .C(n_58132), .D(n_56803), .Z
		(n_228479785));
	notech_or4 i_29852(.A(n_101413114), .B(n_54709), .C(instrc[121]), .D(n_58479
		), .Z(n_228579786));
	notech_nao3 i_29851(.A(n_26828), .B(n_56443), .C(n_54709), .Z(n_228679787
		));
	notech_nand2 i_29849(.A(n_54718), .B(n_26828), .Z(n_228779788));
	notech_and2 i_29601(.A(n_229779798), .B(n_229679797), .Z(n_228879789));
	notech_nao3 i_4758444(.A(n_60292), .B(opa[1]), .C(n_3852), .Z(n_229179792
		));
	notech_nand3 i_5758434(.A(n_2988), .B(n_60292), .C(opb[1]), .Z(n_229279793
		));
	notech_or4 i_29953(.A(n_54727), .B(n_57078), .C(instrc[116]), .D(n_26807
		), .Z(n_229379794));
	notech_nand2 i_29950(.A(n_54718), .B(n_56482), .Z(n_229479795));
	notech_and3 i_191256638(.A(n_276234718), .B(n_229179792), .C(n_229279793
		), .Z(n_229679797));
	notech_ao4 i_191056640(.A(n_58432), .B(n_60024), .C(n_58391), .D(n_29678
		), .Z(n_229779798));
	notech_ao4 i_184656703(.A(n_31492), .B(n_184768864), .C(n_302491799), .D
		(n_184668863), .Z(n_230079801));
	notech_ao4 i_184456705(.A(n_58376), .B(n_27996), .C(n_31456), .D(n_54678
		), .Z(n_230279803));
	notech_and4 i_184856701(.A(n_230279803), .B(n_230079801), .C(n_227879779
		), .D(n_228179782), .Z(n_230479805));
	notech_ao4 i_184156708(.A(nbus_11295[11]), .B(n_26823), .C(n_57809), .D(\nbus_11307[11] 
		), .Z(n_230579806));
	notech_and4 i_184356706(.A(n_187368889), .B(n_227279773), .C(n_230579806
		), .D(n_227579776), .Z(n_230879809));
	notech_ao4 i_183456715(.A(n_54678), .B(n_31411), .C(n_56636), .D(n_187568890
		), .Z(n_230979810));
	notech_ao4 i_183356716(.A(nbus_11295[10]), .B(n_26823), .C(n_57809), .D(\nbus_11307[10] 
		), .Z(n_231179812));
	notech_ao4 i_183056719(.A(n_31433), .B(n_57473), .C(n_57807), .D(\nbus_11358[10] 
		), .Z(n_231379814));
	notech_and4 i_183256717(.A(n_187968894), .B(n_231379814), .C(n_226379764
		), .D(n_226679767), .Z(n_231679817));
	notech_ao4 i_181756732(.A(n_56190), .B(n_228679787), .C(n_302491799), .D
		(n_228579786), .Z(n_231779818));
	notech_ao4 i_181556734(.A(\nbus_11358[11] ), .B(n_26855), .C(\nbus_11307[11] 
		), .D(n_26856), .Z(n_231979820));
	notech_and4 i_181956730(.A(n_231979820), .B(n_231779818), .C(n_225979760
		), .D(n_226279763), .Z(n_232179822));
	notech_ao4 i_181256737(.A(n_30528), .B(n_56662), .C(n_27996), .D(n_58375
		), .Z(n_232279823));
	notech_ao4 i_181056739(.A(n_30088), .B(n_323080731), .C(n_31476), .D(n_322780728
		), .Z(n_232479825));
	notech_and4 i_181456735(.A(n_187368889), .B(n_232479825), .C(n_232279823
		), .D(n_225679757), .Z(n_232679827));
	notech_ao4 i_180756742(.A(n_87532846), .B(n_323080731), .C(n_187568890),
		 .D(n_56662), .Z(n_232779828));
	notech_ao4 i_180556744(.A(\nbus_11307[10] ), .B(n_26856), .C(n_322980730
		), .D(n_56145), .Z(n_232979830));
	notech_and4 i_180956740(.A(n_232979830), .B(n_232779828), .C(n_224879749
		), .D(n_225179752), .Z(n_233179832));
	notech_ao4 i_180256747(.A(n_58375), .B(n_27993), .C(n_31411), .D(n_58479
		), .Z(n_233279833));
	notech_and4 i_180456745(.A(n_187968894), .B(n_224279743), .C(n_233279833
		), .D(n_224579746), .Z(n_233579836));
	notech_ao4 i_179956750(.A(n_56046), .B(n_57249), .C(n_56037), .D(n_57316
		), .Z(n_233679837));
	notech_ao4 i_179656753(.A(n_56028), .B(n_211879619), .C(n_26807), .D(n_211779618
		), .Z(n_233879839));
	notech_ao4 i_179556754(.A(n_291363180), .B(n_143071910), .C(n_175062033)
		, .D(n_229479795), .Z(n_234079841));
	notech_ao4 i_179256757(.A(n_59993), .B(n_143571915), .C(n_143471914), .D
		(n_59187), .Z(n_234279843));
	notech_and4 i_179456755(.A(n_152275466), .B(n_223179732), .C(n_234279843
		), .D(n_223479735), .Z(n_234579846));
	notech_ao4 i_177956769(.A(n_31492), .B(n_184468861), .C(n_302491799), .D
		(n_184368860), .Z(n_234679847));
	notech_ao4 i_177756771(.A(n_57181), .B(\nbus_11358[11] ), .C(\nbus_11307[11] 
		), .D(n_26607), .Z(n_234879849));
	notech_and4 i_178156767(.A(n_234879849), .B(n_223079731), .C(n_234679847
		), .D(n_222779728), .Z(n_235079851));
	notech_ao4 i_177456774(.A(n_30528), .B(n_56649), .C(n_27996), .D(n_58374
		), .Z(n_235179852));
	notech_and4 i_177656772(.A(n_187368889), .B(n_222479725), .C(n_235179852
		), .D(n_222179722), .Z(n_235479855));
	notech_ao4 i_177056778(.A(n_87532846), .B(n_313270143), .C(n_187568890),
		 .D(n_56649), .Z(n_235579856));
	notech_ao4 i_176956779(.A(\nbus_11307[10] ), .B(n_26607), .C(n_319970210
		), .D(n_56145), .Z(n_235779858));
	notech_ao4 i_176656782(.A(n_31411), .B(n_54736), .C(n_57181), .D(\nbus_11358[10] 
		), .Z(n_235979860));
	notech_and4 i_176856780(.A(n_187968894), .B(n_235979860), .C(n_221279713
		), .D(n_221579716), .Z(n_236279863));
	notech_ao4 i_176456784(.A(n_56046), .B(n_57322), .C(n_56037), .D(n_151731932
		), .Z(n_236479865));
	notech_ao4 i_176056788(.A(n_58486), .B(n_211479615), .C(n_266380164), .D
		(n_211379614), .Z(n_236579866));
	notech_ao4 i_175956789(.A(n_147171951), .B(n_59187), .C(n_175062033), .D
		(n_247579976), .Z(n_236779868));
	notech_ao4 i_175656792(.A(n_291363180), .B(n_178472264), .C(n_59993), .D
		(n_147271952), .Z(n_236979870));
	notech_and4 i_175856790(.A(n_152275466), .B(n_236979870), .C(n_220379704
		), .D(n_220079701), .Z(n_237279873));
	notech_ao4 i_171856830(.A(n_31492), .B(n_228379784), .C(n_56190), .D(n_228279783
		), .Z(n_237379874));
	notech_ao4 i_171656832(.A(\nbus_11358[11] ), .B(n_26853), .C(\nbus_11307[11] 
		), .D(n_26854), .Z(n_237579876));
	notech_and4 i_172056828(.A(n_237579876), .B(n_237379874), .C(n_219679697
		), .D(n_219979700), .Z(n_237779878));
	notech_ao4 i_171356835(.A(n_30528), .B(n_56914), .C(n_27996), .D(n_58372
		), .Z(n_237879879));
	notech_ao4 i_171156837(.A(n_30088), .B(n_58041), .C(n_31476), .D(n_322580726
		), .Z(n_238079881));
	notech_and4 i_171556833(.A(n_187368889), .B(n_238079881), .C(n_237879879
		), .D(n_219379694), .Z(n_238279883));
	notech_ao4 i_170856840(.A(n_87532846), .B(n_58041), .C(n_187568890), .D(n_56914
		), .Z(n_238379884));
	notech_ao4 i_170656842(.A(\nbus_11307[10] ), .B(n_26854), .C(n_322680727
		), .D(n_56145), .Z(n_238579886));
	notech_and4 i_171056838(.A(n_238579886), .B(n_218879689), .C(n_238379884
		), .D(n_218579686), .Z(n_238779888));
	notech_ao4 i_170356845(.A(n_58372), .B(n_27993), .C(n_31411), .D(n_56803
		), .Z(n_238879889));
	notech_and4 i_170556843(.A(n_187968894), .B(n_217979680), .C(n_238879889
		), .D(n_218279683), .Z(n_239179892));
	notech_ao4 i_169156857(.A(n_181679320), .B(n_56190), .C(n_302491799), .D
		(n_181779321), .Z(n_239279893));
	notech_ao4 i_168956859(.A(n_31456), .B(n_58481), .C(n_58052), .D(\nbus_11358[11] 
		), .Z(n_239479895));
	notech_and4 i_169356855(.A(n_239479895), .B(n_239279893), .C(n_217579676
		), .D(n_217879679), .Z(n_239679897));
	notech_ao4 i_168656862(.A(n_31476), .B(n_57765), .C(n_30528), .D(n_56498
		), .Z(n_239779898));
	notech_and4 i_168856860(.A(n_187368889), .B(n_239779898), .C(n_216979670
		), .D(n_217279673), .Z(n_240079901));
	notech_ao4 i_168256866(.A(n_87532846), .B(n_58038), .C(n_187568890), .D(n_56498
		), .Z(n_240179902));
	notech_ao4 i_168156867(.A(n_57625), .B(n_26851), .C(n_197279473), .D(n_56145
		), .Z(n_240379904));
	notech_ao4 i_167856870(.A(n_31411), .B(n_58481), .C(n_58052), .D(\nbus_11358[10] 
		), .Z(n_240579906));
	notech_and4 i_168056868(.A(n_187968894), .B(n_216079661), .C(n_240579906
		), .D(n_216379664), .Z(n_240879909));
	notech_ao3 i_139157150(.A(n_215979660), .B(n_26777), .C(n_215779658), .Z
		(n_241079911));
	notech_ao4 i_138857153(.A(n_56046), .B(n_284880349), .C(n_284580346), .D
		(n_59187), .Z(n_241179912));
	notech_ao4 i_138557156(.A(n_291163178), .B(n_57915), .C(n_178572265), .D
		(n_291363180), .Z(n_241479915));
	notech_and4 i_138757154(.A(n_152275466), .B(n_241479915), .C(n_215079651
		), .D(n_215379654), .Z(n_241779918));
	notech_ao4 i_134857193(.A(n_25875), .B(n_302491799), .C(n_31492), .D(n_25874
		), .Z(n_241879919));
	notech_ao4 i_134657195(.A(n_302291801), .B(n_56181), .C(n_57635), .D(n_27293
		), .Z(n_242079921));
	notech_and4 i_135057191(.A(n_242079921), .B(n_214979650), .C(n_241879919
		), .D(n_214679647), .Z(n_242279923));
	notech_ao4 i_134257198(.A(n_30528), .B(n_56601), .C(n_27996), .D(n_302391800
		), .Z(n_242379924));
	notech_and4 i_134457196(.A(n_242379924), .B(n_187368889), .C(n_214079641
		), .D(n_214379644), .Z(n_242679927));
	notech_ao4 i_133757202(.A(n_87532846), .B(n_301991804), .C(n_187568890),
		 .D(n_56601), .Z(n_242779928));
	notech_ao4 i_133557204(.A(n_57625), .B(n_27293), .C(n_322480725), .D(n_56145
		), .Z(n_242979930));
	notech_and4 i_134057200(.A(n_242979930), .B(n_242779928), .C(n_213679637
		), .D(n_213979640), .Z(n_243179932));
	notech_ao4 i_133257207(.A(n_302391800), .B(n_27993), .C(n_31411), .D(n_54934
		), .Z(n_243279933));
	notech_and4 i_133457205(.A(n_54667), .B(n_243279933), .C(n_187968894), .D
		(n_213379634), .Z(n_243579936));
	notech_ao4 i_132857211(.A(n_27293), .B(n_57613), .C(n_189962171), .D(n_210879609
		), .Z(n_243679937));
	notech_ao4 i_132757212(.A(n_302291801), .B(n_56136), .C(n_60016), .D(n_25875
		), .Z(n_243879939));
	notech_ao4 i_132457215(.A(n_25884), .B(n_291963186), .C(n_56601), .D(n_58106
		), .Z(n_244079941));
	notech_and4 i_132657213(.A(n_200065529), .B(n_244079941), .C(n_212279623
		), .D(n_212579626), .Z(n_244379944));
	notech_and3 i_10055417(.A(n_246279963), .B(n_246179962), .C(n_58610), .Z
		(n_244479945));
	notech_ao3 i_10155416(.A(n_244979950), .B(n_245779958), .C(n_245879959),
		 .Z(n_244579946));
	notech_ao4 i_10355414(.A(n_62892), .B(n_2480), .C(n_56822), .D(n_32299),
		 .Z(n_244679947));
	notech_nao3 i_40355122(.A(n_58806), .B(n_56809), .C(n_175062033), .Z(n_244979950
		));
	notech_or4 i_40155124(.A(n_58132), .B(n_56903), .C(n_56028), .D(n_314360224
		), .Z(n_245779958));
	notech_ao4 i_40255123(.A(n_56979), .B(n_26627), .C(n_26904), .D(n_26793)
		, .Z(n_245879959));
	notech_nand3 i_39955126(.A(n_56903), .B(\opa_12[0] ), .C(n_26790), .Z(n_246179962
		));
	notech_or4 i_40055125(.A(n_58132), .B(n_56046), .C(n_32326), .D(n_32339)
		, .Z(n_246279963));
	notech_or2 i_42855097(.A(n_57154), .B(n_56010), .Z(n_246779968));
	notech_nand3 i_42555100(.A(n_26792), .B(n_26805), .C(\opa_12[1] ), .Z(n_247079971
		));
	notech_or4 i_42255103(.A(n_54756), .B(n_280073280), .C(n_32331), .D(n_57542
		), .Z(n_247379974));
	notech_or2 i_30295(.A(n_54765), .B(n_266380164), .Z(n_247479975));
	notech_nand2 i_30292(.A(n_54765), .B(n_26806), .Z(n_247579976));
	notech_nand2 i_30272(.A(n_26792), .B(n_26805), .Z(n_247679977));
	notech_ao4 i_88954694(.A(n_147271952), .B(n_59992), .C(n_147171951), .D(n_59241
		), .Z(n_247779978));
	notech_ao4 i_88754696(.A(n_247579976), .B(n_297866507), .C(n_297966508),
		 .D(n_247479975), .Z(n_247979980));
	notech_and4 i_89154692(.A(n_247979980), .B(n_247779978), .C(n_247079971)
		, .D(n_247379974), .Z(n_248179982));
	notech_ao4 i_88354699(.A(n_57141), .B(n_298066509), .C(n_60024), .D(n_57084
		), .Z(n_248279983));
	notech_ao4 i_88154701(.A(n_58486), .B(n_297666505), .C(n_297766506), .D(n_266380164
		), .Z(n_248479985));
	notech_and4 i_88654697(.A(n_228879789), .B(n_248479985), .C(n_248279983)
		, .D(n_246779968), .Z(n_248679987));
	notech_nand2 i_84754732(.A(n_56903), .B(opa[0]), .Z(n_249079991));
	notech_ao4 i_84654733(.A(n_58806), .B(n_291263179), .C(n_58132), .D(n_249079991
		), .Z(n_249179992));
	notech_ao4 i_83954736(.A(n_244679947), .B(n_244579946), .C(n_26804), .D(n_244479945
		), .Z(n_249379994));
	notech_ao4 i_83854737(.A(n_57773), .B(n_56914), .C(n_56356), .D(nbus_11295
		[0]), .Z(n_249479995));
	notech_ao4 i_83654739(.A(n_291163178), .B(n_257980080), .C(n_147471954),
		 .D(n_291363180), .Z(n_249679997));
	notech_ao3 i_10950557(.A(tsc[24]), .B(n_55820), .C(n_59469), .Z(n_249879999
		));
	notech_or2 i_10850558(.A(n_59124), .B(nbus_11295[24]), .Z(n_250180002)
		);
	notech_or2 i_10550561(.A(n_60001), .B(n_151428791), .Z(n_250480005));
	notech_or2 i_10250564(.A(n_289027272), .B(n_151128788), .Z(n_250780008)
		);
	notech_nor2 i_37350295(.A(n_57868), .B(n_57742), .Z(n_250880009));
	notech_or2 i_36850300(.A(n_289227274), .B(n_154831963), .Z(n_251580016)
		);
	notech_ao3 i_80149886(.A(n_32304), .B(opd[22]), .C(n_56688), .Z(n_251680017
		));
	notech_nand2 i_79649891(.A(n_287027252), .B(\regs_13_14[22] ), .Z(n_252380024
		));
	notech_ao3 i_81749870(.A(n_32304), .B(opd[24]), .C(n_56688), .Z(n_252480025
		));
	notech_nand2 i_81249875(.A(n_287027252), .B(\regs_13_14[24] ), .Z(n_253180032
		));
	notech_or2 i_85749830(.A(n_57867), .B(n_57751), .Z(n_253280033));
	notech_or2 i_85649831(.A(n_57865), .B(n_56347), .Z(n_253580036));
	notech_or2 i_85149836(.A(n_289127273), .B(n_305624320), .Z(n_254080041)
		);
	notech_ao4 i_177248935(.A(n_58007), .B(n_225665785), .C(n_222565754), .D
		(n_58008), .Z(n_254180042));
	notech_ao4 i_177148936(.A(n_29765), .B(n_26937), .C(n_58423), .D(n_28008
		), .Z(n_254380044));
	notech_ao4 i_176848939(.A(n_60002), .B(n_58138), .C(n_57726), .D(n_28149
		), .Z(n_254580046));
	notech_and4 i_177048937(.A(n_254580046), .B(n_253280033), .C(n_253580036
		), .D(n_26618), .Z(n_254880049));
	notech_ao4 i_173748970(.A(n_286927251), .B(n_221065739), .C(n_286827250)
		, .D(n_225565784), .Z(n_254980050));
	notech_ao4 i_173648971(.A(n_57861), .B(n_57761), .C(n_287827260), .D(n_289027272
		), .Z(n_255180052));
	notech_nand3 i_173948968(.A(n_254980050), .B(n_255180052), .C(n_253180032
		), .Z(n_255280053));
	notech_ao4 i_173448973(.A(n_58139), .B(n_60001), .C(n_57863), .D(n_56475
		), .Z(n_255380054));
	notech_ao4 i_172348984(.A(n_286927251), .B(n_224065769), .C(n_286827250)
		, .D(n_225765786), .Z(n_255680057));
	notech_ao4 i_172248985(.A(n_57861), .B(n_57742), .C(n_287827260), .D(n_289227274
		), .Z(n_255880059));
	notech_nand3 i_172548982(.A(n_255680057), .B(n_255880059), .C(n_252380024
		), .Z(n_255980060));
	notech_ao4 i_172048987(.A(n_58139), .B(n_60003), .C(n_57863), .D(n_56338
		), .Z(n_256080061));
	notech_ao4 i_132549374(.A(n_225765786), .B(n_151931934), .C(n_224065769)
		, .D(n_58084), .Z(n_256380064));
	notech_ao4 i_132449375(.A(n_29708), .B(n_26929), .C(n_58429), .D(n_28007
		), .Z(n_256580066));
	notech_nand3 i_132749372(.A(n_256380064), .B(n_256580066), .C(n_251580016
		), .Z(n_256680067));
	notech_ao4 i_132249377(.A(n_57875), .B(n_56338), .C(n_60003), .D(n_58147
		), .Z(n_256780068));
	notech_ao4 i_109549600(.A(n_225565784), .B(n_311391710), .C(n_221065739)
		, .D(n_311491709), .Z(n_257080071));
	notech_ao4 i_109349602(.A(n_29769), .B(n_26696), .C(n_311291711), .D(n_28009
		), .Z(n_257280073));
	notech_and4 i_109749598(.A(n_257280073), .B(n_257080071), .C(n_250480005
		), .D(n_250780008), .Z(n_257480075));
	notech_ao4 i_109049605(.A(n_311091713), .B(n_57761), .C(n_311191712), .D
		(n_56475), .Z(n_257580076));
	notech_nand2 i_109149604(.A(n_257580076), .B(n_250180002), .Z(n_257680077
		));
	notech_or4 i_116955586(.A(n_57026), .B(n_56863), .C(n_26804), .D(n_57033
		), .Z(n_257980080));
	notech_or2 i_116246575(.A(n_54765), .B(n_258180082), .Z(n_258080081));
	notech_and3 i_186155564(.A(n_56843), .B(n_187762157), .C(n_54736), .Z(n_258180082
		));
	notech_or4 i_116746570(.A(n_57026), .B(n_56863), .C(n_57033), .D(n_57827
		), .Z(n_258280083));
	notech_or4 i_28847412(.A(n_54954), .B(n_3845), .C(n_58020), .D(n_56302),
		 .Z(n_258580086));
	notech_or4 i_28547415(.A(n_56824), .B(n_56946), .C(n_56601), .D(n_28003)
		, .Z(n_258880089));
	notech_or4 i_28247418(.A(n_3845), .B(n_26767), .C(n_60926), .D(nbus_11295
		[18]), .Z(n_259180092));
	notech_or2 i_68947034(.A(n_56356), .B(nbus_11295[16]), .Z(n_259280093)
		);
	notech_or4 i_68847035(.A(n_58132), .B(n_58493), .C(n_56903), .D(\nbus_11358[16] 
		), .Z(n_259580096));
	notech_or4 i_68547038(.A(n_56822), .B(n_56979), .C(n_56914), .D(n_313747721
		), .Z(n_259880099));
	notech_or4 i_68247041(.A(n_62858), .B(n_58493), .C(n_62788), .D(\nbus_11365[16] 
		), .Z(n_260180102));
	notech_nor2 i_70947014(.A(n_56356), .B(nbus_11295[18]), .Z(n_260280103)
		);
	notech_or4 i_70847015(.A(n_56822), .B(n_56946), .C(n_56914), .D(n_28003)
		, .Z(n_260580106));
	notech_or2 i_70547018(.A(n_58143), .B(n_3864), .Z(n_260880109));
	notech_or2 i_70247021(.A(n_286869880), .B(n_57698), .Z(n_261180112));
	notech_nand2 i_32634(.A(n_312491699), .B(n_27102), .Z(n_261280113));
	notech_ao4 i_171346047(.A(n_306124325), .B(n_77522039), .C(n_305924323),
		 .D(n_3861), .Z(n_261380114));
	notech_ao4 i_171146049(.A(n_58085), .B(n_95222216), .C(n_60121865), .D(n_58493
		), .Z(n_261580116));
	notech_and4 i_171546045(.A(n_261580116), .B(n_261380114), .C(n_260880109
		), .D(n_261180112), .Z(n_261780118));
	notech_ao4 i_170846052(.A(n_57877), .B(n_56302), .C(n_26902), .D(n_29711
		), .Z(n_261880119));
	notech_nand2 i_170946051(.A(n_261880119), .B(n_260580106), .Z(n_261980120
		));
	notech_ao4 i_169346065(.A(n_311224366), .B(n_56914), .C(n_286869880), .D
		(\nbus_11365[16] ), .Z(n_262280123));
	notech_ao4 i_169146067(.A(n_254466073), .B(n_266280163), .C(n_252966058)
		, .D(n_58085), .Z(n_262480125));
	notech_and4 i_169546063(.A(n_262480125), .B(n_262280123), .C(n_259880099
		), .D(n_260180102), .Z(n_262680127));
	notech_ao4 i_168846070(.A(n_29710), .B(n_26902), .C(n_60009), .D(n_58143
		), .Z(n_262780128));
	notech_and4 i_169046068(.A(n_194675885), .B(n_262780128), .C(n_259280093
		), .D(n_259580096), .Z(n_263080131));
	notech_nand2 i_5047649(.A(n_26670), .B(n_27029), .Z(n_263180132));
	notech_ao4 i_135846386(.A(n_60121865), .B(n_3845), .C(n_263180132), .D(n_57698
		), .Z(n_263280133));
	notech_ao4 i_135646388(.A(n_3861), .B(n_3837), .C(n_77522039), .D(n_3843
		), .Z(n_263480135));
	notech_and4 i_136046384(.A(n_258880089), .B(n_263480135), .C(n_263280133
		), .D(n_259180092), .Z(n_263680137));
	notech_ao4 i_135346391(.A(n_3864), .B(n_148228759), .C(n_29711), .D(n_26642
		), .Z(n_263780138));
	notech_and4 i_135546389(.A(n_54667), .B(n_263780138), .C(n_258580086), .D
		(n_26621), .Z(n_264080141));
	notech_and2 i_14744349(.A(n_92619108), .B(n_264380144), .Z(n_264180142)
		);
	notech_ao4 i_14844348(.A(n_26895), .B(n_57592), .C(n_56082), .D(n_57758)
		, .Z(n_264280143));
	notech_nao3 i_46544035(.A(n_56367), .B(\opa_12[6] ), .C(n_58184), .Z(n_264380144
		));
	notech_and2 i_14044356(.A(n_313291691), .B(n_52335319), .Z(n_264680147)
		);
	notech_ao4 i_14144355(.A(n_27349), .B(n_29619), .C(n_303791786), .D(\nbus_11365[31] 
		), .Z(n_264780148));
	notech_and2 i_14244354(.A(n_27348), .B(n_265280153), .Z(n_264880149));
	notech_nand3 i_54043967(.A(n_312491699), .B(n_30946), .C(n_2026), .Z(n_265280153
		));
	notech_nand3 i_66343853(.A(n_60127), .B(n_60246), .C(read_data[31]), .Z(n_265380154
		));
	notech_ao4 i_5544439(.A(n_26810), .B(n_59223), .C(n_308721251), .D(n_56675
		), .Z(n_265480155));
	notech_ao4 i_5444440(.A(n_26810), .B(n_59205), .C(n_308621250), .D(n_56675
		), .Z(n_265780158));
	notech_and2 i_150447762(.A(n_257980080), .B(n_258280083), .Z(n_266280163
		));
	notech_and4 i_187155563(.A(n_56843), .B(n_58494), .C(n_187762157), .D(n_54736
		), .Z(n_266380164));
	notech_nao3 i_125043312(.A(n_57730), .B(n_32344), .C(n_58184), .Z(n_266680167
		));
	notech_or2 i_44444053(.A(n_57982), .B(\nbus_11358[3] ), .Z(n_266780168)
		);
	notech_or4 i_44344054(.A(n_62858), .B(n_26812), .C(n_62788), .D(n_29728)
		, .Z(n_267080171));
	notech_or2 i_44044057(.A(n_265480155), .B(n_56485), .Z(n_267380174));
	notech_nao3 i_43744060(.A(n_26811), .B(\opa_12[3] ), .C(n_26812), .Z(n_267680177
		));
	notech_or2 i_45744043(.A(n_57982), .B(\nbus_11358[5] ), .Z(n_267780178)
		);
	notech_or4 i_45644044(.A(n_62858), .B(n_26812), .C(n_62788), .D(n_29651)
		, .Z(n_268080181));
	notech_or2 i_45344047(.A(n_56485), .B(n_265780158), .Z(n_268380184));
	notech_nao3 i_45044050(.A(n_26811), .B(\opa_12[5] ), .C(n_26812), .Z(n_268680187
		));
	notech_or4 i_46444036(.A(n_26812), .B(n_58802), .C(n_60926), .D(n_28131)
		, .Z(n_268780188));
	notech_nand3 i_53543971(.A(n_54834), .B(n_7344), .C(n_56172), .Z(n_269480195
		));
	notech_nand3 i_53443972(.A(n_7343), .B(n_56163), .C(n_54834), .Z(n_269780198
		));
	notech_nand3 i_53143975(.A(n_27340), .B(n_62788), .C(opc[31]), .Z(n_270080201
		));
	notech_or2 i_52743978(.A(n_313491689), .B(n_264780148), .Z(n_270380204)
		);
	notech_or4 i_67843838(.A(n_58133), .B(n_26906), .C(n_32322), .D(\nbus_11307[3] 
		), .Z(n_270480205));
	notech_or4 i_67743839(.A(n_62860), .B(n_58489), .C(n_62824), .D(n_29728)
		, .Z(n_270780208));
	notech_nao3 i_67443842(.A(n_318891635), .B(n_318791636), .C(n_265480155)
		, .Z(n_271080211));
	notech_nao3 i_67143845(.A(n_26813), .B(\opa_12[3] ), .C(n_58489), .Z(n_271380214
		));
	notech_or4 i_71843806(.A(n_58133), .B(n_26906), .C(n_32322), .D(\nbus_11307[5] 
		), .Z(n_271480215));
	notech_or4 i_71743807(.A(n_62856), .B(n_58489), .C(n_62788), .D(n_29651)
		, .Z(n_271780218));
	notech_nao3 i_71343810(.A(n_318891635), .B(n_318791636), .C(n_265780158)
		, .Z(n_272080221));
	notech_nao3 i_70843813(.A(n_26813), .B(\opa_12[5] ), .C(n_58489), .Z(n_272380224
		));
	notech_nao3 i_76743759(.A(n_26824), .B(\opa_12[3] ), .C(n_26804), .Z(n_272880229
		));
	notech_nao3 i_76443762(.A(n_58078), .B(opd[3]), .C(n_56914), .Z(n_273180232
		));
	notech_nao3 i_78243747(.A(n_26824), .B(\opa_12[5] ), .C(n_26804), .Z(n_274080241
		));
	notech_nao3 i_77943750(.A(n_58078), .B(opd[5]), .C(n_56914), .Z(n_274380244
		));
	notech_nand2 i_82243708(.A(\regs_13_14[31] ), .B(n_58144), .Z(n_274880249
		));
	notech_or2 i_82143709(.A(n_56356), .B(nbus_11295[31]), .Z(n_275180252)
		);
	notech_nao3 i_81643714(.A(n_62826), .B(opc_10[31]), .C(n_266280163), .Z(n_275680257
		));
	notech_or4 i_88543655(.A(n_54756), .B(n_280073280), .C(n_32331), .D(\nbus_11307[3] 
		), .Z(n_276180262));
	notech_or2 i_88043658(.A(n_308721251), .B(n_147271952), .Z(n_276480265)
		);
	notech_or4 i_87743661(.A(n_54765), .B(n_266380164), .C(nbus_11295[3]), .D
		(n_60926), .Z(n_276780268));
	notech_or4 i_89643644(.A(n_54756), .B(n_280073280), .C(n_32331), .D(\nbus_11307[5] 
		), .Z(n_277280273));
	notech_or2 i_89343647(.A(n_308621250), .B(n_147271952), .Z(n_277580276)
		);
	notech_or4 i_89043650(.A(n_54765), .B(n_266380164), .C(nbus_11295[5]), .D
		(n_60926), .Z(n_277880279));
	notech_and2 i_93243609(.A(n_26675), .B(\regs_13_14[31] ), .Z(n_277980280
		));
	notech_nao3 i_92743614(.A(n_62826), .B(opc_10[31]), .C(n_57116), .Z(n_278680287
		));
	notech_or4 i_94143600(.A(n_54709), .B(n_26807), .C(n_32332), .D(\nbus_11307[3] 
		), .Z(n_279180292));
	notech_or2 i_93843603(.A(n_308721251), .B(n_143571915), .Z(n_279480295)
		);
	notech_or4 i_93543606(.A(n_54718), .B(n_26807), .C(nbus_11295[3]), .D(n_60926
		), .Z(n_279780298));
	notech_or4 i_95243589(.A(n_58100), .B(n_26807), .C(n_32332), .D(n_57583)
		, .Z(n_280280303));
	notech_or2 i_94943592(.A(n_308621250), .B(n_143571915), .Z(n_280580306)
		);
	notech_or4 i_94643595(.A(n_58817), .B(n_26807), .C(nbus_11295[5]), .D(n_60924
		), .Z(n_280880309));
	notech_or4 i_100143544(.A(n_58087), .B(n_56529), .C(n_32338), .D(n_57563
		), .Z(n_281380314));
	notech_or2 i_99843547(.A(n_308721251), .B(n_124271722), .Z(n_281680317)
		);
	notech_nao3 i_99543550(.A(opc[3]), .B(n_62824), .C(n_123971719), .Z(n_281980320
		));
	notech_or4 i_101643529(.A(n_58087), .B(n_56529), .C(n_32338), .D(n_57583
		), .Z(n_282480325));
	notech_or4 i_101343532(.A(n_56822), .B(n_56979), .C(n_56636), .D(n_308621250
		), .Z(n_282780328));
	notech_or4 i_101043535(.A(n_282066349), .B(n_56863), .C(n_245362720), .D
		(n_56529), .Z(n_283080331));
	notech_or2 i_119843363(.A(n_122428501), .B(n_28157), .Z(n_283380334));
	notech_nao3 i_119543366(.A(n_19065), .B(read_data[31]), .C(n_59100), .Z(n_283680337
		));
	notech_or2 i_119243369(.A(n_122528502), .B(n_314791676), .Z(n_283980340)
		);
	notech_nand2 i_118943372(.A(add_len_pc[31]), .B(n_26766), .Z(n_284280343
		));
	notech_nao3 i_9944395(.A(n_56367), .B(n_58164), .C(n_58184), .Z(n_284380344
		));
	notech_nand2 i_9444400(.A(n_58802), .B(n_58164), .Z(n_284480345));
	notech_or2 i_33266(.A(n_56485), .B(n_26810), .Z(n_284580346));
	notech_or4 i_7944415(.A(n_26852), .B(n_57078), .C(n_57051), .D(n_54916),
		 .Z(n_284680347));
	notech_or2 i_9344401(.A(n_26812), .B(n_58419), .Z(n_284780348));
	notech_or2 i_8144413(.A(n_26812), .B(n_57758), .Z(n_284880349));
	notech_or2 i_7844416(.A(n_58489), .B(n_58421), .Z(n_284980350));
	notech_or4 i_7744417(.A(n_60854), .B(n_58133), .C(n_58489), .D(n_26735),
		 .Z(n_285080351));
	notech_ao4 i_211642474(.A(n_124328520), .B(n_314391680), .C(n_309391730)
		, .D(n_96519147), .Z(n_285180352));
	notech_ao4 i_211442476(.A(n_308991734), .B(\nbus_11365[31] ), .C(n_60127
		), .D(n_27269), .Z(n_285380354));
	notech_and4 i_211842472(.A(n_285380354), .B(n_285180352), .C(n_283980340
		), .D(n_284280343), .Z(n_285580356));
	notech_ao4 i_211142479(.A(n_121628493), .B(n_28016), .C(n_309091733), .D
		(\nbus_11358[31] ), .Z(n_285680357));
	notech_ao4 i_210942481(.A(n_26765), .B(n_29619), .C(n_56091), .D(n_30031
		), .Z(n_285880359));
	notech_and4 i_211342477(.A(n_285880359), .B(n_285680357), .C(n_283380334
		), .D(n_283680337), .Z(n_286080361));
	notech_ao4 i_198742602(.A(n_281966348), .B(n_56529), .C(n_281866347), .D
		(n_124171721), .Z(n_286180362));
	notech_ao4 i_198542604(.A(n_282266351), .B(n_58488), .C(n_282166350), .D
		(n_153979043), .Z(n_286380364));
	notech_and4 i_198942600(.A(n_286380364), .B(n_286180362), .C(n_282780328
		), .D(n_283080331), .Z(n_286580366));
	notech_ao4 i_198242607(.A(n_58044), .B(n_56073), .C(n_123771717), .D(n_59205
		), .Z(n_286680367));
	notech_ao4 i_198042609(.A(n_60020), .B(n_57470), .C(n_154079044), .D(n_29651
		), .Z(n_286880369));
	notech_and4 i_198442605(.A(n_216276101), .B(n_286880369), .C(n_286680367
		), .D(n_282480325), .Z(n_287080371));
	notech_ao4 i_197442615(.A(n_124171721), .B(n_306670077), .C(n_56529), .D
		(n_306570076), .Z(n_287180372));
	notech_ao4 i_197242617(.A(n_306970080), .B(n_58488), .C(n_306870079), .D
		(n_153979043), .Z(n_287380374));
	notech_and4 i_197642613(.A(n_287380374), .B(n_287180372), .C(n_281680317
		), .D(n_281980320), .Z(n_287580376));
	notech_ao4 i_196942620(.A(n_58044), .B(\nbus_11358[3] ), .C(n_123771717)
		, .D(n_59223), .Z(n_287680377));
	notech_ao4 i_196742622(.A(n_60022), .B(n_57470), .C(n_154079044), .D(n_29728
		), .Z(n_287880379));
	notech_and4 i_197142618(.A(n_216676105), .B(n_287880379), .C(n_287680377
		), .D(n_281380314), .Z(n_288080381));
	notech_ao4 i_193942650(.A(n_281966348), .B(n_26807), .C(n_281866347), .D
		(n_229479795), .Z(n_288180382));
	notech_ao4 i_193742652(.A(n_282266351), .B(n_26816), .C(n_282166350), .D
		(n_57139), .Z(n_288380384));
	notech_and4 i_194142648(.A(n_288380384), .B(n_288180382), .C(n_280580306
		), .D(n_280880309), .Z(n_288580386));
	notech_ao4 i_193442655(.A(n_56073), .B(n_57573), .C(n_143471914), .D(n_59205
		), .Z(n_288680387));
	notech_ao4 i_193242657(.A(n_60020), .B(n_301180512), .C(n_153879042), .D
		(n_29651), .Z(n_288880389));
	notech_and4 i_193642653(.A(n_216276101), .B(n_288880389), .C(n_288680387
		), .D(n_280280303), .Z(n_289080391));
	notech_ao4 i_192942660(.A(n_306670077), .B(n_229479795), .C(n_306570076)
		, .D(n_26807), .Z(n_289180392));
	notech_ao4 i_192742662(.A(n_306970080), .B(n_26816), .C(n_306870079), .D
		(n_57139), .Z(n_289380394));
	notech_and4 i_193142658(.A(n_289380394), .B(n_289180392), .C(n_279480295
		), .D(n_279780298), .Z(n_289580396));
	notech_ao4 i_192442665(.A(n_57573), .B(n_55983), .C(n_143471914), .D(n_59223
		), .Z(n_289680397));
	notech_ao4 i_192242667(.A(n_60022), .B(n_301180512), .C(n_29728), .D(n_153879042
		), .Z(n_289880399));
	notech_and4 i_192642663(.A(n_216676105), .B(n_289880399), .C(n_289680397
		), .D(n_279180292), .Z(n_290080401));
	notech_ao4 i_191942670(.A(n_96519147), .B(n_307124335), .C(n_306221226),
		 .D(n_56649), .Z(n_290180402));
	notech_ao4 i_191842671(.A(n_314047718), .B(\nbus_11365[31] ), .C(n_314391680
		), .D(n_147271952), .Z(n_290380404));
	notech_nand3 i_192142668(.A(n_290180402), .B(n_290380404), .C(n_278680287
		), .Z(n_290480405));
	notech_ao4 i_191642673(.A(n_57864), .B(\nbus_11358[31] ), .C(n_58141), .D
		(n_314791676), .Z(n_290580406));
	notech_ao4 i_189442695(.A(n_281966348), .B(n_266380164), .C(n_281866347)
		, .D(n_247579976), .Z(n_290880409));
	notech_ao4 i_189242697(.A(n_282266351), .B(n_58486), .C(n_282166350), .D
		(n_57141), .Z(n_291080411));
	notech_and4 i_189642693(.A(n_291080411), .B(n_290880409), .C(n_277580276
		), .D(n_277880279), .Z(n_291280413));
	notech_ao4 i_188942700(.A(n_56073), .B(n_57154), .C(n_147171951), .D(n_59205
		), .Z(n_291380414));
	notech_ao4 i_188742702(.A(n_60020), .B(n_57084), .C(n_247679977), .D(n_29651
		), .Z(n_291580416));
	notech_and4 i_189142698(.A(n_216276101), .B(n_291580416), .C(n_291380414
		), .D(n_277280273), .Z(n_291780418));
	notech_ao4 i_188442705(.A(n_306670077), .B(n_247579976), .C(n_306570076)
		, .D(n_266380164), .Z(n_291880419));
	notech_ao4 i_188242707(.A(n_306970080), .B(n_58486), .C(n_306870079), .D
		(n_57141), .Z(n_292080421));
	notech_and4 i_188642703(.A(n_292080421), .B(n_291880419), .C(n_276480265
		), .D(n_276780268), .Z(n_292280423));
	notech_ao4 i_187942710(.A(n_57154), .B(n_55983), .C(n_147171951), .D(n_59223
		), .Z(n_292380424));
	notech_ao4 i_187742712(.A(n_60022), .B(n_57084), .C(n_29728), .D(n_247679977
		), .Z(n_292580426));
	notech_and4 i_188142708(.A(n_216676105), .B(n_292580426), .C(n_292380424
		), .D(n_276180262), .Z(n_292780428));
	notech_ao4 i_183642753(.A(n_96519147), .B(n_58085), .C(n_306221226), .D(n_56916
		), .Z(n_292880429));
	notech_ao4 i_183542754(.A(n_57870), .B(\nbus_11365[31] ), .C(n_314391680
		), .D(n_153779041), .Z(n_293080431));
	notech_ao4 i_183242757(.A(n_57877), .B(\nbus_11358[31] ), .C(n_314791676
		), .D(n_58143), .Z(n_293280433));
	notech_and4 i_183442755(.A(n_293280433), .B(n_274880249), .C(n_275180252
		), .D(n_26710), .Z(n_293580436));
	notech_ao4 i_180742782(.A(n_281966348), .B(n_58162), .C(n_281866347), .D
		(n_153379037), .Z(n_293680437));
	notech_ao4 i_180642783(.A(n_282166350), .B(n_257980080), .C(n_282066349)
		, .D(n_153279036), .Z(n_293780438));
	notech_ao4 i_180442785(.A(n_153779041), .B(n_308621250), .C(n_26804), .D
		(n_282266351), .Z(n_293980440));
	notech_and4 i_180942780(.A(n_293980440), .B(n_293780438), .C(n_293680437
		), .D(n_274380244), .Z(n_294180442));
	notech_ao4 i_180142788(.A(n_57583), .B(n_153479038), .C(n_58047), .D(n_56073
		), .Z(n_294280443));
	notech_ao4 i_179842790(.A(n_56356), .B(nbus_11295[5]), .C(n_60020), .D(n_153579039
		), .Z(n_294480445));
	notech_and4 i_180342786(.A(n_216276101), .B(n_294480445), .C(n_294280443
		), .D(n_274080241), .Z(n_294680447));
	notech_ao4 i_179542793(.A(n_306670077), .B(n_153379037), .C(n_306570076)
		, .D(n_58162), .Z(n_294780448));
	notech_ao4 i_179442794(.A(n_306870079), .B(n_257980080), .C(n_306770078)
		, .D(n_153279036), .Z(n_294880449));
	notech_ao4 i_179242796(.A(n_153779041), .B(n_308721251), .C(n_26804), .D
		(n_306970080), .Z(n_295080451));
	notech_and4 i_179742791(.A(n_295080451), .B(n_294880449), .C(n_294780448
		), .D(n_273180232), .Z(n_295280453));
	notech_ao4 i_178942799(.A(n_153479038), .B(n_57563), .C(n_58047), .D(n_55983
		), .Z(n_295380454));
	notech_ao4 i_178742801(.A(n_56356), .B(nbus_11295[3]), .C(n_60022), .D(n_153579039
		), .Z(n_295580456));
	notech_and4 i_179142797(.A(n_216676105), .B(n_295580456), .C(n_295380454
		), .D(n_272880229), .Z(n_295780458));
	notech_ao4 i_176042828(.A(n_281866347), .B(n_303873518), .C(n_282066349)
		, .D(n_303773517), .Z(n_295880459));
	notech_ao4 i_175842830(.A(n_304173521), .B(n_56073), .C(n_60020), .D(n_285080351
		), .Z(n_296080461));
	notech_and4 i_176242826(.A(n_296080461), .B(n_295880459), .C(n_272080221
		), .D(n_272380224), .Z(n_296280463));
	notech_ao4 i_175542833(.A(n_282166350), .B(n_57923), .C(n_281966348), .D
		(n_26906), .Z(n_296380464));
	notech_and4 i_175742831(.A(n_216276101), .B(n_296380464), .C(n_271480215
		), .D(n_271780218), .Z(n_296680467));
	notech_ao4 i_168842900(.A(n_306670077), .B(n_303873518), .C(n_306770078)
		, .D(n_303773517), .Z(n_296780468));
	notech_ao4 i_168642902(.A(n_304173521), .B(n_55983), .C(n_60022), .D(n_285080351
		), .Z(n_296980470));
	notech_and4 i_169042898(.A(n_296980470), .B(n_296780468), .C(n_271080211
		), .D(n_271380214), .Z(n_297180472));
	notech_ao4 i_168342905(.A(n_306870079), .B(n_57923), .C(n_306570076), .D
		(n_26906), .Z(n_297280473));
	notech_and4 i_168542903(.A(n_216676105), .B(n_297280473), .C(n_270480205
		), .D(n_270780208), .Z(n_297580476));
	notech_and2 i_8344411(.A(n_38618568), .B(n_265380154), .Z(n_297680477)
		);
	notech_or2 i_159342994(.A(n_303791786), .B(n_26815), .Z(n_297780478));
	notech_ao4 i_159042997(.A(n_314791676), .B(n_264680147), .C(\nbus_11358[31] 
		), .D(n_297780478), .Z(n_297880479));
	notech_ao4 i_158842999(.A(n_314591678), .B(n_56542), .C(n_83019012), .D(n_264880149
		), .Z(n_298080481));
	notech_and4 i_159242995(.A(n_298080481), .B(n_297880479), .C(n_270080201
		), .D(n_270380204), .Z(n_298280483));
	notech_ao4 i_158443002(.A(n_261280113), .B(n_29619), .C(n_60127), .D(n_27217
		), .Z(n_298380484));
	notech_and2 i_158243003(.A(n_297680477), .B(n_269480195), .Z(n_298580486
		));
	notech_ao4 i_153743047(.A(n_26852), .B(n_264280143), .C(n_26812), .D(n_264180142
		), .Z(n_298780488));
	notech_ao4 i_153643048(.A(n_284680347), .B(n_26802), .C(n_3874), .D(n_284880349
		), .Z(n_298880489));
	notech_ao4 i_153443050(.A(n_92519107), .B(n_178572265), .C(n_56485), .D(n_302621190
		), .Z(n_299080491));
	notech_and3 i_153543049(.A(n_311173591), .B(n_299080491), .C(n_268780188
		), .Z(n_299280493));
	notech_ao4 i_153043054(.A(n_281866347), .B(n_284480345), .C(n_57583), .D
		(n_284380344), .Z(n_299380494));
	notech_ao4 i_152843056(.A(n_284680347), .B(n_282066349), .C(n_60020), .D
		(n_284880349), .Z(n_299580496));
	notech_and4 i_153243052(.A(n_299580496), .B(n_299380494), .C(n_268380184
		), .D(n_268680187), .Z(n_299780498));
	notech_ao4 i_152543059(.A(n_282166350), .B(n_57915), .C(n_281966348), .D
		(n_26852), .Z(n_299880499));
	notech_and4 i_152743057(.A(n_299880499), .B(n_216276101), .C(n_267780178
		), .D(n_268080181), .Z(n_300180502));
	notech_ao4 i_152143063(.A(n_306670077), .B(n_284480345), .C(n_284380344)
		, .D(n_57563), .Z(n_300280503));
	notech_ao4 i_151943065(.A(n_306770078), .B(n_284680347), .C(n_60022), .D
		(n_284880349), .Z(n_300480505));
	notech_and4 i_152343061(.A(n_300480505), .B(n_300280503), .C(n_267380174
		), .D(n_267680177), .Z(n_300680507));
	notech_ao4 i_151643068(.A(n_306870079), .B(n_57915), .C(n_306570076), .D
		(n_26852), .Z(n_300780508));
	notech_and4 i_151843066(.A(n_300780508), .B(n_216676105), .C(n_266780168
		), .D(n_267080171), .Z(n_301080511));
	notech_or4 i_200264473(.A(n_101413114), .B(n_54709), .C(instrc[121]), .D
		(n_26816), .Z(n_301180512));
	notech_and2 i_1841238(.A(n_58646), .B(n_301680517), .Z(n_301280513));
	notech_and2 i_1941237(.A(n_332480825), .B(n_58610), .Z(n_301380514));
	notech_or2 i_61540676(.A(n_318991634), .B(n_59742), .Z(n_301680517));
	notech_mux2 i_2241234(.S(n_32365), .A(n_56037), .B(n_60025), .Z(n_301780518
		));
	notech_ao3 i_62240669(.A(n_32365), .B(opb[0]), .C(n_317391650), .Z(n_302080521
		));
	notech_nand3 i_78940515(.A(n_32393), .B(n_62824), .C(n_26832), .Z(n_302180522
		));
	notech_or4 i_98440338(.A(n_59387), .B(n_59275), .C(n_4011), .D(n_29178),
		 .Z(n_303880539));
	notech_nao3 i_98940333(.A(n_56925), .B(n_318791636), .C(n_4011), .Z(n_304080541
		));
	notech_nao3 i_99040332(.A(n_190062172), .B(n_58171), .C(n_56863), .Z(n_304180542
		));
	notech_nand2 i_5841199(.A(n_58097), .B(opb[8]), .Z(n_304680547));
	notech_nand3 i_5541202(.A(n_27179), .B(n_26941), .C(\opa_12[8] ), .Z(n_304980550
		));
	notech_nao3 i_5241205(.A(n_318791636), .B(n_246991940), .C(n_325270263),
		 .Z(n_305280553));
	notech_or4 i_46640812(.A(n_54954), .B(n_54934), .C(n_5933), .D(n_58020),
		 .Z(n_305580556));
	notech_or2 i_46140815(.A(n_302391800), .B(n_27991), .Z(n_305880559));
	notech_or4 i_45740818(.A(n_26767), .B(n_28134), .C(n_60924), .D(n_54934)
		, .Z(n_306180562));
	notech_or2 i_54440741(.A(n_5933), .B(n_181779321), .Z(n_306280563));
	notech_nand3 i_54340742(.A(n_26813), .B(n_26821), .C(\opa_12[8] ), .Z(n_306580566
		));
	notech_or4 i_53840747(.A(n_54814), .B(n_28134), .C(n_60924), .D(n_58481)
		, .Z(n_307080571));
	notech_or2 i_55440731(.A(n_56356), .B(nbus_11295[8]), .Z(n_307180572));
	notech_nand2 i_55340732(.A(opb[8]), .B(n_58050), .Z(n_307480575));
	notech_or4 i_55040735(.A(n_58132), .B(n_56803), .C(n_5933), .D(n_56903),
		 .Z(n_307780578));
	notech_or4 i_54740738(.A(n_58806), .B(n_28134), .C(n_60926), .D(n_56803)
		, .Z(n_308080581));
	notech_or2 i_57340713(.A(n_5933), .B(n_57025), .Z(n_308180582));
	notech_or2 i_57240714(.A(n_57181), .B(\nbus_11358[8] ), .Z(n_308480585)
		);
	notech_nao3 i_56740719(.A(n_319091633), .B(n_56925), .C(n_325270263), .Z
		(n_308980590));
	notech_or2 i_58340703(.A(n_5933), .B(n_228579786), .Z(n_309080591));
	notech_nand2 i_58240704(.A(opb[8]), .B(n_57179), .Z(n_309380594));
	notech_nand3 i_57940707(.A(n_26828), .B(n_26827), .C(\opa_12[8] ), .Z(n_309680597
		));
	notech_or4 i_57640710(.A(n_54718), .B(n_28134), .C(n_60926), .D(n_58479)
		, .Z(n_309980600));
	notech_or2 i_59240694(.A(n_5933), .B(n_57299), .Z(n_310080601));
	notech_or2 i_59140695(.A(n_57807), .B(\nbus_11358[8] ), .Z(n_310380604)
		);
	notech_nao3 i_58640700(.A(opc_10[8]), .B(n_62814), .C(n_57473), .Z(n_310880609
		));
	notech_or4 i_59540691(.A(n_308891735), .B(n_32382), .C(n_60263), .D(n_29787
		), .Z(n_311380614));
	notech_or4 i_61440677(.A(n_317391650), .B(n_316591658), .C(n_56396), .D(n_56028
		), .Z(n_311680617));
	notech_nand2 i_60840680(.A(sav_epc[0]), .B(n_61145), .Z(n_311980620));
	notech_or2 i_60440683(.A(n_58406), .B(n_59187), .Z(n_312280623));
	notech_ao4 i_60040686(.A(n_26818), .B(n_26817), .C(n_302080521), .D(n_26830
		), .Z(n_312580626));
	notech_nao3 i_67840626(.A(n_11411), .B(n_32272), .C(n_2868), .Z(n_313280633
		));
	notech_nand2 i_67540629(.A(sav_epc[8]), .B(n_61145), .Z(n_313580636));
	notech_or4 i_67240632(.A(n_62860), .B(n_62814), .C(n_29787), .D(n_316891655
		), .Z(n_313880639));
	notech_nao3 i_70740597(.A(n_11412), .B(n_32272), .C(n_2868), .Z(n_314580646
		));
	notech_nand2 i_70440600(.A(sav_epc[9]), .B(n_61143), .Z(n_314880649));
	notech_or4 i_70140603(.A(n_62860), .B(n_62814), .C(n_29743), .D(n_316891655
		), .Z(n_315180652));
	notech_nao3 i_72040584(.A(n_11413), .B(n_32272), .C(n_2868), .Z(n_315880659
		));
	notech_nand2 i_71740587(.A(sav_epc[10]), .B(n_61143), .Z(n_316180662));
	notech_or4 i_71440590(.A(n_62856), .B(n_62814), .C(n_56145), .D(n_316891655
		), .Z(n_316480665));
	notech_nao3 i_73440570(.A(n_11414), .B(n_32272), .C(n_2868), .Z(n_317180672
		));
	notech_nand2 i_72740577(.A(opa[11]), .B(n_290918108), .Z(n_317880679));
	notech_nao3 i_76140543(.A(n_11416), .B(n_32272), .C(n_2868), .Z(n_318580686
		));
	notech_nand2 i_75440550(.A(opa[13]), .B(n_290918108), .Z(n_319280693));
	notech_nao3 i_77540529(.A(n_11417), .B(n_32272), .C(n_2868), .Z(n_319980700
		));
	notech_nand2 i_76840536(.A(opa[14]), .B(n_290918108), .Z(n_320680707));
	notech_nao3 i_78840516(.A(n_11418), .B(n_32272), .C(n_2868), .Z(n_321380714
		));
	notech_nand2 i_78540519(.A(sav_epc[15]), .B(n_61143), .Z(n_321680717));
	notech_or4 i_78240522(.A(n_62860), .B(n_62814), .C(n_56266), .D(n_316891655
		), .Z(n_321980720));
	notech_nand2 i_34056(.A(n_27029), .B(n_26669), .Z(n_322480725));
	notech_or4 i_30907(.A(n_57020), .B(n_56863), .C(n_57033), .D(n_56803), .Z
		(n_322580726));
	notech_nand2 i_30904(.A(n_26825), .B(n_26824), .Z(n_322680727));
	notech_or4 i_29841(.A(n_54727), .B(n_57078), .C(n_57064), .D(n_58479), .Z
		(n_322780728));
	notech_nao3 i_29840(.A(n_62826), .B(n_26826), .C(n_54718), .Z(n_322880729
		));
	notech_nand2 i_29834(.A(n_26828), .B(n_26827), .Z(n_322980730));
	notech_nao3 i_29833(.A(n_30945), .B(n_56471), .C(n_54727), .Z(n_323080731
		));
	notech_or2 i_29369(.A(n_54678), .B(n_57505), .Z(n_323180732));
	notech_or4 i_14164(.A(n_101413114), .B(n_54709), .C(n_58503), .D(instrc[
		121]), .Z(n_323280733));
	notech_and4 i_32441306(.A(n_57020), .B(n_30945), .C(instrc[119]), .D(n_62814
		), .Z(n_323480735));
	notech_nand2 i_154341253(.A(n_27196), .B(n_26818), .Z(n_323580736));
	notech_nand3 i_151541254(.A(n_246591944), .B(n_57051), .C(n_26818), .Z(n_323680737
		));
	notech_ao4 i_181739573(.A(n_298466513), .B(n_323680737), .C(n_56266), .D
		(n_323580736), .Z(n_323780738));
	notech_ao4 i_181639574(.A(n_290818107), .B(nbus_11295[15]), .C(n_290718106
		), .D(n_56275), .Z(n_323880739));
	notech_ao4 i_181439576(.A(n_28000), .B(n_291718116), .C(\nbus_11307[15] 
		), .D(n_26857), .Z(n_324180742));
	notech_and4 i_181939571(.A(n_324180742), .B(n_323880739), .C(n_323780738
		), .D(n_321980720), .Z(n_324380744));
	notech_ao4 i_181139579(.A(n_315591668), .B(n_59962), .C(n_122628503), .D
		(n_29552), .Z(n_324480745));
	notech_ao4 i_180939581(.A(n_309291731), .B(n_28104), .C(n_60010), .D(n_316791656
		), .Z(n_324680747));
	notech_and4 i_181339577(.A(n_321380714), .B(n_324680747), .C(n_324480745
		), .D(n_321680717), .Z(n_324880749));
	notech_or2 i_206141244(.A(n_32393), .B(n_316891655), .Z(n_324980750));
	notech_nand3 i_205841245(.A(n_56396), .B(n_27194), .C(n_26818), .Z(n_325180752
		));
	notech_ao4 i_180339586(.A(n_56257), .B(n_325180752), .C(n_298366512), .D
		(n_324980750), .Z(n_325280753));
	notech_ao4 i_180239587(.A(n_298266511), .B(n_323680737), .C(n_60011), .D
		(n_316791656), .Z(n_325580756));
	notech_ao4 i_180039589(.A(n_290818107), .B(nbus_11295[14]), .C(n_290718106
		), .D(\nbus_11358[14] ), .Z(n_325780758));
	notech_and4 i_180639584(.A(n_325780758), .B(n_325580756), .C(n_325280753
		), .D(n_320680707), .Z(n_325980760));
	notech_ao4 i_179739592(.A(n_298166510), .B(n_316891655), .C(n_291718116)
		, .D(n_27999), .Z(n_326080761));
	notech_ao4 i_179639593(.A(n_315591668), .B(n_59963), .C(n_122628503), .D
		(n_29551), .Z(n_326180762));
	notech_ao4 i_179439595(.A(n_309291731), .B(n_28103), .C(n_60127), .D(n_27255
		), .Z(n_326380764));
	notech_and4 i_179939590(.A(n_326380764), .B(n_326180762), .C(n_326080761
		), .D(n_319980700), .Z(n_326580766));
	notech_ao4 i_179139598(.A(n_325180752), .B(n_56239), .C(n_31576), .D(n_324980750
		), .Z(n_326680767));
	notech_ao4 i_179039599(.A(n_31560), .B(n_323680737), .C(n_302091803), .D
		(n_316791656), .Z(n_326780768));
	notech_ao4 i_178839601(.A(nbus_11295[13]), .B(n_290818107), .C(\nbus_11358[13] 
		), .D(n_290718106), .Z(n_326980770));
	notech_and4 i_179339596(.A(n_326980770), .B(n_326780768), .C(n_326680767
		), .D(n_319280693), .Z(n_327180772));
	notech_ao4 i_178539604(.A(n_122628503), .B(n_29550), .C(n_291718116), .D
		(n_27998), .Z(n_327280773));
	notech_ao4 i_178439605(.A(n_301691807), .B(n_315591668), .C(n_316891655)
		, .D(n_31540), .Z(n_327380774));
	notech_ao4 i_178239607(.A(n_309291731), .B(n_28102), .C(n_60127), .D(n_27254
		), .Z(n_327580776));
	notech_and4 i_178739602(.A(n_327580776), .B(n_327380774), .C(n_327280773
		), .D(n_318580686), .Z(n_327780778));
	notech_ao4 i_176739621(.A(n_325180752), .B(n_56190), .C(n_31492), .D(n_324980750
		), .Z(n_327880779));
	notech_ao4 i_176539622(.A(n_31476), .B(n_323680737), .C(n_302491799), .D
		(n_316791656), .Z(n_327980780));
	notech_ao4 i_176339624(.A(n_290818107), .B(nbus_11295[11]), .C(n_290718106
		), .D(n_56181), .Z(n_328180782));
	notech_and4 i_177039619(.A(n_328180782), .B(n_327980780), .C(n_327880779
		), .D(n_317880679), .Z(n_328380784));
	notech_ao4 i_176039627(.A(n_31456), .B(n_316891655), .C(n_291718116), .D
		(n_27996), .Z(n_328480785));
	notech_ao4 i_175939628(.A(n_302891795), .B(n_315591668), .C(n_122628503)
		, .D(n_29548), .Z(n_328580786));
	notech_ao4 i_175739630(.A(n_309291731), .B(n_28100), .C(n_60127), .D(n_27253
		), .Z(n_328780788));
	notech_and4 i_176239625(.A(n_328780788), .B(n_328580786), .C(n_328480785
		), .D(n_317180672), .Z(n_328980790));
	notech_ao4 i_175439633(.A(n_31433), .B(n_323680737), .C(n_323580736), .D
		(n_29684), .Z(n_329080791));
	notech_ao4 i_175339634(.A(n_290818107), .B(nbus_11295[10]), .C(n_290718106
		), .D(n_56154), .Z(n_329180792));
	notech_ao4 i_175139636(.A(n_291718116), .B(n_27993), .C(n_57625), .D(n_26857
		), .Z(n_329380794));
	notech_and4 i_175639631(.A(n_329380794), .B(n_329180792), .C(n_329080791
		), .D(n_316480665), .Z(n_329580796));
	notech_ao4 i_174839639(.A(n_3851), .B(n_315591668), .C(n_122628503), .D(n_29547
		), .Z(n_329680797));
	notech_ao4 i_174639641(.A(n_309291731), .B(n_28099), .C(n_3850), .D(n_316791656
		), .Z(n_329880799));
	notech_and4 i_175039637(.A(n_315880659), .B(n_329880799), .C(n_329680797
		), .D(n_316180662), .Z(n_330080801));
	notech_ao4 i_174339644(.A(n_291963186), .B(n_323680737), .C(n_323580736)
		, .D(n_56127), .Z(n_330180802));
	notech_ao4 i_174239645(.A(n_290818107), .B(nbus_11295[9]), .C(n_290718106
		), .D(n_56136), .Z(n_330280803));
	notech_ao4 i_174039647(.A(n_291718116), .B(n_27992), .C(n_57613), .D(n_26857
		), .Z(n_330480805));
	notech_and4 i_174539642(.A(n_330480805), .B(n_330280803), .C(n_330180802
		), .D(n_315180652), .Z(n_330680807));
	notech_ao4 i_173739650(.A(n_315591668), .B(n_59968), .C(n_122628503), .D
		(n_29546), .Z(n_330780808));
	notech_ao4 i_173539652(.A(n_309291731), .B(n_28098), .C(n_60016), .D(n_316791656
		), .Z(n_330980810));
	notech_and4 i_173939648(.A(n_314580646), .B(n_330980810), .C(n_330780808
		), .D(n_314880649), .Z(n_331180812));
	notech_ao4 i_171839669(.A(n_308066609), .B(n_323680737), .C(n_323580736)
		, .D(n_29787), .Z(n_331280813));
	notech_ao4 i_171739670(.A(n_290818107), .B(nbus_11295[8]), .C(n_290718106
		), .D(\nbus_11358[8] ), .Z(n_331380814));
	notech_ao4 i_171539672(.A(n_291718116), .B(n_27991), .C(\nbus_11307[8] )
		, .D(n_26857), .Z(n_331580816));
	notech_and4 i_172039667(.A(n_331580816), .B(n_331380814), .C(n_331280813
		), .D(n_313880639), .Z(n_331780818));
	notech_ao4 i_171239675(.A(n_122628503), .B(n_29545), .C(n_315591668), .D
		(n_293018129), .Z(n_331880819));
	notech_ao4 i_171039677(.A(n_309291731), .B(n_28097), .C(n_5933), .D(n_316791656
		), .Z(n_332080821));
	notech_and4 i_171439673(.A(n_313280633), .B(n_332080821), .C(n_331880819
		), .D(n_313580636), .Z(n_332280823));
	notech_ao4 i_168239705(.A(n_32309), .B(nbus_11295[0]), .C(n_315891665), 
		.D(n_59742), .Z(n_332380824));
	notech_ao4 i_168339704(.A(n_32393), .B(n_291363180), .C(n_317391650), .D
		(n_301780518), .Z(n_332480825));
	notech_ao4 i_167839708(.A(n_317091653), .B(n_301380514), .C(n_316591658)
		, .D(n_301280513), .Z(n_332580826));
	notech_ao4 i_167639710(.A(n_309391730), .B(n_291263179), .C(n_286163128)
		, .D(n_291163178), .Z(n_332780828));
	notech_and4 i_168139706(.A(n_332780828), .B(n_332580826), .C(n_312280623
		), .D(n_26831), .Z(n_332980830));
	notech_ao4 i_167339713(.A(n_317991644), .B(n_59993), .C(n_122628503), .D
		(n_29538), .Z(n_333080831));
	notech_ao4 i_166939715(.A(n_56091), .B(n_30032), .C(n_309291731), .D(n_28089
		), .Z(n_333280833));
	notech_and4 i_167539711(.A(n_333280833), .B(n_333080831), .C(n_311680617
		), .D(n_311980620), .Z(n_333480835));
	notech_ao4 i_166339721(.A(n_54678), .B(n_308166610), .C(n_325270263), .D
		(n_56636), .Z(n_333580836));
	notech_ao4 i_166239722(.A(n_58376), .B(n_27991), .C(n_29787), .D(n_323180732
		), .Z(n_333780838));
	notech_ao4 i_165939725(.A(nbus_11295[8]), .B(n_26823), .C(n_57809), .D(\nbus_11307[8] 
		), .Z(n_333980840));
	notech_ao4 i_166739717(.A(n_30569), .B(\nbus_11358[8] ), .C(n_30568), .D
		(\nbus_11307[8] ), .Z(n_334180842));
	notech_ao4 i_166639718(.A(n_30565), .B(n_5933), .C(n_60303), .D(n_28097)
		, .Z(n_334380844));
	notech_and3 i_65941274(.A(n_334180842), .B(n_334380844), .C(n_311380614)
		, .Z(n_334480845));
	notech_and4 i_166139723(.A(n_334480845), .B(n_310080601), .C(n_333980840
		), .D(n_310380604), .Z(n_334680847));
	notech_ao4 i_165539729(.A(n_308166610), .B(n_58479), .C(n_325270263), .D
		(n_56662), .Z(n_334780848));
	notech_ao4 i_165339731(.A(n_322880729), .B(nbus_11295[8]), .C(n_309666625
		), .D(n_323080731), .Z(n_334980850));
	notech_and4 i_165739727(.A(n_334980850), .B(n_309980600), .C(n_334780848
		), .D(n_309680597), .Z(n_335180852));
	notech_ao4 i_165039734(.A(\nbus_11307[8] ), .B(n_26856), .C(n_58375), .D
		(n_27991), .Z(n_335280853));
	notech_and4 i_165239732(.A(n_334480845), .B(n_309080591), .C(n_335280853
		), .D(n_309380594), .Z(n_335580856));
	notech_ao4 i_164639738(.A(n_57604), .B(n_26607), .C(n_309666625), .D(n_313270143
		), .Z(n_335680857));
	notech_ao4 i_164539739(.A(n_308066609), .B(n_319870209), .C(n_308166610)
		, .D(n_54736), .Z(n_335880859));
	notech_ao4 i_164239742(.A(n_58374), .B(n_27991), .C(n_319970210), .D(n_29787
		), .Z(n_336080861));
	notech_and4 i_164439740(.A(n_334480845), .B(n_308180582), .C(n_336080861
		), .D(n_308480585), .Z(n_336380864));
	notech_ao4 i_163039754(.A(n_308166610), .B(n_58477), .C(n_325270263), .D
		(n_56916), .Z(n_336480865));
	notech_ao4 i_162839756(.A(n_322680727), .B(n_29787), .C(n_309666625), .D
		(n_58041), .Z(n_336680867));
	notech_and4 i_163239752(.A(n_307780578), .B(n_336680867), .C(n_308080581
		), .D(n_336480865), .Z(n_336880869));
	notech_ao4 i_162539759(.A(n_57604), .B(n_26854), .C(n_58372), .D(n_27991
		), .Z(n_336980870));
	notech_and4 i_162739757(.A(n_334480845), .B(n_336980870), .C(n_307180572
		), .D(n_307480575), .Z(n_337280873));
	notech_ao4 i_162139763(.A(n_308166610), .B(n_58481), .C(n_325270263), .D
		(n_56498), .Z(n_337380874));
	notech_ao4 i_162039764(.A(n_57604), .B(n_26851), .C(n_309666625), .D(n_58038
		), .Z(n_337580876));
	notech_ao4 i_161739767(.A(n_58052), .B(n_56118), .C(n_27991), .D(n_26850
		), .Z(n_337780878));
	notech_and4 i_161939765(.A(n_334480845), .B(n_306280563), .C(n_337780878
		), .D(n_306580566), .Z(n_338080881));
	notech_ao4 i_148839890(.A(n_308166610), .B(n_54934), .C(n_325270263), .D
		(n_56601), .Z(n_338180882));
	notech_ao4 i_148639892(.A(n_322480725), .B(n_29787), .C(n_309666625), .D
		(n_301991804), .Z(n_338380884));
	notech_and4 i_149039888(.A(n_338380884), .B(n_306180562), .C(n_338180882
		), .D(n_305880559), .Z(n_338580886));
	notech_ao4 i_148339895(.A(n_302291801), .B(n_56118), .C(n_57604), .D(n_27293
		), .Z(n_338680887));
	notech_and4 i_148539893(.A(n_54667), .B(n_334480845), .C(n_305580556), .D
		(n_338680887), .Z(n_338980890));
	notech_ao4 i_104440289(.A(n_309666625), .B(n_312970140), .C(n_54638), .D
		(n_28950), .Z(n_339080891));
	notech_ao4 i_104240291(.A(n_308066609), .B(n_319670207), .C(n_308166610)
		, .D(n_23512), .Z(n_339280893));
	notech_and4 i_104640287(.A(n_339280893), .B(n_339080891), .C(n_304980550
		), .D(n_305280553), .Z(n_339480895));
	notech_ao4 i_103940294(.A(n_26819), .B(n_57604), .C(n_58408), .D(n_27991
		), .Z(n_339580896));
	notech_ao4 i_103740296(.A(n_59124), .B(nbus_11295[8]), .C(n_5933), .D(n_316691657
		), .Z(n_339780898));
	notech_and4 i_104140292(.A(n_339780898), .B(n_339580896), .C(n_334480845
		), .D(n_304680547), .Z(n_339980900));
	notech_or2 i_136532765(.A(instrc[126]), .B(instrc[125]), .Z(n_340380904)
		);
	notech_nand2 i_102432705(.A(instrc[126]), .B(instrc[127]), .Z(n_340480905
		));
	notech_nand3 i_160832699(.A(n_56888), .B(n_3751), .C(n_29628), .Z(n_340580906
		));
	notech_ao4 i_9532644(.A(n_317591648), .B(n_60841), .C(n_347280973), .D(n_26898
		), .Z(n_341080911));
	notech_and4 i_32832462(.A(n_30905), .B(n_3828), .C(n_3829), .D(n_27035),
		 .Z(n_341180912));
	notech_and2 i_32932461(.A(n_347380974), .B(n_27034), .Z(n_341280913));
	notech_ao4 i_26832509(.A(n_60964), .B(n_60953), .C(n_26991), .D(n_26837)
		, .Z(n_341380914));
	notech_and2 i_67832160(.A(n_3835), .B(n_341780918), .Z(n_341680917));
	notech_nand2 i_24832526(.A(n_58088), .B(n_27641), .Z(n_341780918));
	notech_or4 i_68032158(.A(n_3730), .B(instrc[122]), .C(n_32334), .D(n_26894
		), .Z(n_341880919));
	notech_nand2 i_51032317(.A(sav_epc[30]), .B(n_61143), .Z(n_342180922));
	notech_nand2 i_50732320(.A(n_122228499), .B(\regs_13_14[30] ), .Z(n_342480925
		));
	notech_or2 i_50332323(.A(n_121628493), .B(n_28015), .Z(n_342780928));
	notech_nao3 i_50032326(.A(n_11433), .B(n_32272), .C(n_2868), .Z(n_343080931
		));
	notech_nand2 i_29685(.A(instrc[127]), .B(n_3813), .Z(n_343180932));
	notech_nao3 i_66532170(.A(n_29640), .B(n_29631), .C(n_344680947), .Z(n_343780938
		));
	notech_or2 i_66232173(.A(n_26888), .B(n_344880949), .Z(n_344080941));
	notech_or4 i_65732178(.A(n_26887), .B(n_26894), .C(instrc[98]), .D(n_340580906
		), .Z(n_344180942));
	notech_or4 i_65832177(.A(n_57462), .B(instrc[100]), .C(instrc[103]), .D(n_6588872
		), .Z(n_344280943));
	notech_or4 i_65932176(.A(n_57064), .B(n_345480955), .C(instrc[119]), .D(n_57078
		), .Z(n_344380944));
	notech_ao4 i_35200(.A(n_61117), .B(n_341680917), .C(n_32263), .D(n_59469
		), .Z(n_344480945));
	notech_nand2 i_31088(.A(n_58122), .B(n_29179), .Z(n_344580946));
	notech_or4 i_31406(.A(n_6368850), .B(instrc[88]), .C(n_314663413), .D(instrc
		[90]), .Z(n_344680947));
	notech_or4 i_31089(.A(n_57369), .B(instrc[105]), .C(n_26894), .D(n_26728
		), .Z(n_344880949));
	notech_nor2 i_31081(.A(n_340380904), .B(n_32747), .Z(n_345280953));
	notech_or4 i_30346(.A(n_30359), .B(n_30344), .C(n_57020), .D(n_314663413
		), .Z(n_345480955));
	notech_nor2 i_30345(.A(n_30344), .B(n_57020), .Z(n_345580956));
	notech_nand3 i_98832881(.A(instrc[127]), .B(n_3830), .C(instrc[124]), .Z
		(n_345680957));
	notech_or2 i_29650(.A(n_345880959), .B(n_29641), .Z(n_345780958));
	notech_nao3 i_29649(.A(instrc[99]), .B(n_26858), .C(n_30359), .Z(n_345880959
		));
	notech_nand2 i_29664(.A(n_27031), .B(n_29179), .Z(n_345980960));
	notech_nand2 i_29665(.A(n_29631), .B(instrc[91]), .Z(n_346080961));
	notech_or4 i_29676(.A(instrc[105]), .B(n_26728), .C(n_26894), .D(n_29736
		), .Z(n_346180962));
	notech_or4 i_29605(.A(n_61143), .B(n_60303), .C(n_26900), .D(n_29638), .Z
		(n_346280963));
	notech_and3 i_121931663(.A(n_344180942), .B(n_344380944), .C(n_344280943
		), .Z(n_347180972));
	notech_or4 i_124531638(.A(instrc[126]), .B(instrc[125]), .C(n_316191662)
		, .D(n_32747), .Z(n_347280973));
	notech_ao4 i_124231641(.A(n_30905), .B(n_60926), .C(n_32408), .D(n_26839
		), .Z(n_347380974));
	notech_ao4 i_121631666(.A(n_26942), .B(n_341280913), .C(n_341180912), .D
		(n_341080911), .Z(n_347480975));
	notech_ao4 i_121331669(.A(n_26959), .B(n_40675), .C(n_56579), .D(n_3829)
		, .Z(n_347780978));
	notech_ao4 i_121131671(.A(n_32343), .B(n_344580946), .C(n_26956), .D(n_340380904
		), .Z(n_348180982));
	notech_and4 i_121531667(.A(n_344480945), .B(n_348180982), .C(n_343780938
		), .D(n_347780978), .Z(n_348380984));
	notech_ao4 i_93931925(.A(n_309291731), .B(n_28121), .C(n_309391730), .D(n_32252
		), .Z(n_348480985));
	notech_ao4 i_93731927(.A(n_308991734), .B(n_57828), .C(n_309091733), .D(\nbus_11358[30] 
		), .Z(n_348680987));
	notech_and4 i_94131923(.A(n_348680987), .B(n_348480985), .C(n_342780928)
		, .D(n_343080931), .Z(n_348880989));
	notech_ao4 i_93431930(.A(n_124328520), .B(n_303091793), .C(n_122628503),
		 .D(n_29554), .Z(n_348980990));
	notech_ao4 i_93231932(.A(n_122528502), .B(n_302991794), .C(n_122428501),
		 .D(n_28156), .Z(n_349180992));
	notech_and4 i_93631928(.A(n_349180992), .B(n_348980990), .C(n_342180922)
		, .D(n_342480925), .Z(n_349380994));
	notech_nand2 i_117878(.A(n_114078644), .B(n_113978643), .Z(write_data_25
		[0]));
	notech_or4 i_179462709(.A(n_3730), .B(instrc[122]), .C(n_32334), .D(n_29179
		), .Z(n_142261705));
	notech_or4 i_179162712(.A(n_139361676), .B(n_139461677), .C(n_139261675)
		, .D(n_139561678), .Z(n_142161704));
	notech_ao3 i_33867441(.A(n_1874), .B(n_19086), .C(n_32476), .Z(n_349480995
		));
	notech_or2 i_173067438(.A(n_118078684), .B(n_127078774), .Z(n_349580996)
		);
	notech_and4 i_173167437(.A(n_127278776), .B(n_127178775), .C(n_118778691
		), .D(n_118478688), .Z(n_349680997100234));
	notech_or4 i_39079(.A(n_29737), .B(n_57369), .C(n_29734), .D(instrc[104]
		), .Z(n_349780998));
	notech_or4 i_39081(.A(instrc[105]), .B(n_29736), .C(n_114178645), .D(n_30937
		), .Z(n_349880999));
	notech_nand2 i_39085(.A(n_3914), .B(n_114278646), .Z(n_349981000));
	notech_nand2 i_162332766(.A(n_29635), .B(n_29665), .Z(n_57462));
	notech_nand2 i_33336(.A(n_29640), .B(n_29631), .Z(n_190010112));
	notech_xor2 i_110938300(.A(n_28049), .B(opz[1]), .Z(n_57940));
	notech_or4 i_55262(.A(n_26736), .B(n_158179085), .C(n_161479118), .D(n_26740
		), .Z(\nbus_11373[0] ));
	notech_or4 i_55009(.A(n_157479078), .B(n_162579129), .C(n_26741), .D(n_26742
		), .Z(\nbus_11372[0] ));
	notech_or4 i_51972(.A(n_156279066), .B(n_164079144), .C(n_26743), .D(n_26744
		), .Z(\nbus_11335[0] ));
	notech_and4 i_51718(.A(n_165579159), .B(n_166279166), .C(n_155179055), .D
		(n_165479158), .Z(\nbus_11334[0] ));
	notech_and4 i_85564499(.A(n_56843), .B(n_56803), .C(n_125961542), .D(n_58493
		), .Z(n_58162));
	notech_and2 i_100264496(.A(n_57877), .B(n_133278836), .Z(n_58047));
	notech_and3 i_122264488(.A(n_56843), .B(n_125961542), .C(n_56803), .Z(n_57827
		));
	notech_and4 i_1620773(.A(n_166679170), .B(n_166879172), .C(n_167379177),
		 .D(n_153079034), .Z(n_24520));
	notech_nand2 i_520762(.A(n_168279186), .B(n_167879182), .Z(n_24454));
	notech_nand2 i_220759(.A(n_169179195), .B(n_168779191), .Z(n_24436));
	notech_and4 i_120758(.A(n_169779201), .B(n_169679200), .C(n_152275466), 
		.D(n_149478998), .Z(n_24430));
	notech_nand2 i_1020863(.A(n_170879212), .B(n_170479208), .Z(n_24136));
	notech_nand2 i_520858(.A(n_171879222), .B(n_171379217), .Z(n_24106));
	notech_nand2 i_220855(.A(n_172879232), .B(n_172379227), .Z(n_24088));
	notech_nand2 i_520986(.A(n_173879242), .B(n_173379237), .Z(n_23758));
	notech_and4 i_1021087(.A(n_173979243), .B(n_174179245), .C(n_174679250),
		 .D(n_145078954), .Z(n_18883));
	notech_nand2 i_521082(.A(n_175679260), .B(n_175179255), .Z(n_18853));
	notech_nand2 i_221079(.A(n_176679270), .B(n_176179265), .Z(n_18835));
	notech_and4 i_1021183(.A(n_176779271), .B(n_176979273), .C(n_177479278),
		 .D(n_141978923), .Z(n_18534));
	notech_nand2 i_521178(.A(n_178479288), .B(n_177979283), .Z(n_18504));
	notech_nand2 i_221175(.A(n_179479298), .B(n_178979293), .Z(n_18486));
	notech_nand2 i_521626(.A(n_180479308), .B(n_179979303), .Z(n_17804));
	notech_nand2 i_221623(.A(n_181479318), .B(n_180979313), .Z(n_17786));
	notech_ao4 i_2064433(.A(n_59992), .B(n_56675), .C(n_26810), .D(n_59241),
		 .Z(n_253640554));
	notech_or4 i_2764426(.A(n_32579), .B(n_32567), .C(n_60303), .D(n_30361),
		 .Z(n_252940547));
	notech_and2 i_5464399(.A(n_57470), .B(n_132978833), .Z(n_250240520));
	notech_ao4 i_5564398(.A(n_59441), .B(n_26829), .C(n_254240560), .D(n_26808
		), .Z(n_250140519));
	notech_or4 i_178362720(.A(n_138661669), .B(n_26980), .C(n_138761670), .D
		(n_26979), .Z(n_141261695));
	notech_ao4 i_178062723(.A(n_129361576), .B(n_54794), .C(instrc[126]), .D
		(n_141061693), .Z(n_141161694));
	notech_nao3 i_180362700(.A(instrc[125]), .B(n_29632), .C(n_343180932), .Z
		(n_141061693));
	notech_or2 i_4064413(.A(n_175162034), .B(n_32319), .Z(n_140661689));
	notech_or4 i_180862695(.A(n_3812), .B(n_18981), .C(n_19057), .D(n_3807),
		 .Z(n_140461687));
	notech_and3 i_30713(.A(instrc[99]), .B(n_29667), .C(instrc[97]), .Z(n_139861681
		));
	notech_nand2 i_64061830(.A(n_321438009), .B(n_182379327), .Z(n_58377));
	notech_ao4 i_99661823(.A(n_59441), .B(n_26813), .C(n_58172), .D(n_26921)
		, .Z(n_58053));
	notech_and2 i_99761822(.A(n_57873), .B(n_58192), .Z(n_58052));
	notech_and2 i_101161821(.A(n_58082), .B(n_182279326), .Z(n_58038));
	notech_and4 i_105063430(.A(n_57051), .B(instrc[119]), .C(n_57078), .D(n_345580956
		), .Z(n_139561678));
	notech_and4 i_104963431(.A(n_30366), .B(n_29634), .C(instrc[95]), .D(n_76238782
		), .Z(n_139461677));
	notech_and4 i_105263428(.A(n_56888), .B(n_3751), .C(n_29641), .D(n_139861681
		), .Z(n_139361676));
	notech_and4 i_3120788(.A(n_197579476), .B(n_197779478), .C(n_197179472),
		 .D(n_198279483), .Z(n_24610));
	notech_nand2 i_1420771(.A(n_199179492), .B(n_198779488), .Z(n_24508));
	notech_nand2 i_1620869(.A(n_200079501), .B(n_199679497), .Z(n_24172));
	notech_nand2 i_1420867(.A(n_201079511), .B(n_200579506), .Z(n_24160));
	notech_and4 i_1620997(.A(n_201179512), .B(n_201379514), .C(n_201879519),
		 .D(n_192979432), .Z(n_23824));
	notech_nand2 i_1420995(.A(n_202779528), .B(n_202379524), .Z(n_23812));
	notech_nand2 i_1621093(.A(n_203679537), .B(n_203279533), .Z(n_18919));
	notech_nand2 i_1421091(.A(n_204679547), .B(n_204179542), .Z(n_18907));
	notech_and4 i_1621189(.A(n_204779548), .B(n_204979550), .C(n_205479555),
		 .D(n_188879392), .Z(n_18570));
	notech_nand2 i_1421187(.A(n_206379564), .B(n_205979560), .Z(n_18558));
	notech_and4 i_3121876(.A(n_206479565), .B(n_206679567), .C(n_207179572),
		 .D(n_186979373), .Z(n_20798));
	notech_and4 i_1621861(.A(n_207279573), .B(n_207479575), .C(n_207979580),
		 .D(n_186179365), .Z(n_20708));
	notech_and4 i_3121940(.A(n_208579586), .B(n_208779588), .C(n_208479585),
		 .D(n_184679350), .Z(n_17612));
	notech_or4 i_3117620(.A(n_117868195), .B(n_183479338), .C(n_209579596), 
		.D(n_26764), .Z(n_16886));
	notech_nand2 i_1417603(.A(n_210779608), .B(n_210379604), .Z(n_16784));
	notech_and4 i_105163429(.A(instrc[105]), .B(n_30301), .C(n_29736), .D(n_26844
		), .Z(n_139261675));
	notech_nand2 i_1220769(.A(n_230879809), .B(n_230479805), .Z(n_24496));
	notech_and4 i_1120768(.A(n_230979810), .B(n_231179812), .C(n_231679817),
		 .D(n_227179772), .Z(n_24490));
	notech_nand2 i_1220865(.A(n_232679827), .B(n_232179822), .Z(n_24148));
	notech_nand2 i_1120864(.A(n_233579836), .B(n_233179832), .Z(n_24142));
	notech_and4 i_120854(.A(n_233879839), .B(n_234079841), .C(n_234579846), 
		.D(n_26772), .Z(n_24082));
	notech_nand2 i_1220993(.A(n_235479855), .B(n_235079851), .Z(n_23800));
	notech_and4 i_1120992(.A(n_235579856), .B(n_235779858), .C(n_236279863),
		 .D(n_222079721), .Z(n_23794));
	notech_and4 i_120982(.A(n_236579866), .B(n_236779868), .C(n_220879709), 
		.D(n_237279873), .Z(n_23734));
	notech_nand2 i_1221089(.A(n_238279883), .B(n_237779878), .Z(n_18895));
	notech_nand2 i_1121088(.A(n_239179892), .B(n_238779888), .Z(n_18889));
	notech_nand2 i_1221185(.A(n_240079901), .B(n_239679897), .Z(n_18546));
	notech_and4 i_1121184(.A(n_240179902), .B(n_240379904), .C(n_240879909),
		 .D(n_216879669), .Z(n_18540));
	notech_and4 i_121622(.A(n_215679657), .B(n_241179912), .C(n_241779918), 
		.D(n_241079911), .Z(n_17780));
	notech_nand2 i_1221857(.A(n_242679927), .B(n_242279923), .Z(n_20684));
	notech_nand2 i_1121856(.A(n_243579936), .B(n_243179932), .Z(n_20678));
	notech_and4 i_1021855(.A(n_243679937), .B(n_243879939), .C(n_244379944),
		 .D(n_213079631), .Z(n_20672));
	notech_and4 i_105663424(.A(n_30973), .B(n_29668), .C(n_29642), .D(n_3811
		), .Z(n_138961672));
	notech_ao3 i_105563425(.A(n_29665), .B(n_29633), .C(n_29256), .Z(n_138861671
		));
	notech_ao3 i_104063440(.A(instrc[121]), .B(n_32367), .C(n_58692), .Z(n_138761670
		));
	notech_and4 i_103963441(.A(n_62868), .B(n_76638786), .C(n_129261575), .D
		(n_26849), .Z(n_138661669));
	notech_or4 i_103863442(.A(n_27068), .B(n_32476), .C(n_140461687), .D(n_29655
		), .Z(n_138561668));
	notech_nand2 i_220983(.A(n_248679987), .B(n_248179982), .Z(n_23740));
	notech_and4 i_121078(.A(n_186962151), .B(n_249679997), .C(n_249479995), 
		.D(n_249379994), .Z(n_18829));
	notech_and4 i_2420781(.A(n_254180042), .B(n_254380044), .C(n_254880049),
		 .D(n_254080041), .Z(n_24568));
	notech_or4 i_2520878(.A(n_257669588), .B(n_252480025), .C(n_255280053), 
		.D(n_26794), .Z(n_24226));
	notech_or4 i_2320876(.A(n_258469596), .B(n_251680017), .C(n_255980060), 
		.D(n_26795), .Z(n_24214));
	notech_or4 i_2321644(.A(n_258469596), .B(n_250880009), .C(n_256680067), 
		.D(n_26797), .Z(n_17912));
	notech_or4 i_2517614(.A(n_249879999), .B(n_257669588), .C(n_257680077), 
		.D(n_26798), .Z(n_16850));
	notech_and2 i_197647748(.A(n_57141), .B(n_258080081), .Z(n_57116));
	notech_or4 i_1921096(.A(n_288369895), .B(n_260280103), .C(n_261980120), 
		.D(n_26801), .Z(n_18937));
	notech_nand2 i_1721094(.A(n_263080131), .B(n_262680127), .Z(n_18925));
	notech_nand2 i_1921864(.A(n_264080141), .B(n_263680137), .Z(n_20726));
	notech_and2 i_106744547(.A(n_57329), .B(n_266680167), .Z(n_57982));
	notech_or2 i_85344546(.A(n_57730), .B(n_26662), .Z(n_58164));
	notech_mux2 i_3211701(.S(n_60550), .A(regs_14[31]), .B(add_len_pc32[31])
		, .Z(add_len_pc[31]));
	notech_and3 i_104563435(.A(n_318891635), .B(n_319091633), .C(n_26836), .Z
		(n_138061663));
	notech_nand2 i_3220725(.A(n_286080361), .B(n_285580356), .Z(n_24942));
	notech_nand2 i_620763(.A(n_287080371), .B(n_286580366), .Z(n_24460));
	notech_nand2 i_420761(.A(n_288080381), .B(n_287580376), .Z(n_24448));
	notech_nand2 i_620859(.A(n_289080391), .B(n_288580386), .Z(n_24112));
	notech_nand2 i_420857(.A(n_290080401), .B(n_289580396), .Z(n_24100));
	notech_or4 i_3221013(.A(n_215876097), .B(n_277980280), .C(n_290480405), 
		.D(n_26814), .Z(n_23920));
	notech_nand2 i_620987(.A(n_291780418), .B(n_291280413), .Z(n_23764));
	notech_nand2 i_420985(.A(n_292780428), .B(n_292280423), .Z(n_23752));
	notech_and4 i_3221109(.A(n_292880429), .B(n_293080431), .C(n_275680257),
		 .D(n_293580436), .Z(n_19015));
	notech_nand2 i_621083(.A(n_294680447), .B(n_294180442), .Z(n_18859));
	notech_nand2 i_421081(.A(n_295780458), .B(n_295280453), .Z(n_18847));
	notech_nand2 i_621179(.A(n_296680467), .B(n_296280463), .Z(n_18510));
	notech_nand2 i_421177(.A(n_297580476), .B(n_297180472), .Z(n_18498));
	notech_and4 i_3221557(.A(n_298380484), .B(n_298580486), .C(n_298280483),
		 .D(n_269780198), .Z(n_18318));
	notech_nand3 i_721628(.A(n_298880489), .B(n_298780488), .C(n_299280493),
		 .Z(n_17816));
	notech_nand2 i_621627(.A(n_300180502), .B(n_299780498), .Z(n_17810));
	notech_nand2 i_421625(.A(n_301080511), .B(n_300680507), .Z(n_17798));
	notech_ao4 i_5344441(.A(n_27989), .B(n_26810), .C(n_3868), .D(n_56675), 
		.Z(n_302621190));
	notech_and2 i_29610(.A(n_26964), .B(n_26999), .Z(n_137961662));
	notech_and2 i_34487(.A(n_25386), .B(n_125761540), .Z(n_137861661));
	notech_nand2 i_90663570(.A(n_2683), .B(n_27641), .Z(n_137661659));
	notech_and2 i_100841344(.A(n_58085), .B(n_304180542), .Z(n_58041));
	notech_nand2 i_99941343(.A(n_57877), .B(n_58190), .Z(n_58050));
	notech_ao4 i_99841342(.A(n_59441), .B(n_26824), .C(n_58171), .D(n_26800)
		, .Z(n_58051));
	notech_and2 i_64541341(.A(n_58427), .B(n_304080541), .Z(n_58372));
	notech_nand3 i_191241335(.A(n_57863), .B(n_301180512), .C(n_323280733), 
		.Z(n_57179));
	notech_ao4 i_191141334(.A(n_59441), .B(n_26827), .C(n_56471), .D(n_26826
		), .Z(n_57180));
	notech_and2 i_64241333(.A(n_58424), .B(n_303880539), .Z(n_58375));
	notech_mux2 i_111670(.S(n_60550), .A(n_5160), .B(add_len_pc32[0]), .Z(add_len_pc
		[0]));
	notech_mux2 i_911678(.S(n_60550), .A(n_5168), .B(add_len_pc32[8]), .Z(add_len_pc
		[8]));
	notech_mux2 i_1011679(.S(n_60550), .A(n_5169), .B(add_len_pc32[9]), .Z(add_len_pc
		[9]));
	notech_mux2 i_1111680(.S(n_60550), .A(n_5170), .B(add_len_pc32[10]), .Z(add_len_pc
		[10]));
	notech_mux2 i_1211681(.S(n_60550), .A(n_5171), .B(add_len_pc32[11]), .Z(add_len_pc
		[11]));
	notech_mux2 i_1411683(.S(n_60537), .A(n_5173), .B(add_len_pc32[13]), .Z(add_len_pc
		[13]));
	notech_mux2 i_1511684(.S(n_60537), .A(n_5174), .B(add_len_pc32[14]), .Z(add_len_pc
		[14]));
	notech_mux2 i_1611685(.S(n_60537), .A(n_5175), .B(add_len_pc32[15]), .Z(add_len_pc
		[15]));
	notech_or4 i_89563581(.A(n_27917), .B(n_61117), .C(n_60868), .D(n_27896)
		, .Z(n_136961652));
	notech_or4 i_39014(.A(n_58815), .B(n_17107), .C(n_26945), .D(n_26769), .Z
		(n_136861651));
	notech_nand2 i_1620709(.A(n_324880749), .B(n_324380744), .Z(n_24846));
	notech_nand2 i_1520708(.A(n_326580766), .B(n_325980760), .Z(n_24840));
	notech_nand2 i_1420707(.A(n_327780778), .B(n_327180772), .Z(n_24834));
	notech_nand2 i_1220705(.A(n_328980790), .B(n_328380784), .Z(n_24822));
	notech_nand2 i_1120704(.A(n_330080801), .B(n_329580796), .Z(n_24816));
	notech_nand2 i_1020703(.A(n_331180812), .B(n_330680807), .Z(n_24810));
	notech_nand2 i_920702(.A(n_332280823), .B(n_331780818), .Z(n_24804));
	notech_nand2 i_120694(.A(n_333480835), .B(n_332980830), .Z(n_24756));
	notech_and4 i_920766(.A(n_310880609), .B(n_333580836), .C(n_333780838), 
		.D(n_334680847), .Z(n_24478));
	notech_nand2 i_920862(.A(n_335580856), .B(n_335180852), .Z(n_24130));
	notech_and4 i_920990(.A(n_335680857), .B(n_335880859), .C(n_336380864), 
		.D(n_308980590), .Z(n_23782));
	notech_nand2 i_921086(.A(n_337280873), .B(n_336880869), .Z(n_18877));
	notech_and4 i_921182(.A(n_307080571), .B(n_337380874), .C(n_337580876), 
		.D(n_338080881), .Z(n_18528));
	notech_nand2 i_921854(.A(n_338980890), .B(n_338580886), .Z(n_20666));
	notech_nand2 i_917598(.A(n_339980900), .B(n_339480895), .Z(n_16754));
	notech_and3 i_60541276(.A(n_317991644), .B(n_318691637), .C(n_121628493)
		, .Z(n_291718116));
	notech_ao4 i_105541268(.A(n_59441), .B(n_27196), .C(n_2417), .D(n_26832)
		, .Z(n_290918108));
	notech_and2 i_105641267(.A(n_315991664), .B(n_302180522), .Z(n_290818107
		));
	notech_and3 i_105741266(.A(n_318191642), .B(n_316991654), .C(n_309091733
		), .Z(n_290718106));
	notech_or4 i_39011(.A(n_57020), .B(n_29658), .C(n_57064), .D(n_57033), .Z
		(n_136761650));
	notech_nand3 i_39009(.A(n_54929), .B(n_54794), .C(n_125661539), .Z(n_136661649
		));
	notech_nao3 i_30415(.A(n_32386), .B(n_32287), .C(n_56822), .Z(n_136561648
		));
	notech_or2 i_9364360(.A(n_285463121), .B(n_297363240), .Z(n_136461647)
		);
	notech_or2 i_9064363(.A(n_275363020), .B(n_26945), .Z(n_136361646));
	notech_or2 i_8764366(.A(n_275363020), .B(n_54794), .Z(n_136261645));
	notech_or2 i_30625(.A(n_285463121), .B(n_26945), .Z(n_136161644));
	notech_nao3 i_11064343(.A(n_126061543), .B(n_56414), .C(n_175162034), .Z
		(n_136061643));
	notech_or4 i_30635(.A(n_59387), .B(n_29178), .C(n_27192), .D(n_26810), .Z
		(n_135961642));
	notech_nao3 i_72363750(.A(opc[9]), .B(n_62814), .C(n_152461807), .Z(n_135861641
		));
	notech_xor2 i_133938298(.A(n_28051), .B(n_307215148), .Z(n_57710));
	notech_and4 i_50417(.A(n_344080941), .B(n_347480975), .C(n_348380984), .D
		(n_347180972), .Z(\nbus_11329[0] ));
	notech_or4 i_32532929(.A(tcmp), .B(n_26602), .C(n_61117), .D(instrc[122]
		), .Z(n_58692));
	notech_nand2 i_89532911(.A(n_58692), .B(n_341880919), .Z(n_58122));
	notech_mux2 i_3111700(.S(n_60537), .A(regs_14[30]), .B(add_len_pc32[30])
		, .Z(add_len_pc[30]));
	notech_nand2 i_19274(.A(n_29636), .B(n_29666), .Z(n_40675));
	notech_nand2 i_3120724(.A(n_349380994), .B(n_348880989), .Z(n_24936));
	notech_or2 i_72863745(.A(n_60016), .B(n_285563122), .Z(n_135161634));
	notech_or4 i_71163762(.A(n_62860), .B(n_136361646), .C(n_60935), .D(n_57957
		), .Z(n_134861631));
	notech_or4 i_71463759(.A(n_285463121), .B(n_60935), .C(n_28133), .D(n_54794
		), .Z(n_134561628));
	notech_or4 i_71763756(.A(n_62860), .B(n_285463121), .C(n_62814), .D(n_29614
		), .Z(n_134261625));
	notech_ao3 i_71863755(.A(n_318891635), .B(n_319091633), .C(n_57947), .Z(n_133961622
		));
	notech_or4 i_70163772(.A(n_62856), .B(n_136361646), .C(n_60935), .D(n_57574
		), .Z(n_133861621));
	notech_or2 i_70463769(.A(n_5743), .B(n_296863235), .Z(n_133561618));
	notech_or2 i_70763766(.A(n_275463021), .B(n_56064), .Z(n_133261615));
	notech_or4 i_70863765(.A(n_62860), .B(n_285463121), .C(n_62814), .D(n_29725
		), .Z(n_132961612));
	notech_or4 i_69163782(.A(n_62860), .B(n_136361646), .C(n_60935), .D(n_57542
		), .Z(n_132861611));
	notech_or2 i_69463779(.A(n_60024), .B(n_296863235), .Z(n_132561608));
	notech_or2 i_69763776(.A(n_275463021), .B(n_56010), .Z(n_132261605));
	notech_or4 i_69863775(.A(n_62840), .B(n_285463121), .C(n_62814), .D(n_56019
		), .Z(n_131961602));
	notech_nand3 i_68663786(.A(opc[0]), .B(n_62814), .C(n_26945), .Z(n_131661599
		));
	notech_nao3 i_67763795(.A(n_126361546), .B(n_56809), .C(n_126161544), .Z
		(n_131561598));
	notech_ao4 i_67663796(.A(n_305291771), .B(n_127561558), .C(n_26905), .D(n_126461547
		), .Z(n_131461597));
	notech_or4 i_67563797(.A(n_175062033), .B(n_126161544), .C(n_26789), .D(n_26945
		), .Z(n_131361596));
	notech_nao3 i_68263790(.A(n_318891635), .B(n_319091633), .C(n_57773), .Z
		(n_130861591));
	notech_nand2 i_106063421(.A(n_3825), .B(n_56625), .Z(n_130461587));
	notech_ao4 i_6364390(.A(n_56946), .B(n_3695), .C(n_30910), .D(n_32287), 
		.Z(n_130361586));
	notech_nand3 i_7164382(.A(n_27035), .B(n_30905), .C(n_130461587), .Z(n_130161584
		));
	notech_and2 i_104863432(.A(n_56625), .B(n_26836), .Z(n_129861581));
	notech_nand2 i_104663434(.A(n_56625), .B(n_341380914), .Z(n_129661579)
		);
	notech_or4 i_13264322(.A(n_138961672), .B(n_138861671), .C(n_142161704),
		 .D(n_26977), .Z(n_129561578));
	notech_nor2 i_13164323(.A(n_129861581), .B(n_26883), .Z(n_129461577));
	notech_and3 i_13064324(.A(n_184658942), .B(n_27034), .C(n_129661579), .Z
		(n_129361576));
	notech_ao4 i_10564348(.A(n_59440), .B(n_26833), .C(n_130161584), .D(n_26982
		), .Z(n_129261575));
	notech_or4 i_98563492(.A(n_32579), .B(n_26975), .C(n_143561718), .D(n_60303
		), .Z(n_129161574));
	notech_and3 i_10864345(.A(n_58020), .B(n_58009), .C(n_57976), .Z(n_128761570
		));
	notech_nand2 i_90163575(.A(n_26776), .B(n_57839), .Z(n_128361566));
	notech_and4 i_16664288(.A(n_146061743), .B(n_145761740), .C(n_2654), .D(n_145961742
		), .Z(n_128261565));
	notech_ao4 i_16564289(.A(n_26965), .B(n_60845), .C(n_23036), .D(n_128761570
		), .Z(n_128161564));
	notech_and2 i_16464290(.A(n_144861731), .B(n_128361566), .Z(n_128061563)
		);
	notech_ao4 i_4264411(.A(n_27907), .B(n_59435), .C(n_59419), .D(n_27904),
		 .Z(n_127961562));
	notech_ao3 i_86963607(.A(n_32386), .B(n_56625), .C(n_56829), .Z(n_127561558
		));
	notech_or4 i_86563611(.A(n_2938), .B(n_2937), .C(n_56829), .D(n_32287), 
		.Z(n_127161554));
	notech_nao3 i_86263614(.A(n_276163028), .B(n_32319), .C(n_175162034), .Z
		(n_127061553));
	notech_or2 i_86163615(.A(n_287163138), .B(n_54794), .Z(n_126961552));
	notech_and2 i_15764297(.A(n_58285), .B(n_147761760), .Z(n_126661549));
	notech_ao3 i_68363789(.A(n_56414), .B(\opa_12[0] ), .C(n_175162034), .Z(n_126461547
		));
	notech_nand3 i_15964295(.A(n_58646), .B(n_150661789), .C(n_131661599), .Z
		(n_126361546));
	notech_ao4 i_964441(.A(n_2480), .B(n_62892), .C(n_56829), .D(n_32287), .Z
		(n_126161544));
	notech_nand3 i_1864435(.A(n_54774), .B(n_146961752), .C(n_281263079), .Z
		(n_126061543));
	notech_or4 i_9764356(.A(n_2938), .B(n_2937), .C(n_56829), .D(n_32299), .Z
		(n_125961542));
	notech_or4 i_5264401(.A(calc_sz[3]), .B(n_2938), .C(n_25385), .D(calc_sz
		[2]), .Z(n_125761540));
	notech_or2 i_3964414(.A(n_58815), .B(n_26769), .Z(n_125661539));
	notech_or4 i_2564428(.A(instrc[122]), .B(n_175162034), .C(n_29179), .D(n_26735
		), .Z(n_125561538));
	notech_or4 i_112964452(.A(n_61138), .B(n_60263), .C(n_62814), .D(n_60910
		), .Z(n_125461537));
	notech_or4 i_35264454(.A(n_32563), .B(n_32548), .C(n_144761730), .D(n_32580
		), .Z(n_125361536));
	notech_and4 i_118266246(.A(n_124761530), .B(n_123061513), .C(n_123161514
		), .D(n_123261515), .Z(n_125061533));
	notech_and4 i_117966249(.A(n_124561528), .B(n_124461527), .C(n_124261525
		), .D(n_124161524), .Z(n_124761530));
	notech_ao4 i_117666252(.A(n_1895), .B(n_60263), .C(n_58768), .D(n_29740)
		, .Z(n_124561528));
	notech_ao4 i_117566253(.A(n_53341148), .B(nbus_11295[3]), .C(n_53641151)
		, .D(n_57563), .Z(n_124461527));
	notech_ao4 i_117466254(.A(n_53841153), .B(n_29739), .C(n_54141156), .D(n_29738
		), .Z(n_124261525));
	notech_ao4 i_117366255(.A(n_40241017), .B(n_29089), .C(n_39041005), .D(n_28929
		), .Z(n_124161524));
	notech_or4 i_109766331(.A(n_61175), .B(n_61165), .C(n_3792), .D(n_19101)
		, .Z(n_124061523));
	notech_or4 i_33367402(.A(n_55524), .B(n_26964), .C(n_19079), .D(n_19101)
		, .Z(n_24540860));
	notech_or4 i_5367348(.A(n_55508), .B(n_59241), .C(n_59187), .D(n_59259),
		 .Z(n_25140866));
	notech_mux2 i_110466324(.S(opd[2]), .A(n_55508), .B(n_27040885), .Z(n_123661519
		));
	notech_mux2 i_2167379(.S(opd[0]), .A(n_55508), .B(n_27040885), .Z(n_123561518
		));
	notech_nand3 i_31867403(.A(n_19109), .B(n_60263), .C(n_19101), .Z(n_27040885
		));
	notech_nao3 i_3167369(.A(n_56662), .B(n_190262174), .C(n_329763514), .Z(n_83341448
		));
	notech_and4 i_412921(.A(n_123361516), .B(n_125061533), .C(n_330063517), 
		.D(n_122161504), .Z(n_25963));
	notech_or2 i_116966259(.A(n_24540860), .B(n_28092), .Z(n_123361516));
	notech_nand2 i_117066258(.A(add_src[3]), .B(n_26723), .Z(n_123261515));
	notech_or2 i_116866260(.A(n_329363510), .B(n_29741), .Z(n_123161514));
	notech_or2 i_117266256(.A(n_25140866), .B(opd[3]), .Z(n_123061513));
	notech_nand2 i_117166257(.A(opd[3]), .B(n_329563512), .Z(n_122161504));
	notech_and3 i_109166337(.A(n_19109), .B(n_330363520), .C(n_60373), .Z(n_121261495
		));
	notech_nao3 i_39967028(.A(n_60095), .B(n_318891635), .C(n_246791942), .Z
		(n_121161494));
	notech_nand2 i_40067027(.A(n_329263509), .B(imm[3]), .Z(n_121061493));
	notech_ao4 i_127168591(.A(n_136861651), .B(n_28126), .C(n_136761650), .D
		(n_27730), .Z(n_120861491));
	notech_ao4 i_127268590(.A(n_136661649), .B(n_27768), .C(n_54929), .D(n_27426
		), .Z(n_120761490));
	notech_nand2 i_27416(.A(n_26964), .B(n_60263), .Z(n_32559));
	notech_or2 i_50488(.A(n_27037), .B(n_26757), .Z(n_19072));
	notech_or4 i_50481(.A(fsm[0]), .B(fsm[3]), .C(n_26757), .D(n_27717), .Z(n_19109
		));
	notech_and4 i_50478(.A(fsm[0]), .B(n_2885), .C(fsm[1]), .D(n_27720), .Z(n_19127
		));
	notech_and4 i_9582203(.A(n_57552), .B(n_3787), .C(n_57563), .D(n_57574),
		 .Z(n_27885));
	notech_or2 i_50503(.A(n_2896), .B(n_3790), .Z(n_18998));
	notech_nor2 i_50505(.A(n_3790), .B(n_3792), .Z(n_18989));
	notech_or4 i_155182202(.A(n_32566), .B(n_19022), .C(n_19014), .D(n_19036
		), .Z(n_32563));
	notech_and3 i_134082201(.A(fsm[0]), .B(n_27717), .C(fsm[3]), .Z(n_32562)
		);
	notech_and3 i_50496(.A(n_61165), .B(n_61175), .C(n_3794), .Z(n_19036));
	notech_or4 i_117882200(.A(n_32569), .B(n_3804), .C(n_19050), .D(n_19036)
		, .Z(n_32565));
	notech_nao3 i_22782199(.A(n_32586), .B(n_60127), .C(n_32581), .Z(n_32579
		));
	notech_nand3 i_22582198(.A(n_19093), .B(n_60372), .C(n_32586), .Z(n_32580
		));
	notech_and4 i_22382197(.A(n_19109), .B(n_19117), .C(n_26761), .D(n_19137
		), .Z(n_32586));
	notech_nand2 i_50476(.A(n_2885), .B(n_3794), .Z(n_19137));
	notech_or4 i_50479(.A(fsm[3]), .B(fsm[0]), .C(fsm[1]), .D(n_26757), .Z(n_19117
		));
	notech_and4 i_50482(.A(fsm[0]), .B(n_27720), .C(fsm[1]), .D(n_32605), .Z
		(n_19101));
	notech_nand2 i_50484(.A(n_2885), .B(n_3796), .Z(n_19093));
	notech_ao3 i_50491(.A(n_61165), .B(n_272491901), .C(n_61175), .Z(n_19057
		));
	notech_ao3 i_50493(.A(n_61165), .B(n_3794), .C(n_61175), .Z(n_19050));
	notech_and4 i_50499(.A(fsm[0]), .B(n_27720), .C(fsm[1]), .D(n_2880), .Z(n_19022
		));
	notech_ao3 i_50502(.A(n_61167), .B(n_32562), .C(fsm[2]), .Z(n_19006));
	notech_ao3 i_50506(.A(n_61167), .B(fsm[2]), .C(n_27037), .Z(n_18981));
	notech_and4 i_50509(.A(fsm[3]), .B(fsm[0]), .C(fsm[1]), .D(n_32605), .Z(n_18964
		));
	notech_and3 i_50508(.A(n_61167), .B(fsm[2]), .C(n_32562), .Z(n_18972));
	notech_nor2 i_27424(.A(n_3806), .B(n_32579), .Z(n_32551));
	notech_or4 i_27422(.A(n_32555), .B(n_19057), .C(n_60303), .D(n_19006), .Z
		(n_32553));
	notech_or4 i_27409(.A(n_3804), .B(n_19086), .C(n_19079), .D(n_19050), .Z
		(n_32566));
	notech_nao3 i_27408(.A(n_26983), .B(n_26985), .C(n_3804), .Z(n_32567));
	notech_nand2 i_27406(.A(n_26983), .B(n_26985), .Z(n_32569));
	notech_nand2 i_27394(.A(n_19093), .B(n_60372), .Z(n_32581));
	notech_or2 i_28832495(.A(n_30312), .B(n_56463), .Z(n_3925));
	notech_or4 i_26232515(.A(n_32555), .B(n_32559), .C(n_32579), .D(n_3698),
		 .Z(n_5968810));
	notech_nand2 i_163382191(.A(n_18998), .B(n_26989), .Z(n_32596));
	notech_or2 i_20432566(.A(n_3730), .B(n_32334), .Z(n_30315));
	notech_and4 i_15832584(.A(n_3668), .B(n_3767), .C(n_3667), .D(n_27039), 
		.Z(n_3923));
	notech_ao3 i_50722(.A(instrc[126]), .B(n_30930), .C(instrc[125]), .Z(n_3922
		));
	notech_or4 i_50725(.A(instrc[101]), .B(n_29665), .C(instrc[100]), .D(instrc
		[103]), .Z(n_3921));
	notech_or4 i_50727(.A(instrc[97]), .B(n_29667), .C(instrc[99]), .D(instrc
		[96]), .Z(n_3920));
	notech_and4 i_50728(.A(n_29636), .B(instrc[94]), .C(n_29634), .D(n_29638
		), .Z(n_3919));
	notech_or4 i_50730(.A(instrc[89]), .B(n_29668), .C(instrc[91]), .D(instrc
		[88]), .Z(n_3918));
	notech_and4 i_111532761(.A(n_3925), .B(n_3910), .C(n_3760), .D(n_3639), 
		.Z(n_3917));
	notech_nand2 i_32402(.A(n_3590), .B(n_27714), .Z(n_3916));
	notech_and2 i_193932764(.A(instrc[125]), .B(instrc[126]), .Z(n_28120));
	notech_nand2 i_164932767(.A(instrc[104]), .B(instrc[107]), .Z(n_30303)
		);
	notech_and2 i_194432768(.A(instrc[127]), .B(instrc[124]), .Z(n_30322));
	notech_and2 i_25649(.A(n_3826), .B(n_30910), .Z(n_3915));
	notech_and2 i_164732773(.A(instrc[105]), .B(n_57369), .Z(n_30933));
	notech_or4 i_830224(.A(instrc[105]), .B(n_29736), .C(instrc[107]), .D(instrc
		[104]), .Z(n_3914));
	notech_and2 i_120132774(.A(n_29737), .B(n_57369), .Z(n_30939));
	notech_and2 i_175132698(.A(instrc[101]), .B(instrc[103]), .Z(n_30952));
	notech_and2 i_184432777(.A(instrc[93]), .B(instrc[94]), .Z(n_30966));
	notech_and2 i_185232697(.A(instrc[89]), .B(instrc[91]), .Z(n_30973));
	notech_nand2 i_26921(.A(n_27853), .B(all_cnt[0]), .Z(n_3913));
	notech_and2 i_25215(.A(all_cnt[1]), .B(all_cnt[0]), .Z(n_32420));
	notech_and3 i_197532816(.A(all_cnt[1]), .B(all_cnt[2]), .C(all_cnt[0]), 
		.Z(n_32421));
	notech_or4 i_22132549(.A(n_2893), .B(n_60935), .C(n_60910), .D(reps[2]),
		 .Z(n_32452));
	notech_or4 i_22232548(.A(fsm[2]), .B(n_61167), .C(n_2896), .D(n_32476), 
		.Z(n_3912));
	notech_or4 i_13032611(.A(n_32581), .B(n_26900), .C(n_61131), .D(n_60303)
		, .Z(n_32476));
	notech_or2 i_12332618(.A(n_18981), .B(n_18972), .Z(n_32548));
	notech_and2 i_21532555(.A(n_27580), .B(n_27377), .Z(n_3911));
	notech_or2 i_11716(.A(n_3911), .B(n_26702), .Z(n_3910));
	notech_or4 i_29682(.A(n_59322), .B(n_30294), .C(n_26900), .D(n_30359), .Z
		(n_3908));
	notech_and4 i_50487(.A(fsm[3]), .B(fsm[0]), .C(n_2885), .D(fsm[1]), .Z(n_19079
		));
	notech_and3 i_56140(.A(n_27570), .B(n_26992), .C(n_3636), .Z(n_3907));
	notech_and4 i_55746(.A(n_318091643), .B(n_3739), .C(n_3737), .D(n_3696),
		 .Z(n_3906));
	notech_nao3 i_182332910(.A(n_2885), .B(n_3794), .C(n_59322), .Z(n_107111189
		));
	notech_or4 i_9539(.A(n_61154), .B(n_320063467), .C(n_26757), .D(n_19127)
		, .Z(n_3905));
	notech_xor2 i_2535075(.A(n_341791456), .B(n_341591458), .Z(n_3904));
	notech_or4 i_119035091(.A(fsm[2]), .B(n_61167), .C(n_61154), .D(n_1871),
		 .Z(n_3903));
	notech_or4 i_118935092(.A(fsm[2]), .B(n_61167), .C(n_61154), .D(n_1870),
		 .Z(n_3902));
	notech_or4 i_42435097(.A(n_59419), .B(n_25629), .C(n_60263), .D(n_57957)
		, .Z(n_3901));
	notech_and4 i_317752(.A(n_3586), .B(n_3579), .C(n_357091303), .D(n_356491309
		), .Z(n_3900));
	notech_and4 i_417753(.A(n_355491319), .B(n_354891325), .C(n_354191332), 
		.D(n_353591338), .Z(n_3899));
	notech_and4 i_517754(.A(n_352591348), .B(n_351991354), .C(n_351291361), 
		.D(n_350691367), .Z(n_3898));
	notech_and4 i_717756(.A(n_349691377), .B(n_349091383), .C(n_348391390), 
		.D(n_347791396), .Z(n_3897));
	notech_and4 i_817757(.A(n_346791406), .B(n_346191412), .C(n_345391420), 
		.D(n_344791426), .Z(n_3896));
	notech_or4 i_321368(.A(n_338091493), .B(n_342391450), .C(n_343591438), .D
		(n_27057), .Z(n_3895));
	notech_or4 i_28135114(.A(n_25615), .B(n_62848), .C(n_62814), .D(n_60263)
		, .Z(n_25329));
	notech_or4 i_169135119(.A(fsm[2]), .B(n_61167), .C(n_61154), .D(n_32446)
		, .Z(n_3894));
	notech_nao3 i_163532901(.A(n_2885), .B(n_2896), .C(n_3792), .Z(n_25397)
		);
	notech_and2 i_157735133(.A(n_32263), .B(n_308012096), .Z(n_3893));
	notech_or4 i_151635116(.A(n_25629), .B(n_62848), .C(n_62814), .D(n_60263
		), .Z(n_3892));
	notech_or4 i_40435115(.A(fsm[2]), .B(n_61167), .C(n_61154), .D(n_58046),
		 .Z(n_3889));
	notech_ao4 i_2338211(.A(n_58046), .B(n_60263), .C(n_58220), .D(n_330763524
		), .Z(n_34012440));
	notech_ao4 i_159438220(.A(n_19117), .B(n_25641), .C(mask8b[2]), .D(n_25640
		), .Z(n_3888));
	notech_ao4 i_81038225(.A(n_54912649), .B(n_59344), .C(n_58746), .D(n_308860169
		), .Z(n_3887));
	notech_and2 i_45138228(.A(n_296060041), .B(n_3888), .Z(n_3886));
	notech_or4 i_180938235(.A(n_60893), .B(n_25625), .C(n_28081), .D(n_60263
		), .Z(n_54512645));
	notech_and4 i_38738239(.A(n_3892), .B(n_337091503), .C(n_34012440), .D(n_309660177
		), .Z(n_388560287));
	notech_and2 i_38138240(.A(n_296860049), .B(n_25613), .Z(n_388360286));
	notech_ao4 i_35738248(.A(n_2895), .B(n_60263), .C(n_308760168), .D(n_309060171
		), .Z(n_3882));
	notech_nand3 i_316216(.A(n_311060191), .B(n_310560186), .C(n_312160202),
		 .Z(n_3881));
	notech_and2 i_141738257(.A(n_25629), .B(n_58220), .Z(n_3880));
	notech_nand3 i_84341361(.A(n_211359194), .B(n_56843), .C(n_3853), .Z(n_3879
		));
	notech_or2 i_118341390(.A(n_183858934), .B(n_3845), .Z(n_3878));
	notech_nao3 i_117541392(.A(n_32335), .B(n_26670), .C(n_54954), .Z(n_3877
		));
	notech_nao3 i_82141397(.A(n_3879), .B(n_32335), .C(n_54954), .Z(n_3876)
		);
	notech_and4 i_91738294(.A(n_306960150), .B(n_306860149), .C(n_306460145)
		, .D(n_306760148), .Z(n_3874));
	notech_ao4 i_6444430(.A(n_3874), .B(n_58432), .C(n_58530), .D(n_56082), 
		.Z(n_3873));
	notech_nand3 i_44944492(.A(n_60910), .B(n_62814), .C(\opa_12[6] ), .Z(n_92519107
		));
	notech_or4 i_44544494(.A(n_60964), .B(n_60953), .C(n_62848), .D(n_29723)
		, .Z(n_92619108));
	notech_and4 i_417017(.A(n_292160002), .B(n_292060001), .C(n_291960000), 
		.D(n_292560006), .Z(n_3872));
	notech_and4 i_617019(.A(n_290759988), .B(n_290659987), .C(n_290559986), 
		.D(n_291159992), .Z(n_3871));
	notech_nand2 i_717020(.A(n_289859979), .B(n_289259973), .Z(n_3870));
	notech_or4 i_721372(.A(n_283259913), .B(n_287559956), .C(n_288559966), .D
		(n_27072), .Z(n_3869));
	notech_and4 i_142944499(.A(n_286959950), .B(n_286859949), .C(n_286459945
		), .D(n_286759948), .Z(n_3868));
	notech_or4 i_130244507(.A(n_27925), .B(n_32643), .C(n_59419), .D(n_60263
		), .Z(n_3867));
	notech_or2 i_19597(.A(n_277459855), .B(n_276159842), .Z(n_3866));
	notech_or2 i_153844573(.A(n_3867), .B(n_27025), .Z(n_125828535));
	notech_ao4 i_121544578(.A(n_32382), .B(n_27076), .C(n_56979), .D(n_3633)
		, .Z(n_3865));
	notech_and4 i_92938282(.A(n_305560136), .B(n_305460135), .C(n_305060131)
		, .D(n_305360134), .Z(n_3864));
	notech_and4 i_1717030(.A(n_275659837), .B(n_275559836), .C(n_275459835),
		 .D(n_275959840), .Z(n_3863));
	notech_nand2 i_1917032(.A(n_274659827), .B(n_274159822), .Z(n_3862));
	notech_and4 i_144147709(.A(n_273359814), .B(n_273259813), .C(n_272859809
		), .D(n_273159812), .Z(n_3861));
	notech_and4 i_317016(.A(n_266759748), .B(n_266659747), .C(n_266559746), 
		.D(n_267159752), .Z(n_3860));
	notech_nand2 i_2317036(.A(n_265659737), .B(n_265159732), .Z(n_3859));
	notech_ao4 i_86744551(.A(n_59440), .B(n_27029), .C(n_3879), .D(n_26669),
		 .Z(n_148128758));
	notech_and2 i_86844552(.A(n_3876), .B(n_25875), .Z(n_148228759));
	notech_or4 i_96658533(.A(n_55581), .B(n_57051), .C(n_29658), .D(n_3845),
		 .Z(n_3858));
	notech_or4 i_58758553(.A(n_59355), .B(n_56829), .C(n_27192), .D(n_56946)
		, .Z(n_3857));
	notech_nand2 i_202153909(.A(read_data[26]), .B(n_60263), .Z(n_3884));
	notech_or4 i_3399(.A(n_32643), .B(n_27123), .C(n_60868), .D(n_27125), .Z
		(n_3986));
	notech_nand2 i_3117044(.A(n_213859219), .B(n_213359214), .Z(n_3856));
	notech_ao4 i_51055530(.A(n_32352), .B(n_32284), .C(n_56854), .D(n_26962)
		, .Z(n_26055));
	notech_ao3 i_19355532(.A(n_57064), .B(n_57078), .C(n_55581), .Z(n_26061)
		);
	notech_ao4 i_53455625(.A(n_56813), .B(n_32284), .C(n_56854), .D(n_32382)
		, .Z(n_26054));
	notech_ao4 i_83455574(.A(n_62826), .B(n_60910), .C(n_60893), .D(n_26061)
		, .Z(n_3854));
	notech_ao4 i_52655629(.A(n_56675), .B(n_32284), .C(n_56854), .D(n_56979)
		, .Z(n_3853));
	notech_and2 i_23555640(.A(n_30821), .B(n_30470), .Z(n_3852));
	notech_and4 i_143341319(.A(n_295460035), .B(n_295360034), .C(n_294960030
		), .D(n_295260033), .Z(n_3851));
	notech_and4 i_92138290(.A(n_308360164), .B(n_308260163), .C(n_307860159)
		, .D(n_308160162), .Z(n_3850));
	notech_or2 i_8458407(.A(n_3867), .B(n_3596), .Z(n_3849));
	notech_nand2 i_1117024(.A(n_211159192), .B(n_210559186), .Z(n_3848));
	notech_and4 i_521914(.A(n_209559176), .B(n_209459175), .C(n_209359174), 
		.D(n_209859179), .Z(n_3847));
	notech_ao4 i_260558502(.A(calc_sz[1]), .B(n_56970), .C(n_32386), .D(n_26627
		), .Z(n_3846));
	notech_ao4 i_51855632(.A(n_56688), .B(n_32284), .C(n_56854), .D(n_56946)
		, .Z(n_3845));
	notech_or2 i_162755529(.A(n_54954), .B(n_32335), .Z(n_3844));
	notech_or4 i_108061761(.A(n_55581), .B(n_57051), .C(n_29658), .D(n_192159008
		), .Z(n_3843));
	notech_nand2 i_217015(.A(n_206159142), .B(n_205459135), .Z(n_3842));
	notech_nand2 i_1317026(.A(n_204759128), .B(n_204159122), .Z(n_3841));
	notech_and4 i_1417027(.A(n_203059111), .B(n_202959110), .C(n_202859109),
		 .D(n_203459115), .Z(n_3840));
	notech_and4 i_1517028(.A(n_201659097), .B(n_201559096), .C(n_201459095),
		 .D(n_202059101), .Z(n_3839));
	notech_nand2 i_2217035(.A(n_200759088), .B(n_200259083), .Z(n_3838));
	notech_nao3 i_33932(.A(n_57988), .B(n_319091633), .C(n_59355), .Z(n_3837
		));
	notech_ao4 i_193361789(.A(n_306791756), .B(n_305891765), .C(n_30821), .D
		(n_61115), .Z(n_3836));
	notech_or4 i_35632898(.A(n_27925), .B(n_59419), .C(n_32643), .D(n_3595),
		 .Z(n_3835));
	notech_ao4 i_60058552(.A(n_54954), .B(n_32335), .C(n_59419), .D(n_26061)
		, .Z(n_3834));
	notech_nand2 i_30030(.A(n_26991), .B(n_62784), .Z(n_3833));
	notech_ao4 i_94832913(.A(n_26894), .B(n_27045), .C(n_30312), .D(n_3753),
		 .Z(n_3832));
	notech_nand2 i_2578(.A(n_3908), .B(n_26838), .Z(n_3830));
	notech_and2 i_8264371(.A(n_29734), .B(instrc[104]), .Z(n_28132));
	notech_and2 i_7764376(.A(n_29639), .B(instrc[96]), .Z(n_28130));
	notech_and3 i_1364437(.A(n_3826), .B(n_30910), .C(n_3827), .Z(n_3829));
	notech_and2 i_1264438(.A(n_29663), .B(instrc[124]), .Z(n_28122));
	notech_or2 i_31532827(.A(n_56944), .B(n_3695), .Z(n_3828));
	notech_and3 i_664443(.A(n_3828), .B(n_27035), .C(n_30905), .Z(n_74438764
		));
	notech_or4 i_25650(.A(n_32378), .B(n_7298943), .C(n_32730), .D(n_306391760
		), .Z(n_3827));
	notech_or4 i_27432771(.A(n_32378), .B(n_7298943), .C(n_32730), .D(n_56959
		), .Z(n_3826));
	notech_nand2 i_464444(.A(n_3826), .B(n_3827), .Z(n_3825));
	notech_ao3 i_264445(.A(n_27034), .B(n_3833), .C(n_183058926), .Z(n_3824)
		);
	notech_nor2 i_113632902(.A(n_3594), .B(n_60935), .Z(n_3823));
	notech_and2 i_164446(.A(n_184658942), .B(n_27034), .Z(n_251040528));
	notech_nor2 i_31432826(.A(n_3695), .B(n_56959), .Z(n_3822));
	notech_nand2 i_161064464(.A(fecx), .B(n_61131), .Z(n_3821));
	notech_or4 i_12026(.A(n_61117), .B(n_27917), .C(n_62848), .D(n_62824), .Z
		(n_3820));
	notech_nor2 i_28732820(.A(n_6258839), .B(n_27052), .Z(n_3819));
	notech_and3 i_47552(.A(n_184758943), .B(n_184858944), .C(n_26992), .Z(n_3818
		));
	notech_and4 i_52154(.A(n_340991464), .B(n_340891465), .C(n_340791466), .D
		(n_191859005), .Z(n_3817));
	notech_and4 i_53131(.A(n_191058997), .B(n_191759004), .C(n_185858954), .D
		(n_190958996), .Z(n_3816));
	notech_and4 i_51465(.A(n_189858988), .B(n_3821), .C(n_189758987), .D(n_189358984
		), .Z(n_3815));
	notech_or2 i_121658506(.A(n_26611), .B(n_3846), .Z(n_3814));
	notech_nor2 i_50500(.A(n_27037), .B(n_3790), .Z(n_19014));
	notech_nor2 i_30432479(.A(n_3593), .B(n_7298943), .Z(n_3813));
	notech_or2 i_14932592(.A(n_26602), .B(tcmp), .Z(n_30312));
	notech_or4 i_30696(.A(n_32596), .B(n_19014), .C(n_29282), .D(n_19006), .Z
		(n_3812));
	notech_and4 i_20532565(.A(all_cnt[0]), .B(n_3914), .C(all_cnt[1]), .D(n_320191622
		), .Z(n_30301));
	notech_or4 i_43432712(.A(all_cnt[2]), .B(all_cnt[1]), .C(n_27042), .D(n_3922
		), .Z(n_30294));
	notech_nor2 i_194232772(.A(instrc[125]), .B(n_29664), .Z(n_30931));
	notech_ao3 i_44132707(.A(n_32421), .B(n_3918), .C(all_cnt[3]), .Z(n_3811
		));
	notech_ao3 i_44032708(.A(n_27090), .B(n_6858899), .C(n_27042), .Z(n_30366
		));
	notech_and4 i_43832710(.A(all_cnt[2]), .B(n_3921), .C(n_27853), .D(n_3724
		), .Z(n_3810));
	notech_and2 i_195032778(.A(n_29631), .B(instrc[90]), .Z(n_30976));
	notech_nand2 i_22153(.A(n_29636), .B(instrc[94]), .Z(n_30969));
	notech_and2 i_194832775(.A(n_29635), .B(instrc[102]), .Z(n_30955));
	notech_and2 i_1467386(.A(n_32434), .B(n_32432), .Z(n_268643294));
	notech_or4 i_30697(.A(n_32567), .B(n_19050), .C(n_19036), .D(n_19043), .Z
		(n_3807));
	notech_or4 i_10082141(.A(n_32555), .B(n_32559), .C(n_32563), .D(n_19006)
		, .Z(n_3806));
	notech_nand2 i_51982140(.A(n_19072), .B(n_19065), .Z(n_3804));
	notech_nao3 i_22482139(.A(n_19029), .B(n_26963), .C(n_32559), .Z(n_3803)
		);
	notech_ao3 i_162282132(.A(n_27717), .B(fsm[3]), .C(fsm[0]), .Z(n_3796)
		);
	notech_and3 i_183082130(.A(fsm[0]), .B(n_27717), .C(n_27720), .Z(n_3794)
		);
	notech_nand3 i_179982128(.A(fsm[0]), .B(fsm[3]), .C(fsm[1]), .Z(n_3792)
		);
	notech_nand2 i_137082126(.A(n_61167), .B(n_27719), .Z(n_3790));
	notech_or4 i_100782125(.A(opa[0]), .B(opa[1]), .C(opa[2]), .D(opa[3]), .Z
		(n_3789));
	notech_nand3 i_96082124(.A(\nbus_11307[0] ), .B(n_57542), .C(n_57552), .Z
		(n_3788));
	notech_and2 i_78082123(.A(\nbus_11307[0] ), .B(n_57542), .Z(n_3787));
	notech_nao3 i_111031762(.A(n_32605), .B(n_26761), .C(n_61154), .Z(n_3786
		));
	notech_or4 i_122231660(.A(\nbus_11307[0] ), .B(opa[1]), .C(opa[3]), .D(opa
		[4]), .Z(n_3784));
	notech_or4 i_122731655(.A(n_3633), .B(opa[6]), .C(opa[7]), .D(n_27046), 
		.Z(n_3781));
	notech_or4 i_23732536(.A(n_32580), .B(n_32555), .C(n_32559), .D(n_61131)
		, .Z(n_3777));
	notech_or4 i_22974(.A(n_3641), .B(n_3640), .C(n_3646), .D(n_3645), .Z(n_3776
		));
	notech_ao4 i_127931605(.A(n_26601), .B(n_30344), .C(n_29256), .D(n_3766)
		, .Z(n_3767));
	notech_nand2 i_128131603(.A(instrc[100]), .B(instrc[102]), .Z(n_3766));
	notech_ao4 i_126331621(.A(n_3916), .B(n_32378), .C(n_3911), .D(n_26643),
		 .Z(n_3760));
	notech_or4 i_126731617(.A(n_29663), .B(n_29632), .C(n_26891), .D(n_32747
		), .Z(n_3759));
	notech_ao4 i_28232499(.A(n_304591778), .B(n_56941), .C(n_59435), .D(n_32380
		), .Z(n_3758));
	notech_or4 i_25932518(.A(n_3806), .B(n_32579), .C(n_32596), .D(n_32548),
		 .Z(n_6258839));
	notech_nand3 i_130631579(.A(instrc[122]), .B(n_60127), .C(n_60303), .Z(n_3753
		));
	notech_nand2 i_20632564(.A(n_3811), .B(n_26841), .Z(n_6368850));
	notech_and4 i_44167(.A(all_cnt[0]), .B(n_27853), .C(all_cnt[2]), .D(n_27856
		), .Z(n_3751));
	notech_or4 i_22732543(.A(n_59322), .B(n_26900), .C(n_30359), .D(n_26724)
		, .Z(n_6588872));
	notech_or4 i_133731548(.A(n_19022), .B(n_32555), .C(n_19057), .D(n_19050
		), .Z(n_3742));
	notech_ao4 i_134131544(.A(n_60122), .B(n_27246), .C(n_3829), .D(n_56592)
		, .Z(n_3739));
	notech_ao4 i_134331542(.A(n_3701), .B(n_3624), .C(n_61115), .D(n_3623), 
		.Z(n_3737));
	notech_ao4 i_134831537(.A(n_30315), .B(n_56396), .C(n_3729), .D(n_3690),
		 .Z(n_3731));
	notech_nand3 i_5317(.A(all_cnt[0]), .B(n_27853), .C(n_320191622), .Z(n_3730
		));
	notech_or4 i_7232667(.A(all_cnt[0]), .B(all_cnt[1]), .C(n_27070), .D(n_3922
		), .Z(n_3729));
	notech_and2 i_201232688(.A(n_27852), .B(n_27856), .Z(n_3724));
	notech_and4 i_5336(.A(all_cnt[0]), .B(all_cnt[1]), .C(all_cnt[2]), .D(n_27856
		), .Z(n_6888902));
	notech_ao3 i_135131534(.A(n_3686), .B(n_3685), .C(n_3683), .Z(n_3720));
	notech_or4 i_7132668(.A(all_cnt[0]), .B(n_27070), .C(n_27853), .D(n_17107
		), .Z(n_3714));
	notech_and3 i_6632673(.A(instrc[98]), .B(instrc[99]), .C(instrc[97]), .Z
		(n_3706));
	notech_or4 i_20332567(.A(n_32555), .B(n_3698), .C(n_314463411), .D(n_314663413
		), .Z(n_3701));
	notech_or4 i_11732624(.A(n_27037), .B(n_3790), .C(n_19022), .D(n_32565),
		 .Z(n_3698));
	notech_ao4 i_134431541(.A(n_3622), .B(n_3621), .C(n_314663413), .D(n_3688
		), .Z(n_3696));
	notech_or4 i_26032517(.A(tcmp), .B(n_61115), .C(n_32378), .D(\opcode[3] 
		), .Z(n_3695));
	notech_nand3 i_200532689(.A(n_60122), .B(n_60303), .C(n_27714), .Z(n_7298943
		));
	notech_nao3 i_138431505(.A(instrc[125]), .B(n_29632), .C(n_340480905), .Z
		(n_3690));
	notech_nao3 i_138831501(.A(n_60372), .B(n_19093), .C(n_266891921), .Z(n_3688
		));
	notech_or4 i_31032473(.A(n_32378), .B(n_7298943), .C(n_32730), .D(n_56941
		), .Z(n_30910));
	notech_or4 i_74732098(.A(all_cnt[3]), .B(all_cnt[1]), .C(n_3625), .D(n_27854
		), .Z(n_3686));
	notech_nand3 i_74532099(.A(n_30933), .B(n_26844), .C(n_30301), .Z(n_3685
		));
	notech_and4 i_74332100(.A(n_57020), .B(n_57078), .C(n_27043), .D(n_159379097
		), .Z(n_3683));
	notech_and2 i_29021(.A(n_29633), .B(n_29637), .Z(n_30954));
	notech_or4 i_29614(.A(n_27037), .B(n_3790), .C(n_3742), .D(n_19036), .Z(n_30361
		));
	notech_and3 i_31132472(.A(n_3810), .B(n_30352), .C(instrc[100]), .Z(n_30350
		));
	notech_ao3 i_29633(.A(n_57020), .B(n_30352), .C(n_30344), .Z(n_30342));
	notech_ao3 i_29618(.A(n_30366), .B(instrc[92]), .C(n_30359), .Z(n_30357)
		);
	notech_and3 i_31832469(.A(n_26841), .B(n_26760), .C(n_30301), .Z(n_30300
		));
	notech_and2 i_29000(.A(n_29640), .B(n_29642), .Z(n_3673));
	notech_nao3 i_30732476(.A(n_26841), .B(instrc[90]), .C(n_26727), .Z(n_30306
		));
	notech_ao3 i_30932474(.A(instrc[122]), .B(n_56391), .C(n_3730), .Z(n_3672
		));
	notech_and4 i_29643(.A(n_60122), .B(n_60263), .C(n_32586), .D(instrc[98]
		), .Z(n_30332));
	notech_nand3 i_30719(.A(instrc[101]), .B(instrc[103]), .C(n_3810), .Z(n_29256
		));
	notech_or4 i_70232137(.A(n_26891), .B(n_30294), .C(n_29663), .D(n_29632)
		, .Z(n_3668));
	notech_nao3 i_70132138(.A(n_30933), .B(n_30301), .C(n_30303), .Z(n_3667)
		);
	notech_and4 i_69832141(.A(n_30366), .B(instrc[92]), .C(instrc[95]), .D(n_30966
		), .Z(n_3646));
	notech_and4 i_69732142(.A(instrc[123]), .B(instrc[120]), .C(instrc[121])
		, .D(n_3672), .Z(n_3645));
	notech_and4 i_70032139(.A(n_30973), .B(n_3811), .C(instrc[88]), .D(instrc
		[90]), .Z(n_3641));
	notech_and4 i_69932140(.A(n_56888), .B(n_3751), .C(instrc[96]), .D(n_3706
		), .Z(n_3640));
	notech_or2 i_70932130(.A(n_26602), .B(n_27377), .Z(n_3639));
	notech_ao4 i_32405(.A(n_3598), .B(n_61131), .C(n_27377), .D(n_3912), .Z(n_27570
		));
	notech_or2 i_69632143(.A(n_3923), .B(n_5968810), .Z(n_3636));
	notech_nao3 i_30632477(.A(n_30366), .B(n_29634), .C(n_30359), .Z(n_29954
		));
	notech_or4 i_33016(.A(n_59322), .B(n_29954), .C(n_26900), .D(instrc[95])
		, .Z(n_26959));
	notech_nao3 i_33019(.A(n_29632), .B(n_3830), .C(instrc[127]), .Z(n_26956
		));
	notech_or4 i_79053915(.A(opa[8]), .B(opa[9]), .C(n_241659497), .D(n_241559496
		), .Z(n_3633));
	notech_and4 i_80353978(.A(n_241159492), .B(n_240859489), .C(n_240459485)
		, .D(n_240159482), .Z(n_3632));
	notech_and3 i_30008(.A(n_3810), .B(n_30352), .C(n_29633), .Z(n_29967));
	notech_nand2 i_30693(.A(n_19029), .B(n_26755), .Z(n_29282));
	notech_nao3 i_75632091(.A(n_62868), .B(n_27044), .C(n_3690), .Z(n_3630)
		);
	notech_or4 i_75532092(.A(n_26889), .B(instrc[92]), .C(n_29638), .D(n_26725
		), .Z(n_3629));
	notech_and4 i_75432093(.A(n_30973), .B(n_6888902), .C(n_29642), .D(instrc
		[90]), .Z(n_3628));
	notech_and4 i_75332094(.A(n_56888), .B(n_3706), .C(all_cnt[0]), .D(n_29641
		), .Z(n_3627));
	notech_and4 i_75232095(.A(n_29633), .B(n_30952), .C(n_27852), .D(instrc[
		102]), .Z(n_3626));
	notech_nor2 i_14732594(.A(n_3627), .B(n_3626), .Z(n_3625));
	notech_and4 i_32132466(.A(n_3731), .B(n_3629), .C(n_3720), .D(n_27041), 
		.Z(n_3624));
	notech_and4 i_32032467(.A(n_32446), .B(n_27085), .C(n_30987), .D(n_16879899
		), .Z(n_3623));
	notech_and4 i_31932468(.A(n_30905), .B(n_3828), .C(n_27035), .D(n_3829),
		 .Z(n_3622));
	notech_and3 i_12132620(.A(n_32309), .B(n_3630), .C(n_32361), .Z(n_3621)
		);
	notech_nao3 i_73632107(.A(calc_sz[1]), .B(n_314191682), .C(n_56970), .Z(n_3620
		));
	notech_or2 i_71432125(.A(n_306891755), .B(n_32380), .Z(n_3615));
	notech_and2 i_30332480(.A(n_3758), .B(n_3615), .Z(n_3613));
	notech_nao3 i_13532606(.A(n_319191632), .B(n_62892), .C(n_246791942), .Z
		(n_3610));
	notech_ao4 i_22957(.A(n_26601), .B(n_60933), .C(n_3613), .D(n_3759), .Z(n_3609
		));
	notech_or4 i_29432489(.A(n_60893), .B(n_2893), .C(reps[2]), .D(n_27377),
		 .Z(n_3603));
	notech_and2 i_70632133(.A(n_3917), .B(n_3603), .Z(n_3602));
	notech_ao4 i_70532134(.A(n_3602), .B(n_60257), .C(n_27753), .D(n_27580),
		 .Z(n_3598));
	notech_or4 i_33632456(.A(opa[2]), .B(opa[5]), .C(n_3784), .D(n_3781), .Z
		(n_3597));
	notech_ao3 i_6730025(.A(n_3632), .B(n_277959860), .C(n_3633), .Z(n_3596)
		);
	notech_and2 i_67932159(.A(n_3597), .B(n_27025), .Z(n_3595));
	notech_and2 i_67432164(.A(n_3828), .B(n_27035), .Z(n_3594));
	notech_and3 i_15532586(.A(n_26702), .B(n_3852), .C(n_3620), .Z(n_3593)
		);
	notech_and2 i_27232506(.A(n_29734), .B(n_29735), .Z(n_30937));
	notech_or4 i_198132691(.A(tcmp), .B(n_26891), .C(n_29632), .D(n_29663), 
		.Z(n_27580));
	notech_nand3 i_15632585(.A(n_3609), .B(n_27746), .C(n_3610), .Z(n_3590)
		);
	notech_or2 i_31232828(.A(n_56979), .B(n_3695), .Z(n_3589));
	notech_or4 i_31332829(.A(calc_sz[3]), .B(calc_sz[2]), .C(n_2938), .D(n_3695
		), .Z(n_3588));
	notech_and2 i_25675(.A(n_29639), .B(n_29641), .Z(n_30961));
	notech_and2 i_25660(.A(n_29632), .B(n_29663), .Z(n_30930));
	notech_and4 i_25212(.A(n_60122), .B(n_60257), .C(n_32586), .D(n_26841), 
		.Z(n_30352));
	notech_or4 i_43632711(.A(all_cnt[2]), .B(n_27042), .C(n_17107), .D(n_27853
		), .Z(n_30344));
	notech_or4 i_36232713(.A(n_32569), .B(n_32581), .C(n_30361), .D(n_3804),
		 .Z(n_30359));
	notech_and4 i_123733903(.A(n_3584), .B(n_3582), .C(n_3580), .D(n_316960250
		), .Z(n_3586));
	notech_ao4 i_123233908(.A(n_22309), .B(n_28627), .C(n_28076), .D(n_29005
		), .Z(n_3584));
	notech_ao4 i_123433906(.A(n_22594), .B(n_28772), .C(n_22591), .D(n_28740
		), .Z(n_3582));
	notech_ao4 i_123533905(.A(n_22590), .B(n_29732), .C(n_22582), .D(n_28637
		), .Z(n_3580));
	notech_and4 i_124333897(.A(n_357591298), .B(n_357391300), .C(n_357291301
		), .D(n_317660257), .Z(n_3579));
	notech_ao4 i_123833902(.A(n_22585), .B(n_28911), .C(n_22572), .D(n_28652
		), .Z(n_357591298));
	notech_ao4 i_124033900(.A(n_22571), .B(n_56302), .C(n_23040), .D(n_28685
		), .Z(n_357391300));
	notech_ao4 i_124133899(.A(n_55773), .B(n_29731), .C(n_57920), .D(n_27694
		), .Z(n_357291301));
	notech_and4 i_125033890(.A(n_356891305), .B(n_356691307), .C(n_356591308
		), .D(n_318360264), .Z(n_357091303));
	notech_ao4 i_124533895(.A(n_55764), .B(n_27655), .C(n_57859), .D(n_28681
		), .Z(n_356891305));
	notech_ao4 i_124733893(.A(n_27781), .B(n_28720), .C(n_57512), .D(n_28804
		), .Z(n_356691307));
	notech_ao4 i_124833892(.A(n_57121), .B(n_28835), .C(n_57155), .D(n_56154
		), .Z(n_356591308));
	notech_and4 i_125733883(.A(n_356291311), .B(n_356191312), .C(n_355991314
		), .D(n_355891315), .Z(n_356491309));
	notech_ao4 i_125133889(.A(n_57165), .B(n_57625), .C(n_57848), .D(n_55992
		), .Z(n_356291311));
	notech_ao4 i_125233888(.A(n_57498), .B(n_29733), .C(n_22313), .D(n_59259
		), .Z(n_356191312));
	notech_ao4 i_125433886(.A(n_23059), .B(n_27899), .C(n_57533), .D(nbus_11295
		[2]), .Z(n_355991314));
	notech_ao4 i_125533885(.A(n_57552), .B(n_312560206), .C(n_22322), .D(n_355691317
		), .Z(n_355891315));
	notech_ao4 i_125933881(.A(n_22322), .B(n_27038), .C(n_57143), .D(nbus_11310
		[2]), .Z(n_355791316));
	notech_nand2 i_126033880(.A(n_57552), .B(n_27038), .Z(n_355691317));
	notech_and4 i_126733874(.A(n_355291321), .B(n_355091323), .C(n_354991324
		), .D(n_320060281), .Z(n_355491319));
	notech_ao4 i_126133879(.A(n_22309), .B(n_28628), .C(n_22313), .D(n_59223
		), .Z(n_355291321));
	notech_ao4 i_126433877(.A(n_28076), .B(n_29006), .C(n_22594), .D(n_28773
		), .Z(n_355091323));
	notech_ao4 i_126533876(.A(n_22591), .B(n_28741), .C(n_22590), .D(n_29730
		), .Z(n_354991324));
	notech_and4 i_127333868(.A(n_354691327), .B(n_354491329), .C(n_354391330
		), .D(n_321691616), .Z(n_354891325));
	notech_ao4 i_126833873(.A(n_22579), .B(n_28880), .C(n_22585), .D(n_28912
		), .Z(n_354691327));
	notech_ao4 i_127033871(.A(n_22572), .B(n_28653), .C(n_22571), .D(n_56311
		), .Z(n_354491329));
	notech_ao4 i_127133870(.A(n_23040), .B(n_28686), .C(n_55773), .D(n_29729
		), .Z(n_354391330));
	notech_and4 i_128133861(.A(n_353991334), .B(n_353791336), .C(n_353691337
		), .D(n_324291609), .Z(n_354191332));
	notech_ao4 i_127533866(.A(n_23031), .B(n_27678), .C(n_55764), .D(n_27656
		), .Z(n_353991334));
	notech_ao4 i_127833864(.A(n_57859), .B(n_27513), .C(n_27781), .D(n_28723
		), .Z(n_353791336));
	notech_ao4 i_127933863(.A(n_57848), .B(n_55983), .C(n_57512), .D(n_28805
		), .Z(n_353691337));
	notech_and4 i_128833854(.A(n_353391340), .B(n_353291341), .C(n_353091343
		), .D(n_352991344), .Z(n_353591338));
	notech_ao4 i_128233860(.A(n_57498), .B(n_29728), .C(n_57121), .D(n_28836
		), .Z(n_353391340));
	notech_ao4 i_128333859(.A(n_57155), .B(n_56181), .C(n_57165), .D(n_57635
		), .Z(n_353291341));
	notech_ao4 i_128533857(.A(n_57524), .B(n_27901), .C(n_57533), .D(nbus_11295
		[3]), .Z(n_353091343));
	notech_ao4 i_128633856(.A(n_57563), .B(n_312660207), .C(n_22322), .D(n_352791346
		), .Z(n_352991344));
	notech_ao4 i_129033852(.A(n_3788), .B(n_22322), .C(n_57143), .D(nbus_11310
		[3]), .Z(n_352891345));
	notech_nand2 i_129133851(.A(n_57563), .B(n_3788), .Z(n_352791346));
	notech_and4 i_129733845(.A(n_352391350), .B(n_352191352), .C(n_352091353
		), .D(n_328191592), .Z(n_352591348));
	notech_ao4 i_129233850(.A(n_22309), .B(n_28629), .C(n_22313), .D(n_27986
		), .Z(n_352391350));
	notech_ao4 i_129433848(.A(n_28076), .B(n_29007), .C(n_22594), .D(n_28774
		), .Z(n_352191352));
	notech_ao4 i_129533847(.A(n_22591), .B(n_28742), .C(n_22590), .D(n_29727
		), .Z(n_352091353));
	notech_and4 i_130333839(.A(n_351791356), .B(n_351591358), .C(n_351491359
		), .D(n_328891585), .Z(n_351991354));
	notech_ao4 i_129833844(.A(n_22579), .B(n_28881), .C(n_22585), .D(n_28913
		), .Z(n_351791356));
	notech_ao4 i_130033842(.A(n_22572), .B(n_28654), .C(n_22571), .D(n_56320
		), .Z(n_351591358));
	notech_ao4 i_130133841(.A(n_23040), .B(n_28687), .C(n_55773), .D(n_29726
		), .Z(n_351491359));
	notech_and4 i_131033832(.A(n_351091363), .B(n_350891365), .C(n_350791366
		), .D(n_329591578), .Z(n_351291361));
	notech_ao4 i_130533837(.A(n_23031), .B(n_27679), .C(n_55764), .D(n_27657
		), .Z(n_351091363));
	notech_ao4 i_130733835(.A(n_57859), .B(n_27514), .C(n_27781), .D(n_28725
		), .Z(n_350891365));
	notech_ao4 i_130833834(.A(n_57848), .B(n_56064), .C(n_57512), .D(n_28806
		), .Z(n_350791366));
	notech_and4 i_131733825(.A(n_350491369), .B(n_350391370), .C(n_350191372
		), .D(n_350091373), .Z(n_350691367));
	notech_ao4 i_131133831(.A(n_57498), .B(n_56055), .C(n_57121), .D(n_28837
		), .Z(n_350491369));
	notech_ao4 i_131233830(.A(n_57155), .B(n_56221), .C(n_57165), .D(n_57644
		), .Z(n_350391370));
	notech_ao4 i_131433828(.A(n_57524), .B(n_27902), .C(n_57533), .D(nbus_11295
		[4]), .Z(n_350191372));
	notech_ao4 i_131533827(.A(n_57574), .B(n_312760208), .C(n_22322), .D(n_349891375
		), .Z(n_350091373));
	notech_ao4 i_131933823(.A(n_3789), .B(n_22322), .C(n_57143), .D(nbus_11310
		[4]), .Z(n_349991374));
	notech_nand2 i_132033822(.A(n_57574), .B(n_3789), .Z(n_349891375));
	notech_and4 i_132633816(.A(n_349491379), .B(n_349291381), .C(n_349191382
		), .D(n_331291561), .Z(n_349691377));
	notech_ao4 i_132133821(.A(n_22309), .B(n_28632), .C(n_22313), .D(n_27989
		), .Z(n_349491379));
	notech_ao4 i_132333819(.A(n_28076), .B(n_29008), .C(n_22594), .D(n_28776
		), .Z(n_349291381));
	notech_ao4 i_132433818(.A(n_22591), .B(n_28744), .C(n_22590), .D(n_29724
		), .Z(n_349191382));
	notech_and4 i_133433810(.A(n_348891385), .B(n_348691387), .C(n_348591388
		), .D(n_331991554), .Z(n_349091383));
	notech_ao4 i_132733815(.A(n_22579), .B(n_28883), .C(n_22585), .D(n_28915
		), .Z(n_348891385));
	notech_ao4 i_132933813(.A(n_22572), .B(n_28658), .C(n_22571), .D(n_56338
		), .Z(n_348691387));
	notech_ao4 i_133033812(.A(n_23040), .B(n_28688), .C(n_57533), .D(nbus_11295
		[6]), .Z(n_348591388));
	notech_and4 i_134133803(.A(n_348191392), .B(n_347991394), .C(n_347891395
		), .D(n_332691547), .Z(n_348391390));
	notech_ao4 i_133633808(.A(n_57920), .B(n_27695), .C(n_23031), .D(n_27681
		), .Z(n_348191392));
	notech_ao4 i_133833806(.A(n_55764), .B(n_27658), .C(n_57859), .D(n_27515
		), .Z(n_347991394));
	notech_ao4 i_133933805(.A(n_27781), .B(n_28726), .C(n_57848), .D(n_56082
		), .Z(n_347891395));
	notech_and4 i_134833796(.A(n_347591398), .B(n_347491399), .C(n_347291401
		), .D(n_347191402), .Z(n_347791396));
	notech_ao4 i_134233802(.A(n_57512), .B(n_28807), .C(n_57498), .D(n_29723
		), .Z(n_347591398));
	notech_ao4 i_134333801(.A(n_57121), .B(n_28838), .C(n_57155), .D(n_56248
		), .Z(n_347491399));
	notech_ao4 i_134533799(.A(n_57165), .B(n_57662), .C(n_57524), .D(n_27909
		), .Z(n_347291401));
	notech_ao4 i_134633798(.A(n_57592), .B(n_312860209), .C(n_341191462), .D
		(n_346991404), .Z(n_347191402));
	notech_ao4 i_135033794(.A(nbus_11310[6]), .B(n_57143), .C(n_22322), .D(n_27060
		), .Z(n_347091403));
	notech_or2 i_135133793(.A(n_22322), .B(opa[6]), .Z(n_346991404));
	notech_and4 i_135733787(.A(n_57948), .B(n_346591408), .C(n_346391410), .D
		(n_346291411), .Z(n_346791406));
	notech_ao4 i_135233792(.A(n_27782), .B(n_28670), .C(n_22309), .D(n_28634
		), .Z(n_346591408));
	notech_ao4 i_135433790(.A(n_22313), .B(n_56100), .C(n_28076), .D(n_29009
		), .Z(n_346391410));
	notech_ao4 i_135533789(.A(n_22594), .B(n_28777), .C(n_22591), .D(n_28745
		), .Z(n_346291411));
	notech_and4 i_136433780(.A(n_345991414), .B(n_345891415), .C(n_345691417
		), .D(n_345591418), .Z(n_346191412));
	notech_ao4 i_135833786(.A(n_22590), .B(n_29722), .C(n_22582), .D(n_28639
		), .Z(n_345991414));
	notech_ao4 i_135933785(.A(n_22579), .B(n_28884), .C(n_22585), .D(n_28916
		), .Z(n_345891415));
	notech_ao4 i_136133783(.A(n_22572), .B(n_28659), .C(n_22571), .D(n_56347
		), .Z(n_345691417));
	notech_ao4 i_136233782(.A(n_23040), .B(n_28689), .C(n_55773), .D(n_29721
		), .Z(n_345591418));
	notech_and4 i_137133773(.A(n_345191422), .B(n_344991424), .C(n_344891425
		), .D(n_335791516), .Z(n_345391420));
	notech_ao4 i_136633778(.A(n_23031), .B(n_27682), .C(n_55764), .D(n_27659
		), .Z(n_345191422));
	notech_ao4 i_136833776(.A(n_57859), .B(n_27516), .C(n_27781), .D(n_28727
		), .Z(n_344991424));
	notech_ao4 i_136933775(.A(n_57512), .B(n_28808), .C(n_57498), .D(n_29614
		), .Z(n_344891425));
	notech_and4 i_137833766(.A(n_344591428), .B(n_344491429), .C(n_344291431
		), .D(n_344191432), .Z(n_344791426));
	notech_ao4 i_137233772(.A(n_57121), .B(n_28839), .C(n_57848), .D(n_56109
		), .Z(n_344591428));
	notech_ao4 i_137333771(.A(n_57533), .B(nbus_11295[7]), .C(n_57155), .D(n_56275
		), .Z(n_344491429));
	notech_ao4 i_137533769(.A(n_57165), .B(n_57671), .C(n_57524), .D(n_27910
		), .Z(n_344291431));
	notech_ao4 i_137633768(.A(n_313060211), .B(n_57957), .C(n_312960210), .D
		(n_343791436), .Z(n_344191432));
	notech_ao4 i_138133763(.A(nbus_11310[7]), .B(n_57143), .C(n_22322), .D(n_27062
		), .Z(n_343891435));
	notech_or4 i_138333761(.A(n_32384), .B(n_27879), .C(n_26782), .D(opa[7])
		, .Z(n_343791436));
	notech_and3 i_10035010(.A(n_57524), .B(n_3902), .C(n_3903), .Z(n_81910939
		));
	notech_nand3 i_200833145(.A(n_343291441), .B(n_343491439), .C(n_337791496
		), .Z(n_343591438));
	notech_ao4 i_200533148(.A(n_211169123), .B(n_59991), .C(n_308091743), .D
		(n_28091), .Z(n_343491439));
	notech_ao4 i_200633147(.A(n_58444), .B(n_55992), .C(n_343270443), .D(n_344366972
		), .Z(n_343291441));
	notech_ao4 i_200933144(.A(n_57552), .B(n_313460215), .C(n_313360214), .D
		(n_313260213), .Z(n_342991444));
	notech_ao4 i_201433139(.A(n_56463), .B(n_344466973), .C(n_59435), .D(n_29733
		), .Z(n_342591448));
	notech_ao4 i_201533138(.A(n_27757), .B(n_315160232), .C(n_315060231), .D
		(n_32327), .Z(n_342491449));
	notech_nand3 i_201233141(.A(n_338291491), .B(n_338191492), .C(n_338391490
		), .Z(n_342391450));
	notech_nand3 i_201733136(.A(n_60303), .B(n_1904), .C(\opa_12[2] ), .Z(n_341891455
		));
	notech_xor2 i_133135089(.A(opa[6]), .B(n_341691457), .Z(n_341791456));
	notech_xor2 i_5435056(.A(opa[5]), .B(opa[7]), .Z(n_341691457));
	notech_xor2 i_71635095(.A(n_341491459), .B(n_341391460), .Z(n_341591458)
		);
	notech_xor2 i_15634955(.A(opa[3]), .B(opa[4]), .Z(n_341491459));
	notech_xor2 i_1335079(.A(n_57552), .B(n_307947775), .Z(n_341391460));
	notech_and2 i_4235068(.A(n_27885), .B(n_57583), .Z(n_341191462));
	notech_ao4 i_206433089(.A(n_320063467), .B(n_3786), .C(n_32263), .D(n_26965
		), .Z(n_340991464));
	notech_ao4 i_206533088(.A(n_107111189), .B(n_29655), .C(n_58220), .D(n_3893
		), .Z(n_340891465));
	notech_and4 i_207033083(.A(n_339491479), .B(n_340691467), .C(n_339391480
		), .D(n_339591478), .Z(n_340791466));
	notech_ao4 i_206733086(.A(n_61115), .B(n_316660247), .C(n_25397), .D(n_340391470
		), .Z(n_340691467));
	notech_ao4 i_207233081(.A(n_303991784), .B(n_25619), .C(n_1864), .D(n_305047803
		), .Z(n_340491469));
	notech_nao3 i_207333080(.A(instrc[107]), .B(n_32612), .C(n_116368180), .Z
		(n_340391470));
	notech_or4 i_111534020(.A(n_27925), .B(n_32643), .C(n_125461537), .D(n_27641
		), .Z(n_339591478));
	notech_or4 i_111434021(.A(n_60893), .B(n_61117), .C(n_1868), .D(n_25625)
		, .Z(n_339491479));
	notech_nao3 i_111334022(.A(n_26776), .B(n_316560246), .C(n_59322), .Z(n_339391480
		));
	notech_ao4 i_34287(.A(n_305047803), .B(n_27105), .C(n_25615), .D(n_330763524
		), .Z(n_25613));
	notech_or4 i_106934066(.A(calc_sz[1]), .B(n_56970), .C(n_60263), .D(n_26634
		), .Z(n_338791486));
	notech_or2 i_105034085(.A(n_56979), .B(n_313160212), .Z(n_338391490));
	notech_or4 i_104934086(.A(n_32446), .B(n_60263), .C(n_57772), .D(n_3904)
		, .Z(n_338291491));
	notech_or4 i_104834087(.A(n_26789), .B(n_56829), .C(n_56513), .D(n_59259
		), .Z(n_338191492));
	notech_ao4 i_105334082(.A(n_27058), .B(n_27059), .C(n_305291771), .D(n_1448
		), .Z(n_338091493));
	notech_nand2 i_105634079(.A(nPF), .B(n_26593), .Z(n_337791496));
	notech_or4 i_9378(.A(n_25615), .B(n_62824), .C(n_60910), .D(n_60263), .Z
		(n_337091503));
	notech_nao3 i_40534723(.A(n_2950), .B(\nbus_14520[7] ), .C(n_57933), .Z(n_335791516
		));
	notech_nao3 i_37134754(.A(n_2947), .B(n_10907), .C(n_19093), .Z(n_332691547
		));
	notech_nao3 i_37834747(.A(n_295591839), .B(nbus_163[6]), .C(n_27907), .Z
		(n_331991554));
	notech_nand3 i_38534740(.A(n_27784), .B(n_2944), .C(nbus_158[6]), .Z(n_331291561
		));
	notech_nao3 i_33834785(.A(n_2950), .B(\nbus_14520[4] ), .C(n_57933), .Z(n_329591578
		));
	notech_nao3 i_34534778(.A(n_295591839), .B(nbus_163[4]), .C(n_27907), .Z
		(n_328891585));
	notech_nand3 i_35334771(.A(n_27784), .B(n_2944), .C(nbus_158[4]), .Z(n_328191592
		));
	notech_nao3 i_30634816(.A(n_2950), .B(\nbus_14520[3] ), .C(n_57933), .Z(n_324291609
		));
	notech_nao3 i_31334809(.A(n_295591839), .B(nbus_163[3]), .C(n_27907), .Z
		(n_321691616));
	notech_nand3 i_32034802(.A(n_27784), .B(n_2944), .C(nbus_158[3]), .Z(n_320060281
		));
	notech_nao3 i_27034847(.A(cr2_reg[2]), .B(n_57992), .C(n_2949), .Z(n_318360264
		));
	notech_nao3 i_27734840(.A(nbus_162[2]), .B(n_2956), .C(n_59451), .Z(n_317660257
		));
	notech_nand3 i_28734833(.A(n_27784), .B(n_2944), .C(nbus_158[2]), .Z(n_316960250
		));
	notech_and4 i_15534956(.A(n_2895), .B(n_304784038), .C(n_340491469), .D(n_137861661
		), .Z(n_316660247));
	notech_nand2 i_8935021(.A(n_5380), .B(n_26779), .Z(n_316560246));
	notech_ao4 i_8435026(.A(n_312447734), .B(n_56463), .C(n_59419), .D(n_29733
		), .Z(n_315160232));
	notech_ao4 i_8535025(.A(n_312347735), .B(n_27757), .C(n_60868), .D(n_29733
		), .Z(n_315060231));
	notech_nand3 i_106634069(.A(n_62826), .B(opc[2]), .C(n_27757), .Z(n_314760228
		));
	notech_or4 i_106534070(.A(n_62856), .B(n_60933), .C(n_57552), .D(n_27757
		), .Z(n_314660227));
	notech_and3 i_10235008(.A(n_314760228), .B(n_58316), .C(n_314660227), .Z
		(n_314560226));
	notech_ao3 i_10335007(.A(n_56959), .B(n_56941), .C(n_32384), .Z(n_314360224
		));
	notech_ao4 i_3635074(.A(n_27746), .B(n_55992), .C(n_57552), .D(n_306991754
		), .Z(n_314260223));
	notech_ao4 i_8635024(.A(n_26602), .B(n_60023), .C(n_32459), .D(n_29733),
		 .Z(n_313860219));
	notech_and3 i_12034990(.A(n_26606), .B(n_338791486), .C(n_57314), .Z(n_313460215
		));
	notech_ao4 i_11934991(.A(n_314560226), .B(n_26789), .C(n_314260223), .D(n_314360224
		), .Z(n_313360214));
	notech_ao4 i_235086(.A(n_2480), .B(n_62892), .C(n_56829), .D(n_32294), .Z
		(n_313260213));
	notech_ao4 i_11834992(.A(n_313860219), .B(n_27754), .C(n_57823), .D(n_341891455
		), .Z(n_313160212));
	notech_and4 i_14734964(.A(n_337091503), .B(n_343891435), .C(n_3889), .D(n_81910939
		), .Z(n_313060211));
	notech_and2 i_6435046(.A(n_57592), .B(n_341191462), .Z(n_312960210));
	notech_and2 i_14834963(.A(n_347091403), .B(n_1884), .Z(n_312860209));
	notech_and2 i_14934962(.A(n_1884), .B(n_349991374), .Z(n_312760208));
	notech_and2 i_15034961(.A(n_1884), .B(n_352891345), .Z(n_312660207));
	notech_and2 i_15134960(.A(n_1884), .B(n_355791316), .Z(n_312560206));
	notech_and4 i_126537037(.A(n_311760198), .B(n_311960200), .C(n_311660197
		), .D(n_297460055), .Z(n_312160202));
	notech_ao4 i_125637046(.A(n_54912649), .B(n_101413114), .C(n_55886), .D(nbus_11295
		[10]), .Z(n_311960200));
	notech_ao4 i_125737045(.A(n_60023), .B(n_53612636), .C(n_53412634), .D(n_29169
		), .Z(n_311760198));
	notech_and4 i_126437038(.A(n_311460195), .B(n_311260193), .C(n_297760058
		), .D(n_298060061), .Z(n_311660197));
	notech_ao4 i_126037042(.A(n_54212642), .B(n_57552), .C(n_54012640), .D(n_29252
		), .Z(n_311460195));
	notech_ao4 i_126237040(.A(n_388560287), .B(n_55992), .C(n_33012430), .D(n_28989
		), .Z(n_311260193));
	notech_and4 i_127037032(.A(n_310860189), .B(n_298660067), .C(n_310660187
		), .D(n_298360064), .Z(n_311060191));
	notech_ao4 i_126637036(.A(n_33312433), .B(n_29010), .C(n_54512645), .D(n_56154
		), .Z(n_310860189));
	notech_ao4 i_126837034(.A(n_26948), .B(n_28107), .C(n_19312293), .D(n_28115
		), .Z(n_310660187));
	notech_and4 i_127537027(.A(n_310360184), .B(n_310160182), .C(n_298960070
		), .D(n_299260073), .Z(n_310560186));
	notech_ao4 i_127137031(.A(n_3886), .B(n_28091), .C(n_3887), .D(n_29054),
		 .Z(n_310360184));
	notech_ao4 i_127337029(.A(n_8812188), .B(n_29736), .C(n_54912649), .D(n_295860039
		), .Z(n_310160182));
	notech_nao3 i_4238192(.A(instrc[107]), .B(n_295760038), .C(n_296760048),
		 .Z(n_8812188));
	notech_ao4 i_127737025(.A(n_60841), .B(n_28051), .C(n_57710), .D(n_58009
		), .Z(n_310060181));
	notech_nao3 i_131038221(.A(instrc[107]), .B(n_295960040), .C(n_296760048
		), .Z(n_17012270));
	notech_ao4 i_138036924(.A(n_330763524), .B(n_305047803), .C(n_27105), .D
		(n_296160042), .Z(n_309660177));
	notech_and3 i_44638231(.A(mask8b[1]), .B(n_309160172), .C(n_27541), .Z(n_18912289
		));
	notech_nand3 i_44838230(.A(mask8b[1]), .B(n_309160172), .C(mask8b[0]), .Z
		(n_19312293));
	notech_and2 i_138336921(.A(mask8b[1]), .B(mask8b[0]), .Z(n_309460175));
	notech_ao3 i_45038229(.A(mask8b[0]), .B(n_309160172), .C(mask8b[1]), .Z(n_19512295
		));
	notech_and4 i_3338201(.A(mask8b[2]), .B(n_2885), .C(n_3794), .D(n_61154)
		, .Z(n_309160172));
	notech_or4 i_39338238(.A(n_27917), .B(n_59435), .C(n_60263), .D(n_26782)
		, .Z(n_33012430));
	notech_or4 i_39738236(.A(n_62826), .B(n_60910), .C(n_60263), .D(n_26965)
		, .Z(n_33312433));
	notech_or4 i_42138232(.A(n_27917), .B(n_59435), .C(n_60268), .D(n_27896)
		, .Z(n_33412434));
	notech_or4 i_39638237(.A(n_25349), .B(n_60933), .C(n_60910), .D(n_60268)
		, .Z(n_33512435));
	notech_nand2 i_170436602(.A(n_27052), .B(n_27056), .Z(n_309060171));
	notech_or4 i_36938247(.A(n_27917), .B(n_62832), .C(n_62824), .D(n_60268)
		, .Z(n_52112621));
	notech_or4 i_37738244(.A(n_25619), .B(n_62824), .C(n_60910), .D(n_60268)
		, .Z(n_53412634));
	notech_or4 i_37838243(.A(n_305047803), .B(n_62824), .C(n_60910), .D(n_60268
		), .Z(n_53512635));
	notech_or2 i_37538246(.A(instrc[107]), .B(n_296760048), .Z(n_53612636)
		);
	notech_nao3 i_38038241(.A(n_57899), .B(n_27052), .C(n_308760168), .Z(n_54012640
		));
	notech_and2 i_170536601(.A(n_57899), .B(n_27052), .Z(n_308960170));
	notech_or4 i_37938242(.A(n_25619), .B(n_62832), .C(n_60933), .D(n_60268)
		, .Z(n_54212642));
	notech_nand2 i_170636600(.A(n_19137), .B(n_19117), .Z(n_308860169));
	notech_nand2 i_37638245(.A(instrc[107]), .B(n_27071), .Z(n_54912649));
	notech_nao3 i_2538209(.A(n_19117), .B(n_26985), .C(n_25641), .Z(n_308760168
		));
	notech_ao4 i_194736361(.A(n_57976), .B(n_28299), .C(n_60841), .D(n_28493
		), .Z(n_308360164));
	notech_ao4 i_194836360(.A(n_58009), .B(n_27868), .C(n_56463), .D(n_56163
		), .Z(n_308260163));
	notech_and2 i_195236356(.A(n_308060161), .B(n_307960160), .Z(n_308160162
		));
	notech_ao4 i_195036358(.A(n_56396), .B(n_28168), .C(n_56391), .D(n_28397
		), .Z(n_308060161));
	notech_ao4 i_195136357(.A(n_59344), .B(n_28528), .C(n_56367), .D(n_28333
		), .Z(n_307960160));
	notech_and4 i_196036348(.A(n_307660157), .B(n_307560156), .C(n_307360154
		), .D(n_307260153), .Z(n_307860159));
	notech_ao4 i_195436354(.A(n_56452), .B(n_28267), .C(n_58020), .D(n_28461
		), .Z(n_307660157));
	notech_ao4 i_195536353(.A(n_56443), .B(n_28233), .C(n_56432), .D(n_28200
		), .Z(n_307560156));
	notech_ao4 i_195736351(.A(n_56903), .B(n_29720), .C(n_56423), .D(n_28365
		), .Z(n_307360154));
	notech_ao4 i_195836350(.A(n_56414), .B(n_28429), .C(n_56405), .D(n_28571
		), .Z(n_307260153));
	notech_and2 i_26367158(.A(n_60537), .B(n_349480995), .Z(n_108582086));
	notech_nao3 i_50693(.A(n_116778671), .B(n_126078764), .C(n_108582086), .Z
		(\nbus_11330[16] ));
	notech_ao4 i_48388(.A(n_315963426), .B(n_29793), .C(n_57966), .D(n_135041965
		), .Z(\nbus_11301[0] ));
	notech_or4 i_27267149(.A(n_60964), .B(n_60953), .C(n_62832), .D(n_3880),
		 .Z(n_108782088));
	notech_and4 i_6367338(.A(n_304084031), .B(n_313884129), .C(n_112441739),
		 .D(n_108782088), .Z(n_108982090));
	notech_ao4 i_49425(.A(n_29793), .B(n_121282213), .C(n_108982090), .D(n_135041965
		), .Z(\nbus_11313[16] ));
	notech_and4 i_6467337(.A(n_2676), .B(n_23627), .C(n_310084091), .D(n_60051
		), .Z(n_109382094));
	notech_ao4 i_49423(.A(n_109382094), .B(n_135041965), .C(n_29793), .D(n_326684257
		), .Z(\nbus_11313[5] ));
	notech_nor2 i_7656(.A(n_32476), .B(n_57403), .Z(n_109482095));
	notech_and3 i_31767104(.A(n_18981), .B(n_32551), .C(read_ack), .Z(n_109582096
		));
	notech_or4 i_56293(.A(n_109582096), .B(n_121682217), .C(n_121582216), .D
		(n_109482095), .Z(\nbus_11377[0] ));
	notech_nao3 i_5997(.A(over_seg[5]), .B(n_60542), .C(n_58683), .Z(n_109682097
		));
	notech_nor2 i_33567088(.A(n_322984220), .B(n_29655), .Z(n_109782098));
	notech_or2 i_33667087(.A(n_26860), .B(sema_rw), .Z(n_109882099));
	notech_or4 i_53810(.A(n_109782098), .B(n_61131), .C(n_122182222), .D(n_26988
		), .Z(n_21582));
	notech_and2 i_40967018(.A(imm[6]), .B(n_329263509), .Z(n_109982100));
	notech_and2 i_41167016(.A(imm[7]), .B(n_329863515), .Z(n_110082101));
	notech_and4 i_41367014(.A(n_59408), .B(n_59397), .C(n_246991940), .D(imm
		[8]), .Z(n_110182102));
	notech_and4 i_41567012(.A(n_59408), .B(n_59398), .C(n_246991940), .D(imm
		[9]), .Z(n_110282103));
	notech_and4 i_41767010(.A(n_59408), .B(n_59398), .C(n_246991940), .D(imm
		[11]), .Z(n_110382104));
	notech_and4 i_41967008(.A(n_59408), .B(n_59398), .C(n_246991940), .D(imm
		[12]), .Z(n_110482105));
	notech_and4 i_42167006(.A(n_59408), .B(n_59397), .C(n_246991940), .D(imm
		[13]), .Z(n_110582106));
	notech_and4 i_42367004(.A(n_59408), .B(n_59397), .C(n_246991940), .D(imm
		[14]), .Z(n_110682107));
	notech_and4 i_42567002(.A(n_59407), .B(n_59397), .C(n_246991940), .D(imm
		[15]), .Z(n_110782108));
	notech_and4 i_43966988(.A(n_59407), .B(n_59397), .C(n_246991940), .D(imm
		[22]), .Z(n_110882109));
	notech_ao4 i_80866619(.A(n_179382794), .B(n_26781), .C(n_56205), .D(n_110882109
		), .Z(n_110982110));
	notech_nand2 i_2312940(.A(n_123082231), .B(n_26861), .Z(n_26058));
	notech_ao4 i_92866499(.A(n_56205), .B(n_110782108), .C(n_330363520), .D(n_26781
		), .Z(n_111882119));
	notech_or4 i_92766500(.A(n_60312), .B(n_26964), .C(n_19079), .D(n_28104)
		, .Z(n_112782128));
	notech_or4 i_1612933(.A(n_111882119), .B(n_123782238), .C(n_26863), .D(n_26862
		), .Z(n_26023));
	notech_ao4 i_94766480(.A(n_56205), .B(n_110682107), .C(n_330363520), .D(n_26781
		), .Z(n_112882129));
	notech_or4 i_94666481(.A(n_60312), .B(n_26964), .C(n_19079), .D(n_28103)
		, .Z(n_113782138));
	notech_or4 i_1512932(.A(n_112882129), .B(n_124582246), .C(n_26865), .D(n_26864
		), .Z(n_26018));
	notech_ao4 i_96666461(.A(n_56205), .B(n_110582106), .C(n_330363520), .D(n_26781
		), .Z(n_113882139));
	notech_or4 i_96566462(.A(n_60292), .B(n_26964), .C(n_19079), .D(n_28102)
		, .Z(n_114782148));
	notech_or4 i_1412931(.A(n_113882139), .B(n_125382254), .C(n_26867), .D(n_26866
		), .Z(n_26013));
	notech_ao4 i_98666442(.A(n_56205), .B(n_110482105), .C(n_330363520), .D(n_26781
		), .Z(n_114882149));
	notech_or4 i_98566443(.A(n_60312), .B(n_26964), .C(n_19079), .D(n_28101)
		, .Z(n_115782158));
	notech_or4 i_1312930(.A(n_114882149), .B(n_126182262), .C(n_26869), .D(n_26868
		), .Z(n_26008));
	notech_ao4 i_100566423(.A(n_56205), .B(n_110382104), .C(n_330363520), .D
		(n_26781), .Z(n_115882159));
	notech_or4 i_100466424(.A(n_60312), .B(n_26964), .C(n_19079), .D(n_28100
		), .Z(n_116782168));
	notech_or4 i_1212929(.A(n_115882159), .B(n_126982270), .C(n_26871), .D(n_26870
		), .Z(n_26003));
	notech_ao4 i_102466404(.A(n_56204), .B(n_110282103), .C(n_330363520), .D
		(n_26781), .Z(n_116882169));
	notech_or4 i_102366405(.A(n_60312), .B(n_26964), .C(n_19079), .D(n_28098
		), .Z(n_117782178));
	notech_or4 i_1012927(.A(n_116882169), .B(n_127782278), .C(n_26873), .D(n_26872
		), .Z(n_25993));
	notech_ao4 i_104366385(.A(n_56204), .B(n_110182102), .C(n_330363520), .D
		(n_26781), .Z(n_117882179));
	notech_or4 i_104266386(.A(n_60312), .B(n_26964), .C(n_19079), .D(n_28097
		), .Z(n_118782188));
	notech_or4 i_912926(.A(n_117882179), .B(n_128582286), .C(n_26875), .D(n_26874
		), .Z(n_25988));
	notech_ao4 i_106266366(.A(n_56204), .B(n_110082101), .C(n_330363520), .D
		(n_26781), .Z(n_118882189));
	notech_or4 i_106166367(.A(n_60312), .B(n_26964), .C(n_19079), .D(n_28096
		), .Z(n_119782198));
	notech_or4 i_812925(.A(n_118882189), .B(n_129382294), .C(n_26877), .D(n_26876
		), .Z(n_25983));
	notech_ao4 i_108166347(.A(n_83341448), .B(n_109982100), .C(n_330363520),
		 .D(n_26781), .Z(n_119882199));
	notech_or4 i_108066348(.A(n_60292), .B(n_26964), .C(n_19079), .D(n_28095
		), .Z(n_120782208));
	notech_or4 i_712924(.A(n_119882199), .B(n_130182302), .C(n_26879), .D(n_26878
		), .Z(n_25978));
	notech_ao4 i_222685(.A(n_27895), .B(n_130382304), .C(n_60292), .D(n_19043
		), .Z(n_22451));
	notech_nand3 i_24067405(.A(n_60127), .B(n_60292), .C(n_61560), .Z(n_135041965
		));
	notech_and4 i_2967371(.A(n_313784128), .B(n_32656), .C(n_60051), .D(n_60074
		), .Z(n_112441739));
	notech_nand3 i_27767144(.A(n_130882309), .B(n_60127), .C(n_60268), .Z(n_121282213
		));
	notech_nand3 i_32167101(.A(n_58664), .B(n_58662), .C(n_58683), .Z(n_121582216
		));
	notech_nand3 i_32067102(.A(n_309384084), .B(n_187310085), .C(n_26860), .Z
		(n_121682217));
	notech_nand3 i_34067084(.A(n_58664), .B(n_309384084), .C(n_109882099), .Z
		(n_122182222));
	notech_ao4 i_80966618(.A(n_54141156), .B(n_30033), .C(n_328184272), .D(n_29076
		), .Z(n_122482225));
	notech_ao4 i_81066617(.A(n_53341148), .B(nbus_11295[22]), .C(n_53841153)
		, .D(n_30034), .Z(n_122582226));
	notech_ao4 i_81166616(.A(n_58773), .B(n_29108), .C(n_58768), .D(n_30035)
		, .Z(n_122782228));
	notech_ao4 i_81266615(.A(n_52741142), .B(n_28111), .C(n_53641151), .D(n_57742
		), .Z(n_122882229));
	notech_and4 i_81566612(.A(n_122882229), .B(n_122782228), .C(n_122582226)
		, .D(n_122482225), .Z(n_123082231));
	notech_ao4 i_93066497(.A(n_54141156), .B(n_30036), .C(n_40241017), .D(n_29101
		), .Z(n_123182232));
	notech_ao4 i_93166496(.A(n_53641151), .B(n_57671), .C(n_53841153), .D(n_30037
		), .Z(n_123282233));
	notech_ao4 i_93266495(.A(n_58768), .B(n_30039), .C(n_53341148), .D(nbus_11295
		[15]), .Z(n_123482235));
	notech_ao4 i_92966498(.A(n_39041005), .B(n_28941), .C(n_180682807), .D(n_29067
		), .Z(n_123582236));
	notech_nand3 i_93566492(.A(n_112782128), .B(n_123582236), .C(n_123482235
		), .Z(n_123782238));
	notech_ao4 i_94966478(.A(n_54141156), .B(n_30040), .C(n_40241017), .D(n_29100
		), .Z(n_123982240));
	notech_ao4 i_95066477(.A(n_53341148), .B(nbus_11295[14]), .C(n_53841153)
		, .D(n_30041), .Z(n_124082241));
	notech_ao4 i_95166476(.A(n_53641151), .B(n_57662), .C(n_58768), .D(n_30042
		), .Z(n_124282243));
	notech_ao4 i_94866479(.A(n_39041005), .B(n_28940), .C(n_180682807), .D(n_29066
		), .Z(n_124382244));
	notech_nand3 i_95466473(.A(n_113782138), .B(n_124382244), .C(n_124282243
		), .Z(n_124582246));
	notech_ao4 i_96866459(.A(n_54141156), .B(n_30043), .C(n_40241017), .D(n_29099
		), .Z(n_124782248));
	notech_ao4 i_96966458(.A(n_53641151), .B(n_57653), .C(n_53841153), .D(n_30044
		), .Z(n_124882249));
	notech_ao4 i_97066457(.A(n_58768), .B(n_30045), .C(n_53341148), .D(nbus_11295
		[13]), .Z(n_125082251));
	notech_ao4 i_96766460(.A(n_39041005), .B(n_28939), .C(n_180682807), .D(n_29065
		), .Z(n_125182252));
	notech_nand3 i_97366454(.A(n_114782148), .B(n_125182252), .C(n_125082251
		), .Z(n_125382254));
	notech_ao4 i_98866440(.A(n_54141156), .B(n_30046), .C(n_40241017), .D(n_29098
		), .Z(n_125582256));
	notech_ao4 i_98966439(.A(n_53341148), .B(nbus_11295[12]), .C(n_53841153)
		, .D(n_30047), .Z(n_125682257));
	notech_ao4 i_99066438(.A(n_53641151), .B(\nbus_11307[12] ), .C(n_58768),
		 .D(n_30048), .Z(n_125882259));
	notech_ao4 i_98766441(.A(n_39041005), .B(n_28938), .C(n_180682807), .D(n_29064
		), .Z(n_125982260));
	notech_nand3 i_99366435(.A(n_115782158), .B(n_125982260), .C(n_125882259
		), .Z(n_126182262));
	notech_ao4 i_100766421(.A(n_54141156), .B(n_30050), .C(n_40241017), .D(n_29097
		), .Z(n_126382264));
	notech_ao4 i_100866420(.A(n_53341148), .B(nbus_11295[11]), .C(n_53841153
		), .D(n_30051), .Z(n_126482265));
	notech_ao4 i_100966419(.A(n_53641151), .B(n_57635), .C(n_58768), .D(n_30052
		), .Z(n_126682267));
	notech_ao4 i_100666422(.A(n_39041005), .B(n_28937), .C(n_180682807), .D(n_29063
		), .Z(n_126782268));
	notech_nand3 i_101266416(.A(n_116782168), .B(n_126782268), .C(n_126682267
		), .Z(n_126982270));
	notech_ao4 i_102666402(.A(n_54141156), .B(n_30053), .C(n_40241017), .D(n_29095
		), .Z(n_127182272));
	notech_ao4 i_102766401(.A(n_53341148), .B(nbus_11295[9]), .C(n_53841153)
		, .D(n_30054), .Z(n_127282273));
	notech_ao4 i_102866400(.A(n_53641151), .B(n_57613), .C(n_58768), .D(n_30055
		), .Z(n_127482275));
	notech_ao4 i_102566403(.A(n_39041005), .B(n_28935), .C(n_180682807), .D(n_29062
		), .Z(n_127582276));
	notech_nand3 i_103166397(.A(n_117782178), .B(n_127582276), .C(n_127482275
		), .Z(n_127782278));
	notech_ao4 i_104566383(.A(n_54141156), .B(n_30056), .C(n_40241017), .D(n_29094
		), .Z(n_127982280));
	notech_ao4 i_104666382(.A(n_53341148), .B(nbus_11295[8]), .C(n_53841153)
		, .D(n_30057), .Z(n_128082281));
	notech_ao4 i_104766381(.A(n_53641151), .B(n_57604), .C(n_58768), .D(n_30058
		), .Z(n_128282283));
	notech_ao4 i_104466384(.A(n_39041005), .B(n_28934), .C(n_180682807), .D(n_29061
		), .Z(n_128382284));
	notech_nand3 i_105066378(.A(n_118782188), .B(n_128382284), .C(n_128282283
		), .Z(n_128582286));
	notech_ao4 i_106466364(.A(n_54141156), .B(n_30059), .C(n_40241017), .D(n_29093
		), .Z(n_128782288));
	notech_ao4 i_106566363(.A(n_53341148), .B(nbus_11295[7]), .C(n_53841153)
		, .D(n_30060), .Z(n_128882289));
	notech_ao4 i_106666362(.A(n_53641151), .B(n_57957), .C(n_58768), .D(n_30061
		), .Z(n_129082291));
	notech_ao4 i_106366365(.A(n_39041005), .B(n_28933), .C(n_180682807), .D(n_29060
		), .Z(n_129182292));
	notech_nand3 i_106966359(.A(n_119782198), .B(n_129182292), .C(n_129082291
		), .Z(n_129382294));
	notech_ao4 i_108366345(.A(n_55200), .B(n_30062), .C(n_40241017), .D(n_29092
		), .Z(n_129582296));
	notech_ao4 i_108466344(.A(n_55220), .B(n_57592), .C(n_55209), .D(n_30063
		), .Z(n_129682297));
	notech_ao4 i_108566343(.A(n_58768), .B(n_30064), .C(n_53341148), .D(nbus_11295
		[6]), .Z(n_129882299));
	notech_ao4 i_108266346(.A(n_39041005), .B(n_28932), .C(n_180682807), .D(n_29056
		), .Z(n_129982300));
	notech_nand3 i_108866340(.A(n_120782208), .B(n_129982300), .C(n_129882299
		), .Z(n_130182302));
	notech_nand2 i_155165878(.A(n_56979), .B(n_304184032), .Z(n_130382304)
		);
	notech_nand2 i_15064304(.A(n_313484125), .B(n_130782308), .Z(n_130482305
		));
	notech_nand2 i_27564186(.A(divr_1[19]), .B(n_60268), .Z(n_130582306));
	notech_nand3 i_85063625(.A(n_130882309), .B(n_60122), .C(n_60268), .Z(n_130782308
		));
	notech_or4 i_49409(.A(n_138682387), .B(n_138882389), .C(n_138782388), .D
		(n_26778), .Z(n_130882309));
	notech_or4 i_168267440(.A(n_61154), .B(n_3790), .C(n_32567), .D(n_29655)
		, .Z(n_57403));
	notech_and4 i_85463621(.A(n_59407), .B(n_59397), .C(n_246991940), .D(imm
		[31]), .Z(n_130982310));
	notech_and4 i_85663620(.A(n_59407), .B(n_59398), .C(n_246991940), .D(imm
		[30]), .Z(n_131082311));
	notech_and4 i_85763619(.A(n_59407), .B(n_59398), .C(n_246991940), .D(imm
		[26]), .Z(n_131182312));
	notech_and4 i_85863618(.A(n_59407), .B(n_59398), .C(n_246991940), .D(imm
		[25]), .Z(n_131282313));
	notech_ao4 i_10764346(.A(n_59440), .B(n_26880), .C(n_131982320), .D(n_26881
		), .Z(n_131382314));
	notech_ao4 i_14664308(.A(n_3824), .B(n_26939), .C(n_3829), .D(n_24996), 
		.Z(n_131482315));
	notech_nand3 i_7364380(.A(n_27035), .B(n_30905), .C(n_132282323), .Z(n_131982320
		));
	notech_ao4 i_6664387(.A(n_56941), .B(n_3695), .C(n_30910), .D(n_32295), 
		.Z(n_132182322));
	notech_nand2 i_92563552(.A(n_3825), .B(n_56527), .Z(n_132282323));
	notech_ao3 i_14364311(.A(n_184658942), .B(n_27034), .C(n_132782328), .Z(n_132482325
		));
	notech_and2 i_95963518(.A(n_341380914), .B(n_56485), .Z(n_132782328));
	notech_ao4 i_96063517(.A(n_59275), .B(n_59355), .C(n_26837), .D(n_26991)
		, .Z(n_132882329));
	notech_and4 i_96163516(.A(n_62868), .B(n_28122), .C(n_30931), .D(n_57602
		), .Z(n_132982330));
	notech_nao3 i_13864316(.A(n_184658942), .B(n_133382334), .C(n_3823), .Z(n_133082331
		));
	notech_nand2 i_100463475(.A(n_56566), .B(n_27033), .Z(n_133382334));
	notech_ao4 i_100663474(.A(n_246791942), .B(n_59355), .C(n_26837), .D(n_26991
		), .Z(n_133482335));
	notech_and4 i_100763473(.A(n_62868), .B(n_28122), .C(n_27301), .D(n_28120
		), .Z(n_133582336));
	notech_or4 i_17364281(.A(n_25625), .B(n_25617), .C(n_190710119), .D(\nbus_11365[25] 
		), .Z(n_134482345));
	notech_or4 i_18264272(.A(n_25625), .B(n_25617), .C(n_190710119), .D(\nbus_11365[26] 
		), .Z(n_135382354));
	notech_or4 i_19164263(.A(n_25625), .B(n_25617), .C(n_190710119), .D(n_57828
		), .Z(n_136282363));
	notech_nao3 i_20764248(.A(n_9369), .B(n_55820), .C(n_59451), .Z(n_136782368
		));
	notech_nao3 i_20464251(.A(nbus_166[31]), .B(n_55820), .C(n_27917), .Z(n_137082371
		));
	notech_ao4 i_20064254(.A(n_56204), .B(n_130982310), .C(n_179382794), .D(n_26781
		), .Z(n_137382374));
	notech_nao3 i_74863725(.A(opc[9]), .B(n_62824), .C(n_313270143), .Z(n_137682377
		));
	notech_or2 i_74763726(.A(n_60016), .B(n_57025), .Z(n_137982380));
	notech_nao3 i_74263731(.A(n_319091633), .B(n_56925), .C(n_58106), .Z(n_138482385
		));
	notech_nand2 i_19731(.A(n_61559), .B(n_130482305), .Z(n_138582386));
	notech_nor2 i_85363622(.A(n_32580), .B(n_57403), .Z(n_138682387));
	notech_and4 i_85163624(.A(n_26776), .B(n_57839), .C(n_26759), .D(n_27056
		), .Z(n_138782388));
	notech_and3 i_85263623(.A(n_19101), .B(n_32586), .C(n_5221), .Z(n_138882389
		));
	notech_or4 i_91463563(.A(n_57042), .B(n_57064), .C(n_345480955), .D(n_57011
		), .Z(n_139782398));
	notech_and4 i_90763569(.A(n_62868), .B(n_131382314), .C(n_76638786), .D(n_30930
		), .Z(n_140082401));
	notech_or4 i_90963568(.A(instrc[103]), .B(n_29635), .C(n_26899), .D(instrc
		[102]), .Z(n_140182402));
	notech_nor2 i_95663521(.A(n_56485), .B(n_3829), .Z(n_140682407));
	notech_or2 i_95163526(.A(n_58802), .B(n_132482325), .Z(n_140782408));
	notech_ao4 i_95263525(.A(n_26883), .B(n_132882329), .C(n_132982330), .D(n_26882
		), .Z(n_140882409));
	notech_or2 i_95363524(.A(n_66438684), .B(n_26968), .Z(n_140982410));
	notech_and4 i_94863529(.A(n_26858), .B(instrc[98]), .C(n_28130), .D(n_30352
		), .Z(n_141082411));
	notech_and4 i_94963528(.A(n_30350), .B(instrc[102]), .C(n_29635), .D(n_29637
		), .Z(n_141182412));
	notech_and4 i_95063527(.A(n_57011), .B(n_57064), .C(n_57033), .D(n_30342
		), .Z(n_141282413));
	notech_and4 i_100063478(.A(n_30350), .B(n_29637), .C(instrc[101]), .D(instrc
		[102]), .Z(n_141782418));
	notech_and4 i_99563483(.A(n_57064), .B(n_57078), .C(n_30946), .D(n_133082331
		), .Z(n_141882419));
	notech_ao4 i_99663482(.A(n_133482335), .B(n_26883), .C(n_133582336), .D(n_28546
		), .Z(n_141982420));
	notech_ao3 i_99763481(.A(instrc[125]), .B(instrc[126]), .C(n_66438684), 
		.Z(n_142082421));
	notech_and4 i_99363485(.A(n_29639), .B(instrc[96]), .C(n_77638796), .D(n_30332
		), .Z(n_142182422));
	notech_ao3 i_99463484(.A(instrc[121]), .B(n_27031), .C(n_32614), .Z(n_142282423
		));
	notech_and4 i_99163487(.A(n_57078), .B(n_57033), .C(n_57064), .D(n_30342
		), .Z(n_142382424));
	notech_and4 i_99263486(.A(n_30301), .B(n_30352), .C(n_30933), .D(n_28132
		), .Z(n_142482425));
	notech_or4 i_173962764(.A(n_142182422), .B(n_142482425), .C(n_142382424)
		, .D(n_142282423), .Z(n_143182432));
	notech_or4 i_174062763(.A(n_141982420), .B(n_141882419), .C(n_143182432)
		, .D(n_142082421), .Z(n_143582436));
	notech_ao4 i_173262771(.A(n_65638676), .B(n_316384154), .C(n_26889), .D(n_65738677
		), .Z(n_143682437));
	notech_ao4 i_173062773(.A(n_56566), .B(n_3829), .C(n_61117), .D(n_28532)
		, .Z(n_143882439));
	notech_nand2 i_173162772(.A(n_3821), .B(n_143882439), .Z(n_143982440));
	notech_nao3 i_168462818(.A(n_140782408), .B(n_140982410), .C(n_140882409
		), .Z(n_144982450));
	notech_or4 i_168762815(.A(n_141182412), .B(n_141082411), .C(n_141282413)
		, .D(n_144982450), .Z(n_145082451));
	notech_ao4 i_168062822(.A(n_26892), .B(n_346180962), .C(n_65738677), .D(n_30969
		), .Z(n_145182452));
	notech_ao4 i_167962823(.A(n_316384154), .B(n_190010112), .C(n_345980960)
		, .D(n_32614), .Z(n_145382454));
	notech_ao4 i_165762845(.A(n_74838768), .B(n_26888), .C(n_131482315), .D(n_32295
		), .Z(n_145882459));
	notech_ao3 i_165962843(.A(n_140182402), .B(n_145882459), .C(n_140082401)
		, .Z(n_145982460));
	notech_ao4 i_165562847(.A(n_77438794), .B(n_26887), .C(n_32343), .D(n_74738767
		), .Z(n_146082461));
	notech_ao4 i_165262850(.A(n_26959), .B(n_26886), .C(n_65638676), .D(n_344680947
		), .Z(n_146382464));
	notech_ao4 i_165162851(.A(n_74438764), .B(n_24996), .C(n_26939), .D(n_251040528
		), .Z(n_146482465));
	notech_ao4 i_164962853(.A(n_3829), .B(n_56527), .C(n_26885), .D(n_26956)
		, .Z(n_146682467));
	notech_and4 i_165462848(.A(n_344480945), .B(n_146682467), .C(n_146482465
		), .D(n_146382464), .Z(n_146882469));
	notech_ao4 i_147863016(.A(n_147271952), .B(n_27992), .C(n_58608), .D(n_54736
		), .Z(n_147482475));
	notech_ao4 i_147763017(.A(n_57181), .B(n_56136), .C(n_26607), .D(\nbus_11307[9] 
		), .Z(n_147682477));
	notech_ao4 i_147463020(.A(n_319970210), .B(n_56127), .C(n_291963186), .D
		(n_319870209), .Z(n_147882479));
	notech_and4 i_147663018(.A(n_200065529), .B(n_147882479), .C(n_137982380
		), .D(n_137682377), .Z(n_148182482));
	notech_or4 i_6964384(.A(fsm[2]), .B(n_61167), .C(n_61154), .D(n_60074), 
		.Z(n_148282483));
	notech_or2 i_25164457(.A(n_148282483), .B(\nbus_11358[31] ), .Z(n_148382484
		));
	notech_or2 i_24164458(.A(n_148282483), .B(nbus_11295[31]), .Z(n_148482485
		));
	notech_ao4 i_118263304(.A(n_55564), .B(n_30080), .C(n_55549), .D(\nbus_11365[19] 
		), .Z(n_148582486));
	notech_ao4 i_115863326(.A(n_55564), .B(opb[31]), .C(n_148382484), .D(opc
		[31]), .Z(n_148682487));
	notech_ao4 i_115663328(.A(n_55220), .B(\nbus_11365[31] ), .C(n_55229), .D
		(nbus_11295[31]), .Z(n_148882489));
	notech_and4 i_116063324(.A(n_148882489), .B(n_148682487), .C(n_137082371
		), .D(n_26901), .Z(n_149082491));
	notech_ao4 i_115363331(.A(n_55209), .B(n_30079), .C(n_58768), .D(n_30078
		), .Z(n_149182492));
	notech_ao4 i_115263332(.A(n_328184272), .B(n_29085), .C(n_52741142), .D(n_28123
		), .Z(n_149382494));
	notech_ao4 i_114963335(.A(n_55229), .B(nbus_11295[30]), .C(n_30077), .D(n_328284273
		), .Z(n_149582496));
	notech_ao4 i_114763336(.A(n_58768), .B(n_30076), .C(n_58773), .D(n_29115
		), .Z(n_149782498));
	notech_and3 i_115163333(.A(n_149582496), .B(n_149782498), .C(n_136282363
		), .Z(n_149882499));
	notech_ao4 i_114563338(.A(n_55200), .B(n_30075), .C(n_55209), .D(n_30074
		), .Z(n_149982500));
	notech_ao4 i_114463339(.A(n_328184272), .B(n_29084), .C(n_52741142), .D(n_28121
		), .Z(n_150082501));
	notech_ao4 i_114163342(.A(n_55229), .B(nbus_11295[26]), .C(n_30073), .D(n_328284273
		), .Z(n_150282503));
	notech_ao4 i_114063343(.A(n_55632), .B(n_30072), .C(n_58773), .D(n_29112
		), .Z(n_150482505));
	notech_and3 i_114363340(.A(n_150282503), .B(n_150482505), .C(n_135382354
		), .Z(n_150582506));
	notech_ao4 i_113863345(.A(n_55200), .B(n_30071), .C(n_55209), .D(n_30070
		), .Z(n_150682507));
	notech_ao4 i_113763346(.A(n_328184272), .B(n_29080), .C(n_52741142), .D(n_28115
		), .Z(n_150782508));
	notech_ao4 i_113463349(.A(n_55229), .B(nbus_11295[25]), .C(n_30068), .D(n_328284273
		), .Z(n_150982510));
	notech_ao4 i_113363350(.A(n_55632), .B(n_30067), .C(n_58773), .D(n_29111
		), .Z(n_151182512));
	notech_and3 i_113663347(.A(n_150982510), .B(n_151182512), .C(n_134482345
		), .Z(n_151282513));
	notech_ao4 i_113163352(.A(n_55200), .B(n_30066), .C(n_55209), .D(n_30065
		), .Z(n_151382514));
	notech_ao4 i_113063353(.A(n_328184272), .B(n_29079), .C(n_52741142), .D(n_28114
		), .Z(n_151482515));
	notech_or2 i_97460787(.A(n_56356), .B(nbus_11295[30]), .Z(n_151682517)
		);
	notech_nao3 i_97360788(.A(n_62822), .B(opc_10[30]), .C(n_306124325), .Z(n_151982520
		));
	notech_or4 i_96860793(.A(n_58132), .B(n_58493), .C(n_56903), .D(n_55929)
		, .Z(n_152482525));
	notech_ao3 i_107460704(.A(n_62798), .B(opc_10[30]), .C(n_306624330), .Z(n_152582526
		));
	notech_or4 i_106960709(.A(n_54756), .B(n_58494), .C(n_56432), .D(n_55929
		), .Z(n_153282533));
	notech_nao3 i_112760656(.A(n_62776), .B(opc_10[30]), .C(n_286827250), .Z
		(n_153382534));
	notech_or4 i_112260661(.A(n_54709), .B(n_58495), .C(n_56443), .D(n_55929
		), .Z(n_154082541));
	notech_ao4 i_219059648(.A(n_58139), .B(n_302991794), .C(n_57861), .D(n_57828
		), .Z(n_154182542));
	notech_ao4 i_218959649(.A(n_287827260), .B(n_303091793), .C(n_26615), .D
		(n_29591), .Z(n_154382544));
	notech_ao4 i_218759651(.A(n_286927251), .B(n_32252), .C(n_58424), .D(n_28015
		), .Z(n_154582546));
	notech_and3 i_218859650(.A(n_153382534), .B(n_154582546), .C(n_26604), .Z
		(n_154782548));
	notech_ao4 i_214759691(.A(n_58141), .B(n_302991794), .C(n_314047718), .D
		(n_57828), .Z(n_154882549));
	notech_ao4 i_214659692(.A(n_306824332), .B(n_303091793), .C(n_307324337)
		, .D(n_29591), .Z(n_155082551));
	notech_nand3 i_214959689(.A(n_154882549), .B(n_155082551), .C(n_153282533
		), .Z(n_155182552));
	notech_ao4 i_214459694(.A(n_307124335), .B(n_32252), .C(n_58425), .D(n_28015
		), .Z(n_155282553));
	notech_ao4 i_207359765(.A(n_302991794), .B(n_58143), .C(n_57870), .D(n_57828
		), .Z(n_155582556));
	notech_ao4 i_207259766(.A(n_303091793), .B(n_305924323), .C(n_29591), .D
		(n_26902), .Z(n_155782558));
	notech_ao4 i_206959769(.A(n_32252), .B(n_58085), .C(n_58427), .D(n_28015
		), .Z(n_155982560));
	notech_and4 i_207159767(.A(n_155982560), .B(n_151682517), .C(n_151982520
		), .D(n_26604), .Z(n_156282563));
	notech_and2 i_14958344(.A(n_58646), .B(n_156682567), .Z(n_156382564));
	notech_and2 i_15058343(.A(n_158082581), .B(n_58610), .Z(n_156482565));
	notech_nand3 i_15158342(.A(n_181779321), .B(n_57873), .C(n_157682577), .Z
		(n_156582566));
	notech_nao3 i_79657721(.A(n_56423), .B(opa[0]), .C(n_58133), .Z(n_156682567
		));
	notech_or4 i_79557722(.A(n_54814), .B(n_26906), .C(nbus_11295[0]), .D(n_60933
		), .Z(n_156782568));
	notech_or4 i_79457723(.A(n_58489), .B(n_54814), .C(n_28124), .D(n_60933)
		, .Z(n_157082571));
	notech_nand2 i_78957728(.A(opb[0]), .B(n_156582566), .Z(n_157582576));
	notech_or4 i_79957718(.A(n_60854), .B(n_58133), .C(n_58505), .D(n_26735)
		, .Z(n_157682577));
	notech_ao4 i_167656872(.A(n_56046), .B(n_58325), .C(n_56037), .D(n_295921141
		), .Z(n_158082581));
	notech_ao4 i_167256876(.A(n_58489), .B(n_156482565), .C(n_26906), .D(n_156382564
		), .Z(n_158182582));
	notech_ao4 i_167156877(.A(n_303973519), .B(n_59187), .C(n_175062033), .D
		(n_303873518), .Z(n_158382584));
	notech_ao4 i_166856880(.A(n_291363180), .B(n_304073520), .C(n_304273522)
		, .D(n_59993), .Z(n_158582586));
	notech_and4 i_167056878(.A(n_152275466), .B(n_156782568), .C(n_157082571
		), .D(n_158582586), .Z(n_158882589));
	notech_or2 i_18455336(.A(n_58750), .B(n_27997), .Z(n_159182592));
	notech_or4 i_18155339(.A(n_25617), .B(n_27573), .C(n_303747815), .D(nbus_11295
		[12]), .Z(n_159482595));
	notech_nao3 i_17855342(.A(n_11280), .B(n_60292), .C(n_1893), .Z(n_159782598
		));
	notech_or2 i_17555345(.A(n_58788), .B(n_28399), .Z(n_160082601));
	notech_or2 i_19955324(.A(n_58750), .B(n_27998), .Z(n_160382604));
	notech_or4 i_19655327(.A(n_25617), .B(n_303747815), .C(n_27573), .D(nbus_11295
		[13]), .Z(n_160682607));
	notech_nao3 i_19255330(.A(n_11282), .B(n_60292), .C(n_1893), .Z(n_160982610
		));
	notech_or2 i_18755333(.A(n_58788), .B(n_28400), .Z(n_161282613));
	notech_or2 i_21155312(.A(n_58750), .B(n_27999), .Z(n_161582616));
	notech_or4 i_20855315(.A(n_25617), .B(n_27573), .C(n_303747815), .D(nbus_11295
		[14]), .Z(n_161882619));
	notech_nao3 i_20555318(.A(n_11284), .B(n_60292), .C(n_1893), .Z(n_162182622
		));
	notech_or2 i_20255321(.A(n_58788), .B(n_28401), .Z(n_162482625));
	notech_or2 i_22355300(.A(n_58750), .B(n_28000), .Z(n_162782628));
	notech_or4 i_22055303(.A(n_25617), .B(n_27573), .C(n_303747815), .D(nbus_11295
		[15]), .Z(n_163082631));
	notech_nao3 i_21755306(.A(n_11286), .B(n_60292), .C(n_1893), .Z(n_163382634
		));
	notech_or2 i_21455309(.A(n_58788), .B(n_28402), .Z(n_163682637));
	notech_or2 i_23655288(.A(n_58750), .B(n_28001), .Z(n_163982640));
	notech_or4 i_23255291(.A(n_25617), .B(n_27573), .C(n_303747815), .D(nbus_11295
		[16]), .Z(n_164282643));
	notech_nao3 i_22955294(.A(n_11288), .B(n_60292), .C(n_1893), .Z(n_164582646
		));
	notech_or2 i_22655297(.A(n_58788), .B(n_28403), .Z(n_164882649));
	notech_or2 i_24855276(.A(n_58750), .B(n_28002), .Z(n_165182652));
	notech_or4 i_24555279(.A(n_25617), .B(n_27573), .C(n_303747815), .D(nbus_11295
		[17]), .Z(n_165482655));
	notech_nao3 i_24255282(.A(n_11290), .B(n_60292), .C(n_1893), .Z(n_165782658
		));
	notech_or2 i_23955285(.A(n_58788), .B(n_28404), .Z(n_166082661));
	notech_or2 i_26055264(.A(n_58750), .B(n_28003), .Z(n_166382664));
	notech_or4 i_25755267(.A(n_25617), .B(n_27573), .C(n_303747815), .D(nbus_11295
		[18]), .Z(n_166682667));
	notech_nao3 i_25455270(.A(n_11292), .B(n_60303), .C(n_1893), .Z(n_166982670
		));
	notech_or2 i_25155273(.A(n_58788), .B(n_28405), .Z(n_167282673));
	notech_or2 i_27255252(.A(n_58750), .B(n_28004), .Z(n_167582676));
	notech_or4 i_26955255(.A(n_25617), .B(n_27573), .C(n_303747815), .D(nbus_11295
		[19]), .Z(n_167882679));
	notech_nao3 i_26655258(.A(n_11294), .B(n_60294), .C(n_1893), .Z(n_168182682
		));
	notech_or2 i_26355261(.A(n_58788), .B(n_28406), .Z(n_168482685));
	notech_or2 i_28455240(.A(n_58750), .B(n_28013), .Z(n_168782688));
	notech_or4 i_28155243(.A(n_25617), .B(n_27573), .C(n_303747815), .D(nbus_11295
		[28]), .Z(n_169082691));
	notech_nao3 i_27855246(.A(n_11312), .B(n_60294), .C(n_1893), .Z(n_169382694
		));
	notech_or2 i_27555249(.A(n_58788), .B(n_28415), .Z(n_169682697));
	notech_ao4 i_64154915(.A(n_58789), .B(n_28621), .C(n_58791), .D(n_29374)
		, .Z(n_169782698));
	notech_ao4 i_63954917(.A(n_27065), .B(n_29343), .C(n_59153), .D(n_29312)
		, .Z(n_169982700));
	notech_and4 i_64354913(.A(n_169982700), .B(n_169782698), .C(n_169382694)
		, .D(n_169682697), .Z(n_170182702));
	notech_ao4 i_63654920(.A(n_310247754), .B(n_30099), .C(n_330563522), .D(n_27831
		), .Z(n_170282703));
	notech_ao4 i_63454922(.A(n_58751), .B(\nbus_11358[28] ), .C(n_310447752)
		, .D(n_30098), .Z(n_170482705));
	notech_and4 i_63854918(.A(n_170482705), .B(n_170282703), .C(n_168782688)
		, .D(n_169082691), .Z(n_170682707));
	notech_ao4 i_63154925(.A(n_58789), .B(n_28612), .C(n_58791), .D(n_29365)
		, .Z(n_170782708));
	notech_ao4 i_62954927(.A(n_27065), .B(n_29334), .C(n_59152), .D(n_29303)
		, .Z(n_170982710));
	notech_and4 i_63354923(.A(n_170982710), .B(n_170782708), .C(n_168182682)
		, .D(n_168482685), .Z(n_171182712));
	notech_ao4 i_62654930(.A(n_310247754), .B(n_30097), .C(n_330563522), .D(n_27822
		), .Z(n_171282713));
	notech_ao4 i_62454932(.A(n_58751), .B(n_56311), .C(n_310447752), .D(n_30096
		), .Z(n_171482715));
	notech_and4 i_62854928(.A(n_171482715), .B(n_171282713), .C(n_167582676)
		, .D(n_167882679), .Z(n_171682717));
	notech_ao4 i_62154935(.A(n_58789), .B(n_28611), .C(n_58791), .D(n_29364)
		, .Z(n_171782718));
	notech_ao4 i_61954937(.A(n_27065), .B(n_29333), .C(n_59152), .D(n_29302)
		, .Z(n_171982720));
	notech_and4 i_62354933(.A(n_171982720), .B(n_171782718), .C(n_166982670)
		, .D(n_167282673), .Z(n_172182722));
	notech_ao4 i_61654940(.A(n_310247754), .B(n_30095), .C(n_330563522), .D(n_27821
		), .Z(n_172282723));
	notech_ao4 i_61454942(.A(n_58751), .B(n_56302), .C(n_310447752), .D(n_30094
		), .Z(n_172482725));
	notech_and4 i_61854938(.A(n_172482725), .B(n_172282723), .C(n_166382664)
		, .D(n_166682667), .Z(n_172682727));
	notech_ao4 i_61154945(.A(n_58789), .B(n_28610), .C(n_58791), .D(n_29363)
		, .Z(n_172782728));
	notech_ao4 i_60954947(.A(n_27065), .B(n_29332), .C(n_59152), .D(n_29301)
		, .Z(n_172982730));
	notech_and4 i_61354943(.A(n_172982730), .B(n_172782728), .C(n_165782658)
		, .D(n_166082661), .Z(n_173182732));
	notech_ao4 i_60654950(.A(n_310247754), .B(n_30093), .C(n_330563522), .D(n_27820
		), .Z(n_173282733));
	notech_ao4 i_60354952(.A(n_58751), .B(n_56293), .C(n_310447752), .D(n_30092
		), .Z(n_173482735));
	notech_and4 i_60854948(.A(n_173482735), .B(n_173282733), .C(n_165182652)
		, .D(n_165482655), .Z(n_173682737));
	notech_ao4 i_59954955(.A(n_58789), .B(n_28609), .C(n_58791), .D(n_29362)
		, .Z(n_173782738));
	notech_ao4 i_59654957(.A(n_27065), .B(n_29331), .C(n_59152), .D(n_29300)
		, .Z(n_173982740));
	notech_and4 i_60154953(.A(n_173982740), .B(n_173782738), .C(n_164582646)
		, .D(n_164882649), .Z(n_174182742));
	notech_ao4 i_59354960(.A(n_310247754), .B(n_30091), .C(n_330563522), .D(n_27819
		), .Z(n_174282743));
	notech_ao4 i_59154962(.A(n_58751), .B(n_56284), .C(n_310447752), .D(n_30090
		), .Z(n_174482745));
	notech_and4 i_59554958(.A(n_174482745), .B(n_174282743), .C(n_163982640)
		, .D(n_164282643), .Z(n_174682747));
	notech_ao4 i_58754965(.A(n_58789), .B(n_28608), .C(n_58791), .D(n_29361)
		, .Z(n_174782748));
	notech_ao4 i_58354967(.A(n_27065), .B(n_29330), .C(n_59152), .D(n_29299)
		, .Z(n_174982750));
	notech_and4 i_59054963(.A(n_174982750), .B(n_174782748), .C(n_163382634)
		, .D(n_163682637), .Z(n_175182752));
	notech_ao4 i_58054970(.A(n_310247754), .B(n_30089), .C(n_330563522), .D(n_27818
		), .Z(n_175282753));
	notech_ao4 i_57854972(.A(n_58751), .B(n_56275), .C(n_310447752), .D(n_30087
		), .Z(n_175482755));
	notech_and4 i_58254968(.A(n_175482755), .B(n_175282753), .C(n_162782628)
		, .D(n_163082631), .Z(n_175682757));
	notech_ao4 i_57554975(.A(n_58789), .B(n_28607), .C(n_58791), .D(n_29360)
		, .Z(n_175782758));
	notech_ao4 i_57354977(.A(n_27065), .B(n_29329), .C(n_59152), .D(n_29298)
		, .Z(n_175982760));
	notech_and4 i_57754973(.A(n_175982760), .B(n_175782758), .C(n_162182622)
		, .D(n_162482625), .Z(n_176182762));
	notech_ao4 i_57054980(.A(n_310247754), .B(n_30086), .C(n_330563522), .D(n_27817
		), .Z(n_176282763));
	notech_ao4 i_56854982(.A(n_58751), .B(n_56248), .C(n_310447752), .D(n_30085
		), .Z(n_176482765));
	notech_and4 i_57254978(.A(n_176482765), .B(n_176282763), .C(n_161582616)
		, .D(n_161882619), .Z(n_176682767));
	notech_ao4 i_56454985(.A(n_58789), .B(n_28606), .C(n_58791), .D(n_29359)
		, .Z(n_176782768));
	notech_ao4 i_56254987(.A(n_27065), .B(n_29328), .C(n_59152), .D(n_29297)
		, .Z(n_176982770));
	notech_and4 i_56654983(.A(n_176982770), .B(n_176782768), .C(n_160982610)
		, .D(n_161282613), .Z(n_177182772));
	notech_ao4 i_55954990(.A(n_310247754), .B(n_30084), .C(n_330563522), .D(n_27816
		), .Z(n_177282773));
	notech_ao4 i_55754992(.A(n_58751), .B(\nbus_11358[13] ), .C(n_310447752)
		, .D(n_30083), .Z(n_177482775));
	notech_and4 i_56154988(.A(n_177482775), .B(n_177282773), .C(n_160382604)
		, .D(n_160682607), .Z(n_177682777));
	notech_ao4 i_55454995(.A(n_58789), .B(n_28605), .C(n_58791), .D(n_29358)
		, .Z(n_177782778));
	notech_ao4 i_55254997(.A(n_27065), .B(n_29327), .C(n_59152), .D(n_29296)
		, .Z(n_177982780));
	notech_and4 i_55654993(.A(n_177982780), .B(n_177782778), .C(n_159782598)
		, .D(n_160082601), .Z(n_178182782));
	notech_ao4 i_54855000(.A(n_310247754), .B(n_30082), .C(n_330563522), .D(n_27815
		), .Z(n_178282783));
	notech_ao4 i_54655002(.A(n_58751), .B(n_56221), .C(n_310447752), .D(n_30081
		), .Z(n_178482785));
	notech_and4 i_55154998(.A(n_178482785), .B(n_178282783), .C(n_159182592)
		, .D(n_159482595), .Z(n_178682787));
	notech_nand3 i_5953853(.A(n_60113), .B(n_60294), .C(n_178982790), .Z(n_178882789
		));
	notech_nand3 i_1653893(.A(n_3986), .B(n_205183042), .C(n_212969141), .Z(n_178982790
		));
	notech_nand3 i_47592(.A(n_328484275), .B(n_205383044), .C(n_178882789), 
		.Z(n_12057));
	notech_and3 i_16953766(.A(n_318891635), .B(n_318791636), .C(imm[7]), .Z(n_179182792
		));
	notech_and4 i_17153764(.A(n_59408), .B(n_59398), .C(n_246991940), .D(imm
		[10]), .Z(n_179282793));
	notech_and3 i_17353762(.A(n_60268), .B(n_26999), .C(n_26985), .Z(n_179382794
		));
	notech_and4 i_17853757(.A(n_59408), .B(n_59398), .C(n_59286), .D(imm[27]
		), .Z(n_179582796));
	notech_or2 i_177652201(.A(n_328184272), .B(n_29081), .Z(n_179682797));
	notech_nao3 i_177252205(.A(nbus_166[27]), .B(n_55820), .C(n_59460), .Z(n_180382804
		));
	notech_ao4 i_177752200(.A(n_56204), .B(n_179582796), .C(n_179382794), .D
		(n_55191), .Z(n_180482805));
	notech_nao3 i_2812945(.A(n_206483055), .B(n_179682797), .C(n_180482805),
		 .Z(n_26083));
	notech_and2 i_180252175(.A(add_src[10]), .B(n_26910), .Z(n_180582806));
	notech_ao4 i_89253969(.A(n_26985), .B(n_60294), .C(n_180782808), .D(n_56566
		), .Z(n_180682807));
	notech_or2 i_21653968(.A(n_179282793), .B(n_56205), .Z(\nbus_11317[10] )
		);
	notech_nor2 i_24653967(.A(n_330363520), .B(n_55191), .Z(n_180782808));
	notech_ao3 i_180752170(.A(n_9264), .B(n_55820), .C(n_59451), .Z(n_181082811
		));
	notech_ao3 i_180152176(.A(n_9265), .B(n_27855), .C(n_319691627), .Z(n_181382814
		));
	notech_ao4 i_180352174(.A(n_55191), .B(n_330363520), .C(n_56205), .D(n_179282793
		), .Z(n_181682817));
	notech_or4 i_1112928(.A(n_181682817), .B(n_180582806), .C(n_207183062), 
		.D(n_26912), .Z(n_25998));
	notech_nand3 i_3218997(.A(n_207583066), .B(n_207483065), .C(n_208383074)
		, .Z(n_25674));
	notech_nand3 i_3118996(.A(n_208583076), .B(n_208483075), .C(n_209383084)
		, .Z(n_25668));
	notech_nand3 i_2718992(.A(n_209583086), .B(n_209483085), .C(n_210383094)
		, .Z(n_25644));
	notech_nand3 i_2618991(.A(n_210583096), .B(n_210483095), .C(n_211383104)
		, .Z(n_25638));
	notech_nand3 i_2518990(.A(n_211583106), .B(n_211483105), .C(n_212383114)
		, .Z(n_25632));
	notech_nand3 i_2418989(.A(n_212583116), .B(n_212483115), .C(n_213383124)
		, .Z(n_25626));
	notech_nand3 i_2318988(.A(n_213583126), .B(n_213483125), .C(n_214383134)
		, .Z(n_25620));
	notech_nand3 i_2218987(.A(n_214583136), .B(n_214483135), .C(n_215383144)
		, .Z(n_25614));
	notech_nand3 i_2118986(.A(n_215583146), .B(n_215483145), .C(n_216383154)
		, .Z(n_25608));
	notech_nand3 i_1118976(.A(n_216583156), .B(n_216483155), .C(n_217383164)
		, .Z(n_25548));
	notech_or4 i_210951872(.A(n_27988), .B(n_59435), .C(n_60268), .D(n_27990
		), .Z(n_195982950));
	notech_and4 i_1018975(.A(n_195982950), .B(n_217583166), .C(n_217483165),
		 .D(n_218483175), .Z(n_25542));
	notech_or4 i_213451847(.A(n_27988), .B(n_59435), .C(n_60268), .D(n_27989
		), .Z(n_197282963));
	notech_and4 i_918974(.A(n_197282963), .B(n_218683177), .C(n_218583176), 
		.D(n_219583186), .Z(n_25536));
	notech_or4 i_216051822(.A(n_59435), .B(n_27988), .C(n_60268), .D(n_59205
		), .Z(n_198582976));
	notech_and4 i_818973(.A(n_198582976), .B(n_219783188), .C(n_219683187), 
		.D(n_220683197), .Z(n_25530));
	notech_or4 i_218651797(.A(n_27988), .B(n_59435), .C(n_60268), .D(n_27986
		), .Z(n_199882989));
	notech_and4 i_718972(.A(n_199882989), .B(n_220883199), .C(n_220783198), 
		.D(n_221783208), .Z(n_25524));
	notech_or4 i_221151772(.A(n_27988), .B(n_59434), .C(n_60263), .D(n_27985
		), .Z(n_201183002));
	notech_and4 i_618971(.A(n_201183002), .B(n_221983210), .C(n_221883209), 
		.D(n_222883219), .Z(n_25518));
	notech_or4 i_223651747(.A(n_59429), .B(n_27988), .C(n_60268), .D(n_59259
		), .Z(n_202483015));
	notech_and4 i_518970(.A(n_202483015), .B(n_223083221), .C(n_222983220), 
		.D(n_223983230), .Z(n_25512));
	notech_or4 i_226151722(.A(n_27988), .B(n_59429), .C(n_60268), .D(n_27983
		), .Z(n_203783028));
	notech_and4 i_418969(.A(n_203783028), .B(n_224183232), .C(n_224083231), 
		.D(n_225083241), .Z(n_25506));
	notech_or4 i_228651697(.A(n_27988), .B(n_59424), .C(n_60268), .D(n_59187
		), .Z(n_205083041));
	notech_and4 i_318968(.A(n_205083041), .B(n_225283243), .C(n_225183242), 
		.D(n_226183252), .Z(n_25500));
	notech_ao4 i_5853854(.A(n_59460), .B(n_303991784), .C(n_2895), .D(1'b0),
		 .Z(n_205183042));
	notech_and3 i_6153851(.A(n_3820), .B(n_248240500), .C(n_326184252), .Z(n_205383044
		));
	notech_or4 i_101753913(.A(n_32304), .B(n_26783), .C(n_179182792), .D(n_329763514
		), .Z(n_81541430));
	notech_nand3 i_29653923(.A(n_19050), .B(n_60268), .C(n_26985), .Z(n_52741142
		));
	notech_or4 i_37775(.A(n_2885), .B(n_61156), .C(n_3790), .D(n_19079), .Z(n_205883049
		));
	notech_ao4 i_178052197(.A(n_55200), .B(n_30102), .C(n_55632), .D(n_30101
		), .Z(n_205983050));
	notech_ao4 i_178152196(.A(n_55220), .B(n_57792), .C(n_55229), .D(n_57881
		), .Z(n_206183052));
	notech_ao4 i_178252195(.A(n_52741142), .B(n_28116), .C(n_55209), .D(n_30103
		), .Z(n_206283053));
	notech_and4 i_178552192(.A(n_206283053), .B(n_206183052), .C(n_205983050
		), .D(n_180382804), .Z(n_206483055));
	notech_ao4 i_181252165(.A(n_40241017), .B(n_29096), .C(n_39041005), .D(n_28936
		), .Z(n_206683057));
	notech_ao4 i_181052167(.A(n_55220), .B(n_57625), .C(n_55229), .D(nbus_11295
		[10]), .Z(n_206783058));
	notech_ao4 i_180852169(.A(n_28099), .B(n_205883049), .C(n_55632), .D(n_30104
		), .Z(n_206883059));
	notech_or4 i_181452164(.A(n_181082811), .B(n_181382814), .C(n_26915), .D
		(n_26913), .Z(n_207183062));
	notech_ao4 i_183452144(.A(n_58788), .B(n_28418), .C(n_59152), .D(n_29315
		), .Z(n_207483065));
	notech_ao4 i_183552143(.A(n_58791), .B(n_29377), .C(n_58789), .D(n_28624
		), .Z(n_207583066));
	notech_ao4 i_183052148(.A(n_58751), .B(\nbus_11358[31] ), .C(n_58750), .D
		(n_28016), .Z(n_207783068));
	notech_ao4 i_183152147(.A(n_310347753), .B(nbus_11295[31]), .C(n_310447752
		), .D(n_30105), .Z(n_207883069));
	notech_ao4 i_183252146(.A(n_330563522), .B(n_27834), .C(n_30106), .D(n_310247754
		), .Z(n_208083071));
	notech_ao4 i_183352145(.A(n_27065), .B(n_29346), .C(n_1887), .D(n_30107)
		, .Z(n_208183072));
	notech_and4 i_183952139(.A(n_208183072), .B(n_208083071), .C(n_207883069
		), .D(n_207783068), .Z(n_208383074));
	notech_ao4 i_185752121(.A(n_58788), .B(n_28417), .C(n_59152), .D(n_29314
		), .Z(n_208483075));
	notech_ao4 i_185852120(.A(n_58791), .B(n_29376), .C(n_58789), .D(n_28623
		), .Z(n_208583076));
	notech_ao4 i_185352125(.A(n_58751), .B(n_55929), .C(n_58750), .D(n_28015
		), .Z(n_208783078));
	notech_ao4 i_185452124(.A(n_310347753), .B(nbus_11295[30]), .C(n_310447752
		), .D(n_30108), .Z(n_208883079));
	notech_ao4 i_185552123(.A(n_330563522), .B(n_27833), .C(n_310247754), .D
		(n_30110), .Z(n_209083081));
	notech_ao4 i_185652122(.A(n_27065), .B(n_29345), .C(n_1887), .D(n_30111)
		, .Z(n_209183082));
	notech_and4 i_186252116(.A(n_209183082), .B(n_209083081), .C(n_208883079
		), .D(n_208783078), .Z(n_209383084));
	notech_ao4 i_192652052(.A(n_58751), .B(\nbus_11358[26] ), .C(n_310347753
		), .D(nbus_11295[26]), .Z(n_209483085));
	notech_ao4 i_192752051(.A(n_58788), .B(n_28413), .C(n_58750), .D(n_28011
		), .Z(n_209583086));
	notech_ao4 i_192252056(.A(n_310247754), .B(n_30113), .C(n_310447752), .D
		(n_30112), .Z(n_209783088));
	notech_ao4 i_192352055(.A(n_1887), .B(n_30114), .C(n_330563522), .D(n_27829
		), .Z(n_209883089));
	notech_ao4 i_192452054(.A(n_59152), .B(n_29310), .C(n_27065), .D(n_29341
		), .Z(n_210083091));
	notech_ao4 i_192552053(.A(n_58789), .B(n_28619), .C(n_58791), .D(n_29372
		), .Z(n_210183092));
	notech_and4 i_193152047(.A(n_210183092), .B(n_210083091), .C(n_209883089
		), .D(n_209783088), .Z(n_210383094));
	notech_ao4 i_194952029(.A(n_58788), .B(n_28412), .C(n_59153), .D(n_29309
		), .Z(n_210483095));
	notech_ao4 i_195052028(.A(n_58791), .B(n_29371), .C(n_58789), .D(n_28618
		), .Z(n_210583096));
	notech_ao4 i_194552033(.A(n_58751), .B(n_55965), .C(n_58750), .D(n_28010
		), .Z(n_210783098));
	notech_ao4 i_194652032(.A(n_310347753), .B(nbus_11295[25]), .C(n_310447752
		), .D(n_30115), .Z(n_210883099));
	notech_ao4 i_194752031(.A(n_330563522), .B(n_27828), .C(n_310247754), .D
		(n_30116), .Z(n_211083101));
	notech_ao4 i_194852030(.A(n_27065), .B(n_29340), .C(n_1887), .D(n_30117)
		, .Z(n_211183102));
	notech_and4 i_195452024(.A(n_211183102), .B(n_211083101), .C(n_210883099
		), .D(n_210783098), .Z(n_211383104));
	notech_ao4 i_197252006(.A(n_58788), .B(n_28411), .C(n_59153), .D(n_29308
		), .Z(n_211483105));
	notech_ao4 i_197352005(.A(n_58791), .B(n_29370), .C(n_58789), .D(n_28617
		), .Z(n_211583106));
	notech_ao4 i_196852010(.A(n_58751), .B(n_56475), .C(n_58750), .D(n_28009
		), .Z(n_211783108));
	notech_ao4 i_196952009(.A(n_310347753), .B(nbus_11295[24]), .C(n_310447752
		), .D(n_30118), .Z(n_211883109));
	notech_ao4 i_197052008(.A(n_330563522), .B(n_27827), .C(n_310247754), .D
		(n_30119), .Z(n_212083111));
	notech_ao4 i_197152007(.A(n_27065), .B(n_29339), .C(n_1887), .D(n_30120)
		, .Z(n_212183112));
	notech_and4 i_197752001(.A(n_212183112), .B(n_212083111), .C(n_211883109
		), .D(n_211783108), .Z(n_212383114));
	notech_ao4 i_199551983(.A(n_58788), .B(n_28410), .C(n_59153), .D(n_29307
		), .Z(n_212483115));
	notech_ao4 i_199651982(.A(n_58791), .B(n_29369), .C(n_58789), .D(n_28616
		), .Z(n_212583116));
	notech_ao4 i_199151987(.A(n_55429), .B(n_56347), .C(n_55400), .D(n_28008
		), .Z(n_212783118));
	notech_ao4 i_199251986(.A(n_310347753), .B(nbus_11295[23]), .C(n_55420),
		 .D(n_30121), .Z(n_212883119));
	notech_ao4 i_199351985(.A(n_59176), .B(n_27826), .C(n_310247754), .D(n_30122
		), .Z(n_213083121));
	notech_ao4 i_199451984(.A(n_59335), .B(n_29338), .C(n_1887), .D(n_30125)
		, .Z(n_213183122));
	notech_and4 i_200051978(.A(n_213183122), .B(n_213083121), .C(n_212883119
		), .D(n_212783118), .Z(n_213383124));
	notech_ao4 i_201851960(.A(n_55367), .B(n_28409), .C(n_59153), .D(n_29306
		), .Z(n_213483125));
	notech_ao4 i_201951959(.A(n_55378), .B(n_29368), .C(n_55389), .D(n_28615
		), .Z(n_213583126));
	notech_ao4 i_201451964(.A(n_55429), .B(n_56338), .C(n_55400), .D(n_28007
		), .Z(n_213783128));
	notech_ao4 i_201551963(.A(n_310347753), .B(nbus_11295[22]), .C(n_55420),
		 .D(n_30127), .Z(n_213883129));
	notech_ao4 i_201651962(.A(n_59176), .B(n_27825), .C(n_55409), .D(n_30128
		), .Z(n_214083131));
	notech_ao4 i_201751961(.A(n_59335), .B(n_29337), .C(n_1887), .D(n_30129)
		, .Z(n_214183132));
	notech_and4 i_202451955(.A(n_214183132), .B(n_214083131), .C(n_213883129
		), .D(n_213783128), .Z(n_214383134));
	notech_ao4 i_204251937(.A(n_55367), .B(n_28408), .C(n_59153), .D(n_29305
		), .Z(n_214483135));
	notech_ao4 i_204351936(.A(n_55378), .B(n_29367), .C(n_55389), .D(n_28614
		), .Z(n_214583136));
	notech_ao4 i_203851941(.A(n_55429), .B(n_56329), .C(n_55400), .D(n_28006
		), .Z(n_214783138));
	notech_ao4 i_203951940(.A(n_310347753), .B(nbus_11295[21]), .C(n_55420),
		 .D(n_30130), .Z(n_214883139));
	notech_ao4 i_204051939(.A(n_59176), .B(n_27824), .C(n_55409), .D(n_30131
		), .Z(n_215083141));
	notech_ao4 i_204151938(.A(n_59335), .B(n_29336), .C(n_1887), .D(n_30132)
		, .Z(n_215183142));
	notech_and4 i_204851932(.A(n_215183142), .B(n_215083141), .C(n_214883139
		), .D(n_214783138), .Z(n_215383144));
	notech_ao4 i_206751914(.A(n_55367), .B(n_28407), .C(n_59153), .D(n_29304
		), .Z(n_215483145));
	notech_ao4 i_206851913(.A(n_55378), .B(n_29366), .C(n_55389), .D(n_28613
		), .Z(n_215583146));
	notech_ao4 i_206351918(.A(n_55429), .B(n_56320), .C(n_55400), .D(n_28005
		), .Z(n_215783148));
	notech_ao4 i_206451917(.A(n_310347753), .B(nbus_11295[20]), .C(n_55420),
		 .D(n_30133), .Z(n_215883149));
	notech_ao4 i_206551916(.A(n_59176), .B(n_27823), .C(n_55409), .D(n_30136
		), .Z(n_216083151));
	notech_ao4 i_206651915(.A(n_59335), .B(n_29335), .C(n_1887), .D(n_30137)
		, .Z(n_216183152));
	notech_and4 i_207251909(.A(n_216183152), .B(n_216083151), .C(n_215883149
		), .D(n_215783148), .Z(n_216383154));
	notech_ao4 i_209051891(.A(n_55389), .B(n_28603), .C(n_55367), .D(n_28397
		), .Z(n_216483155));
	notech_ao4 i_209151890(.A(n_310347753), .B(nbus_11295[10]), .C(n_55378),
		 .D(n_29356), .Z(n_216583156));
	notech_ao4 i_208651895(.A(n_55429), .B(n_56154), .C(n_55400), .D(n_27993
		), .Z(n_216783158));
	notech_ao4 i_208751894(.A(n_55409), .B(n_30140), .C(n_55420), .D(n_30139
		), .Z(n_216883159));
	notech_ao4 i_208851893(.A(n_1887), .B(n_30144), .C(n_59176), .D(n_27813)
		, .Z(n_217083161));
	notech_ao4 i_208951892(.A(n_59153), .B(n_29294), .C(n_59335), .D(n_29326
		), .Z(n_217183162));
	notech_and4 i_209551886(.A(n_217183162), .B(n_217083161), .C(n_216883159
		), .D(n_216783158), .Z(n_217383164));
	notech_ao4 i_211551866(.A(n_55378), .B(n_29355), .C(n_55389), .D(n_28602
		), .Z(n_217483165));
	notech_ao4 i_211051871(.A(n_55429), .B(n_56136), .C(n_55400), .D(n_27992
		), .Z(n_217583166));
	notech_ao4 i_211151870(.A(n_55347), .B(nbus_11295[9]), .C(n_55420), .D(n_30145
		), .Z(n_217883169));
	notech_ao4 i_211251869(.A(n_59176), .B(n_27812), .C(n_55409), .D(n_30146
		), .Z(n_217983170));
	notech_ao4 i_211351868(.A(n_59335), .B(n_29325), .C(n_59167), .D(n_30147
		), .Z(n_218183172));
	notech_ao4 i_211451867(.A(n_55367), .B(n_28396), .C(n_59153), .D(n_29293
		), .Z(n_218283173));
	notech_and4 i_212051861(.A(n_218283173), .B(n_218183172), .C(n_217983170
		), .D(n_217883169), .Z(n_218483175));
	notech_ao4 i_214051841(.A(n_55378), .B(n_29354), .C(n_55389), .D(n_28601
		), .Z(n_218583176));
	notech_ao4 i_213551846(.A(n_55429), .B(n_56118), .C(n_55400), .D(n_27991
		), .Z(n_218683177));
	notech_ao4 i_213651845(.A(n_55347), .B(nbus_11295[8]), .C(n_55420), .D(n_30148
		), .Z(n_218983180));
	notech_ao4 i_213751844(.A(n_59176), .B(n_27811), .C(n_55409), .D(n_30149
		), .Z(n_219083181));
	notech_ao4 i_213851843(.A(n_59335), .B(n_29324), .C(n_59167), .D(n_30150
		), .Z(n_219283183));
	notech_ao4 i_213951842(.A(n_55367), .B(n_28395), .C(n_59153), .D(n_29292
		), .Z(n_219383184));
	notech_and4 i_214551836(.A(n_219383184), .B(n_219283183), .C(n_219083181
		), .D(n_218983180), .Z(n_219583186));
	notech_ao4 i_216751816(.A(n_55378), .B(n_29353), .C(n_55389), .D(n_28600
		), .Z(n_219683187));
	notech_ao4 i_216151821(.A(n_55429), .B(n_56109), .C(n_55400), .D(n_56100
		), .Z(n_219783188));
	notech_ao4 i_216251820(.A(n_55347), .B(nbus_11295[7]), .C(n_55420), .D(n_30151
		), .Z(n_220083191));
	notech_ao4 i_216451819(.A(n_59176), .B(n_27810), .C(n_55409), .D(n_30152
		), .Z(n_220183192));
	notech_ao4 i_216551818(.A(n_59335), .B(n_29323), .C(n_59167), .D(n_30153
		), .Z(n_220383194));
	notech_ao4 i_216651817(.A(n_55367), .B(n_28394), .C(n_59153), .D(n_29291
		), .Z(n_220483195));
	notech_and4 i_217251811(.A(n_220483195), .B(n_220383194), .C(n_220183192
		), .D(n_220083191), .Z(n_220683197));
	notech_ao4 i_219251791(.A(n_55378), .B(n_29352), .C(n_55389), .D(n_28599
		), .Z(n_220783198));
	notech_ao4 i_218751796(.A(n_55429), .B(n_56082), .C(n_55400), .D(n_27989
		), .Z(n_220883199));
	notech_ao4 i_218851795(.A(n_55347), .B(nbus_11295[6]), .C(n_55420), .D(n_30154
		), .Z(n_221183202));
	notech_ao4 i_218951794(.A(n_59176), .B(n_27809), .C(n_55409), .D(n_30155
		), .Z(n_221283203));
	notech_ao4 i_219051793(.A(n_59335), .B(n_29322), .C(n_59167), .D(n_30156
		), .Z(n_221483205));
	notech_ao4 i_219151792(.A(n_55367), .B(n_28393), .C(n_59153), .D(n_29290
		), .Z(n_221583206));
	notech_and4 i_219751786(.A(n_221583206), .B(n_221483205), .C(n_221283203
		), .D(n_221183202), .Z(n_221783208));
	notech_ao4 i_221751766(.A(n_55378), .B(n_29351), .C(n_55389), .D(n_28598
		), .Z(n_221883209));
	notech_ao4 i_221251771(.A(n_55429), .B(n_56073), .C(n_55400), .D(n_59205
		), .Z(n_221983210));
	notech_ao4 i_221351770(.A(n_55347), .B(nbus_11295[5]), .C(n_55420), .D(n_30157
		), .Z(n_222283213));
	notech_ao4 i_221451769(.A(n_59176), .B(n_27808), .C(n_55409), .D(n_30158
		), .Z(n_222383214));
	notech_ao4 i_221551768(.A(n_59335), .B(n_29321), .C(n_59167), .D(n_30159
		), .Z(n_222583216));
	notech_ao4 i_221651767(.A(n_55367), .B(n_28392), .C(n_59153), .D(n_29289
		), .Z(n_222683217));
	notech_and4 i_222251761(.A(n_222683217), .B(n_222583216), .C(n_222383214
		), .D(n_222283213), .Z(n_222883219));
	notech_ao4 i_224251741(.A(n_55378), .B(n_29350), .C(n_55389), .D(n_28597
		), .Z(n_222983220));
	notech_ao4 i_223751746(.A(n_55429), .B(n_56064), .C(n_55400), .D(n_27986
		), .Z(n_223083221));
	notech_ao4 i_223851745(.A(n_55347), .B(nbus_11295[4]), .C(n_55420), .D(n_30160
		), .Z(n_223383224));
	notech_ao4 i_223951744(.A(n_59176), .B(n_27807), .C(n_55409), .D(n_30161
		), .Z(n_223483225));
	notech_ao4 i_224051743(.A(n_59335), .B(n_29320), .C(n_59167), .D(n_30162
		), .Z(n_223683227));
	notech_ao4 i_224151742(.A(n_55367), .B(n_28391), .C(n_59153), .D(n_29288
		), .Z(n_223783228));
	notech_and4 i_224751736(.A(n_223783228), .B(n_223683227), .C(n_223483225
		), .D(n_223383224), .Z(n_223983230));
	notech_ao4 i_226751716(.A(n_55378), .B(n_29349), .C(n_55389), .D(n_28596
		), .Z(n_224083231));
	notech_ao4 i_226251721(.A(n_55429), .B(n_55983), .C(n_55400), .D(n_59223
		), .Z(n_224183232));
	notech_ao4 i_226351720(.A(n_55347), .B(nbus_11295[3]), .C(n_55420), .D(n_30163
		), .Z(n_224483235));
	notech_ao4 i_226451719(.A(n_59176), .B(n_27806), .C(n_55409), .D(n_30164
		), .Z(n_224583236));
	notech_ao4 i_226551718(.A(n_27065), .B(n_29319), .C(n_59167), .D(n_30165
		), .Z(n_224783238));
	notech_ao4 i_226651717(.A(n_55367), .B(n_28390), .C(n_59153), .D(n_29287
		), .Z(n_224883239));
	notech_and4 i_227251711(.A(n_224883239), .B(n_224783238), .C(n_224583236
		), .D(n_224483235), .Z(n_225083241));
	notech_ao4 i_229251691(.A(n_55378), .B(n_29348), .C(n_55389), .D(n_28595
		), .Z(n_225183242));
	notech_ao4 i_228751696(.A(n_55429), .B(n_55992), .C(n_55400), .D(n_59259
		), .Z(n_225283243));
	notech_ao4 i_228851695(.A(n_310347753), .B(nbus_11295[2]), .C(n_55420), 
		.D(n_30166), .Z(n_225583246));
	notech_ao4 i_228951694(.A(n_59176), .B(n_27805), .C(n_55409), .D(n_30167
		), .Z(n_225683247));
	notech_ao4 i_229051693(.A(n_59335), .B(n_29318), .C(n_59167), .D(n_30168
		), .Z(n_225883249));
	notech_ao4 i_229151692(.A(n_55367), .B(n_28389), .C(n_59153), .D(n_29286
		), .Z(n_225983250));
	notech_and4 i_229751686(.A(n_225983250), .B(n_225883249), .C(n_225683247
		), .D(n_225583246), .Z(n_226183252));
	notech_or4 i_40247307(.A(n_58184), .B(n_58498), .C(n_56367), .D(n_56284)
		, .Z(n_226283253));
	notech_or2 i_40147308(.A(n_60009), .B(n_58147), .Z(n_226583256));
	notech_or4 i_39647313(.A(n_62856), .B(n_58498), .C(n_62824), .D(n_57680)
		, .Z(n_227083261));
	notech_or2 i_64047079(.A(n_138168398), .B(n_57680), .Z(n_227183262));
	notech_or4 i_63947080(.A(n_58133), .B(n_58497), .C(n_56423), .D(n_56284)
		, .Z(n_227483265));
	notech_or4 i_63447085(.A(n_58497), .B(n_54814), .C(nbus_11295[16]), .D(n_60933
		), .Z(n_227983270));
	notech_or4 i_79246932(.A(n_54756), .B(n_58494), .C(n_56432), .D(n_56284)
		, .Z(n_228083271));
	notech_or2 i_79146933(.A(n_60009), .B(n_58141), .Z(n_228383274));
	notech_nand2 i_78646938(.A(\regs_13_14[16] ), .B(n_26675), .Z(n_228883279
		));
	notech_or2 i_83546889(.A(n_57861), .B(n_57680), .Z(n_228983280));
	notech_nand3 i_83046894(.A(opc_10[16]), .B(n_62824), .C(n_57115), .Z(n_229683287
		));
	notech_or2 i_88046848(.A(n_60009), .B(n_58138), .Z(n_229783288));
	notech_or2 i_87846849(.A(n_57867), .B(n_57680), .Z(n_230083291));
	notech_or4 i_87046854(.A(n_56863), .B(n_54727), .C(n_254466073), .D(n_58504
		), .Z(n_230583296));
	notech_ao4 i_186245902(.A(n_58008), .B(n_252966058), .C(n_56636), .D(n_311224366
		), .Z(n_230683297));
	notech_ao4 i_186145903(.A(n_29710), .B(n_26937), .C(n_124271722), .D(n_313747721
		), .Z(n_230883299));
	notech_ao4 i_185845906(.A(n_57865), .B(n_56284), .C(n_57726), .D(n_28142
		), .Z(n_231083301));
	notech_and4 i_186045904(.A(n_194675885), .B(n_231083301), .C(n_229783288
		), .D(n_230083291), .Z(n_231383304));
	notech_ao4 i_182545938(.A(n_252966058), .B(n_286927251), .C(n_56662), .D
		(n_311224366), .Z(n_231483305));
	notech_ao4 i_182445939(.A(n_29710), .B(n_26615), .C(n_143571915), .D(n_313747721
		), .Z(n_231683307));
	notech_ao4 i_182245941(.A(n_57863), .B(n_56284), .C(n_60009), .D(n_58139
		), .Z(n_231883309));
	notech_and3 i_182345940(.A(n_194675885), .B(n_231883309), .C(n_228983280
		), .Z(n_232083311));
	notech_ao4 i_178445976(.A(n_252966058), .B(n_307124335), .C(n_241472894)
		, .D(n_57680), .Z(n_232183312));
	notech_ao4 i_178345977(.A(n_58494), .B(n_312324377), .C(n_311224366), .D
		(n_56649), .Z(n_232383314));
	notech_ao4 i_178045980(.A(n_313747721), .B(n_147271952), .C(n_254466073)
		, .D(n_57116), .Z(n_232583316));
	notech_and4 i_178245978(.A(n_194675885), .B(n_232583316), .C(n_228083271
		), .D(n_228383274), .Z(n_232883319));
	notech_ao4 i_165346105(.A(n_58497), .B(n_312324377), .C(n_56498), .D(n_311224366
		), .Z(n_232983320));
	notech_ao4 i_165246106(.A(n_313747721), .B(n_304273522), .C(n_254466073)
		, .D(n_57596), .Z(n_233183322));
	notech_ao4 i_164946109(.A(n_60009), .B(n_58145), .C(n_26918), .D(n_29710
		), .Z(n_233383324));
	notech_and4 i_165146107(.A(n_194675885), .B(n_233383324), .C(n_227183262
		), .D(n_227483265), .Z(n_233683327));
	notech_ao4 i_145746293(.A(n_311224366), .B(n_56485), .C(n_241372893), .D
		(n_57680), .Z(n_233783328));
	notech_ao4 i_145646294(.A(n_254466073), .B(n_235883349), .C(n_252966058)
		, .D(n_58084), .Z(n_233983330));
	notech_ao4 i_145346297(.A(n_29710), .B(n_26929), .C(n_313747721), .D(n_303673516
		), .Z(n_234183332));
	notech_and4 i_145546295(.A(n_234183332), .B(n_194675885), .C(n_226283253
		), .D(n_226583256), .Z(n_234483335));
	notech_and4 i_9144403(.A(n_56843), .B(n_23512), .C(n_234983340), .D(n_27024
		), .Z(n_234583336));
	notech_ao4 i_16744329(.A(n_29619), .B(n_316191662), .C(n_314791676), .D(n_23507
		), .Z(n_234683337));
	notech_or2 i_22044276(.A(n_4011), .B(n_32408), .Z(n_234983340));
	notech_and4 i_9044404(.A(n_56843), .B(n_25010), .C(n_235783348), .D(n_27024
		), .Z(n_235083341));
	notech_ao4 i_15944337(.A(n_311891705), .B(n_29619), .C(n_311991704), .D(\nbus_11365[31] 
		), .Z(n_235183342));
	notech_ao4 i_16044336(.A(n_24996), .B(n_311991704), .C(n_60268), .D(n_26984
		), .Z(n_235283343));
	notech_or2 i_32744169(.A(n_4011), .B(n_32295), .Z(n_235783348));
	notech_and2 i_148844545(.A(n_57915), .B(n_236083351), .Z(n_235883349));
	notech_or2 i_75643769(.A(n_56675), .B(n_314391680), .Z(n_235983350));
	notech_or4 i_124943313(.A(n_57078), .B(n_57051), .C(n_54916), .D(n_236183352
		), .Z(n_236083351));
	notech_and3 i_10644389(.A(n_56843), .B(n_188562161), .C(n_58482), .Z(n_236183352
		));
	notech_ao3 i_21744279(.A(tsc[31]), .B(n_55820), .C(n_59469), .Z(n_236283353
		));
	notech_or4 i_21044286(.A(n_60935), .B(n_28157), .C(n_26942), .D(n_234583336
		), .Z(n_236783358));
	notech_nand3 i_21144285(.A(opc[31]), .B(n_60298), .C(n_58088), .Z(n_236883359
		));
	notech_or2 i_21244284(.A(n_234683337), .B(n_316391660), .Z(n_236983360)
		);
	notech_ao3 i_32244174(.A(tsc[63]), .B(n_55820), .C(n_59469), .Z(n_237083361
		));
	notech_or4 i_31644180(.A(n_26939), .B(n_60935), .C(n_28157), .D(n_235083341
		), .Z(n_237583366));
	notech_or4 i_31744179(.A(n_314891675), .B(n_311891705), .C(n_314791676),
		 .D(n_57976), .Z(n_237683367));
	notech_or4 i_36844128(.A(n_54954), .B(n_3845), .C(n_58020), .D(n_57837),
		 .Z(n_237783368));
	notech_nao3 i_36344133(.A(n_62822), .B(opc_10[31]), .C(n_57595), .Z(n_238483375
		));
	notech_nand2 i_47544026(.A(\regs_13_14[31] ), .B(n_58148), .Z(n_238583376
		));
	notech_or2 i_105243495(.A(n_57726), .B(n_28157), .Z(n_239283383));
	notech_nand2 i_105143496(.A(\regs_13_14[31] ), .B(n_57569), .Z(n_239583386
		));
	notech_nao3 i_104643501(.A(n_62820), .B(opc_10[31]), .C(n_58007), .Z(n_240083391
		));
	notech_ao4 i_201142579(.A(n_96519147), .B(n_58008), .C(n_56636), .D(n_306221226
		), .Z(n_240183392));
	notech_ao4 i_201042580(.A(n_57867), .B(n_59726), .C(n_314391680), .D(n_124271722
		), .Z(n_240383394));
	notech_ao4 i_200742583(.A(n_57865), .B(n_57837), .C(n_314791676), .D(n_58138
		), .Z(n_240583396));
	notech_and4 i_200942581(.A(n_240583396), .B(n_26710), .C(n_239283383), .D
		(n_239583386), .Z(n_240883399));
	notech_ao4 i_154443041(.A(n_96519147), .B(n_58084), .C(n_56485), .D(n_303721201
		), .Z(n_240983400));
	notech_ao4 i_154343042(.A(n_57868), .B(n_59726), .C(n_83019012), .D(n_235883349
		), .Z(n_241083401));
	notech_ao4 i_154143044(.A(n_57875), .B(n_57837), .C(n_314791676), .D(n_58147
		), .Z(n_241283403));
	notech_and3 i_154243043(.A(n_241283403), .B(n_26710), .C(n_238583376), .Z
		(n_241483405));
	notech_ao4 i_144743124(.A(n_3858), .B(n_96519147), .C(n_306221226), .D(n_56601
		), .Z(n_241583406));
	notech_ao4 i_144643125(.A(n_26642), .B(n_29619), .C(n_314391680), .D(n_147671956
		), .Z(n_241783408));
	notech_ao4 i_144443127(.A(n_3878), .B(n_59726), .C(n_148228759), .D(n_314791676
		), .Z(n_241983410));
	notech_and3 i_144543126(.A(n_241983410), .B(n_26710), .C(n_237783368), .Z
		(n_242183412));
	notech_ao4 i_140643161(.A(n_235283343), .B(n_57837), .C(n_235183342), .D
		(n_312291701), .Z(n_242783418));
	notech_nand3 i_140843159(.A(n_237683367), .B(n_237583366), .C(n_242783418
		), .Z(n_242883419));
	notech_ao4 i_140443163(.A(n_310891715), .B(n_96519147), .C(n_56532), .D(n_303721201
		), .Z(n_242983420));
	notech_ao4 i_130943254(.A(n_96519147), .B(n_311491709), .C(n_56579), .D(n_303721201
		), .Z(n_243783428));
	notech_and4 i_131243251(.A(n_236783358), .B(n_243783428), .C(n_236883359
		), .D(n_236983360), .Z(n_243883429));
	notech_ao4 i_130743256(.A(n_311191712), .B(n_57837), .C(n_311091713), .D
		(n_59726), .Z(n_243983430));
	notech_nao3 i_16441096(.A(n_60298), .B(mul64[24]), .C(n_2647), .Z(n_244683437
		));
	notech_or4 i_16141099(.A(n_60893), .B(n_60268), .C(n_26965), .D(nbus_11295
		[16]), .Z(n_244983440));
	notech_ao4 i_113640206(.A(n_55886), .B(n_56028), .C(n_57367), .D(n_56118
		), .Z(n_245483445));
	notech_ao4 i_113540207(.A(n_227976218), .B(n_30171), .C(n_60372), .D(n_29386
		), .Z(n_245583446));
	notech_ao4 i_113340209(.A(n_308084071), .B(nbus_11328[8]), .C(n_307884069
		), .D(n_30170), .Z(n_245783448));
	notech_and4 i_113840204(.A(n_245783448), .B(n_245583446), .C(n_245483445
		), .D(n_244983440), .Z(n_245983450));
	notech_ao4 i_113040212(.A(n_307584066), .B(n_28113), .C(n_3892), .D(nbus_11295
		[24]), .Z(n_246083451));
	notech_ao4 i_112840214(.A(n_307484065), .B(n_30169), .C(n_58651), .D(n_28134
		), .Z(n_246283453));
	notech_and4 i_113240210(.A(n_307384064), .B(n_246283453), .C(n_246083451
		), .D(n_244683437), .Z(n_246483455));
	notech_or4 i_2238212(.A(instrc[122]), .B(n_32614), .C(instrc[121]), .D(n_58813
		), .Z(n_246583456));
	notech_ao4 i_5438187(.A(n_32614), .B(n_32342), .C(n_246883459), .D(n_28049
		), .Z(n_246683457));
	notech_and2 i_4138193(.A(n_58009), .B(n_60841), .Z(n_246883459));
	notech_and2 i_5238188(.A(n_299783988), .B(n_56391), .Z(n_246983460));
	notech_and2 i_5038190(.A(n_276383754), .B(n_247183462), .Z(n_247083461)
		);
	notech_or4 i_25837985(.A(instrc[122]), .B(n_54912649), .C(n_29179), .D(n_26735
		), .Z(n_247183462));
	notech_ao4 i_39137863(.A(n_330763524), .B(n_305047803), .C(n_25629), .D(n_27105
		), .Z(n_247283463));
	notech_or4 i_60537661(.A(n_60854), .B(n_54912649), .C(n_26735), .D(n_29022
		), .Z(n_247583466));
	notech_or4 i_61937647(.A(instrc[122]), .B(n_32339), .C(instrc[121]), .D(n_29736
		), .Z(n_247683467));
	notech_and3 i_2938205(.A(n_248283473), .B(n_248183472), .C(n_248083471),
		 .Z(n_247983470));
	notech_or4 i_62237644(.A(n_2888), .B(n_59419), .C(n_32443), .D(n_56109),
		 .Z(n_248083471));
	notech_or4 i_62337643(.A(n_62856), .B(n_58220), .C(n_60935), .D(n_56275)
		, .Z(n_248183472));
	notech_or4 i_62437642(.A(n_25625), .B(n_25617), .C(n_60894), .D(n_56109)
		, .Z(n_248283473));
	notech_nand2 i_10438138(.A(resb_shiftbox[0]), .B(n_27003), .Z(n_248683477
		));
	notech_or4 i_10138141(.A(n_25625), .B(n_25617), .C(n_303747815), .D(n_59187
		), .Z(n_248983480));
	notech_or2 i_9838144(.A(n_388360286), .B(nbus_11295[0]), .Z(n_249283483)
		);
	notech_or2 i_9538147(.A(n_33512435), .B(n_28001), .Z(n_249583486));
	notech_nao3 i_9238150(.A(nbus_160[0]), .B(n_26782), .C(n_52112621), .Z(n_249883489
		));
	notech_nand2 i_8938153(.A(read_data[8]), .B(n_19512295), .Z(n_250183492)
		);
	notech_nao3 i_8638156(.A(n_295960040), .B(imm[0]), .C(n_54912649), .Z(n_250483495
		));
	notech_nand2 i_12838115(.A(resb_shiftbox[1]), .B(n_27003), .Z(n_250883499
		));
	notech_or4 i_12538118(.A(n_25625), .B(n_59478), .C(n_57132), .D(n_59241)
		, .Z(n_251183502));
	notech_or2 i_12238121(.A(n_388360286), .B(nbus_11295[1]), .Z(n_251483505
		));
	notech_or2 i_11838124(.A(n_33512435), .B(n_28002), .Z(n_251783508));
	notech_nao3 i_11538127(.A(nbus_160[1]), .B(n_26782), .C(n_52112621), .Z(n_252083511
		));
	notech_nand2 i_11238130(.A(read_data[9]), .B(n_19512295), .Z(n_252383514
		));
	notech_nao3 i_10938133(.A(imm[1]), .B(n_295960040), .C(n_54912649), .Z(n_252683517
		));
	notech_nand2 i_17538068(.A(resb_shiftbox[3]), .B(n_27003), .Z(n_253283523
		));
	notech_or4 i_17238071(.A(n_25625), .B(n_59478), .C(n_57132), .D(n_59223)
		, .Z(n_253583526));
	notech_or2 i_16938074(.A(n_388360286), .B(nbus_11295[3]), .Z(n_253883529
		));
	notech_or2 i_16438079(.A(n_54512645), .B(n_56181), .Z(n_254383534));
	notech_nand3 i_16138082(.A(n_309160172), .B(n_309460175), .C(read_data[
		27]), .Z(n_254683537));
	notech_nand2 i_15838085(.A(add_src[3]), .B(n_27001), .Z(n_254983540));
	notech_nand2 i_19638047(.A(resb_shiftbox[4]), .B(n_27003), .Z(n_255383544
		));
	notech_or4 i_19338050(.A(n_58086), .B(n_59478), .C(n_57132), .D(n_27986)
		, .Z(n_255683547));
	notech_or2 i_19038053(.A(n_388360286), .B(nbus_11295[4]), .Z(n_255983550
		));
	notech_or2 i_18538058(.A(n_54512645), .B(n_56221), .Z(n_256483555));
	notech_nand3 i_18238061(.A(n_309160172), .B(read_data[28]), .C(n_309460175
		), .Z(n_256783558));
	notech_nand2 i_17938064(.A(add_src[4]), .B(n_27001), .Z(n_257083561));
	notech_nand2 i_21638027(.A(resb_shiftbox[5]), .B(n_27003), .Z(n_257483565
		));
	notech_nao3 i_21138032(.A(n_308960170), .B(resb_shift4box[5]), .C(n_308760168
		), .Z(n_257983570));
	notech_nao3 i_20638037(.A(imm[37]), .B(n_25374), .C(n_57132), .Z(n_258483575
		));
	notech_nand2 i_20338040(.A(read_data[21]), .B(n_18912289), .Z(n_258783578
		));
	notech_nand2 i_20038043(.A(read_data[5]), .B(n_27002), .Z(n_259083581)
		);
	notech_or2 i_3038204(.A(n_54912649), .B(n_308815164), .Z(n_259183582));
	notech_nand2 i_23638007(.A(resb_shiftbox[6]), .B(n_27003), .Z(n_259583586
		));
	notech_nao3 i_23138012(.A(n_308960170), .B(resb_shift4box[6]), .C(n_308760168
		), .Z(n_260083591));
	notech_nao3 i_22638017(.A(imm[38]), .B(n_25374), .C(n_57132), .Z(n_260583596
		));
	notech_nand2 i_22338020(.A(read_data[22]), .B(n_18912289), .Z(n_260883599
		));
	notech_nand2 i_22038023(.A(n_27002), .B(read_data[6]), .Z(n_261183602)
		);
	notech_or2 i_25737986(.A(n_55886), .B(nbus_11295[15]), .Z(n_261283603)
		);
	notech_nand2 i_25637987(.A(resb_shiftbox[7]), .B(n_27003), .Z(n_261583606
		));
	notech_nao3 i_25137992(.A(resb_shift4box[7]), .B(n_308960170), .C(n_308760168
		), .Z(n_262083611));
	notech_ao3 i_24637997(.A(imm[39]), .B(n_25374), .C(n_57132), .Z(n_262583616
		));
	notech_nand2 i_24138002(.A(read_data[7]), .B(n_27002), .Z(n_263083621)
		);
	notech_or2 i_27837966(.A(n_55886), .B(n_56475), .Z(n_263183622));
	notech_nor2 i_27337971(.A(n_53512635), .B(n_27991), .Z(n_263883629));
	notech_nand2 i_26337980(.A(n_27001), .B(add_src[8]), .Z(n_264783638));
	notech_or2 i_29537949(.A(n_55886), .B(\nbus_11358[25] ), .Z(n_264883639)
		);
	notech_nor2 i_29037954(.A(n_53512635), .B(n_27992), .Z(n_265583646));
	notech_nand2 i_28137963(.A(n_27001), .B(add_src[9]), .Z(n_266483655));
	notech_or2 i_31237932(.A(n_55885), .B(\nbus_11358[26] ), .Z(n_266583656)
		);
	notech_nor2 i_30737937(.A(n_53512635), .B(n_27993), .Z(n_267283663));
	notech_nand2 i_29837946(.A(add_src[10]), .B(n_27001), .Z(n_268183672));
	notech_or2 i_32937915(.A(n_55885), .B(n_55938), .Z(n_268283673));
	notech_or4 i_32437920(.A(n_58086), .B(n_59478), .C(n_57132), .D(n_27996)
		, .Z(n_268983680));
	notech_nand2 i_31537929(.A(n_27001), .B(add_src[11]), .Z(n_269883689));
	notech_or2 i_36437881(.A(n_55885), .B(\nbus_11358[29] ), .Z(n_269983690)
		);
	notech_or4 i_35937886(.A(n_58086), .B(n_59478), .C(n_57132), .D(n_27998)
		, .Z(n_270683697));
	notech_nand2 i_34937895(.A(n_27001), .B(add_src[13]), .Z(n_271583706));
	notech_or2 i_39037864(.A(n_55885), .B(n_55929), .Z(n_271683707));
	notech_nor2 i_38437869(.A(n_53512635), .B(n_27999), .Z(n_272383714));
	notech_nand2 i_36737878(.A(n_27001), .B(add_src[14]), .Z(n_273283723));
	notech_or4 i_39237862(.A(n_58220), .B(n_62834), .C(n_60938), .D(n_60252)
		, .Z(n_273383724));
	notech_or2 i_41537844(.A(n_55885), .B(n_57837), .Z(n_273483725));
	notech_nor2 i_41037849(.A(n_53512635), .B(n_28000), .Z(n_274183732));
	notech_or2 i_40537854(.A(n_33512435), .B(n_28016), .Z(n_274683737));
	notech_or2 i_40037859(.A(n_3888), .B(n_28104), .Z(n_275083741));
	notech_or2 i_45837808(.A(n_3864), .B(n_53612636), .Z(n_275583746));
	notech_or2 i_45537811(.A(n_54212642), .B(n_57698), .Z(n_275883749));
	notech_or2 i_94638224(.A(n_54912649), .B(n_56405), .Z(n_276383754));
	notech_or4 i_170336603(.A(n_25629), .B(n_60935), .C(n_60910), .D(n_60252
		), .Z(n_276483755));
	notech_ao4 i_39938233(.A(n_247983470), .B(n_60252), .C(n_276483755), .D(n_56275
		), .Z(n_276883759));
	notech_and3 i_2038214(.A(n_276883759), .B(n_259183582), .C(n_247583466),
		 .Z(n_277183762));
	notech_ao4 i_155436751(.A(n_276383754), .B(n_29046), .C(n_3888), .D(n_28107
		), .Z(n_277283763));
	notech_ao4 i_155336752(.A(n_310315179), .B(n_56302), .C(n_3887), .D(n_29072
		), .Z(n_277383764));
	notech_ao4 i_155136754(.A(n_54012640), .B(n_29270), .C(n_388360286), .D(nbus_11295
		[18]), .Z(n_277583766));
	notech_and4 i_155636749(.A(n_277583766), .B(n_277383764), .C(n_277283763
		), .D(n_275883749), .Z(n_277783768));
	notech_ao4 i_154836757(.A(n_53412634), .B(n_29668), .C(n_53512635), .D(n_28003
		), .Z(n_277883769));
	notech_ao4 i_154636759(.A(n_3882), .B(n_29235), .C(n_52112621), .D(n_29198
		), .Z(n_278083771));
	notech_and4 i_155036755(.A(n_277183762), .B(n_278083771), .C(n_277883769
		), .D(n_275583746), .Z(n_278283773));
	notech_ao4 i_151336792(.A(n_34012440), .B(n_56275), .C(n_60252), .D(n_247983470
		), .Z(n_278383774));
	notech_ao4 i_151236793(.A(n_3887), .B(n_29067), .C(n_276383754), .D(n_29028
		), .Z(n_278583776));
	notech_nand3 i_151536790(.A(n_278383774), .B(n_278583776), .C(n_275083741
		), .Z(n_278683777));
	notech_ao4 i_150936796(.A(n_33312433), .B(n_29045), .C(n_33412434), .D(n_29194
		), .Z(n_278783778));
	notech_ao4 i_150836797(.A(n_388360286), .B(nbus_11295[15]), .C(n_33012430
		), .D(n_29002), .Z(n_278983780));
	notech_nand3 i_151136794(.A(n_278783778), .B(n_278983780), .C(n_274683737
		), .Z(n_279083781));
	notech_ao4 i_150436801(.A(n_54212642), .B(n_57671), .C(n_54012640), .D(n_29267
		), .Z(n_279283783));
	notech_ao4 i_150336802(.A(n_60010), .B(n_53612636), .C(n_53412634), .D(n_29649
		), .Z(n_279483785));
	notech_nao3 i_150636799(.A(n_279283783), .B(n_279483785), .C(n_274183732
		), .Z(n_279583786));
	notech_ao4 i_150136804(.A(n_3892), .B(nbus_11295[7]), .C(n_3882), .D(n_29232
		), .Z(n_279683787));
	notech_ao4 i_3938195(.A(n_54912649), .B(n_328270293), .C(n_54512645), .D
		(n_56275), .Z(n_279783788));
	notech_nand3 i_150236803(.A(n_279783788), .B(n_279683787), .C(n_273483725
		), .Z(n_279983790));
	notech_ao4 i_149536810(.A(n_276383754), .B(n_29027), .C(n_3888), .D(n_28103
		), .Z(n_280183792));
	notech_ao4 i_149436811(.A(n_33412434), .B(n_29192), .C(n_309615172), .D(n_56248
		), .Z(n_280483795));
	notech_and3 i_149736808(.A(n_280183792), .B(n_280483795), .C(n_273283723
		), .Z(n_280583796));
	notech_ao4 i_149236813(.A(n_33512435), .B(n_28015), .C(n_33312433), .D(n_29044
		), .Z(n_280683797));
	notech_ao4 i_149136814(.A(n_388360286), .B(nbus_11295[14]), .C(n_33012430
		), .D(n_29001), .Z(n_280783798));
	notech_ao4 i_148736818(.A(n_54212642), .B(n_57662), .C(n_54012640), .D(n_29266
		), .Z(n_281083801));
	notech_ao4 i_148636819(.A(n_60011), .B(n_53612636), .C(n_53412634), .D(n_29648
		), .Z(n_281283803));
	notech_ao3 i_148936816(.A(n_281083801), .B(n_281283803), .C(n_272383714)
		, .Z(n_281383804));
	notech_ao4 i_148436821(.A(n_3892), .B(nbus_11295[6]), .C(n_3882), .D(n_29231
		), .Z(n_281483805));
	notech_and3 i_3238202(.A(n_259183582), .B(n_247583466), .C(n_309515171),
		 .Z(n_281583806));
	notech_and4 i_149036815(.A(n_281583806), .B(n_281483805), .C(n_281383804
		), .D(n_271683707), .Z(n_281883809));
	notech_ao4 i_147936826(.A(n_276383754), .B(n_29026), .C(n_3888), .D(n_28102
		), .Z(n_281983810));
	notech_ao4 i_147836827(.A(n_33412434), .B(n_29191), .C(n_309615172), .D(\nbus_11358[13] 
		), .Z(n_282183812));
	notech_and3 i_148136824(.A(n_281983810), .B(n_282183812), .C(n_271583706
		), .Z(n_282283813));
	notech_ao4 i_147636829(.A(n_33512435), .B(n_28014), .C(n_33312433), .D(n_29043
		), .Z(n_282383814));
	notech_ao4 i_147536830(.A(n_388360286), .B(nbus_11295[13]), .C(n_33012430
		), .D(n_29000), .Z(n_282483815));
	notech_ao4 i_147136834(.A(n_54212642), .B(n_57653), .C(n_54012640), .D(n_29265
		), .Z(n_282783818));
	notech_ao4 i_147036835(.A(n_302091803), .B(n_53612636), .C(n_53412634), 
		.D(n_29650), .Z(n_282983820));
	notech_and3 i_147336832(.A(n_282783818), .B(n_282983820), .C(n_270683697
		), .Z(n_283083821));
	notech_ao4 i_146836837(.A(n_3892), .B(nbus_11295[5]), .C(n_3882), .D(n_29229
		), .Z(n_283183822));
	notech_and4 i_147436831(.A(n_281583806), .B(n_283183822), .C(n_269983690
		), .D(n_283083821), .Z(n_283483825));
	notech_ao4 i_144736858(.A(n_276383754), .B(n_29025), .C(n_3888), .D(n_28100
		), .Z(n_283583826));
	notech_ao4 i_144636859(.A(n_33412434), .B(n_29189), .C(n_309615172), .D(n_56181
		), .Z(n_283783828));
	notech_and3 i_144936856(.A(n_283583826), .B(n_283783828), .C(n_269883689
		), .Z(n_283883829));
	notech_ao4 i_144436861(.A(n_33512435), .B(n_28012), .C(n_33312433), .D(n_29042
		), .Z(n_283983830));
	notech_ao4 i_144336862(.A(n_388360286), .B(nbus_11295[11]), .C(n_33012430
		), .D(n_28998), .Z(n_284083831));
	notech_ao4 i_143936866(.A(n_54212642), .B(n_57635), .C(n_54012640), .D(n_29263
		), .Z(n_284383834));
	notech_ao4 i_143836867(.A(n_302491799), .B(n_53612636), .C(n_53412634), 
		.D(n_29646), .Z(n_284583836));
	notech_and3 i_144136864(.A(n_284383834), .B(n_284583836), .C(n_268983680
		), .Z(n_284683837));
	notech_ao4 i_143636869(.A(n_3892), .B(n_57909), .C(n_3882), .D(n_29227),
		 .Z(n_284783838));
	notech_and4 i_144236863(.A(n_342670437), .B(n_284783838), .C(n_268283673
		), .D(n_284683837), .Z(n_285083841));
	notech_ao4 i_143136874(.A(n_276383754), .B(n_29033), .C(n_3888), .D(n_28099
		), .Z(n_285183842));
	notech_ao4 i_143036875(.A(n_33412434), .B(n_29188), .C(n_309615172), .D(n_56154
		), .Z(n_285383844));
	notech_and3 i_143336872(.A(n_285183842), .B(n_285383844), .C(n_268183672
		), .Z(n_285483845));
	notech_ao4 i_142836877(.A(n_33512435), .B(n_28011), .C(n_33312433), .D(n_29041
		), .Z(n_285583846));
	notech_ao4 i_142736878(.A(n_388360286), .B(nbus_11295[10]), .C(n_33012430
		), .D(n_28997), .Z(n_285683847));
	notech_ao4 i_142336882(.A(n_54212642), .B(n_57625), .C(n_54012640), .D(n_29261
		), .Z(n_285983850));
	notech_ao4 i_142236883(.A(n_3850), .B(n_53612636), .C(n_53412634), .D(n_29644
		), .Z(n_286183852));
	notech_ao3 i_142536880(.A(n_285983850), .B(n_286183852), .C(n_267283663)
		, .Z(n_286283853));
	notech_ao4 i_142036885(.A(n_3892), .B(nbus_11295[2]), .C(n_3882), .D(n_29226
		), .Z(n_286383854));
	notech_and4 i_142636879(.A(n_281583806), .B(n_286383854), .C(n_286283853
		), .D(n_266583656), .Z(n_286683857));
	notech_ao4 i_141436890(.A(n_55791), .B(n_29024), .C(n_55782), .D(n_28098
		), .Z(n_286783858));
	notech_ao4 i_141336891(.A(n_33412434), .B(n_29187), .C(n_309615172), .D(n_56136
		), .Z(n_286983860));
	notech_and3 i_141636888(.A(n_286783858), .B(n_286983860), .C(n_266483655
		), .Z(n_287083861));
	notech_ao4 i_141136893(.A(n_33512435), .B(n_28010), .C(n_33312433), .D(n_29040
		), .Z(n_287183862));
	notech_ao4 i_141036894(.A(n_55809), .B(nbus_11295[9]), .C(n_33012430), .D
		(n_28996), .Z(n_287283863));
	notech_ao4 i_140636898(.A(n_54212642), .B(n_57613), .C(n_54012640), .D(n_29258
		), .Z(n_287583866));
	notech_ao4 i_140536899(.A(n_53612636), .B(n_60016), .C(n_53412634), .D(n_29643
		), .Z(n_287783868));
	notech_ao3 i_140836896(.A(n_287583866), .B(n_287783868), .C(n_265583646)
		, .Z(n_287883869));
	notech_ao4 i_140336901(.A(n_3892), .B(nbus_11295[1]), .C(n_3882), .D(n_29222
		), .Z(n_287983870));
	notech_and4 i_140936895(.A(n_287983870), .B(n_281583806), .C(n_287883869
		), .D(n_264883639), .Z(n_288283873));
	notech_ao4 i_139836906(.A(n_55791), .B(n_29023), .C(n_55782), .D(n_28097
		), .Z(n_288383874));
	notech_ao4 i_139736907(.A(n_33412434), .B(n_29186), .C(n_309615172), .D(n_56118
		), .Z(n_288583876));
	notech_and3 i_140036904(.A(n_288383874), .B(n_288583876), .C(n_264783638
		), .Z(n_288683877));
	notech_ao4 i_139536909(.A(n_33512435), .B(n_28009), .C(n_33312433), .D(n_29039
		), .Z(n_288783878));
	notech_ao4 i_139436910(.A(n_55809), .B(nbus_11295[8]), .C(n_33012430), .D
		(n_28995), .Z(n_288883879));
	notech_ao4 i_139036914(.A(n_54212642), .B(n_57604), .C(n_54012640), .D(n_29255
		), .Z(n_289183882));
	notech_ao4 i_138936915(.A(n_5933), .B(n_53612636), .C(n_53412634), .D(n_29645
		), .Z(n_289383884));
	notech_ao3 i_139236912(.A(n_289183882), .B(n_289383884), .C(n_263883629)
		, .Z(n_289483885));
	notech_ao4 i_138736917(.A(n_3892), .B(n_59717), .C(n_55891), .D(n_29218)
		, .Z(n_289583886));
	notech_and4 i_139336911(.A(n_342670437), .B(n_289583886), .C(n_289483885
		), .D(n_263183622), .Z(n_289883889));
	notech_ao4 i_137536929(.A(n_3887), .B(n_29060), .C(n_247083461), .D(n_29022
		), .Z(n_289983890));
	notech_ao4 i_137436930(.A(n_28123), .B(n_19312293), .C(n_26949), .D(n_28104
		), .Z(n_290183892));
	notech_ao4 i_137136933(.A(n_33412434), .B(n_29185), .C(n_26948), .D(n_28112
		), .Z(n_290383894));
	notech_ao4 i_137036934(.A(n_33012430), .B(n_28994), .C(n_33512435), .D(n_28008
		), .Z(n_290583896));
	notech_ao3 i_137336931(.A(n_290383894), .B(n_290583896), .C(n_262583616)
		, .Z(n_290683897));
	notech_and4 i_137836926(.A(n_289983890), .B(n_290183892), .C(n_263083621
		), .D(n_290683897), .Z(n_290783898));
	notech_ao4 i_136636938(.A(n_55809), .B(nbus_11295[7]), .C(n_388560287), 
		.D(n_56109), .Z(n_290883899));
	notech_ao4 i_136536939(.A(n_53512635), .B(n_56100), .C(n_54212642), .D(n_57957
		), .Z(n_291083901));
	notech_and3 i_136836936(.A(n_290883899), .B(n_291083901), .C(n_262083611
		), .Z(n_291183902));
	notech_ao4 i_136236942(.A(n_303191792), .B(n_53612636), .C(n_53412634), 
		.D(n_29174), .Z(n_291283903));
	notech_and4 i_136436940(.A(n_279783788), .B(n_291283903), .C(n_261283603
		), .D(n_261583606), .Z(n_291583906));
	notech_ao4 i_135636948(.A(n_3887), .B(n_29056), .C(n_17012270), .D(n_29021
		), .Z(n_291783908));
	notech_ao4 i_135436950(.A(n_19312293), .B(n_28121), .C(n_26949), .D(n_28103
		), .Z(n_291983910));
	notech_and4 i_135836946(.A(n_291983910), .B(n_291783908), .C(n_260883599
		), .D(n_261183602), .Z(n_292183912));
	notech_ao4 i_135136953(.A(n_54512645), .B(n_56248), .C(n_33412434), .D(n_29184
		), .Z(n_292283913));
	notech_ao4 i_135036954(.A(n_33012430), .B(n_28993), .C(n_33512435), .D(n_28007
		), .Z(n_292483915));
	notech_and3 i_135336951(.A(n_292283913), .B(n_292483915), .C(n_260583596
		), .Z(n_292583916));
	notech_ao4 i_134636958(.A(n_55809), .B(nbus_11295[6]), .C(n_388560287), 
		.D(n_56082), .Z(n_292783918));
	notech_ao4 i_134536959(.A(n_55829), .B(n_27989), .C(n_55869), .D(n_57592
		), .Z(n_292983920));
	notech_and3 i_134836956(.A(n_292783918), .B(n_292983920), .C(n_260083591
		), .Z(n_293083921));
	notech_ao4 i_134236962(.A(n_3874), .B(n_55849), .C(n_55838), .D(n_29173)
		, .Z(n_293183922));
	notech_ao4 i_134136963(.A(n_55885), .B(nbus_11295[14]), .C(n_55909), .D(n_308815164
		), .Z(n_293383924));
	notech_and4 i_134936955(.A(n_293183922), .B(n_293383924), .C(n_259583586
		), .D(n_293083921), .Z(n_293583926));
	notech_ao4 i_133636967(.A(n_3887), .B(n_29055), .C(n_17012270), .D(n_29017
		), .Z(n_293683927));
	notech_ao4 i_133436969(.A(n_19312293), .B(n_28118), .C(n_26949), .D(n_28102
		), .Z(n_293883929));
	notech_and4 i_133836965(.A(n_293883929), .B(n_293683927), .C(n_258783578
		), .D(n_259083581), .Z(n_294083931));
	notech_ao4 i_133136972(.A(n_54512645), .B(n_56230), .C(n_33412434), .D(n_29183
		), .Z(n_294183932));
	notech_ao4 i_133036973(.A(n_33012430), .B(n_28992), .C(n_33512435), .D(n_28006
		), .Z(n_294383934));
	notech_and3 i_133336970(.A(n_294183932), .B(n_294383934), .C(n_258483575
		), .Z(n_294483935));
	notech_ao4 i_132636977(.A(n_55809), .B(nbus_11295[5]), .C(n_388560287), 
		.D(n_56073), .Z(n_294683937));
	notech_ao4 i_132536978(.A(n_55829), .B(n_27987), .C(n_55869), .D(n_57583
		), .Z(n_294883939));
	notech_and3 i_132836975(.A(n_294683937), .B(n_294883939), .C(n_257983570
		), .Z(n_294983940));
	notech_ao4 i_132236981(.A(n_60020), .B(n_55849), .C(n_55838), .D(n_29172
		), .Z(n_295083941));
	notech_ao4 i_132136982(.A(n_55909), .B(n_308815164), .C(n_55886), .D(nbus_11295
		[13]), .Z(n_295283943));
	notech_and4 i_132936974(.A(n_295083941), .B(n_295283943), .C(n_257483565
		), .D(n_294983940), .Z(n_295483945));
	notech_or4 i_132036983(.A(opz[0]), .B(opz[1]), .C(n_28051), .D(n_56396),
		 .Z(n_295583946));
	notech_ao4 i_131636987(.A(n_17012270), .B(n_29016), .C(n_55909), .D(n_295583946
		), .Z(n_295683947));
	notech_ao4 i_131436989(.A(n_26949), .B(n_28101), .C(n_3886), .D(n_28093)
		, .Z(n_295883949));
	notech_and4 i_131836985(.A(n_295883949), .B(n_295683947), .C(n_257083561
		), .D(n_256783558), .Z(n_296083951));
	notech_ao4 i_131136992(.A(n_33412434), .B(n_29182), .C(n_26948), .D(n_28109
		), .Z(n_296183952));
	notech_ao4 i_130936993(.A(n_33512435), .B(n_28005), .C(n_33312433), .D(n_29038
		), .Z(n_296383954));
	notech_and4 i_131936984(.A(n_296183952), .B(n_296383954), .C(n_296083951
		), .D(n_256483555), .Z(n_296583956));
	notech_ao4 i_130536997(.A(n_388560287), .B(n_56064), .C(n_33012430), .D(n_28991
		), .Z(n_296683957));
	notech_ao4 i_130336999(.A(n_55869), .B(n_57574), .C(n_55860), .D(n_29254
		), .Z(n_296883959));
	notech_and4 i_130736995(.A(n_296883959), .B(n_296683957), .C(n_255683547
		), .D(n_255983550), .Z(n_297083961));
	notech_ao4 i_130037002(.A(n_5743), .B(n_55849), .C(n_55838), .D(n_29171)
		, .Z(n_297183962));
	notech_ao4 i_129937003(.A(n_55909), .B(n_308815164), .C(n_55886), .D(nbus_11295
		[12]), .Z(n_297383964));
	notech_and3 i_130237000(.A(n_297183962), .B(n_297383964), .C(n_255383544
		), .Z(n_297483965));
	notech_nao3 i_129837004(.A(n_60095), .B(instrc[121]), .C(n_101413114), .Z
		(n_297683967));
	notech_ao4 i_129437008(.A(n_17012270), .B(n_29011), .C(n_55909), .D(n_297683967
		), .Z(n_297783968));
	notech_ao4 i_129237010(.A(n_26949), .B(n_28100), .C(n_3886), .D(n_28092)
		, .Z(n_297983970));
	notech_and4 i_129637006(.A(n_297983970), .B(n_297783968), .C(n_254983540
		), .D(n_254683537), .Z(n_298183972));
	notech_ao4 i_128937013(.A(n_33412434), .B(n_29181), .C(n_26948), .D(n_28108
		), .Z(n_298283973));
	notech_ao4 i_128837014(.A(n_33512435), .B(n_28004), .C(n_33312433), .D(n_29037
		), .Z(n_298483975));
	notech_and4 i_129737005(.A(n_298283973), .B(n_298483975), .C(n_298183972
		), .D(n_254383534), .Z(n_298683977));
	notech_ao4 i_128437018(.A(n_388560287), .B(n_55983), .C(n_33012430), .D(n_28990
		), .Z(n_298783978));
	notech_ao4 i_128237020(.A(n_55869), .B(\nbus_11307[3] ), .C(n_55860), .D
		(n_29253), .Z(n_298983980));
	notech_and4 i_128637016(.A(n_298983980), .B(n_298783978), .C(n_253583526
		), .D(n_253883529), .Z(n_299183982));
	notech_ao4 i_127937023(.A(n_60022), .B(n_55849), .C(n_55838), .D(n_29170
		), .Z(n_299283983));
	notech_ao4 i_127837024(.A(n_55909), .B(n_308815164), .C(n_55886), .D(nbus_11295
		[11]), .Z(n_299483985));
	notech_and3 i_128137021(.A(n_299283983), .B(n_299483985), .C(n_253283523
		), .Z(n_299583986));
	notech_ao4 i_125537047(.A(n_60841), .B(n_28050), .C(n_57940), .D(n_58009
		), .Z(n_299783988));
	notech_ao4 i_125137051(.A(n_8812188), .B(n_29737), .C(n_55909), .D(n_246983460
		), .Z(n_299883989));
	notech_ao4 i_124937053(.A(n_3886), .B(n_28090), .C(n_3887), .D(n_29053),
		 .Z(n_300083991));
	notech_and4 i_125337049(.A(n_300083991), .B(n_299883989), .C(n_252383514
		), .D(n_252683517), .Z(n_300283993));
	notech_ao4 i_124637056(.A(n_26948), .B(n_28106), .C(n_19312293), .D(n_28114
		), .Z(n_300383994));
	notech_ao4 i_124437058(.A(n_33312433), .B(n_29036), .C(n_54512645), .D(n_56136
		), .Z(n_300583996));
	notech_and4 i_124837054(.A(n_300583996), .B(n_252083511), .C(n_300383994
		), .D(n_251783508), .Z(n_300783998));
	notech_ao4 i_124037062(.A(n_388560287), .B(n_56010), .C(n_33012430), .D(n_28986
		), .Z(n_300984000));
	notech_ao4 i_123837064(.A(n_55869), .B(n_57542), .C(n_55860), .D(n_29251
		), .Z(n_301184002));
	notech_and4 i_124237060(.A(n_301184002), .B(n_300984000), .C(n_251183502
		), .D(n_251483505), .Z(n_301384004));
	notech_ao4 i_123537067(.A(n_60024), .B(n_55849), .C(n_55838), .D(n_29168
		), .Z(n_301484005));
	notech_ao4 i_123437068(.A(n_54912649), .B(n_101413114), .C(n_55886), .D(nbus_11295
		[9]), .Z(n_301684007));
	notech_and4 i_124337059(.A(n_301484005), .B(n_301684007), .C(n_301384004
		), .D(n_250883499), .Z(n_301884009));
	notech_ao4 i_123037072(.A(n_8812188), .B(n_29735), .C(n_55909), .D(n_246683457
		), .Z(n_301984010));
	notech_ao4 i_122837074(.A(n_3886), .B(n_28089), .C(n_55800), .D(n_29052)
		, .Z(n_302184012));
	notech_and4 i_123237070(.A(n_302184012), .B(n_301984010), .C(n_250183492
		), .D(n_250483495), .Z(n_302384014));
	notech_ao4 i_122537077(.A(n_26948), .B(n_28105), .C(n_19312293), .D(n_28113
		), .Z(n_302484015));
	notech_ao4 i_122337079(.A(n_33312433), .B(n_29035), .C(n_54512645), .D(n_56118
		), .Z(n_302684017));
	notech_and4 i_122737075(.A(n_302684017), .B(n_249883489), .C(n_302484015
		), .D(n_249583486), .Z(n_302884019));
	notech_ao4 i_121937083(.A(n_388560287), .B(n_56028), .C(n_33012430), .D(n_28985
		), .Z(n_303084021));
	notech_ao4 i_121737085(.A(n_55869), .B(n_59742), .C(n_55860), .D(n_29250
		), .Z(n_303284023));
	notech_and4 i_122137081(.A(n_303284023), .B(n_303084021), .C(n_248983480
		), .D(n_249283483), .Z(n_303484025));
	notech_ao4 i_121437088(.A(n_56046), .B(n_55849), .C(n_55838), .D(n_29167
		), .Z(n_303584026));
	notech_ao4 i_121337089(.A(n_55909), .B(n_101413114), .C(n_55886), .D(nbus_11295
		[8]), .Z(n_303784028));
	notech_and4 i_122237080(.A(n_303584026), .B(n_303784028), .C(n_303484025
		), .D(n_248683477), .Z(n_303984030));
	notech_ao4 i_151335088(.A(n_59419), .B(n_305047803), .C(n_25615), .D(n_306884059
		), .Z(n_304084031));
	notech_nand2 i_33035151(.A(n_59153), .B(n_308484075), .Z(n_304184032));
	notech_or2 i_1535077(.A(n_276483755), .B(nbus_11295[15]), .Z(n_304284033
		));
	notech_and2 i_5035060(.A(n_304984040), .B(n_304484035), .Z(n_304384034)
		);
	notech_or4 i_4535065(.A(n_32259), .B(n_59419), .C(n_62870), .D(n_62892),
		 .Z(n_304484035));
	notech_or4 i_6735043(.A(n_58220), .B(n_59424), .C(n_60252), .D(n_308784078
		), .Z(n_304584036));
	notech_or4 i_7735033(.A(n_61156), .B(n_3790), .C(n_32476), .D(n_32567), 
		.Z(n_304684037));
	notech_and3 i_10135009(.A(n_32656), .B(n_304084031), .C(n_304884039), .Z
		(n_304784038));
	notech_or4 i_7035040(.A(n_2875), .B(n_28081), .C(n_32443), .D(n_59429), 
		.Z(n_304884039));
	notech_or4 i_10435006(.A(n_32259), .B(n_32747), .C(n_32730), .D(n_59429)
		, .Z(n_304984040));
	notech_ao4 i_11234998(.A(n_59451), .B(n_330763524), .C(n_1897), .D(n_60252
		), .Z(n_306084051));
	notech_and2 i_11134999(.A(n_318563452), .B(n_305987333), .Z(n_306484055)
		);
	notech_or4 i_111234023(.A(n_62856), .B(n_61117), .C(n_27857), .D(n_62824
		), .Z(n_306684057));
	notech_xor2 i_15734954(.A(n_60935), .B(n_60910), .Z(n_306884059));
	notech_and3 i_17494(.A(calc_sz[1]), .B(n_56970), .C(n_304184032), .Z(n_307084061
		));
	notech_and2 i_37483(.A(n_309184082), .B(n_304684037), .Z(n_307184062));
	notech_and3 i_35991(.A(n_304584036), .B(n_304284033), .C(n_57948), .Z(n_307384064
		));
	notech_or4 i_10635004(.A(n_32581), .B(n_19057), .C(n_60294), .D(n_18964)
		, .Z(n_307484065));
	notech_nao3 i_35969(.A(n_19093), .B(n_60372), .C(n_23755), .Z(n_307584066
		));
	notech_or4 i_35966(.A(fsm[2]), .B(n_61167), .C(n_61156), .D(n_2647), .Z(n_307684067
		));
	notech_or2 i_35812(.A(n_55773), .B(n_19101), .Z(n_307884069));
	notech_or4 i_35806(.A(n_2875), .B(n_59478), .C(n_32443), .D(n_330763524)
		, .Z(n_307984070));
	notech_or2 i_35805(.A(n_57533), .B(n_19101), .Z(n_308084071));
	notech_mux2 i_206033093(.S(n_60294), .A(n_26963), .B(n_306484055), .Z(n_308484075
		));
	notech_or4 i_205933094(.A(n_32580), .B(n_32559), .C(n_32567), .D(n_61131
		), .Z(n_308584076));
	notech_nao3 i_7835032(.A(n_26964), .B(n_60252), .C(n_32581), .Z(n_308684077
		));
	notech_mux2 i_735083(.S(n_32384), .A(n_59726), .B(n_57671), .Z(n_308784078
		));
	notech_ao4 i_203733116(.A(n_1878), .B(n_27069), .C(n_32579), .D(n_319991624
		), .Z(n_309184082));
	notech_nao3 i_5927(.A(n_60113), .B(n_60294), .C(n_311984110), .Z(n_309384084
		));
	notech_or2 i_24732527(.A(n_1869), .B(cond_1), .Z(n_309784088));
	notech_or4 i_25132523(.A(n_2875), .B(n_59478), .C(n_32443), .D(n_60894),
		 .Z(n_309884089));
	notech_and4 i_49292(.A(n_325884249), .B(n_313884129), .C(n_304784038), .D
		(n_57966), .Z(n_310084091));
	notech_and3 i_27032508(.A(n_32434), .B(n_2419), .C(n_53745), .Z(n_310384094
		));
	notech_and2 i_34132452(.A(n_326684257), .B(n_313484125), .Z(n_310584096)
		);
	notech_and4 i_34232451(.A(n_58697), .B(n_27056), .C(n_312984120), .D(n_57406
		), .Z(n_310784098));
	notech_nand2 i_33032460(.A(n_23627), .B(n_311284103), .Z(n_310884099));
	notech_ao4 i_33132459(.A(n_60283), .B(n_26985), .C(n_2896), .D(n_26757),
		 .Z(n_310984100));
	notech_and2 i_33332458(.A(n_28533), .B(n_322284213), .Z(n_311084101));
	notech_nor2 i_33532457(.A(n_320584196), .B(n_322084211), .Z(n_311184102)
		);
	notech_or4 i_63332201(.A(n_2884), .B(n_57514), .C(n_62850), .D(n_62824),
		 .Z(n_311284103));
	notech_and2 i_30132482(.A(n_311484105), .B(n_322184212), .Z(n_311384104)
		);
	notech_nao3 i_63532199(.A(n_32730), .B(n_27641), .C(n_62870), .Z(n_311484105
		));
	notech_or4 i_64032195(.A(n_4978711), .B(n_32643), .C(n_32655), .D(n_59429
		), .Z(n_311784108));
	notech_nand2 i_64332192(.A(n_23006), .B(n_26984), .Z(n_311884109));
	notech_and4 i_64432191(.A(n_4758689), .B(n_1893), .C(n_314984140), .D(n_304384034
		), .Z(n_311984110));
	notech_and2 i_64532190(.A(n_27988), .B(n_28533), .Z(n_312084111));
	notech_or4 i_64632189(.A(n_27925), .B(n_62870), .C(n_62892), .D(n_27084)
		, .Z(n_312184112));
	notech_ao4 i_11632625(.A(n_56941), .B(n_3695), .C(n_30910), .D(n_32298),
		 .Z(n_312284113));
	notech_ao3 i_32232465(.A(n_58573), .B(n_57076), .C(n_316484155), .Z(n_312384114
		));
	notech_and3 i_12032621(.A(n_58573), .B(n_57076), .C(n_312684117), .Z(n_312484115
		));
	notech_and4 i_32432464(.A(n_30905), .B(n_27035), .C(n_3826), .D(n_3827),
		 .Z(n_312584116));
	notech_or4 i_73232111(.A(n_340480905), .B(instrc[125]), .C(n_29632), .D(n_317284163
		), .Z(n_312684117));
	notech_nand2 i_53932288(.A(rep_en5), .B(n_27053), .Z(n_312984120));
	notech_or4 i_53832289(.A(n_19093), .B(n_59322), .C(n_19101), .D(n_26900)
		, .Z(n_313084121));
	notech_or4 i_53532292(.A(n_6258839), .B(n_57899), .C(n_26967), .D(n_26779
		), .Z(n_313184122));
	notech_or4 i_53632291(.A(n_5380), .B(n_27069), .C(n_32596), .D(n_32548),
		 .Z(n_313284123));
	notech_or4 i_53732290(.A(n_59322), .B(n_26900), .C(n_60372), .D(n_29656)
		, .Z(n_313384124));
	notech_ao4 i_36054(.A(n_61117), .B(n_310084091), .C(n_55632), .D(n_61131
		), .Z(n_313484125));
	notech_ao4 i_200336305(.A(n_57976), .B(n_28295), .C(n_60841), .D(n_28489
		), .Z(n_306960150));
	notech_or4 i_35659(.A(n_32643), .B(n_2875), .C(n_2877), .D(n_59429), .Z(n_313784128
		));
	notech_and4 i_35953(.A(n_25386), .B(n_125761540), .C(n_309884089), .D(n_313984130
		), .Z(n_313884129));
	notech_or4 i_15132590(.A(n_252140539), .B(n_2888), .C(n_1864), .D(n_2877
		), .Z(n_313984130));
	notech_or2 i_63132203(.A(n_17779989), .B(n_311184102), .Z(n_314284133)
		);
	notech_nao3 i_62732207(.A(n_18559), .B(n_32272), .C(n_27500), .Z(n_314384134
		));
	notech_nand3 i_62832206(.A(n_60113), .B(n_60294), .C(n_310884099), .Z(n_314484135
		));
	notech_or4 i_62532209(.A(n_32263), .B(n_27501), .C(n_18559), .D(n_32729)
		, .Z(n_314584136));
	notech_nao3 i_62632208(.A(n_17189930), .B(n_27052), .C(n_6258839), .Z(n_314684137
		));
	notech_nor2 i_65632179(.A(writeio_ack), .B(readio_ack), .Z(n_314784138)
		);
	notech_or4 i_19832572(.A(n_60964), .B(n_60953), .C(n_62850), .D(n_312084111
		), .Z(n_314984140));
	notech_ao3 i_72832115(.A(instrc[98]), .B(n_26760), .C(n_345780958), .Z(n_315684147
		));
	notech_ao3 i_72532118(.A(instrc[104]), .B(instrc[107]), .C(n_346180962),
		 .Z(n_315984150));
	notech_and4 i_71632123(.A(n_29635), .B(instrc[102]), .C(instrc[103]), .D
		(n_30350), .Z(n_316084151));
	notech_or4 i_71732122(.A(n_57078), .B(n_57051), .C(n_57033), .D(n_26971)
		, .Z(n_316184152));
	notech_nao3 i_71832121(.A(n_30357), .B(n_26847), .C(n_30969), .Z(n_316284153
		));
	notech_or4 i_29671(.A(n_59322), .B(n_30306), .C(n_26900), .D(n_29642), .Z
		(n_316384154));
	notech_and4 i_73132112(.A(n_62868), .B(n_58632), .C(n_30931), .D(n_30322
		), .Z(n_316484155));
	notech_nao3 i_129231592(.A(n_316284153), .B(n_316184152), .C(n_316084151
		), .Z(n_316984160));
	notech_nand2 i_131831567(.A(n_62868), .B(n_58632), .Z(n_317284163));
	notech_ao4 i_128931595(.A(n_312584116), .B(n_312484115), .C(n_312284113)
		, .D(n_312384114), .Z(n_317784168));
	notech_ao4 i_128631598(.A(n_32339), .B(n_345980960), .C(n_346080961), .D
		(n_316384154), .Z(n_318084171));
	notech_ao4 i_128531599(.A(n_56640), .B(n_3829), .C(n_345680957), .D(n_26968
		), .Z(n_318284173));
	notech_nao3 i_128831596(.A(n_318084171), .B(n_318284173), .C(n_315684147
		), .Z(n_318384174));
	notech_and4 i_110531767(.A(n_314384134), .B(n_314584136), .C(n_314484135
		), .D(n_314684137), .Z(n_319084181));
	notech_or4 i_119931681(.A(opb[1]), .B(opb[2]), .C(opb[3]), .D(opb[0]), .Z
		(n_319384184));
	notech_or4 i_119631684(.A(opb[6]), .B(opb[7]), .C(opb[4]), .D(opb[5]), .Z
		(n_319684187));
	notech_or4 i_119131688(.A(opb[10]), .B(opb[11]), .C(opb[8]), .D(opb[9]),
		 .Z(n_320084191));
	notech_or4 i_118831691(.A(opb[15]), .B(opb[16]), .C(opb[12]), .D(opb[14]
		), .Z(n_320384194));
	notech_or4 i_120231679(.A(n_320384194), .B(n_320084191), .C(n_319684187)
		, .D(n_319384184), .Z(n_320584196));
	notech_or4 i_118331696(.A(opb[19]), .B(opb[20]), .C(opb[17]), .D(opb[18]
		), .Z(n_320884199));
	notech_or4 i_118031699(.A(opb[23]), .B(opb[24]), .C(opb[21]), .D(opb[22]
		), .Z(n_321184202));
	notech_or4 i_117631703(.A(opb[28]), .B(opb[29]), .C(opb[25]), .D(opb[26]
		), .Z(n_321584206));
	notech_or4 i_117231706(.A(opb[27]), .B(opb[30]), .C(opb[13]), .D(opb[31]
		), .Z(n_321884209));
	notech_or4 i_118531694(.A(n_321884209), .B(n_321584206), .C(n_321184202)
		, .D(n_320884199), .Z(n_322084211));
	notech_ao4 i_27132507(.A(n_18559), .B(n_1868), .C(n_32729), .D(n_27641),
		 .Z(n_322184212));
	notech_ao4 i_120431677(.A(n_27925), .B(n_1868), .C(n_27501), .D(n_311384104
		), .Z(n_322284213));
	notech_ao4 i_110131771(.A(n_308012096), .B(n_311084101), .C(n_32476), .D
		(n_310984100), .Z(n_322384214));
	notech_and3 i_109931773(.A(n_3912), .B(n_313084121), .C(n_17669978), .Z(n_322784218
		));
	notech_and3 i_34832737(.A(n_307184062), .B(n_57716), .C(n_107111189), .Z
		(n_322984220));
	notech_nand3 i_116631712(.A(n_27132), .B(n_27123), .C(n_32747), .Z(n_323084221
		));
	notech_ao4 i_116231716(.A(n_3777), .B(n_3698), .C(n_61117), .D(n_57912),
		 .Z(n_323384224));
	notech_and3 i_148932700(.A(n_318591638), .B(n_60136), .C(n_323384224), .Z
		(n_323584226));
	notech_and4 i_110031772(.A(n_320263469), .B(n_323584226), .C(n_322984220
		), .D(n_322784218), .Z(n_323884229));
	notech_and4 i_110731765(.A(n_322384214), .B(n_319084181), .C(n_323884229
		), .D(n_314284133), .Z(n_323984230));
	notech_and4 i_109131779(.A(n_187410086), .B(n_187310085), .C(n_309384084
		), .D(n_26860), .Z(n_324384234));
	notech_and4 i_109231778(.A(n_58664), .B(n_187610088), .C(n_57285), .D(n_324384234
		), .Z(n_324684237));
	notech_ao3 i_108631784(.A(n_3905), .B(n_27379), .C(n_27097), .Z(n_325184242
		));
	notech_and4 i_108731783(.A(n_59763), .B(n_58683), .C(n_60113), .D(n_325184242
		), .Z(n_325484245));
	notech_or4 i_22032550(.A(n_18981), .B(n_288827270), .C(n_18972), .D(n_27052
		), .Z(n_325684247));
	notech_ao4 i_106231807(.A(n_252140539), .B(n_2647), .C(n_59424), .D(n_58220
		), .Z(n_325884249));
	notech_or2 i_141132762(.A(n_6258839), .B(n_26779), .Z(n_326184252));
	notech_ao4 i_102931839(.A(n_319963466), .B(n_314663413), .C(n_32476), .D
		(n_57403), .Z(n_326584256));
	notech_and4 i_33932750(.A(n_326584256), .B(n_313284123), .C(n_313184122)
		, .D(n_313384124), .Z(n_326684257));
	notech_nao3 i_26732510(.A(n_57839), .B(n_61559), .C(n_6258839), .Z(n_326784258
		));
	notech_or2 i_159067432(.A(n_109982100), .B(n_83341448), .Z(n_327084261)
		);
	notech_or2 i_21867431(.A(n_110082101), .B(n_56205), .Z(n_327184262));
	notech_or2 i_20267430(.A(n_110182102), .B(n_56205), .Z(n_327284263));
	notech_or2 i_21467429(.A(n_110282103), .B(n_56205), .Z(n_327384264));
	notech_or2 i_19667428(.A(n_110382104), .B(n_56205), .Z(n_327484265));
	notech_or2 i_20367427(.A(n_110482105), .B(n_56205), .Z(n_327584266));
	notech_or2 i_20867426(.A(n_110582106), .B(n_56205), .Z(n_327684267));
	notech_or2 i_21167425(.A(n_110682107), .B(n_56205), .Z(n_327784268));
	notech_or2 i_19767424(.A(n_110782108), .B(n_56205), .Z(n_327884269));
	notech_or2 i_21267417(.A(n_110882109), .B(n_56205), .Z(n_327984270));
	notech_or4 i_33432866(.A(tcmp), .B(n_61131), .C(n_60252), .D(n_1881), .Z
		(n_58683));
	notech_or4 i_19242(.A(n_58220), .B(n_10157), .C(n_58009), .D(n_32323), .Z
		(n_328084271));
	notech_ao4 i_37599(.A(n_61117), .B(n_310384094), .C(n_32405), .D(n_32403
		), .Z(n_187310085));
	notech_ao4 i_200436304(.A(n_58009), .B(n_27864), .C(n_56463), .D(n_29718
		), .Z(n_306860149));
	notech_ao4 i_85753966(.A(n_60294), .B(n_26985), .C(n_328284273), .D(n_56566
		), .Z(n_328184272));
	notech_nor2 i_23753964(.A(n_179382794), .B(n_55191), .Z(n_328284273));
	notech_or4 i_53658(.A(n_141782418), .B(n_143582436), .C(n_143982440), .D
		(n_26893), .Z(\nbus_11350[0] ));
	notech_or4 i_51208(.A(n_145082451), .B(n_140682407), .C(n_26896), .D(n_26897
		), .Z(\nbus_11332[0] ));
	notech_and4 i_50955(.A(n_139782398), .B(n_146082461), .C(n_146882469), .D
		(n_145982460), .Z(\nbus_11331[0] ));
	notech_or2 i_21564469(.A(n_56205), .B(n_131282313), .Z(\nbus_11317[25] )
		);
	notech_or2 i_21764468(.A(n_56204), .B(n_131182312), .Z(\nbus_11317[26] )
		);
	notech_or2 i_21364467(.A(n_56199), .B(n_131082311), .Z(\nbus_11317[30] )
		);
	notech_or2 i_20164466(.A(n_130982310), .B(n_56199), .Z(\nbus_11317[31] )
		);
	notech_and4 i_1020991(.A(n_147482475), .B(n_147682477), .C(n_148182482),
		 .D(n_138482385), .Z(n_23788));
	notech_nand2 i_2027371(.A(n_148582486), .B(n_130582306), .Z(n_21765));
	notech_and4 i_3212949(.A(n_149182492), .B(n_149382494), .C(n_149082491),
		 .D(n_136782368), .Z(n_26103));
	notech_nand3 i_3112948(.A(n_150082501), .B(n_149982500), .C(n_149882499)
		, .Z(n_26098));
	notech_nand3 i_2712944(.A(n_150782508), .B(n_150682507), .C(n_150582506)
		, .Z(n_26078));
	notech_nand3 i_2612943(.A(n_151482515), .B(n_151382514), .C(n_151282513)
		, .Z(n_26073));
	notech_and2 i_200836300(.A(n_306660147), .B(n_306560146), .Z(n_306760148
		));
	notech_ao4 i_200636302(.A(n_56396), .B(n_28164), .C(n_56391), .D(n_28393
		), .Z(n_306660147));
	notech_ao4 i_172264449(.A(n_313784128), .B(n_60252), .C(n_148282483), .D
		(opc[31]), .Z(n_255640574));
	notech_or4 i_8064373(.A(fsm[2]), .B(n_61167), .C(n_61156), .D(n_313784128
		), .Z(n_247640494));
	notech_ao4 i_200736301(.A(n_59344), .B(n_28522), .C(n_56367), .D(n_28328
		), .Z(n_306560146));
	notech_and4 i_201636292(.A(n_306260143), .B(n_306160142), .C(n_305960140
		), .D(n_305860139), .Z(n_306460145));
	notech_ao4 i_201036298(.A(n_56452), .B(n_28263), .C(n_58020), .D(n_28457
		), .Z(n_306260143));
	notech_and4 i_3120884(.A(n_154182542), .B(n_154382544), .C(n_154082541),
		 .D(n_154782548), .Z(n_24262));
	notech_or4 i_3121012(.A(n_117868195), .B(n_152582526), .C(n_155182552), 
		.D(n_26903), .Z(n_23914));
	notech_and4 i_3121108(.A(n_155582556), .B(n_155782558), .C(n_156282563),
		 .D(n_152482525), .Z(n_19009));
	notech_and4 i_121174(.A(n_158182582), .B(n_158382584), .C(n_158882589), 
		.D(n_157582576), .Z(n_18480));
	notech_nand2 i_2918994(.A(n_170682707), .B(n_170182702), .Z(n_25656));
	notech_nand2 i_2018985(.A(n_171682717), .B(n_171182712), .Z(n_25602));
	notech_nand2 i_1918984(.A(n_172682727), .B(n_172182722), .Z(n_25596));
	notech_nand2 i_1818983(.A(n_173682737), .B(n_173182732), .Z(n_25590));
	notech_nand2 i_1718982(.A(n_174682747), .B(n_174182742), .Z(n_25584));
	notech_nand2 i_1618981(.A(n_175682757), .B(n_175182752), .Z(n_25578));
	notech_nand2 i_1518980(.A(n_176682767), .B(n_176182762), .Z(n_25572));
	notech_nand2 i_1418979(.A(n_177682777), .B(n_177182772), .Z(n_25566));
	notech_nand2 i_1318978(.A(n_178682787), .B(n_178182782), .Z(n_25560));
	notech_ao4 i_22635137(.A(n_60294), .B(n_26964), .C(n_32553), .D(n_18989)
		, .Z(n_58791));
	notech_ao4 i_22835138(.A(n_32559), .B(n_26963), .C(n_32434), .D(n_60252)
		, .Z(n_58789));
	notech_ao4 i_22935139(.A(n_32559), .B(n_26580), .C(n_32432), .D(n_60252)
		, .Z(n_58788));
	notech_ao4 i_201136297(.A(n_56443), .B(n_28229), .C(n_56432), .D(n_28196
		), .Z(n_306160142));
	notech_ao4 i_201336295(.A(n_56908), .B(n_29719), .C(n_56423), .D(n_28361
		), .Z(n_305960140));
	notech_ao4 i_26635140(.A(n_28533), .B(n_190710119), .C(n_27063), .D(n_57440
		), .Z(n_58751));
	notech_ao4 i_26735141(.A(n_58786), .B(n_60246), .C(n_27063), .D(n_306084051
		), .Z(n_58750));
	notech_or2 i_20053965(.A(n_179582796), .B(n_56199), .Z(n_328384274));
	notech_nao3 i_22153938(.A(n_60113), .B(n_60294), .C(n_58072), .Z(n_328484275
		));
	notech_ao4 i_201436294(.A(n_56414), .B(n_28425), .C(n_56405), .D(n_28566
		), .Z(n_305860139));
	notech_ao4 i_214936159(.A(n_57976), .B(n_28308), .C(n_60841), .D(n_28501
		), .Z(n_305560136));
	notech_ao4 i_215036158(.A(n_58009), .B(n_27876), .C(n_56463), .D(n_29712
		), .Z(n_305460135));
	notech_and2 i_215436154(.A(n_305260133), .B(n_305160132), .Z(n_305360134
		));
	notech_ao4 i_215236156(.A(n_56400), .B(n_28176), .C(n_56391), .D(n_28405
		), .Z(n_305260133));
	notech_ao4 i_215336155(.A(n_59344), .B(n_28539), .C(n_56371), .D(n_28341
		), .Z(n_305160132));
	notech_and4 i_1720774(.A(n_230683297), .B(n_230883299), .C(n_231383304),
		 .D(n_230583296), .Z(n_24526));
	notech_and4 i_1720870(.A(n_231483305), .B(n_231683307), .C(n_232083311),
		 .D(n_229683287), .Z(n_24178));
	notech_and4 i_1720998(.A(n_232183312), .B(n_232383314), .C(n_232883319),
		 .D(n_228883279), .Z(n_23830));
	notech_and4 i_1721190(.A(n_232983320), .B(n_233183322), .C(n_233683327),
		 .D(n_227983270), .Z(n_18576));
	notech_and4 i_1721638(.A(n_233783328), .B(n_233983330), .C(n_234483335),
		 .D(n_227083261), .Z(n_17876));
	notech_nand2 i_96144582(.A(n_319591628), .B(n_319491629), .Z(n_58088));
	notech_and4 i_3220789(.A(n_240183392), .B(n_240383394), .C(n_240883399),
		 .D(n_240083391), .Z(n_24616));
	notech_nand3 i_3221653(.A(n_241083401), .B(n_240983400), .C(n_241483405)
		, .Z(n_17966));
	notech_and4 i_3221877(.A(n_241583406), .B(n_241783408), .C(n_242183412),
		 .D(n_238483375), .Z(n_20804));
	notech_or4 i_3221941(.A(n_237083361), .B(n_215876097), .C(n_242883419), 
		.D(n_26940), .Z(n_17618));
	notech_or4 i_3217621(.A(n_215876097), .B(n_236283353), .C(n_26944), .D(n_26943
		), .Z(n_16892));
	notech_and2 i_4144453(.A(n_306221226), .B(n_235983350), .Z(n_303721201)
		);
	notech_nand2 i_917182(.A(n_246483455), .B(n_245983450), .Z(n_15061));
	notech_and2 i_171935136(.A(n_25613), .B(n_55632), .Z(n_57367));
	notech_and4 i_216236146(.A(n_304860129), .B(n_304760128), .C(n_304560126
		), .D(n_304460125), .Z(n_305060131));
	notech_ao4 i_215636152(.A(n_56452), .B(n_28275), .C(n_58024), .D(n_28469
		), .Z(n_304860129));
	notech_ao4 i_215736151(.A(n_56443), .B(n_28243), .C(n_56432), .D(n_28208
		), .Z(n_304760128));
	notech_ao4 i_36635135(.A(n_32656), .B(n_60252), .C(n_27052), .D(n_308684077
		), .Z(n_58651));
	notech_ao4 i_215936149(.A(n_56908), .B(n_29713), .C(n_56423), .D(n_28373
		), .Z(n_304560126));
	notech_ao4 i_216036148(.A(n_56414), .B(n_28437), .C(n_56405), .D(n_28579
		), .Z(n_304460125));
	notech_or4 i_27138258(.A(fsm[2]), .B(n_61167), .C(n_3792), .D(n_60294), 
		.Z(n_58746));
	notech_nand2 i_1916232(.A(n_278283773), .B(n_277783768), .Z(n_19214));
	notech_or4 i_1616229(.A(n_279983790), .B(n_279583786), .C(n_279083781), 
		.D(n_278683777), .Z(n_19196));
	notech_and4 i_1516228(.A(n_280783798), .B(n_280683797), .C(n_280583796),
		 .D(n_281883809), .Z(n_19190));
	notech_and4 i_1416227(.A(n_282483815), .B(n_282383814), .C(n_282283813),
		 .D(n_283483825), .Z(n_19184));
	notech_and4 i_1216225(.A(n_284083831), .B(n_283983830), .C(n_285083841),
		 .D(n_283883829), .Z(n_19172));
	notech_and4 i_1116224(.A(n_285683847), .B(n_285583846), .C(n_285483845),
		 .D(n_286683857), .Z(n_19166));
	notech_and4 i_1016223(.A(n_287283863), .B(n_287183862), .C(n_287083861),
		 .D(n_288283873), .Z(n_19160));
	notech_and4 i_916222(.A(n_288883879), .B(n_288783878), .C(n_289883889), 
		.D(n_288683877), .Z(n_19154));
	notech_nand3 i_816221(.A(n_291583906), .B(n_290783898), .C(n_291183902),
		 .Z(n_19148));
	notech_nand3 i_716220(.A(n_292183912), .B(n_293583926), .C(n_292583916),
		 .Z(n_19142));
	notech_nand3 i_616219(.A(n_294083931), .B(n_295483945), .C(n_294483935),
		 .Z(n_19136));
	notech_nand3 i_516218(.A(n_297083961), .B(n_296583956), .C(n_297483965),
		 .Z(n_19130));
	notech_nand3 i_416217(.A(n_299183982), .B(n_298683977), .C(n_299583986),
		 .Z(n_19124));
	notech_nand3 i_216215(.A(n_300783998), .B(n_300283993), .C(n_301884009),
		 .Z(n_19112));
	notech_nand3 i_116214(.A(n_302884019), .B(n_302384014), .C(n_303984030),
		 .Z(n_19106));
	notech_and3 i_45238227(.A(n_273383724), .B(n_34012440), .C(n_54512645), 
		.Z(n_309615172));
	notech_or2 i_45338226(.A(n_247283463), .B(n_56109), .Z(n_309515171));
	notech_and3 i_938219(.A(n_56443), .B(n_247683467), .C(n_246583456), .Z(n_308815164
		));
	notech_or4 i_3438200(.A(instrc[122]), .B(instrc[121]), .C(n_26735), .D(n_29022
		), .Z(n_306915145));
	notech_and2 i_39838234(.A(n_54512645), .B(n_3892), .Z(n_310315179));
	notech_and4 i_52155(.A(n_340991464), .B(n_340891465), .C(n_306684057), .D
		(n_340791466), .Z(\nbus_11337[16] ));
	notech_nand2 i_54849(.A(n_311187385), .B(n_109682097), .Z(n_23569));
	notech_ao4 i_133335148(.A(n_27068), .B(n_27069), .C(n_308584076), .D(n_26999
		), .Z(n_57716));
	notech_or4 i_21344(.A(n_2884), .B(n_62824), .C(n_60910), .D(n_60246), .Z
		(n_38609));
	notech_nao3 i_79735118(.A(n_2825), .B(n_27132), .C(n_27994), .Z(n_58220)
		);
	notech_or4 i_164535117(.A(n_59460), .B(n_60935), .C(n_60910), .D(n_60246
		), .Z(n_57440));
	notech_or4 i_38066(.A(fsm[2]), .B(n_61167), .C(n_61156), .D(n_304384034)
		, .Z(n_310447752));
	notech_or4 i_38070(.A(n_60868), .B(n_59478), .C(n_60246), .D(n_27573), .Z
		(n_310347753));
	notech_or4 i_38071(.A(n_3790), .B(n_32562), .C(n_3792), .D(n_3803), .Z(n_310247754
		));
	notech_or4 i_55515(.A(n_315984150), .B(n_316984160), .C(n_318384174), .D
		(n_26974), .Z(\nbus_11374[0] ));
	notech_nao3 i_52472(.A(n_325484245), .B(n_324684237), .C(n_26978), .Z(\nbus_11340[0] 
		));
	notech_or2 i_3429(.A(n_4958709), .B(n_323084221), .Z(n_60055));
	notech_or4 i_48800(.A(n_60894), .B(n_61110), .C(n_2839), .D(n_2888), .Z(n_60123
		));
	notech_or4 i_32632915(.A(n_18964), .B(n_60094), .C(n_6258839), .D(n_17189930
		), .Z(n_58691));
	notech_or4 i_5935(.A(n_2884), .B(n_61103), .C(n_60935), .D(n_60910), .Z(n_53748
		));
	notech_nand2 i_5940(.A(nZF), .B(n_311884109), .Z(n_53745));
	notech_and2 i_113732897(.A(n_311784108), .B(n_60055), .Z(n_57912));
	notech_nao3 i_80232865(.A(n_60113), .B(n_60294), .C(n_57308), .Z(n_58215
		));
	notech_or4 i_35132864(.A(n_19072), .B(n_32476), .C(n_32569), .D(n_314784138
		), .Z(n_58666));
	notech_ao4 i_19613(.A(n_310784098), .B(n_326784258), .C(n_310584096), .D
		(n_29793), .Z(\nbus_11313[0] ));
	notech_and4 i_27732819(.A(n_26702), .B(n_26643), .C(n_59708), .D(n_32452
		), .Z(n_58740));
	notech_nao3 i_178332818(.A(reps[2]), .B(n_27922), .C(n_60868), .Z(n_57308
		));
	notech_nand2 i_169832763(.A(n_312184112), .B(n_58691), .Z(n_14570));
	notech_and2 i_108332752(.A(n_313784128), .B(n_60074), .Z(n_57966));
	notech_ao4 i_37585(.A(n_61103), .B(n_16879899), .C(n_26992), .D(n_29771)
		, .Z(n_187610088));
	notech_and2 i_37596(.A(n_53748), .B(n_60123), .Z(n_187410086));
	notech_and2 i_20832562(.A(n_58740), .B(n_309784088), .Z(n_16879899));
	notech_nao3 i_13438109(.A(n_295960040), .B(imm[2]), .C(n_55909), .Z(n_299260073
		));
	notech_nand2 i_13738106(.A(n_19512295), .B(read_data[10]), .Z(n_298960070
		));
	notech_nao3 i_14038103(.A(nbus_160[2]), .B(n_26782), .C(n_52112621), .Z(n_298660067
		));
	notech_or2 i_14338100(.A(n_33512435), .B(n_28003), .Z(n_298360064));
	notech_or2 i_14638097(.A(n_55809), .B(nbus_11295[2]), .Z(n_298060061));
	notech_or4 i_14938094(.A(n_58086), .B(n_59478), .C(n_57132), .D(n_59259)
		, .Z(n_297760058));
	notech_nand2 i_15238091(.A(resb_shiftbox[2]), .B(n_27003), .Z(n_297460055
		));
	notech_or4 i_63037636(.A(n_60868), .B(n_27925), .C(n_32643), .D(n_60252)
		, .Z(n_296860049));
	notech_ao4 i_62937637(.A(n_32656), .B(n_60252), .C(n_308760168), .D(n_27052
		), .Z(n_296760048));
	notech_and3 i_5638186(.A(n_25629), .B(n_58220), .C(n_26965), .Z(n_296160042
		));
	notech_nao3 i_25937984(.A(n_309160172), .B(n_27541), .C(mask8b[1]), .Z(n_296060041
		));
	notech_nand3 i_23838005(.A(n_56427), .B(n_56414), .C(n_56405), .Z(n_295960040
		));
	notech_and2 i_5138189(.A(n_310060181), .B(n_56371), .Z(n_295860039));
	notech_nand2 i_1738217(.A(n_56432), .B(n_56908), .Z(n_295760038));
	notech_ao4 i_193439465(.A(n_56666), .B(n_28233), .C(n_56653), .D(n_28200
		), .Z(n_295460035));
	notech_ao4 i_193539464(.A(n_56916), .B(n_29720), .C(n_56640), .D(n_28267
		), .Z(n_295360034));
	notech_and2 i_193939460(.A(n_295160032), .B(n_295060031), .Z(n_295260033
		));
	notech_ao4 i_193739462(.A(n_28299), .B(n_56532), .C(n_56513), .D(n_56163
		), .Z(n_295160032));
	notech_ao4 i_193839461(.A(n_56502), .B(n_28365), .C(n_56489), .D(n_28333
		), .Z(n_295060031));
	notech_and4 i_194739452(.A(n_294760028), .B(n_294660027), .C(n_294460025
		), .D(n_294360024), .Z(n_294960030));
	notech_ao4 i_194139458(.A(n_56627), .B(n_28429), .C(n_56614), .D(n_28397
		), .Z(n_294760028));
	notech_ao4 i_194239457(.A(n_56601), .B(n_28461), .C(n_56592), .D(n_28168
		), .Z(n_294660027));
	notech_ao4 i_194439455(.A(n_56579), .B(n_28493), .C(n_56566), .D(n_28528
		), .Z(n_294460025));
	notech_ao4 i_194539454(.A(n_56553), .B(n_27868), .C(n_56542), .D(n_28571
		), .Z(n_294360024));
	notech_nand2 i_28542(.A(n_62798), .B(opc_10[10]), .Z(n_31433));
	notech_or4 i_28564(.A(n_60964), .B(n_60953), .C(n_62850), .D(n_56145), .Z
		(n_31411));
	notech_and3 i_131743246(.A(n_281259893), .B(n_292360004), .C(n_278059861
		), .Z(n_292560006));
	notech_ao4 i_131643247(.A(n_29717), .B(n_151761800), .C(n_60022), .D(n_58004
		), .Z(n_292360004));
	notech_ao4 i_131843245(.A(n_58003), .B(n_29728), .C(n_58409), .D(n_59223
		), .Z(n_292160002));
	notech_ao4 i_132043244(.A(n_59095), .B(n_28092), .C(n_60113), .D(n_27120
		), .Z(n_292060001));
	notech_and4 i_133243235(.A(n_291759998), .B(n_291659997), .C(n_291459995
		), .D(n_291359994), .Z(n_291960000));
	notech_ao4 i_132443241(.A(n_57889), .B(n_57563), .C(n_57890), .D(n_55983
		), .Z(n_291759998));
	notech_ao4 i_132543240(.A(n_308721251), .B(n_306091763), .C(n_306970080)
		, .D(n_24583), .Z(n_291659997));
	notech_ao4 i_132943238(.A(n_306870079), .B(n_57841), .C(n_306770078), .D
		(n_151961802), .Z(n_291459995));
	notech_ao4 i_133043237(.A(n_306570076), .B(n_26774), .C(n_306670077), .D
		(n_281363080), .Z(n_291359994));
	notech_and3 i_133543232(.A(n_281259893), .B(n_290959990), .C(n_279559876
		), .Z(n_291159992));
	notech_ao4 i_133443233(.A(n_151761800), .B(n_29716), .C(n_60020), .D(n_58004
		), .Z(n_290959990));
	notech_ao4 i_133643231(.A(n_58003), .B(n_29651), .C(n_58409), .D(n_59205
		), .Z(n_290759988));
	notech_ao4 i_133743230(.A(n_59095), .B(n_28094), .C(n_60113), .D(n_27122
		), .Z(n_290659987));
	notech_and4 i_134643221(.A(n_290359984), .B(n_290259983), .C(n_290059981
		), .D(n_289959980), .Z(n_290559986));
	notech_ao4 i_134043227(.A(\nbus_11307[5] ), .B(n_57889), .C(n_57890), .D
		(n_56073), .Z(n_290359984));
	notech_ao4 i_134143226(.A(n_308621250), .B(n_306091763), .C(n_282266351)
		, .D(n_24583), .Z(n_290259983));
	notech_ao4 i_134343224(.A(n_57841), .B(n_282166350), .C(n_282066349), .D
		(n_151961802), .Z(n_290059981));
	notech_ao4 i_134443223(.A(n_281966348), .B(n_26774), .C(n_281866347), .D
		(n_281363080), .Z(n_289959980));
	notech_and4 i_135243215(.A(n_281259893), .B(n_289659977), .C(n_289459975
		), .D(n_289359974), .Z(n_289859979));
	notech_ao4 i_134743220(.A(n_151861801), .B(n_29715), .C(n_151761800), .D
		(n_29714), .Z(n_289659977));
	notech_ao4 i_134943218(.A(n_59095), .B(n_28095), .C(n_58409), .D(n_27989
		), .Z(n_289459975));
	notech_ao4 i_135043217(.A(n_3874), .B(n_58004), .C(n_60113), .D(n_27124)
		, .Z(n_289359974));
	notech_and4 i_135943208(.A(n_289059971), .B(n_288959970), .C(n_288759968
		), .D(n_288659967), .Z(n_289259973));
	notech_ao4 i_135343214(.A(n_3868), .B(n_306091763), .C(n_151961802), .D(n_26802
		), .Z(n_289059971));
	notech_ao4 i_135443213(.A(n_92619108), .B(n_24583), .C(n_92019102), .D(n_57841
		), .Z(n_288959970));
	notech_ao4 i_135643211(.A(n_92519107), .B(n_281463081), .C(n_276459845),
		 .D(n_29723), .Z(n_288759968));
	notech_ao4 i_135743210(.A(n_276359844), .B(n_56082), .C(n_57592), .D(n_276259843
		), .Z(n_288659967));
	notech_nand3 i_161742970(.A(n_288259963), .B(n_288459965), .C(n_282959910
		), .Z(n_288559966));
	notech_ao4 i_161442973(.A(n_307091753), .B(n_27641), .C(n_55726), .D(n_28095
		), .Z(n_288459965));
	notech_ao4 i_161542972(.A(n_343270443), .B(n_92019102), .C(n_3873), .D(eval_flag
		), .Z(n_288259963));
	notech_ao4 i_161842969(.A(n_57592), .B(n_276859849), .C(n_276759848), .D
		(n_56508), .Z(n_287959960));
	notech_ao4 i_162542962(.A(n_26789), .B(n_26606), .C(n_304591778), .D(n_56508
		), .Z(n_287859959));
	notech_ao4 i_162442963(.A(n_27746), .B(n_3874), .C(n_92519107), .D(n_27757
		), .Z(n_287659957));
	notech_nand3 i_162142966(.A(n_283459915), .B(n_283359914), .C(n_283559916
		), .Z(n_287559956));
	notech_ao4 i_208142509(.A(n_28229), .B(n_56666), .C(n_28196), .D(n_56653
		), .Z(n_286959950));
	notech_ao4 i_208242508(.A(n_56916), .B(n_29719), .C(n_28263), .D(n_56640
		), .Z(n_286859949));
	notech_and2 i_208642504(.A(n_286659947), .B(n_286559946), .Z(n_286759948
		));
	notech_ao4 i_208442506(.A(n_28295), .B(n_56532), .C(n_56502), .D(n_28361
		), .Z(n_286659947));
	notech_ao4 i_208542505(.A(n_56489), .B(n_28328), .C(n_28425), .D(n_56627
		), .Z(n_286559946));
	notech_and4 i_209442496(.A(n_286259943), .B(n_286159942), .C(n_285959940
		), .D(n_285859939), .Z(n_286459945));
	notech_ao4 i_208842502(.A(n_56614), .B(n_28393), .C(n_56605), .D(n_28457
		), .Z(n_286259943));
	notech_ao4 i_208942501(.A(n_56592), .B(n_28164), .C(n_28489), .D(n_56579
		), .Z(n_286159942));
	notech_ao4 i_209142499(.A(n_56566), .B(n_28522), .C(n_56553), .D(n_27864
		), .Z(n_285959940));
	notech_ao4 i_209242498(.A(n_56547), .B(n_28566), .C(n_56513), .D(n_29718
		), .Z(n_285859939));
	notech_and2 i_10444496(.A(n_62820), .B(opc[6]), .Z(n_91719099));
	notech_nand2 i_44744493(.A(n_62820), .B(opc_10[6]), .Z(n_92019102));
	notech_nao3 i_58243925(.A(n_56463), .B(\opa_12[6] ), .C(n_1433), .Z(n_283659917
		));
	notech_nao3 i_56743940(.A(n_60294), .B(n_276659847), .C(n_32446), .Z(n_283559916
		));
	notech_nao3 i_56643941(.A(n_27075), .B(\opa_12[6] ), .C(n_56979), .Z(n_283459915
		));
	notech_nao3 i_56543942(.A(opd[6]), .B(n_58078), .C(n_56513), .Z(n_283359914
		));
	notech_and2 i_57043937(.A(n_276959850), .B(n_27061), .Z(n_283259913));
	notech_or4 i_57343934(.A(n_56829), .B(n_56979), .C(n_56513), .D(n_3868),
		 .Z(n_282959910));
	notech_nao3 i_60455613(.A(n_60113), .B(n_60294), .C(n_212859209), .Z(n_281259893
		));
	notech_nand3 i_25044246(.A(n_310991714), .B(\regs_1[5] ), .C(n_28680), .Z
		(n_279559876));
	notech_nand3 i_23544261(.A(n_310991714), .B(\regs_1[3] ), .C(n_28680), .Z
		(n_278059861));
	notech_and3 i_79153914(.A(n_57592), .B(n_341191462), .C(n_57957), .Z(n_277959860
		));
	notech_ao4 i_121643346(.A(n_58062), .B(n_2937), .C(n_27896), .D(n_27046)
		, .Z(n_277459855));
	notech_nand3 i_13944357(.A(n_92619108), .B(n_287659957), .C(n_283659917)
		, .Z(n_276959850));
	notech_and2 i_13844358(.A(n_57314), .B(n_287859959), .Z(n_276859849));
	notech_ao4 i_13744359(.A(n_27746), .B(n_56082), .C(n_26601), .D(n_26802)
		, .Z(n_276759848));
	notech_nand2 i_13644360(.A(n_3866), .B(n_3865), .Z(n_276659847));
	notech_ao4 i_16644330(.A(n_305991764), .B(n_24583), .C(n_61103), .D(n_30825
		), .Z(n_276459845));
	notech_and2 i_16544331(.A(n_57615), .B(n_28222), .Z(n_276359844));
	notech_and2 i_16444332(.A(n_298991830), .B(n_26773), .Z(n_276259843));
	notech_nao3 i_127953972(.A(n_57957), .B(n_312960210), .C(n_3633), .Z(n_276159842
		));
	notech_ao3 i_123246508(.A(n_296969981), .B(n_281259893), .C(n_267959760)
		, .Z(n_275959840));
	notech_ao4 i_123346507(.A(n_59095), .B(n_28105), .C(n_308591738), .D(n_28001
		), .Z(n_275659837));
	notech_ao4 i_123446506(.A(n_305491769), .B(n_56284), .C(n_2990), .D(n_57680
		), .Z(n_275559836));
	notech_and4 i_124246498(.A(n_275259833), .B(n_275059831), .C(n_274759828
		), .D(n_268659767), .Z(n_275459835));
	notech_ao4 i_123746503(.A(n_313747721), .B(n_150228779), .C(n_307891745)
		, .D(n_252966058), .Z(n_275259833));
	notech_ao4 i_123946501(.A(n_254466073), .B(n_267659757), .C(n_306791756)
		, .D(n_267559756), .Z(n_275059831));
	notech_ao4 i_124446496(.A(n_305891765), .B(n_57680), .C(n_24590), .D(n_56284
		), .Z(n_274859829));
	notech_ao4 i_124046500(.A(n_29710), .B(n_27080), .C(n_60009), .D(n_187592028
		), .Z(n_274759828));
	notech_and4 i_126046481(.A(n_281259893), .B(n_274459825), .C(n_274259823
		), .D(n_269859779), .Z(n_274659827));
	notech_ao4 i_125646485(.A(n_26648), .B(n_29709), .C(n_3836), .D(n_57698)
		, .Z(n_274459825));
	notech_ao4 i_125846483(.A(n_150728784), .B(n_3864), .C(n_150628783), .D(n_29711
		), .Z(n_274259823));
	notech_and4 i_126646475(.A(n_273959820), .B(n_273759818), .C(n_273659817
		), .D(n_270159782), .Z(n_274159822));
	notech_ao4 i_126146480(.A(n_308591738), .B(n_28003), .C(n_60113), .D(n_27138
		), .Z(n_273959820));
	notech_ao4 i_126346478(.A(n_150228779), .B(n_3861), .C(n_308791736), .D(n_77522039
		), .Z(n_273759818));
	notech_ao4 i_126446477(.A(n_307891745), .B(n_95222216), .C(n_60121865), 
		.D(n_306791756), .Z(n_273659817));
	notech_or4 i_30947695(.A(n_60964), .B(n_60953), .C(n_62850), .D(n_57698)
		, .Z(n_60121865));
	notech_nand2 i_1847704(.A(n_62820), .B(opc_10[18]), .Z(n_77522039));
	notech_ao4 i_205145732(.A(n_56666), .B(n_28243), .C(n_56653), .D(n_28208
		), .Z(n_273359814));
	notech_ao4 i_205245731(.A(n_56916), .B(n_29713), .C(n_56640), .D(n_28275
		), .Z(n_273259813));
	notech_and2 i_205645727(.A(n_273059811), .B(n_272959810), .Z(n_273159812
		));
	notech_ao4 i_205445729(.A(n_56532), .B(n_28308), .C(n_56518), .D(n_29712
		), .Z(n_273059811));
	notech_ao4 i_205545728(.A(n_56502), .B(n_28373), .C(n_56489), .D(n_28341
		), .Z(n_272959810));
	notech_and4 i_206445719(.A(n_272659807), .B(n_272559806), .C(n_272359804
		), .D(n_272259803), .Z(n_272859809));
	notech_ao4 i_205845725(.A(n_56627), .B(n_28437), .C(n_56614), .D(n_28405
		), .Z(n_272659807));
	notech_ao4 i_205945724(.A(n_56605), .B(n_28469), .C(n_56592), .D(n_28176
		), .Z(n_272559806));
	notech_ao4 i_206145722(.A(n_56583), .B(n_28501), .C(n_56553), .D(n_27876
		), .Z(n_272359804));
	notech_ao4 i_206245721(.A(n_56547), .B(n_28579), .C(n_56566), .D(n_28539
		), .Z(n_272259803));
	notech_nand2 i_29147700(.A(n_62820), .B(opc[18]), .Z(n_95222216));
	notech_or4 i_18447516(.A(n_61131), .B(n_60298), .C(n_60283), .D(n_28107)
		, .Z(n_270159782));
	notech_or2 i_18747513(.A(n_150528782), .B(n_56302), .Z(n_269859779));
	notech_or4 i_16547535(.A(n_55581), .B(n_24582), .C(n_57078), .D(n_57051)
		, .Z(n_269159772));
	notech_nand2 i_15547545(.A(sav_ecx[16]), .B(n_61133), .Z(n_268659767));
	notech_and4 i_16047540(.A(\regs_1_0[16] ), .B(n_60113), .C(n_60252), .D(n_60283
		), .Z(n_267959760));
	notech_and3 i_8947610(.A(n_57799), .B(n_57841), .C(n_269159772), .Z(n_267659757
		));
	notech_and2 i_8847611(.A(n_312324377), .B(n_274859829), .Z(n_267559756)
		);
	notech_ao4 i_8747612(.A(n_59440), .B(n_27079), .C(n_26775), .D(n_27274),
		 .Z(n_267459755));
	notech_and3 i_110949586(.A(n_281259893), .B(n_230865837), .C(n_266959750
		), .Z(n_267159752));
	notech_ao4 i_110849587(.A(n_151861801), .B(n_29707), .C(n_151761800), .D
		(n_29706), .Z(n_266959750));
	notech_ao4 i_111049585(.A(n_344366972), .B(n_57841), .C(n_57889), .D(n_57552
		), .Z(n_266759748));
	notech_ao4 i_111149584(.A(\nbus_11358[2] ), .B(n_57890), .C(n_58409), .D
		(n_59259), .Z(n_266659747));
	notech_and4 i_112049575(.A(n_266359744), .B(n_266259743), .C(n_266059741
		), .D(n_265959740), .Z(n_266559746));
	notech_ao4 i_111449581(.A(n_28091), .B(n_59095), .C(n_60113), .D(n_27118
		), .Z(n_266359744));
	notech_ao4 i_111549580(.A(n_59991), .B(n_306091763), .C(n_26774), .D(n_58316
		), .Z(n_266259743));
	notech_ao4 i_111749578(.A(n_152472004), .B(n_151961802), .C(n_152572005)
		, .D(n_281363080), .Z(n_266059741));
	notech_ao4 i_111849577(.A(n_261759698), .B(n_281463081), .C(n_24583), .D
		(n_261659697), .Z(n_265959740));
	notech_mux2 i_112149574(.S(n_32316), .A(n_312347735), .B(n_312447734), .Z
		(n_265859739));
	notech_mux2 i_112349573(.S(n_32316), .A(n_312147737), .B(n_344466973), .Z
		(n_265759738));
	notech_and4 i_112849568(.A(n_281259893), .B(n_265459735), .C(n_265259733
		), .D(n_264059721), .Z(n_265659737));
	notech_ao4 i_112449572(.A(n_26648), .B(n_29705), .C(n_150428781), .D(n_57742
		), .Z(n_265459735));
	notech_ao4 i_112649570(.A(n_150728784), .B(n_60003), .C(n_150628783), .D
		(n_29708), .Z(n_265259733));
	notech_and4 i_113349563(.A(n_264959730), .B(n_264759728), .C(n_264359724
		), .D(n_264659727), .Z(n_265159732));
	notech_ao4 i_112949567(.A(n_308591738), .B(n_28007), .C(n_60113), .D(n_27144
		), .Z(n_264959730));
	notech_ao4 i_113149565(.A(n_308791736), .B(n_225765786), .C(n_307891745)
		, .D(n_224065769), .Z(n_264759728));
	notech_or2 i_14150526(.A(n_150228779), .B(n_289227274), .Z(n_264659727)
		);
	notech_or4 i_14450523(.A(n_61133), .B(n_60298), .C(n_60283), .D(n_28111)
		, .Z(n_264359724));
	notech_or2 i_14750520(.A(n_150528782), .B(n_56338), .Z(n_264059721));
	notech_and2 i_5550611(.A(n_58717), .B(n_265859739), .Z(n_261759698));
	notech_and2 i_5450612(.A(n_265759738), .B(n_58714), .Z(n_261659697));
	notech_and4 i_188552093(.A(n_261359694), .B(n_261259693), .C(n_261059691
		), .D(n_260959690), .Z(n_261559696));
	notech_ao4 i_187952099(.A(n_55389), .B(n_28622), .C(n_55378), .D(n_29375
		), .Z(n_261359694));
	notech_ao4 i_187852100(.A(n_59153), .B(n_29313), .C(n_59335), .D(n_29344
		), .Z(n_261259693));
	notech_ao4 i_187752101(.A(n_59167), .B(n_29704), .C(n_59176), .D(n_27832
		), .Z(n_261059691));
	notech_ao4 i_187652102(.A(n_55409), .B(n_29702), .C(n_55420), .D(n_29701
		), .Z(n_260959690));
	notech_ao4 i_188152097(.A(n_55367), .B(n_28416), .C(n_55400), .D(n_28014
		), .Z(n_260759688));
	notech_ao4 i_188052098(.A(n_55429), .B(n_55956), .C(n_55347), .D(nbus_11295
		[29]), .Z(n_260659687));
	notech_ao4 i_168452292(.A(n_172792106), .B(n_311491709), .C(n_174492092)
		, .D(n_311391710), .Z(n_260459685));
	notech_and4 i_168252294(.A(n_260059681), .B(n_259959680), .C(n_259759678
		), .D(n_238059461), .Z(n_260259683));
	notech_ao4 i_167952297(.A(n_29662), .B(n_26696), .C(n_130528582), .D(n_151428791
		), .Z(n_260059681));
	notech_ao4 i_167852298(.A(n_311191712), .B(\nbus_11358[28] ), .C(n_311091713
		), .D(\nbus_11365[28] ), .Z(n_259959680));
	notech_ao4 i_167752299(.A(n_59124), .B(nbus_11295[28]), .C(n_54638), .D(n_28959
		), .Z(n_259759678));
	notech_nand3 i_164352333(.A(n_258859669), .B(n_258759668), .C(n_259359674
		), .Z(n_259459675));
	notech_and4 i_164252334(.A(n_281259893), .B(n_259059671), .C(n_236959450
		), .D(n_236259443), .Z(n_259359674));
	notech_ao4 i_163952337(.A(n_308591738), .B(n_28011), .C(n_59095), .D(n_28115
		), .Z(n_259059671));
	notech_ao4 i_163852338(.A(n_150628783), .B(n_29660), .C(n_133728614), .D
		(n_150728784), .Z(n_258859669));
	notech_ao4 i_163752339(.A(n_150528782), .B(n_55947), .C(n_150428781), .D
		(\nbus_11365[26] ), .Z(n_258759668));
	notech_and4 i_162252354(.A(n_258059661), .B(n_257859659), .C(n_257759658
		), .D(n_258359664), .Z(n_258559666));
	notech_and3 i_161952357(.A(n_281259893), .B(n_258259663), .C(n_235059431
		), .Z(n_258359664));
	notech_ao4 i_161552361(.A(n_150428781), .B(n_57792), .C(n_310091723), .D
		(n_308791736), .Z(n_258259663));
	notech_ao4 i_161852358(.A(n_60113), .B(n_27149), .C(n_308591738), .D(n_28012
		), .Z(n_258059661));
	notech_ao4 i_161752359(.A(n_59095), .B(n_28116), .C(n_150628783), .D(n_29661
		), .Z(n_257859659));
	notech_ao4 i_161652360(.A(n_131228589), .B(n_150728784), .C(n_150528782)
		, .D(n_55938), .Z(n_257759658));
	notech_nand3 i_157852398(.A(n_256859649), .B(n_256759648), .C(n_257359654
		), .Z(n_257459655));
	notech_and4 i_157752399(.A(n_281259893), .B(n_257059651), .C(n_234559426
		), .D(n_233859419), .Z(n_257359654));
	notech_ao4 i_157452402(.A(n_308591738), .B(n_28014), .C(n_59095), .D(n_28118
		), .Z(n_257059651));
	notech_ao4 i_157352403(.A(n_150628783), .B(n_29659), .C(n_128228559), .D
		(n_150728784), .Z(n_256859649));
	notech_ao4 i_157252404(.A(n_150528782), .B(n_55956), .C(n_150428781), .D
		(\nbus_11365[29] ), .Z(n_256759648));
	notech_and4 i_155652420(.A(n_256159642), .B(n_256059641), .C(n_255959640
		), .D(n_3884), .Z(n_256459645));
	notech_ao4 i_155252424(.A(n_133728614), .B(n_149128768), .C(n_149428771)
		, .D(n_55947), .Z(n_256159642));
	notech_ao4 i_155152425(.A(n_149328770), .B(n_57783), .C(n_54638), .D(n_28980
		), .Z(n_256059641));
	notech_ao4 i_155352423(.A(n_310691717), .B(n_28011), .C(n_149228769), .D
		(n_29660), .Z(n_255959640));
	notech_and4 i_151952457(.A(n_255359634), .B(n_255259633), .C(n_255159632
		), .D(n_232359404), .Z(n_255659637));
	notech_ao4 i_151552461(.A(n_130528582), .B(n_149128768), .C(n_149428771)
		, .D(n_55974), .Z(n_255359634));
	notech_ao4 i_151452462(.A(n_149328770), .B(\nbus_11365[28] ), .C(n_54638
		), .D(n_28983), .Z(n_255259633));
	notech_ao4 i_151652460(.A(n_310691717), .B(n_28013), .C(n_149228769), .D
		(n_29662), .Z(n_255159632));
	notech_ao4 i_144652525(.A(n_172792106), .B(n_3858), .C(n_174492092), .D(n_3843
		), .Z(n_254959630));
	notech_and4 i_144452527(.A(n_54667), .B(n_254559626), .C(n_254359624), .D
		(n_230859389), .Z(n_254759628));
	notech_ao4 i_144152530(.A(n_130528582), .B(n_148228759), .C(n_3877), .D(n_55974
		), .Z(n_254559626));
	notech_ao4 i_144252529(.A(n_3857), .B(n_28013), .C(n_29662), .D(n_26642)
		, .Z(n_254359624));
	notech_and4 i_136152609(.A(n_253359614), .B(n_253259613), .C(n_230459385
		), .D(n_253959620), .Z(n_254159622));
	notech_and3 i_135952611(.A(n_253759618), .B(n_253659617), .C(n_253559616
		), .Z(n_253959620));
	notech_ao4 i_135352617(.A(n_146928746), .B(\nbus_11365[28] ), .C(n_54865
		), .D(n_29700), .Z(n_253759618));
	notech_ao4 i_135252618(.A(n_54883), .B(n_28621), .C(n_54894), .D(n_27481
		), .Z(n_253659617));
	notech_ao4 i_135652614(.A(n_60113), .B(n_27185), .C(n_310391720), .D(n_28013
		), .Z(n_253559616));
	notech_ao4 i_135552615(.A(n_54874), .B(n_28117), .C(n_147128748), .D(n_29662
		), .Z(n_253359614));
	notech_ao4 i_135452616(.A(n_130528582), .B(n_147228749), .C(n_147028747)
		, .D(n_55974), .Z(n_253259613));
	notech_and4 i_133652634(.A(n_252259603), .B(n_252159602), .C(n_229059371
		), .D(n_252859609), .Z(n_253059611));
	notech_and3 i_133452636(.A(n_252659607), .B(n_252559606), .C(n_252459605
		), .Z(n_252859609));
	notech_ao4 i_132852642(.A(n_146928746), .B(n_57815), .C(n_54865), .D(n_29699
		), .Z(n_252659607));
	notech_ao4 i_132752643(.A(n_54883), .B(n_28622), .C(n_54894), .D(n_27483
		), .Z(n_252559606));
	notech_ao4 i_133152639(.A(n_60117), .B(n_27186), .C(n_310391720), .D(n_28014
		), .Z(n_252459605));
	notech_ao4 i_133052640(.A(n_54874), .B(n_28118), .C(n_147128748), .D(n_29659
		), .Z(n_252259603));
	notech_ao4 i_132952641(.A(n_128228559), .B(n_147228749), .C(n_147028747)
		, .D(n_55956), .Z(n_252159602));
	notech_nand3 i_119852770(.A(n_251259593), .B(n_251159592), .C(n_251759598
		), .Z(n_251859599));
	notech_and3 i_119752771(.A(n_251559596), .B(n_251459595), .C(n_227559356
		), .Z(n_251759598));
	notech_ao4 i_119152777(.A(n_54658), .B(n_29698), .C(n_27334), .D(n_29697
		), .Z(n_251559596));
	notech_ao4 i_119452774(.A(n_27319), .B(n_28013), .C(n_59322), .D(n_28117
		), .Z(n_251459595));
	notech_ao4 i_119352775(.A(n_145028727), .B(n_29662), .C(n_130528582), .D
		(n_145128728), .Z(n_251259593));
	notech_ao4 i_119252776(.A(n_144928726), .B(n_55974), .C(n_144828725), .D
		(n_57802), .Z(n_251159592));
	notech_nand3 i_117552793(.A(n_250259583), .B(n_250159582), .C(n_250759588
		), .Z(n_250859589));
	notech_and3 i_117452794(.A(n_250559586), .B(n_250459585), .C(n_226359344
		), .Z(n_250759588));
	notech_ao4 i_116852800(.A(n_27335), .B(n_29696), .C(n_27334), .D(n_29695
		), .Z(n_250559586));
	notech_ao4 i_117152797(.A(n_27319), .B(n_28014), .C(n_59322), .D(n_28118
		), .Z(n_250459585));
	notech_ao4 i_117052798(.A(n_145028727), .B(n_29659), .C(n_128228559), .D
		(n_145128728), .Z(n_250259583));
	notech_ao4 i_116952799(.A(n_144928726), .B(n_55956), .C(n_144828725), .D
		(n_57815), .Z(n_250159582));
	notech_and4 i_102852938(.A(n_249459575), .B(n_249759578), .C(n_225359334
		), .D(n_225059331), .Z(n_249959580));
	notech_ao4 i_102652940(.A(n_308547770), .B(n_27100), .C(n_224559326), .D
		(n_27857), .Z(n_249759578));
	notech_ao4 i_100952955(.A(n_27105), .B(n_29116), .C(n_57132), .D(n_28925
		), .Z(n_249659577));
	notech_ao4 i_102452942(.A(n_27781), .B(n_29693), .C(n_27782), .D(n_28679
		), .Z(n_249459575));
	notech_ao4 i_99752967(.A(n_222259303), .B(n_27850), .C(n_1889), .D(n_29692
		), .Z(n_249159572));
	notech_ao4 i_99152973(.A(n_27105), .B(n_28942), .C(n_57132), .D(n_28668)
		, .Z(n_249059571));
	notech_and4 i_98652978(.A(n_248459565), .B(n_248359564), .C(n_248159562)
		, .D(n_248059561), .Z(n_248659567));
	notech_ao4 i_98052984(.A(n_57542), .B(n_27898), .C(n_57563), .D(n_27901)
		, .Z(n_248459565));
	notech_ao4 i_97952985(.A(n_57552), .B(n_27899), .C(n_57583), .D(n_27905)
		, .Z(n_248359564));
	notech_ao4 i_97852986(.A(n_57574), .B(n_27902), .C(n_57957), .D(n_27910)
		, .Z(n_248159562));
	notech_ao4 i_97752987(.A(n_57592), .B(n_27909), .C(n_57613), .D(n_27912)
		, .Z(n_248059561));
	notech_and4 i_98552979(.A(n_247759558), .B(n_247659557), .C(n_247459555)
		, .D(n_247359554), .Z(n_247959560));
	notech_ao4 i_97652988(.A(n_57604), .B(n_27911), .C(n_57635), .D(n_27914)
		, .Z(n_247759558));
	notech_ao4 i_97552989(.A(\nbus_11307[10] ), .B(n_27913), .C(n_57653), .D
		(n_27916), .Z(n_247659557));
	notech_ao4 i_97452990(.A(n_57644), .B(n_27915), .C(\nbus_11307[15] ), .D
		(n_27923), .Z(n_247459555));
	notech_ao4 i_97352991(.A(n_57662), .B(n_27918), .C(\nbus_11365[17] ), .D
		(n_27927), .Z(n_247359554));
	notech_and4 i_95553008(.A(n_246959550), .B(n_246859549), .C(n_246659547)
		, .D(n_246559546), .Z(n_247159552));
	notech_ao4 i_94953014(.A(n_57815), .B(n_27939), .C(n_57802), .D(n_27938)
		, .Z(n_246959550));
	notech_ao4 i_94853015(.A(n_57792), .B(n_27937), .C(n_57783), .D(n_27936)
		, .Z(n_246859549));
	notech_ao4 i_94753016(.A(n_57680), .B(n_27926), .C(n_57707), .D(n_27929)
		, .Z(n_246659547));
	notech_ao4 i_94653017(.A(\nbus_11365[18] ), .B(n_27928), .C(n_57733), .D
		(n_27931), .Z(n_246559546));
	notech_and4 i_95453009(.A(n_246259543), .B(n_246159542), .C(n_245959540)
		, .D(n_245859539), .Z(n_246459545));
	notech_ao4 i_94553018(.A(n_57720), .B(n_27930), .C(n_57751), .D(n_27933)
		, .Z(n_246259543));
	notech_ao4 i_94453019(.A(n_57742), .B(n_27932), .C(n_57771), .D(n_27935)
		, .Z(n_246159542));
	notech_ao4 i_94353020(.A(n_57761), .B(n_27934), .C(n_59726), .D(n_27941)
		, .Z(n_245959540));
	notech_ao4 i_94253021(.A(n_57828), .B(n_27940), .C(n_59742), .D(n_27897)
		, .Z(n_245859539));
	notech_ao4 i_100552959(.A(n_223159312), .B(n_26638), .C(CFOF_mul), .D(n_3986
		), .Z(n_245759538));
	notech_nand3 i_87153090(.A(n_244859529), .B(n_244759528), .C(n_245359534
		), .Z(n_245459535));
	notech_and3 i_87053091(.A(n_245159532), .B(n_245059531), .C(n_218359264)
		, .Z(n_245359534));
	notech_ao4 i_86453097(.A(n_54649), .B(n_29691), .C(n_28527), .D(n_29690)
		, .Z(n_245159532));
	notech_ao4 i_86753094(.A(n_303591788), .B(n_28013), .C(n_59322), .D(n_28117
		), .Z(n_245059531));
	notech_ao4 i_86653095(.A(n_140328680), .B(n_29662), .C(n_130528582), .D(n_140428681
		), .Z(n_244859529));
	notech_ao4 i_86553096(.A(n_140228679), .B(n_55974), .C(n_140128678), .D(n_57802
		), .Z(n_244759528));
	notech_nand3 i_84653113(.A(n_243859519), .B(n_243759518), .C(n_244359524
		), .Z(n_244459525));
	notech_and3 i_84553114(.A(n_244159522), .B(n_244059521), .C(n_217059251)
		, .Z(n_244359524));
	notech_ao4 i_83953120(.A(n_54649), .B(n_29689), .C(n_28527), .D(n_29687)
		, .Z(n_244159522));
	notech_ao4 i_84253117(.A(n_303591788), .B(n_28014), .C(n_59326), .D(n_28118
		), .Z(n_244059521));
	notech_ao4 i_84153118(.A(n_140328680), .B(n_29659), .C(n_128228559), .D(n_140428681
		), .Z(n_243859519));
	notech_ao4 i_84053119(.A(n_140228679), .B(n_55956), .C(n_140128678), .D(n_57815
		), .Z(n_243759518));
	notech_and4 i_68153272(.A(n_215759238), .B(n_243159512), .C(n_243059511)
		, .D(n_3884), .Z(n_243459515));
	notech_ao4 i_67753276(.A(n_251362780), .B(n_55947), .C(n_250962776), .D(n_57783
		), .Z(n_243159512));
	notech_ao4 i_67853275(.A(n_29660), .B(n_251162778), .C(n_133728614), .D(n_251262779
		), .Z(n_243059511));
	notech_and4 i_64953304(.A(n_214859229), .B(n_242459505), .C(n_242359504)
		, .D(n_232359404), .Z(n_242759508));
	notech_ao4 i_64553308(.A(n_251362780), .B(n_55974), .C(n_250962776), .D(n_57802
		), .Z(n_242459505));
	notech_ao4 i_64653307(.A(n_251162778), .B(n_29662), .C(n_130528582), .D(n_251262779
		), .Z(n_242359504));
	notech_and3 i_68453917(.A(n_242059501), .B(n_241959500), .C(n_232359404)
		, .Z(n_242259503));
	notech_ao4 i_42753523(.A(n_309591728), .B(n_29662), .C(n_130528582), .D(n_30803
		), .Z(n_242059501));
	notech_ao4 i_42653524(.A(n_304691777), .B(n_55974), .C(n_309491729), .D(n_57802
		), .Z(n_241959500));
	notech_nand2 i_13353780(.A(n_57635), .B(n_57625), .Z(n_241659497));
	notech_or4 i_15753778(.A(opa[13]), .B(opa[12]), .C(opa[15]), .D(opa[14])
		, .Z(n_241559496));
	notech_and4 i_11953794(.A(n_57815), .B(n_57802), .C(n_57792), .D(n_57783
		), .Z(n_241159492));
	notech_and4 i_11853795(.A(n_57680), .B(n_57689), .C(n_57698), .D(n_57707
		), .Z(n_240859489));
	notech_and4 i_11753796(.A(n_57720), .B(n_57733), .C(n_57742), .D(n_57751
		), .Z(n_240459485));
	notech_and4 i_11653797(.A(\nbus_11365[24] ), .B(n_57771), .C(n_57828), .D
		(n_59726), .Z(n_240159482));
	notech_nand3 i_3018995(.A(n_260759688), .B(n_260659687), .C(n_261559696)
		, .Z(n_239659477));
	notech_and4 i_2917618(.A(n_260259683), .B(n_260459685), .C(n_242259503),
		 .D(n_237359454), .Z(n_238359464));
	notech_or4 i_167352303(.A(n_56829), .B(n_56941), .C(n_56583), .D(n_28013
		), .Z(n_238059461));
	notech_or2 i_167452302(.A(n_151128788), .B(n_3982), .Z(n_237359454));
	notech_or4 i_2717040(.A(n_237059451), .B(n_237159452), .C(n_236159442), 
		.D(n_259459675), .Z(n_237259453));
	notech_ao3 i_163552341(.A(opc[26]), .B(n_62812), .C(n_307891745), .Z(n_237159452
		));
	notech_ao3 i_163452342(.A(opc_10[26]), .B(n_62812), .C(n_308791736), .Z(n_237059451
		));
	notech_nand2 i_163252344(.A(sav_ecx[26]), .B(n_61133), .Z(n_236959450)
		);
	notech_nao3 i_162552351(.A(\regs_1_0[26] ), .B(n_60283), .C(n_59326), .Z
		(n_236259443));
	notech_nor2 i_163352343(.A(n_3983), .B(n_150228779), .Z(n_236159442));
	notech_nand3 i_2817041(.A(n_258559666), .B(n_235959440), .C(n_234959430)
		, .Z(n_236059441));
	notech_nao3 i_161352363(.A(opc[27]), .B(n_62812), .C(n_307891745), .Z(n_235959440
		));
	notech_nao3 i_160352373(.A(\regs_1_0[27] ), .B(n_60283), .C(n_59326), .Z
		(n_235059431));
	notech_or2 i_161252364(.A(n_4016), .B(n_150228779), .Z(n_234959430));
	notech_or4 i_3017043(.A(n_234659427), .B(n_234759428), .C(n_233759418), 
		.D(n_257459655), .Z(n_234859429));
	notech_ao3 i_157052406(.A(opc[29]), .B(n_62812), .C(n_307891745), .Z(n_234759428
		));
	notech_ao3 i_156952407(.A(opc_10[29]), .B(n_62812), .C(n_308791736), .Z(n_234659427
		));
	notech_nand2 i_156752409(.A(sav_ecx[29]), .B(n_61133), .Z(n_234559426)
		);
	notech_nao3 i_156052416(.A(\regs_1_0[29] ), .B(n_60283), .C(n_59326), .Z
		(n_233859419));
	notech_nor2 i_156852408(.A(n_3981), .B(n_150228779), .Z(n_233759418));
	notech_or4 i_2721936(.A(n_233459415), .B(n_233559416), .C(n_232759408), 
		.D(n_27082), .Z(n_233659417));
	notech_ao3 i_155052426(.A(opc[26]), .B(n_62812), .C(n_310891715), .Z(n_233559416
		));
	notech_ao3 i_154952427(.A(opc_10[26]), .B(n_62812), .C(n_310791716), .Z(n_233459415
		));
	notech_nor2 i_154852428(.A(n_148728764), .B(n_3983), .Z(n_232759408));
	notech_or4 i_2921938(.A(n_232459405), .B(n_232559406), .C(n_231659397), 
		.D(n_27083), .Z(n_232659407));
	notech_ao3 i_151352463(.A(opc[28]), .B(n_62812), .C(n_310891715), .Z(n_232559406
		));
	notech_ao3 i_151252464(.A(opc_10[28]), .B(n_62812), .C(n_310791716), .Z(n_232459405
		));
	notech_nand2 i_206053907(.A(read_data[28]), .B(n_60252), .Z(n_232359404)
		);
	notech_nor2 i_151152465(.A(n_148728764), .B(n_3982), .Z(n_231659397));
	notech_and4 i_2921874(.A(n_242259503), .B(n_254759628), .C(n_254959630),
		 .D(n_230759388), .Z(n_231559396));
	notech_or2 i_143252539(.A(n_3878), .B(n_57802), .Z(n_230859389));
	notech_or2 i_143752534(.A(n_3982), .B(n_3837), .Z(n_230759388));
	notech_nand3 i_2921810(.A(n_254159622), .B(n_230559386), .C(n_229359374)
		, .Z(n_230659387));
	notech_or4 i_135152619(.A(n_312191702), .B(nbus_11295[28]), .C(n_60935),
		 .D(n_54929), .Z(n_230559386));
	notech_nao3 i_135052620(.A(opc_10[28]), .B(n_62812), .C(n_301791806), .Z
		(n_230459385));
	notech_or2 i_134952621(.A(n_146428741), .B(n_3982), .Z(n_229359374));
	notech_nand3 i_3021811(.A(n_253059611), .B(n_229159372), .C(n_227959360)
		, .Z(n_229259373));
	notech_or4 i_132652644(.A(n_312191702), .B(nbus_11295[29]), .C(n_60935),
		 .D(n_54929), .Z(n_229159372));
	notech_nao3 i_132552645(.A(opc_10[29]), .B(n_62812), .C(n_301791806), .Z
		(n_229059371));
	notech_or2 i_132452646(.A(n_146428741), .B(n_3981), .Z(n_227959360));
	notech_or4 i_2921554(.A(n_227659357), .B(n_251859599), .C(n_227759358), 
		.D(n_226759348), .Z(n_227859359));
	notech_and3 i_119052778(.A(opc[28]), .B(n_62812), .C(n_27340), .Z(n_227759358
		));
	notech_ao3 i_118952779(.A(opc_10[28]), .B(n_62812), .C(n_27329), .Z(n_227659357
		));
	notech_nand2 i_118752781(.A(sav_esi[28]), .B(n_61133), .Z(n_227559356)
		);
	notech_nor2 i_118852780(.A(n_144428721), .B(n_3982), .Z(n_226759348));
	notech_or4 i_3021555(.A(n_226459345), .B(n_250859589), .C(n_226559346), 
		.D(n_225559336), .Z(n_226659347));
	notech_and3 i_116752801(.A(opc[29]), .B(n_62812), .C(n_27340), .Z(n_226559346
		));
	notech_ao3 i_116652802(.A(opc_10[29]), .B(n_62812), .C(n_27329), .Z(n_226459345
		));
	notech_nand2 i_116452804(.A(sav_esi[29]), .B(n_61133), .Z(n_226359344)
		);
	notech_nor2 i_116552803(.A(n_144428721), .B(n_3981), .Z(n_225559336));
	notech_and4 i_7720(.A(n_222359304), .B(n_249159572), .C(n_249959580), .D
		(n_224359324), .Z(n_225459335));
	notech_nao3 i_102252944(.A(n_27096), .B(n_276159842), .C(n_27879), .Z(n_225359334
		));
	notech_nand2 i_102052946(.A(n_224659327), .B(n_60252), .Z(n_225059331)
		);
	notech_mux2 i_2353886(.S(n_26782), .A(nbus_163[16]), .B(nbus_162[32]), .Z
		(n_224759328));
	notech_mux2 i_2453885(.S(n_57899), .A(nCF_shiftbox), .B(nCF_shift4box), 
		.Z(n_224659327));
	notech_and2 i_2553884(.A(n_249659577), .B(n_223659317), .Z(n_224559326)
		);
	notech_and2 i_2953883(.A(n_223259313), .B(n_245759538), .Z(n_224459325)
		);
	notech_or4 i_101852948(.A(fsm[2]), .B(n_61165), .C(n_61156), .D(n_224459325
		), .Z(n_224359324));
	notech_nand3 i_100852956(.A(nbus_160[32]), .B(n_59440), .C(n_60298), .Z(n_223659317
		));
	notech_ao4 i_3053882(.A(n_277959860), .B(n_27096), .C(n_27896), .D(n_3632
		), .Z(n_223359314));
	notech_or4 i_100452960(.A(n_27573), .B(n_59419), .C(n_223359314), .D(n_28081
		), .Z(n_223259313));
	notech_ao4 i_3153881(.A(n_27096), .B(n_28635), .C(n_27896), .D(n_28802),
		 .Z(n_223159312));
	notech_and4 i_3953873(.A(n_248659567), .B(n_247959560), .C(n_247159552),
		 .D(n_246459545), .Z(n_222459305));
	notech_or4 i_99452970(.A(n_315291671), .B(n_60868), .C(n_222459305), .D(n_60257
		), .Z(n_222359304));
	notech_and2 i_3853874(.A(n_249059571), .B(n_221959300), .Z(n_222259303)
		);
	notech_nand3 i_99052974(.A(nbus_161[16]), .B(n_59441), .C(n_60298), .Z(n_221959300
		));
	notech_or4 i_2921362(.A(n_218459265), .B(n_245459535), .C(n_218559266), 
		.D(n_217459255), .Z(n_218659267));
	notech_and3 i_86353098(.A(opc[28]), .B(n_62768), .C(n_309791726), .Z(n_218559266
		));
	notech_ao3 i_86253099(.A(opc_10[28]), .B(n_62812), .C(n_309691727), .Z(n_218459265
		));
	notech_nand2 i_86053101(.A(sav_edi[28]), .B(n_61133), .Z(n_218359264));
	notech_nor2 i_86153100(.A(n_139728674), .B(n_3982), .Z(n_217459255));
	notech_or4 i_3021363(.A(n_217159252), .B(n_244459525), .C(n_217259253), 
		.D(n_216159242), .Z(n_217359254));
	notech_and3 i_83853121(.A(opc[29]), .B(n_62770), .C(n_309791726), .Z(n_217259253
		));
	notech_ao3 i_83753122(.A(opc_10[29]), .B(n_62792), .C(n_309691727), .Z(n_217159252
		));
	notech_nand2 i_83553124(.A(sav_edi[29]), .B(n_61133), .Z(n_217059251));
	notech_nor2 i_83653123(.A(n_139728674), .B(n_3981), .Z(n_216159242));
	notech_or4 i_2721040(.A(n_215859239), .B(n_215959240), .C(n_215259233), 
		.D(n_27098), .Z(n_216059241));
	notech_and3 i_67653277(.A(opc[26]), .B(n_62792), .C(n_26762), .Z(n_215959240
		));
	notech_ao3 i_67553278(.A(opc_10[26]), .B(n_62792), .C(n_316537960), .Z(n_215859239
		));
	notech_or4 i_67353280(.A(n_56832), .B(n_56941), .C(n_56627), .D(n_28011)
		, .Z(n_215759238));
	notech_nor2 i_67453279(.A(n_322438019), .B(n_3983), .Z(n_215259233));
	notech_or4 i_2921042(.A(n_214959230), .B(n_215059231), .C(n_214359224), 
		.D(n_27099), .Z(n_215159232));
	notech_and3 i_64453309(.A(opc[28]), .B(n_62792), .C(n_26762), .Z(n_215059231
		));
	notech_ao3 i_64353310(.A(opc_10[28]), .B(n_62792), .C(n_316537960), .Z(n_214959230
		));
	notech_or4 i_64153312(.A(n_56832), .B(n_56941), .C(n_56627), .D(n_28013)
		, .Z(n_214859229));
	notech_nor2 i_64253311(.A(n_322438019), .B(n_3982), .Z(n_214359224));
	notech_and4 i_64854908(.A(n_281259893), .B(n_213659217), .C(n_213459215)
		, .D(n_212159202), .Z(n_213859219));
	notech_ao4 i_64454912(.A(n_59095), .B(n_28121), .C(n_26648), .D(n_29685)
		, .Z(n_213659217));
	notech_ao4 i_64654910(.A(n_150228779), .B(n_303091793), .C(n_150428781),
		 .D(\nbus_11365[30] ), .Z(n_213459215));
	notech_and4 i_65354903(.A(n_213159212), .B(n_212959210), .C(n_212459205)
		, .D(n_212759208), .Z(n_213359214));
	notech_ao4 i_64954907(.A(n_150628783), .B(n_29591), .C(n_150728784), .D(n_302991794
		), .Z(n_213159212));
	notech_ao4 i_65154905(.A(n_308591738), .B(n_28015), .C(n_308791736), .D(n_30809
		), .Z(n_212959210));
	notech_or4 i_97854610(.A(n_27925), .B(n_32643), .C(n_59413), .D(n_27025)
		, .Z(n_212859209));
	notech_nao3 i_28755237(.A(n_62798), .B(opc[30]), .C(n_307891745), .Z(n_212759208
		));
	notech_or2 i_29055234(.A(n_150528782), .B(n_55929), .Z(n_212459205));
	notech_nand2 i_29355231(.A(sav_ecx[30]), .B(n_61133), .Z(n_212159202));
	notech_or4 i_47555050(.A(n_58062), .B(n_2937), .C(n_56829), .D(n_32284),
		 .Z(n_211359194));
	notech_or4 i_129255531(.A(instrc[122]), .B(n_32614), .C(n_54954), .D(n_29179
		), .Z(n_26060));
	notech_and4 i_119157341(.A(n_281259893), .B(n_210959190), .C(n_210759188
		), .D(n_210659187), .Z(n_211159192));
	notech_ao4 i_118657346(.A(n_151861801), .B(n_29683), .C(n_151761800), .D
		(n_29682), .Z(n_210959190));
	notech_ao4 i_118857344(.A(n_305791766), .B(n_3851), .C(n_57799), .D(n_31433
		), .Z(n_210759188));
	notech_ao4 i_118957343(.A(n_58381), .B(n_27993), .C(n_31411), .D(n_24589
		), .Z(n_210659187));
	notech_and4 i_119757335(.A(n_210359184), .B(n_210159182), .C(n_210059181
		), .D(n_207159152), .Z(n_210559186));
	notech_ao4 i_119257340(.A(n_57984), .B(n_57625), .C(n_57936), .D(n_56145
		), .Z(n_210359184));
	notech_ao4 i_119457338(.A(n_57937), .B(n_3850), .C(n_59095), .D(n_28099)
		, .Z(n_210159182));
	notech_ao4 i_119557337(.A(n_60117), .B(n_27130), .C(n_87532846), .D(n_152061803
		), .Z(n_210059181));
	notech_and3 i_122657308(.A(n_3849), .B(n_207659157), .C(n_276134717), .Z
		(n_209859179));
	notech_ao4 i_122757307(.A(n_291663183), .B(n_305970070), .C(n_5723), .D(n_311791706
		), .Z(n_209559176));
	notech_ao4 i_122957306(.A(n_291863185), .B(n_306270073), .C(n_291763184)
		, .D(n_306170072), .Z(n_209459175));
	notech_and4 i_123757298(.A(n_209159172), .B(n_208959170), .C(n_208859169
		), .D(n_208359164), .Z(n_209359174));
	notech_ao4 i_123257303(.A(n_58410), .B(n_27986), .C(n_291463181), .D(n_24994
		), .Z(n_209159172));
	notech_ao4 i_123457301(.A(n_57891), .B(n_57574), .C(n_57938), .D(n_56055
		), .Z(n_208959170));
	notech_ao4 i_123557300(.A(n_5743), .B(n_57619), .C(n_57882), .D(n_56064)
		, .Z(n_208859169));
	notech_nand2 i_3658484(.A(n_62820), .B(opc[10]), .Z(n_87532846));
	notech_or4 i_35658138(.A(n_62844), .B(n_26697), .C(n_62792), .D(n_57574)
		, .Z(n_208359164));
	notech_nao3 i_36158133(.A(tsc[36]), .B(n_55820), .C(n_59469), .Z(n_207659157
		));
	notech_or2 i_31658177(.A(n_57983), .B(n_56154), .Z(n_207159152));
	notech_and4 i_129560502(.A(n_205959140), .B(n_205859139), .C(n_205659137
		), .D(n_205559136), .Z(n_206159142));
	notech_ao4 i_128960508(.A(n_61103), .B(n_212859209), .C(n_59095), .D(n_28090
		), .Z(n_205959140));
	notech_ao4 i_129060507(.A(n_281363080), .B(n_297866507), .C(n_57889), .D
		(n_57542), .Z(n_205859139));
	notech_ao4 i_129260505(.A(n_57890), .B(n_56010), .C(n_24583), .D(n_297666505
		), .Z(n_205659137));
	notech_ao4 i_129360504(.A(n_306091763), .B(n_59992), .C(n_57841), .D(n_298066509
		), .Z(n_205559136));
	notech_and4 i_130260495(.A(n_205259133), .B(n_205159132), .C(n_204959130
		), .D(n_204859129), .Z(n_205459135));
	notech_ao4 i_129660501(.A(n_60117), .B(n_27117), .C(n_58409), .D(n_59241
		), .Z(n_205259133));
	notech_ao4 i_129760500(.A(n_26774), .B(n_297766506), .C(n_58004), .D(n_60024
		), .Z(n_205159132));
	notech_ao4 i_129960498(.A(n_58003), .B(n_56019), .C(n_151761800), .D(n_29677
		), .Z(n_204959130));
	notech_ao4 i_130060497(.A(n_151861801), .B(n_29676), .C(n_151961802), .D
		(n_297966508), .Z(n_204859129));
	notech_and4 i_136060440(.A(n_281259893), .B(n_204559126), .C(n_204359124
		), .D(n_204259123), .Z(n_204759128));
	notech_ao4 i_135460445(.A(n_320070211), .B(n_24589), .C(n_59095), .D(n_28101
		), .Z(n_204559126));
	notech_ao4 i_135660443(.A(n_305791766), .B(n_59965), .C(n_57799), .D(n_320170212
		), .Z(n_204359124));
	notech_ao4 i_135760442(.A(n_60117), .B(n_27133), .C(n_58381), .D(n_27997
		), .Z(n_204259123));
	notech_and4 i_136660434(.A(n_203959120), .B(n_203759118), .C(n_203659117
		), .D(n_194659033), .Z(n_204159122));
	notech_ao4 i_136160439(.A(n_57983), .B(n_56221), .C(n_57937), .D(n_60013
		), .Z(n_203959120));
	notech_ao4 i_136360437(.A(n_57936), .B(n_29679), .C(n_151761800), .D(n_29675
		), .Z(n_203759118));
	notech_ao4 i_136460436(.A(n_151861801), .B(n_29674), .C(n_152061803), .D
		(n_156768584), .Z(n_203659117));
	notech_and3 i_136960431(.A(n_281259893), .B(n_111364642), .C(n_203259113
		), .Z(n_203459115));
	notech_ao4 i_136860432(.A(n_31540), .B(n_24589), .C(n_59100), .D(n_28102
		), .Z(n_203259113));
	notech_ao4 i_137060430(.A(n_305791766), .B(n_301691807), .C(n_57799), .D
		(n_31560), .Z(n_203059111));
	notech_ao4 i_137160429(.A(n_60117), .B(n_27134), .C(n_58381), .D(n_27998
		), .Z(n_202959110));
	notech_and4 i_138060420(.A(n_202659107), .B(n_202559106), .C(n_202359104
		), .D(n_202259103), .Z(n_202859109));
	notech_ao4 i_137460426(.A(n_57984), .B(n_57653), .C(n_57983), .D(n_56230
		), .Z(n_202659107));
	notech_ao4 i_137560425(.A(n_175262035), .B(n_31576), .C(n_151761800), .D
		(n_29673), .Z(n_202559106));
	notech_ao4 i_137760423(.A(n_151861801), .B(n_29672), .C(n_152061803), .D
		(n_30109), .Z(n_202359104));
	notech_ao4 i_137860422(.A(n_188857101), .B(n_302091803), .C(n_169761980)
		, .D(n_56239), .Z(n_202259103));
	notech_and3 i_138360417(.A(n_281259893), .B(n_164365172), .C(n_201859099
		), .Z(n_202059101));
	notech_ao4 i_138260418(.A(n_298166510), .B(n_24589), .C(n_59095), .D(n_28103
		), .Z(n_201859099));
	notech_ao4 i_138460416(.A(n_305791766), .B(n_59963), .C(n_57799), .D(n_298266511
		), .Z(n_201659097));
	notech_ao4 i_138560415(.A(n_60117), .B(n_27135), .C(n_58381), .D(n_27999
		), .Z(n_201559096));
	notech_and4 i_139460406(.A(n_201259093), .B(n_201159092), .C(n_200959090
		), .D(n_200859089), .Z(n_201459095));
	notech_ao4 i_138860412(.A(n_57984), .B(n_57662), .C(n_57983), .D(n_56248
		), .Z(n_201259093));
	notech_ao4 i_138960411(.A(n_298366512), .B(n_175262035), .C(n_151761800)
		, .D(n_29671), .Z(n_201159092));
	notech_ao4 i_139160409(.A(n_151861801), .B(n_29670), .C(n_152061803), .D
		(n_157165100), .Z(n_200959090));
	notech_ao4 i_139260408(.A(n_60011), .B(n_188857101), .C(n_56257), .D(n_169761980
		), .Z(n_200859089));
	notech_and4 i_141560386(.A(n_281259893), .B(n_200559086), .C(n_200359084
		), .D(n_198859070), .Z(n_200759088));
	notech_ao4 i_141160390(.A(n_26648), .B(n_29669), .C(n_59095), .D(n_28110
		), .Z(n_200559086));
	notech_nor2 i_20091(.A(n_55508), .B(n_29536), .Z(n_101485291));
	notech_and3 i_5467347(.A(n_32656), .B(n_1869), .C(n_138785664), .Z(n_101785294
		));
	notech_ao4 i_53844(.A(n_101785294), .B(n_61103), .C(n_288827270), .D(n_26992
		), .Z(\nbus_11351[0] ));
	notech_ao3 i_5667345(.A(n_3821), .B(n_26992), .C(n_26993), .Z(n_101985296
		));
	notech_and3 i_5567346(.A(n_32446), .B(n_58740), .C(n_57308), .Z(n_102185298
		));
	notech_ao4 i_48535(.A(n_102185298), .B(n_135041965), .C(n_101985296), .D
		(n_29793), .Z(n_13782));
	notech_and4 i_5767344(.A(n_32434), .B(n_32432), .C(n_32446), .D(n_58740)
		, .Z(n_102385300));
	notech_ao4 i_48930(.A(n_6258839), .B(n_27052), .C(n_102385300), .D(n_61103
		), .Z(n_14391));
	notech_and3 i_8867313(.A(n_60117), .B(n_60303), .C(n_7148928), .Z(n_102485301
		));
	notech_or4 i_48487(.A(n_26993), .B(n_26612), .C(n_102485301), .D(n_3819)
		, .Z(n_13726));
	notech_or4 i_9467307(.A(n_61130), .B(n_60257), .C(n_29793), .D(n_138785664
		), .Z(n_102585302));
	notech_nand2 i_48178(.A(n_139285669), .B(n_102585302), .Z(\nbus_11299[0] 
		));
	notech_nand2 i_52677(.A(n_46630), .B(n_26992), .Z(n_19896));
	notech_or2 i_52706(.A(n_349480995), .B(n_3819), .Z(n_19928));
	notech_or4 i_49041(.A(n_27106), .B(n_61130), .C(n_60303), .D(n_19928), .Z
		(\nbus_11308[0] ));
	notech_ao4 i_4067361(.A(n_2883), .B(n_2877), .C(n_59460), .D(n_27896), .Z
		(n_102785304));
	notech_or4 i_28767134(.A(n_60964), .B(n_60953), .C(n_305047803), .D(n_62850
		), .Z(n_102885305));
	notech_or4 i_28867133(.A(n_2875), .B(n_28081), .C(n_32443), .D(n_60868),
		 .Z(n_102985306));
	notech_or2 i_28967132(.A(n_102785304), .B(n_59413), .Z(n_103085307));
	notech_or4 i_29767124(.A(n_61130), .B(n_60257), .C(n_29793), .D(n_103485311
		), .Z(n_103385310));
	notech_and4 i_6667335(.A(n_329163508), .B(n_112441739), .C(n_103085307),
		 .D(n_139685673), .Z(n_103485311));
	notech_ao4 i_6567336(.A(n_32548), .B(n_139985676), .C(n_26999), .D(n_319791626
		), .Z(n_103585312));
	notech_or4 i_29867123(.A(n_32579), .B(n_32559), .C(n_103585312), .D(n_29793
		), .Z(n_103685313));
	notech_or4 i_29967122(.A(n_32476), .B(n_25397), .C(n_29793), .D(n_56570)
		, .Z(n_103785314));
	notech_nand3 i_56534(.A(n_103785314), .B(n_103685313), .C(n_103385310), 
		.Z(\nbus_11380[16] ));
	notech_and3 i_30467117(.A(n_60054), .B(n_103985316), .C(n_1894), .Z(n_103885315
		));
	notech_or4 i_4267359(.A(n_4958709), .B(tss_esp0), .C(n_62870), .D(n_32655
		), .Z(n_103985316));
	notech_or4 i_10641(.A(n_61130), .B(n_60257), .C(n_29793), .D(n_103885315
		), .Z(n_104085317));
	notech_or4 i_30767114(.A(n_27069), .B(n_29655), .C(n_29793), .D(n_27068)
		, .Z(n_104185318));
	notech_nand2 i_52834(.A(n_104085317), .B(n_104185318), .Z(\nbus_11346[0] 
		));
	notech_nao3 i_31167110(.A(n_104685323), .B(n_61560), .C(n_61109), .Z(n_104285319
		));
	notech_nand2 i_56415(.A(n_140585682), .B(n_104285319), .Z(\nbus_11378[0] 
		));
	notech_nand3 i_32667096(.A(n_60117), .B(n_60303), .C(n_104685323), .Z(n_104585322
		));
	notech_nand3 i_3067370(.A(n_32434), .B(n_2419), .C(n_53745), .Z(n_104685323
		));
	notech_or4 i_32567097(.A(n_19057), .B(n_32579), .C(n_317791646), .D(n_60303
		), .Z(n_104785324));
	notech_and4 i_54290(.A(n_58683), .B(n_26992), .C(n_104785324), .D(n_104585322
		), .Z(\nbus_11357[0] ));
	notech_or4 i_33067092(.A(n_61109), .B(n_310587379), .C(n_59424), .D(n_32747
		), .Z(n_104885325));
	notech_nand2 i_53981(.A(n_26992), .B(n_104885325), .Z(n_22030));
	notech_and2 i_34767078(.A(write_ack), .B(n_105085327), .Z(n_104985326)
		);
	notech_nand2 i_6767334(.A(n_57285), .B(n_318591638), .Z(n_105085327));
	notech_nor2 i_34567079(.A(n_27063), .B(n_58683), .Z(n_105185328));
	notech_or4 i_49250(.A(n_105185328), .B(n_61130), .C(n_140985686), .D(n_104985326
		), .Z(n_14840));
	notech_nao3 i_35267073(.A(n_60117), .B(n_60298), .C(n_1880), .Z(n_105285329
		));
	notech_nand3 i_49205(.A(n_53731), .B(n_187610088), .C(n_105285329), .Z(n_14789
		));
	notech_nand2 i_48057(.A(n_187410086), .B(n_26992), .Z(\nbus_11298[0] )
		);
	notech_nao3 i_35767068(.A(n_60113), .B(n_60298), .C(n_30987), .Z(n_105385330
		));
	notech_or4 i_35667069(.A(n_27501), .B(n_3893), .C(\opcode[0] ), .D(n_32730
		), .Z(n_105485331));
	notech_nand3 i_47880(.A(n_26992), .B(n_105485331), .C(n_105385330), .Z(n_12360
		));
	notech_and4 i_42767000(.A(n_59408), .B(n_59398), .C(n_59286), .D(imm[16]
		), .Z(n_105585332));
	notech_and4 i_42966998(.A(n_59408), .B(n_59398), .C(n_59286), .D(imm[17]
		), .Z(n_105685333));
	notech_and4 i_43166996(.A(n_59408), .B(n_59398), .C(n_59286), .D(imm[18]
		), .Z(n_105785334));
	notech_and4 i_43366994(.A(n_59408), .B(n_59398), .C(n_59286), .D(imm[19]
		), .Z(n_105885335));
	notech_and4 i_43566992(.A(n_59408), .B(n_59398), .C(n_59286), .D(imm[20]
		), .Z(n_105985336));
	notech_and4 i_43766990(.A(n_59408), .B(n_59398), .C(n_59286), .D(imm[21]
		), .Z(n_106085337));
	notech_and4 i_44166986(.A(n_59408), .B(n_59393), .C(n_59286), .D(imm[23]
		), .Z(n_106185338));
	notech_and4 i_44366984(.A(n_59408), .B(n_59393), .C(n_59286), .D(imm[24]
		), .Z(n_106285339));
	notech_and4 i_44566982(.A(n_59408), .B(n_59393), .C(n_59286), .D(imm[28]
		), .Z(n_106385340));
	notech_and4 i_44766980(.A(n_59408), .B(n_59393), .C(n_59286), .D(imm[29]
		), .Z(n_106485341));
	notech_ao4 i_44966978(.A(n_4958709), .B(n_323084221), .C(n_60894), .D(n_27509
		), .Z(n_106585342));
	notech_ao4 i_4467357(.A(n_62844), .B(n_62792), .C(n_59413), .D(mul64[7])
		, .Z(n_106985346));
	notech_or4 i_47666951(.A(n_143685713), .B(n_143385710), .C(n_144585722),
		 .D(n_143085707), .Z(n_107085347));
	notech_ao4 i_367392(.A(n_60894), .B(mul64[31]), .C(n_62792), .D(n_60910)
		, .Z(n_107185348));
	notech_nao3 i_47466953(.A(n_5187), .B(mul64[31]), .C(n_60894), .Z(n_107285349
		));
	notech_nao3 i_47566952(.A(n_5183), .B(mul64[7]), .C(n_59413), .Z(n_107385350
		));
	notech_nand2 i_47366954(.A(n_5179), .B(n_27007), .Z(n_107485351));
	notech_or4 i_51566912(.A(n_2875), .B(n_28081), .C(n_2877), .D(n_107885355
		), .Z(n_107785354));
	notech_and4 i_7067331(.A(n_107085347), .B(n_107385350), .C(n_107285349),
		 .D(n_107485351), .Z(n_107885355));
	notech_mux2 i_6967332(.S(mul64[15]), .A(n_30202), .B(n_30201), .Z(n_107985356
		));
	notech_nand2 i_7661(.A(n_107785354), .B(n_145185728), .Z(n_12393));
	notech_ao4 i_3215669(.A(n_62041235), .B(n_28123), .C(n_317887452), .D(n_28418
		), .Z(n_22875));
	notech_ao4 i_3115668(.A(n_62041235), .B(n_28121), .C(n_317887452), .D(n_28417
		), .Z(n_22870));
	notech_ao4 i_3015667(.A(n_62041235), .B(n_28118), .C(n_317887452), .D(n_28416
		), .Z(n_22865));
	notech_ao4 i_2915666(.A(n_62041235), .B(n_28117), .C(n_317887452), .D(n_28415
		), .Z(n_22860));
	notech_ao4 i_2815665(.A(n_62041235), .B(n_28116), .C(n_317887452), .D(n_28414
		), .Z(n_22855));
	notech_ao4 i_2715664(.A(n_62041235), .B(n_28115), .C(n_317887452), .D(n_28413
		), .Z(n_22850));
	notech_ao4 i_2615663(.A(n_62041235), .B(n_28114), .C(n_317887452), .D(n_28412
		), .Z(n_22845));
	notech_ao4 i_2515662(.A(n_62041235), .B(n_28113), .C(n_317887452), .D(n_28411
		), .Z(n_22840));
	notech_ao4 i_2415661(.A(n_62041235), .B(n_28112), .C(n_317887452), .D(n_28410
		), .Z(n_22835));
	notech_ao4 i_2315660(.A(n_62041235), .B(n_28111), .C(n_317887452), .D(n_28409
		), .Z(n_22830));
	notech_ao4 i_2215659(.A(n_62041235), .B(n_28110), .C(n_317887452), .D(n_28408
		), .Z(n_22825));
	notech_ao4 i_2115658(.A(n_62041235), .B(n_28109), .C(n_317887452), .D(n_28407
		), .Z(n_22820));
	notech_ao4 i_2015657(.A(n_62041235), .B(n_28108), .C(n_317887452), .D(n_28406
		), .Z(n_22815));
	notech_ao4 i_1915656(.A(n_62041235), .B(n_28107), .C(n_317887452), .D(n_28405
		), .Z(n_22810));
	notech_ao4 i_1815655(.A(n_54409), .B(n_28106), .C(n_54400), .D(n_28404),
		 .Z(n_22805));
	notech_ao4 i_1715654(.A(n_54409), .B(n_28105), .C(n_54400), .D(n_28403),
		 .Z(n_22800));
	notech_ao4 i_1615653(.A(n_54409), .B(n_28104), .C(n_54400), .D(n_28402),
		 .Z(n_22795));
	notech_ao4 i_1515652(.A(n_54409), .B(n_28103), .C(n_54400), .D(n_28401),
		 .Z(n_22790));
	notech_ao4 i_1415651(.A(n_54409), .B(n_28102), .C(n_54400), .D(n_28400),
		 .Z(n_22785));
	notech_ao4 i_1315650(.A(n_54409), .B(n_28101), .C(n_54400), .D(n_28399),
		 .Z(n_22780));
	notech_ao4 i_1215649(.A(n_54409), .B(n_28100), .C(n_54400), .D(n_28398),
		 .Z(n_22775));
	notech_ao4 i_1115648(.A(n_54409), .B(n_28099), .C(n_54400), .D(n_28397),
		 .Z(n_22770));
	notech_ao4 i_1015647(.A(n_54409), .B(n_28098), .C(n_54400), .D(n_28396),
		 .Z(n_22765));
	notech_ao4 i_915646(.A(n_54409), .B(n_28097), .C(n_54400), .D(n_28395), 
		.Z(n_22760));
	notech_ao4 i_815645(.A(n_54409), .B(n_28096), .C(n_317887452), .D(n_28394
		), .Z(n_22755));
	notech_ao4 i_715644(.A(n_54409), .B(n_28095), .C(n_54400), .D(n_28393), 
		.Z(n_22750));
	notech_ao4 i_515642(.A(n_54409), .B(n_28093), .C(n_54400), .D(n_28391), 
		.Z(n_22740));
	notech_ao4 i_415641(.A(n_28092), .B(n_54409), .C(n_28390), .D(n_54400), 
		.Z(n_22735));
	notech_ao4 i_215639(.A(n_54409), .B(n_28090), .C(n_54400), .D(n_28388), 
		.Z(n_22725));
	notech_ao4 i_115638(.A(n_54409), .B(n_28089), .C(n_54400), .D(n_28387), 
		.Z(n_22720));
	notech_ao4 i_223101(.A(n_209986373), .B(n_59241), .C(n_57440), .D(n_56010
		), .Z(n_16495));
	notech_ao4 i_123100(.A(n_209986373), .B(n_59187), .C(n_56028), .D(n_57440
		), .Z(n_16489));
	notech_ao4 i_74066687(.A(n_56199), .B(n_106485341), .C(n_179382794), .D(n_55191
		), .Z(n_114785424));
	notech_or2 i_21067413(.A(n_106485341), .B(n_56199), .Z(\nbus_11317[29] )
		);
	notech_nand2 i_3012947(.A(n_145885735), .B(n_27008), .Z(n_26093));
	notech_ao4 i_75766670(.A(n_56199), .B(n_106385340), .C(n_179382794), .D(n_55191
		), .Z(n_115685433));
	notech_or2 i_20767414(.A(n_106385340), .B(n_56199), .Z(\nbus_11317[28] )
		);
	notech_nand2 i_2912946(.A(n_146585742), .B(n_27009), .Z(n_26088));
	notech_ao4 i_77466653(.A(n_56199), .B(n_106285339), .C(n_179382794), .D(n_55191
		), .Z(n_116585442));
	notech_or2 i_20667415(.A(n_106285339), .B(n_56199), .Z(\nbus_11317[24] )
		);
	notech_nand2 i_2512942(.A(n_147285749), .B(n_27010), .Z(n_26068));
	notech_ao4 i_79166636(.A(n_56199), .B(n_106185338), .C(n_179382794), .D(n_55191
		), .Z(n_117485451));
	notech_or2 i_19967416(.A(n_106185338), .B(n_56199), .Z(\nbus_11317[23] )
		);
	notech_nand2 i_2412941(.A(n_147985756), .B(n_27012), .Z(n_26063));
	notech_ao4 i_82566602(.A(n_56204), .B(n_106085337), .C(n_179382794), .D(n_55191
		), .Z(n_118385460));
	notech_or2 i_20967418(.A(n_106085337), .B(n_56204), .Z(\nbus_11317[21] )
		);
	notech_nand2 i_2212939(.A(n_148685763), .B(n_27013), .Z(n_26053));
	notech_ao4 i_84266585(.A(n_56204), .B(n_105985336), .C(n_179382794), .D(n_26781
		), .Z(n_119285469));
	notech_or2 i_20567419(.A(n_105985336), .B(n_56204), .Z(\nbus_11317[20] )
		);
	notech_nand2 i_2112938(.A(n_149385770), .B(n_27014), .Z(n_26048));
	notech_ao4 i_85966568(.A(n_56204), .B(n_105885335), .C(n_179382794), .D(n_55191
		), .Z(n_120185478));
	notech_or2 i_19867420(.A(n_105885335), .B(n_56204), .Z(\nbus_11317[19] )
		);
	notech_nand2 i_2012937(.A(n_150085777), .B(n_27016), .Z(n_26043));
	notech_ao4 i_87666551(.A(n_56204), .B(n_105785334), .C(n_179382794), .D(n_55191
		), .Z(n_121085487));
	notech_or2 i_158067421(.A(n_105785334), .B(n_56204), .Z(\nbus_11317[18] 
		));
	notech_nand2 i_1912936(.A(n_150785784), .B(n_27017), .Z(n_26038));
	notech_ao4 i_89366534(.A(n_56204), .B(n_105685333), .C(n_179382794), .D(n_55191
		), .Z(n_121985496));
	notech_or2 i_157967422(.A(n_105685333), .B(n_56204), .Z(\nbus_11317[17] 
		));
	notech_nand2 i_1812935(.A(n_151485791), .B(n_27018), .Z(n_26033));
	notech_ao4 i_91066517(.A(n_105585332), .B(n_56204), .C(n_179382794), .D(n_55191
		), .Z(n_122885505));
	notech_or2 i_20467423(.A(n_105585332), .B(n_56204), .Z(\nbus_11317[16] )
		);
	notech_nand2 i_1712934(.A(n_152185798), .B(n_27021), .Z(n_26028));
	notech_nand2 i_126466164(.A(write_data_33[31]), .B(n_60257), .Z(n_124185518
		));
	notech_nand3 i_3218837(.A(n_152385800), .B(n_152285799), .C(n_124185518)
		, .Z(n_25859));
	notech_nand2 i_127366155(.A(write_data_33[30]), .B(n_60257), .Z(n_124685523
		));
	notech_nand3 i_3118836(.A(n_152685803), .B(n_152585802), .C(n_124685523)
		, .Z(n_25854));
	notech_nand2 i_128266146(.A(write_data_33[29]), .B(n_60257), .Z(n_125185528
		));
	notech_nand3 i_3018835(.A(n_152985806), .B(n_152885805), .C(n_125185528)
		, .Z(n_25849));
	notech_nand2 i_129166137(.A(write_data_33[28]), .B(n_60257), .Z(n_125685533
		));
	notech_nand3 i_2918834(.A(n_153285809), .B(n_153185808), .C(n_125685533)
		, .Z(n_25844));
	notech_nand2 i_130066128(.A(write_data_33[27]), .B(n_60257), .Z(n_126185538
		));
	notech_nand3 i_2818833(.A(n_153585812), .B(n_153485811), .C(n_126185538)
		, .Z(n_25839));
	notech_nand2 i_130966119(.A(write_data_33[26]), .B(n_60257), .Z(n_126685543
		));
	notech_nand3 i_2718832(.A(n_153885815), .B(n_153785814), .C(n_126685543)
		, .Z(n_25834));
	notech_nand2 i_131866110(.A(write_data_33[25]), .B(n_60257), .Z(n_127185548
		));
	notech_nand3 i_2618831(.A(n_154185818), .B(n_154085817), .C(n_127185548)
		, .Z(n_25829));
	notech_nand2 i_132766101(.A(write_data_33[24]), .B(n_60257), .Z(n_127685553
		));
	notech_nand3 i_2518830(.A(n_154485821), .B(n_154385820), .C(n_127685553)
		, .Z(n_25824));
	notech_nand2 i_133666092(.A(write_data_33[23]), .B(n_60257), .Z(n_128185558
		));
	notech_nand3 i_2418829(.A(n_154785824), .B(n_154685823), .C(n_128185558)
		, .Z(n_25819));
	notech_nand2 i_134666083(.A(write_data_33[22]), .B(n_60252), .Z(n_128685563
		));
	notech_nand3 i_2318828(.A(n_155085827), .B(n_154985826), .C(n_128685563)
		, .Z(n_25814));
	notech_nand2 i_135566074(.A(write_data_33[21]), .B(n_60252), .Z(n_129185568
		));
	notech_nand3 i_2218827(.A(n_155385830), .B(n_155285829), .C(n_129185568)
		, .Z(n_25809));
	notech_nand2 i_136466065(.A(write_data_33[20]), .B(n_60252), .Z(n_129685573
		));
	notech_nand3 i_2118826(.A(n_155685833), .B(n_155585832), .C(n_129685573)
		, .Z(n_25804));
	notech_nand2 i_137366056(.A(write_data_33[19]), .B(n_60257), .Z(n_130185578
		));
	notech_nand3 i_2018825(.A(n_155985836), .B(n_155885835), .C(n_130185578)
		, .Z(n_25799));
	notech_nand2 i_138266047(.A(write_data_33[18]), .B(n_60257), .Z(n_130685583
		));
	notech_nand3 i_1918824(.A(n_156285839), .B(n_156185838), .C(n_130685583)
		, .Z(n_25794));
	notech_nand2 i_139166038(.A(write_data_33[17]), .B(n_60257), .Z(n_131185588
		));
	notech_nand3 i_1818823(.A(n_156585842), .B(n_156485841), .C(n_131185588)
		, .Z(n_25789));
	notech_nand2 i_140066029(.A(write_data_33[16]), .B(n_60257), .Z(n_131685593
		));
	notech_nand3 i_1718822(.A(n_156885845), .B(n_156785844), .C(n_131685593)
		, .Z(n_25784));
	notech_nand2 i_140966020(.A(write_data_33[15]), .B(n_60257), .Z(n_132185598
		));
	notech_nand3 i_1618821(.A(n_157185848), .B(n_157085847), .C(n_132185598)
		, .Z(n_25779));
	notech_nand2 i_141866011(.A(write_data_33[14]), .B(n_60171), .Z(n_132685603
		));
	notech_nand3 i_1518820(.A(n_157485851), .B(n_157385850), .C(n_132685603)
		, .Z(n_25774));
	notech_nand2 i_142766002(.A(write_data_33[13]), .B(n_60171), .Z(n_133185608
		));
	notech_nand3 i_1418819(.A(n_157785854), .B(n_157685853), .C(n_133185608)
		, .Z(n_25769));
	notech_nand2 i_143665993(.A(write_data_33[12]), .B(n_60171), .Z(n_133685613
		));
	notech_nand3 i_1318818(.A(n_158085857), .B(n_157985856), .C(n_133685613)
		, .Z(n_25764));
	notech_nand2 i_144565984(.A(write_data_33[11]), .B(n_60171), .Z(n_134185618
		));
	notech_nand3 i_1218817(.A(n_158385860), .B(n_158285859), .C(n_134185618)
		, .Z(n_25759));
	notech_nand2 i_145465975(.A(write_data_33[10]), .B(n_60171), .Z(n_134685623
		));
	notech_nand3 i_1118816(.A(n_158685863), .B(n_158585862), .C(n_134685623)
		, .Z(n_25754));
	notech_nand2 i_146365966(.A(write_data_33[9]), .B(n_60171), .Z(n_135185628
		));
	notech_nand3 i_1018815(.A(n_158985866), .B(n_158885865), .C(n_135185628)
		, .Z(n_25749));
	notech_nand2 i_147265957(.A(write_data_33[8]), .B(n_60171), .Z(n_135685633
		));
	notech_nand3 i_918814(.A(n_159285869), .B(n_159185868), .C(n_135685633),
		 .Z(n_25744));
	notech_nand2 i_148165948(.A(write_data_33[7]), .B(n_60171), .Z(n_136185638
		));
	notech_nand3 i_818813(.A(n_159585872), .B(n_159485871), .C(n_136185638),
		 .Z(n_25739));
	notech_nand2 i_149065939(.A(write_data_33[6]), .B(n_60171), .Z(n_136685643
		));
	notech_nand3 i_718812(.A(n_159885875), .B(n_159785874), .C(n_136685643),
		 .Z(n_25734));
	notech_nand2 i_150865921(.A(write_data_33[4]), .B(n_60171), .Z(n_137185648
		));
	notech_nand3 i_518810(.A(n_160185878), .B(n_160085877), .C(n_137185648),
		 .Z(n_25724));
	notech_nand2 i_151765912(.A(write_data_33[3]), .B(n_60171), .Z(n_137685653
		));
	notech_nand3 i_418809(.A(n_160485881), .B(n_160385880), .C(n_137685653),
		 .Z(n_25719));
	notech_nand2 i_153565894(.A(write_data_33[1]), .B(n_60184), .Z(n_138185658
		));
	notech_nand3 i_218807(.A(n_160785884), .B(n_160685883), .C(n_138185658),
		 .Z(n_25709));
	notech_nand2 i_154465885(.A(write_data_33[0]), .B(n_60184), .Z(n_138685663
		));
	notech_nand3 i_118806(.A(n_161085887), .B(n_160985886), .C(n_138685663),
		 .Z(n_25704));
	notech_and2 i_2767373(.A(n_60054), .B(n_57912), .Z(n_138785664));
	notech_or4 i_3967362(.A(n_32580), .B(n_32559), .C(n_61130), .D(n_29793),
		 .Z(n_139185668));
	notech_ao4 i_9667305(.A(n_5968810), .B(n_29793), .C(n_139185668), .D(n_317791646
		), .Z(n_139285669));
	notech_and4 i_29167130(.A(n_1894), .B(n_1895), .C(n_102885305), .D(n_102985306
		), .Z(n_139685673));
	notech_or4 i_29667125(.A(n_3812), .B(n_5380), .C(n_32565), .D(n_19043), 
		.Z(n_139985676));
	notech_ao4 i_31367108(.A(n_32405), .B(n_139185668), .C(n_58683), .D(n_29793
		), .Z(n_140585682));
	notech_nand2 i_34867077(.A(n_187310085), .B(n_53739), .Z(n_140985686));
	notech_or4 i_2667374(.A(n_60969), .B(n_60958), .C(n_61109), .D(n_60910),
		 .Z(n_10157));
	notech_or4 i_49766930(.A(mul64[42]), .B(mul64[43]), .C(mul64[41]), .D(mul64
		[40]), .Z(n_141885695));
	notech_or4 i_49866929(.A(mul64[46]), .B(mul64[47]), .C(mul64[44]), .D(mul64
		[45]), .Z(n_142185698));
	notech_or4 i_49966928(.A(mul64[50]), .B(mul64[51]), .C(mul64[48]), .D(mul64
		[49]), .Z(n_142585702));
	notech_or4 i_50066927(.A(mul64[54]), .B(mul64[55]), .C(mul64[52]), .D(mul64
		[53]), .Z(n_142885705));
	notech_or4 i_50866919(.A(n_142885705), .B(n_142585702), .C(n_142185698),
		 .D(n_141885695), .Z(n_143085707));
	notech_or4 i_50166926(.A(mul64[58]), .B(mul64[59]), .C(mul64[56]), .D(mul64
		[57]), .Z(n_143385710));
	notech_or4 i_50266925(.A(mul64[62]), .B(mul64[63]), .C(mul64[60]), .D(mul64
		[61]), .Z(n_143685713));
	notech_and4 i_49566932(.A(n_30197), .B(n_30198), .C(n_30196), .D(n_30199
		), .Z(n_144085717));
	notech_or4 i_49666931(.A(mul64[38]), .B(mul64[37]), .C(mul64[39]), .D(mul64
		[36]), .Z(n_144385720));
	notech_nao3 i_50766920(.A(n_27040), .B(n_144085717), .C(n_107185348), .Z
		(n_144585722));
	notech_ao4 i_51766910(.A(n_1900), .B(n_107985356), .C(n_1899), .D(n_30202
		), .Z(n_145185728));
	notech_nand2 i_37467399(.A(n_19014), .B(n_60184), .Z(n_62041235));
	notech_ao4 i_74166686(.A(n_55200), .B(n_30203), .C(n_328184272), .D(n_29083
		), .Z(n_145285729));
	notech_ao4 i_74266685(.A(n_55220), .B(n_57815), .C(n_55209), .D(n_30204)
		, .Z(n_145385730));
	notech_ao4 i_74366684(.A(n_55632), .B(n_30205), .C(n_55229), .D(nbus_11295
		[29]), .Z(n_145585732));
	notech_ao4 i_74466683(.A(n_52741142), .B(n_28118), .C(n_58773), .D(n_29114
		), .Z(n_145685733));
	notech_and4 i_74766680(.A(n_145685733), .B(n_145585732), .C(n_145385730)
		, .D(n_145285729), .Z(n_145885735));
	notech_ao4 i_75866669(.A(n_55200), .B(n_30206), .C(n_328184272), .D(n_29082
		), .Z(n_145985736));
	notech_ao4 i_75966668(.A(n_55220), .B(\nbus_11365[28] ), .C(n_55209), .D
		(n_30207), .Z(n_146085737));
	notech_ao4 i_76066667(.A(n_55632), .B(n_30208), .C(n_55229), .D(nbus_11295
		[28]), .Z(n_146285739));
	notech_ao4 i_76166666(.A(n_52741142), .B(n_28117), .C(n_58773), .D(n_29113
		), .Z(n_146385740));
	notech_and4 i_76466663(.A(n_146385740), .B(n_146285739), .C(n_146085737)
		, .D(n_145985736), .Z(n_146585742));
	notech_ao4 i_77566652(.A(n_55200), .B(n_30209), .C(n_328184272), .D(n_29078
		), .Z(n_146685743));
	notech_ao4 i_77666651(.A(n_55229), .B(nbus_11295[24]), .C(n_55209), .D(n_30210
		), .Z(n_146785744));
	notech_ao4 i_77766650(.A(n_58773), .B(n_29110), .C(n_55632), .D(n_30211)
		, .Z(n_146985746));
	notech_ao4 i_77866649(.A(n_28113), .B(n_52741142), .C(n_55220), .D(n_57761
		), .Z(n_147085747));
	notech_and4 i_78166646(.A(n_147085747), .B(n_146985746), .C(n_146785744)
		, .D(n_146685743), .Z(n_147285749));
	notech_ao4 i_79266635(.A(n_55200), .B(n_30212), .C(n_328184272), .D(n_29077
		), .Z(n_147385750));
	notech_ao4 i_79366634(.A(n_55229), .B(nbus_11295[23]), .C(n_55209), .D(n_30213
		), .Z(n_147485751));
	notech_ao4 i_79466633(.A(n_58773), .B(n_29109), .C(n_55632), .D(n_30214)
		, .Z(n_147685753));
	notech_ao4 i_79566632(.A(n_52741142), .B(n_28112), .C(n_55220), .D(n_57751
		), .Z(n_147785754));
	notech_and4 i_79866629(.A(n_147785754), .B(n_147685753), .C(n_147485751)
		, .D(n_147385750), .Z(n_147985756));
	notech_ao4 i_82666601(.A(n_55200), .B(n_30215), .C(n_328184272), .D(n_29075
		), .Z(n_148085757));
	notech_ao4 i_82766600(.A(n_53341148), .B(nbus_11295[21]), .C(n_55209), .D
		(n_30216), .Z(n_148185758));
	notech_ao4 i_82866599(.A(n_58773), .B(n_29107), .C(n_58768), .D(n_30217)
		, .Z(n_148385760));
	notech_ao4 i_82966598(.A(n_52741142), .B(n_28110), .C(n_55220), .D(n_57733
		), .Z(n_148485761));
	notech_and4 i_83266595(.A(n_148485761), .B(n_148385760), .C(n_148185758)
		, .D(n_148085757), .Z(n_148685763));
	notech_ao4 i_84366584(.A(n_55200), .B(n_30218), .C(n_328184272), .D(n_29074
		), .Z(n_148785764));
	notech_ao4 i_84466583(.A(n_55220), .B(n_57720), .C(n_55209), .D(n_30219)
		, .Z(n_148885765));
	notech_ao4 i_84566582(.A(n_55632), .B(n_30220), .C(n_55229), .D(nbus_11295
		[20]), .Z(n_149085767));
	notech_ao4 i_84666581(.A(n_52741142), .B(n_28109), .C(n_58773), .D(n_29106
		), .Z(n_149185768));
	notech_and4 i_84966578(.A(n_149185768), .B(n_149085767), .C(n_148885765)
		, .D(n_148785764), .Z(n_149385770));
	notech_ao4 i_86066567(.A(n_55200), .B(n_30221), .C(n_328184272), .D(n_29073
		), .Z(n_149485771));
	notech_ao4 i_86166566(.A(n_55229), .B(nbus_11295[19]), .C(n_55209), .D(n_30222
		), .Z(n_149585772));
	notech_ao4 i_86266565(.A(n_58773), .B(n_29105), .C(n_55632), .D(n_30223)
		, .Z(n_149785774));
	notech_ao4 i_86366564(.A(n_52741142), .B(n_28108), .C(n_55220), .D(n_57707
		), .Z(n_149885775));
	notech_and4 i_86666561(.A(n_149885775), .B(n_149785774), .C(n_149585772)
		, .D(n_149485771), .Z(n_150085777));
	notech_ao4 i_87766550(.A(n_55200), .B(n_30224), .C(n_328184272), .D(n_29072
		), .Z(n_150185778));
	notech_ao4 i_87866549(.A(n_55229), .B(nbus_11295[18]), .C(n_55209), .D(n_30225
		), .Z(n_150285779));
	notech_ao4 i_87966548(.A(n_58773), .B(n_29104), .C(n_55632), .D(n_30226)
		, .Z(n_150485781));
	notech_ao4 i_88066547(.A(n_52741142), .B(n_28107), .C(n_55220), .D(n_57698
		), .Z(n_150585782));
	notech_and4 i_88366544(.A(n_150585782), .B(n_150485781), .C(n_150285779)
		, .D(n_150185778), .Z(n_150785784));
	notech_ao4 i_89466533(.A(n_55200), .B(n_30227), .C(n_328184272), .D(n_29070
		), .Z(n_150885785));
	notech_ao4 i_89566532(.A(n_55229), .B(nbus_11295[17]), .C(n_55209), .D(n_30228
		), .Z(n_150985786));
	notech_ao4 i_89666531(.A(n_58773), .B(n_29103), .C(n_55632), .D(n_30229)
		, .Z(n_151185788));
	notech_ao4 i_89766530(.A(n_52741142), .B(n_28106), .C(n_55220), .D(n_57689
		), .Z(n_151285789));
	notech_and4 i_90066527(.A(n_151285789), .B(n_151185788), .C(n_150985786)
		, .D(n_150885785), .Z(n_151485791));
	notech_ao4 i_91166516(.A(n_55200), .B(n_30230), .C(n_328184272), .D(n_29069
		), .Z(n_151585792));
	notech_ao4 i_91266515(.A(n_55229), .B(nbus_11295[16]), .C(n_55209), .D(n_30231
		), .Z(n_151685793));
	notech_ao4 i_91366514(.A(n_58773), .B(n_29102), .C(n_55632), .D(n_30232)
		, .Z(n_151885795));
	notech_ao4 i_91466513(.A(n_52741142), .B(n_28105), .C(n_55220), .D(n_57680
		), .Z(n_151985796));
	notech_and4 i_91766510(.A(n_151985796), .B(n_151885795), .C(n_151685793)
		, .D(n_151585792), .Z(n_152185798));
	notech_ao4 i_126666162(.A(n_318291641), .B(n_57837), .C(n_318391640), .D
		(nbus_11295[31]), .Z(n_152285799));
	notech_ao4 i_126566163(.A(n_315391670), .B(n_27893), .C(n_59142), .D(n_28482
		), .Z(n_152385800));
	notech_ao4 i_127566153(.A(n_318291641), .B(n_55929), .C(n_318391640), .D
		(nbus_11295[30]), .Z(n_152585802));
	notech_ao4 i_127466154(.A(n_315391670), .B(n_27892), .C(n_59142), .D(n_28481
		), .Z(n_152685803));
	notech_ao4 i_128466144(.A(n_318291641), .B(n_55956), .C(n_318391640), .D
		(nbus_11295[29]), .Z(n_152885805));
	notech_ao4 i_128366145(.A(n_315391670), .B(n_27891), .C(n_59142), .D(n_28480
		), .Z(n_152985806));
	notech_ao4 i_129366135(.A(n_318291641), .B(n_55974), .C(n_318391640), .D
		(nbus_11295[28]), .Z(n_153185808));
	notech_ao4 i_129266136(.A(n_315391670), .B(n_27890), .C(n_59142), .D(n_28479
		), .Z(n_153285809));
	notech_ao4 i_130266126(.A(n_318291641), .B(n_55938), .C(n_318391640), .D
		(n_57881), .Z(n_153485811));
	notech_ao4 i_130166127(.A(n_315391670), .B(n_27889), .C(n_59147), .D(n_28478
		), .Z(n_153585812));
	notech_ao4 i_131166117(.A(n_318291641), .B(n_55947), .C(n_318391640), .D
		(nbus_11295[26]), .Z(n_153785814));
	notech_ao4 i_131066118(.A(n_315391670), .B(n_27888), .C(n_59147), .D(n_28477
		), .Z(n_153885815));
	notech_ao4 i_132066108(.A(n_318291641), .B(n_55965), .C(n_318391640), .D
		(nbus_11295[25]), .Z(n_154085817));
	notech_ao4 i_131966109(.A(n_315391670), .B(n_27887), .C(n_59142), .D(n_28476
		), .Z(n_154185818));
	notech_ao4 i_132966099(.A(n_318291641), .B(n_56475), .C(n_318391640), .D
		(nbus_11295[24]), .Z(n_154385820));
	notech_ao4 i_132866100(.A(n_315391670), .B(n_27886), .C(n_59142), .D(n_28475
		), .Z(n_154485821));
	notech_ao4 i_133866090(.A(n_318291641), .B(n_56347), .C(n_318391640), .D
		(nbus_11295[23]), .Z(n_154685823));
	notech_ao4 i_133766091(.A(n_315391670), .B(n_27884), .C(n_59142), .D(n_28474
		), .Z(n_154785824));
	notech_ao4 i_134866081(.A(n_318291641), .B(n_56338), .C(n_318391640), .D
		(nbus_11295[22]), .Z(n_154985826));
	notech_ao4 i_134766082(.A(n_315391670), .B(n_27883), .C(n_59142), .D(n_28473
		), .Z(n_155085827));
	notech_ao4 i_135766072(.A(n_318291641), .B(n_56329), .C(n_318391640), .D
		(nbus_11295[21]), .Z(n_155285829));
	notech_ao4 i_135666073(.A(n_315391670), .B(n_27882), .C(n_59142), .D(n_28472
		), .Z(n_155385830));
	notech_ao4 i_136666063(.A(n_318291641), .B(n_56320), .C(n_318391640), .D
		(nbus_11295[20]), .Z(n_155585832));
	notech_ao4 i_136566064(.A(n_315391670), .B(n_27881), .C(n_59142), .D(n_28471
		), .Z(n_155685833));
	notech_ao4 i_137566054(.A(n_318291641), .B(n_56311), .C(n_318391640), .D
		(nbus_11295[19]), .Z(n_155885835));
	notech_ao4 i_137466055(.A(n_315391670), .B(n_27878), .C(n_59142), .D(n_28470
		), .Z(n_155985836));
	notech_ao4 i_138466045(.A(n_318291641), .B(n_56302), .C(n_318391640), .D
		(nbus_11295[18]), .Z(n_156185838));
	notech_ao4 i_138366046(.A(n_315391670), .B(n_27876), .C(n_59142), .D(n_28469
		), .Z(n_156285839));
	notech_ao4 i_139366036(.A(n_318291641), .B(n_56293), .C(n_318391640), .D
		(nbus_11295[17]), .Z(n_156485841));
	notech_ao4 i_139266037(.A(n_59133), .B(n_27875), .C(n_59142), .D(n_28468
		), .Z(n_156585842));
	notech_ao4 i_140266027(.A(n_59106), .B(\nbus_11358[16] ), .C(n_59115), .D
		(nbus_11295[16]), .Z(n_156785844));
	notech_ao4 i_140166028(.A(n_59133), .B(n_27874), .C(n_59142), .D(n_28467
		), .Z(n_156885845));
	notech_ao4 i_141166018(.A(n_59106), .B(\nbus_11358[15] ), .C(n_59115), .D
		(nbus_11295[15]), .Z(n_157085847));
	notech_ao4 i_141066019(.A(n_59133), .B(n_27873), .C(n_59142), .D(n_28466
		), .Z(n_157185848));
	notech_ao4 i_142066009(.A(n_59106), .B(n_56248), .C(n_59115), .D(nbus_11295
		[14]), .Z(n_157385850));
	notech_ao4 i_141966010(.A(n_59133), .B(n_27872), .C(n_59147), .D(n_28465
		), .Z(n_157485851));
	notech_ao4 i_142966000(.A(n_59106), .B(n_56230), .C(n_59115), .D(nbus_11295
		[13]), .Z(n_157685853));
	notech_ao4 i_142866001(.A(n_59133), .B(n_27871), .C(n_59147), .D(n_28464
		), .Z(n_157785854));
	notech_ao4 i_143865991(.A(n_59106), .B(n_56221), .C(n_59115), .D(nbus_11295
		[12]), .Z(n_157985856));
	notech_ao4 i_143765992(.A(n_59133), .B(n_27870), .C(n_59147), .D(n_28463
		), .Z(n_158085857));
	notech_ao4 i_144765982(.A(n_59106), .B(n_56181), .C(n_59115), .D(nbus_11295
		[11]), .Z(n_158285859));
	notech_ao4 i_144665983(.A(n_59133), .B(n_27869), .C(n_59147), .D(n_28462
		), .Z(n_158385860));
	notech_ao4 i_145665973(.A(n_59106), .B(n_56154), .C(n_59115), .D(nbus_11295
		[10]), .Z(n_158585862));
	notech_ao4 i_145565974(.A(n_59133), .B(n_27868), .C(n_59152), .D(n_28461
		), .Z(n_158685863));
	notech_ao4 i_146565964(.A(n_59106), .B(n_56136), .C(n_59115), .D(nbus_11295
		[9]), .Z(n_158885865));
	notech_ao4 i_146465965(.A(n_59133), .B(n_27867), .C(n_59152), .D(n_28460
		), .Z(n_158985866));
	notech_ao4 i_147465955(.A(n_59106), .B(\nbus_11358[8] ), .C(n_59115), .D
		(nbus_11295[8]), .Z(n_159185868));
	notech_ao4 i_147365956(.A(n_59133), .B(n_27866), .C(n_59147), .D(n_28459
		), .Z(n_159285869));
	notech_ao4 i_148365946(.A(n_59106), .B(n_56109), .C(n_59115), .D(nbus_11295
		[7]), .Z(n_159485871));
	notech_ao4 i_148265947(.A(n_59133), .B(n_27865), .C(n_59147), .D(n_28458
		), .Z(n_159585872));
	notech_ao4 i_149265937(.A(n_318291641), .B(\nbus_11358[6] ), .C(n_318391640
		), .D(nbus_11295[6]), .Z(n_159785874));
	notech_ao4 i_149165938(.A(n_59133), .B(n_27864), .C(n_59147), .D(n_28457
		), .Z(n_159885875));
	notech_ao4 i_151065919(.A(n_59106), .B(n_56064), .C(n_59115), .D(nbus_11295
		[4]), .Z(n_160085877));
	notech_ao4 i_150965920(.A(n_59133), .B(n_27862), .C(n_59147), .D(n_28455
		), .Z(n_160185878));
	notech_ao4 i_151965910(.A(n_59106), .B(\nbus_11358[3] ), .C(n_59115), .D
		(n_57909), .Z(n_160385880));
	notech_ao4 i_151865911(.A(n_59133), .B(n_27861), .C(n_59147), .D(n_28454
		), .Z(n_160485881));
	notech_ao4 i_153765892(.A(n_59106), .B(n_56010), .C(n_59115), .D(nbus_11295
		[1]), .Z(n_160685883));
	notech_ao4 i_153665893(.A(n_59133), .B(n_27859), .C(n_59147), .D(n_28452
		), .Z(n_160785884));
	notech_ao4 i_154665883(.A(n_59106), .B(\nbus_11358[0] ), .C(n_59115), .D
		(n_59717), .Z(n_160985886));
	notech_ao4 i_154565884(.A(n_59133), .B(n_27858), .C(n_59147), .D(n_28451
		), .Z(n_161085887));
	notech_nao3 i_36064509(.A(n_2885), .B(n_106585342), .C(n_61156), .Z(n_161285889
		));
	notech_xor2 i_16764287(.A(pipe_mul[1]), .B(pipe_mul[0]), .Z(n_161385890)
		);
	notech_nand2 i_21264243(.A(divr_1[0]), .B(n_60184), .Z(n_161485891));
	notech_nand2 i_21864240(.A(divr_1[1]), .B(n_60184), .Z(n_161585892));
	notech_nand2 i_22164237(.A(divr_1[2]), .B(n_60171), .Z(n_161685893));
	notech_nand2 i_22464234(.A(divr_1[3]), .B(n_60171), .Z(n_161785894));
	notech_nand2 i_22764231(.A(divr_1[4]), .B(n_60171), .Z(n_161885895));
	notech_nand2 i_23064228(.A(divr_1[5]), .B(n_60184), .Z(n_161985896));
	notech_nand2 i_23364225(.A(divr_1[6]), .B(n_60171), .Z(n_162085897));
	notech_nand2 i_23664222(.A(divr_1[7]), .B(n_60195), .Z(n_162185898));
	notech_nand2 i_23964219(.A(divr_1[8]), .B(n_60195), .Z(n_162285899));
	notech_nand2 i_24364216(.A(divr_1[9]), .B(n_60195), .Z(n_162385900));
	notech_nand2 i_24664213(.A(divr_1[10]), .B(n_60195), .Z(n_162485901));
	notech_nand2 i_24964210(.A(divr_1[11]), .B(n_60195), .Z(n_162585902));
	notech_nand2 i_25364207(.A(divr_1[12]), .B(n_60193), .Z(n_162685903));
	notech_nand2 i_25664204(.A(divr_1[13]), .B(n_60193), .Z(n_162785904));
	notech_nand2 i_25964201(.A(divr_1[14]), .B(n_60193), .Z(n_162885905));
	notech_nand2 i_26264198(.A(divr_1[15]), .B(n_60195), .Z(n_162985906));
	notech_nand2 i_26664195(.A(divr_1[16]), .B(n_60193), .Z(n_163085907));
	notech_nand2 i_26964192(.A(divr_1[17]), .B(n_60195), .Z(n_163185908));
	notech_nand2 i_27264189(.A(divr_1[18]), .B(n_60195), .Z(n_163285909));
	notech_nand2 i_27864183(.A(divr_1[20]), .B(n_60195), .Z(n_163385910));
	notech_nand2 i_28164180(.A(divr_1[21]), .B(n_60195), .Z(n_163485911));
	notech_nand2 i_28464177(.A(divr_1[22]), .B(n_60171), .Z(n_163585912));
	notech_nand2 i_28864174(.A(divr_1[23]), .B(n_60195), .Z(n_163685913));
	notech_nand2 i_29164171(.A(divr_1[24]), .B(n_60195), .Z(n_163785914));
	notech_nand2 i_29464168(.A(divr_1[25]), .B(n_60195), .Z(n_163885915));
	notech_nand2 i_29764165(.A(divr_1[26]), .B(n_60195), .Z(n_163985916));
	notech_nand2 i_30064162(.A(divr_1[27]), .B(n_60195), .Z(n_164085917));
	notech_nand2 i_30364159(.A(divr_1[28]), .B(n_60195), .Z(n_164185918));
	notech_nand2 i_30664156(.A(divr_1[29]), .B(n_60173), .Z(n_164285919));
	notech_nand2 i_30964153(.A(divr_1[30]), .B(n_60173), .Z(n_164385920));
	notech_nand2 i_31264150(.A(divr_1[31]), .B(n_60173), .Z(n_164485921));
	notech_nand2 i_31564147(.A(divr_1[32]), .B(n_60173), .Z(n_164585922));
	notech_nand2 i_31864144(.A(divr_1[33]), .B(n_60173), .Z(n_164685923));
	notech_nand2 i_32164141(.A(divr_1[34]), .B(n_60178), .Z(n_164785924));
	notech_nand2 i_32464138(.A(divr_1[35]), .B(n_60178), .Z(n_164885925));
	notech_nand2 i_32764135(.A(divr_1[36]), .B(n_60178), .Z(n_164985926));
	notech_nand2 i_33064132(.A(divr_1[37]), .B(n_60178), .Z(n_165085927));
	notech_nand2 i_33364129(.A(divr_1[38]), .B(n_60178), .Z(n_165185928));
	notech_nand2 i_33664126(.A(divr_1[39]), .B(n_60173), .Z(n_165285929));
	notech_nand2 i_33964123(.A(divr_1[40]), .B(n_60173), .Z(n_165385930));
	notech_nand2 i_34264120(.A(divr_1[41]), .B(n_60173), .Z(n_165485931));
	notech_nand2 i_34564117(.A(divr_1[42]), .B(n_60173), .Z(n_165585932));
	notech_nand2 i_34864114(.A(divr_1[43]), .B(n_60173), .Z(n_165685933));
	notech_nand2 i_35164111(.A(divr_1[44]), .B(n_60173), .Z(n_165785934));
	notech_nand2 i_35564108(.A(divr_1[45]), .B(n_60173), .Z(n_165885935));
	notech_nand2 i_35864105(.A(divr_1[46]), .B(n_60173), .Z(n_165985936));
	notech_nand2 i_36264102(.A(divr_1[47]), .B(n_60173), .Z(n_166085937));
	notech_nand2 i_36564099(.A(divr_1[48]), .B(n_60173), .Z(n_166185938));
	notech_nand2 i_36864096(.A(divr_1[49]), .B(n_60173), .Z(n_166285939));
	notech_nand2 i_37164093(.A(divr_1[50]), .B(n_60184), .Z(n_166385940));
	notech_nand2 i_37464090(.A(divr_1[51]), .B(n_60184), .Z(n_166485941));
	notech_nand2 i_37764087(.A(divr_1[52]), .B(n_60184), .Z(n_166585942));
	notech_nand2 i_38064084(.A(divr_1[53]), .B(n_60184), .Z(n_166685943));
	notech_nand2 i_38364081(.A(divr_1[54]), .B(n_60184), .Z(n_166785944));
	notech_nand2 i_38664078(.A(divr_1[55]), .B(n_60184), .Z(n_166885945));
	notech_nand2 i_38964075(.A(divr_1[56]), .B(n_60184), .Z(n_166985946));
	notech_nand2 i_39264072(.A(divr_1[57]), .B(n_60184), .Z(n_167085947));
	notech_nand2 i_39564069(.A(divr_1[58]), .B(n_60184), .Z(n_167185948));
	notech_nand2 i_39864066(.A(divr_1[59]), .B(n_60184), .Z(n_167285949));
	notech_nand2 i_40164063(.A(divr_1[60]), .B(n_60178), .Z(n_167385950));
	notech_nand2 i_40464060(.A(divr_1[61]), .B(n_60178), .Z(n_167485951));
	notech_nand2 i_40764057(.A(divr_1[62]), .B(n_60178), .Z(n_167585952));
	notech_nand2 i_41164053(.A(divr_1[63]), .B(n_60178), .Z(n_167685953));
	notech_or2 i_41464050(.A(n_55524), .B(n_29475), .Z(n_167785954));
	notech_ao4 i_26564456(.A(n_313784128), .B(n_60178), .C(n_148282483), .D(opb
		[31]), .Z(n_167885955));
	notech_or2 i_55263918(.A(n_55525), .B(n_29507), .Z(n_168085957));
	notech_and2 i_17960(.A(n_161285889), .B(regs_10[17]), .Z(n_168285959));
	notech_ao3 i_23300(.A(n_1891), .B(n_60298), .C(pipe_mul[0]), .Z(n_194086214
		));
	notech_and3 i_23301(.A(n_161385890), .B(n_1891), .C(n_60298), .Z(n_194186215
		));
	notech_ao4 i_130063190(.A(n_55508), .B(n_29505), .C(n_148382484), .D(n_30372
		), .Z(n_194286216));
	notech_ao4 i_129963191(.A(n_148382484), .B(n_30371), .C(n_247640494), .D
		(n_57837), .Z(n_194386217));
	notech_ao4 i_129863192(.A(n_55524), .B(n_29506), .C(n_55508), .D(n_29504
		), .Z(n_194486218));
	notech_ao4 i_129763193(.A(n_148382484), .B(n_30369), .C(n_167885955), .D
		(n_55929), .Z(n_194586219));
	notech_ao4 i_129663194(.A(n_55508), .B(n_29503), .C(n_55524), .D(n_29505
		), .Z(n_194686220));
	notech_ao4 i_129563195(.A(n_148382484), .B(n_30368), .C(n_167885955), .D
		(n_55956), .Z(n_194786221));
	notech_ao4 i_129463196(.A(n_55524), .B(n_29504), .C(n_55508), .D(n_29502
		), .Z(n_194886222));
	notech_ao4 i_129363197(.A(n_148382484), .B(n_30367), .C(n_167885955), .D
		(\nbus_11358[28] ), .Z(n_194986223));
	notech_ao4 i_129263198(.A(n_55524), .B(n_29503), .C(n_55508), .D(n_29501
		), .Z(n_195086224));
	notech_ao4 i_129163199(.A(n_148382484), .B(n_30364), .C(n_167885955), .D
		(\nbus_11358[27] ), .Z(n_195186225));
	notech_ao4 i_129063200(.A(n_55524), .B(n_29502), .C(n_55508), .D(n_29500
		), .Z(n_195286226));
	notech_ao4 i_128963201(.A(n_148382484), .B(n_30363), .C(n_167885955), .D
		(n_55947), .Z(n_195386227));
	notech_ao4 i_128863202(.A(n_55524), .B(n_29501), .C(n_55508), .D(n_29499
		), .Z(n_195486228));
	notech_ao4 i_128763203(.A(n_148382484), .B(n_30362), .C(n_167885955), .D
		(n_55965), .Z(n_195586229));
	notech_ao4 i_128663204(.A(n_55524), .B(n_29500), .C(n_55508), .D(n_29498
		), .Z(n_195686230));
	notech_ao4 i_128563205(.A(n_148382484), .B(n_30360), .C(n_167885955), .D
		(n_56475), .Z(n_195786231));
	notech_ao4 i_128463206(.A(n_55524), .B(n_29499), .C(n_55509), .D(n_29497
		), .Z(n_195886232));
	notech_ao4 i_128263207(.A(n_148382484), .B(n_30358), .C(n_167885955), .D
		(n_56347), .Z(n_195986233));
	notech_ao4 i_128163208(.A(n_55524), .B(n_29498), .C(n_55509), .D(n_29496
		), .Z(n_196086234));
	notech_ao4 i_128063209(.A(n_148382484), .B(n_30356), .C(n_167885955), .D
		(n_56338), .Z(n_196186235));
	notech_ao4 i_127963210(.A(n_55524), .B(n_29497), .C(n_55509), .D(n_29495
		), .Z(n_196286236));
	notech_ao4 i_127863211(.A(n_148382484), .B(n_30355), .C(n_167885955), .D
		(n_56329), .Z(n_196386237));
	notech_ao4 i_127763212(.A(n_55525), .B(n_29496), .C(n_55509), .D(n_29494
		), .Z(n_196486238));
	notech_ao4 i_127663213(.A(n_148382484), .B(n_30354), .C(n_167885955), .D
		(n_56320), .Z(n_196586239));
	notech_ao4 i_127563214(.A(n_55525), .B(n_29495), .C(n_55509), .D(n_29493
		), .Z(n_196686240));
	notech_ao4 i_127463215(.A(n_148382484), .B(n_30353), .C(n_167885955), .D
		(n_56311), .Z(n_196786241));
	notech_ao4 i_127363216(.A(n_55525), .B(n_29494), .C(n_55509), .D(n_29492
		), .Z(n_196886242));
	notech_ao4 i_127263217(.A(n_148382484), .B(n_30351), .C(n_167885955), .D
		(n_56302), .Z(n_196986243));
	notech_ao4 i_127163218(.A(n_55525), .B(n_29493), .C(n_55509), .D(n_29491
		), .Z(n_197086244));
	notech_ao4 i_127063219(.A(n_148382484), .B(n_30349), .C(n_167885955), .D
		(n_56293), .Z(n_197186245));
	notech_ao4 i_126963220(.A(n_55525), .B(n_29492), .C(n_55509), .D(n_29490
		), .Z(n_197286246));
	notech_ao4 i_126863221(.A(n_55489), .B(n_30348), .C(n_167885955), .D(n_56284
		), .Z(n_197386247));
	notech_ao4 i_126763222(.A(n_55525), .B(n_29491), .C(n_55509), .D(n_29489
		), .Z(n_197486248));
	notech_ao4 i_126663223(.A(n_55489), .B(n_30347), .C(n_167885955), .D(n_56275
		), .Z(n_197586249));
	notech_ao4 i_126563224(.A(n_55525), .B(n_29490), .C(n_55509), .D(n_29488
		), .Z(n_197686250));
	notech_ao4 i_126463225(.A(n_55489), .B(n_30346), .C(n_55480), .D(\nbus_11358[14] 
		), .Z(n_197786251));
	notech_ao4 i_126363226(.A(n_55525), .B(n_29489), .C(n_55509), .D(n_29487
		), .Z(n_197886252));
	notech_ao4 i_126263227(.A(n_55489), .B(n_30345), .C(n_55480), .D(n_56230
		), .Z(n_197986253));
	notech_ao4 i_126163228(.A(n_55525), .B(n_29488), .C(n_55509), .D(n_29486
		), .Z(n_198086254));
	notech_ao4 i_126063229(.A(n_55489), .B(n_30343), .C(n_55480), .D(n_56221
		), .Z(n_198186255));
	notech_ao4 i_125963230(.A(n_55525), .B(n_29487), .C(n_55509), .D(n_29485
		), .Z(n_198286256));
	notech_ao4 i_125863231(.A(n_55489), .B(n_30341), .C(n_55480), .D(n_56181
		), .Z(n_198386257));
	notech_ao4 i_125763232(.A(n_55525), .B(n_29486), .C(n_55509), .D(n_29484
		), .Z(n_198486258));
	notech_ao4 i_125663233(.A(n_55489), .B(n_30340), .C(n_55480), .D(n_56154
		), .Z(n_198586259));
	notech_ao4 i_125563234(.A(n_55525), .B(n_29485), .C(n_55509), .D(n_29483
		), .Z(n_198686260));
	notech_ao4 i_125463235(.A(n_55489), .B(n_30339), .C(n_55480), .D(n_56136
		), .Z(n_198786261));
	notech_ao4 i_125363236(.A(n_55525), .B(n_29484), .C(n_55509), .D(n_29482
		), .Z(n_198886262));
	notech_ao4 i_125263237(.A(n_55489), .B(n_30338), .C(n_55480), .D(n_56118
		), .Z(n_198986263));
	notech_ao4 i_125163238(.A(n_55525), .B(n_29483), .C(n_55509), .D(n_29481
		), .Z(n_199086264));
	notech_ao4 i_125063239(.A(n_55489), .B(n_30337), .C(n_55480), .D(n_56109
		), .Z(n_199186265));
	notech_ao4 i_124963240(.A(n_55525), .B(n_29482), .C(n_55509), .D(n_29480
		), .Z(n_199286266));
	notech_ao4 i_124863241(.A(n_55489), .B(n_30336), .C(n_55480), .D(n_56082
		), .Z(n_199386267));
	notech_ao4 i_124763242(.A(n_55525), .B(n_29481), .C(n_55498), .D(n_29479
		), .Z(n_199486268));
	notech_ao4 i_124663243(.A(n_148382484), .B(n_30335), .C(n_55480), .D(\nbus_11358[5] 
		), .Z(n_199586269));
	notech_ao4 i_124563244(.A(n_55525), .B(n_29480), .C(n_55498), .D(n_29478
		), .Z(n_199686270));
	notech_ao4 i_124463245(.A(n_55489), .B(n_30334), .C(n_55480), .D(n_56064
		), .Z(n_199786271));
	notech_ao4 i_124363246(.A(n_55524), .B(n_29479), .C(n_55498), .D(n_29477
		), .Z(n_199886272));
	notech_ao4 i_124263247(.A(n_55489), .B(n_30333), .C(n_55480), .D(n_55983
		), .Z(n_199986273));
	notech_ao4 i_124163248(.A(n_55514), .B(n_29478), .C(n_55498), .D(n_29476
		), .Z(n_200086274));
	notech_ao4 i_124063249(.A(n_55489), .B(n_30331), .C(n_55480), .D(n_55992
		), .Z(n_200186275));
	notech_ao4 i_123963250(.A(n_55514), .B(n_29477), .C(n_55498), .D(n_29475
		), .Z(n_200286276));
	notech_ao4 i_123863251(.A(n_55489), .B(n_30330), .C(n_55480), .D(\nbus_11358[1] 
		), .Z(n_200386277));
	notech_ao4 i_123763252(.A(n_29476), .B(n_55514), .C(n_55498), .D(n_29474
		), .Z(n_200486278));
	notech_ao4 i_122963259(.A(n_55489), .B(n_30327), .C(n_55480), .D(n_56028
		), .Z(n_200586279));
	notech_ao4 i_122863260(.A(n_55564), .B(n_30326), .C(n_247640494), .D(nbus_11295
		[31]), .Z(n_200686280));
	notech_ao4 i_122763261(.A(n_55564), .B(n_30324), .C(n_55549), .D(nbus_11295
		[30]), .Z(n_200786281));
	notech_ao4 i_122663262(.A(n_55565), .B(n_30323), .C(n_55549), .D(nbus_11295
		[29]), .Z(n_200886282));
	notech_ao4 i_122563263(.A(n_55565), .B(n_30321), .C(n_55549), .D(nbus_11295
		[28]), .Z(n_200986283));
	notech_ao4 i_122463264(.A(n_55564), .B(n_30320), .C(n_55549), .D(n_57881
		), .Z(n_201086284));
	notech_ao4 i_122363265(.A(n_55564), .B(n_30319), .C(n_55549), .D(nbus_11295
		[26]), .Z(n_201186285));
	notech_ao4 i_122163266(.A(n_55564), .B(n_30318), .C(n_55549), .D(nbus_11295
		[25]), .Z(n_201286286));
	notech_ao4 i_122063267(.A(n_55564), .B(n_30317), .C(n_55549), .D(nbus_11295
		[24]), .Z(n_201386287));
	notech_ao4 i_121963268(.A(n_55564), .B(n_30316), .C(n_55545), .D(nbus_11295
		[23]), .Z(n_201486288));
	notech_ao4 i_121863269(.A(n_55564), .B(n_30314), .C(n_55545), .D(nbus_11295
		[22]), .Z(n_201586289));
	notech_ao4 i_121763270(.A(n_55564), .B(n_30313), .C(n_55545), .D(nbus_11295
		[21]), .Z(n_201686290));
	notech_ao4 i_121663271(.A(n_55564), .B(n_30309), .C(n_55549), .D(nbus_11295
		[20]), .Z(n_201786291));
	notech_ao4 i_121563272(.A(n_55564), .B(n_30308), .C(n_55549), .D(nbus_11295
		[19]), .Z(n_201886292));
	notech_ao4 i_121463273(.A(n_55564), .B(n_30307), .C(n_55549), .D(nbus_11295
		[18]), .Z(n_201986293));
	notech_ao4 i_121363274(.A(n_55565), .B(n_30304), .C(n_55549), .D(nbus_11295
		[17]), .Z(n_202086294));
	notech_ao4 i_121263275(.A(n_55565), .B(n_30302), .C(n_55549), .D(nbus_11295
		[16]), .Z(n_202186295));
	notech_ao4 i_121163276(.A(n_55565), .B(n_30298), .C(n_55550), .D(nbus_11295
		[15]), .Z(n_202286296));
	notech_ao4 i_120963277(.A(n_55565), .B(n_30297), .C(n_55550), .D(nbus_11295
		[14]), .Z(n_202386297));
	notech_ao4 i_120863278(.A(n_55565), .B(n_30296), .C(n_55550), .D(nbus_11295
		[13]), .Z(n_202486298));
	notech_ao4 i_120763279(.A(n_55565), .B(n_30295), .C(n_55550), .D(nbus_11295
		[12]), .Z(n_202586299));
	notech_ao4 i_120663280(.A(n_55565), .B(n_30293), .C(n_55550), .D(nbus_11295
		[11]), .Z(n_202686300));
	notech_ao4 i_120563281(.A(n_55565), .B(n_30292), .C(n_55550), .D(nbus_11295
		[10]), .Z(n_202786301));
	notech_ao4 i_120463282(.A(n_55565), .B(n_30291), .C(n_55550), .D(nbus_11295
		[9]), .Z(n_202886302));
	notech_ao4 i_120363283(.A(n_55565), .B(n_30289), .C(n_55550), .D(nbus_11295
		[8]), .Z(n_202986303));
	notech_ao4 i_120263284(.A(n_55565), .B(n_30288), .C(n_55550), .D(nbus_11295
		[7]), .Z(n_203086304));
	notech_ao4 i_120163285(.A(n_55565), .B(n_30287), .C(n_55550), .D(nbus_11295
		[6]), .Z(n_203186305));
	notech_ao4 i_120063286(.A(n_55565), .B(n_30286), .C(n_55549), .D(nbus_11295
		[5]), .Z(n_203286306));
	notech_ao4 i_119963287(.A(n_55565), .B(n_30285), .C(n_55550), .D(nbus_11295
		[4]), .Z(n_203386307));
	notech_ao4 i_119863288(.A(n_55565), .B(n_30284), .C(n_55550), .D(n_57909
		), .Z(n_203486308));
	notech_ao4 i_119763289(.A(n_55565), .B(n_30283), .C(n_55550), .D(nbus_11295
		[2]), .Z(n_203586309));
	notech_ao4 i_119663290(.A(n_55564), .B(n_30282), .C(n_55550), .D(nbus_11295
		[1]), .Z(n_203686310));
	notech_ao4 i_119563291(.A(n_55559), .B(n_30281), .C(n_55545), .D(n_59717
		), .Z(n_203786311));
	notech_ao4 i_119463292(.A(n_55559), .B(n_30280), .C(n_55542), .D(n_59726
		), .Z(n_203886312));
	notech_ao4 i_119363293(.A(n_55554), .B(n_30279), .C(n_55542), .D(n_57828
		), .Z(n_203986313));
	notech_ao4 i_119263294(.A(n_55554), .B(n_30277), .C(n_55542), .D(n_57815
		), .Z(n_204086314));
	notech_ao4 i_119163295(.A(n_55559), .B(n_30276), .C(n_55542), .D(n_57802
		), .Z(n_204186315));
	notech_ao4 i_119063296(.A(n_55559), .B(n_30275), .C(n_55542), .D(n_57792
		), .Z(n_204286316));
	notech_ao4 i_118963297(.A(n_55559), .B(n_30271), .C(n_55542), .D(n_57783
		), .Z(n_204386317));
	notech_ao4 i_118863298(.A(n_55559), .B(n_30267), .C(n_55542), .D(n_57771
		), .Z(n_204486318));
	notech_ao4 i_118763299(.A(n_55554), .B(n_30265), .C(n_55542), .D(n_57761
		), .Z(n_204586319));
	notech_ao4 i_118663300(.A(n_55554), .B(n_30263), .C(n_55541), .D(n_57751
		), .Z(n_204686320));
	notech_ao4 i_118563301(.A(n_55554), .B(n_30262), .C(n_55541), .D(n_57742
		), .Z(n_204786321));
	notech_ao4 i_118463302(.A(n_55554), .B(n_30260), .C(n_55541), .D(n_57733
		), .Z(n_204886322));
	notech_ao4 i_118363303(.A(n_55554), .B(n_30259), .C(n_55541), .D(n_57720
		), .Z(n_204986323));
	notech_ao4 i_118163305(.A(n_55554), .B(n_30257), .C(n_55541), .D(n_57698
		), .Z(n_205086324));
	notech_ao4 i_118063306(.A(n_55554), .B(n_30255), .C(n_55541), .D(n_57689
		), .Z(n_205186325));
	notech_ao4 i_117963307(.A(n_55554), .B(n_30253), .C(n_55541), .D(n_57680
		), .Z(n_205286326));
	notech_ao4 i_117863308(.A(n_55559), .B(n_30252), .C(n_55542), .D(n_57671
		), .Z(n_205386327));
	notech_ao4 i_117763309(.A(n_55559), .B(n_30250), .C(n_55545), .D(n_57662
		), .Z(n_205486328));
	notech_ao4 i_117663310(.A(n_55559), .B(n_30249), .C(n_55545), .D(n_57653
		), .Z(n_205586329));
	notech_ao4 i_117563311(.A(n_55559), .B(n_30248), .C(n_55545), .D(n_57644
		), .Z(n_205686330));
	notech_ao4 i_117463312(.A(n_55564), .B(n_30247), .C(n_55545), .D(n_57635
		), .Z(n_205786331));
	notech_ao4 i_117363313(.A(n_55564), .B(n_30245), .C(n_55545), .D(n_57625
		), .Z(n_205886332));
	notech_ao4 i_117163314(.A(n_55559), .B(n_30243), .C(n_55545), .D(n_57613
		), .Z(n_205986333));
	notech_ao4 i_117063315(.A(n_55559), .B(n_30242), .C(n_55545), .D(n_57604
		), .Z(n_206086334));
	notech_ao4 i_116963316(.A(n_55559), .B(n_30241), .C(n_55545), .D(\nbus_11307[7] 
		), .Z(n_206186335));
	notech_ao4 i_116763317(.A(n_55559), .B(n_30240), .C(n_55542), .D(n_57592
		), .Z(n_206286336));
	notech_ao4 i_116663318(.A(n_55559), .B(n_30239), .C(n_55542), .D(n_57583
		), .Z(n_206386337));
	notech_ao4 i_116563319(.A(n_55559), .B(n_30238), .C(n_55542), .D(n_57574
		), .Z(n_206486338));
	notech_ao4 i_116463320(.A(n_55559), .B(n_30237), .C(n_55542), .D(n_57563
		), .Z(n_206586339));
	notech_ao4 i_116363321(.A(n_55559), .B(n_30236), .C(n_55545), .D(n_57552
		), .Z(n_206686340));
	notech_ao4 i_116263322(.A(n_55559), .B(n_30235), .C(n_55545), .D(n_57542
		), .Z(n_206786341));
	notech_ao4 i_116163323(.A(n_55559), .B(n_30234), .C(n_55542), .D(n_59742
		), .Z(n_206886342));
	notech_nand2 i_123855513(.A(n_58786), .B(n_207086344), .Z(n_206986343)
		);
	notech_or4 i_17255348(.A(n_60868), .B(n_2884), .C(n_27063), .D(n_27047),
		 .Z(n_207086344));
	notech_nao3 i_15955361(.A(n_11255), .B(n_60298), .C(n_304384034), .Z(n_207486348
		));
	notech_nao3 i_15655364(.A(n_11256), .B(n_60298), .C(n_1893), .Z(n_207786351
		));
	notech_or2 i_15355367(.A(n_55367), .B(n_28387), .Z(n_208086354));
	notech_nand3 i_14855372(.A(n_206986343), .B(opd[0]), .C(n_60298), .Z(n_208186355
		));
	notech_or4 i_14955371(.A(n_28533), .B(n_59424), .C(n_60178), .D(n_56028)
		, .Z(n_208286356));
	notech_or4 i_15055370(.A(n_59478), .B(n_27573), .C(n_57132), .D(n_59717)
		, .Z(n_208386357));
	notech_nao3 i_17155349(.A(n_11257), .B(n_60298), .C(n_304384034), .Z(n_208686360
		));
	notech_nao3 i_16855352(.A(Daddrgs[1]), .B(n_27063), .C(n_326591251), .Z(n_208986363
		));
	notech_nao3 i_16555355(.A(Daddrs_8[1]), .B(n_60298), .C(n_319591628), .Z
		(n_209286366));
	notech_nand3 i_16055360(.A(opd[1]), .B(n_60312), .C(n_206986343), .Z(n_209386367
		));
	notech_or4 i_16155359(.A(n_28533), .B(n_59424), .C(n_60178), .D(n_56010)
		, .Z(n_209486368));
	notech_nand2 i_16255358(.A(Daddrs_1[1]), .B(n_27066), .Z(n_209586369));
	notech_or4 i_112555514(.A(instrc[110]), .B(instrc[111]), .C(n_29175), .D
		(n_29176), .Z(n_209886372));
	notech_ao4 i_100055528(.A(n_59451), .B(n_330763524), .C(n_38609), .D(n_209886372
		), .Z(n_209986373));
	notech_and3 i_53855006(.A(n_209486368), .B(n_209386367), .C(n_209586369)
		, .Z(n_210386377));
	notech_ao4 i_53355009(.A(n_55367), .B(n_28388), .C(n_55389), .D(n_28594)
		, .Z(n_210486378));
	notech_ao4 i_52855012(.A(n_59167), .B(n_30376), .C(n_59335), .D(n_29317)
		, .Z(n_210786381));
	notech_ao4 i_52455014(.A(n_55347), .B(nbus_11295[1]), .C(n_55409), .D(n_30375
		), .Z(n_210986383));
	notech_and4 i_53055010(.A(n_210986383), .B(n_210786381), .C(n_208686360)
		, .D(n_208986363), .Z(n_211186385));
	notech_and3 i_52055017(.A(n_208286356), .B(n_208186355), .C(n_208386357)
		, .Z(n_211486388));
	notech_ao4 i_51455020(.A(n_55389), .B(n_28593), .C(n_55378), .D(n_29347)
		, .Z(n_211586389));
	notech_ao4 i_50955023(.A(n_59335), .B(n_29316), .C(n_59147), .D(n_29285)
		, .Z(n_211886392));
	notech_ao4 i_50755025(.A(n_55409), .B(n_30373), .C(n_59176), .D(n_27804)
		, .Z(n_212086394));
	notech_and4 i_51355021(.A(n_212086394), .B(n_211886392), .C(n_207486348)
		, .D(n_207786351), .Z(n_212286396));
	notech_ao4 i_53863(.A(n_57818), .B(n_116568182), .C(n_3986), .D(n_61109)
		, .Z(n_21651));
	notech_xor2 i_5750609(.A(vliw_pc[1]), .B(vliw_pc[0]), .Z(n_212486398));
	notech_xor2 i_5850608(.A(n_32843), .B(vliw_pc[2]), .Z(n_212586399));
	notech_xor2 i_5950607(.A(vliw_pc[3]), .B(n_32834), .Z(n_212686400));
	notech_xor2 i_6050606(.A(vliw_pc[4]), .B(n_214786421), .Z(n_212786401)
		);
	notech_ao4 i_24350672(.A(n_59095), .B(n_18964), .C(n_61109), .D(n_27048)
		, .Z(n_212886402));
	notech_or4 i_5650610(.A(n_27501), .B(n_60894), .C(n_59478), .D(n_27980),
		 .Z(n_213886412));
	notech_and2 i_18280(.A(n_212486398), .B(n_27049), .Z(n_214286416));
	notech_and2 i_18281(.A(n_27049), .B(n_212586399), .Z(n_214386417));
	notech_and2 i_18282(.A(n_27049), .B(n_212686400), .Z(n_214486418));
	notech_and2 i_18283(.A(n_212786401), .B(n_27049), .Z(n_214586419));
	notech_and4 i_6150605(.A(vliw_pc[3]), .B(vliw_pc[0]), .C(vliw_pc[1]), .D
		(vliw_pc[2]), .Z(n_214786421));
	notech_ao4 i_106349630(.A(n_5380), .B(n_59095), .C(vliw_pc[0]), .D(n_212886402
		), .Z(n_214886422));
	notech_mux2 i_3641221(.S(n_57899), .A(n_215186425), .B(n_59717), .Z(n_214986423
		));
	notech_and2 i_3741220(.A(n_276487038), .B(n_215486428), .Z(n_215186425)
		);
	notech_and3 i_3841219(.A(n_57406), .B(n_58675), .C(n_58697), .Z(n_215386427
		));
	notech_nand2 i_7741180(.A(\opc_1[0] ), .B(rep_en1), .Z(n_215486428));
	notech_xor2 i_3341223(.A(opc[1]), .B(n_59735), .Z(n_215586429));
	notech_and3 i_3541222(.A(n_271686990), .B(n_55886), .C(n_220686480), .Z(n_215686430
		));
	notech_and3 i_3141225(.A(n_55886), .B(n_216286436), .C(n_215986433), .Z(n_215786431
		));
	notech_and2 i_3241224(.A(n_271686990), .B(n_273487008), .Z(n_215886432)
		);
	notech_nao3 i_10841149(.A(n_291218111), .B(n_27050), .C(n_271086984), .Z
		(n_215986433));
	notech_and3 i_2941227(.A(n_55886), .B(n_271786991), .C(n_216286436), .Z(n_216086434
		));
	notech_and2 i_3041226(.A(n_271686990), .B(n_271486988), .Z(n_216186435)
		);
	notech_nao3 i_13041128(.A(n_291418113), .B(n_269686970), .C(n_271086984)
		, .Z(n_216286436));
	notech_mux2 i_2341233(.S(n_57899), .A(n_216786441), .B(n_216586439), .Z(n_216386437
		));
	notech_xor2 i_2441232(.A(opc[4]), .B(n_27959), .Z(n_216586439));
	notech_and2 i_2541231(.A(n_269886972), .B(n_269786971), .Z(n_216786441)
		);
	notech_xor2 i_2641230(.A(opc[4]), .B(n_269586969), .Z(n_216986443));
	notech_xor2 i_2741229(.A(n_291118110), .B(opc[4]), .Z(n_217086444));
	notech_ao4 i_23641287(.A(n_32656), .B(n_60178), .C(n_32559), .D(n_248786761
		), .Z(n_217486448));
	notech_or4 i_40640865(.A(n_59413), .B(n_25629), .C(n_60178), .D(n_57957)
		, .Z(n_217586449));
	notech_or4 i_7041187(.A(n_60894), .B(n_60178), .C(n_26965), .D(nbus_11295
		[24]), .Z(n_218186455));
	notech_nao3 i_6741190(.A(mul64[32]), .B(n_60319), .C(n_314563412), .Z(n_218486458
		));
	notech_or2 i_9241165(.A(n_58651), .B(n_28125), .Z(n_219186465));
	notech_nao3 i_9341164(.A(n_27050), .B(n_59717), .C(n_271086984), .Z(n_220686480
		));
	notech_or2 i_12741131(.A(n_58651), .B(n_28127), .Z(n_222386497));
	notech_ao3 i_11341144(.A(\opc_1[3] ), .B(rep_en1), .C(n_271086984), .Z(n_223886512
		));
	notech_or4 i_14041118(.A(n_60894), .B(n_60178), .C(n_26965), .D(nbus_11295
		[28]), .Z(n_224586519));
	notech_or2 i_13741121(.A(n_55886), .B(nbus_11295[4]), .Z(n_224886522));
	notech_nao3 i_17641084(.A(n_60319), .B(mul64[25]), .C(n_2647), .Z(n_226186535
		));
	notech_or4 i_17341087(.A(n_60894), .B(n_60193), .C(n_26965), .D(nbus_11295
		[17]), .Z(n_226486538));
	notech_nao3 i_18841072(.A(n_60321), .B(mul64[26]), .C(n_2647), .Z(n_227386547
		));
	notech_or4 i_18541075(.A(n_60894), .B(n_60218), .C(n_26965), .D(nbus_11295
		[18]), .Z(n_227686550));
	notech_nao3 i_20041060(.A(n_60321), .B(mul64[27]), .C(n_2647), .Z(n_228586559
		));
	notech_or4 i_19741063(.A(n_60894), .B(n_60218), .C(n_26965), .D(nbus_11295
		[19]), .Z(n_228886562));
	notech_nao3 i_21241048(.A(n_60319), .B(mul64[28]), .C(n_2647), .Z(n_229786571
		));
	notech_or4 i_20941051(.A(n_60894), .B(n_60218), .C(n_26965), .D(nbus_11295
		[20]), .Z(n_230086574));
	notech_nao3 i_22441036(.A(n_60319), .B(mul64[29]), .C(n_2647), .Z(n_230986583
		));
	notech_or4 i_22141039(.A(n_60894), .B(n_60218), .C(n_26965), .D(nbus_11295
		[21]), .Z(n_231286586));
	notech_nao3 i_23741024(.A(n_60319), .B(mul64[30]), .C(n_2647), .Z(n_232186595
		));
	notech_or4 i_23341027(.A(n_60894), .B(n_60218), .C(n_26965), .D(nbus_11295
		[22]), .Z(n_232486598));
	notech_or4 i_24941012(.A(n_60894), .B(n_60218), .C(n_26965), .D(nbus_11295
		[23]), .Z(n_233386607));
	notech_or2 i_24641015(.A(n_55886), .B(n_56109), .Z(n_233686610));
	notech_or2 i_26041001(.A(n_57367), .B(n_56284), .Z(n_234186615));
	notech_nao3 i_25941002(.A(n_60373), .B(divr[16]), .C(n_57537), .Z(n_234486618
		));
	notech_or4 i_25441007(.A(n_60894), .B(n_60218), .C(n_26965), .D(nbus_11295
		[8]), .Z(n_234986623));
	notech_or2 i_27140992(.A(n_57367), .B(n_56293), .Z(n_235086624));
	notech_nao3 i_27040993(.A(n_60373), .B(divr[17]), .C(n_57537), .Z(n_235386627
		));
	notech_or4 i_26440998(.A(n_60893), .B(n_60218), .C(n_26965), .D(nbus_11295
		[9]), .Z(n_235886632));
	notech_or2 i_28040983(.A(n_57367), .B(n_56302), .Z(n_235986633));
	notech_nao3 i_27940984(.A(n_60373), .B(divr[18]), .C(n_57537), .Z(n_236286636
		));
	notech_or4 i_27440989(.A(n_60883), .B(n_60218), .C(n_26965), .D(nbus_11295
		[10]), .Z(n_236786641));
	notech_or2 i_29040974(.A(n_57367), .B(n_56311), .Z(n_236886642));
	notech_nao3 i_28940975(.A(n_60373), .B(divr[19]), .C(n_57537), .Z(n_237186645
		));
	notech_or4 i_28440980(.A(n_60883), .B(n_60218), .C(n_58033), .D(nbus_11295
		[11]), .Z(n_237686650));
	notech_or2 i_29940965(.A(n_57367), .B(n_56320), .Z(n_237786651));
	notech_nao3 i_29840966(.A(n_60373), .B(divr[20]), .C(n_57537), .Z(n_238086654
		));
	notech_or4 i_29340971(.A(n_60883), .B(n_60212), .C(n_58033), .D(nbus_11295
		[12]), .Z(n_238586659));
	notech_or2 i_30840956(.A(n_57367), .B(n_56329), .Z(n_238686660));
	notech_nao3 i_30740957(.A(n_60373), .B(divr[21]), .C(n_57533), .Z(n_238986663
		));
	notech_or4 i_30240962(.A(n_60212), .B(n_60883), .C(n_58033), .D(nbus_11295
		[13]), .Z(n_239486668));
	notech_or2 i_31740947(.A(n_57367), .B(n_56338), .Z(n_239586669));
	notech_nao3 i_31640948(.A(n_60373), .B(divr[22]), .C(n_57533), .Z(n_239886672
		));
	notech_or4 i_31140953(.A(n_60883), .B(n_60212), .C(n_58033), .D(nbus_11295
		[14]), .Z(n_240386677));
	notech_or2 i_32840938(.A(n_57367), .B(n_56347), .Z(n_240486678));
	notech_nao3 i_32740939(.A(n_60373), .B(divr[23]), .C(n_57533), .Z(n_240786681
		));
	notech_or4 i_32140944(.A(n_60888), .B(n_60212), .C(n_58033), .D(nbus_11295
		[15]), .Z(n_241286686));
	notech_or2 i_33740929(.A(n_57367), .B(n_56475), .Z(n_241386687));
	notech_nao3 i_33640930(.A(n_60373), .B(divr[24]), .C(n_57537), .Z(n_241686690
		));
	notech_or4 i_33140935(.A(n_60883), .B(n_60212), .C(n_58033), .D(nbus_11295
		[0]), .Z(n_242186695));
	notech_or4 i_34740920(.A(n_60883), .B(n_60212), .C(n_58033), .D(nbus_11295
		[1]), .Z(n_242286696));
	notech_or2 i_34640921(.A(n_57367), .B(n_55965), .Z(n_242586699));
	notech_nand2 i_34040926(.A(opc_14[25]), .B(n_19101), .Z(n_243086704));
	notech_or4 i_35640911(.A(n_60883), .B(n_60212), .C(n_58033), .D(nbus_11295
		[2]), .Z(n_243186705));
	notech_or2 i_35540912(.A(n_57367), .B(n_55947), .Z(n_243486708));
	notech_nand2 i_35040917(.A(opc_14[26]), .B(n_19101), .Z(n_243986713));
	notech_or4 i_36540902(.A(n_60883), .B(n_60212), .C(n_58033), .D(n_57909)
		, .Z(n_244086714));
	notech_or2 i_36440903(.A(n_57367), .B(n_55938), .Z(n_244386717));
	notech_nand2 i_35940908(.A(opc_14[27]), .B(n_19101), .Z(n_244886722));
	notech_or4 i_37540893(.A(n_60883), .B(n_60212), .C(n_58033), .D(nbus_11295
		[4]), .Z(n_244986723));
	notech_or2 i_37440894(.A(n_57367), .B(n_55974), .Z(n_245286726));
	notech_nand2 i_36840899(.A(opc_14[28]), .B(n_19101), .Z(n_245786731));
	notech_or4 i_38540884(.A(n_60883), .B(n_60212), .C(n_58033), .D(nbus_11295
		[5]), .Z(n_245886732));
	notech_or2 i_38340885(.A(n_57367), .B(n_55956), .Z(n_246186735));
	notech_nand2 i_37840890(.A(opc_14[29]), .B(n_19101), .Z(n_246686740));
	notech_or4 i_39640875(.A(n_60883), .B(n_60212), .C(n_26965), .D(nbus_11295
		[6]), .Z(n_246786741));
	notech_or2 i_39440876(.A(n_57367), .B(n_55929), .Z(n_247086744));
	notech_nand2 i_38840881(.A(opc_14[30]), .B(n_19101), .Z(n_247586749));
	notech_or4 i_40540866(.A(n_60883), .B(n_60223), .C(n_58033), .D(nbus_11295
		[7]), .Z(n_247686750));
	notech_or2 i_40440867(.A(n_55592), .B(\nbus_11358[31] ), .Z(n_247986753)
		);
	notech_nand2 i_39940872(.A(opc_14[31]), .B(n_19101), .Z(n_248486758));
	notech_or4 i_26141286(.A(n_32581), .B(n_19057), .C(n_60319), .D(n_18964)
		, .Z(n_248686760));
	notech_nand3 i_136539997(.A(n_19093), .B(n_60373), .C(n_18964), .Z(n_248786761
		));
	notech_ao4 i_136140001(.A(n_217486448), .B(n_28157), .C(n_248686760), .D
		(n_30438), .Z(n_248886762));
	notech_ao4 i_136040002(.A(n_55886), .B(nbus_11295[31]), .C(n_227976218),
		 .D(n_30172), .Z(n_249086764));
	notech_ao4 i_135740005(.A(n_308084071), .B(nbus_11328[31]), .C(n_307884069
		), .D(n_30437), .Z(n_249286766));
	notech_and3 i_28241285(.A(n_304584036), .B(n_217586449), .C(n_304284033)
		, .Z(n_249586769));
	notech_and4 i_135940003(.A(n_249586769), .B(n_249286766), .C(n_247686750
		), .D(n_247986753), .Z(n_249786771));
	notech_ao4 i_135240009(.A(n_217486448), .B(n_28156), .C(n_248686760), .D
		(n_30436), .Z(n_249886772));
	notech_ao4 i_135140010(.A(n_55886), .B(nbus_11295[30]), .C(n_227976218),
		 .D(n_30173), .Z(n_250086774));
	notech_ao4 i_134840013(.A(n_308084071), .B(nbus_11328[30]), .C(n_307884069
		), .D(n_30435), .Z(n_250286776));
	notech_and4 i_135040011(.A(n_249586769), .B(n_250286776), .C(n_246786741
		), .D(n_247086744), .Z(n_250586779));
	notech_ao4 i_134440017(.A(n_217486448), .B(n_28155), .C(n_248686760), .D
		(n_30434), .Z(n_250686780));
	notech_ao4 i_134340018(.A(n_55880), .B(nbus_11295[29]), .C(n_227976218),
		 .D(n_30174), .Z(n_250886782));
	notech_ao4 i_134040021(.A(n_308084071), .B(nbus_11328[29]), .C(n_307884069
		), .D(n_30433), .Z(n_251086784));
	notech_and4 i_134240019(.A(n_249586769), .B(n_251086784), .C(n_245886732
		), .D(n_246186735), .Z(n_251386787));
	notech_ao4 i_133640025(.A(n_217486448), .B(n_28154), .C(n_248686760), .D
		(n_30432), .Z(n_251486788));
	notech_ao4 i_133540026(.A(n_55880), .B(nbus_11295[28]), .C(n_227976218),
		 .D(n_30175), .Z(n_251686790));
	notech_ao4 i_133240029(.A(n_308084071), .B(nbus_11328[28]), .C(n_307884069
		), .D(n_30431), .Z(n_251886792));
	notech_and4 i_133440027(.A(n_249586769), .B(n_251886792), .C(n_244986723
		), .D(n_245286726), .Z(n_252186795));
	notech_ao4 i_132840033(.A(n_217486448), .B(n_28153), .C(n_248686760), .D
		(n_30430), .Z(n_252286796));
	notech_ao4 i_132740034(.A(n_55880), .B(n_57881), .C(n_227976218), .D(n_30176
		), .Z(n_252486798));
	notech_ao4 i_132440037(.A(n_308084071), .B(nbus_11328[27]), .C(n_307884069
		), .D(n_30429), .Z(n_252686800));
	notech_and4 i_132640035(.A(n_249586769), .B(n_252686800), .C(n_244086714
		), .D(n_244386717), .Z(n_252986803));
	notech_ao4 i_132040041(.A(n_217486448), .B(n_28152), .C(n_248686760), .D
		(n_30428), .Z(n_253086804));
	notech_ao4 i_131940042(.A(n_55880), .B(nbus_11295[26]), .C(n_57379), .D(n_30177
		), .Z(n_253286806));
	notech_ao4 i_131640045(.A(n_308084071), .B(nbus_11328[26]), .C(n_307884069
		), .D(n_30427), .Z(n_253486808));
	notech_and4 i_131840043(.A(n_249586769), .B(n_253486808), .C(n_243186705
		), .D(n_243486708), .Z(n_253786811));
	notech_ao4 i_131240049(.A(n_217486448), .B(n_28151), .C(n_248686760), .D
		(n_30426), .Z(n_253886812));
	notech_ao4 i_131140050(.A(n_55880), .B(nbus_11295[25]), .C(n_57375), .D(n_30178
		), .Z(n_254086814));
	notech_ao4 i_130840053(.A(n_308084071), .B(nbus_11328[25]), .C(n_307884069
		), .D(n_30425), .Z(n_254286816));
	notech_and4 i_131040051(.A(n_249586769), .B(n_254286816), .C(n_242586699
		), .D(n_242286696), .Z(n_254586819));
	notech_ao4 i_130340057(.A(n_217486448), .B(n_28150), .C(n_248686760), .D
		(n_30424), .Z(n_254686820));
	notech_ao4 i_130240058(.A(n_57375), .B(n_30179), .C(n_60373), .D(n_29402
		), .Z(n_254886822));
	notech_ao4 i_129940061(.A(n_307884069), .B(n_30423), .C(n_55880), .D(nbus_11295
		[24]), .Z(n_255086824));
	notech_and4 i_130140059(.A(n_249586769), .B(n_255086824), .C(n_241386687
		), .D(n_241686690), .Z(n_255386827));
	notech_ao4 i_129440065(.A(n_217486448), .B(n_28149), .C(n_248686760), .D
		(n_30422), .Z(n_255486828));
	notech_ao4 i_129340066(.A(n_57375), .B(n_30180), .C(n_60373), .D(n_29401
		), .Z(n_255686830));
	notech_ao4 i_129040069(.A(n_307884069), .B(n_30421), .C(n_55880), .D(nbus_11295
		[23]), .Z(n_255886832));
	notech_and4 i_129240067(.A(n_249586769), .B(n_255886832), .C(n_240486678
		), .D(n_240786681), .Z(n_256186835));
	notech_ao4 i_128440073(.A(n_217486448), .B(n_28148), .C(n_248686760), .D
		(n_30420), .Z(n_256286836));
	notech_ao4 i_128340074(.A(n_57379), .B(n_30181), .C(n_60367), .D(n_29400
		), .Z(n_256486838));
	notech_ao4 i_128040077(.A(n_307884069), .B(n_30419), .C(n_55880), .D(nbus_11295
		[22]), .Z(n_256686840));
	notech_and4 i_128240075(.A(n_249586769), .B(n_256686840), .C(n_239586669
		), .D(n_239886672), .Z(n_256986843));
	notech_ao4 i_127640081(.A(n_217486448), .B(n_28147), .C(n_248686760), .D
		(n_30418), .Z(n_257086844));
	notech_ao4 i_127540082(.A(n_57375), .B(n_30182), .C(n_60367), .D(n_29399
		), .Z(n_257286846));
	notech_ao4 i_127240085(.A(n_307884069), .B(n_30417), .C(n_55880), .D(nbus_11295
		[21]), .Z(n_257486848));
	notech_and4 i_127440083(.A(n_249586769), .B(n_257486848), .C(n_238686660
		), .D(n_238986663), .Z(n_257786851));
	notech_ao4 i_126840089(.A(n_217486448), .B(n_28146), .C(n_248686760), .D
		(n_30416), .Z(n_257886852));
	notech_ao4 i_126740090(.A(n_57375), .B(n_30183), .C(n_60367), .D(n_29398
		), .Z(n_258086854));
	notech_ao4 i_126340093(.A(n_307884069), .B(n_30414), .C(n_55880), .D(nbus_11295
		[20]), .Z(n_258286856));
	notech_and4 i_126540091(.A(n_249586769), .B(n_258286856), .C(n_237786651
		), .D(n_238086654), .Z(n_258586859));
	notech_ao4 i_125840097(.A(n_217486448), .B(n_28145), .C(n_248686760), .D
		(n_30413), .Z(n_258686860));
	notech_ao4 i_125740098(.A(n_57375), .B(n_30184), .C(n_60367), .D(n_29397
		), .Z(n_258886862));
	notech_ao4 i_125440101(.A(n_307884069), .B(n_30412), .C(n_55880), .D(nbus_11295
		[19]), .Z(n_259086864));
	notech_and4 i_125640099(.A(n_249586769), .B(n_259086864), .C(n_236886642
		), .D(n_237186645), .Z(n_259386867));
	notech_ao4 i_125040105(.A(n_217486448), .B(n_28144), .C(n_248686760), .D
		(n_30411), .Z(n_259486868));
	notech_ao4 i_124940106(.A(n_57375), .B(n_30185), .C(n_60367), .D(n_29396
		), .Z(n_259686870));
	notech_ao4 i_124640109(.A(n_307884069), .B(n_30410), .C(n_55880), .D(nbus_11295
		[18]), .Z(n_259886872));
	notech_and4 i_124840107(.A(n_249586769), .B(n_259886872), .C(n_235986633
		), .D(n_236286636), .Z(n_260186875));
	notech_ao4 i_123940113(.A(n_217486448), .B(n_28143), .C(n_248686760), .D
		(n_30409), .Z(n_260286876));
	notech_ao4 i_123840114(.A(n_57375), .B(n_30186), .C(n_60367), .D(n_29395
		), .Z(n_260486878));
	notech_ao4 i_123540117(.A(n_307884069), .B(n_30408), .C(n_55885), .D(nbus_11295
		[17]), .Z(n_260686880));
	notech_and4 i_123740115(.A(n_249586769), .B(n_260686880), .C(n_235086624
		), .D(n_235386627), .Z(n_260986883));
	notech_ao4 i_123140121(.A(n_217486448), .B(n_28142), .C(n_248686760), .D
		(n_30407), .Z(n_261086884));
	notech_ao4 i_123040122(.A(n_57375), .B(n_30187), .C(n_60367), .D(n_29394
		), .Z(n_261286886));
	notech_ao4 i_122740125(.A(n_55612), .B(n_30406), .C(n_55885), .D(nbus_11295
		[16]), .Z(n_261486888));
	notech_and4 i_122940123(.A(n_249586769), .B(n_261486888), .C(n_234186615
		), .D(n_234486618), .Z(n_261786891));
	notech_ao4 i_122040129(.A(n_217486448), .B(n_28141), .C(n_248686760), .D
		(n_30405), .Z(n_261886892));
	notech_ao4 i_121740130(.A(n_60367), .B(n_29393), .C(n_55592), .D(n_56275
		), .Z(n_261986893));
	notech_ao4 i_121540132(.A(n_3892), .B(nbus_11295[31]), .C(n_57375), .D(n_30188
		), .Z(n_262186895));
	notech_and4 i_122240127(.A(n_262186895), .B(n_261986893), .C(n_261886892
		), .D(n_233686610), .Z(n_262386897));
	notech_ao4 i_121240135(.A(n_308084071), .B(nbus_11328[15]), .C(n_55612),
		 .D(n_30404), .Z(n_262486898));
	notech_ao4 i_121040137(.A(n_307684067), .B(n_30017), .C(n_307584066), .D
		(n_28123), .Z(n_262686900));
	notech_and4 i_121440133(.A(n_249586769), .B(n_262686900), .C(n_262486898
		), .D(n_233386607), .Z(n_262886902));
	notech_ao4 i_120740140(.A(n_60367), .B(n_29392), .C(n_55592), .D(n_56248
		), .Z(n_262986903));
	notech_ao4 i_120640141(.A(n_55885), .B(n_56082), .C(n_57379), .D(n_30189
		), .Z(n_263086904));
	notech_ao4 i_120440143(.A(n_308084071), .B(nbus_11328[14]), .C(n_55612),
		 .D(n_30403), .Z(n_263286906));
	notech_and4 i_120940138(.A(n_263286906), .B(n_263086904), .C(n_262986903
		), .D(n_232486598), .Z(n_263486908));
	notech_ao4 i_120140146(.A(n_307584066), .B(n_28121), .C(n_3892), .D(nbus_11295
		[30]), .Z(n_263586909));
	notech_ao4 i_119940148(.A(n_307484065), .B(n_30402), .C(n_58651), .D(n_28140
		), .Z(n_263786911));
	notech_and4 i_120340144(.A(n_307384064), .B(n_263786911), .C(n_263586909
		), .D(n_232186595), .Z(n_263986913));
	notech_ao4 i_119640151(.A(n_60367), .B(n_29391), .C(n_55592), .D(n_56230
		), .Z(n_264086914));
	notech_ao4 i_119540152(.A(n_55885), .B(n_56073), .C(n_57379), .D(n_30190
		), .Z(n_264186915));
	notech_ao4 i_119340154(.A(n_308084071), .B(nbus_11328[13]), .C(n_55612),
		 .D(n_30401), .Z(n_264386917));
	notech_and4 i_119840149(.A(n_264386917), .B(n_264186915), .C(n_264086914
		), .D(n_231286586), .Z(n_264586919));
	notech_ao4 i_119040157(.A(n_28118), .B(n_307584066), .C(n_55900), .D(nbus_11295
		[29]), .Z(n_264686920));
	notech_ao4 i_118840159(.A(n_307484065), .B(n_30400), .C(n_58651), .D(n_28139
		), .Z(n_264886922));
	notech_and4 i_119240155(.A(n_307384064), .B(n_264886922), .C(n_264686920
		), .D(n_230986583), .Z(n_265086924));
	notech_ao4 i_118540162(.A(n_55885), .B(n_56064), .C(n_55592), .D(n_56221
		), .Z(n_265186925));
	notech_ao4 i_118440163(.A(n_57379), .B(n_30191), .C(n_60367), .D(n_29390
		), .Z(n_265286926));
	notech_ao4 i_118140165(.A(n_308084071), .B(nbus_11328[12]), .C(n_55612),
		 .D(n_30399), .Z(n_265486928));
	notech_and4 i_118740160(.A(n_265486928), .B(n_265286926), .C(n_265186925
		), .D(n_230086574), .Z(n_265686930));
	notech_ao4 i_117740168(.A(n_307584066), .B(n_28117), .C(n_55900), .D(nbus_11295
		[28]), .Z(n_265786931));
	notech_ao4 i_117440170(.A(n_307484065), .B(n_30398), .C(n_58651), .D(n_28138
		), .Z(n_265986933));
	notech_and4 i_118040166(.A(n_307384064), .B(n_265986933), .C(n_265786931
		), .D(n_229786571), .Z(n_266186935));
	notech_ao4 i_117140173(.A(n_60367), .B(n_29389), .C(n_55592), .D(n_56181
		), .Z(n_266286936));
	notech_ao4 i_117040174(.A(n_55885), .B(n_55983), .C(n_57379), .D(n_30192
		), .Z(n_266386937));
	notech_ao4 i_116840176(.A(n_55623), .B(nbus_11328[11]), .C(n_55612), .D(n_30397
		), .Z(n_266586939));
	notech_and4 i_117340171(.A(n_266586939), .B(n_266386937), .C(n_266286936
		), .D(n_228886562), .Z(n_266786941));
	notech_ao4 i_116540179(.A(n_307584066), .B(n_28116), .C(n_55900), .D(n_57881
		), .Z(n_266886942));
	notech_ao4 i_116340181(.A(n_307484065), .B(n_30396), .C(n_58651), .D(n_28137
		), .Z(n_267086944));
	notech_and4 i_116740177(.A(n_307384064), .B(n_267086944), .C(n_266886942
		), .D(n_228586559), .Z(n_267286946));
	notech_ao4 i_116040184(.A(n_60372), .B(n_29388), .C(n_55592), .D(n_56154
		), .Z(n_267386947));
	notech_ao4 i_115940185(.A(n_55885), .B(n_55992), .C(n_57379), .D(n_30193
		), .Z(n_267486948));
	notech_ao4 i_115740187(.A(n_55623), .B(nbus_11328[10]), .C(n_55612), .D(n_30395
		), .Z(n_267686950));
	notech_and4 i_116240182(.A(n_267686950), .B(n_267486948), .C(n_267386947
		), .D(n_227686550), .Z(n_267886952));
	notech_ao4 i_115240190(.A(n_307584066), .B(n_28115), .C(n_55900), .D(nbus_11295
		[26]), .Z(n_267986953));
	notech_ao4 i_115040192(.A(n_307484065), .B(n_30394), .C(n_58651), .D(n_28136
		), .Z(n_268186955));
	notech_and4 i_115640188(.A(n_307384064), .B(n_268186955), .C(n_267986953
		), .D(n_227386547), .Z(n_268386957));
	notech_ao4 i_114740195(.A(n_55885), .B(n_56010), .C(n_55592), .D(n_56136
		), .Z(n_268486958));
	notech_ao4 i_114640196(.A(n_57379), .B(n_30194), .C(n_60372), .D(n_29387
		), .Z(n_268586959));
	notech_ao4 i_114440198(.A(n_55623), .B(nbus_11328[9]), .C(n_55612), .D(n_30393
		), .Z(n_268786961));
	notech_and4 i_114940193(.A(n_268786961), .B(n_268586959), .C(n_268486958
		), .D(n_226486538), .Z(n_268986963));
	notech_ao4 i_114140201(.A(n_307584066), .B(n_28114), .C(n_55900), .D(nbus_11295
		[25]), .Z(n_269086964));
	notech_ao4 i_113940203(.A(n_307484065), .B(n_30392), .C(n_58651), .D(n_28135
		), .Z(n_269286966));
	notech_and4 i_114340199(.A(n_307384064), .B(n_269286966), .C(n_269086964
		), .D(n_226186535), .Z(n_269486968));
	notech_or4 i_2841228(.A(nbus_11295[1]), .B(n_59717), .C(nbus_11295[2]), 
		.D(n_57909), .Z(n_269586969));
	notech_nand2 i_88241280(.A(n_57406), .B(n_58675), .Z(n_269686970));
	notech_ao4 i_112740215(.A(n_217086444), .B(n_27055), .C(n_58697), .D(n_216986443
		), .Z(n_269786971));
	notech_ao4 i_112640216(.A(n_30391), .B(n_27378), .C(n_314863415), .D(n_30390
		), .Z(n_269886972));
	notech_ao4 i_112340219(.A(n_217486448), .B(n_28128), .C(n_248686760), .D
		(n_216386437), .Z(n_269986973));
	notech_ao4 i_112240220(.A(n_55592), .B(n_56064), .C(n_55900), .D(n_56221
		), .Z(n_270086974));
	notech_ao4 i_112040222(.A(n_57379), .B(n_30195), .C(n_60372), .D(n_29382
		), .Z(n_270286976));
	notech_and4 i_112540217(.A(n_270286976), .B(n_270086974), .C(n_269986973
		), .D(n_224886522), .Z(n_270486978));
	notech_ao4 i_111740225(.A(n_55623), .B(nbus_11328[4]), .C(n_55612), .D(n_30388
		), .Z(n_270586979));
	notech_ao4 i_111540227(.A(n_307684067), .B(n_29996), .C(n_307584066), .D
		(n_28109), .Z(n_270786981));
	notech_and4 i_111940223(.A(n_270786981), .B(n_270586979), .C(n_249586769
		), .D(n_224586519), .Z(n_270986983));
	notech_or4 i_128741261(.A(n_314463411), .B(n_60321), .C(n_18964), .D(n_27877
		), .Z(n_271086984));
	notech_or2 i_176641250(.A(n_271086984), .B(n_27378), .Z(n_271186985));
	notech_or2 i_45641282(.A(n_271086984), .B(n_58697), .Z(n_271286986));
	notech_or2 i_111440228(.A(n_271286986), .B(opc[3]), .Z(n_271386987));
	notech_or2 i_46241279(.A(n_271086984), .B(n_27055), .Z(n_271486988));
	notech_or4 i_46041281(.A(n_314463411), .B(n_60321), .C(n_18964), .D(n_27056
		), .Z(n_271686990));
	notech_ao4 i_111340229(.A(n_271286986), .B(n_27051), .C(n_216186435), .D
		(nbus_11295[2]), .Z(n_271786991));
	notech_ao4 i_110940233(.A(nbus_11295[3]), .B(n_216086434), .C(n_271386987
		), .D(n_290618105), .Z(n_271886992));
	notech_or2 i_46341278(.A(n_271086984), .B(n_314863415), .Z(n_272086994)
		);
	notech_ao4 i_110840234(.A(n_272086994), .B(n_30386), .C(n_271486988), .D
		(n_291118110), .Z(n_272186995));
	notech_ao3 i_111140231(.A(n_271886992), .B(n_272186995), .C(n_223886512)
		, .Z(n_272286996));
	notech_ao4 i_110640236(.A(n_55900), .B(\nbus_11358[11] ), .C(n_271686990
		), .D(n_27959), .Z(n_272386997));
	notech_ao4 i_110540237(.A(n_57379), .B(n_30196), .C(n_60372), .D(n_29381
		), .Z(n_272486998));
	notech_and3 i_111240230(.A(n_272486998), .B(n_272386997), .C(n_272286996
		), .Z(n_272687000));
	notech_ao4 i_110240240(.A(n_55623), .B(nbus_11328[3]), .C(n_30385), .D(n_55612
		), .Z(n_272787001));
	notech_ao4 i_110140241(.A(n_307984070), .B(n_57881), .C(n_55592), .D(n_55983
		), .Z(n_272887002));
	notech_ao4 i_109640243(.A(n_307684067), .B(n_29994), .C(n_307584066), .D
		(n_28108), .Z(n_273087004));
	notech_and3 i_109740242(.A(n_307384064), .B(n_273087004), .C(n_222386497
		), .Z(n_273287006));
	notech_ao4 i_109240245(.A(n_271486988), .B(n_291418113), .C(n_271286986)
		, .D(n_291218111), .Z(n_273487008));
	notech_mux2 i_108940248(.S(opc[2]), .A(n_215886432), .B(n_215786431), .Z
		(n_273587009));
	notech_ao4 i_108840249(.A(n_272086994), .B(n_30384), .C(n_271186985), .D
		(n_30383), .Z(n_273687010));
	notech_ao4 i_108640251(.A(n_60372), .B(n_29380), .C(n_55900), .D(n_56154
		), .Z(n_273887012));
	notech_ao4 i_108540252(.A(n_55612), .B(n_30382), .C(n_57379), .D(n_30197
		), .Z(n_273987013));
	notech_and4 i_109140246(.A(n_273987013), .B(n_273887012), .C(n_273687010
		), .D(n_273587009), .Z(n_274187015));
	notech_ao4 i_108140255(.A(n_55592), .B(n_55992), .C(nbus_11328[2]), .D(n_55623
		), .Z(n_274287016));
	notech_ao4 i_108040256(.A(n_307584066), .B(n_28107), .C(n_307984070), .D
		(nbus_11295[26]), .Z(n_274387017));
	notech_ao4 i_107840258(.A(n_58651), .B(n_28126), .C(n_307684067), .D(n_29988
		), .Z(n_274587019));
	notech_and4 i_108340253(.A(n_274587019), .B(n_274387017), .C(n_274287016
		), .D(n_307384064), .Z(n_274787021));
	notech_nand2 i_107740259(.A(nbus_11295[1]), .B(n_59735), .Z(n_274887022)
		);
	notech_ao4 i_107340263(.A(n_271486988), .B(n_215586429), .C(n_271286986)
		, .D(n_274887022), .Z(n_274987023));
	notech_ao4 i_107240264(.A(n_271186985), .B(n_30381), .C(n_215686430), .D
		(nbus_11295[1]), .Z(n_275187025));
	notech_ao4 i_107040266(.A(n_55900), .B(n_56136), .C(n_272086994), .D(n_30380
		), .Z(n_275387027));
	notech_ao4 i_106940267(.A(n_60372), .B(n_29379), .C(n_55592), .D(n_56010
		), .Z(n_275487028));
	notech_and4 i_107540261(.A(n_275487028), .B(n_275387027), .C(n_275187025
		), .D(n_274987023), .Z(n_275687030));
	notech_ao4 i_106640270(.A(n_55612), .B(n_30379), .C(n_57379), .D(n_30198
		), .Z(n_275787031));
	notech_ao4 i_106540271(.A(n_307984070), .B(nbus_11295[25]), .C(n_55623),
		 .D(nbus_11328[1]), .Z(n_275887032));
	notech_ao4 i_106340273(.A(n_307684067), .B(n_29986), .C(n_307584066), .D
		(n_28106), .Z(n_276087034));
	notech_and3 i_106440272(.A(n_307384064), .B(n_276087034), .C(n_219186465
		), .Z(n_276287036));
	notech_ao4 i_106140275(.A(n_30378), .B(n_314863415), .C(n_59735), .D(n_215386427
		), .Z(n_276487038));
	notech_ao4 i_105840278(.A(n_217486448), .B(n_28124), .C(n_248686760), .D
		(n_214986423), .Z(n_276587039));
	notech_ao4 i_105440279(.A(n_3892), .B(n_56118), .C(n_55885), .D(n_59717)
		, .Z(n_276687040));
	notech_ao4 i_105240281(.A(n_60372), .B(n_29378), .C(n_55592), .D(n_56028
		), .Z(n_276887042));
	notech_and2 i_105340280(.A(n_276887042), .B(n_218486458), .Z(n_276987043
		));
	notech_ao4 i_104940284(.A(n_55623), .B(nbus_11328[0]), .C(n_55612), .D(n_30377
		), .Z(n_277187045));
	notech_ao4 i_104740286(.A(n_307684067), .B(n_29983), .C(n_307584066), .D
		(n_28105), .Z(n_277387047));
	notech_and4 i_105140282(.A(n_277387047), .B(n_249586769), .C(n_277187045
		), .D(n_218186455), .Z(n_277587049));
	notech_nao3 i_6438178(.A(mul64[37]), .B(n_60321), .C(n_314563412), .Z(n_278487058
		));
	notech_nao3 i_7738165(.A(mul64[38]), .B(n_60321), .C(n_314563412), .Z(n_279787071
		));
	notech_or2 i_42837832(.A(n_55849), .B(n_60009), .Z(n_280687080));
	notech_or2 i_42537835(.A(n_55869), .B(n_57680), .Z(n_280987083));
	notech_or2 i_50637760(.A(n_60003), .B(n_55849), .Z(n_281887092));
	notech_or2 i_50337763(.A(n_55869), .B(n_57742), .Z(n_282187095));
	notech_or2 i_51837748(.A(n_60002), .B(n_55849), .Z(n_283087104));
	notech_or2 i_51537751(.A(n_55869), .B(n_57751), .Z(n_283387107));
	notech_or2 i_53037736(.A(n_60001), .B(n_55849), .Z(n_284287116));
	notech_or2 i_52737739(.A(n_55869), .B(n_57761), .Z(n_284587119));
	notech_or2 i_55437712(.A(n_133728614), .B(n_55849), .Z(n_285487128));
	notech_or2 i_55137715(.A(n_55869), .B(n_57783), .Z(n_285787131));
	notech_or2 i_56637700(.A(n_131228589), .B(n_55849), .Z(n_286687140));
	notech_or2 i_56337703(.A(n_55869), .B(n_57792), .Z(n_286987143));
	notech_or2 i_57837688(.A(n_130528582), .B(n_55849), .Z(n_287887152));
	notech_or2 i_57537691(.A(n_55869), .B(n_57802), .Z(n_288187155));
	notech_or2 i_59037676(.A(n_128228559), .B(n_55849), .Z(n_289087164));
	notech_or2 i_58737679(.A(n_55869), .B(\nbus_11365[29] ), .Z(n_289387167)
		);
	notech_or2 i_60237664(.A(n_302991794), .B(n_55849), .Z(n_290287176));
	notech_or2 i_59937667(.A(n_55869), .B(n_57828), .Z(n_290587179));
	notech_or2 i_61537651(.A(n_314791676), .B(n_55849), .Z(n_291487188));
	notech_or2 i_61237654(.A(n_55869), .B(n_59726), .Z(n_291787191));
	notech_ao4 i_169836608(.A(n_55791), .B(n_29030), .C(n_55782), .D(n_28123
		), .Z(n_292287196));
	notech_ao4 i_169736609(.A(n_310315179), .B(n_57837), .C(n_55800), .D(n_29085
		), .Z(n_292387197));
	notech_ao4 i_169536611(.A(n_55860), .B(n_29284), .C(n_55809), .D(nbus_11295
		[31]), .Z(n_292587199));
	notech_and4 i_170036606(.A(n_292587199), .B(n_292387197), .C(n_292287196
		), .D(n_291787191), .Z(n_292787201));
	notech_ao4 i_169236614(.A(n_55838), .B(n_29637), .C(n_55829), .D(n_28016
		), .Z(n_292887202));
	notech_and2 i_1938215(.A(n_276883759), .B(n_309115167), .Z(n_293087204)
		);
	notech_ao4 i_169036616(.A(n_55891), .B(n_29249), .C(n_52112621), .D(n_29217
		), .Z(n_293187205));
	notech_and4 i_169436612(.A(n_293087204), .B(n_293187205), .C(n_292887202
		), .D(n_291487188), .Z(n_293387207));
	notech_ao4 i_168736619(.A(n_55791), .B(n_29031), .C(n_55782), .D(n_28121
		), .Z(n_293487208));
	notech_ao4 i_168636620(.A(n_310315179), .B(n_55929), .C(n_55800), .D(n_29084
		), .Z(n_293587209));
	notech_ao4 i_168436622(.A(n_55860), .B(n_29283), .C(n_55809), .D(nbus_11295
		[30]), .Z(n_293787211));
	notech_and4 i_168936617(.A(n_293787211), .B(n_293587209), .C(n_293487208
		), .D(n_290587179), .Z(n_293987213));
	notech_ao4 i_168136625(.A(n_55838), .B(n_29665), .C(n_55829), .D(n_28015
		), .Z(n_294087214));
	notech_ao4 i_167936627(.A(n_55891), .B(n_29248), .C(n_52112621), .D(n_29216
		), .Z(n_294287216));
	notech_and4 i_168336623(.A(n_277183762), .B(n_294287216), .C(n_294087214
		), .D(n_290287176), .Z(n_294487218));
	notech_ao4 i_167636630(.A(n_55791), .B(n_29051), .C(n_55782), .D(n_28118
		), .Z(n_294587219));
	notech_ao4 i_167536631(.A(n_310315179), .B(\nbus_11358[29] ), .C(n_55800
		), .D(n_29083), .Z(n_294687220));
	notech_ao4 i_167336633(.A(n_55860), .B(n_29281), .C(n_55809), .D(nbus_11295
		[29]), .Z(n_294887222));
	notech_and4 i_167836628(.A(n_294887222), .B(n_294687220), .C(n_294587219
		), .D(n_289387167), .Z(n_295087224));
	notech_ao4 i_167036636(.A(n_55838), .B(n_29635), .C(n_55829), .D(n_28014
		), .Z(n_295187225));
	notech_ao4 i_166836638(.A(n_55891), .B(n_29247), .C(n_52112621), .D(n_29214
		), .Z(n_295387227));
	notech_and4 i_167236634(.A(n_277183762), .B(n_295387227), .C(n_295187225
		), .D(n_289087164), .Z(n_295587229));
	notech_ao4 i_166536641(.A(n_55791), .B(n_29050), .C(n_55782), .D(n_28117
		), .Z(n_295687230));
	notech_ao4 i_166436642(.A(n_310315179), .B(n_55974), .C(n_55800), .D(n_29082
		), .Z(n_295787231));
	notech_ao4 i_166236644(.A(n_55860), .B(n_29280), .C(n_55809), .D(nbus_11295
		[28]), .Z(n_295987233));
	notech_and4 i_166736639(.A(n_295987233), .B(n_295787231), .C(n_295687230
		), .D(n_288187155), .Z(n_296187235));
	notech_ao4 i_165936647(.A(n_55838), .B(n_29633), .C(n_55829), .D(n_28013
		), .Z(n_296287236));
	notech_ao4 i_165736649(.A(n_55891), .B(n_29246), .C(n_52112621), .D(n_29213
		), .Z(n_296487238));
	notech_and4 i_166136645(.A(n_293087204), .B(n_296487238), .C(n_296287236
		), .D(n_287887152), .Z(n_296687240));
	notech_ao4 i_165436652(.A(n_55791), .B(n_29034), .C(n_55782), .D(n_28116
		), .Z(n_296787241));
	notech_ao4 i_165336653(.A(n_310315179), .B(n_55938), .C(n_55800), .D(n_29081
		), .Z(n_296887242));
	notech_ao4 i_165136655(.A(n_55860), .B(n_29279), .C(n_55809), .D(n_57881
		), .Z(n_297087244));
	notech_and4 i_165636650(.A(n_297087244), .B(n_296887242), .C(n_296787241
		), .D(n_286987143), .Z(n_297287246));
	notech_ao4 i_164836658(.A(n_55838), .B(n_29639), .C(n_55829), .D(n_28012
		), .Z(n_297387247));
	notech_ao4 i_164636660(.A(n_55891), .B(n_29245), .C(n_52112621), .D(n_29211
		), .Z(n_297587249));
	notech_and4 i_165036656(.A(n_293087204), .B(n_297587249), .C(n_297387247
		), .D(n_286687140), .Z(n_297787251));
	notech_ao4 i_164336663(.A(n_55791), .B(n_29032), .C(n_55782), .D(n_28115
		), .Z(n_297887252));
	notech_ao4 i_164236664(.A(n_310315179), .B(n_55947), .C(n_55800), .D(n_29080
		), .Z(n_297987253));
	notech_ao4 i_164036666(.A(n_55860), .B(n_29278), .C(n_55809), .D(nbus_11295
		[26]), .Z(n_298187255));
	notech_and4 i_164536661(.A(n_298187255), .B(n_297987253), .C(n_297887252
		), .D(n_285787131), .Z(n_298387257));
	notech_ao4 i_163736669(.A(n_55838), .B(n_29667), .C(n_55829), .D(n_28011
		), .Z(n_298487258));
	notech_ao4 i_163536671(.A(n_55891), .B(n_29244), .C(n_52112621), .D(n_29210
		), .Z(n_298687260));
	notech_and4 i_163936667(.A(n_277183762), .B(n_298687260), .C(n_298487258
		), .D(n_285487128), .Z(n_298887262));
	notech_ao4 i_162136685(.A(n_55791), .B(n_29049), .C(n_55782), .D(n_28113
		), .Z(n_298987263));
	notech_ao4 i_162036686(.A(n_310315179), .B(n_56475), .C(n_55800), .D(n_29078
		), .Z(n_299087264));
	notech_ao4 i_161836688(.A(n_55860), .B(n_29276), .C(n_55809), .D(nbus_11295
		[24]), .Z(n_299287266));
	notech_and4 i_162336683(.A(n_299287266), .B(n_299087264), .C(n_298987263
		), .D(n_284587119), .Z(n_299487268));
	notech_ao4 i_161536691(.A(n_55838), .B(n_29641), .C(n_55829), .D(n_28009
		), .Z(n_299587269));
	notech_ao4 i_161336693(.A(n_55891), .B(n_29242), .C(n_52112621), .D(n_29206
		), .Z(n_299787271));
	notech_and4 i_161736689(.A(n_293087204), .B(n_299787271), .C(n_299587269
		), .D(n_284287116), .Z(n_299987273));
	notech_ao4 i_161036696(.A(n_55791), .B(n_29048), .C(n_55782), .D(n_28112
		), .Z(n_300087274));
	notech_ao4 i_160936697(.A(n_310315179), .B(n_56347), .C(n_55800), .D(n_29077
		), .Z(n_300187275));
	notech_ao4 i_160736699(.A(n_55860), .B(n_29275), .C(n_55809), .D(nbus_11295
		[23]), .Z(n_300387277));
	notech_and4 i_161236694(.A(n_300387277), .B(n_300187275), .C(n_300087274
		), .D(n_283387107), .Z(n_300587279));
	notech_ao4 i_160436702(.A(n_55838), .B(n_29638), .C(n_55829), .D(n_28008
		), .Z(n_300687280));
	notech_ao4 i_160236704(.A(n_55891), .B(n_29241), .C(n_52112621), .D(n_29205
		), .Z(n_300887282));
	notech_and4 i_160636700(.A(n_293087204), .B(n_300887282), .C(n_300687280
		), .D(n_283087104), .Z(n_301087284));
	notech_ao4 i_159936707(.A(n_55791), .B(n_29029), .C(n_55782), .D(n_28111
		), .Z(n_301187285));
	notech_ao4 i_159836708(.A(n_310315179), .B(n_56338), .C(n_55800), .D(n_29076
		), .Z(n_301287286));
	notech_ao4 i_159636710(.A(n_55860), .B(n_29274), .C(n_55809), .D(nbus_11295
		[22]), .Z(n_301487288));
	notech_and4 i_160136705(.A(n_301487288), .B(n_301287286), .C(n_301187285
		), .D(n_282187095), .Z(n_301687290));
	notech_ao4 i_159236713(.A(n_55838), .B(n_29666), .C(n_55829), .D(n_28007
		), .Z(n_301787291));
	notech_ao4 i_159036715(.A(n_55891), .B(n_29239), .C(n_52112621), .D(n_29203
		), .Z(n_301987293));
	notech_and4 i_159536711(.A(n_277183762), .B(n_301987293), .C(n_301787291
		), .D(n_281887092), .Z(n_302187295));
	notech_ao4 i_153236773(.A(n_55791), .B(n_29047), .C(n_55782), .D(n_28105
		), .Z(n_302287296));
	notech_ao4 i_153136774(.A(n_310315179), .B(n_56284), .C(n_55800), .D(n_29069
		), .Z(n_302387297));
	notech_ao4 i_152936776(.A(n_55860), .B(n_29268), .C(n_55809), .D(nbus_11295
		[16]), .Z(n_302587299));
	notech_and4 i_153436771(.A(n_302587299), .B(n_302387297), .C(n_302287296
		), .D(n_280987083), .Z(n_302787301));
	notech_ao4 i_152636779(.A(n_55838), .B(n_29642), .C(n_55829), .D(n_28001
		), .Z(n_302887302));
	notech_ao4 i_152436781(.A(n_55891), .B(n_29233), .C(n_52112621), .D(n_29195
		), .Z(n_303087304));
	notech_and4 i_152836777(.A(n_303087304), .B(n_302887302), .C(n_293087204
		), .D(n_280687080), .Z(n_303287306));
	notech_ao4 i_121037092(.A(n_307984070), .B(nbus_11295[30]), .C(n_55900),
		 .D(n_56248), .Z(n_303387307));
	notech_ao4 i_120937093(.A(n_55885), .B(nbus_11295[6]), .C(n_307584066), 
		.D(n_28111), .Z(n_303487308));
	notech_ao4 i_120737095(.A(n_60372), .B(n_29384), .C(n_55592), .D(n_56082
		), .Z(n_303687310));
	notech_and4 i_121237090(.A(n_303687310), .B(n_303487308), .C(n_303387307
		), .D(n_279787071), .Z(n_303887312));
	notech_ao4 i_120437098(.A(n_55623), .B(nbus_11328[6]), .C(n_55612), .D(n_30445
		), .Z(n_303987313));
	notech_ao4 i_120337099(.A(n_307684067), .B(n_30000), .C(n_58651), .D(n_28131
		), .Z(n_304087314));
	notech_ao4 i_120137101(.A(n_309987373), .B(n_30444), .C(n_309887372), .D
		(n_30443), .Z(n_304287316));
	notech_and4 i_120637096(.A(n_307384064), .B(n_304287316), .C(n_304087314
		), .D(n_303987313), .Z(n_304487318));
	notech_ao4 i_119837104(.A(n_307984070), .B(nbus_11295[29]), .C(n_55900),
		 .D(n_56230), .Z(n_304587319));
	notech_ao4 i_119737105(.A(n_55885), .B(nbus_11295[5]), .C(n_307584066), 
		.D(n_28110), .Z(n_304687320));
	notech_ao4 i_119537107(.A(n_60372), .B(n_29383), .C(n_55592), .D(n_56073
		), .Z(n_304887322));
	notech_and4 i_120037102(.A(n_304887322), .B(n_304687320), .C(n_304587319
		), .D(n_278487058), .Z(n_305087324));
	notech_ao4 i_119237110(.A(n_55623), .B(nbus_11328[5]), .C(n_55612), .D(n_30441
		), .Z(n_305187325));
	notech_ao4 i_119137111(.A(n_307684067), .B(n_29998), .C(n_58651), .D(n_28129
		), .Z(n_305287326));
	notech_ao4 i_118937113(.A(n_309987373), .B(n_30440), .C(n_309887372), .D
		(n_30439), .Z(n_305487328));
	notech_and4 i_119437108(.A(n_307384064), .B(n_305487328), .C(n_305287326
		), .D(n_305187325), .Z(n_305687330));
	notech_and2 i_15834953(.A(n_32446), .B(n_306187335), .Z(n_305787331));
	notech_and3 i_15434957(.A(n_304984040), .B(n_304484035), .C(n_305987333)
		, .Z(n_305887332));
	notech_or4 i_19034921(.A(n_2839), .B(n_2888), .C(n_60868), .D(n_58812), 
		.Z(n_305987333));
	notech_or4 i_102434111(.A(n_27994), .B(n_2839), .C(n_1864), .D(n_3866), 
		.Z(n_306087334));
	notech_or4 i_107934056(.A(n_27994), .B(n_2839), .C(n_60863), .D(n_57818)
		, .Z(n_306187335));
	notech_or2 i_112734008(.A(n_306587339), .B(n_27063), .Z(n_306487338));
	notech_ao4 i_3935071(.A(n_61103), .B(n_25651), .C(n_59451), .D(n_308012096
		), .Z(n_306587339));
	notech_nao3 i_17334938(.A(Daddrs_3[11]), .B(n_32562), .C(n_3790), .Z(n_307087344
		));
	notech_nao3 i_17034941(.A(n_11278), .B(n_60321), .C(n_1893), .Z(n_307387347
		));
	notech_or2 i_16734944(.A(n_55367), .B(n_28398), .Z(n_307687350));
	notech_nao3 i_16434947(.A(n_11277), .B(n_60321), .C(n_304384034), .Z(n_307987353
		));
	notech_or4 i_102234113(.A(n_32729), .B(n_27573), .C(n_59424), .D(n_30448
		), .Z(n_308287356));
	notech_or2 i_102334112(.A(n_2985), .B(n_3865), .Z(n_308387357));
	notech_or4 i_103134104(.A(n_60883), .B(n_60223), .C(n_58033), .D(nbus_11295
		[31]), .Z(n_309287366));
	notech_nor2 i_23146(.A(n_3904), .B(n_305787331), .Z(n_309787371));
	notech_or4 i_36068(.A(n_18964), .B(n_314463411), .C(n_60321), .D(n_27378
		), .Z(n_309887372));
	notech_or4 i_36066(.A(n_314463411), .B(n_18964), .C(n_60321), .D(rep_en1
		), .Z(n_309987373));
	notech_or4 i_111034025(.A(n_60883), .B(n_61103), .C(n_27988), .D(n_27880
		), .Z(n_310087374));
	notech_or4 i_111134024(.A(n_32747), .B(n_62892), .C(n_27573), .D(n_27084
		), .Z(n_310187375));
	notech_or4 i_112534010(.A(n_60888), .B(n_61103), .C(n_310587379), .D(\opcode[0] 
		), .Z(n_310287376));
	notech_ao3 i_112634009(.A(mask8b[2]), .B(read_ack), .C(n_107111189), .Z(n_310387377
		));
	notech_or4 i_208133072(.A(n_27170), .B(n_32443), .C(n_32695), .D(n_32730
		), .Z(n_310587379));
	notech_ao4 i_7335037(.A(n_61103), .B(n_1893), .C(n_306587339), .D(n_58812
		), .Z(n_311187385));
	notech_ao4 i_195033203(.A(n_309887372), .B(n_30452), .C(n_57379), .D(n_30200
		), .Z(n_311287386));
	notech_ao4 i_194933204(.A(n_307584066), .B(n_28112), .C(n_309987373), .D
		(n_30450), .Z(n_311387387));
	notech_ao4 i_194733206(.A(n_55612), .B(n_30449), .C(n_307684067), .D(n_30002
		), .Z(n_311587389));
	notech_and4 i_195233201(.A(n_311587389), .B(n_311387387), .C(n_311287386
		), .D(n_309287366), .Z(n_311787391));
	notech_ao4 i_194433209(.A(n_55885), .B(nbus_11295[7]), .C(n_55623), .D(nbus_11328
		[7]), .Z(n_311887392));
	notech_ao4 i_194333210(.A(n_58651), .B(n_28133), .C(n_55900), .D(n_56275
		), .Z(n_311987393));
	notech_ao4 i_194133212(.A(n_60372), .B(n_29385), .C(n_55592), .D(n_56109
		), .Z(n_312187395));
	notech_and4 i_194633207(.A(n_307384064), .B(n_312187395), .C(n_311987393
		), .D(n_311887392), .Z(n_312387397));
	notech_ao4 i_117233964(.A(n_57716), .B(read_ack), .C(n_61103), .D(n_305887332
		), .Z(n_312687400));
	notech_ao4 i_115033986(.A(n_55347), .B(nbus_11295[11]), .C(n_55409), .D(n_30446
		), .Z(n_312987403));
	notech_ao4 i_114833988(.A(n_55389), .B(n_28604), .C(n_55378), .D(n_29357
		), .Z(n_313187405));
	notech_and4 i_115233984(.A(n_313187405), .B(n_312987403), .C(n_307687350
		), .D(n_307987353), .Z(n_313387407));
	notech_ao4 i_114533991(.A(n_55400), .B(n_27996), .C(n_55429), .D(n_56181
		), .Z(n_313487408));
	notech_ao4 i_114333993(.A(n_59147), .B(n_29295), .C(n_59176), .D(n_27814
		), .Z(n_313687410));
	notech_and4 i_114733989(.A(n_313687410), .B(n_313487408), .C(n_307087344
		), .D(n_307387347), .Z(n_313887412));
	notech_and4 i_35932440(.A(n_32458), .B(n_1869), .C(n_331163528), .D(n_18906874
		), .Z(n_313987413));
	notech_ao4 i_36032439(.A(n_27037), .B(n_27145), .C(read_ack), .D(n_27068
		), .Z(n_314087414));
	notech_nand3 i_32732463(.A(n_316087434), .B(n_316787441), .C(n_316187435
		), .Z(n_314287416));
	notech_mux2 i_25432520(.S(all_cnt[0]), .A(n_3921), .B(n_56888), .Z(n_314387417
		));
	notech_mux4 i_29632487(.S0(all_cnt[1]), .S1(all_cnt[0]), .A(n_27107), .B
		(n_54929), .C(n_56391), .D(n_3914), .Z(n_314487418));
	notech_and4 i_37467(.A(n_60136), .B(n_323384224), .C(n_320491619), .D(n_318591638
		), .Z(n_315787431));
	notech_and4 i_68132157(.A(read_ack), .B(n_18981), .C(n_61560), .D(n_32551
		), .Z(n_315887432));
	notech_nao3 i_68232156(.A(n_61560), .B(n_314287416), .C(n_5968810), .Z(n_315987433
		));
	notech_or4 i_68532153(.A(all_cnt[0]), .B(all_cnt[3]), .C(n_27090), .D(n_27113
		), .Z(n_316087434));
	notech_nand3 i_68632152(.A(n_6888902), .B(n_30976), .C(n_3673), .Z(n_316187435
		));
	notech_nao3 i_125831626(.A(all_cnt[2]), .B(n_27853), .C(all_cnt[3]), .Z(n_316687440
		));
	notech_ao4 i_125731627(.A(n_314487418), .B(n_27070), .C(n_314387417), .D
		(n_316687440), .Z(n_316787441));
	notech_ao4 i_79832049(.A(n_27069), .B(n_314087414), .C(n_61103), .D(n_313987413
		), .Z(n_317087444));
	notech_and4 i_79632051(.A(n_53731), .B(n_315787431), .C(n_17779989), .D(n_320263469
		), .Z(n_317587449));
	notech_ao4 i_141360388(.A(n_308591738), .B(n_28006), .C(n_150228779), .D
		(n_59980), .Z(n_200359084));
	notech_or4 i_17461(.A(n_61103), .B(n_310587379), .C(n_60888), .D(n_32747
		), .Z(n_317687450));
	notech_or4 i_17837(.A(n_60863), .B(n_61103), .C(n_69641311), .D(n_32747)
		, .Z(n_317787451));
	notech_and4 i_142160380(.A(n_200059081), .B(n_199859079), .C(n_199759078
		), .D(n_199159073), .Z(n_200259083));
	notech_mux2 i_35867400(.S(n_60321), .A(n_19014), .B(n_106585342), .Z(n_317887452
		));
	notech_ao3 i_17463(.A(n_2885), .B(opb[1]), .C(n_61156), .Z(n_317987453)
		);
	notech_ao3 i_17465(.A(n_2885), .B(opb[3]), .C(n_61156), .Z(n_318087454)
		);
	notech_ao3 i_17466(.A(n_2885), .B(opb[4]), .C(n_61156), .Z(n_318187455)
		);
	notech_ao3 i_17468(.A(n_2885), .B(opb[6]), .C(n_61156), .Z(n_318287456)
		);
	notech_ao3 i_17469(.A(n_2885), .B(opb[7]), .C(n_61156), .Z(n_318387457)
		);
	notech_ao3 i_17470(.A(n_2885), .B(opb[8]), .C(n_61156), .Z(n_318487458)
		);
	notech_ao3 i_17471(.A(n_2885), .B(opb[9]), .C(n_61156), .Z(n_318587459)
		);
	notech_ao3 i_17472(.A(n_2885), .B(opb[10]), .C(n_61156), .Z(n_318687460)
		);
	notech_ao3 i_17473(.A(n_60378), .B(opb[11]), .C(n_61156), .Z(n_318787461
		));
	notech_ao3 i_17474(.A(n_60378), .B(opb[12]), .C(n_61149), .Z(n_318887462
		));
	notech_ao3 i_17475(.A(n_60378), .B(opb[13]), .C(n_61149), .Z(n_318987463
		));
	notech_ao3 i_17476(.A(n_60378), .B(opb[14]), .C(n_61149), .Z(n_319087464
		));
	notech_ao3 i_17477(.A(n_60378), .B(opb[15]), .C(n_61149), .Z(n_319187465
		));
	notech_and2 i_17942(.A(regs_10[0]), .B(n_161285889), .Z(n_319287466));
	notech_and2 i_17944(.A(n_161285889), .B(regs_10[1]), .Z(n_319387467));
	notech_and2 i_17945(.A(n_161285889), .B(regs_10[2]), .Z(n_319487468));
	notech_and2 i_17946(.A(n_161285889), .B(regs_10[3]), .Z(n_319587469));
	notech_and2 i_17947(.A(n_161285889), .B(regs_10[4]), .Z(n_319687470));
	notech_and2 i_17948(.A(n_161285889), .B(regs_10[5]), .Z(n_319787471));
	notech_and2 i_17949(.A(n_161285889), .B(regs_10[6]), .Z(n_319887472));
	notech_and2 i_17950(.A(n_161285889), .B(regs_10[7]), .Z(n_319987473));
	notech_and2 i_17951(.A(n_161285889), .B(regs_10[8]), .Z(n_320087474));
	notech_and2 i_17952(.A(n_161285889), .B(regs_10[9]), .Z(n_320187475));
	notech_and2 i_17953(.A(n_161285889), .B(regs_10[10]), .Z(n_320287476));
	notech_and2 i_17954(.A(n_161285889), .B(regs_10[11]), .Z(n_320387477));
	notech_and2 i_17955(.A(n_161285889), .B(regs_10[12]), .Z(n_320487478));
	notech_and2 i_17956(.A(n_161285889), .B(regs_10[13]), .Z(n_320587479));
	notech_and2 i_17957(.A(n_161285889), .B(regs_10[14]), .Z(n_320687480));
	notech_and2 i_17958(.A(n_53259), .B(regs_10[15]), .Z(n_320787481));
	notech_and2 i_17959(.A(n_53259), .B(regs_10[16]), .Z(n_320887482));
	notech_and2 i_17961(.A(n_53259), .B(regs_10[18]), .Z(n_320987483));
	notech_and2 i_17962(.A(n_53259), .B(regs_10[19]), .Z(n_321087484));
	notech_and2 i_17963(.A(n_53259), .B(regs_10[20]), .Z(n_321187485));
	notech_and2 i_17964(.A(n_53259), .B(regs_10[21]), .Z(n_321287486));
	notech_and2 i_17965(.A(n_53259), .B(regs_10[22]), .Z(n_321387487));
	notech_and2 i_17966(.A(n_53259), .B(regs_10[23]), .Z(n_321487488));
	notech_and2 i_17967(.A(n_53259), .B(regs_10[24]), .Z(n_321587489));
	notech_and2 i_17968(.A(n_53259), .B(regs_10[25]), .Z(n_321687490));
	notech_and2 i_17969(.A(n_53259), .B(regs_10[26]), .Z(n_321787491));
	notech_and2 i_17970(.A(n_53259), .B(regs_10[27]), .Z(n_321887492));
	notech_and2 i_17971(.A(n_53259), .B(regs_10[28]), .Z(n_321987493));
	notech_and2 i_17972(.A(n_53259), .B(regs_10[29]), .Z(n_322087494));
	notech_and2 i_17973(.A(n_53259), .B(regs_10[30]), .Z(n_322187495));
	notech_and2 i_17974(.A(n_53259), .B(regs_10[31]), .Z(n_322287496));
	notech_nor2 i_26926(.A(n_268643294), .B(n_60223), .Z(n_322387497));
	notech_ao3 i_26931(.A(n_60113), .B(n_60319), .C(n_330463521), .Z(n_322487498
		));
	notech_nand2 i_3327512(.A(n_194286216), .B(n_168085957), .Z(n_13531));
	notech_nand2 i_3227511(.A(n_194486218), .B(n_194386217), .Z(n_13526));
	notech_nand2 i_3127510(.A(n_194686220), .B(n_194586219), .Z(n_13521));
	notech_nand2 i_3027509(.A(n_194886222), .B(n_194786221), .Z(n_13516));
	notech_nand2 i_2927508(.A(n_195086224), .B(n_194986223), .Z(n_13511));
	notech_nand2 i_2827507(.A(n_195286226), .B(n_195186225), .Z(n_13506));
	notech_nand2 i_2727506(.A(n_195486228), .B(n_195386227), .Z(n_13501));
	notech_nand2 i_2627505(.A(n_195686230), .B(n_195586229), .Z(n_13496));
	notech_nand2 i_2527504(.A(n_195886232), .B(n_195786231), .Z(n_13491));
	notech_nand2 i_2427503(.A(n_196086234), .B(n_195986233), .Z(n_13486));
	notech_nand2 i_2327502(.A(n_196286236), .B(n_196186235), .Z(n_13481));
	notech_nand2 i_2227501(.A(n_196486238), .B(n_196386237), .Z(n_13476));
	notech_nand2 i_2127500(.A(n_196686240), .B(n_196586239), .Z(n_13471));
	notech_nand2 i_2027499(.A(n_196886242), .B(n_196786241), .Z(n_13466));
	notech_nand2 i_1927498(.A(n_197086244), .B(n_196986243), .Z(n_13461));
	notech_nand2 i_1827497(.A(n_197286246), .B(n_197186245), .Z(n_13456));
	notech_nand2 i_1727496(.A(n_197486248), .B(n_197386247), .Z(n_13451));
	notech_nand2 i_1627495(.A(n_197686250), .B(n_197586249), .Z(n_13446));
	notech_nand2 i_1527494(.A(n_197886252), .B(n_197786251), .Z(n_13441));
	notech_nand2 i_1427493(.A(n_198086254), .B(n_197986253), .Z(n_13436));
	notech_nand2 i_1327492(.A(n_198286256), .B(n_198186255), .Z(n_13431));
	notech_nand2 i_1227491(.A(n_198486258), .B(n_198386257), .Z(n_13426));
	notech_nand2 i_1127490(.A(n_198686260), .B(n_198586259), .Z(n_13421));
	notech_nand2 i_1027489(.A(n_198886262), .B(n_198786261), .Z(n_13416));
	notech_nand2 i_927488(.A(n_199086264), .B(n_198986263), .Z(n_13411));
	notech_nand2 i_827487(.A(n_199286266), .B(n_199186265), .Z(n_13406));
	notech_nand2 i_727486(.A(n_199486268), .B(n_199386267), .Z(n_13401));
	notech_nand2 i_627485(.A(n_199686270), .B(n_199586269), .Z(n_13396));
	notech_nand2 i_527484(.A(n_199886272), .B(n_199786271), .Z(n_13391));
	notech_nand2 i_427483(.A(n_200086274), .B(n_199986273), .Z(n_13386));
	notech_nand2 i_327482(.A(n_200286276), .B(n_200186275), .Z(n_13381));
	notech_nand2 i_227481(.A(n_200486278), .B(n_200386277), .Z(n_13376));
	notech_nand2 i_127480(.A(n_200586279), .B(n_167785954), .Z(n_13371));
	notech_nand2 i_6427415(.A(n_200686280), .B(n_167685953), .Z(n_21985));
	notech_nand2 i_6327414(.A(n_200786281), .B(n_167585952), .Z(n_21980));
	notech_nand2 i_6227413(.A(n_200886282), .B(n_167485951), .Z(n_21975));
	notech_nand2 i_6127412(.A(n_200986283), .B(n_167385950), .Z(n_21970));
	notech_nand2 i_6027411(.A(n_201086284), .B(n_167285949), .Z(n_21965));
	notech_nand2 i_5927410(.A(n_201186285), .B(n_167185948), .Z(n_21960));
	notech_nand2 i_5827409(.A(n_201286286), .B(n_167085947), .Z(n_21955));
	notech_nand2 i_5727408(.A(n_201386287), .B(n_166985946), .Z(n_21950));
	notech_nand2 i_5627407(.A(n_201486288), .B(n_166885945), .Z(n_21945));
	notech_nand2 i_5527406(.A(n_201586289), .B(n_166785944), .Z(n_21940));
	notech_nand2 i_5427405(.A(n_201686290), .B(n_166685943), .Z(n_21935));
	notech_nand2 i_5327404(.A(n_201786291), .B(n_166585942), .Z(n_21930));
	notech_nand2 i_5227403(.A(n_201886292), .B(n_166485941), .Z(n_21925));
	notech_nand2 i_5127402(.A(n_201986293), .B(n_166385940), .Z(n_21920));
	notech_nand2 i_5027401(.A(n_202086294), .B(n_166285939), .Z(n_21915));
	notech_nand2 i_4927400(.A(n_202186295), .B(n_166185938), .Z(n_21910));
	notech_nand2 i_4827399(.A(n_202286296), .B(n_166085937), .Z(n_21905));
	notech_nand2 i_4727398(.A(n_202386297), .B(n_165985936), .Z(n_21900));
	notech_nand2 i_4627397(.A(n_202486298), .B(n_165885935), .Z(n_21895));
	notech_nand2 i_4527396(.A(n_202586299), .B(n_165785934), .Z(n_21890));
	notech_nand2 i_4427395(.A(n_202686300), .B(n_165685933), .Z(n_21885));
	notech_nand2 i_4327394(.A(n_202786301), .B(n_165585932), .Z(n_21880));
	notech_nand2 i_4227393(.A(n_202886302), .B(n_165485931), .Z(n_21875));
	notech_nand2 i_4127392(.A(n_202986303), .B(n_165385930), .Z(n_21870));
	notech_nand2 i_4027391(.A(n_203086304), .B(n_165285929), .Z(n_21865));
	notech_nand2 i_3927390(.A(n_203186305), .B(n_165185928), .Z(n_21860));
	notech_nand2 i_3827389(.A(n_203286306), .B(n_165085927), .Z(n_21855));
	notech_nand2 i_3727388(.A(n_203386307), .B(n_164985926), .Z(n_21850));
	notech_nand2 i_3627387(.A(n_203486308), .B(n_164885925), .Z(n_21845));
	notech_nand2 i_3527386(.A(n_203586309), .B(n_164785924), .Z(n_21840));
	notech_nand2 i_3427385(.A(n_203686310), .B(n_164685923), .Z(n_21835));
	notech_nand2 i_3327384(.A(n_203786311), .B(n_164585922), .Z(n_21830));
	notech_nand2 i_3227383(.A(n_203886312), .B(n_164485921), .Z(n_21825));
	notech_nand2 i_3127382(.A(n_203986313), .B(n_164385920), .Z(n_21820));
	notech_nand2 i_3027381(.A(n_204086314), .B(n_164285919), .Z(n_21815));
	notech_nand2 i_2927380(.A(n_204186315), .B(n_164185918), .Z(n_21810));
	notech_nand2 i_2827379(.A(n_204286316), .B(n_164085917), .Z(n_21805));
	notech_nand2 i_2727378(.A(n_204386317), .B(n_163985916), .Z(n_21800));
	notech_nand2 i_2627377(.A(n_204486318), .B(n_163885915), .Z(n_21795));
	notech_nand2 i_2527376(.A(n_204586319), .B(n_163785914), .Z(n_21790));
	notech_nand2 i_2427375(.A(n_204686320), .B(n_163685913), .Z(n_21785));
	notech_nand2 i_2327374(.A(n_204786321), .B(n_163585912), .Z(n_21780));
	notech_nand2 i_2227373(.A(n_204886322), .B(n_163485911), .Z(n_21775));
	notech_nand2 i_2127372(.A(n_204986323), .B(n_163385910), .Z(n_21770));
	notech_nand2 i_1927370(.A(n_205086324), .B(n_163285909), .Z(n_21760));
	notech_nand2 i_1827369(.A(n_205186325), .B(n_163185908), .Z(n_21755));
	notech_nand2 i_1727368(.A(n_205286326), .B(n_163085907), .Z(n_21750));
	notech_nand2 i_1627367(.A(n_205386327), .B(n_162985906), .Z(n_21745));
	notech_nand2 i_1527366(.A(n_205486328), .B(n_162885905), .Z(n_21740));
	notech_nand2 i_1427365(.A(n_205586329), .B(n_162785904), .Z(n_21735));
	notech_nand2 i_1327364(.A(n_205686330), .B(n_162685903), .Z(n_21730));
	notech_nand2 i_1227363(.A(n_205786331), .B(n_162585902), .Z(n_21725));
	notech_nand2 i_1127362(.A(n_205886332), .B(n_162485901), .Z(n_21720));
	notech_nand2 i_1027361(.A(n_205986333), .B(n_162385900), .Z(n_21715));
	notech_nand2 i_927360(.A(n_206086334), .B(n_162285899), .Z(n_21710));
	notech_nand2 i_827359(.A(n_206186335), .B(n_162185898), .Z(n_21705));
	notech_nand2 i_727358(.A(n_206286336), .B(n_162085897), .Z(n_21700));
	notech_nand2 i_627357(.A(n_206386337), .B(n_161985896), .Z(n_21695));
	notech_nand2 i_527356(.A(n_206486338), .B(n_161885895), .Z(n_21690));
	notech_nand2 i_427355(.A(n_206586339), .B(n_161785894), .Z(n_21685));
	notech_nand2 i_327354(.A(n_206686340), .B(n_161685893), .Z(n_21680));
	notech_nand2 i_227353(.A(n_206786341), .B(n_161585892), .Z(n_21675));
	notech_nand2 i_127352(.A(n_206886342), .B(n_161485891), .Z(n_21670));
	notech_ao4 i_141660385(.A(n_150528782), .B(n_56329), .C(n_150728784), .D
		(n_60004), .Z(n_200059081));
	notech_ao4 i_141860383(.A(n_60117), .B(n_27141), .C(n_3836), .D(n_57733)
		, .Z(n_199859079));
	notech_ao4 i_141960382(.A(n_308791736), .B(n_110964638), .C(n_306791756)
		, .D(n_111164640), .Z(n_199759078));
	notech_nand2 i_323102(.A(n_57440), .B(n_209986373), .Z(n_16501));
	notech_and4 i_218967(.A(n_210486378), .B(n_211186385), .C(n_209286366), 
		.D(n_210386377), .Z(n_25494));
	notech_and4 i_118966(.A(n_211586389), .B(n_212286396), .C(n_208086354), 
		.D(n_211486388), .Z(n_25488));
	notech_nand2 i_126970(.A(n_214886422), .B(n_26648), .Z(n_14515));
	notech_and4 i_3217205(.A(n_248886762), .B(n_249086764), .C(n_249786771),
		 .D(n_248486758), .Z(n_15176));
	notech_and4 i_3117204(.A(n_249886772), .B(n_250086774), .C(n_250586779),
		 .D(n_247586749), .Z(n_15171));
	notech_and4 i_3017203(.A(n_250686780), .B(n_250886782), .C(n_251386787),
		 .D(n_246686740), .Z(n_15166));
	notech_and4 i_2917202(.A(n_251486788), .B(n_251686790), .C(n_252186795),
		 .D(n_245786731), .Z(n_15161));
	notech_and4 i_2817201(.A(n_252286796), .B(n_252486798), .C(n_252986803),
		 .D(n_244886722), .Z(n_15156));
	notech_and4 i_2717200(.A(n_253086804), .B(n_253286806), .C(n_253786811),
		 .D(n_243986713), .Z(n_15151));
	notech_and4 i_2617199(.A(n_253886812), .B(n_254086814), .C(n_254586819),
		 .D(n_243086704), .Z(n_15146));
	notech_and4 i_2517198(.A(n_254686820), .B(n_254886822), .C(n_255386827),
		 .D(n_242186695), .Z(n_15141));
	notech_and4 i_2417197(.A(n_255486828), .B(n_255686830), .C(n_256186835),
		 .D(n_241286686), .Z(n_15136));
	notech_and4 i_2317196(.A(n_256286836), .B(n_256486838), .C(n_256986843),
		 .D(n_240386677), .Z(n_15131));
	notech_and4 i_2217195(.A(n_257086844), .B(n_257286846), .C(n_257786851),
		 .D(n_239486668), .Z(n_15126));
	notech_and4 i_2117194(.A(n_257886852), .B(n_258086854), .C(n_258586859),
		 .D(n_238586659), .Z(n_15121));
	notech_and4 i_2017193(.A(n_258686860), .B(n_258886862), .C(n_259386867),
		 .D(n_237686650), .Z(n_15116));
	notech_and4 i_1917192(.A(n_259486868), .B(n_259686870), .C(n_260186875),
		 .D(n_236786641), .Z(n_15111));
	notech_and4 i_1817191(.A(n_260286876), .B(n_260486878), .C(n_260986883),
		 .D(n_235886632), .Z(n_15106));
	notech_and4 i_1717190(.A(n_261086884), .B(n_261286886), .C(n_261786891),
		 .D(n_234986623), .Z(n_15101));
	notech_nand2 i_1617189(.A(n_262886902), .B(n_262386897), .Z(n_15096));
	notech_nand2 i_1517188(.A(n_263986913), .B(n_263486908), .Z(n_15091));
	notech_nand2 i_1417187(.A(n_265086924), .B(n_264586919), .Z(n_15086));
	notech_nand2 i_1317186(.A(n_266186935), .B(n_265686930), .Z(n_15081));
	notech_nand2 i_1217185(.A(n_267286946), .B(n_266786941), .Z(n_15076));
	notech_nand2 i_1117184(.A(n_268386957), .B(n_267886952), .Z(n_15071));
	notech_nand2 i_1017183(.A(n_269486968), .B(n_268986963), .Z(n_15066));
	notech_nand2 i_517178(.A(n_270986983), .B(n_270486978), .Z(n_15041));
	notech_and4 i_417177(.A(n_272887002), .B(n_272787001), .C(n_272687000), 
		.D(n_273287006), .Z(n_15036));
	notech_nand2 i_317176(.A(n_274787021), .B(n_274187015), .Z(n_15031));
	notech_and4 i_217175(.A(n_275887032), .B(n_275787031), .C(n_275687030), 
		.D(n_276287036), .Z(n_15026));
	notech_and4 i_117174(.A(n_276687040), .B(n_276587039), .C(n_277587049), 
		.D(n_276987043), .Z(n_15021));
	notech_or2 i_22961499(.A(n_150628783), .B(n_29681), .Z(n_199159073));
	notech_nand2 i_3216245(.A(n_293387207), .B(n_292787201), .Z(n_19292));
	notech_nand2 i_3116244(.A(n_294487218), .B(n_293987213), .Z(n_19286));
	notech_nand2 i_3016243(.A(n_295587229), .B(n_295087224), .Z(n_19280));
	notech_nand2 i_2916242(.A(n_296687240), .B(n_296187235), .Z(n_19274));
	notech_nand2 i_2816241(.A(n_297787251), .B(n_297287246), .Z(n_19268));
	notech_nand2 i_2716240(.A(n_298887262), .B(n_298387257), .Z(n_19262));
	notech_nand2 i_2516238(.A(n_299987273), .B(n_299487268), .Z(n_19250));
	notech_nand2 i_2416237(.A(n_301087284), .B(n_300587279), .Z(n_19244));
	notech_nand2 i_2316236(.A(n_302187295), .B(n_301687290), .Z(n_19238));
	notech_nand2 i_1716230(.A(n_303287306), .B(n_302787301), .Z(n_19202));
	notech_nand2 i_717180(.A(n_304487318), .B(n_303887312), .Z(n_15051));
	notech_nand2 i_617179(.A(n_305687330), .B(n_305087324), .Z(n_15046));
	notech_nao3 i_50210(.A(n_310287376), .B(n_306487338), .C(n_310387377), .Z
		(\nbus_11326[0] ));
	notech_nand3 i_53952(.A(n_310187375), .B(n_58219), .C(n_310087374), .Z(n_21998
		));
	notech_nand3 i_8397(.A(n_308287356), .B(n_306087334), .C(n_308387357), .Z
		(n_22001));
	notech_nand2 i_817181(.A(n_312387397), .B(n_311787391), .Z(n_15056));
	notech_and4 i_526954(.A(n_315787431), .B(n_311187385), .C(n_312687400), 
		.D(n_307184062), .Z(n_19671));
	notech_nand2 i_1218977(.A(n_313887412), .B(n_313387407), .Z(n_25554));
	notech_nao3 i_23261496(.A(opc[21]), .B(n_62792), .C(n_307891745), .Z(n_198859070
		));
	notech_nao3 i_54455(.A(n_104085317), .B(n_315987433), .C(n_315887432), .Z
		(\nbus_11363[0] ));
	notech_and4 i_326952(.A(n_324463483), .B(n_317087444), .C(n_317587449), 
		.D(n_17539965), .Z(n_19659));
	notech_or2 i_17261556(.A(n_57984), .B(n_57644), .Z(n_194659033));
	notech_and4 i_118960602(.A(n_211359194), .B(n_56843), .C(n_3853), .D(n_54934
		), .Z(n_192159008));
	notech_ao4 i_166362839(.A(n_59460), .B(n_27084), .C(n_125461537), .D(n_58033
		), .Z(n_191859005));
	notech_and4 i_166962833(.A(n_191559002), .B(n_191359000), .C(n_185258948
		), .D(n_185358949), .Z(n_191759004));
	notech_ao4 i_166462838(.A(n_61103), .B(n_3835), .C(n_26060), .D(n_74438764
		), .Z(n_191559002));
	notech_ao4 i_166762835(.A(n_74738767), .B(n_32614), .C(n_74838768), .D(n_26892
		), .Z(n_191359000));
	notech_ao4 i_167062832(.A(n_26885), .B(n_66438684), .C(n_75738777), .D(n_65638676
		), .Z(n_191058997));
	notech_and4 i_167462828(.A(n_185958955), .B(n_183458930), .C(n_186158957
		), .D(n_27101), .Z(n_190958996));
	notech_ao4 i_169362809(.A(n_26956), .B(n_26891), .C(n_26959), .D(n_26889
		), .Z(n_189858988));
	notech_ao3 i_169662806(.A(n_186558961), .B(n_186658962), .C(n_186458960)
		, .Z(n_189758987));
	notech_and4 i_170362799(.A(n_186958964), .B(n_186758963), .C(n_187258965
		), .D(n_188758979), .Z(n_189358984));
	notech_and4 i_170262800(.A(n_187458967), .B(n_187358966), .C(n_187658969
		), .D(n_187558968), .Z(n_188758979));
	notech_nand2 i_8164372(.A(n_29640), .B(instrc[89]), .Z(n_65638676));
	notech_or4 i_11764337(.A(n_59326), .B(n_26900), .C(instrc[95]), .D(n_26972
		), .Z(n_65738677));
	notech_nao3 i_11964335(.A(n_3830), .B(instrc[124]), .C(instrc[127]), .Z(n_66438684
		));
	notech_nand2 i_11464339(.A(n_58122), .B(n_60915), .Z(n_74738767));
	notech_nao3 i_11564338(.A(instrc[105]), .B(n_30300), .C(n_57369), .Z(n_74838768
		));
	notech_or4 i_12064334(.A(n_6368850), .B(instrc[90]), .C(n_29642), .D(n_314663413
		), .Z(n_75738777));
	notech_and2 i_4764406(.A(n_29666), .B(instrc[93]), .Z(n_76238782));
	notech_and2 i_164364450(.A(instrc[125]), .B(n_29664), .Z(n_76638786));
	notech_nand3 i_10964344(.A(n_77638796), .B(n_29667), .C(n_26760), .Z(n_77438794
		));
	notech_and4 i_45964453(.A(n_56888), .B(n_3751), .C(instrc[97]), .D(n_26841
		), .Z(n_77638796));
	notech_and2 i_3164422(.A(n_3588), .B(n_3589), .Z(n_30905));
	notech_or4 i_96363514(.A(n_65638676), .B(instrc[88]), .C(n_314663413), .D
		(n_30306), .Z(n_187658969));
	notech_or4 i_96263515(.A(n_57011), .B(n_57042), .C(n_57064), .D(n_26971)
		, .Z(n_187558968));
	notech_nao3 i_96563512(.A(n_30332), .B(n_77638796), .C(n_26887), .Z(n_187458967
		));
	notech_or4 i_96463513(.A(instrc[103]), .B(n_29635), .C(n_29665), .D(n_26899
		), .Z(n_187358966));
	notech_nao3 i_96863509(.A(n_30946), .B(n_2026), .C(n_3824), .Z(n_187258965
		));
	notech_nao3 i_96763510(.A(n_30300), .B(n_30933), .C(n_26888), .Z(n_186958964
		));
	notech_or4 i_96663511(.A(instrc[123]), .B(instrc[120]), .C(n_3832), .D(n_29179
		), .Z(n_186758963));
	notech_or4 i_97163506(.A(instrc[115]), .B(n_59387), .C(n_246791942), .D(n_3829
		), .Z(n_186658962));
	notech_nao3 i_97063507(.A(n_60117), .B(n_60331), .C(n_304091783), .Z(n_186558961
		));
	notech_ao4 i_96963508(.A(n_26883), .B(n_26836), .C(n_184458940), .D(n_27344
		), .Z(n_186458960));
	notech_or4 i_92963548(.A(n_57042), .B(n_345480955), .C(n_57011), .D(n_57051
		), .Z(n_186158957));
	notech_and4 i_92863549(.A(n_62868), .B(n_76638786), .C(n_183358929), .D(n_28122
		), .Z(n_186058956));
	notech_or4 i_93063547(.A(instrc[103]), .B(n_29635), .C(instrc[102]), .D(n_26970
		), .Z(n_185958955));
	notech_nao3 i_93463543(.A(n_29666), .B(instrc[93]), .C(n_65738677), .Z(n_185858954
		));
	notech_nao3 i_93763540(.A(n_29639), .B(instrc[96]), .C(n_77438794), .Z(n_185358949
		));
	notech_nao3 i_94163536(.A(n_319091633), .B(n_26836), .C(n_59355), .Z(n_185258948
		));
	notech_nao3 i_88763589(.A(n_60117), .B(n_60319), .C(n_183158927), .Z(n_184858944
		));
	notech_or4 i_88663590(.A(n_27925), .B(n_32643), .C(n_125461537), .D(nZF)
		, .Z(n_184758943));
	notech_nand2 i_108463397(.A(n_26840), .B(n_62792), .Z(n_184658942));
	notech_and4 i_97663501(.A(n_62868), .B(n_28120), .C(n_30930), .D(n_27102
		), .Z(n_184458940));
	notech_nand2 i_6564388(.A(n_3828), .B(n_30910), .Z(n_184158937));
	notech_and4 i_7264381(.A(n_3827), .B(n_3826), .C(n_27035), .D(n_30905), 
		.Z(n_183958935));
	notech_and2 i_2364430(.A(n_59424), .B(n_3834), .Z(n_183858934));
	notech_ao4 i_14564309(.A(n_3824), .B(n_26767), .C(n_3829), .D(n_26060), 
		.Z(n_183458930));
	notech_ao4 i_10664347(.A(n_59441), .B(n_27029), .C(n_184158937), .D(n_27103
		), .Z(n_183358929));
	notech_or4 i_88863588(.A(n_25617), .B(n_27925), .C(n_60863), .D(nZF), .Z
		(n_183258928));
	notech_and4 i_14864306(.A(n_32656), .B(n_1869), .C(n_2941), .D(n_183258928
		), .Z(n_183158927));
	notech_ao4 i_10264351(.A(n_26840), .B(n_26837), .C(n_60969), .D(n_60958)
		, .Z(n_183058926));
	notech_and4 i_20067206(.A(n_177058866), .B(n_182558921), .C(n_177158867)
		, .D(n_177258868), .Z(n_182858924));
	notech_and4 i_19367209(.A(n_176758863), .B(n_312991694), .C(n_176958865)
		, .D(n_176858864), .Z(n_182558921));
	notech_or4 i_13967263(.A(temp_sp[0]), .B(temp_sp[1]), .C(n_181658912), .D
		(n_181358909), .Z(n_181858914));
	notech_nao3 i_12767275(.A(n_319391630), .B(n_27487), .C(temp_sp[30]), .Z
		(n_181658912));
	notech_or4 i_13467268(.A(temp_sp[3]), .B(temp_sp[4]), .C(temp_sp[5]), .D
		(temp_sp[2]), .Z(n_181358909));
	notech_or4 i_13367269(.A(temp_sp[6]), .B(temp_sp[7]), .C(temp_sp[8]), .D
		(temp_sp[9]), .Z(n_180958905));
	notech_or4 i_13267270(.A(temp_sp[10]), .B(temp_sp[11]), .C(temp_sp[12]),
		 .D(temp_sp[13]), .Z(n_180658902));
	notech_or4 i_14067262(.A(n_180158897), .B(n_179858894), .C(n_179458890),
		 .D(n_179158887), .Z(n_180358899));
	notech_or4 i_13167271(.A(temp_sp[14]), .B(temp_sp[16]), .C(temp_sp[17]),
		 .D(temp_sp[15]), .Z(n_180158897));
	notech_or4 i_13067272(.A(temp_sp[18]), .B(temp_sp[19]), .C(temp_sp[20]),
		 .D(temp_sp[21]), .Z(n_179858894));
	notech_or4 i_12967273(.A(temp_sp[22]), .B(temp_sp[23]), .C(temp_sp[24]),
		 .D(temp_sp[25]), .Z(n_179458890));
	notech_or4 i_12867274(.A(temp_sp[26]), .B(temp_sp[27]), .C(temp_sp[28]),
		 .D(temp_sp[29]), .Z(n_179158887));
	notech_ao4 i_14867254(.A(n_26611), .B(n_3846), .C(n_54930), .D(n_60935),
		 .Z(n_178658882));
	notech_nao3 i_17867224(.A(n_19029), .B(n_19014), .C(n_19022), .Z(n_178158877
		));
	notech_and2 i_17267230(.A(n_175858854), .B(n_175758853), .Z(n_178058876)
		);
	notech_nand2 i_17767225(.A(n_18981), .B(n_26780), .Z(n_177658872));
	notech_nor2 i_267393(.A(n_32403), .B(n_3807), .Z(n_177558871));
	notech_ao3 i_53401(.A(n_177358869), .B(n_182858924), .C(n_176458860), .Z
		(n_177458870));
	notech_or4 i_18367219(.A(tcmp), .B(n_174958845), .C(n_61130), .D(n_176358859
		), .Z(n_177358869));
	notech_nao3 i_18267220(.A(n_177558871), .B(n_176258858), .C(n_19029), .Z
		(n_177258868));
	notech_nand3 i_18567217(.A(n_60117), .B(n_60319), .C(n_176658862), .Z(n_177158867
		));
	notech_or4 i_18767215(.A(tcmp), .B(n_56614), .C(n_56829), .D(n_61130), .Z
		(n_177058866));
	notech_or4 i_18667216(.A(instrc[127]), .B(n_26968), .C(n_26838), .D(instrc
		[124]), .Z(n_176958865));
	notech_nand2 i_18167221(.A(fesp), .B(n_61130), .Z(n_176858864));
	notech_or4 i_18067222(.A(n_19057), .B(n_32579), .C(n_317791646), .D(n_60331
		), .Z(n_176758863));
	notech_nand3 i_5967342(.A(n_32434), .B(n_176158857), .C(n_32432), .Z(n_176658862
		));
	notech_ao4 i_6067341(.A(n_178058876), .B(n_178158877), .C(n_177658872), 
		.D(n_29655), .Z(n_176558861));
	notech_nor2 i_18467218(.A(n_176558861), .B(n_27108), .Z(n_176458860));
	notech_ao3 i_6167340(.A(n_178658882), .B(n_175658852), .C(n_175358849), 
		.Z(n_176358859));
	notech_or4 i_6267339(.A(n_180958905), .B(n_180658902), .C(n_181858914), 
		.D(n_180358899), .Z(n_176258858));
	notech_or2 i_17967223(.A(n_30312), .B(n_56391), .Z(n_176158857));
	notech_or4 i_15667246(.A(instrc[123]), .B(instrc[120]), .C(n_60915), .D(n_27045
		), .Z(n_175858854));
	notech_or4 i_15167251(.A(n_30344), .B(n_57082), .C(n_57064), .D(n_54916)
		, .Z(n_175758853));
	notech_nao3 i_14567257(.A(n_32334), .B(n_26626), .C(n_2351), .Z(n_175658852
		));
	notech_ao4 i_3567366(.A(n_59441), .B(n_27110), .C(n_56939), .D(n_32380),
		 .Z(n_175458850));
	notech_and4 i_14667256(.A(n_62868), .B(n_30930), .C(n_175458850), .D(n_30931
		), .Z(n_175358849));
	notech_ao4 i_067394(.A(n_2480), .B(n_62892), .C(n_56829), .D(n_32286), .Z
		(n_174958845));
	notech_or4 i_99(.A(n_62844), .B(n_27904), .C(n_60935), .D(n_60223), .Z(n_27879
		));
	notech_nand2 i_1979(.A(n_27132), .B(n_27123), .Z(n_32655));
	notech_or2 i_1743(.A(n_293591841), .B(n_27056), .Z(n_23040));
	notech_nand2 i_1624(.A(n_27123), .B(n_62892), .Z(n_32462));
	notech_nao3 i_1616(.A(n_62870), .B(n_32730), .C(n_58086), .Z(n_25349));
	notech_ao4 i_1571(.A(n_60863), .B(n_25615), .C(n_25629), .D(n_59413), .Z
		(n_25386));
	notech_nao3 i_1520(.A(n_32747), .B(n_62892), .C(n_58086), .Z(n_25619));
	notech_ao4 i_1458(.A(n_60863), .B(n_25349), .C(n_60888), .D(n_25615), .Z
		(n_23007));
	notech_nao3 i_1301(.A(n_60874), .B(n_32730), .C(n_27925), .Z(n_27924));
	notech_or4 i_1262(.A(n_26638), .B(n_26782), .C(n_60223), .D(n_26962), .Z
		(n_27782));
	notech_or4 i_1261(.A(n_26638), .B(n_26782), .C(n_60223), .D(n_32384), .Z
		(n_22309));
	notech_nao3 i_1248(.A(n_60874), .B(n_62892), .C(n_27501), .Z(n_27500));
	notech_and2 i_1202(.A(n_2676), .B(n_23627), .Z(n_23625));
	notech_nand2 i_1171(.A(n_2825), .B(n_27132), .Z(n_32443));
	notech_nor2 i_1141(.A(n_61161), .B(n_27719), .Z(n_32605));
	notech_or4 i_1029(.A(n_60863), .B(n_59451), .C(n_60223), .D(n_26782), .Z
		(n_22582));
	notech_or4 i_1028(.A(n_60863), .B(n_59451), .C(n_60223), .D(n_27896), .Z
		(n_22579));
	notech_or4 i_796(.A(n_60274), .B(n_32443), .C(n_60874), .D(n_62892), .Z(n_25615
		));
	notech_or4 i_794(.A(n_2825), .B(n_60274), .C(n_59478), .D(n_27132), .Z(n_27917
		));
	notech_nao3 i_789(.A(n_27170), .B(n_32695), .C(n_32443), .Z(n_32259));
	notech_or4 i_782(.A(n_2825), .B(n_2838), .C(n_32695), .D(n_2864), .Z(n_27501
		));
	notech_nand2 i_752(.A(n_60874), .B(n_62892), .Z(n_32643));
	notech_nao3 i_742(.A(n_27170), .B(n_32695), .C(n_2839), .Z(n_25625));
	notech_nao3 i_433(.A(n_57976), .B(n_58009), .C(n_57933), .Z(n_23029));
	notech_or4 i_432(.A(instrc[123]), .B(instrc[120]), .C(n_32342), .D(n_57933
		), .Z(n_23031));
	notech_or4 i_430(.A(n_60223), .B(n_60841), .C(n_59424), .D(n_58033), .Z(n_23019
		));
	notech_ao3 i_386(.A(n_59441), .B(n_27896), .C(n_59451), .Z(n_27784));
	notech_ao4 i_322(.A(n_60863), .B(n_27924), .C(n_59424), .D(n_27095), .Z(n_23627
		));
	notech_or4 i_37224(.A(n_61171), .B(n_61161), .C(n_61149), .D(n_1892), .Z
		(n_22313));
	notech_nao3 i_891(.A(n_26962), .B(n_57967), .C(n_27879), .Z(n_22322));
	notech_or4 i_37002(.A(n_25619), .B(n_62850), .C(n_62792), .D(n_60223), .Z
		(n_22571));
	notech_or4 i_37001(.A(n_60863), .B(n_59460), .C(n_60223), .D(n_26782), .Z
		(n_22572));
	notech_or4 i_36990(.A(n_60863), .B(n_59460), .C(n_60218), .D(n_57967), .Z
		(n_22585));
	notech_or4 i_36986(.A(calc_sz[3]), .B(n_58062), .C(n_27879), .D(calc_sz[
		2]), .Z(n_22590));
	notech_or4 i_36985(.A(n_59413), .B(n_27904), .C(n_60218), .D(n_57967), .Z
		(n_22591));
	notech_or4 i_36983(.A(n_27907), .B(n_59429), .C(n_60218), .D(n_57967), .Z
		(n_22594));
	notech_nao3 i_2873(.A(n_62820), .B(n_62850), .C(n_2884), .Z(n_22995));
	notech_or4 i_36638(.A(n_61171), .B(n_61161), .C(n_61149), .D(n_2530), .Z
		(n_23003));
	notech_or4 i_36633(.A(n_59451), .B(n_62850), .C(n_62792), .D(n_60218), .Z
		(n_23009));
	notech_or4 i_36621(.A(instrc[122]), .B(n_32614), .C(n_57933), .D(n_60915
		), .Z(n_23023));
	notech_or4 i_36610(.A(n_60274), .B(n_59478), .C(n_32443), .D(n_32323), .Z
		(n_23036));
	notech_or4 i_36603(.A(n_319691627), .B(n_62792), .C(n_60899), .D(n_60218
		), .Z(n_23045));
	notech_or4 i_1206(.A(n_32729), .B(n_58086), .C(n_59413), .D(n_60218), .Z
		(n_23049));
	notech_or4 i_1014(.A(n_25619), .B(n_60935), .C(n_60899), .D(n_60218), .Z
		(n_23052));
	notech_or4 i_413(.A(n_315291671), .B(n_62850), .C(n_60933), .D(n_60218),
		 .Z(n_23059));
	notech_nao3 i_35811(.A(n_60378), .B(n_2947), .C(n_27037), .Z(n_23940));
	notech_or4 i_35804(.A(n_61171), .B(n_61161), .C(n_27037), .D(n_2947), .Z
		(n_23947));
	notech_ao3 i_792(.A(n_2825), .B(n_27132), .C(n_2883), .Z(n_25374));
	notech_ao4 i_1457(.A(n_59413), .B(n_25615), .C(n_25629), .D(n_60888), .Z
		(n_25385));
	notech_nao3 i_800(.A(n_2825), .B(n_27132), .C(n_2888), .Z(n_25629));
	notech_nao3 i_32466(.A(n_60874), .B(n_32730), .C(n_32259), .Z(n_27509)
		);
	notech_or4 i_32194(.A(n_61171), .B(n_61161), .C(n_61149), .D(n_58072), .Z
		(n_27781));
	notech_or2 i_32125(.A(n_27917), .B(n_26782), .Z(n_27850));
	notech_or2 i_1282(.A(n_59460), .B(n_57967), .Z(n_27857));
	notech_and2 i_210006(.A(rep_en2), .B(n_1886), .Z(n_27877));
	notech_and2 i_18656(.A(n_26962), .B(n_57967), .Z(n_27880));
	notech_ao3 i_3091(.A(n_60899), .B(n_62792), .C(n_27904), .Z(n_27903));
	notech_ao3 i_2994(.A(n_60899), .B(n_60931), .C(n_59451), .Z(n_27906));
	notech_ao3 i_32053(.A(n_62868), .B(n_32730), .C(n_27925), .Z(n_27922));
	notech_nand2 i_904(.A(n_57909), .B(nbus_11295[2]), .Z(n_27959));
	notech_nao3 i_31899(.A(n_60378), .B(n_1891), .C(n_61149), .Z(n_28076));
	notech_and2 i_828(.A(n_60863), .B(n_60888), .Z(n_1864));
	notech_or4 i_31896(.A(n_28081), .B(n_2877), .C(n_27123), .D(n_27170), .Z
		(n_28079));
	notech_ao4 i_1195(.A(n_59413), .B(n_2893), .C(n_2868), .D(n_59429), .Z(n_30987
		));
	notech_and3 i_972(.A(n_26702), .B(n_26643), .C(n_59708), .Z(n_32458));
	notech_ao4 i_900(.A(n_59413), .B(n_2868), .C(n_2873), .D(n_2872), .Z(n_32459
		));
	notech_and2 i_27323(.A(n_32656), .B(n_1869), .Z(n_32652));
	notech_or4 i_2827(.A(n_60969), .B(n_60958), .C(n_2884), .D(n_62850), .Z(n_32656
		));
	notech_and3 i_1938(.A(vliw_pc[0]), .B(vliw_pc[1]), .C(vliw_pc[2]), .Z(n_32834
		));
	notech_and2 i_1913(.A(vliw_pc[0]), .B(vliw_pc[1]), .Z(n_32843));
	notech_and2 i_901(.A(n_32729), .B(n_28081), .Z(n_1868));
	notech_or4 i_3505(.A(n_2825), .B(n_2838), .C(n_32695), .D(n_27170), .Z(n_1869
		));
	notech_or4 i_3126(.A(n_58086), .B(n_28081), .C(n_62850), .D(n_60931), .Z
		(n_1870));
	notech_or4 i_3113(.A(n_58086), .B(n_28081), .C(n_62792), .D(n_60899), .Z
		(n_1871));
	notech_or4 i_5970(.A(n_2839), .B(n_2883), .C(n_60931), .D(n_60904), .Z(n_1872
		));
	notech_nand2 i_5(.A(n_2659), .B(n_27352), .Z(n_18559));
	notech_and3 i_2350(.A(reps[2]), .B(n_2666), .C(n_2663), .Z(n_1874));
	notech_ao4 i_359(.A(n_293591841), .B(n_57899), .C(n_2895), .D(n_60218), 
		.Z(n_18756873));
	notech_ao4 i_361(.A(n_27052), .B(n_293491842), .C(n_32656), .D(n_60218),
		 .Z(n_1876));
	notech_mux2 i_363(.S(n_60331), .A(n_19072), .B(n_22995), .Z(n_1877));
	notech_ao4 i_1196(.A(n_2896), .B(n_3790), .C(n_27145), .D(n_27037), .Z(n_1878
		));
	notech_and3 i_316(.A(n_30987), .B(n_32446), .C(n_2658), .Z(n_1880));
	notech_or4 i_2835(.A(n_60274), .B(n_28081), .C(n_2839), .D(n_60863), .Z(n_1881
		));
	notech_or4 i_1309(.A(n_61171), .B(n_61161), .C(n_61149), .D(n_2653), .Z(n_1884
		));
	notech_nand3 i_1710(.A(n_57909), .B(nbus_11295[2]), .C(nbus_11295[4]), .Z
		(n_1886));
	notech_or4 i_248(.A(n_61171), .B(n_61161), .C(n_61149), .D(n_1893), .Z(n_1887
		));
	notech_or4 i_1557(.A(n_61171), .B(n_61160), .C(n_61149), .D(n_2895), .Z(n_1889
		));
	notech_nao3 i_3579(.A(n_62820), .B(n_62850), .C(n_2893), .Z(n_18906874)
		);
	notech_nand3 i_1280(.A(n_1899), .B(n_1900), .C(n_28079), .Z(n_1891));
	notech_and2 i_389(.A(n_1906), .B(n_1907), .Z(n_1892));
	notech_and2 i_1198(.A(n_1894), .B(n_1895), .Z(n_1893));
	notech_nao3 i_3323(.A(n_62844), .B(n_62790), .C(n_27509), .Z(n_1894));
	notech_or4 i_2845(.A(n_60969), .B(n_60958), .C(n_2884), .D(n_60899), .Z(n_1897
		));
	notech_nao3 i_2934(.A(n_62820), .B(n_62850), .C(n_59460), .Z(n_1898));
	notech_or4 i_3035(.A(n_32729), .B(n_60274), .C(n_2877), .D(n_59429), .Z(n_1899
		));
	notech_or4 i_3052(.A(n_32729), .B(n_60274), .C(n_59413), .D(n_2877), .Z(n_1900
		));
	notech_or4 i_3099(.A(n_58086), .B(n_28081), .C(n_62850), .D(n_62816), .Z
		(n_1906));
	notech_or4 i_3106(.A(n_60969), .B(n_60958), .C(n_25349), .D(n_62834), .Z
		(n_1907));
	notech_and4 i_127960(.A(n_2789), .B(n_2798), .C(n_2575), .D(n_2562), .Z(n_32747
		));
	notech_and4 i_827967(.A(n_2840), .B(n_2849), .C(n_2603), .D(n_2590), .Z(n_32695
		));
	notech_and3 i_1592(.A(n_2676), .B(n_23627), .C(n_2685), .Z(n_22035));
	notech_and4 i_329(.A(n_32656), .B(n_1869), .C(n_2939), .D(n_1872), .Z(n_22024
		));
	notech_and3 i_37503(.A(n_2529), .B(n_59167), .C(n_2531), .Z(n_22015));
	notech_nand3 i_50490(.A(n_2881), .B(fsm[3]), .C(n_32605), .Z(n_19065));
	notech_ao3 i_1304(.A(n_2838), .B(n_27170), .C(n_2825), .Z(n_32470));
	notech_ao4 i_1035(.A(n_60863), .B(n_2884), .C(n_60893), .D(n_59460), .Z(n_25651
		));
	notech_nor2 i_1330436(.A(n_330963526), .B(n_2946), .Z(n_1862));
	notech_or4 i_23932535(.A(n_2366), .B(n_32579), .C(n_19057), .D(n_60331),
		 .Z(n_320491619));
	notech_and3 i_22332547(.A(n_18998), .B(n_18989), .C(n_32551), .Z(n_320391620
		));
	notech_nand2 i_16232580(.A(n_18998), .B(n_18989), .Z(n_320291621));
	notech_or4 i_50497(.A(fsm[0]), .B(fsm[3]), .C(n_27145), .D(n_27717), .Z(n_19029
		));
	notech_and3 i_50494(.A(n_61160), .B(n_61171), .C(n_272491901), .Z(n_19043
		));
	notech_nao3 i_762(.A(n_27123), .B(n_2864), .C(n_32443), .Z(n_27925));
	notech_or4 i_795(.A(n_32643), .B(n_60274), .C(n_2825), .D(n_27132), .Z(n_27907
		));
	notech_and4 i_8532654(.A(n_60899), .B(n_60931), .C(n_60138), .D(n_60331)
		, .Z(n_32272));
	notech_and2 i_119332703(.A(n_27854), .B(n_27856), .Z(n_320191622));
	notech_and4 i_126950(.A(n_320491619), .B(n_2526), .C(n_2525), .D(n_26860
		), .Z(n_320091623));
	notech_and4 i_830221(.A(n_57020), .B(n_57011), .C(n_57051), .D(n_57033),
		 .Z(n_17107));
	notech_and2 i_27932741(.A(n_26755), .B(n_59335), .Z(n_319991624));
	notech_or4 i_21132559(.A(instrc[122]), .B(n_32343), .C(n_60915), .D(n_317591648
		), .Z(n_23507));
	notech_ao4 i_105932745(.A(n_317591648), .B(n_32323), .C(n_59418), .D(n_23510
		), .Z(n_319891625));
	notech_ao3 i_19232746(.A(n_57011), .B(n_57055), .C(n_55581), .Z(n_23510)
		);
	notech_ao4 i_48832748(.A(n_56854), .B(n_26962), .C(n_32352), .D(n_32408)
		, .Z(n_23513));
	notech_ao4 i_49232749(.A(n_56854), .B(n_56979), .C(n_56675), .D(n_32408)
		, .Z(n_23514));
	notech_nand2 i_129732751(.A(n_60207), .B(n_19057), .Z(n_23755));
	notech_or4 i_35948(.A(n_3804), .B(n_60283), .C(n_19079), .D(n_29655), .Z
		(n_319791626));
	notech_or4 i_80632753(.A(n_59478), .B(n_2877), .C(n_27123), .D(n_27170),
		 .Z(n_319691627));
	notech_or4 i_3499(.A(n_32729), .B(n_62816), .C(n_60899), .D(n_27573), .Z
		(n_319591628));
	notech_nand2 i_725(.A(n_62868), .B(n_32730), .Z(n_32729));
	notech_or4 i_3495(.A(n_60969), .B(n_60958), .C(n_27904), .D(n_60899), .Z
		(n_319491629));
	notech_mux2 i_2137(.S(n_2488), .A(n_2376), .B(n_3848598), .Z(n_319391630
		));
	notech_nand2 i_27420(.A(n_19029), .B(n_26963), .Z(n_32555));
	notech_ao4 i_59932756(.A(n_2351), .B(n_32334), .C(n_59418), .D(n_17107),
		 .Z(n_319291631));
	notech_or2 i_21332557(.A(n_2351), .B(n_56391), .Z(n_26611));
	notech_ao4 i_74632758(.A(n_32351), .B(n_32286), .C(n_56843), .D(n_61131)
		, .Z(n_26613));
	notech_ao4 i_74432759(.A(n_32355), .B(n_32286), .C(n_61131), .D(n_27024)
		, .Z(n_26614));
	notech_or4 i_13432607(.A(n_60274), .B(n_2839), .C(n_62870), .D(n_60986),
		 .Z(n_27988));
	notech_and2 i_197432692(.A(n_57011), .B(n_57055), .Z(n_30945));
	notech_and2 i_29029(.A(n_57020), .B(n_57033), .Z(n_30946));
	notech_or4 i_125632779(.A(n_62844), .B(n_60931), .C(n_61131), .D(n_60207
		), .Z(n_32263));
	notech_and2 i_18018(.A(n_59387), .B(instrc[115]), .Z(n_319191632));
	notech_and2 i_132791(.A(n_59402), .B(n_29177), .Z(n_319091633));
	notech_nand3 i_23532538(.A(n_246591944), .B(n_57055), .C(n_62816), .Z(n_32309
		));
	notech_nor2 i_830276(.A(n_58062), .B(n_2937), .Z(n_32384));
	notech_nao3 i_16032582(.A(n_60915), .B(n_27194), .C(n_101413114), .Z(n_32361
		));
	notech_ao4 i_38832805(.A(n_317391650), .B(n_32365), .C(n_32393), .D(n_59418
		), .Z(n_318991634));
	notech_nao3 i_72332806(.A(n_32380), .B(n_60138), .C(n_56829), .Z(n_32370
		));
	notech_nao3 i_22432546(.A(n_60319), .B(n_62892), .C(n_32378), .Z(n_32372
		));
	notech_nor2 i_194532694(.A(n_59387), .B(n_29178), .Z(n_318891635));
	notech_nao3 i_197132809(.A(n_60319), .B(n_60986), .C(n_32378), .Z(n_32376
		));
	notech_and4 i_15732813(.A(n_57020), .B(n_57042), .C(n_57082), .D(n_57055
		), .Z(n_32393));
	notech_or4 i_12532616(.A(n_32581), .B(n_32559), .C(n_26900), .D(n_61131)
		, .Z(n_32403));
	notech_or4 i_14132600(.A(n_32569), .B(n_3804), .C(n_19050), .D(n_26963),
		 .Z(n_32405));
	notech_nor2 i_032814(.A(n_59402), .B(n_59393), .Z(n_318791636));
	notech_ao4 i_851(.A(n_59429), .B(n_2870), .C(n_60863), .D(n_2868), .Z(n_32446
		));
	notech_nand2 i_123232817(.A(n_32446), .B(n_27085), .Z(n_7148928));
	notech_or4 i_16330(.A(n_59387), .B(n_246791942), .C(n_32351), .D(n_59364
		), .Z(n_318691637));
	notech_and4 i_427963(.A(n_2801), .B(n_2810), .C(n_2589), .D(n_2576), .Z(n_32730
		));
	notech_or4 i_3327(.A(n_32259), .B(n_60893), .C(n_60874), .D(\opcode[3] )
		, .Z(n_1895));
	notech_or4 i_5990(.A(n_32403), .B(n_19043), .C(n_26756), .D(n_32566), .Z
		(n_318591638));
	notech_or4 i_32332867(.A(n_27988), .B(n_62836), .C(n_62816), .D(n_60207)
		, .Z(n_318491639));
	notech_or4 i_25632868(.A(n_61171), .B(n_61160), .C(n_61149), .D(n_23006)
		, .Z(n_318391640));
	notech_or4 i_25732869(.A(n_61171), .B(n_61160), .C(n_61149), .D(n_2368),
		 .Z(n_318291641));
	notech_or4 i_16322(.A(n_101413114), .B(n_29179), .C(n_317391650), .D(n_32350
		), .Z(n_318191642));
	notech_nao3 i_16334(.A(n_60138), .B(n_60319), .C(n_32257), .Z(n_318091643
		));
	notech_or4 i_67232823(.A(n_59387), .B(n_246791942), .C(n_32355), .D(n_59364
		), .Z(n_317991644));
	notech_or4 i_7522(.A(n_59393), .B(n_59402), .C(n_304291781), .D(n_27577)
		, .Z(n_317891645));
	notech_or2 i_34332899(.A(n_32405), .B(n_3848598), .Z(n_317791646));
	notech_nand2 i_185832904(.A(n_27177), .B(n_60845), .Z(n_317691647));
	notech_ao4 i_83632906(.A(n_62820), .B(n_60899), .C(n_60888), .D(n_23510)
		, .Z(n_317591648));
	notech_ao4 i_98932908(.A(n_62798), .B(n_60899), .C(n_60888), .D(n_32393)
		, .Z(n_317391650));
	notech_ao3 i_183832909(.A(n_60931), .B(n_62836), .C(n_2893), .Z(n_317291651
		));
	notech_or2 i_167332916(.A(n_2351), .B(n_32334), .Z(n_317191652));
	notech_ao4 i_48332799(.A(n_32355), .B(n_32373), .C(n_61131), .D(n_27024)
		, .Z(n_317091653));
	notech_or4 i_154732922(.A(n_101413114), .B(n_317091653), .C(n_29179), .D
		(n_317391650), .Z(n_316991654));
	notech_ao4 i_48532871(.A(n_32347), .B(n_32373), .C(n_305391770), .D(n_61131
		), .Z(n_316891655));
	notech_or4 i_154432923(.A(n_101413114), .B(n_29179), .C(n_317391650), .D
		(n_316891655), .Z(n_316791656));
	notech_ao4 i_49432747(.A(n_56854), .B(n_56959), .C(n_56813), .D(n_32408)
		, .Z(n_23512));
	notech_or4 i_137832924(.A(n_60854), .B(n_32343), .C(n_317591648), .D(n_23512
		), .Z(n_316691657));
	notech_ao4 i_48632925(.A(n_32370), .B(n_32373), .C(n_305091773), .D(n_61131
		), .Z(n_316591658));
	notech_ao4 i_49032926(.A(n_56858), .B(n_56941), .C(n_56684), .D(n_32408)
		, .Z(n_316491659));
	notech_and3 i_86232927(.A(n_23513), .B(n_23514), .C(n_23512), .Z(n_316391660
		));
	notech_nand3 i_81332930(.A(n_2414), .B(n_27177), .C(n_32323), .Z(n_316291661
		));
	notech_and2 i_148032893(.A(n_59434), .B(n_319891625), .Z(n_316191662));
	notech_nand3 i_81532932(.A(n_32393), .B(n_2417), .C(n_62816), .Z(n_315991664
		));
	notech_and2 i_199332872(.A(n_59434), .B(n_318991634), .Z(n_315891665));
	notech_or4 i_66932934(.A(n_59393), .B(n_59402), .C(n_56675), .D(n_27577)
		, .Z(n_315691667));
	notech_or4 i_66632935(.A(n_59387), .B(n_246791942), .C(n_32347), .D(n_59364
		), .Z(n_315591668));
	notech_or4 i_23832937(.A(n_61171), .B(n_61160), .C(n_61149), .D(n_319591628
		), .Z(n_315491669));
	notech_or4 i_25832938(.A(n_61171), .B(n_61160), .C(n_61149), .D(n_319491629
		), .Z(n_315391670));
	notech_nand2 i_724(.A(n_60874), .B(n_60986), .Z(n_28081));
	notech_nao3 i_3463(.A(n_62844), .B(n_60931), .C(n_59469), .Z(n_23006));
	notech_or4 i_31981(.A(n_62870), .B(n_60986), .C(n_27123), .D(n_27170), .Z
		(n_27994));
	notech_or4 i_31982(.A(n_60274), .B(n_2877), .C(n_62870), .D(n_60986), .Z
		(n_315291671));
	notech_and3 i_32120(.A(n_60899), .B(n_62816), .C(n_60319), .Z(n_27855)
		);
	notech_or4 i_2860(.A(n_4958709), .B(n_27123), .C(n_27132), .D(n_60874), 
		.Z(n_32432));
	notech_or4 i_2853(.A(n_4958709), .B(n_27123), .C(n_27132), .D(n_62870), 
		.Z(n_32434));
	notech_nor2 i_930428(.A(n_60854), .B(n_32343), .Z(n_32323));
	notech_ao3 i_1338260(.A(n_60915), .B(n_32367), .C(n_60975), .Z(n_32319)
		);
	notech_ao3 i_1438261(.A(n_29179), .B(n_32367), .C(n_60975), .Z(n_32322)
		);
	notech_or2 i_1326(.A(n_60975), .B(n_60915), .Z(n_32326));
	notech_ao3 i_4338262(.A(instrc[120]), .B(instrc[123]), .C(n_60854), .Z(n_32325
		));
	notech_ao3 i_4538263(.A(instrc[120]), .B(instrc[123]), .C(n_32342), .Z(n_32331
		));
	notech_and3 i_4638264(.A(n_60975), .B(n_32367), .C(n_29179), .Z(n_32332)
		);
	notech_or2 i_27633(.A(n_60975), .B(n_29179), .Z(n_32342));
	notech_and4 i_5338266(.A(n_60975), .B(instrc[120]), .C(instrc[123]), .D(n_29179
		), .Z(n_32338));
	notech_ao3 i_5538267(.A(n_60975), .B(n_29179), .C(n_32614), .Z(n_32344)
		);
	notech_nand2 i_27361(.A(instrc[120]), .B(n_29180), .Z(n_32614));
	notech_or2 i_1230(.A(instrc[120]), .B(instrc[123]), .Z(n_32343));
	notech_ao3 i_21717(.A(n_60975), .B(n_29179), .C(n_32343), .Z(n_32334));
	notech_and3 i_4938304(.A(n_60975), .B(n_32367), .C(n_60915), .Z(n_32365)
		);
	notech_ao4 i_49341299(.A(n_56858), .B(n_56983), .C(n_56675), .D(n_32295)
		, .Z(n_24994));
	notech_nor2 i_930492(.A(n_32343), .B(n_32342), .Z(n_32341));
	notech_or4 i_129641300(.A(instrc[123]), .B(instrc[120]), .C(n_32342), .D
		(n_314891675), .Z(n_24996));
	notech_ao4 i_60141301(.A(n_57992), .B(n_314891675), .C(n_59418), .D(n_25007
		), .Z(n_315191672));
	notech_ao3 i_12441303(.A(n_29653), .B(n_2026), .C(n_57020), .Z(n_25007)
		);
	notech_or4 i_50641307(.A(n_61171), .B(n_61160), .C(n_61149), .D(n_30594)
		, .Z(n_30570));
	notech_or2 i_11290(.A(n_300891815), .B(n_313491689), .Z(n_315091673));
	notech_nand2 i_183741385(.A(n_57976), .B(n_27221), .Z(n_314991674));
	notech_ao4 i_83741386(.A(n_62820), .B(n_60899), .C(n_60888), .D(n_25007)
		, .Z(n_314891675));
	notech_and4 i_94238271(.A(n_2343), .B(n_2342), .C(n_2338), .D(n_2341), .Z
		(n_314791676));
	notech_ao4 i_5744437(.A(n_30822), .B(n_57837), .C(n_30821), .D(n_59726),
		 .Z(n_314691677));
	notech_ao4 i_3944455(.A(n_32370), .B(n_28016), .C(n_314091683), .D(n_314391680
		), .Z(n_314591678));
	notech_and4 i_3217045(.A(n_1990), .B(n_1992), .C(n_1998), .D(n_1923), .Z
		(n_314491679));
	notech_and4 i_145444498(.A(n_1983), .B(n_1982), .C(n_1976), .D(n_1981), 
		.Z(n_314391680));
	notech_ao4 i_49541368(.A(n_56858), .B(n_56959), .C(n_56813), .D(n_32295)
		, .Z(n_25010));
	notech_ao4 i_24304(.A(n_58062), .B(n_2937), .C(n_58101), .D(n_56970), .Z
		(n_314291681));
	notech_nand2 i_186041384(.A(n_26643), .B(n_26634), .Z(n_314191682));
	notech_nand2 i_200044520(.A(n_314191682), .B(n_26627), .Z(n_30470));
	notech_nand3 i_191441382(.A(n_314191682), .B(n_56983), .C(n_314291681), 
		.Z(n_30821));
	notech_or4 i_62244521(.A(n_60969), .B(n_60958), .C(n_62836), .D(n_29614)
		, .Z(n_31279));
	notech_and3 i_103744541(.A(n_32351), .B(n_32355), .C(n_32347), .Z(n_314091683
		));
	notech_ao4 i_132244542(.A(n_1903), .B(n_314191682), .C(n_26627), .D(n_32386
		), .Z(n_313991684));
	notech_or4 i_165544570(.A(n_57064), .B(n_57011), .C(n_54916), .D(n_27349
		), .Z(n_27348));
	notech_nand2 i_114644580(.A(n_27163), .B(n_27102), .Z(n_313891685));
	notech_nand2 i_90644583(.A(n_27163), .B(n_27344), .Z(n_313791686));
	notech_and2 i_88344584(.A(n_32351), .B(n_32355), .Z(n_313691687));
	notech_or2 i_50241389(.A(n_306291761), .B(n_56959), .Z(n_313591688));
	notech_and2 i_148144576(.A(n_59429), .B(n_299691827), .Z(n_313491689));
	notech_nand3 i_2147678(.A(n_32352), .B(n_56813), .C(n_32356), .Z(n_313391690
		));
	notech_nand2 i_32636(.A(n_312491699), .B(n_27344), .Z(n_313291691));
	notech_or4 i_68732755(.A(n_59387), .B(n_59275), .C(n_32347), .D(instrc[
		115]), .Z(n_313191692));
	notech_or4 i_10592(.A(n_59382), .B(n_59275), .C(instrc[115]), .D(n_313691687
		), .Z(n_313091693));
	notech_nao3 i_202332858(.A(n_60138), .B(n_60319), .C(n_1895), .Z(n_312991694
		));
	notech_or2 i_10589(.A(n_26616), .B(n_312091703), .Z(n_312891695));
	notech_or2 i_10588(.A(n_26616), .B(n_26611), .Z(n_312791696));
	notech_nao3 i_186647749(.A(n_32334), .B(n_303491789), .C(n_2351), .Z(n_312691697
		));
	notech_nand2 i_186547750(.A(n_303491789), .B(n_27109), .Z(n_312591698)
		);
	notech_nand2 i_170047756(.A(n_300891815), .B(n_27346), .Z(n_312491699)
		);
	notech_and2 i_147847763(.A(n_301891805), .B(n_300391820), .Z(n_104922313
		));
	notech_ao4 i_147647764(.A(n_59441), .B(n_27302), .C(n_28542), .D(n_26683
		), .Z(n_105022314));
	notech_or4 i_139041298(.A(n_32343), .B(n_32342), .C(n_314891675), .D(n_25010
		), .Z(n_312391700));
	notech_and2 i_158641367(.A(n_59429), .B(n_315191672), .Z(n_312291701));
	notech_ao4 i_75032757(.A(n_32370), .B(n_32286), .C(n_305091773), .D(n_61131
		), .Z(n_312191702));
	notech_and2 i_158832885(.A(n_59429), .B(n_319291631), .Z(n_312091703));
	notech_ao4 i_49141302(.A(n_56858), .B(n_56941), .C(n_56684), .D(n_32295)
		, .Z(n_311991704));
	notech_and4 i_264350693(.A(n_56843), .B(n_2004), .C(n_24994), .D(n_25010
		), .Z(n_311891705));
	notech_and2 i_198371097(.A(n_60899), .B(n_60931), .Z(n_32763));
	notech_or4 i_67141312(.A(n_59382), .B(n_56675), .C(instrc[115]), .D(n_27192
		), .Z(n_311791706));
	notech_or4 i_9177(.A(n_59382), .B(n_304291781), .C(instrc[115]), .D(n_27192
		), .Z(n_311691707));
	notech_ao4 i_48032874(.A(n_61103), .B(n_32257), .C(n_56592), .D(n_32370)
		, .Z(n_121628493));
	notech_ao4 i_85932878(.A(n_59441), .B(n_27196), .C(n_2417), .D(n_26818),
		 .Z(n_122228499));
	notech_and2 i_86032879(.A(n_315991664), .B(n_2372), .Z(n_122428501));
	notech_and3 i_86132880(.A(n_318191642), .B(n_316991654), .C(n_316791656)
		, .Z(n_122528502));
	notech_and3 i_50532875(.A(n_2508), .B(n_26648), .C(n_243491968), .Z(n_122628503
		));
	notech_and3 i_54632877(.A(n_318691637), .B(n_315591668), .C(n_317991644)
		, .Z(n_124328520));
	notech_and4 i_94038272(.A(n_2329), .B(n_2328), .C(n_2324), .D(n_2327), .Z
		(n_128228559));
	notech_and4 i_93938273(.A(n_231591988), .B(n_2314), .C(n_2310), .D(n_2313
		), .Z(n_130528582));
	notech_and4 i_93838307(.A(n_2245), .B(n_2244), .C(n_2240), .D(n_2243), .Z
		(n_131228589));
	notech_and4 i_93738274(.A(n_2301), .B(n_2300), .C(n_2296), .D(n_2299), .Z
		(n_133728614));
	notech_and2 i_55347722(.A(n_28502), .B(n_184692037), .Z(n_139728674));
	notech_ao4 i_188847723(.A(n_301091813), .B(n_299891825), .C(n_30821), .D
		(n_61103), .Z(n_140128678));
	notech_ao4 i_188947724(.A(n_61110), .B(n_30822), .C(n_301091813), .D(n_26681
		), .Z(n_140228679));
	notech_and2 i_189947725(.A(n_305591768), .B(n_26700), .Z(n_140328680));
	notech_and3 i_190047726(.A(n_301891805), .B(n_300391820), .C(n_305691767
		), .Z(n_140428681));
	notech_or4 i_113(.A(calc_sz[0]), .B(calc_sz[3]), .C(n_58101), .D(n_27895
		), .Z(n_27896));
	notech_nor2 i_89347772(.A(n_308391740), .B(n_304791776), .Z(n_142728704)
		);
	notech_ao4 i_89447771(.A(n_304991774), .B(n_27746), .C(n_30822), .D(n_27754
		), .Z(n_142828705));
	notech_ao3 i_89847728(.A(n_104722311), .B(n_313591688), .C(n_306491759),
		 .Z(n_142928706));
	notech_and2 i_89947729(.A(n_1865), .B(n_306691757), .Z(n_143028707));
	notech_ao4 i_47532886(.A(n_32432), .B(n_61110), .C(n_319391630), .D(n_27552
		), .Z(n_146228739));
	notech_ao4 i_48232887(.A(n_32434), .B(n_61110), .C(n_59326), .D(n_26963)
		, .Z(n_146328740));
	notech_and2 i_55247735(.A(n_313191692), .B(n_313091693), .Z(n_146428741)
		);
	notech_ao4 i_188450696(.A(n_30821), .B(n_61109), .C(n_312191702), .D(n_312091703
		), .Z(n_146928746));
	notech_and3 i_188547736(.A(n_305491769), .B(n_312991694), .C(n_1857), .Z
		(n_147028747));
	notech_and3 i_189547737(.A(n_305591768), .B(n_312891695), .C(n_312591698
		), .Z(n_147128748));
	notech_and3 i_189647738(.A(n_305691767), .B(n_312791696), .C(n_312691697
		), .Z(n_147228749));
	notech_and2 i_54950719(.A(n_311791706), .B(n_311691707), .Z(n_148728764)
		);
	notech_and3 i_187850702(.A(n_312391700), .B(n_30803), .C(n_184392040), .Z
		(n_149128768));
	notech_ao4 i_187950700(.A(n_56950), .B(n_2510), .C(n_312291701), .D(n_311891705
		), .Z(n_149228769));
	notech_ao4 i_188050699(.A(n_30821), .B(n_60193), .C(n_312291701), .D(n_311991704
		), .Z(n_149328770));
	notech_and4 i_188150697(.A(n_59147), .B(n_59133), .C(n_304691777), .D(n_184292041
		), .Z(n_149428771));
	notech_and2 i_54232754(.A(n_59147), .B(n_59133), .Z(n_151028787));
	notech_and2 i_54832894(.A(n_317891645), .B(n_315691667), .Z(n_151128788)
		);
	notech_ao4 i_86432895(.A(n_59441), .B(n_27179), .C(n_2414), .D(n_26941),
		 .Z(n_151328790));
	notech_and2 i_86532896(.A(n_316691657), .B(n_316291661), .Z(n_151428791)
		);
	notech_and4 i_165135121(.A(n_57967), .B(n_56950), .C(n_60319), .D(n_1904
		), .Z(n_311591708));
	notech_or4 i_36222(.A(n_55581), .B(n_57082), .C(n_57064), .D(n_54974), .Z
		(n_311491709));
	notech_or4 i_36229(.A(n_55581), .B(n_316391660), .C(n_57082), .D(n_57064
		), .Z(n_311391710));
	notech_or4 i_56532742(.A(n_59393), .B(n_59402), .C(n_56684), .D(n_27577)
		, .Z(n_311291711));
	notech_or4 i_113032743(.A(n_60854), .B(n_32343), .C(n_317591648), .D(n_54974
		), .Z(n_311191712));
	notech_or2 i_117332744(.A(n_316191662), .B(n_54974), .Z(n_311091713));
	notech_nand3 i_31732470(.A(n_60138), .B(n_60193), .C(n_26983), .Z(n_32269
		));
	notech_and3 i_54732824(.A(n_60138), .B(n_60207), .C(n_60283), .Z(n_310991714
		));
	notech_or4 i_191650650(.A(n_57020), .B(n_311991704), .C(n_57042), .D(n_27712
		), .Z(n_310891715));
	notech_or4 i_191750649(.A(n_57020), .B(n_311891705), .C(n_57042), .D(n_27712
		), .Z(n_310791716));
	notech_or4 i_56641400(.A(n_56827), .B(n_56944), .C(n_27192), .D(n_27577)
		, .Z(n_310691717));
	notech_or4 i_180541249(.A(n_62844), .B(n_59469), .C(n_60931), .D(n_60207
		), .Z(n_310591718));
	notech_or4 i_3847661(.A(n_312191702), .B(n_57082), .C(n_57068), .D(n_54916
		), .Z(n_310491719));
	notech_or4 i_57532936(.A(n_59382), .B(n_59275), .C(n_32370), .D(instrc[
		115]), .Z(n_310391720));
	notech_nao3 i_33379(.A(n_60138), .B(n_60207), .C(n_32555), .Z(n_310291721
		));
	notech_nand2 i_33397(.A(n_319391630), .B(n_2492), .Z(n_310191722));
	notech_ao3 i_4347656(.A(n_30946), .B(n_2026), .C(n_303791786), .Z(n_27340
		));
	notech_nand2 i_29213(.A(n_62820), .B(opc_10[27]), .Z(n_310091723));
	notech_or4 i_5647643(.A(n_184892035), .B(n_57068), .C(n_57011), .D(n_54916
		), .Z(n_27329));
	notech_or4 i_62341309(.A(n_60969), .B(n_60958), .C(n_62836), .D(n_29596)
		, .Z(n_31456));
	notech_nao3 i_5547644(.A(n_56925), .B(n_313391690), .C(n_246791942), .Z(n_309891725
		));
	notech_and4 i_4147658(.A(n_57020), .B(n_57033), .C(n_28552), .D(n_26748)
		, .Z(n_309791726));
	notech_or4 i_192547685(.A(n_57055), .B(n_57011), .C(n_26770), .D(n_184992034
		), .Z(n_309691727));
	notech_nand2 i_2070(.A(n_60138), .B(n_60207), .Z(n_32270));
	notech_nao3 i_47832769(.A(n_60319), .B(n_56944), .C(n_308891735), .Z(n_309591728
		));
	notech_nand3 i_47632770(.A(n_60319), .B(n_1901), .C(n_56944), .Z(n_30803
		));
	notech_or4 i_47444591(.A(n_61171), .B(n_61160), .C(n_61151), .D(n_30821)
		, .Z(n_309491729));
	notech_nand3 i_27607(.A(n_246591944), .B(n_57055), .C(n_26832), .Z(n_309391730
		));
	notech_nao3 i_27707(.A(n_19065), .B(n_26983), .C(n_59326), .Z(n_309291731
		));
	notech_or4 i_27704(.A(n_61109), .B(n_2868), .C(n_62836), .D(n_62816), .Z
		(n_309191732));
	notech_or4 i_113532803(.A(n_101413114), .B(n_29179), .C(n_317391650), .D
		(n_316591658), .Z(n_309091733));
	notech_or2 i_137532804(.A(n_315891665), .B(n_316591658), .Z(n_308991734)
		);
	notech_ao3 i_4224(.A(n_29177), .B(n_59286), .C(n_59402), .Z(n_32408));
	notech_and3 i_4885(.A(n_59402), .B(n_59393), .C(n_318891635), .Z(n_32373
		));
	notech_and4 i_4832782(.A(n_59402), .B(n_59382), .C(n_29177), .D(n_59364)
		, .Z(n_32284));
	notech_ao3 i_4239(.A(n_59393), .B(n_59286), .C(n_59402), .Z(n_32286));
	notech_ao3 i_5132783(.A(instrc[115]), .B(n_319091633), .C(n_59382), .Z(n_32287
		));
	notech_ao3 i_5232784(.A(n_59382), .B(n_59364), .C(n_59275), .Z(n_32291)
		);
	notech_ao3 i_5632785(.A(instrc[115]), .B(n_318791636), .C(n_59382), .Z(n_32292
		));
	notech_and3 i_5832787(.A(n_59402), .B(n_29177), .C(n_59286), .Z(n_32295)
		);
	notech_ao3 i_5932788(.A(n_59382), .B(n_59373), .C(n_59275), .Z(n_32298)
		);
	notech_ao3 i_6032789(.A(n_56925), .B(n_29177), .C(n_59402), .Z(n_32299)
		);
	notech_and4 i_6132790(.A(n_59402), .B(n_59382), .C(n_29177), .D(n_59373)
		, .Z(n_32301));
	notech_ao3 i_6232792(.A(n_59393), .B(n_318891635), .C(n_59407), .Z(n_32304
		));
	notech_nand2 i_204453908(.A(read_data[29]), .B(n_60207), .Z(n_3883));
	notech_ao4 i_128153912(.A(n_1567), .B(n_176292077), .C(n_3996), .D(n_176092079
		), .Z(n_3885));
	notech_and4 i_145253929(.A(n_169992130), .B(n_1698), .C(n_169492133), .D
		(n_169792131), .Z(n_3981));
	notech_and4 i_145153930(.A(n_172492109), .B(n_1723), .C(n_171992112), .D
		(n_1722), .Z(n_3982));
	notech_and4 i_144953931(.A(n_173992096), .B(n_173892097), .C(n_173492099
		), .D(n_1737), .Z(n_3983));
	notech_or2 i_32371(.A(n_55735), .B(n_27757), .Z(n_27604));
	notech_or4 i_29447(.A(n_58101), .B(n_56970), .C(n_56827), .D(n_302891795
		), .Z(n_30528));
	notech_mux2 i_3011699(.S(n_60542), .A(regs_14[29]), .B(add_len_pc32[29])
		, .Z(add_len_pc[29]));
	notech_and2 i_7771(.A(n_168792138), .B(n_1479), .Z(n_3996));
	notech_or2 i_11132811(.A(n_58101), .B(n_56970), .Z(n_32382));
	notech_and2 i_85653963(.A(n_27753), .B(n_1478), .Z(n_3997));
	notech_and3 i_171653971(.A(n_1686), .B(n_26606), .C(n_26625), .Z(n_4005)
		);
	notech_ao4 i_114953973(.A(n_55735), .B(n_27746), .C(n_30565), .D(eval_flag
		), .Z(n_4007));
	notech_and3 i_109253974(.A(n_306691757), .B(n_308291741), .C(n_1475), .Z
		(n_4008));
	notech_and2 i_101253975(.A(n_26595), .B(n_1474), .Z(n_4009));
	notech_ao3 i_97053976(.A(n_246591944), .B(n_57068), .C(n_304991774), .Z(n_4010
		));
	notech_and2 i_89753977(.A(n_32352), .B(n_56675), .Z(n_4011));
	notech_and2 i_63853979(.A(n_4014), .B(n_1473), .Z(n_4013));
	notech_or4 i_46632807(.A(n_32378), .B(n_60193), .C(n_60986), .D(n_56944)
		, .Z(n_32371));
	notech_nao3 i_57953980(.A(n_56950), .B(n_32294), .C(n_56827), .Z(n_4014)
		);
	notech_and4 i_145053986(.A(n_168292141), .B(n_168192142), .C(n_167792145
		), .D(n_1680), .Z(n_4016));
	notech_and3 i_189241383(.A(n_26643), .B(n_26634), .C(n_26702), .Z(n_308891735
		));
	notech_and4 i_5732786(.A(n_59382), .B(n_59407), .C(n_59373), .D(n_59397)
		, .Z(n_32294));
	notech_and3 i_832781(.A(n_59382), .B(n_59364), .C(n_318791636), .Z(n_32280
		));
	notech_or4 i_192255508(.A(n_55581), .B(n_57082), .C(n_57055), .D(n_1434)
		, .Z(n_308791736));
	notech_nor2 i_930489(.A(n_32326), .B(n_32614), .Z(n_32316));
	notech_or4 i_47332798(.A(calc_sz[3]), .B(n_58062), .C(n_56858), .D(calc_sz
		[2]), .Z(n_308691737));
	notech_or4 i_56755526(.A(n_56827), .B(n_56553), .C(n_56944), .D(n_61131)
		, .Z(n_308591738));
	notech_or4 i_8792(.A(n_59397), .B(n_59407), .C(n_2479), .D(n_32351), .Z(n_308491739
		));
	notech_and3 i_50485(.A(fsm[3]), .B(n_60378), .C(n_2881), .Z(n_19086));
	notech_nor2 i_11938(.A(n_304991774), .B(n_304591778), .Z(n_308391740));
	notech_or2 i_11937(.A(n_304991774), .B(n_27746), .Z(n_308291741));
	notech_or2 i_136755511(.A(n_1433), .B(n_56463), .Z(n_27746));
	notech_nand2 i_32233(.A(n_26983), .B(n_60193), .Z(n_308091743));
	notech_nao3 i_32366(.A(n_246591944), .B(n_57068), .C(n_55735), .Z(n_307991744
		));
	notech_or4 i_137255510(.A(n_60975), .B(n_32614), .C(n_307691747), .D(n_60915
		), .Z(n_24590));
	notech_or4 i_35219(.A(n_55581), .B(n_306791756), .C(n_57082), .D(n_57051
		), .Z(n_307891745));
	notech_and3 i_189855558(.A(n_307591748), .B(n_305691767), .C(n_188857101
		), .Z(n_150728784));
	notech_and3 i_189755559(.A(n_305591768), .B(n_307291751), .C(n_188357100
		), .Z(n_150628783));
	notech_ao4 i_188755560(.A(n_61110), .B(n_30822), .C(n_306791756), .D(n_24590
		), .Z(n_150528782));
	notech_ao4 i_188655561(.A(n_30821), .B(n_61110), .C(n_307391750), .D(n_306791756
		), .Z(n_150428781));
	notech_and2 i_187555562(.A(n_26702), .B(n_59708), .Z(n_307791746));
	notech_ao3 i_3531(.A(n_60899), .B(n_62816), .C(n_2868), .Z(n_1903));
	notech_ao4 i_84155571(.A(n_62820), .B(n_60899), .C(n_60888), .D(n_24594)
		, .Z(n_307691747));
	notech_and4 i_4438305(.A(n_60975), .B(instrc[120]), .C(instrc[123]), .D(instrc
		[121]), .Z(n_32327));
	notech_or4 i_131555581(.A(n_60854), .B(n_32614), .C(n_307691747), .D(n_307491749
		), .Z(n_307591748));
	notech_and2 i_131655527(.A(n_24582), .B(n_24583), .Z(n_307491749));
	notech_and2 i_158555578(.A(n_59429), .B(n_305891765), .Z(n_307391750));
	notech_or2 i_131455582(.A(n_307391750), .B(n_307491749), .Z(n_307291751)
		);
	notech_mux2 i_123655583(.S(n_60319), .A(n_26983), .B(n_1438), .Z(n_307091753
		));
	notech_or2 i_163755572(.A(n_1433), .B(n_32327), .Z(n_306991754));
	notech_ao4 i_109155589(.A(n_1433), .B(n_32327), .C(n_59418), .D(n_27757)
		, .Z(n_306891755));
	notech_nor2 i_89655594(.A(n_2349), .B(n_1440), .Z(n_306791756));
	notech_or2 i_81955603(.A(n_27746), .B(n_306591758), .Z(n_306691757));
	notech_and3 i_97355591(.A(n_56848), .B(n_1441), .C(n_305191772), .Z(n_306591758
		));
	notech_nor2 i_81855604(.A(n_306591758), .B(n_304591778), .Z(n_306491759)
		);
	notech_ao3 i_10932812(.A(calc_sz[0]), .B(n_58101), .C(n_2937), .Z(n_32386
		));
	notech_and2 i_80855605(.A(n_26962), .B(n_56983), .Z(n_306391760));
	notech_nor2 i_78555606(.A(n_234791985), .B(n_1442), .Z(n_24589));
	notech_ao4 i_78455607(.A(n_56843), .B(n_61133), .C(n_32351), .D(n_32280)
		, .Z(n_24582));
	notech_ao4 i_78355608(.A(n_61136), .B(n_27024), .C(n_32355), .D(n_32280)
		, .Z(n_24583));
	notech_and3 i_199555610(.A(n_26625), .B(n_27753), .C(n_1686), .Z(n_306291761
		));
	notech_nor2 i_3511(.A(n_2873), .B(n_2872), .Z(n_1902));
	notech_ao3 i_66755611(.A(n_27377), .B(n_60321), .C(n_26643), .Z(n_306191762
		));
	notech_or4 i_66555612(.A(n_59397), .B(n_59407), .C(n_59355), .D(n_32355)
		, .Z(n_306091763));
	notech_or2 i_166255570(.A(n_307691747), .B(n_32316), .Z(n_305991764));
	notech_ao4 i_60255614(.A(n_307691747), .B(n_32316), .C(n_59418), .D(n_24594
		), .Z(n_305891765));
	notech_ao3 i_3523(.A(n_60904), .B(n_60931), .C(n_2870), .Z(n_1904));
	notech_or4 i_68955539(.A(n_59397), .B(n_59407), .C(n_59355), .D(n_32347)
		, .Z(n_305791766));
	notech_and3 i_55055619(.A(n_308491739), .B(n_306091763), .C(n_305791766)
		, .Z(n_150228779));
	notech_or4 i_54555620(.A(n_61136), .B(n_60193), .C(n_59708), .D(n_56950)
		, .Z(n_305691767));
	notech_ao3 i_3514(.A(n_62870), .B(n_32470), .C(n_2872), .Z(n_1901));
	notech_and3 i_187032810(.A(n_56959), .B(n_26962), .C(n_56983), .Z(n_32380
		));
	notech_or4 i_54455621(.A(n_308891735), .B(n_61136), .C(n_60193), .D(n_56950
		), .Z(n_305591768));
	notech_nao3 i_54355622(.A(n_60138), .B(n_60316), .C(n_30822), .Z(n_305491769
		));
	notech_or4 i_47232795(.A(n_32378), .B(n_56959), .C(n_60193), .D(\opcode[3] 
		), .Z(n_305391770));
	notech_nor2 i_47032802(.A(n_56854), .B(n_56983), .Z(n_305291771));
	notech_ao4 i_50055634(.A(n_56854), .B(n_56983), .C(n_56675), .D(n_32294)
		, .Z(n_305191772));
	notech_or4 i_47132808(.A(n_32378), .B(n_60193), .C(\opcode[3] ), .D(n_56941
		), .Z(n_305091773));
	notech_ao4 i_49955635(.A(n_56854), .B(n_56941), .C(n_56688), .D(n_32294)
		, .Z(n_304991774));
	notech_and2 i_23130(.A(n_27753), .B(n_26625), .Z(n_304891775));
	notech_ao3 i_47955637(.A(n_56983), .B(n_314291681), .C(n_304891775), .Z(n_304791776
		));
	notech_or4 i_47755638(.A(n_61175), .B(n_61160), .C(n_61151), .D(n_30822)
		, .Z(n_304691777));
	notech_and2 i_38355639(.A(n_306891755), .B(n_59429), .Z(n_304591778));
	notech_nand2 i_199055507(.A(n_29658), .B(n_57068), .Z(n_30854));
	notech_ao3 i_19055642(.A(n_57011), .B(n_57068), .C(n_55581), .Z(n_24594)
		);
	notech_and4 i_12355645(.A(n_57020), .B(n_57042), .C(n_57082), .D(n_57068
		), .Z(n_27757));
	notech_and3 i_732780(.A(n_59407), .B(n_59397), .C(n_59286), .Z(n_32279)
		);
	notech_nand2 i_198271100(.A(n_60931), .B(n_62836), .Z(n_32448));
	notech_nand2 i_198471099(.A(n_62802), .B(n_62836), .Z(n_32467));
	notech_nand2 i_13658357(.A(n_54834), .B(n_56163), .Z(n_27335));
	notech_nand2 i_13558358(.A(n_54834), .B(n_56172), .Z(n_27334));
	notech_and4 i_1032821(.A(n_59407), .B(n_59382), .C(n_59393), .D(n_29178)
		, .Z(n_32616));
	notech_or4 i_11558376(.A(n_28532), .B(n_61136), .C(n_60193), .D(n_56163)
		, .Z(n_28530));
	notech_or4 i_11458377(.A(n_28532), .B(n_61136), .C(n_60193), .D(\eflags[10] 
		), .Z(n_28527));
	notech_nao3 i_793(.A(n_2825), .B(n_2838), .C(n_2883), .Z(n_28533));
	notech_ao4 i_50155633(.A(n_56858), .B(n_56959), .C(n_56813), .D(n_32294)
		, .Z(n_27761));
	notech_nor2 i_134558493(.A(n_304191782), .B(n_59344), .Z(n_28546));
	notech_nand2 i_23413(.A(n_32347), .B(n_32351), .Z(n_304491779));
	notech_nao3 i_11474(.A(n_304491779), .B(n_59286), .C(n_246791942), .Z(n_304391780
		));
	notech_or4 i_46532797(.A(calc_sz[3]), .B(n_2938), .C(n_56827), .D(calc_sz
		[2]), .Z(n_32352));
	notech_or4 i_46732794(.A(n_32378), .B(n_56959), .C(n_60193), .D(n_60986)
		, .Z(n_32348));
	notech_and2 i_259758504(.A(n_32352), .B(n_56813), .Z(n_304291781));
	notech_nor2 i_4738265(.A(n_32614), .B(n_32342), .Z(n_32335));
	notech_ao4 i_85858514(.A(n_62820), .B(n_60904), .C(n_60888), .D(n_28551)
		, .Z(n_304191782));
	notech_ao3 i_1138268(.A(n_60975), .B(n_60915), .C(n_32614), .Z(n_32612)
		);
	notech_or4 i_129458523(.A(n_55581), .B(n_57051), .C(n_57011), .D(n_54934
		), .Z(n_25884));
	notech_nand2 i_119958527(.A(n_303791786), .B(n_27346), .Z(n_27163));
	notech_ao4 i_95558534(.A(n_59418), .B(n_27988), .C(n_60863), .D(n_28533)
		, .Z(n_304091783));
	notech_xor2 i_90558536(.A(n_62776), .B(n_60904), .Z(n_303991784));
	notech_and3 i_84758538(.A(n_28543), .B(n_301091813), .C(n_28545), .Z(n_303891785
		));
	notech_ao4 i_74958539(.A(n_305091773), .B(n_61136), .C(n_32370), .D(n_32279
		), .Z(n_303791786));
	notech_ao4 i_74558541(.A(n_56843), .B(n_61136), .C(n_32351), .D(n_32279)
		, .Z(n_27346));
	notech_or4 i_67058546(.A(n_246791942), .B(n_59355), .C(n_56675), .D(n_61136
		), .Z(n_28502));
	notech_or4 i_66858547(.A(n_59382), .B(n_246791942), .C(n_32355), .D(n_59373
		), .Z(n_303691787));
	notech_or4 i_57458554(.A(n_56827), .B(n_56941), .C(n_61136), .D(n_56570)
		, .Z(n_303591788));
	notech_or4 i_57058555(.A(n_56827), .B(n_56944), .C(n_61138), .D(n_56547)
		, .Z(n_27319));
	notech_or2 i_163658507(.A(n_27353), .B(n_27349), .Z(n_51735313));
	notech_nand2 i_170347755(.A(n_26613), .B(n_26614), .Z(n_303491789));
	notech_ao3 i_1238259(.A(n_60975), .B(n_60915), .C(n_32343), .Z(n_32318)
		);
	notech_and4 i_12558491(.A(n_57020), .B(n_57033), .C(n_57051), .D(n_57078
		), .Z(n_27353));
	notech_and4 i_12158557(.A(n_57020), .B(n_57033), .C(n_57064), .D(n_57078
		), .Z(n_28551));
	notech_nand2 i_198571098(.A(n_60904), .B(n_62816), .Z(n_32650));
	notech_or4 i_29410(.A(n_58101), .B(n_246691943), .C(n_60193), .D(n_59708
		), .Z(n_30565));
	notech_and4 i_143044523(.A(n_1967), .B(n_1966), .C(n_196257103), .D(n_1965
		), .Z(n_303391790));
	notech_and2 i_63558549(.A(n_303591788), .B(n_184692037), .Z(n_303291791)
		);
	notech_and4 i_91838293(.A(n_2273), .B(n_2272), .C(n_2268), .D(n_2271), .Z
		(n_303191792));
	notech_and4 i_145332876(.A(n_2505), .B(n_2504), .C(n_2500), .D(n_2503), 
		.Z(n_303091793));
	notech_and2 i_55147731(.A(n_304391780), .B(n_303691787), .Z(n_144428721)
		);
	notech_ao4 i_189347733(.A(n_56950), .B(n_1452), .C(n_184892035), .D(n_313491689
		), .Z(n_145028727));
	notech_ao4 i_6047639(.A(n_61110), .B(n_30822), .C(n_303791786), .D(n_26815
		), .Z(n_144928726));
	notech_and4 i_94138306(.A(n_2259), .B(n_2258), .C(n_2254), .D(n_2257), .Z
		(n_302991794));
	notech_and3 i_189447734(.A(n_305691767), .B(n_52335319), .C(n_313291691)
		, .Z(n_145128728));
	notech_ao4 i_188247732(.A(n_30821), .B(n_61110), .C(n_313491689), .D(n_303791786
		), .Z(n_144828725));
	notech_nand2 i_29887(.A(n_62798), .B(opc[11]), .Z(n_30088));
	notech_and4 i_143441318(.A(n_2071), .B(n_2070), .C(n_2066), .D(n_2069), 
		.Z(n_302891795));
	notech_and3 i_109441354(.A(n_299591828), .B(n_300791816), .C(n_313791686
		), .Z(n_302791796));
	notech_and3 i_109341353(.A(n_313891685), .B(n_2993), .C(n_315091673), .Z
		(n_302691797));
	notech_and3 i_64841352(.A(n_303691787), .B(n_2025), .C(n_27319), .Z(n_302591798
		));
	notech_and4 i_92238289(.A(n_2287), .B(n_2286), .C(n_2282), .D(n_2285), .Z
		(n_302491799));
	notech_and2 i_64441362(.A(n_3857), .B(n_2000), .Z(n_302391800));
	notech_and2 i_99341364(.A(n_3877), .B(n_3876), .Z(n_302291801));
	notech_ao4 i_99241363(.A(n_59441), .B(n_27029), .C(n_3879), .D(n_26670),
		 .Z(n_302191802));
	notech_and4 i_92438308(.A(n_2231), .B(n_2230), .C(n_2226), .D(n_2229), .Z
		(n_302091803));
	notech_and2 i_101041365(.A(n_3858), .B(n_2001), .Z(n_301991804));
	notech_ao4 i_73858544(.A(n_305391770), .B(n_61138), .C(n_32347), .D(n_32616
		), .Z(n_28545));
	notech_nand2 i_261721(.A(n_26683), .B(n_28546), .Z(n_301891805));
	notech_or4 i_192461726(.A(n_57078), .B(n_57064), .C(n_54916), .D(n_131292192
		), .Z(n_301791806));
	notech_ao4 i_74758540(.A(n_305391770), .B(n_61138), .C(n_32347), .D(n_32279
		), .Z(n_27349));
	notech_and4 i_143641405(.A(n_2054), .B(n_2053), .C(n_2049), .D(n_2052), 
		.Z(n_301691807));
	notech_and4 i_1421859(.A(n_1411), .B(n_1410), .C(n_132092184), .D(n_1414
		), .Z(n_301591808));
	notech_and4 i_1221537(.A(n_1401), .B(n_1400), .C(n_1399), .D(n_1404), .Z
		(n_301491809));
	notech_nand2 i_3121556(.A(n_1392), .B(n_1387), .Z(n_301391810));
	notech_and4 i_821341(.A(n_1378), .B(n_1377), .C(n_1356), .D(n_1381), .Z(n_301291811
		));
	notech_ao4 i_74832889(.A(n_32347), .B(n_32286), .C(n_305391770), .D(n_61138
		), .Z(n_26616));
	notech_and2 i_50437(.A(n_60378), .B(n_272491901), .Z(n_1914992224));
	notech_ao4 i_73958543(.A(n_305091773), .B(n_61138), .C(n_32370), .D(n_32616
		), .Z(n_301091813));
	notech_nand2 i_12542(.A(n_26748), .B(n_28546), .Z(n_300991814));
	notech_ao4 i_73658545(.A(n_61136), .B(n_27024), .C(n_32355), .D(n_32616)
		, .Z(n_28544));
	notech_ao4 i_74358542(.A(n_61136), .B(n_27024), .C(n_32355), .D(n_32279)
		, .Z(n_300891815));
	notech_or2 i_11289(.A(n_300891815), .B(n_26815), .Z(n_300791816));
	notech_or2 i_179158494(.A(n_304191782), .B(n_32612), .Z(n_300591818));
	notech_ao4 i_106061811(.A(n_304191782), .B(n_32612), .C(n_59418), .D(n_28551
		), .Z(n_300491819));
	notech_nand2 i_105361812(.A(n_28542), .B(n_28546), .Z(n_300391820));
	notech_ao4 i_105261813(.A(n_61110), .B(n_30825), .C(n_28544), .D(n_300491819
		), .Z(n_300291821));
	notech_or2 i_12334(.A(n_28544), .B(n_26681), .Z(n_300191822));
	notech_and2 i_105161814(.A(n_300191822), .B(n_2991), .Z(n_300091823));
	notech_nand2 i_91061824(.A(n_28332), .B(n_28546), .Z(n_299991824));
	notech_and2 i_148244575(.A(n_59429), .B(n_300491819), .Z(n_299891825));
	notech_nand2 i_83058492(.A(n_28543), .B(n_301091813), .Z(n_28332));
	notech_nand2 i_90961825(.A(n_28332), .B(n_27301), .Z(n_299791826));
	notech_ao4 i_59761833(.A(n_1416), .B(n_32318), .C(n_59418), .D(n_27353),
		 .Z(n_299691827));
	notech_nand3 i_58361834(.A(n_1476), .B(n_60138), .C(n_60316), .Z(n_299591828
		));
	notech_or4 i_58261835(.A(n_308891735), .B(n_56959), .C(n_61138), .D(n_60193
		), .Z(n_102035816));
	notech_ao4 i_46941401(.A(n_1902), .B(n_1904), .C(n_56950), .D(n_26626), 
		.Z(n_299491829));
	notech_nand3 i_58161836(.A(n_60133), .B(n_60316), .C(n_299491829), .Z(n_2993
		));
	notech_or4 i_58061837(.A(n_58101), .B(n_56970), .C(n_61110), .D(n_59708)
		, .Z(n_102135817));
	notech_or4 i_56961838(.A(n_308891735), .B(n_61136), .C(n_60212), .D(n_56979
		), .Z(n_2992));
	notech_or4 i_56861839(.A(n_61133), .B(n_60212), .C(n_59708), .D(n_56979)
		, .Z(n_2991));
	notech_nao3 i_49655636(.A(n_60138), .B(n_60316), .C(n_30821), .Z(n_2990)
		);
	notech_and2 i_49761840(.A(n_2990), .B(n_131692188), .Z(n_298991830));
	notech_or4 i_889(.A(n_61175), .B(n_61160), .C(n_61151), .D(n_61133), .Z(n_32855
		));
	notech_ao4 i_27835149(.A(n_1903), .B(n_1901), .C(n_26627), .D(n_32380), 
		.Z(n_2988));
	notech_nand3 i_48161841(.A(n_60138), .B(n_60316), .C(n_2988), .Z(n_28222
		));
	notech_and4 i_1019(.A(n_2973), .B(n_2963), .C(n_298557106), .D(n_271791908
		), .Z(n_298691832));
	notech_and4 i_1017(.A(n_271491911), .B(n_2982), .C(n_297891837), .D(n_272091905
		), .Z(n_298557106));
	notech_and4 i_1006(.A(n_297991836), .B(n_2707), .C(n_271291913), .D(n_270491919
		), .Z(n_2982));
	notech_ao4 i_996(.A(n_22579), .B(n_28882), .C(n_22571), .D(n_56329), .Z(n_297991836
		));
	notech_and3 i_1009(.A(n_2976), .B(n_271191914), .C(n_271391912), .Z(n_297891837
		));
	notech_ao4 i_1001(.A(n_22585), .B(n_28914), .C(n_22594), .D(n_28775), .Z
		(n_2976));
	notech_and4 i_1008(.A(n_2970), .B(n_2965), .C(n_2964), .D(n_271091915), 
		.Z(n_2973));
	notech_and4 i_998(.A(n_2966), .B(n_2969), .C(n_2696), .D(n_2697), .Z(n_2970
		));
	notech_ao4 i_995(.A(n_22582), .B(n_28638), .C(n_22572), .D(n_28657), .Z(n_2969
		));
	notech_ao4 i_992(.A(n_55773), .B(n_29627), .C(n_57537), .D(nbus_11295[5]
		), .Z(n_2966));
	notech_ao4 i_997(.A(n_22590), .B(n_29626), .C(n_22591), .D(n_28743), .Z(n_2965
		));
	notech_ao4 i_1003(.A(n_22322), .B(n_2691), .C(n_57155), .D(\nbus_11358[13] 
		), .Z(n_2964));
	notech_ao4 i_1011(.A(n_23031), .B(n_27680), .C(n_56073), .D(n_57848), .Z
		(n_2963));
	notech_ao4 i_1015(.A(n_22309), .B(n_28631), .C(n_27782), .D(n_28669), .Z
		(n_2961));
	notech_and4 i_569(.A(n_62844), .B(n_60931), .C(n_60316), .D(n_26782), .Z
		(n_2956));
	notech_and4 i_568(.A(n_62844), .B(n_60931), .C(n_60316), .D(n_57967), .Z
		(n_295591839));
	notech_and4 i_562(.A(n_60904), .B(n_60933), .C(n_60316), .D(n_32323), .Z
		(n_2952));
	notech_ao4 i_560(.A(n_32343), .B(n_32342), .C(n_60854), .D(n_32614), .Z(n_2950
		));
	notech_or4 i_31(.A(n_58033), .B(n_32323), .C(n_59429), .D(n_60212), .Z(n_2949
		));
	notech_and2 i_87(.A(sign_div), .B(opd[31]), .Z(n_2947));
	notech_nand3 i_546(.A(n_27986), .B(n_59205), .C(n_59187), .Z(n_2946));
	notech_ao3 i_543(.A(n_60378), .B(n_32384), .C(n_61151), .Z(n_2944));
	notech_or4 i_531(.A(n_60274), .B(n_2825), .C(n_27132), .D(\opcode[3] ), 
		.Z(n_2941));
	notech_and4 i_27710(.A(n_18906874), .B(n_26702), .C(n_26643), .D(n_26602
		), .Z(n_2939));
	notech_nand2 i_529(.A(n_58101), .B(n_27894), .Z(n_2938));
	notech_or2 i_27585(.A(calc_sz[3]), .B(calc_sz[2]), .Z(n_2937));
	notech_or2 i_513(.A(n_293491842), .B(n_18964), .Z(n_293591841));
	notech_nand3 i_1205(.A(n_19093), .B(n_19072), .C(n_60207), .Z(n_293491842
		));
	notech_or4 i_489(.A(ecx[17]), .B(ecx[16]), .C(ecx[19]), .D(ecx[18]), .Z(n_2929
		));
	notech_or4 i_488(.A(ecx[21]), .B(ecx[20]), .C(ecx[23]), .D(ecx[22]), .Z(n_2926
		));
	notech_or4 i_487(.A(ecx[25]), .B(ecx[24]), .C(ecx[27]), .D(ecx[26]), .Z(n_2922
		));
	notech_or4 i_486(.A(ecx[30]), .B(ecx[29]), .C(ecx[28]), .D(ecx[31]), .Z(n_291991845
		));
	notech_or4 i_3430135(.A(n_291491850), .B(n_291191853), .C(n_2907), .D(n_290491857
		), .Z(n_291691848));
	notech_or4 i_475(.A(ecx[1]), .B(ecx[0]), .C(ecx[3]), .D(ecx[2]), .Z(n_291491850
		));
	notech_or4 i_474(.A(ecx[7]), .B(ecx[6]), .C(ecx[5]), .D(ecx[4]), .Z(n_291191853
		));
	notech_or4 i_473(.A(ecx[11]), .B(ecx[9]), .C(ecx[8]), .D(ecx[10]), .Z(n_2907
		));
	notech_or4 i_472(.A(ecx[13]), .B(ecx[12]), .C(ecx[15]), .D(ecx[14]), .Z(n_290491857
		));
	notech_and2 i_442(.A(n_1871), .B(n_2654), .Z(n_289791858));
	notech_nao3 i_1811(.A(fsm[1]), .B(fsm[3]), .C(fsm[0]), .Z(n_2896));
	notech_nao3 i_422(.A(n_2649), .B(n_32695), .C(n_27125), .Z(n_2895));
	notech_or4 i_220(.A(n_2877), .B(n_60874), .C(n_2864), .D(n_32462), .Z(n_2893
		));
	notech_or4 i_1784(.A(n_27123), .B(n_27170), .C(n_62870), .D(\opcode[3] )
		, .Z(n_2888));
	notech_nor2 i_1371(.A(n_61160), .B(n_61175), .Z(n_2885));
	notech_or4 i_26997(.A(n_60274), .B(n_2839), .C(n_32747), .D(\opcode[3] )
		, .Z(n_2884));
	notech_or4 i_1668(.A(n_27123), .B(n_27170), .C(n_60874), .D(n_60986), .Z
		(n_2883));
	notech_nor2 i_1535(.A(fsm[0]), .B(n_27717), .Z(n_2881));
	notech_and2 i_1369(.A(n_61160), .B(n_61175), .Z(n_2880));
	notech_or2 i_1364(.A(n_2825), .B(n_2838), .Z(n_2877));
	notech_nand2 i_1528(.A(n_32695), .B(n_2864), .Z(n_2875));
	notech_or4 i_388(.A(n_2825), .B(n_27132), .C(n_2864), .D(n_62870), .Z(n_2873
		));
	notech_or4 i_26939(.A(n_60933), .B(n_60904), .C(n_32695), .D(\opcode[3] 
		), .Z(n_2872));
	notech_or4 i_381(.A(n_2825), .B(n_2869), .C(n_27132), .D(n_2864), .Z(n_2870
		));
	notech_nand3 i_380(.A(n_27123), .B(\opcode[3] ), .C(n_62870), .Z(n_2869)
		);
	notech_or4 i_219(.A(n_32695), .B(n_60986), .C(n_62870), .D(n_27125), .Z(n_2868
		));
	notech_and4 i_627965(.A(n_2852), .B(n_2861), .C(n_2617), .D(n_2604), .Z(n_2864
		));
	notech_ao3 i_310(.A(n_2859), .B(n_2858), .C(n_2614), .Z(n_2861));
	notech_ao4 i_306(.A(n_275591872), .B(n_29132), .C(n_273591890), .D(n_29650
		), .Z(n_2859));
	notech_and4 i_307(.A(n_2855), .B(n_2854), .C(n_2853), .D(n_2613), .Z(n_2858
		));
	notech_ao4 i_302(.A(n_275791870), .B(n_29123), .C(n_29172), .D(n_273791888
		), .Z(n_2855));
	notech_ao4 i_301(.A(n_274891879), .B(n_29156), .C(n_274491883), .D(n_29164
		), .Z(n_2854));
	notech_ao4 i_303(.A(n_275191876), .B(n_29140), .C(n_272791898), .D(n_29636
		), .Z(n_2853));
	notech_ao4 i_309(.A(n_273191894), .B(n_29635), .C(n_275291875), .D(n_29148
		), .Z(n_2852));
	notech_ao3 i_283(.A(n_2847), .B(n_2846), .C(n_2600), .Z(n_2849));
	notech_ao4 i_279(.A(n_275591872), .B(n_29134), .C(n_273591890), .D(n_29649
		), .Z(n_2847));
	notech_and4 i_280(.A(n_2843), .B(n_2842), .C(n_2841), .D(n_2599), .Z(n_2846
		));
	notech_ao4 i_274(.A(n_275791870), .B(n_29125), .C(n_29174), .D(n_273791888
		), .Z(n_2843));
	notech_ao4 i_273(.A(n_274891879), .B(n_29158), .C(n_274491883), .D(n_29166
		), .Z(n_2842));
	notech_ao4 i_276(.A(n_275191876), .B(n_29142), .C(n_272791898), .D(n_29638
		), .Z(n_2841));
	notech_ao4 i_282(.A(n_273191894), .B(n_29637), .C(n_275291875), .D(n_29150
		), .Z(n_2840));
	notech_nand3 i_38870661(.A(instrc[99]), .B(n_139588894), .C(n_94688445),
		 .Z(n_94588444));
	notech_nand2 i_071044(.A(instrc[98]), .B(instrc[97]), .Z(n_94688445));
	notech_ao4 i_90170148(.A(n_154379047), .B(n_27777), .C(n_27107), .D(n_27443
		), .Z(n_132988828));
	notech_ao4 i_90070149(.A(n_154179045), .B(n_56145), .C(n_154279046), .D(n_27739
		), .Z(n_133088829));
	notech_ao4 i_89970150(.A(n_154379047), .B(n_27779), .C(n_27107), .D(n_27445
		), .Z(n_133188830));
	notech_ao4 i_89870151(.A(n_154179045), .B(n_56190), .C(n_154279046), .D(n_27740
		), .Z(n_133288831));
	notech_ao4 i_89770152(.A(n_154379047), .B(n_27780), .C(n_27107), .D(n_27447
		), .Z(n_133388832));
	notech_ao4 i_89670153(.A(n_154179045), .B(n_29679), .C(n_154279046), .D(n_27741
		), .Z(n_133488833));
	notech_ao4 i_89570154(.A(n_154379047), .B(n_27785), .C(n_27107), .D(n_27451
		), .Z(n_133588834));
	notech_ao4 i_89470155(.A(n_154179045), .B(n_56257), .C(n_154279046), .D(n_27743
		), .Z(n_133688835));
	notech_ao4 i_86570184(.A(n_154379047), .B(n_27801), .C(n_27107), .D(n_27483
		), .Z(n_133788836));
	notech_ao4 i_86470185(.A(n_154179045), .B(n_29659), .C(n_154279046), .D(n_27763
		), .Z(n_133888837));
	notech_ao4 i_86370186(.A(n_154379047), .B(n_27802), .C(n_27107), .D(n_27485
		), .Z(n_133988838));
	notech_ao4 i_86270187(.A(n_154179045), .B(n_29591), .C(n_154279046), .D(n_27764
		), .Z(n_134088839));
	notech_ao4 i_86170188(.A(n_154379047), .B(n_27803), .C(n_27107), .D(n_27487
		), .Z(n_134188840));
	notech_ao4 i_86070189(.A(n_154179045), .B(n_29619), .C(n_154279046), .D(n_27765
		), .Z(n_134288841));
	notech_ao4 i_85970190(.A(n_349880999), .B(n_27766), .C(n_3914), .D(n_27422
		), .Z(n_134388842));
	notech_ao4 i_85870191(.A(n_349981000), .B(n_30551), .C(n_349780998), .D(n_27728
		), .Z(n_134488843));
	notech_ao4 i_85770192(.A(n_349880999), .B(n_27767), .C(n_3914), .D(n_27424
		), .Z(n_134588844));
	notech_ao4 i_85670193(.A(n_349981000), .B(n_30550), .C(n_349780998), .D(n_27729
		), .Z(n_134688845));
	notech_ao4 i_85570194(.A(n_349880999), .B(n_27775), .C(n_3914), .D(n_27439
		), .Z(n_134788846));
	notech_ao4 i_85470195(.A(n_349981000), .B(n_30549), .C(n_349780998), .D(n_27737
		), .Z(n_134888847));
	notech_ao4 i_85370196(.A(n_349880999), .B(n_27779), .C(n_3914), .D(n_27445
		), .Z(n_134988848));
	notech_ao4 i_85270197(.A(n_349981000), .B(n_30548), .C(n_349780998), .D(n_27740
		), .Z(n_135088849));
	notech_ao4 i_85170198(.A(n_349880999), .B(n_27780), .C(n_3914), .D(n_27447
		), .Z(n_135188850));
	notech_ao4 i_85070199(.A(n_349981000), .B(n_30547), .C(n_349780998), .D(n_27741
		), .Z(n_135288851));
	notech_ao4 i_84970200(.A(n_349981000), .B(n_30546), .C(n_3914), .D(n_27449
		), .Z(n_135388852));
	notech_ao4 i_84870201(.A(n_349780998), .B(n_27742), .C(n_349880999), .D(n_27783
		), .Z(n_135488853));
	notech_ao4 i_84770202(.A(n_349880999), .B(n_27785), .C(n_3914), .D(n_27451
		), .Z(n_135588854));
	notech_ao4 i_84670203(.A(n_349981000), .B(n_30545), .C(n_349780998), .D(n_27743
		), .Z(n_135688855));
	notech_ao4 i_84570204(.A(n_349880999), .B(n_27786), .C(n_3914), .D(n_27453
		), .Z(n_135788856));
	notech_ao4 i_84470205(.A(n_349981000), .B(n_30544), .C(n_349780998), .D(n_27744
		), .Z(n_135888857));
	notech_ao4 i_84370206(.A(n_349880999), .B(n_27787), .C(n_3914), .D(n_27455
		), .Z(n_135988858));
	notech_ao4 i_84270207(.A(n_349981000), .B(n_30543), .C(n_349780998), .D(n_27745
		), .Z(n_136088859));
	notech_ao4 i_84170208(.A(n_349880999), .B(n_27788), .C(n_3914), .D(n_27457
		), .Z(n_136188860));
	notech_ao4 i_84070209(.A(n_349981000), .B(n_30542), .C(n_349780998), .D(n_27747
		), .Z(n_136288861));
	notech_ao4 i_83970210(.A(n_349880999), .B(n_27789), .C(n_3914), .D(n_27459
		), .Z(n_136388862));
	notech_ao4 i_83870211(.A(n_349981000), .B(n_30541), .C(n_349780998), .D(n_27748
		), .Z(n_136488863));
	notech_ao4 i_83770212(.A(n_349880999), .B(n_27790), .C(n_3914), .D(n_27461
		), .Z(n_136588864));
	notech_ao4 i_83670213(.A(n_349981000), .B(n_30540), .C(n_349780998), .D(n_27749
		), .Z(n_136688865));
	notech_ao4 i_83570214(.A(n_349880999), .B(n_27791), .C(n_3914), .D(n_27463
		), .Z(n_136788866));
	notech_ao4 i_83470215(.A(n_349981000), .B(n_30539), .C(n_349780998), .D(n_27750
		), .Z(n_136888867));
	notech_ao4 i_83370216(.A(n_349880999), .B(n_27792), .C(n_56894), .D(n_27465
		), .Z(n_136988868));
	notech_ao4 i_83270217(.A(n_349981000), .B(n_30538), .C(n_349780998), .D(n_27751
		), .Z(n_137088869));
	notech_ao4 i_83170218(.A(n_349880999), .B(n_27793), .C(n_56894), .D(n_27469
		), .Z(n_137188870));
	notech_ao4 i_83070219(.A(n_349981000), .B(n_30537), .C(n_349780998), .D(n_27752
		), .Z(n_137288871));
	notech_ao4 i_82970220(.A(n_53890), .B(n_27794), .C(n_56894), .D(n_27471)
		, .Z(n_137388872));
	notech_ao4 i_82870221(.A(n_349981000), .B(n_30536), .C(n_53901), .D(n_27755
		), .Z(n_137488873));
	notech_ao4 i_82770222(.A(n_53890), .B(n_27795), .C(n_56894), .D(n_27473)
		, .Z(n_137588874));
	notech_ao4 i_82670223(.A(n_54020), .B(n_30535), .C(n_53901), .D(n_27756)
		, .Z(n_137688875));
	notech_ao4 i_82570224(.A(n_53890), .B(n_27797), .C(n_56894), .D(n_27475)
		, .Z(n_137788876));
	notech_ao4 i_82470225(.A(n_54020), .B(n_30534), .C(n_53901), .D(n_27758)
		, .Z(n_137888877));
	notech_ao4 i_82370226(.A(n_53890), .B(n_27798), .C(n_56894), .D(n_27477)
		, .Z(n_137988878));
	notech_ao4 i_82270227(.A(n_54020), .B(n_30533), .C(n_53901), .D(n_27759)
		, .Z(n_138088879));
	notech_ao4 i_82170228(.A(n_53890), .B(n_27799), .C(n_56894), .D(n_27479)
		, .Z(n_138188880));
	notech_ao4 i_82070229(.A(n_54020), .B(n_30532), .C(n_53901), .D(n_27760)
		, .Z(n_138288881));
	notech_ao4 i_81970230(.A(n_53890), .B(n_27800), .C(n_56894), .D(n_27481)
		, .Z(n_138388882));
	notech_ao4 i_81870231(.A(n_54020), .B(n_30531), .C(n_53901), .D(n_27762)
		, .Z(n_138488883));
	notech_ao4 i_81770232(.A(n_53890), .B(n_27801), .C(n_56894), .D(n_27483)
		, .Z(n_138588884));
	notech_ao4 i_81670233(.A(n_54020), .B(n_30530), .C(n_53901), .D(n_27763)
		, .Z(n_138688885));
	notech_ao4 i_81570234(.A(n_53890), .B(n_27802), .C(n_56894), .D(n_27485)
		, .Z(n_138788886));
	notech_ao4 i_81470235(.A(n_54020), .B(n_30529), .C(n_53901), .D(n_27764)
		, .Z(n_138888887));
	notech_ao4 i_81370236(.A(n_152889027), .B(n_27791), .C(n_3921), .D(n_27463
		), .Z(n_138988888));
	notech_ao4 i_81270237(.A(n_152689025), .B(n_30527), .C(n_152789026), .D(n_27750
		), .Z(n_139088889));
	notech_ao4 i_81170238(.A(n_152889027), .B(n_27792), .C(n_3921), .D(n_27465
		), .Z(n_139188890));
	notech_ao4 i_81070239(.A(n_152689025), .B(n_30526), .C(n_152789026), .D(n_27751
		), .Z(n_139288891));
	notech_or4 i_9371045(.A(n_29628), .B(instrc[98]), .C(n_29639), .D(instrc
		[96]), .Z(n_139488893));
	notech_mux2 i_16722(.S(instrc[97]), .A(instrc[98]), .B(n_29641), .Z(n_139588894
		));
	notech_nand2 i_7871046(.A(n_56888), .B(n_94588444), .Z(n_139788896));
	notech_ao4 i_80670243(.A(n_139788896), .B(n_30525), .C(n_27728), .D(n_139488893
		), .Z(n_139888897));
	notech_or4 i_7271047(.A(instrc[97]), .B(n_29667), .C(n_29639), .D(n_30961
		), .Z(n_140088899));
	notech_ao4 i_80570244(.A(n_56888), .B(n_27422), .C(n_27766), .D(n_140088899
		), .Z(n_140188900));
	notech_ao4 i_80470245(.A(n_139788896), .B(n_30524), .C(n_139488893), .D(n_27729
		), .Z(n_140288901));
	notech_ao4 i_80370246(.A(n_56888), .B(n_27424), .C(n_27767), .D(n_140088899
		), .Z(n_140388902));
	notech_ao4 i_80270247(.A(n_139788896), .B(n_30523), .C(n_139488893), .D(n_27730
		), .Z(n_140488903));
	notech_ao4 i_80170248(.A(n_56888), .B(n_27426), .C(n_27768), .D(n_140088899
		), .Z(n_140588904));
	notech_ao4 i_80070249(.A(n_139788896), .B(n_30522), .C(n_139488893), .D(n_27731
		), .Z(n_140688905));
	notech_ao4 i_79970250(.A(n_56888), .B(n_27428), .C(n_27769), .D(n_140088899
		), .Z(n_140788906));
	notech_ao4 i_79870251(.A(n_139788896), .B(n_30521), .C(n_139488893), .D(n_27732
		), .Z(n_140888907));
	notech_ao4 i_79770252(.A(n_56888), .B(n_27430), .C(n_27770), .D(n_140088899
		), .Z(n_140988908));
	notech_ao4 i_79670253(.A(n_139788896), .B(n_30520), .C(n_139488893), .D(n_27733
		), .Z(n_141088909));
	notech_ao4 i_79570254(.A(n_56888), .B(n_27432), .C(n_27771), .D(n_140088899
		), .Z(n_141188910));
	notech_ao4 i_79470255(.A(n_139788896), .B(n_30519), .C(n_139488893), .D(n_27734
		), .Z(n_141288911));
	notech_ao4 i_79370256(.A(n_56888), .B(n_27434), .C(n_27773), .D(n_140088899
		), .Z(n_141388912));
	notech_ao4 i_79270257(.A(n_139788896), .B(n_30518), .C(n_139488893), .D(n_27735
		), .Z(n_141488913));
	notech_ao4 i_79170258(.A(n_56888), .B(n_27437), .C(n_27774), .D(n_140088899
		), .Z(n_141588914));
	notech_ao4 i_79070259(.A(n_139788896), .B(n_30517), .C(n_139488893), .D(n_27737
		), .Z(n_141688915));
	notech_ao4 i_78970260(.A(n_56888), .B(n_27439), .C(n_27775), .D(n_140088899
		), .Z(n_141788916));
	notech_ao4 i_78870261(.A(n_139788896), .B(n_30516), .C(n_139488893), .D(n_27738
		), .Z(n_141888917));
	notech_ao4 i_78770262(.A(n_56888), .B(n_27441), .C(n_27776), .D(n_140088899
		), .Z(n_141988918));
	notech_ao4 i_78670263(.A(n_139788896), .B(n_30515), .C(n_139488893), .D(n_27739
		), .Z(n_142088919));
	notech_ao4 i_78570264(.A(n_56888), .B(n_27443), .C(n_27777), .D(n_140088899
		), .Z(n_142188920));
	notech_ao4 i_78470265(.A(n_139788896), .B(n_30514), .C(n_139488893), .D(n_27740
		), .Z(n_142288921));
	notech_ao4 i_78370266(.A(n_56888), .B(n_27445), .C(n_27779), .D(n_140088899
		), .Z(n_142388922));
	notech_ao4 i_78270267(.A(n_139788896), .B(n_30513), .C(n_139488893), .D(n_27741
		), .Z(n_142488923));
	notech_ao4 i_78170268(.A(n_56888), .B(n_27447), .C(n_27780), .D(n_140088899
		), .Z(n_142588924));
	notech_ao4 i_78070269(.A(n_139788896), .B(n_30512), .C(n_139488893), .D(n_27742
		), .Z(n_142688925));
	notech_ao4 i_77970270(.A(n_56883), .B(n_27449), .C(n_27783), .D(n_140088899
		), .Z(n_142788926));
	notech_ao4 i_77870271(.A(n_139788896), .B(n_30511), .C(n_139488893), .D(n_27743
		), .Z(n_142888927));
	notech_ao4 i_77770272(.A(n_56883), .B(n_27451), .C(n_27785), .D(n_140088899
		), .Z(n_142988928));
	notech_ao4 i_77670273(.A(n_139788896), .B(n_30510), .C(n_139488893), .D(n_27744
		), .Z(n_143088929));
	notech_ao4 i_77570274(.A(n_56883), .B(n_27453), .C(n_27786), .D(n_140088899
		), .Z(n_143188930));
	notech_ao4 i_77470275(.A(n_53680), .B(n_30509), .C(n_53561), .D(n_27745)
		, .Z(n_143288931));
	notech_ao4 i_77370276(.A(n_56883), .B(n_27455), .C(n_27787), .D(n_53691)
		, .Z(n_143388932));
	notech_ao4 i_77270277(.A(n_53680), .B(n_30508), .C(n_53561), .D(n_27747)
		, .Z(n_143488933));
	notech_ao4 i_77170278(.A(n_56883), .B(n_27457), .C(n_27788), .D(n_53691)
		, .Z(n_143588934));
	notech_ao4 i_77070279(.A(n_53680), .B(n_30507), .C(n_53561), .D(n_27748)
		, .Z(n_143688935));
	notech_ao4 i_76970280(.A(n_56883), .B(n_27459), .C(n_27789), .D(n_53691)
		, .Z(n_143788936));
	notech_ao4 i_76870281(.A(n_53680), .B(n_30506), .C(n_53561), .D(n_27749)
		, .Z(n_143888937));
	notech_ao4 i_76770282(.A(n_56883), .B(n_27461), .C(n_27790), .D(n_53691)
		, .Z(n_143988938));
	notech_ao4 i_76670283(.A(n_53680), .B(n_30505), .C(n_53561), .D(n_27750)
		, .Z(n_144088939));
	notech_ao4 i_76570284(.A(n_56883), .B(n_27463), .C(n_27791), .D(n_53691)
		, .Z(n_144188940));
	notech_ao4 i_76470285(.A(n_53680), .B(n_30504), .C(n_53561), .D(n_27751)
		, .Z(n_144288941));
	notech_ao4 i_76370286(.A(n_56883), .B(n_27465), .C(n_27792), .D(n_53691)
		, .Z(n_144388942));
	notech_ao4 i_76270287(.A(n_53680), .B(n_30503), .C(n_53561), .D(n_27752)
		, .Z(n_144488943));
	notech_ao4 i_76170288(.A(n_56883), .B(n_27469), .C(n_27793), .D(n_53691)
		, .Z(n_144588944));
	notech_ao4 i_76070289(.A(n_53680), .B(n_30502), .C(n_53561), .D(n_27755)
		, .Z(n_144688945));
	notech_ao4 i_75970290(.A(n_56883), .B(n_27471), .C(n_27794), .D(n_53691)
		, .Z(n_144788946));
	notech_ao4 i_75870291(.A(n_53680), .B(n_30501), .C(n_53561), .D(n_27756)
		, .Z(n_144888947));
	notech_ao4 i_75770292(.A(n_56883), .B(n_27473), .C(n_27795), .D(n_53691)
		, .Z(n_144988948));
	notech_ao4 i_75670293(.A(n_53680), .B(n_30500), .C(n_53561), .D(n_27758)
		, .Z(n_145088949));
	notech_ao4 i_75570294(.A(n_56883), .B(n_27475), .C(n_27797), .D(n_53691)
		, .Z(n_145188950));
	notech_ao4 i_75470295(.A(n_53680), .B(n_30499), .C(n_139488893), .D(n_27759
		), .Z(n_145288951));
	notech_ao4 i_75370296(.A(n_56883), .B(n_27477), .C(n_27798), .D(n_140088899
		), .Z(n_145388952));
	notech_ao4 i_75270297(.A(n_53680), .B(n_30498), .C(n_53561), .D(n_27760)
		, .Z(n_145488953));
	notech_ao4 i_75170298(.A(n_56883), .B(n_27479), .C(n_27799), .D(n_53691)
		, .Z(n_145588954));
	notech_ao4 i_75070299(.A(n_53680), .B(n_30496), .C(n_53561), .D(n_27762)
		, .Z(n_145688955));
	notech_ao4 i_74970300(.A(n_56883), .B(n_27481), .C(n_27800), .D(n_53691)
		, .Z(n_145788956));
	notech_ao4 i_74870301(.A(n_53680), .B(n_30495), .C(n_53561), .D(n_27763)
		, .Z(n_145888957));
	notech_ao4 i_74770302(.A(n_56883), .B(n_27483), .C(n_27801), .D(n_53691)
		, .Z(n_145988958));
	notech_ao4 i_74670303(.A(n_53680), .B(n_30494), .C(n_53561), .D(n_27764)
		, .Z(n_146088959));
	notech_ao4 i_74570304(.A(n_56883), .B(n_27485), .C(n_27802), .D(n_53691)
		, .Z(n_146188960));
	notech_ao4 i_74470305(.A(n_53680), .B(n_30493), .C(n_53561), .D(n_27765)
		, .Z(n_146288961));
	notech_ao4 i_74370306(.A(n_56883), .B(n_27487), .C(n_27803), .D(n_53691)
		, .Z(n_146388962));
	notech_ao4 i_74270307(.A(n_324090738), .B(n_27766), .C(n_27090), .D(n_27422
		), .Z(n_146488963));
	notech_ao4 i_74170308(.A(n_324290740), .B(n_30492), .C(n_27728), .D(n_324190739
		), .Z(n_146588964));
	notech_ao4 i_74070309(.A(n_324090738), .B(n_27767), .C(n_27090), .D(n_27424
		), .Z(n_146688965));
	notech_ao4 i_73970310(.A(n_324290740), .B(n_30491), .C(n_27729), .D(n_324190739
		), .Z(n_146788966));
	notech_ao4 i_73870311(.A(n_324090738), .B(n_27768), .C(n_27090), .D(n_27426
		), .Z(n_146888967));
	notech_ao4 i_73770312(.A(n_324290740), .B(n_30490), .C(n_27730), .D(n_324190739
		), .Z(n_146988968));
	notech_ao4 i_73670313(.A(n_324090738), .B(n_27769), .C(n_27090), .D(n_27428
		), .Z(n_147088969));
	notech_ao4 i_73570314(.A(n_324290740), .B(n_30489), .C(n_27731), .D(n_324190739
		), .Z(n_147188970));
	notech_ao4 i_73470315(.A(n_324090738), .B(n_27770), .C(n_27090), .D(n_27430
		), .Z(n_147288971));
	notech_ao4 i_73370316(.A(n_324290740), .B(n_30488), .C(n_27732), .D(n_324190739
		), .Z(n_147388972));
	notech_ao4 i_73270317(.A(n_324090738), .B(n_27771), .C(n_27090), .D(n_27432
		), .Z(n_147488973));
	notech_ao4 i_73170318(.A(n_324290740), .B(n_30487), .C(n_27733), .D(n_324190739
		), .Z(n_147588974));
	notech_ao4 i_73070319(.A(n_324090738), .B(n_27773), .C(n_27090), .D(n_27434
		), .Z(n_147688975));
	notech_ao4 i_72970320(.A(n_324290740), .B(n_30486), .C(n_27734), .D(n_324190739
		), .Z(n_147788976));
	notech_ao4 i_72870321(.A(n_324090738), .B(n_27774), .C(n_27090), .D(n_27437
		), .Z(n_147888977));
	notech_ao4 i_72770322(.A(n_324290740), .B(n_30485), .C(n_27735), .D(n_324190739
		), .Z(n_147988978));
	notech_ao4 i_72670323(.A(n_324090738), .B(n_27775), .C(n_27090), .D(n_27439
		), .Z(n_148088979));
	notech_ao4 i_72570324(.A(n_324290740), .B(n_30484), .C(n_27737), .D(n_324190739
		), .Z(n_148188980));
	notech_ao4 i_72470325(.A(n_324090738), .B(n_27776), .C(n_27090), .D(n_27441
		), .Z(n_148288981));
	notech_ao4 i_72370326(.A(n_324290740), .B(n_30483), .C(n_27738), .D(n_324190739
		), .Z(n_148388982));
	notech_ao4 i_72270327(.A(n_324090738), .B(n_27777), .C(n_27090), .D(n_27443
		), .Z(n_148488983));
	notech_ao4 i_72170328(.A(n_324290740), .B(n_30482), .C(n_27739), .D(n_324190739
		), .Z(n_148588984));
	notech_ao4 i_72070329(.A(n_324090738), .B(n_27779), .C(n_27090), .D(n_27445
		), .Z(n_148688985));
	notech_ao4 i_71970330(.A(n_324290740), .B(n_30480), .C(n_27740), .D(n_324190739
		), .Z(n_148788986));
	notech_ao4 i_71870331(.A(n_324090738), .B(n_27780), .C(n_27090), .D(n_27447
		), .Z(n_148888987));
	notech_ao4 i_71770332(.A(n_324290740), .B(n_30479), .C(n_27741), .D(n_324190739
		), .Z(n_148988988));
	notech_ao4 i_71670333(.A(n_324090738), .B(n_27783), .C(n_27090), .D(n_27449
		), .Z(n_149088989));
	notech_ao4 i_71570334(.A(n_324290740), .B(n_30478), .C(n_27742), .D(n_324190739
		), .Z(n_149188990));
	notech_ao4 i_71470335(.A(n_324090738), .B(n_27785), .C(n_27090), .D(n_27451
		), .Z(n_149288991));
	notech_ao4 i_71370336(.A(n_324290740), .B(n_30477), .C(n_27743), .D(n_324190739
		), .Z(n_149388992));
	notech_ao4 i_71270337(.A(n_324090738), .B(n_27786), .C(n_27090), .D(n_27453
		), .Z(n_149488993));
	notech_ao4 i_71170338(.A(n_324290740), .B(n_30476), .C(n_27744), .D(n_324190739
		), .Z(n_149588994));
	notech_ao4 i_71070339(.A(n_53420), .B(n_27787), .C(n_57002), .D(n_27455)
		, .Z(n_149688995));
	notech_ao4 i_70970340(.A(n_53550), .B(n_30474), .C(n_27745), .D(n_53431)
		, .Z(n_149788996));
	notech_ao4 i_70870341(.A(n_53420), .B(n_27788), .C(n_57002), .D(n_27457)
		, .Z(n_149888997));
	notech_ao4 i_70770342(.A(n_53550), .B(n_30473), .C(n_27747), .D(n_53431)
		, .Z(n_149988998));
	notech_ao4 i_70670343(.A(n_53420), .B(n_27789), .C(n_57002), .D(n_27459)
		, .Z(n_150088999));
	notech_ao4 i_70570344(.A(n_53550), .B(n_30471), .C(n_27748), .D(n_53431)
		, .Z(n_150189000));
	notech_ao4 i_70470345(.A(n_53420), .B(n_27790), .C(n_57002), .D(n_27461)
		, .Z(n_150289001));
	notech_ao4 i_70370346(.A(n_53550), .B(n_30469), .C(n_27749), .D(n_53431)
		, .Z(n_150389002));
	notech_ao4 i_70270347(.A(n_53420), .B(n_27791), .C(n_57002), .D(n_27463)
		, .Z(n_150489003));
	notech_ao4 i_70170348(.A(n_53550), .B(n_30468), .C(n_27750), .D(n_53431)
		, .Z(n_150589004));
	notech_ao4 i_70070349(.A(n_53420), .B(n_27792), .C(n_57002), .D(n_27465)
		, .Z(n_150689005));
	notech_ao4 i_69970350(.A(n_53550), .B(n_30467), .C(n_27751), .D(n_53431)
		, .Z(n_150789006));
	notech_ao4 i_69870351(.A(n_53420), .B(n_27793), .C(n_57002), .D(n_27469)
		, .Z(n_150889007));
	notech_ao4 i_69770352(.A(n_53550), .B(n_30465), .C(n_27752), .D(n_53431)
		, .Z(n_150989008));
	notech_ao4 i_69670353(.A(n_53420), .B(n_27794), .C(n_57002), .D(n_27471)
		, .Z(n_151089009));
	notech_ao4 i_69570354(.A(n_53550), .B(n_30463), .C(n_27755), .D(n_53431)
		, .Z(n_151189010));
	notech_ao4 i_69470355(.A(n_53420), .B(n_27795), .C(n_57002), .D(n_27473)
		, .Z(n_151289011));
	notech_ao4 i_69370356(.A(n_53550), .B(n_30462), .C(n_27756), .D(n_53431)
		, .Z(n_151389012));
	notech_ao4 i_69270357(.A(n_53420), .B(n_27797), .C(n_57002), .D(n_27475)
		, .Z(n_151489013));
	notech_ao4 i_69170358(.A(n_53550), .B(n_30460), .C(n_27758), .D(n_53431)
		, .Z(n_151589014));
	notech_ao4 i_69070359(.A(n_53420), .B(n_27798), .C(n_57002), .D(n_27477)
		, .Z(n_151689015));
	notech_ao4 i_68970360(.A(n_53550), .B(n_30458), .C(n_27759), .D(n_324190739
		), .Z(n_151789016));
	notech_ao4 i_68870361(.A(n_53420), .B(n_27799), .C(n_57002), .D(n_27479)
		, .Z(n_151889017));
	notech_ao4 i_68770362(.A(n_53550), .B(n_30457), .C(n_27760), .D(n_53431)
		, .Z(n_151989018));
	notech_ao4 i_68670363(.A(n_27801), .B(n_53420), .C(n_57002), .D(n_27483)
		, .Z(n_152089019));
	notech_ao4 i_68570364(.A(n_53550), .B(n_30456), .C(n_27763), .D(n_53431)
		, .Z(n_152189020));
	notech_ao4 i_68470365(.A(n_53420), .B(n_27802), .C(n_57002), .D(n_27485)
		, .Z(n_152289021));
	notech_ao4 i_68370366(.A(n_53550), .B(n_30454), .C(n_27764), .D(n_53431)
		, .Z(n_152389022));
	notech_ao4 i_68270367(.A(n_53420), .B(n_27803), .C(n_57002), .D(n_27487)
		, .Z(n_152489023));
	notech_ao4 i_68170368(.A(n_53550), .B(n_30453), .C(n_27765), .D(n_53431)
		, .Z(n_152589024));
	notech_nand2 i_6869872(.A(n_3921), .B(n_153089029), .Z(n_152689025));
	notech_or4 i_7569870(.A(instrc[102]), .B(instrc[100]), .C(n_29635), .D(n_29637
		), .Z(n_152789026));
	notech_or4 i_9969854(.A(instrc[101]), .B(n_29665), .C(n_30954), .D(n_29637
		), .Z(n_152889027));
	notech_nand3 i_15469708(.A(n_314890646), .B(instrc[91]), .C(n_166189160)
		, .Z(n_152989028));
	notech_nand3 i_27569587(.A(n_57462), .B(n_308690584), .C(instrc[103]), .Z
		(n_153089029));
	notech_nand2 i_369839(.A(instrc[90]), .B(instrc[89]), .Z(n_166189160));
	notech_or4 i_9069857(.A(from_acu[3]), .B(from_acu[2]), .C(n_29404), .D(from_acu
		[0]), .Z(n_254690045));
	notech_or4 i_8869859(.A(from_acu[3]), .B(from_acu[2]), .C(n_29404), .D(n_29403
		), .Z(n_254890047));
	notech_ao4 i_172268140(.A(n_53118), .B(n_28451), .C(n_53000), .D(n_28289
		), .Z(n_254990048));
	notech_or4 i_830707(.A(from_acu[1]), .B(from_acu[0]), .C(from_acu[3]), .D
		(from_acu[2]), .Z(n_255190050));
	notech_or4 i_8769860(.A(from_acu[1]), .B(from_acu[0]), .C(from_acu[3]), 
		.D(n_27077), .Z(n_255390052));
	notech_or4 i_8669861(.A(from_acu[1]), .B(from_acu[3]), .C(n_29405), .D(n_29403
		), .Z(n_255690055));
	notech_ao4 i_172168141(.A(n_53138), .B(n_28322), .C(n_53128), .D(n_28387
		), .Z(n_255790056));
	notech_or4 i_8569862(.A(n_29405), .B(from_acu[3]), .C(from_acu[0]), .D(n_29404
		), .Z(n_255990058));
	notech_or4 i_8469863(.A(from_acu[3]), .B(from_acu[2]), .C(n_29403), .D(from_acu
		[1]), .Z(n_256090059));
	notech_ao4 i_171968143(.A(n_53158), .B(n_27858), .C(n_53148), .D(n_28560
		), .Z(n_256190060));
	notech_and4 i_6769873(.A(from_acu[2]), .B(from_acu[1]), .C(from_acu[0]),
		 .D(n_29406), .Z(n_256290061));
	notech_ao4 i_171868144(.A(n_53177), .B(n_28483), .C(n_28516), .D(n_53168
		), .Z(n_256390062));
	notech_ao4 i_171668146(.A(n_53118), .B(n_28452), .C(n_53000), .D(n_28290
		), .Z(n_256590064));
	notech_ao4 i_171568147(.A(n_53138), .B(n_28323), .C(n_53128), .D(n_28388
		), .Z(n_256690065));
	notech_ao4 i_171368149(.A(n_53158), .B(n_27859), .C(n_53148), .D(n_28561
		), .Z(n_256890067));
	notech_ao4 i_171268150(.A(n_53177), .B(n_28484), .C(n_28517), .D(n_53168
		), .Z(n_256990068));
	notech_ao4 i_171068152(.A(n_53118), .B(n_28453), .C(n_53000), .D(n_28291
		), .Z(n_257190070));
	notech_ao4 i_170968153(.A(n_53138), .B(n_28324), .C(n_53128), .D(n_28389
		), .Z(n_257290071));
	notech_ao4 i_170768155(.A(n_53158), .B(n_27860), .C(n_53148), .D(n_28562
		), .Z(n_257490073));
	notech_ao4 i_170668156(.A(n_53177), .B(n_28485), .C(n_28518), .D(n_53168
		), .Z(n_257590074));
	notech_ao4 i_170468158(.A(n_53118), .B(n_28454), .C(n_53000), .D(n_28292
		), .Z(n_257790076));
	notech_ao4 i_170368159(.A(n_28325), .B(n_53138), .C(n_53128), .D(n_28390
		), .Z(n_257890077));
	notech_ao4 i_170168161(.A(n_53158), .B(n_27861), .C(n_53148), .D(n_28563
		), .Z(n_258090079));
	notech_ao4 i_170068162(.A(n_53177), .B(n_28486), .C(n_28519), .D(n_53168
		), .Z(n_258190080));
	notech_ao4 i_169868164(.A(n_53117), .B(n_28455), .C(n_52999), .D(n_28293
		), .Z(n_258390082));
	notech_ao4 i_169768165(.A(n_53137), .B(n_28326), .C(n_53127), .D(n_28391
		), .Z(n_258490083));
	notech_ao4 i_169568167(.A(n_53157), .B(n_27862), .C(n_53147), .D(n_28564
		), .Z(n_258690085));
	notech_ao4 i_169468168(.A(n_53176), .B(n_28487), .C(n_28520), .D(n_53167
		), .Z(n_258790086));
	notech_ao4 i_169268170(.A(n_53117), .B(n_28456), .C(n_52999), .D(n_28294
		), .Z(n_258990088));
	notech_ao4 i_169168171(.A(n_53137), .B(n_28327), .C(n_53127), .D(n_28392
		), .Z(n_259090089));
	notech_ao4 i_168968173(.A(n_53157), .B(n_27863), .C(n_53147), .D(n_28565
		), .Z(n_259290091));
	notech_ao4 i_168868174(.A(n_53176), .B(n_28488), .C(n_28521), .D(n_53167
		), .Z(n_259390092));
	notech_ao4 i_168668176(.A(n_53117), .B(n_28457), .C(n_52999), .D(n_28295
		), .Z(n_259590094));
	notech_ao4 i_168568177(.A(n_53137), .B(n_28328), .C(n_53127), .D(n_28393
		), .Z(n_259690095));
	notech_ao4 i_168368179(.A(n_53157), .B(n_27864), .C(n_53147), .D(n_28566
		), .Z(n_259890097));
	notech_ao4 i_168268180(.A(n_53176), .B(n_28489), .C(n_53167), .D(n_28522
		), .Z(n_259990098));
	notech_ao4 i_168068182(.A(n_53117), .B(n_28458), .C(n_52999), .D(n_28296
		), .Z(n_260190100));
	notech_ao4 i_167968183(.A(n_53137), .B(n_28329), .C(n_53127), .D(n_28394
		), .Z(n_260290101));
	notech_ao4 i_167768185(.A(n_53157), .B(n_27865), .C(n_53147), .D(n_28567
		), .Z(n_260490103));
	notech_ao4 i_167668186(.A(n_53176), .B(n_28490), .C(n_28523), .D(n_53167
		), .Z(n_260590104));
	notech_ao4 i_167468188(.A(n_53120), .B(n_28459), .C(n_53001), .D(n_28297
		), .Z(n_260790106));
	notech_ao4 i_167368189(.A(n_53140), .B(n_28330), .C(n_53129), .D(n_28395
		), .Z(n_260890107));
	notech_ao4 i_167168191(.A(n_53160), .B(n_27866), .C(n_53149), .D(n_28568
		), .Z(n_261090109));
	notech_ao4 i_167068192(.A(n_53178), .B(n_28491), .C(n_28525), .D(n_53169
		), .Z(n_261190110));
	notech_ao4 i_166868194(.A(n_53120), .B(n_28460), .C(n_53001), .D(n_28298
		), .Z(n_261390112));
	notech_ao4 i_166768195(.A(n_53140), .B(n_28331), .C(n_53129), .D(n_28396
		), .Z(n_261490113));
	notech_ao4 i_166568197(.A(n_53160), .B(n_27867), .C(n_53149), .D(n_28570
		), .Z(n_261690115));
	notech_ao4 i_166468198(.A(n_53178), .B(n_28492), .C(n_28526), .D(n_53169
		), .Z(n_261790116));
	notech_ao4 i_166268200(.A(n_53120), .B(n_28461), .C(n_53001), .D(n_28299
		), .Z(n_261990118));
	notech_ao4 i_166168201(.A(n_53140), .B(n_28333), .C(n_53129), .D(n_28397
		), .Z(n_262090119));
	notech_ao4 i_165968203(.A(n_53160), .B(n_27868), .C(n_53149), .D(n_28571
		), .Z(n_262290121));
	notech_ao4 i_165868204(.A(n_53178), .B(n_28493), .C(n_53169), .D(n_28528
		), .Z(n_262390122));
	notech_ao4 i_165668206(.A(n_53120), .B(n_28462), .C(n_53001), .D(n_28301
		), .Z(n_262590124));
	notech_ao4 i_165568207(.A(n_53140), .B(n_28334), .C(n_53129), .D(n_28398
		), .Z(n_262690125));
	notech_ao4 i_165368209(.A(n_53160), .B(n_27869), .C(n_53149), .D(n_28572
		), .Z(n_262890127));
	notech_ao4 i_165268210(.A(n_53178), .B(n_28494), .C(n_53169), .D(n_28529
		), .Z(n_262990128));
	notech_ao4 i_165068212(.A(n_53119), .B(n_28463), .C(n_53000), .D(n_28302
		), .Z(n_263190130));
	notech_ao4 i_164968213(.A(n_53139), .B(n_28335), .C(n_53128), .D(n_28399
		), .Z(n_263290131));
	notech_ao4 i_164768215(.A(n_53159), .B(n_27870), .C(n_53148), .D(n_28573
		), .Z(n_263490133));
	notech_ao4 i_164668216(.A(n_53177), .B(n_28495), .C(n_28531), .D(n_53168
		), .Z(n_263590134));
	notech_ao4 i_164468218(.A(n_53119), .B(n_28464), .C(n_53000), .D(n_28303
		), .Z(n_263790136));
	notech_ao4 i_164368219(.A(n_53139), .B(n_28336), .C(n_53128), .D(n_28400
		), .Z(n_263890137));
	notech_ao4 i_164168221(.A(n_53159), .B(n_27871), .C(n_53148), .D(n_28574
		), .Z(n_264090139));
	notech_ao4 i_164068222(.A(n_53177), .B(n_28496), .C(n_53168), .D(n_28534
		), .Z(n_264190140));
	notech_ao4 i_163868224(.A(n_53119), .B(n_28465), .C(n_53001), .D(n_28304
		), .Z(n_264390142));
	notech_ao4 i_163768225(.A(n_53139), .B(n_28337), .C(n_53129), .D(n_28401
		), .Z(n_264490143));
	notech_ao4 i_163568227(.A(n_53159), .B(n_27872), .C(n_53149), .D(n_28575
		), .Z(n_264690145));
	notech_ao4 i_163468228(.A(n_53178), .B(n_28497), .C(n_53169), .D(n_28535
		), .Z(n_264790146));
	notech_ao4 i_163268230(.A(n_53119), .B(n_28466), .C(n_53001), .D(n_28305
		), .Z(n_264990148));
	notech_ao4 i_163168231(.A(n_53139), .B(n_28338), .C(n_53129), .D(n_28402
		), .Z(n_265090149));
	notech_ao4 i_162968233(.A(n_53159), .B(n_27873), .C(n_53149), .D(n_28576
		), .Z(n_265290151));
	notech_ao4 i_162868234(.A(n_53178), .B(n_28498), .C(n_28536), .D(n_53169
		), .Z(n_265390152));
	notech_ao4 i_162668236(.A(n_53113), .B(n_28467), .C(n_52996), .D(n_28306
		), .Z(n_265590154));
	notech_ao4 i_162568237(.A(n_53133), .B(n_28339), .C(n_53124), .D(n_28403
		), .Z(n_265690155));
	notech_ao4 i_162368239(.A(n_53153), .B(n_27874), .C(n_53144), .D(n_28577
		), .Z(n_265890157));
	notech_ao4 i_162268240(.A(n_53176), .B(n_28499), .C(n_28537), .D(n_53164
		), .Z(n_265990158));
	notech_ao4 i_162068242(.A(n_53113), .B(n_28468), .C(n_52995), .D(n_28307
		), .Z(n_266190160));
	notech_ao4 i_161968243(.A(n_53133), .B(n_28340), .C(n_53123), .D(n_28404
		), .Z(n_266290161));
	notech_ao4 i_161768245(.A(n_53153), .B(n_27875), .C(n_53143), .D(n_28578
		), .Z(n_266490163));
	notech_ao4 i_161668246(.A(n_53173), .B(n_28500), .C(n_28538), .D(n_53163
		), .Z(n_266590164));
	notech_ao4 i_161468248(.A(n_53113), .B(n_28469), .C(n_52996), .D(n_28308
		), .Z(n_266790166));
	notech_ao4 i_161368249(.A(n_53133), .B(n_28341), .C(n_53124), .D(n_28405
		), .Z(n_266890167));
	notech_ao4 i_161168251(.A(n_53153), .B(n_27876), .C(n_53144), .D(n_28579
		), .Z(n_267090169));
	notech_ao4 i_161068252(.A(n_53172), .B(n_28501), .C(n_28539), .D(n_53164
		), .Z(n_267190170));
	notech_ao4 i_160868254(.A(n_53113), .B(n_28470), .C(n_52996), .D(n_28309
		), .Z(n_267390172));
	notech_ao4 i_160768255(.A(n_53133), .B(n_28342), .C(n_53124), .D(n_28406
		), .Z(n_267490173));
	notech_ao4 i_160568257(.A(n_53153), .B(n_27878), .C(n_53144), .D(n_28580
		), .Z(n_267690175));
	notech_ao4 i_160468258(.A(n_53173), .B(n_28503), .C(n_28540), .D(n_53164
		), .Z(n_267790176));
	notech_ao4 i_160268260(.A(n_53112), .B(n_28471), .C(n_52995), .D(n_28310
		), .Z(n_267990178));
	notech_ao4 i_160168261(.A(n_53132), .B(n_28343), .C(n_53123), .D(n_28407
		), .Z(n_268090179));
	notech_ao4 i_159968263(.A(n_53152), .B(n_27881), .C(n_53143), .D(n_28581
		), .Z(n_268290181));
	notech_ao4 i_159868264(.A(n_53173), .B(n_28504), .C(n_28541), .D(n_53163
		), .Z(n_268390182));
	notech_ao4 i_159668266(.A(n_53112), .B(n_28472), .C(n_52995), .D(n_28311
		), .Z(n_268590184));
	notech_ao4 i_159568267(.A(n_53132), .B(n_28344), .C(n_53123), .D(n_28408
		), .Z(n_268690185));
	notech_ao4 i_159368269(.A(n_53152), .B(n_27882), .C(n_53143), .D(n_28582
		), .Z(n_268890187));
	notech_ao4 i_159268270(.A(n_53172), .B(n_28505), .C(n_53163), .D(n_28547
		), .Z(n_268990188));
	notech_ao4 i_159068272(.A(n_53112), .B(n_28473), .C(n_52995), .D(n_28312
		), .Z(n_269190190));
	notech_ao4 i_158968273(.A(n_53132), .B(n_28345), .C(n_53123), .D(n_28409
		), .Z(n_269290191));
	notech_ao4 i_158768275(.A(n_53152), .B(n_27883), .C(n_53143), .D(n_28583
		), .Z(n_269490193));
	notech_ao4 i_158668276(.A(n_53172), .B(n_28506), .C(n_28548), .D(n_53163
		), .Z(n_269590194));
	notech_ao4 i_158468278(.A(n_53112), .B(n_28474), .C(n_52995), .D(n_28313
		), .Z(n_269790196));
	notech_ao4 i_158368279(.A(n_53132), .B(n_28346), .C(n_53123), .D(n_28410
		), .Z(n_269890197));
	notech_ao4 i_158168281(.A(n_53152), .B(n_27884), .C(n_53143), .D(n_28584
		), .Z(n_270090199));
	notech_ao4 i_158068282(.A(n_53172), .B(n_28507), .C(n_28549), .D(n_53163
		), .Z(n_270190200));
	notech_ao4 i_157868284(.A(n_53115), .B(n_28475), .C(n_52997), .D(n_28314
		), .Z(n_270390202));
	notech_ao4 i_157768285(.A(n_53135), .B(n_28347), .C(n_53125), .D(n_28411
		), .Z(n_270490203));
	notech_ao4 i_157568287(.A(n_53155), .B(n_27886), .C(n_53145), .D(n_28585
		), .Z(n_270690205));
	notech_ao4 i_157468288(.A(n_53172), .B(n_28508), .C(n_28550), .D(n_53165
		), .Z(n_270790206));
	notech_ao4 i_157268290(.A(n_53115), .B(n_28476), .C(n_52997), .D(n_28315
		), .Z(n_270990208));
	notech_ao4 i_157168291(.A(n_53135), .B(n_28348), .C(n_53125), .D(n_28412
		), .Z(n_271090209));
	notech_ao4 i_156968293(.A(n_53155), .B(n_27887), .C(n_53145), .D(n_28586
		), .Z(n_271290211));
	notech_ao4 i_156868294(.A(n_53174), .B(n_28509), .C(n_28553), .D(n_53165
		), .Z(n_271390212));
	notech_ao4 i_156668296(.A(n_53115), .B(n_28477), .C(n_52999), .D(n_28316
		), .Z(n_271590214));
	notech_ao4 i_156568297(.A(n_53135), .B(n_28349), .C(n_53127), .D(n_28413
		), .Z(n_271690215));
	notech_ao4 i_156368299(.A(n_53155), .B(n_27888), .C(n_53147), .D(n_28587
		), .Z(n_271890217));
	notech_ao4 i_156268300(.A(n_53174), .B(n_28510), .C(n_28554), .D(n_53167
		), .Z(n_271990218));
	notech_ao4 i_156068302(.A(n_53115), .B(n_28478), .C(n_52997), .D(n_28317
		), .Z(n_272190220));
	notech_ao4 i_155968303(.A(n_53135), .B(n_28350), .C(n_53125), .D(n_28414
		), .Z(n_272290221));
	notech_ao4 i_155768305(.A(n_53155), .B(n_27889), .C(n_53145), .D(n_28588
		), .Z(n_272490223));
	notech_ao4 i_155668306(.A(n_53176), .B(n_28511), .C(n_28555), .D(n_53165
		), .Z(n_272590224));
	notech_ao4 i_155468308(.A(n_53114), .B(n_28479), .C(n_52996), .D(n_28318
		), .Z(n_272790226));
	notech_ao4 i_155368309(.A(n_53134), .B(n_28351), .C(n_53124), .D(n_28415
		), .Z(n_272890227));
	notech_ao4 i_155168311(.A(n_53154), .B(n_27890), .C(n_53144), .D(n_28589
		), .Z(n_273090229));
	notech_ao4 i_155068312(.A(n_53174), .B(n_28512), .C(n_28556), .D(n_53164
		), .Z(n_273190230));
	notech_ao4 i_154868314(.A(n_53114), .B(n_28480), .C(n_52996), .D(n_28319
		), .Z(n_273390232));
	notech_ao4 i_154768315(.A(n_53134), .B(n_28352), .C(n_53124), .D(n_28416
		), .Z(n_273490233));
	notech_ao4 i_154568317(.A(n_53154), .B(n_27891), .C(n_53144), .D(n_28590
		), .Z(n_273690235));
	notech_ao4 i_154468318(.A(n_53173), .B(n_28513), .C(n_28557), .D(n_53164
		), .Z(n_273790236));
	notech_ao4 i_154268320(.A(n_53114), .B(n_28481), .C(n_52997), .D(n_28320
		), .Z(n_273990238));
	notech_ao4 i_154168321(.A(n_53134), .B(n_28353), .C(n_53125), .D(n_28417
		), .Z(n_274090239));
	notech_ao4 i_153968323(.A(n_53154), .B(n_27892), .C(n_53145), .D(n_28591
		), .Z(n_274290241));
	notech_ao4 i_153868324(.A(n_53173), .B(n_28514), .C(n_28558), .D(n_53165
		), .Z(n_274390242));
	notech_ao4 i_153668326(.A(n_53114), .B(n_28482), .C(n_52997), .D(n_28321
		), .Z(n_274590244));
	notech_ao4 i_153568327(.A(n_53134), .B(n_28354), .C(n_53125), .D(n_28418
		), .Z(n_274690245));
	notech_ao4 i_153368329(.A(n_53154), .B(n_27893), .C(n_53145), .D(n_28592
		), .Z(n_274890247));
	notech_ao4 i_153268330(.A(n_53174), .B(n_28515), .C(n_28559), .D(n_53165
		), .Z(n_274990248));
	notech_or4 i_9769855(.A(from_acu[7]), .B(n_29409), .C(n_29408), .D(n_29407
		), .Z(n_275390252));
	notech_or4 i_8369864(.A(from_acu[7]), .B(from_acu[6]), .C(n_29407), .D(from_acu
		[5]), .Z(n_275690255));
	notech_ao4 i_152968333(.A(n_53196), .B(n_27858), .C(n_28516), .D(n_53186
		), .Z(n_275790256));
	notech_or4 i_8269865(.A(from_acu[7]), .B(from_acu[6]), .C(n_29408), .D(from_acu
		[4]), .Z(n_275990258));
	notech_or4 i_8169866(.A(from_acu[7]), .B(from_acu[6]), .C(n_29408), .D(n_29407
		), .Z(n_276090259));
	notech_ao4 i_152868334(.A(n_53216), .B(n_28451), .C(n_53206), .D(n_28289
		), .Z(n_276190260));
	notech_or4 i_830731(.A(from_acu[7]), .B(from_acu[5]), .C(from_acu[4]), .D
		(from_acu[6]), .Z(n_276490263));
	notech_or4 i_7969867(.A(from_acu[5]), .B(from_acu[4]), .C(from_acu[7]), 
		.D(n_27081), .Z(n_276690265));
	notech_or4 i_7769868(.A(from_acu[7]), .B(n_29409), .C(n_29407), .D(from_acu
		[5]), .Z(n_276790266));
	notech_ao4 i_152668336(.A(n_53236), .B(n_28322), .C(n_53226), .D(n_28387
		), .Z(n_276890267));
	notech_or4 i_7669869(.A(from_acu[4]), .B(from_acu[7]), .C(n_29408), .D(n_29409
		), .Z(n_276990268));
	notech_ao4 i_152568337(.A(n_53255), .B(n_28483), .C(n_28560), .D(n_53246
		), .Z(n_277090269));
	notech_ao4 i_152368339(.A(n_53196), .B(n_27859), .C(n_28517), .D(n_53186
		), .Z(n_277290271));
	notech_ao4 i_152268340(.A(n_53216), .B(n_28452), .C(n_53206), .D(n_28290
		), .Z(n_277390272));
	notech_ao4 i_152068342(.A(n_53236), .B(n_28323), .C(n_53226), .D(n_28388
		), .Z(n_277590274));
	notech_ao4 i_151968343(.A(n_53255), .B(n_28484), .C(n_53246), .D(n_28561
		), .Z(n_277690275));
	notech_ao4 i_151768345(.A(n_53196), .B(n_27860), .C(n_28518), .D(n_53186
		), .Z(n_277890277));
	notech_ao4 i_151668346(.A(n_28453), .B(n_53216), .C(n_53206), .D(n_28291
		), .Z(n_277990278));
	notech_ao4 i_151468348(.A(n_53236), .B(n_28324), .C(n_53226), .D(n_28389
		), .Z(n_278190280));
	notech_ao4 i_151368349(.A(n_53255), .B(n_28485), .C(n_53246), .D(n_28562
		), .Z(n_278290281));
	notech_ao4 i_151168351(.A(n_53196), .B(n_27861), .C(n_28519), .D(n_53186
		), .Z(n_278490283));
	notech_ao4 i_151068352(.A(n_53216), .B(n_28454), .C(n_53206), .D(n_28292
		), .Z(n_278590284));
	notech_ao4 i_150868354(.A(n_28325), .B(n_53236), .C(n_53226), .D(n_28390
		), .Z(n_278790286));
	notech_ao4 i_150768355(.A(n_53255), .B(n_28486), .C(n_53246), .D(n_28563
		), .Z(n_278890287));
	notech_ao4 i_150568357(.A(n_53195), .B(n_27862), .C(n_53185), .D(n_28520
		), .Z(n_279090289));
	notech_ao4 i_150468358(.A(n_53215), .B(n_28455), .C(n_53205), .D(n_28293
		), .Z(n_279190290));
	notech_ao4 i_150268360(.A(n_53235), .B(n_28326), .C(n_53225), .D(n_28391
		), .Z(n_279390292));
	notech_ao4 i_150168361(.A(n_53254), .B(n_28487), .C(n_53245), .D(n_28564
		), .Z(n_279490293));
	notech_ao4 i_149968363(.A(n_53195), .B(n_27863), .C(n_28521), .D(n_53185
		), .Z(n_279690295));
	notech_ao4 i_149868364(.A(n_53215), .B(n_28456), .C(n_53205), .D(n_28294
		), .Z(n_279790296));
	notech_ao4 i_149668366(.A(n_53235), .B(n_28327), .C(n_53225), .D(n_28392
		), .Z(n_279990298));
	notech_ao4 i_149568367(.A(n_53254), .B(n_28488), .C(n_53245), .D(n_28565
		), .Z(n_280090299));
	notech_ao4 i_149368369(.A(n_53195), .B(n_27864), .C(n_28522), .D(n_53185
		), .Z(n_280290301));
	notech_ao4 i_149268370(.A(n_53215), .B(n_28457), .C(n_53205), .D(n_28295
		), .Z(n_280390302));
	notech_ao4 i_149068372(.A(n_53235), .B(n_28328), .C(n_53225), .D(n_28393
		), .Z(n_280590304));
	notech_ao4 i_148968373(.A(n_53254), .B(n_28489), .C(n_53245), .D(n_28566
		), .Z(n_280690305));
	notech_ao4 i_148768375(.A(n_53195), .B(n_27865), .C(n_28523), .D(n_53185
		), .Z(n_280890307));
	notech_ao4 i_148668376(.A(n_53215), .B(n_28458), .C(n_53205), .D(n_28296
		), .Z(n_280990308));
	notech_ao4 i_148468378(.A(n_53235), .B(n_28329), .C(n_53225), .D(n_28394
		), .Z(n_281190310));
	notech_ao4 i_148368379(.A(n_53254), .B(n_28490), .C(n_53245), .D(n_28567
		), .Z(n_281290311));
	notech_ao4 i_148168381(.A(n_53198), .B(n_27866), .C(n_28525), .D(n_53187
		), .Z(n_281490313));
	notech_ao4 i_148068382(.A(n_53218), .B(n_28459), .C(n_53207), .D(n_28297
		), .Z(n_281590314));
	notech_ao4 i_147868384(.A(n_53238), .B(n_28330), .C(n_53227), .D(n_28395
		), .Z(n_281790316));
	notech_ao4 i_147768385(.A(n_53256), .B(n_28491), .C(n_53247), .D(n_28568
		), .Z(n_281890317));
	notech_ao4 i_147568387(.A(n_53198), .B(n_27867), .C(n_53187), .D(n_28526
		), .Z(n_282090319));
	notech_ao4 i_147468388(.A(n_53218), .B(n_28460), .C(n_53207), .D(n_28298
		), .Z(n_282190320));
	notech_ao4 i_147268390(.A(n_53238), .B(n_28331), .C(n_53227), .D(n_28396
		), .Z(n_282390322));
	notech_ao4 i_147168391(.A(n_53256), .B(n_28492), .C(n_53247), .D(n_28570
		), .Z(n_282490323));
	notech_ao4 i_146968393(.A(n_53198), .B(n_27868), .C(n_28528), .D(n_53187
		), .Z(n_282690325));
	notech_ao4 i_146868394(.A(n_53218), .B(n_28461), .C(n_53207), .D(n_28299
		), .Z(n_282790326));
	notech_ao4 i_146668396(.A(n_53238), .B(n_28333), .C(n_53227), .D(n_28397
		), .Z(n_282990328));
	notech_ao4 i_146568397(.A(n_53256), .B(n_28493), .C(n_53247), .D(n_28571
		), .Z(n_283090329));
	notech_ao4 i_146368399(.A(n_53198), .B(n_27869), .C(n_28529), .D(n_53187
		), .Z(n_283290331));
	notech_ao4 i_146268400(.A(n_53218), .B(n_28462), .C(n_53207), .D(n_28301
		), .Z(n_283390332));
	notech_ao4 i_146068402(.A(n_53238), .B(n_28334), .C(n_53227), .D(n_28398
		), .Z(n_283590334));
	notech_ao4 i_145968403(.A(n_53256), .B(n_28494), .C(n_53247), .D(n_28572
		), .Z(n_283690335));
	notech_ao4 i_145768405(.A(n_53197), .B(n_27870), .C(n_53186), .D(n_28531
		), .Z(n_283890337));
	notech_ao4 i_145668406(.A(n_53217), .B(n_28463), .C(n_53206), .D(n_28302
		), .Z(n_283990338));
	notech_ao4 i_145468408(.A(n_53237), .B(n_28335), .C(n_53226), .D(n_28399
		), .Z(n_284190340));
	notech_ao4 i_145368409(.A(n_53255), .B(n_28495), .C(n_53246), .D(n_28573
		), .Z(n_284290341));
	notech_ao4 i_145168411(.A(n_53197), .B(n_27871), .C(n_28534), .D(n_53186
		), .Z(n_284490343));
	notech_ao4 i_145068412(.A(n_53217), .B(n_28464), .C(n_53206), .D(n_28303
		), .Z(n_284590344));
	notech_ao4 i_144868414(.A(n_53237), .B(n_28336), .C(n_53226), .D(n_28400
		), .Z(n_284790346));
	notech_ao4 i_144768415(.A(n_53255), .B(n_28496), .C(n_53246), .D(n_28574
		), .Z(n_284890347));
	notech_ao4 i_144568417(.A(n_53197), .B(n_27872), .C(n_28535), .D(n_53187
		), .Z(n_285090349));
	notech_ao4 i_144468418(.A(n_53217), .B(n_28465), .C(n_53207), .D(n_28304
		), .Z(n_285190350));
	notech_ao4 i_144268420(.A(n_53237), .B(n_28337), .C(n_53227), .D(n_28401
		), .Z(n_285390352));
	notech_ao4 i_144168421(.A(n_53256), .B(n_28497), .C(n_53247), .D(n_28575
		), .Z(n_285490353));
	notech_ao4 i_143968423(.A(n_53197), .B(n_27873), .C(n_28536), .D(n_53187
		), .Z(n_285690355));
	notech_ao4 i_143868424(.A(n_53217), .B(n_28466), .C(n_53207), .D(n_28305
		), .Z(n_285790356));
	notech_ao4 i_143668426(.A(n_53237), .B(n_28338), .C(n_53227), .D(n_28402
		), .Z(n_285990358));
	notech_ao4 i_143568427(.A(n_53256), .B(n_28498), .C(n_53247), .D(n_28576
		), .Z(n_286090359));
	notech_ao4 i_143368429(.A(n_53191), .B(n_27874), .C(n_28537), .D(n_53182
		), .Z(n_286290361));
	notech_ao4 i_143268430(.A(n_53211), .B(n_28467), .C(n_53202), .D(n_28306
		), .Z(n_286390362));
	notech_ao4 i_143068432(.A(n_53231), .B(n_28339), .C(n_53222), .D(n_28403
		), .Z(n_286590364));
	notech_ao4 i_142968433(.A(n_53254), .B(n_28499), .C(n_53242), .D(n_28577
		), .Z(n_286690365));
	notech_ao4 i_142768435(.A(n_53191), .B(n_27875), .C(n_28538), .D(n_53181
		), .Z(n_286890367));
	notech_ao4 i_142668436(.A(n_53211), .B(n_28468), .C(n_53201), .D(n_28307
		), .Z(n_286990368));
	notech_ao4 i_142468438(.A(n_53231), .B(n_28340), .C(n_53221), .D(n_28404
		), .Z(n_287190370));
	notech_ao4 i_142368439(.A(n_53251), .B(n_28500), .C(n_53241), .D(n_28578
		), .Z(n_287290371));
	notech_ao4 i_142168441(.A(n_53191), .B(n_27876), .C(n_28539), .D(n_53182
		), .Z(n_287490373));
	notech_ao4 i_142068442(.A(n_53211), .B(n_28469), .C(n_53202), .D(n_28308
		), .Z(n_287590374));
	notech_ao4 i_141868444(.A(n_53231), .B(n_28341), .C(n_53222), .D(n_28405
		), .Z(n_287790376));
	notech_ao4 i_141768445(.A(n_53250), .B(n_28501), .C(n_53242), .D(n_28579
		), .Z(n_287890377));
	notech_ao4 i_141568447(.A(n_53191), .B(n_27878), .C(n_28540), .D(n_53182
		), .Z(n_288090379));
	notech_ao4 i_141468448(.A(n_53211), .B(n_28470), .C(n_53202), .D(n_28309
		), .Z(n_288190380));
	notech_ao4 i_141268450(.A(n_53231), .B(n_28342), .C(n_53222), .D(n_28406
		), .Z(n_288390382));
	notech_ao4 i_141168451(.A(n_53251), .B(n_28503), .C(n_53242), .D(n_28580
		), .Z(n_288490383));
	notech_ao4 i_140968453(.A(n_53190), .B(n_27881), .C(n_28541), .D(n_53181
		), .Z(n_288690385));
	notech_ao4 i_140868454(.A(n_53210), .B(n_28471), .C(n_53201), .D(n_28310
		), .Z(n_288790386));
	notech_ao4 i_140668456(.A(n_53230), .B(n_28343), .C(n_53221), .D(n_28407
		), .Z(n_288990388));
	notech_ao4 i_140568457(.A(n_53251), .B(n_28504), .C(n_53241), .D(n_28581
		), .Z(n_289090389));
	notech_ao4 i_140368459(.A(n_53190), .B(n_27882), .C(n_28547), .D(n_53181
		), .Z(n_289290391));
	notech_ao4 i_140268460(.A(n_53210), .B(n_28472), .C(n_53201), .D(n_28311
		), .Z(n_289390392));
	notech_ao4 i_140068462(.A(n_53230), .B(n_28344), .C(n_53221), .D(n_28408
		), .Z(n_289590394));
	notech_ao4 i_139968463(.A(n_53250), .B(n_28505), .C(n_53241), .D(n_28582
		), .Z(n_289690395));
	notech_ao4 i_139768465(.A(n_53190), .B(n_27883), .C(n_28548), .D(n_53181
		), .Z(n_289890397));
	notech_ao4 i_139668466(.A(n_53210), .B(n_28473), .C(n_53201), .D(n_28312
		), .Z(n_289990398));
	notech_ao4 i_139468468(.A(n_53230), .B(n_28345), .C(n_53221), .D(n_28409
		), .Z(n_290190400));
	notech_ao4 i_139368469(.A(n_53250), .B(n_28506), .C(n_53241), .D(n_28583
		), .Z(n_290290401));
	notech_ao4 i_139168471(.A(n_53190), .B(n_27884), .C(n_28549), .D(n_53181
		), .Z(n_290490403));
	notech_ao4 i_139068472(.A(n_53210), .B(n_28474), .C(n_53201), .D(n_28313
		), .Z(n_290590404));
	notech_ao4 i_138868474(.A(n_53230), .B(n_28346), .C(n_53221), .D(n_28410
		), .Z(n_290790406));
	notech_ao4 i_138768475(.A(n_53250), .B(n_28507), .C(n_53241), .D(n_28584
		), .Z(n_290890407));
	notech_ao4 i_138568477(.A(n_53193), .B(n_27886), .C(n_28550), .D(n_53183
		), .Z(n_291090409));
	notech_ao4 i_138468478(.A(n_53213), .B(n_28475), .C(n_53203), .D(n_28314
		), .Z(n_291190410));
	notech_ao4 i_138268480(.A(n_53233), .B(n_28347), .C(n_53223), .D(n_28411
		), .Z(n_291390412));
	notech_ao4 i_138168481(.A(n_53250), .B(n_28508), .C(n_53243), .D(n_28585
		), .Z(n_291490413));
	notech_ao4 i_137968483(.A(n_53193), .B(n_27887), .C(n_28553), .D(n_53183
		), .Z(n_291690415));
	notech_ao4 i_137868484(.A(n_53213), .B(n_28476), .C(n_53203), .D(n_28315
		), .Z(n_291790416));
	notech_ao4 i_137668486(.A(n_53233), .B(n_28348), .C(n_53223), .D(n_28412
		), .Z(n_291990418));
	notech_ao4 i_137568487(.A(n_53252), .B(n_28509), .C(n_53243), .D(n_28586
		), .Z(n_292090419));
	notech_ao4 i_137368489(.A(n_53193), .B(n_27888), .C(n_28554), .D(n_53185
		), .Z(n_292290421));
	notech_ao4 i_137268490(.A(n_53213), .B(n_28477), .C(n_53205), .D(n_28316
		), .Z(n_292390422));
	notech_ao4 i_137068492(.A(n_53233), .B(n_28349), .C(n_53225), .D(n_28413
		), .Z(n_292590424));
	notech_ao4 i_136968493(.A(n_53252), .B(n_28510), .C(n_53245), .D(n_28587
		), .Z(n_292690425));
	notech_ao4 i_136768495(.A(n_53193), .B(n_27889), .C(n_28555), .D(n_53183
		), .Z(n_292890427));
	notech_ao4 i_136668496(.A(n_53213), .B(n_28478), .C(n_53203), .D(n_28317
		), .Z(n_292990428));
	notech_ao4 i_136468498(.A(n_53233), .B(n_28350), .C(n_53223), .D(n_28414
		), .Z(n_293190430));
	notech_ao4 i_136368499(.A(n_53254), .B(n_28511), .C(n_53243), .D(n_28588
		), .Z(n_293290431));
	notech_ao4 i_136168501(.A(n_53192), .B(n_27890), .C(n_28556), .D(n_53182
		), .Z(n_293490433));
	notech_ao4 i_136068502(.A(n_53212), .B(n_28479), .C(n_53202), .D(n_28318
		), .Z(n_293590434));
	notech_ao4 i_135868504(.A(n_53232), .B(n_28351), .C(n_53222), .D(n_28415
		), .Z(n_293790436));
	notech_ao4 i_135768505(.A(n_53252), .B(n_28512), .C(n_53242), .D(n_28589
		), .Z(n_293890437));
	notech_ao4 i_135568507(.A(n_53192), .B(n_27891), .C(n_28557), .D(n_53182
		), .Z(n_294090439));
	notech_ao4 i_135468508(.A(n_53212), .B(n_28480), .C(n_53202), .D(n_28319
		), .Z(n_294190440));
	notech_ao4 i_135268510(.A(n_53232), .B(n_28352), .C(n_53222), .D(n_28416
		), .Z(n_294390442));
	notech_ao4 i_135168511(.A(n_53251), .B(n_28513), .C(n_53242), .D(n_28590
		), .Z(n_294490443));
	notech_ao4 i_134968513(.A(n_53192), .B(n_27892), .C(n_28558), .D(n_53183
		), .Z(n_294690445));
	notech_ao4 i_134868514(.A(n_53212), .B(n_28481), .C(n_53203), .D(n_28320
		), .Z(n_294790446));
	notech_ao4 i_134668516(.A(n_53232), .B(n_28353), .C(n_53223), .D(n_28417
		), .Z(n_294990448));
	notech_ao4 i_134568517(.A(n_53251), .B(n_28514), .C(n_53243), .D(n_28591
		), .Z(n_295090449));
	notech_ao4 i_134368519(.A(n_53192), .B(n_27893), .C(n_28559), .D(n_53183
		), .Z(n_295290451));
	notech_ao4 i_134268520(.A(n_53212), .B(n_28482), .C(n_53203), .D(n_28321
		), .Z(n_295390452));
	notech_ao4 i_134068522(.A(n_53232), .B(n_28354), .C(n_53223), .D(n_28418
		), .Z(n_295590454));
	notech_ao4 i_133968523(.A(n_53252), .B(n_28515), .C(n_53243), .D(n_28592
		), .Z(n_295690455));
	notech_ao4 i_133868524(.A(n_326990767), .B(n_56046), .C(n_56380), .D(n_27422
		), .Z(n_295890457));
	notech_ao4 i_133768525(.A(n_326790765), .B(n_27728), .C(n_326890766), .D
		(n_27766), .Z(n_295990458));
	notech_ao4 i_133668526(.A(n_60024), .B(n_326990767), .C(n_56380), .D(n_27424
		), .Z(n_296090459));
	notech_ao4 i_133568527(.A(n_326790765), .B(n_27729), .C(n_326890766), .D
		(n_27767), .Z(n_296190460));
	notech_ao4 i_133268530(.A(n_326990767), .B(n_60022), .C(n_56380), .D(n_27428
		), .Z(n_296290461));
	notech_ao4 i_133168531(.A(n_326790765), .B(n_27731), .C(n_326890766), .D
		(n_27769), .Z(n_296390462));
	notech_ao4 i_133068532(.A(n_5743), .B(n_326990767), .C(n_56380), .D(n_27430
		), .Z(n_296490463));
	notech_ao4 i_132968533(.A(n_326790765), .B(n_27732), .C(n_326890766), .D
		(n_27770), .Z(n_296590464));
	notech_ao4 i_132868534(.A(n_326990767), .B(n_60020), .C(n_56380), .D(n_27432
		), .Z(n_296690465));
	notech_ao4 i_132768535(.A(n_326790765), .B(n_27733), .C(n_326890766), .D
		(n_27771), .Z(n_296790466));
	notech_ao4 i_132668536(.A(n_326990767), .B(n_3874), .C(n_56385), .D(n_27434
		), .Z(n_296890467));
	notech_ao4 i_132568537(.A(n_326790765), .B(n_27734), .C(n_326890766), .D
		(n_27773), .Z(n_296990468));
	notech_ao4 i_132468538(.A(n_303191792), .B(n_326990767), .C(n_56380), .D
		(n_27437), .Z(n_297090469));
	notech_ao4 i_132368539(.A(n_326790765), .B(n_27735), .C(n_326890766), .D
		(n_27774), .Z(n_297190470));
	notech_ao4 i_132268540(.A(n_326990767), .B(n_5933), .C(n_56380), .D(n_27439
		), .Z(n_297290471));
	notech_ao4 i_132168541(.A(n_326790765), .B(n_27737), .C(n_326890766), .D
		(n_27775), .Z(n_297390472));
	notech_ao4 i_132068542(.A(n_326990767), .B(n_60016), .C(n_56380), .D(n_27441
		), .Z(n_297490473));
	notech_ao4 i_131968543(.A(n_326790765), .B(n_27738), .C(n_326890766), .D
		(n_27776), .Z(n_297590474));
	notech_ao4 i_131868544(.A(n_3850), .B(n_54062), .C(n_56380), .D(n_27443)
		, .Z(n_297690475));
	notech_ao4 i_131768545(.A(n_54082), .B(n_27739), .C(n_54073), .D(n_27777
		), .Z(n_297790476));
	notech_ao4 i_131668546(.A(n_54062), .B(n_302491799), .C(n_56380), .D(n_27445
		), .Z(n_297890477));
	notech_ao4 i_131568547(.A(n_54082), .B(n_27740), .C(n_54073), .D(n_27779
		), .Z(n_297990478));
	notech_ao4 i_131268550(.A(n_54062), .B(n_302091803), .C(n_56380), .D(n_27449
		), .Z(n_298090479));
	notech_ao4 i_131168551(.A(n_54082), .B(n_27742), .C(n_54073), .D(n_27783
		), .Z(n_298190480));
	notech_ao4 i_131068552(.A(n_54062), .B(n_60011), .C(n_56380), .D(n_27451
		), .Z(n_298290481));
	notech_ao4 i_130968553(.A(n_54082), .B(n_27743), .C(n_54073), .D(n_27785
		), .Z(n_298390482));
	notech_ao4 i_130868554(.A(n_54062), .B(n_60010), .C(n_56380), .D(n_27453
		), .Z(n_298490483));
	notech_ao4 i_130768555(.A(n_54082), .B(n_27744), .C(n_54073), .D(n_27786
		), .Z(n_298690484));
	notech_ao4 i_130668556(.A(n_54062), .B(n_60009), .C(n_56380), .D(n_27455
		), .Z(n_298790485));
	notech_ao4 i_130568557(.A(n_54082), .B(n_27745), .C(n_54073), .D(n_27787
		), .Z(n_298890486));
	notech_ao4 i_129668566(.A(n_54062), .B(n_60003), .C(n_56380), .D(n_27469
		), .Z(n_298990487));
	notech_ao4 i_129568567(.A(n_54082), .B(n_27752), .C(n_54073), .D(n_27793
		), .Z(n_299090488));
	notech_ao4 i_129468568(.A(n_54062), .B(n_60002), .C(n_56380), .D(n_27471
		), .Z(n_299190489));
	notech_ao4 i_129368569(.A(n_54082), .B(n_27755), .C(n_54073), .D(n_27794
		), .Z(n_299290490));
	notech_ao4 i_129268570(.A(n_54062), .B(n_60001), .C(n_56385), .D(n_27473
		), .Z(n_299390491));
	notech_ao4 i_129168571(.A(n_54082), .B(n_27756), .C(n_54073), .D(n_27795
		), .Z(n_299490492));
	notech_ao4 i_128868574(.A(n_54062), .B(n_133728614), .C(n_56385), .D(n_27477
		), .Z(n_299590493));
	notech_ao4 i_128768575(.A(n_54082), .B(n_27759), .C(n_54073), .D(n_27798
		), .Z(n_299690494));
	notech_ao4 i_128668576(.A(n_54062), .B(n_131228589), .C(n_56385), .D(n_27479
		), .Z(n_299790495));
	notech_ao4 i_128568577(.A(n_54082), .B(n_27760), .C(n_326890766), .D(n_27799
		), .Z(n_299890496));
	notech_ao4 i_128468578(.A(n_54062), .B(n_130528582), .C(n_56385), .D(n_27481
		), .Z(n_299990497));
	notech_ao4 i_128368579(.A(n_54082), .B(n_27762), .C(n_54073), .D(n_27800
		), .Z(n_300090498));
	notech_ao4 i_128268580(.A(n_128228559), .B(n_54062), .C(n_56385), .D(n_27483
		), .Z(n_300190499));
	notech_ao4 i_128168581(.A(n_54082), .B(n_27763), .C(n_54073), .D(n_27801
		), .Z(n_300290500));
	notech_ao4 i_128068582(.A(n_302991794), .B(n_54062), .C(n_56385), .D(n_27485
		), .Z(n_300390501));
	notech_ao4 i_127968583(.A(n_54082), .B(n_27764), .C(n_54073), .D(n_27802
		), .Z(n_300490502));
	notech_ao4 i_127868584(.A(n_54062), .B(n_314791676), .C(n_56390), .D(n_27487
		), .Z(n_300590503));
	notech_ao4 i_127768585(.A(n_54082), .B(n_27765), .C(n_54073), .D(n_27803
		), .Z(n_300690504));
	notech_ao4 i_127668586(.A(n_136661649), .B(n_27766), .C(n_54930), .D(n_27422
		), .Z(n_300790505));
	notech_ao4 i_127568587(.A(n_28124), .B(n_136861651), .C(n_136761650), .D
		(n_27728), .Z(n_300890506));
	notech_ao4 i_127468588(.A(n_136661649), .B(n_27767), .C(n_54930), .D(n_27424
		), .Z(n_300990507));
	notech_ao4 i_127368589(.A(n_136861651), .B(n_28125), .C(n_136761650), .D
		(n_27729), .Z(n_301090508));
	notech_ao4 i_127068592(.A(n_136661649), .B(n_27769), .C(n_54930), .D(n_27428
		), .Z(n_301190509));
	notech_ao4 i_126968593(.A(n_136861651), .B(n_28127), .C(n_136761650), .D
		(n_27731), .Z(n_301290510));
	notech_ao4 i_126868594(.A(n_136661649), .B(n_27770), .C(n_54930), .D(n_27430
		), .Z(n_301390511));
	notech_ao4 i_126768595(.A(n_136861651), .B(n_28128), .C(n_136761650), .D
		(n_27732), .Z(n_301490512));
	notech_ao4 i_126668596(.A(n_136661649), .B(n_27773), .C(n_54930), .D(n_27434
		), .Z(n_301590513));
	notech_ao4 i_126568597(.A(n_136861651), .B(n_28131), .C(n_136761650), .D
		(n_27734), .Z(n_301690514));
	notech_ao4 i_126468598(.A(n_136661649), .B(n_27774), .C(n_54930), .D(n_27437
		), .Z(n_301790515));
	notech_ao4 i_126368599(.A(n_136861651), .B(n_28133), .C(n_136761650), .D
		(n_27735), .Z(n_301890516));
	notech_ao4 i_126268600(.A(n_136661649), .B(n_27775), .C(n_54930), .D(n_27439
		), .Z(n_301990517));
	notech_ao4 i_126168601(.A(n_136861651), .B(n_28134), .C(n_136761650), .D
		(n_27737), .Z(n_302090518));
	notech_ao4 i_126068602(.A(n_136661649), .B(n_27776), .C(n_54930), .D(n_27441
		), .Z(n_302190519));
	notech_ao4 i_125968603(.A(n_136861651), .B(n_28135), .C(n_136761650), .D
		(n_27738), .Z(n_302290520));
	notech_ao4 i_125868604(.A(n_136661649), .B(n_27777), .C(n_54930), .D(n_27443
		), .Z(n_302390521));
	notech_ao4 i_125768605(.A(n_136861651), .B(n_28136), .C(n_136761650), .D
		(n_27739), .Z(n_302490522));
	notech_ao4 i_125668606(.A(n_136661649), .B(n_27779), .C(n_54930), .D(n_27445
		), .Z(n_302590523));
	notech_ao4 i_125568607(.A(n_136861651), .B(n_28137), .C(n_136761650), .D
		(n_27740), .Z(n_302690524));
	notech_ao4 i_125468608(.A(n_136661649), .B(n_27780), .C(n_54925), .D(n_27447
		), .Z(n_302790525));
	notech_ao4 i_125368609(.A(n_136861651), .B(n_28138), .C(n_136761650), .D
		(n_27741), .Z(n_302890526));
	notech_ao4 i_125268610(.A(n_136661649), .B(n_27783), .C(n_54925), .D(n_27449
		), .Z(n_302990527));
	notech_ao4 i_125168611(.A(n_136861651), .B(n_28139), .C(n_136761650), .D
		(n_27742), .Z(n_303090528));
	notech_ao4 i_125068612(.A(n_136661649), .B(n_27785), .C(n_54925), .D(n_27451
		), .Z(n_303190529));
	notech_ao4 i_124968613(.A(n_136861651), .B(n_28140), .C(n_136761650), .D
		(n_27743), .Z(n_303290530));
	notech_ao4 i_124868614(.A(n_136661649), .B(n_27786), .C(n_54925), .D(n_27453
		), .Z(n_303390531));
	notech_ao4 i_124768615(.A(n_136861651), .B(n_28141), .C(n_136761650), .D
		(n_27744), .Z(n_303490532));
	notech_ao4 i_124668616(.A(n_136661649), .B(n_27787), .C(n_54925), .D(n_27455
		), .Z(n_303590533));
	notech_ao4 i_124568617(.A(n_136861651), .B(n_28142), .C(n_136761650), .D
		(n_27745), .Z(n_303690534));
	notech_ao4 i_124468618(.A(n_54031), .B(n_27788), .C(n_54925), .D(n_27457
		), .Z(n_303790535));
	notech_ao4 i_124368619(.A(n_54051), .B(n_28143), .C(n_54042), .D(n_27747
		), .Z(n_303890536));
	notech_ao4 i_124268620(.A(n_54042), .B(n_27748), .C(n_54051), .D(n_28144
		), .Z(n_303990537));
	notech_ao4 i_124168621(.A(n_54925), .B(n_27459), .C(n_54031), .D(n_27789
		), .Z(n_304090538));
	notech_ao4 i_124068622(.A(n_54031), .B(n_27790), .C(n_54925), .D(n_27461
		), .Z(n_304190539));
	notech_ao4 i_123968623(.A(n_54051), .B(n_28145), .C(n_54042), .D(n_27749
		), .Z(n_304290540));
	notech_ao4 i_123868624(.A(n_54031), .B(n_27791), .C(n_54925), .D(n_27463
		), .Z(n_304390541));
	notech_ao4 i_123768625(.A(n_54051), .B(n_28146), .C(n_54042), .D(n_27750
		), .Z(n_304490542));
	notech_ao4 i_123668626(.A(n_54031), .B(n_27792), .C(n_54925), .D(n_27465
		), .Z(n_304590543));
	notech_ao4 i_123568627(.A(n_54051), .B(n_28147), .C(n_54042), .D(n_27751
		), .Z(n_304690544));
	notech_ao4 i_123468628(.A(n_54031), .B(n_27793), .C(n_54925), .D(n_27469
		), .Z(n_304790545));
	notech_ao4 i_123368629(.A(n_54051), .B(n_28148), .C(n_54042), .D(n_27752
		), .Z(n_304890546));
	notech_ao4 i_123268630(.A(n_54031), .B(n_27794), .C(n_54929), .D(n_27471
		), .Z(n_304990547));
	notech_ao4 i_123168631(.A(n_54051), .B(n_28149), .C(n_54042), .D(n_27755
		), .Z(n_305090548));
	notech_ao4 i_123068632(.A(n_54031), .B(n_27795), .C(n_54929), .D(n_27473
		), .Z(n_305190549));
	notech_ao4 i_122968633(.A(n_54051), .B(n_28150), .C(n_54042), .D(n_27756
		), .Z(n_305290550));
	notech_ao4 i_122868634(.A(n_54031), .B(n_27797), .C(n_54929), .D(n_27475
		), .Z(n_305390551));
	notech_ao4 i_122768635(.A(n_54051), .B(n_28151), .C(n_54042), .D(n_27758
		), .Z(n_305490552));
	notech_ao4 i_122668636(.A(n_54031), .B(n_27798), .C(n_54929), .D(n_27477
		), .Z(n_305590553));
	notech_ao4 i_122568637(.A(n_54051), .B(n_28152), .C(n_54042), .D(n_27759
		), .Z(n_305690554));
	notech_ao4 i_122468638(.A(n_54031), .B(n_27799), .C(n_54929), .D(n_27479
		), .Z(n_305790555));
	notech_ao4 i_122368639(.A(n_54051), .B(n_28153), .C(n_136761650), .D(n_27760
		), .Z(n_305890556));
	notech_ao4 i_122268640(.A(n_54031), .B(n_27800), .C(n_54925), .D(n_27481
		), .Z(n_305990557));
	notech_ao4 i_122168641(.A(n_54051), .B(n_28154), .C(n_54042), .D(n_27762
		), .Z(n_306090558));
	notech_ao4 i_122068642(.A(n_54031), .B(n_27801), .C(n_54925), .D(n_27483
		), .Z(n_306190559));
	notech_ao4 i_121968643(.A(n_54051), .B(n_28155), .C(n_54042), .D(n_27763
		), .Z(n_306290560));
	notech_ao4 i_121868644(.A(n_54031), .B(n_27802), .C(n_54925), .D(n_27485
		), .Z(n_306390561));
	notech_ao4 i_121768645(.A(n_54051), .B(n_28156), .C(n_54042), .D(n_27764
		), .Z(n_306490562));
	notech_ao4 i_121668646(.A(n_54031), .B(n_27803), .C(n_54929), .D(n_27487
		), .Z(n_306590563));
	notech_ao4 i_121568647(.A(n_54051), .B(n_28157), .C(n_54042), .D(n_27765
		), .Z(n_306690564));
	notech_ao4 i_121468648(.A(n_53890), .B(n_27768), .C(n_56894), .D(n_27426
		), .Z(n_306790565));
	notech_ao4 i_121368649(.A(n_54020), .B(n_30633), .C(n_53901), .D(n_27730
		), .Z(n_306890566));
	notech_ao4 i_121268650(.A(n_53890), .B(n_27770), .C(n_56894), .D(n_27430
		), .Z(n_306990567));
	notech_ao4 i_121168651(.A(n_54020), .B(n_30632), .C(n_53901), .D(n_27732
		), .Z(n_307090568));
	notech_ao4 i_121068652(.A(n_53890), .B(n_27771), .C(n_56894), .D(n_27432
		), .Z(n_307190569));
	notech_ao4 i_120968653(.A(n_54020), .B(n_30631), .C(n_349780998), .D(n_27733
		), .Z(n_307290570));
	notech_ao4 i_120868654(.A(n_53890), .B(n_27773), .C(n_56894), .D(n_27434
		), .Z(n_307390571));
	notech_ao4 i_120768655(.A(n_54020), .B(n_30630), .C(n_53901), .D(n_27734
		), .Z(n_307490572));
	notech_ao4 i_120668656(.A(n_53890), .B(n_27774), .C(n_56894), .D(n_27437
		), .Z(n_307590573));
	notech_ao4 i_120568657(.A(n_54020), .B(n_30629), .C(n_53901), .D(n_27735
		), .Z(n_307690574));
	notech_ao4 i_120468658(.A(n_53890), .B(n_27776), .C(n_56894), .D(n_27441
		), .Z(n_307790575));
	notech_ao4 i_120368659(.A(n_54020), .B(n_30628), .C(n_53901), .D(n_27738
		), .Z(n_307890576));
	notech_ao4 i_120268660(.A(n_53890), .B(n_27777), .C(n_56894), .D(n_27443
		), .Z(n_307990577));
	notech_ao4 i_120168661(.A(n_54020), .B(n_30627), .C(n_53901), .D(n_27739
		), .Z(n_308090578));
	notech_ao4 i_120068662(.A(n_53890), .B(n_27803), .C(n_56894), .D(n_27487
		), .Z(n_308190579));
	notech_ao4 i_119968663(.A(n_54020), .B(n_30626), .C(n_53901), .D(n_27765
		), .Z(n_308290580));
	notech_ao4 i_119568667(.A(n_27728), .B(n_152789026), .C(n_27766), .D(n_152889027
		), .Z(n_308490582));
	notech_ao4 i_119668666(.A(n_29633), .B(n_30955), .C(n_29665), .D(n_29635
		), .Z(n_308690584));
	notech_ao4 i_119468668(.A(n_3921), .B(n_27422), .C(n_152689025), .D(n_30625
		), .Z(n_308790585));
	notech_ao4 i_119368669(.A(n_152789026), .B(n_27729), .C(n_152889027), .D
		(n_27767), .Z(n_308890586));
	notech_ao4 i_119268670(.A(n_3921), .B(n_27424), .C(n_152689025), .D(n_30624
		), .Z(n_308990587));
	notech_ao4 i_119168671(.A(n_152789026), .B(n_27730), .C(n_152889027), .D
		(n_27768), .Z(n_309090588));
	notech_ao4 i_119068672(.A(n_3921), .B(n_27426), .C(n_152689025), .D(n_30623
		), .Z(n_309190589));
	notech_ao4 i_118968673(.A(n_152789026), .B(n_27731), .C(n_152889027), .D
		(n_27769), .Z(n_309290590));
	notech_ao4 i_118868674(.A(n_3921), .B(n_27428), .C(n_152689025), .D(n_30622
		), .Z(n_309390591));
	notech_ao4 i_118768675(.A(n_152789026), .B(n_27732), .C(n_152889027), .D
		(n_27770), .Z(n_309490592));
	notech_ao4 i_118668676(.A(n_3921), .B(n_27430), .C(n_152689025), .D(n_30621
		), .Z(n_309590593));
	notech_ao4 i_118568677(.A(n_152789026), .B(n_27733), .C(n_152889027), .D
		(n_27771), .Z(n_309690594));
	notech_ao4 i_118468678(.A(n_3921), .B(n_27432), .C(n_152689025), .D(n_30620
		), .Z(n_309790595));
	notech_ao4 i_118368679(.A(n_152789026), .B(n_27734), .C(n_152889027), .D
		(n_27773), .Z(n_309890596));
	notech_ao4 i_118268680(.A(n_3921), .B(n_27434), .C(n_152689025), .D(n_30619
		), .Z(n_309990597));
	notech_ao4 i_118168681(.A(n_152789026), .B(n_27735), .C(n_152889027), .D
		(n_27774), .Z(n_310090598));
	notech_ao4 i_118068682(.A(n_3921), .B(n_27437), .C(n_152689025), .D(n_30618
		), .Z(n_310190599));
	notech_ao4 i_117968683(.A(n_152789026), .B(n_27737), .C(n_152889027), .D
		(n_27775), .Z(n_310290600));
	notech_ao4 i_117868684(.A(n_3921), .B(n_27439), .C(n_152689025), .D(n_30617
		), .Z(n_310390601));
	notech_ao4 i_117768685(.A(n_152789026), .B(n_27738), .C(n_152889027), .D
		(n_27776), .Z(n_310490602));
	notech_ao4 i_117668686(.A(n_3921), .B(n_27441), .C(n_152689025), .D(n_30616
		), .Z(n_310590603));
	notech_ao4 i_117568687(.A(n_152789026), .B(n_27739), .C(n_152889027), .D
		(n_27777), .Z(n_310690604));
	notech_ao4 i_117468688(.A(n_3921), .B(n_27443), .C(n_152689025), .D(n_30615
		), .Z(n_310790605));
	notech_ao4 i_117368689(.A(n_152789026), .B(n_27740), .C(n_152889027), .D
		(n_27779), .Z(n_310890606));
	notech_ao4 i_117268690(.A(n_3921), .B(n_27445), .C(n_152689025), .D(n_30614
		), .Z(n_310990607));
	notech_ao4 i_117168691(.A(n_152789026), .B(n_27741), .C(n_152889027), .D
		(n_27780), .Z(n_311090608));
	notech_ao4 i_117068692(.A(n_3921), .B(n_27447), .C(n_152689025), .D(n_30613
		), .Z(n_311190609));
	notech_ao4 i_116968693(.A(n_152789026), .B(n_27742), .C(n_152889027), .D
		(n_27783), .Z(n_311290610));
	notech_ao4 i_116868694(.A(n_56992), .B(n_27449), .C(n_152689025), .D(n_30612
		), .Z(n_311390611));
	notech_ao4 i_116768695(.A(n_53709), .B(n_27743), .C(n_53700), .D(n_27785
		), .Z(n_311490612));
	notech_ao4 i_116668696(.A(n_56992), .B(n_27451), .C(n_53830), .D(n_30611
		), .Z(n_311590613));
	notech_ao4 i_116568697(.A(n_53709), .B(n_27744), .C(n_53700), .D(n_27786
		), .Z(n_311690614));
	notech_ao4 i_116468698(.A(n_56992), .B(n_27453), .C(n_53830), .D(n_30610
		), .Z(n_311790615));
	notech_ao4 i_116368699(.A(n_53709), .B(n_27745), .C(n_53700), .D(n_27787
		), .Z(n_311890616));
	notech_ao4 i_116268700(.A(n_56992), .B(n_27455), .C(n_53830), .D(n_30609
		), .Z(n_311990617));
	notech_ao4 i_116168701(.A(n_53709), .B(n_27747), .C(n_53700), .D(n_27788
		), .Z(n_312090618));
	notech_ao4 i_116068702(.A(n_56992), .B(n_27457), .C(n_53830), .D(n_30608
		), .Z(n_312190619));
	notech_ao4 i_115968703(.A(n_53709), .B(n_27748), .C(n_53700), .D(n_27789
		), .Z(n_312290620));
	notech_ao4 i_115868704(.A(n_56992), .B(n_27459), .C(n_53830), .D(n_30605
		), .Z(n_312390621));
	notech_ao4 i_115768705(.A(n_53709), .B(n_27749), .C(n_53700), .D(n_27790
		), .Z(n_312490622));
	notech_ao4 i_115668706(.A(n_56992), .B(n_27461), .C(n_53830), .D(n_30604
		), .Z(n_312590623));
	notech_ao4 i_115568707(.A(n_53709), .B(n_27752), .C(n_53700), .D(n_27793
		), .Z(n_312690624));
	notech_ao4 i_115468708(.A(n_56992), .B(n_27469), .C(n_53830), .D(n_30603
		), .Z(n_312790625));
	notech_ao4 i_115368709(.A(n_53709), .B(n_27755), .C(n_53700), .D(n_27794
		), .Z(n_312890626));
	notech_ao4 i_115268710(.A(n_56992), .B(n_27471), .C(n_53830), .D(n_30602
		), .Z(n_312990627));
	notech_ao4 i_115168711(.A(n_53709), .B(n_27756), .C(n_53700), .D(n_27795
		), .Z(n_313090628));
	notech_ao4 i_115068712(.A(n_56992), .B(n_27473), .C(n_53830), .D(n_30601
		), .Z(n_313190629));
	notech_ao4 i_114968713(.A(n_53709), .B(n_27758), .C(n_53700), .D(n_27797
		), .Z(n_313290630));
	notech_ao4 i_114868714(.A(n_56992), .B(n_27475), .C(n_53830), .D(n_30600
		), .Z(n_313390631));
	notech_ao4 i_114768715(.A(n_53709), .B(n_27759), .C(n_152889027), .D(n_27798
		), .Z(n_313490632));
	notech_ao4 i_114668716(.A(n_56992), .B(n_27477), .C(n_152689025), .D(n_30599
		), .Z(n_313590633));
	notech_ao4 i_114568717(.A(n_53709), .B(n_27760), .C(n_53700), .D(n_27799
		), .Z(n_313690634));
	notech_ao4 i_114468718(.A(n_56992), .B(n_27479), .C(n_53830), .D(n_30597
		), .Z(n_313790635));
	notech_ao4 i_114368719(.A(n_53709), .B(n_27762), .C(n_53700), .D(n_27800
		), .Z(n_313890636));
	notech_ao4 i_114268720(.A(n_56992), .B(n_27481), .C(n_53830), .D(n_30596
		), .Z(n_313990637));
	notech_ao4 i_114168721(.A(n_53709), .B(n_27763), .C(n_53700), .D(n_27801
		), .Z(n_314090638));
	notech_ao4 i_114068722(.A(n_56992), .B(n_27483), .C(n_30595), .D(n_53830
		), .Z(n_314190639));
	notech_ao4 i_113968723(.A(n_53709), .B(n_27764), .C(n_53700), .D(n_27802
		), .Z(n_314290640));
	notech_ao4 i_113868724(.A(n_56992), .B(n_27485), .C(n_53830), .D(n_30593
		), .Z(n_314390641));
	notech_ao4 i_113768725(.A(n_53709), .B(n_27765), .C(n_53700), .D(n_27803
		), .Z(n_314490642));
	notech_ao4 i_113668726(.A(n_56992), .B(n_27487), .C(n_53830), .D(n_30592
		), .Z(n_314590643));
	notech_or4 i_9169856(.A(instrc[90]), .B(instrc[88]), .C(n_29631), .D(n_29640
		), .Z(n_314690644));
	notech_ao4 i_113468728(.A(n_30976), .B(n_29642), .C(instrc[89]), .D(instrc
		[90]), .Z(n_314890646));
	notech_nand2 i_8969858(.A(n_3918), .B(n_152989028), .Z(n_314990647));
	notech_ao4 i_113268730(.A(n_314990647), .B(n_30591), .C(n_27728), .D(n_314690644
		), .Z(n_315090648));
	notech_or4 i_7169871(.A(n_3673), .B(instrc[89]), .C(n_29668), .D(n_29640
		), .Z(n_315290650));
	notech_ao4 i_113168731(.A(n_3918), .B(n_27422), .C(n_27766), .D(n_315290650
		), .Z(n_315390651));
	notech_ao4 i_113068732(.A(n_314990647), .B(n_30590), .C(n_314690644), .D
		(n_27729), .Z(n_315490652));
	notech_ao4 i_112968733(.A(n_3918), .B(n_27424), .C(n_27767), .D(n_315290650
		), .Z(n_315590653));
	notech_ao4 i_112868734(.A(n_314990647), .B(n_30589), .C(n_314690644), .D
		(n_27730), .Z(n_315690654));
	notech_ao4 i_112768735(.A(n_3918), .B(n_27426), .C(n_27768), .D(n_315290650
		), .Z(n_315790655));
	notech_ao4 i_112668736(.A(n_314990647), .B(n_30587), .C(n_314690644), .D
		(n_27731), .Z(n_315890656));
	notech_ao4 i_112568737(.A(n_3918), .B(n_27428), .C(n_27769), .D(n_315290650
		), .Z(n_315990657));
	notech_ao4 i_112468738(.A(n_314990647), .B(n_30586), .C(n_314690644), .D
		(n_27732), .Z(n_316090658));
	notech_ao4 i_112368739(.A(n_3918), .B(n_27430), .C(n_27770), .D(n_315290650
		), .Z(n_316190659));
	notech_ao4 i_112268740(.A(n_314990647), .B(n_30585), .C(n_314690644), .D
		(n_27733), .Z(n_316290660));
	notech_ao4 i_112168741(.A(n_3918), .B(n_27432), .C(n_27771), .D(n_315290650
		), .Z(n_316390661));
	notech_ao4 i_112068742(.A(n_314990647), .B(n_30581), .C(n_314690644), .D
		(n_27734), .Z(n_316490662));
	notech_ao4 i_111968743(.A(n_3918), .B(n_27434), .C(n_27773), .D(n_315290650
		), .Z(n_316590663));
	notech_ao4 i_111868744(.A(n_314990647), .B(n_30580), .C(n_314690644), .D
		(n_27735), .Z(n_316690664));
	notech_ao4 i_111768745(.A(n_3918), .B(n_27437), .C(n_27774), .D(n_315290650
		), .Z(n_316790665));
	notech_ao4 i_111668746(.A(n_314990647), .B(n_30579), .C(n_314690644), .D
		(n_27737), .Z(n_316890666));
	notech_ao4 i_111568747(.A(n_3918), .B(n_27439), .C(n_27775), .D(n_315290650
		), .Z(n_316990667));
	notech_ao4 i_111468748(.A(n_314990647), .B(n_30578), .C(n_314690644), .D
		(n_27738), .Z(n_317090668));
	notech_ao4 i_111368749(.A(n_3918), .B(n_27441), .C(n_27776), .D(n_315290650
		), .Z(n_317190669));
	notech_ao4 i_111268750(.A(n_314990647), .B(n_30577), .C(n_314690644), .D
		(n_27739), .Z(n_317290670));
	notech_ao4 i_111168751(.A(n_3918), .B(n_27443), .C(n_27777), .D(n_315290650
		), .Z(n_317390671));
	notech_ao4 i_111068752(.A(n_314990647), .B(n_30576), .C(n_314690644), .D
		(n_27740), .Z(n_317490672));
	notech_ao4 i_110968753(.A(n_3918), .B(n_27445), .C(n_27779), .D(n_315290650
		), .Z(n_317590673));
	notech_ao4 i_110868754(.A(n_314990647), .B(n_30575), .C(n_314690644), .D
		(n_27741), .Z(n_317690674));
	notech_ao4 i_110768755(.A(n_3918), .B(n_27447), .C(n_27780), .D(n_315290650
		), .Z(n_317790675));
	notech_ao4 i_110668756(.A(n_314990647), .B(n_30574), .C(n_314690644), .D
		(n_27742), .Z(n_317890676));
	notech_ao4 i_110568757(.A(n_3918), .B(n_27449), .C(n_27783), .D(n_315290650
		), .Z(n_317990677));
	notech_ao4 i_110468758(.A(n_314990647), .B(n_30573), .C(n_314690644), .D
		(n_27743), .Z(n_318090678));
	notech_ao4 i_110368759(.A(n_3918), .B(n_27451), .C(n_27785), .D(n_315290650
		), .Z(n_318190679));
	notech_ao4 i_110268760(.A(n_314990647), .B(n_30572), .C(n_314690644), .D
		(n_27744), .Z(n_318290680));
	notech_ao4 i_110168761(.A(n_57092), .B(n_27453), .C(n_27786), .D(n_315290650
		), .Z(n_318390681));
	notech_ao4 i_110068762(.A(n_53400), .B(n_30571), .C(n_53281), .D(n_27745
		), .Z(n_318490682));
	notech_ao4 i_109968763(.A(n_57092), .B(n_27455), .C(n_27787), .D(n_53411
		), .Z(n_318590683));
	notech_ao4 i_109868764(.A(n_53400), .B(n_30567), .C(n_53281), .D(n_27747
		), .Z(n_318690684));
	notech_ao4 i_109768765(.A(n_57092), .B(n_27457), .C(n_27788), .D(n_53411
		), .Z(n_318790685));
	notech_ao4 i_109668766(.A(n_53400), .B(n_30566), .C(n_53281), .D(n_27748
		), .Z(n_318890686));
	notech_ao4 i_109568767(.A(n_57092), .B(n_27459), .C(n_27789), .D(n_53411
		), .Z(n_318990687));
	notech_ao4 i_109468768(.A(n_53400), .B(n_30564), .C(n_53281), .D(n_27749
		), .Z(n_319090688));
	notech_ao4 i_109368769(.A(n_57092), .B(n_27461), .C(n_27790), .D(n_53411
		), .Z(n_319190689));
	notech_ao4 i_109268770(.A(n_53400), .B(n_30563), .C(n_53281), .D(n_27750
		), .Z(n_319290690));
	notech_ao4 i_109168771(.A(n_57092), .B(n_27463), .C(n_27791), .D(n_53411
		), .Z(n_319390691));
	notech_ao4 i_109068772(.A(n_53400), .B(n_30562), .C(n_53281), .D(n_27751
		), .Z(n_319490692));
	notech_ao4 i_108968773(.A(n_57092), .B(n_27465), .C(n_27792), .D(n_53411
		), .Z(n_319590693));
	notech_ao4 i_108868774(.A(n_53400), .B(n_30561), .C(n_53281), .D(n_27752
		), .Z(n_319690694));
	notech_ao4 i_108768775(.A(n_57092), .B(n_27469), .C(n_27793), .D(n_53411
		), .Z(n_319790695));
	notech_ao4 i_108668776(.A(n_53400), .B(n_30560), .C(n_53281), .D(n_27755
		), .Z(n_319890696));
	notech_ao4 i_108568777(.A(n_57092), .B(n_27471), .C(n_27794), .D(n_53411
		), .Z(n_319990697));
	notech_ao4 i_108468778(.A(n_53400), .B(n_30559), .C(n_53281), .D(n_27756
		), .Z(n_320090698));
	notech_ao4 i_108368779(.A(n_57092), .B(n_27473), .C(n_27795), .D(n_53411
		), .Z(n_320190699));
	notech_ao4 i_108268780(.A(n_53400), .B(n_30558), .C(n_53281), .D(n_27758
		), .Z(n_320290700));
	notech_ao4 i_108168781(.A(n_57092), .B(n_27475), .C(n_27797), .D(n_53411
		), .Z(n_320390701));
	notech_ao4 i_108068782(.A(n_53400), .B(n_30557), .C(n_314690644), .D(n_27759
		), .Z(n_320490702));
	notech_ao4 i_107968783(.A(n_3918), .B(n_27477), .C(n_27798), .D(n_315290650
		), .Z(n_320590703));
	notech_ao4 i_107868784(.A(n_53400), .B(n_30556), .C(n_53281), .D(n_27760
		), .Z(n_320690704));
	notech_ao4 i_107768785(.A(n_57092), .B(n_27479), .C(n_27799), .D(n_53411
		), .Z(n_320790705));
	notech_ao4 i_107668786(.A(n_53400), .B(n_30555), .C(n_53281), .D(n_27762
		), .Z(n_320890706));
	notech_ao4 i_107568787(.A(n_57092), .B(n_27481), .C(n_27800), .D(n_53411
		), .Z(n_320990707));
	notech_ao4 i_107468788(.A(n_53400), .B(n_30554), .C(n_53281), .D(n_27763
		), .Z(n_321090708));
	notech_ao4 i_107368789(.A(n_57092), .B(n_27483), .C(n_27801), .D(n_53411
		), .Z(n_321190709));
	notech_ao4 i_107268790(.A(n_53400), .B(n_30553), .C(n_53281), .D(n_27764
		), .Z(n_321290710));
	notech_ao4 i_107168791(.A(n_57092), .B(n_27485), .C(n_27802), .D(n_53411
		), .Z(n_321390711));
	notech_ao4 i_107068792(.A(n_53400), .B(n_30552), .C(n_53281), .D(n_27765
		), .Z(n_321490712));
	notech_ao4 i_106968793(.A(n_57092), .B(n_27487), .C(n_27803), .D(n_53411
		), .Z(n_321590713));
	notech_ao4 i_49131(.A(n_27085), .B(n_135041965), .C(n_346670477), .D(n_29793
		), .Z(\nbus_11311[0] ));
	notech_or4 i_9867303(.A(n_27925), .B(n_60874), .C(\opcode[3] ), .D(n_27084
		), .Z(n_321890716));
	notech_nand2 i_48961(.A(n_321890716), .B(n_58691), .Z(n_14425));
	notech_ao4 i_53878(.A(n_29656), .B(n_322490722), .C(n_135041965), .D(n_57966
		), .Z(\nbus_11353[0] ));
	notech_or4 i_34367081(.A(n_59418), .B(n_61109), .C(n_32729), .D(n_27573)
		, .Z(n_322190719));
	notech_nand3 i_52736(.A(n_114668163), .B(n_322190719), .C(n_26992), .Z(n_19963
		));
	notech_nand2 i_47674(.A(n_53748), .B(n_58666), .Z(n_12080));
	notech_mux2 i_5252(.S(n_60316), .A(n_19086), .B(n_317291651), .Z(n_13729
		));
	notech_nand3 i_9854(.A(n_19065), .B(n_26983), .C(n_60212), .Z(n_14792)
		);
	notech_or4 i_27067151(.A(n_59322), .B(n_26900), .C(n_60372), .D(n_29793)
		, .Z(n_322490722));
	notech_or2 i_3767364(.A(n_32259), .B(\opcode[3] ), .Z(n_69641311));
	notech_or4 i_46066967(.A(n_32323), .B(n_58024), .C(n_32316), .D(n_57992)
		, .Z(n_323190729));
	notech_or4 i_5764396(.A(n_29638), .B(n_30966), .C(n_323490732), .D(n_27092
		), .Z(n_323390731));
	notech_and2 i_87663600(.A(n_30969), .B(instrc[92]), .Z(n_323490732));
	notech_or4 i_98863490(.A(n_60863), .B(n_27924), .C(n_61133), .D(n_60212)
		, .Z(n_323590733));
	notech_or4 i_39291(.A(instrc[93]), .B(n_29666), .C(n_29638), .D(n_3919),
		 .Z(n_324090738));
	notech_or4 i_39293(.A(n_26886), .B(instrc[92]), .C(n_29638), .D(n_3919),
		 .Z(n_324190739));
	notech_nand2 i_39297(.A(n_57002), .B(n_323390731), .Z(n_324290740));
	notech_ao4 i_161362888(.A(n_154279046), .B(n_27742), .C(n_154379047), .D
		(n_27783), .Z(n_325190749));
	notech_ao4 i_161162889(.A(n_27107), .B(n_27449), .C(n_29592), .D(n_154179045
		), .Z(n_325290750));
	notech_ao4 i_160462894(.A(n_54042), .B(n_27733), .C(n_54051), .D(n_28129
		), .Z(n_325390751));
	notech_ao4 i_160362895(.A(n_54929), .B(n_27432), .C(n_54031), .D(n_27771
		), .Z(n_325490752));
	notech_ao4 i_159862899(.A(n_27762), .B(n_53431), .C(n_53550), .D(n_30634
		), .Z(n_325890756));
	notech_ao4 i_159762900(.A(n_57002), .B(n_27481), .C(n_53420), .D(n_27800
		), .Z(n_325990757));
	notech_nand3 i_3253880(.A(n_212969141), .B(n_3986), .C(n_346770478), .Z(n_326090758
		));
	notech_ao4 i_7782(.A(n_2985), .B(n_3885), .C(n_3986), .D(CFOF_mul), .Z(n_21654
		));
	notech_or4 i_38938(.A(n_60975), .B(n_29179), .C(n_26735), .D(n_32334), .Z
		(n_326790765));
	notech_nand3 i_38940(.A(n_56414), .B(n_56385), .C(n_327090768), .Z(n_326890766
		));
	notech_or4 i_38944(.A(n_32319), .B(n_32334), .C(n_32332), .D(n_32338), .Z
		(n_326990767));
	notech_nand2 i_1638218(.A(n_56447), .B(n_56452), .Z(n_327090768));
	notech_ao4 i_214536163(.A(n_54073), .B(n_27789), .C(n_3864), .D(n_54062)
		, .Z(n_327290770));
	notech_ao4 i_214436164(.A(n_56385), .B(n_27459), .C(n_54082), .D(n_27748
		), .Z(n_327390771));
	notech_or4 i_113034005(.A(n_61109), .B(n_60933), .C(n_60909), .D(n_27095
		), .Z(n_327490772));
	notech_or4 i_113134004(.A(n_61109), .B(n_27924), .C(n_60933), .D(n_60904
		), .Z(n_327590773));
	notech_nand2 i_1117888(.A(n_133088829), .B(n_132988828), .Z(write_data_25
		[10]));
	notech_nand2 i_1217889(.A(n_133288831), .B(n_133188830), .Z(write_data_25
		[11]));
	notech_nand2 i_1317890(.A(n_133488833), .B(n_133388832), .Z(write_data_25
		[12]));
	notech_nand2 i_1517892(.A(n_133688835), .B(n_133588834), .Z(write_data_25
		[14]));
	notech_nand2 i_3017907(.A(n_133888837), .B(n_133788836), .Z(write_data_25
		[29]));
	notech_nand2 i_3117908(.A(n_134088839), .B(n_133988838), .Z(write_data_25
		[30]));
	notech_nand2 i_3217909(.A(n_134288841), .B(n_134188840), .Z(write_data_25
		[31]));
	notech_nand2 i_118262(.A(n_134488843), .B(n_134388842), .Z(write_data_28
		[0]));
	notech_nand2 i_218263(.A(n_134688845), .B(n_134588844), .Z(write_data_28
		[1]));
	notech_nand2 i_918270(.A(n_134888847), .B(n_134788846), .Z(write_data_28
		[8]));
	notech_nand2 i_1218273(.A(n_135088849), .B(n_134988848), .Z(write_data_28
		[11]));
	notech_nand2 i_1318274(.A(n_135288851), .B(n_135188850), .Z(write_data_28
		[12]));
	notech_nand2 i_1418275(.A(n_135488853), .B(n_135388852), .Z(write_data_28
		[13]));
	notech_nand2 i_1518276(.A(n_135688855), .B(n_135588854), .Z(write_data_28
		[14]));
	notech_nand2 i_1618277(.A(n_135888857), .B(n_135788856), .Z(write_data_28
		[15]));
	notech_nand2 i_1718278(.A(n_136088859), .B(n_135988858), .Z(write_data_28
		[16]));
	notech_nand2 i_1818279(.A(n_136288861), .B(n_136188860), .Z(write_data_28
		[17]));
	notech_nand2 i_1918280(.A(n_136488863), .B(n_136388862), .Z(write_data_28
		[18]));
	notech_nand2 i_2018281(.A(n_136688865), .B(n_136588864), .Z(write_data_28
		[19]));
	notech_nand2 i_2118282(.A(n_136888867), .B(n_136788866), .Z(write_data_28
		[20]));
	notech_nand2 i_2218283(.A(n_137088869), .B(n_136988868), .Z(write_data_28
		[21]));
	notech_nand2 i_2318284(.A(n_137288871), .B(n_137188870), .Z(write_data_28
		[22]));
	notech_nand2 i_2418285(.A(n_137488873), .B(n_137388872), .Z(write_data_28
		[23]));
	notech_nand2 i_2518286(.A(n_137688875), .B(n_137588874), .Z(write_data_28
		[24]));
	notech_nand2 i_2618287(.A(n_137888877), .B(n_137788876), .Z(write_data_28
		[25]));
	notech_nand2 i_2718288(.A(n_138088879), .B(n_137988878), .Z(write_data_28
		[26]));
	notech_nand2 i_2818289(.A(n_138288881), .B(n_138188880), .Z(write_data_28
		[27]));
	notech_nand2 i_2918290(.A(n_138488883), .B(n_138388882), .Z(write_data_28
		[28]));
	notech_nand2 i_3018291(.A(n_138688885), .B(n_138588884), .Z(write_data_28
		[29]));
	notech_nand2 i_3118292(.A(n_138888887), .B(n_138788886), .Z(write_data_28
		[30]));
	notech_nand2 i_2118410(.A(n_139088889), .B(n_138988888), .Z(write_data_29
		[20]));
	notech_nand2 i_2218411(.A(n_139288891), .B(n_139188890), .Z(write_data_29
		[21]));
	notech_nand2 i_118518(.A(n_140188900), .B(n_139888897), .Z(write_data_30
		[0]));
	notech_nand2 i_218519(.A(n_140388902), .B(n_140288901), .Z(write_data_30
		[1]));
	notech_nand2 i_318520(.A(n_140588904), .B(n_140488903), .Z(write_data_30
		[2]));
	notech_nand2 i_418521(.A(n_140788906), .B(n_140688905), .Z(write_data_30
		[3]));
	notech_nand2 i_518522(.A(n_140988908), .B(n_140888907), .Z(write_data_30
		[4]));
	notech_nand2 i_618523(.A(n_141188910), .B(n_141088909), .Z(write_data_30
		[5]));
	notech_nand2 i_718524(.A(n_141388912), .B(n_141288911), .Z(write_data_30
		[6]));
	notech_nand2 i_818525(.A(n_141588914), .B(n_141488913), .Z(write_data_30
		[7]));
	notech_nand2 i_918526(.A(n_141788916), .B(n_141688915), .Z(write_data_30
		[8]));
	notech_nand2 i_1018527(.A(n_141988918), .B(n_141888917), .Z(write_data_30
		[9]));
	notech_nand2 i_1118528(.A(n_142188920), .B(n_142088919), .Z(write_data_30
		[10]));
	notech_nand2 i_1218529(.A(n_142388922), .B(n_142288921), .Z(write_data_30
		[11]));
	notech_nand2 i_1318530(.A(n_142588924), .B(n_142488923), .Z(write_data_30
		[12]));
	notech_nand2 i_1418531(.A(n_142788926), .B(n_142688925), .Z(write_data_30
		[13]));
	notech_nand2 i_1518532(.A(n_142988928), .B(n_142888927), .Z(write_data_30
		[14]));
	notech_nand2 i_1618533(.A(n_143188930), .B(n_143088929), .Z(write_data_30
		[15]));
	notech_nand2 i_1718534(.A(n_143388932), .B(n_143288931), .Z(write_data_30
		[16]));
	notech_nand2 i_1818535(.A(n_143588934), .B(n_143488933), .Z(write_data_30
		[17]));
	notech_nand2 i_1918536(.A(n_143788936), .B(n_143688935), .Z(write_data_30
		[18]));
	notech_nand2 i_2018537(.A(n_143988938), .B(n_143888937), .Z(write_data_30
		[19]));
	notech_nand2 i_2118538(.A(n_144188940), .B(n_144088939), .Z(write_data_30
		[20]));
	notech_nand2 i_2218539(.A(n_144388942), .B(n_144288941), .Z(write_data_30
		[21]));
	notech_nand2 i_2318540(.A(n_144588944), .B(n_144488943), .Z(write_data_30
		[22]));
	notech_nand2 i_2418541(.A(n_144788946), .B(n_144688945), .Z(write_data_30
		[23]));
	notech_nand2 i_2518542(.A(n_144988948), .B(n_144888947), .Z(write_data_30
		[24]));
	notech_nand2 i_2618543(.A(n_145188950), .B(n_145088949), .Z(write_data_30
		[25]));
	notech_nand2 i_2718544(.A(n_145388952), .B(n_145288951), .Z(write_data_30
		[26]));
	notech_nand2 i_2818545(.A(n_145588954), .B(n_145488953), .Z(write_data_30
		[27]));
	notech_nand2 i_2918546(.A(n_145788956), .B(n_145688955), .Z(write_data_30
		[28]));
	notech_nand2 i_3018547(.A(n_145988958), .B(n_145888957), .Z(write_data_30
		[29]));
	notech_nand2 i_3118548(.A(n_146188960), .B(n_146088959), .Z(write_data_30
		[30]));
	notech_nand2 i_3218549(.A(n_146388962), .B(n_146288961), .Z(write_data_30
		[31]));
	notech_nand2 i_118646(.A(n_146588964), .B(n_146488963), .Z(write_data_31
		[0]));
	notech_nand2 i_218647(.A(n_146788966), .B(n_146688965), .Z(write_data_31
		[1]));
	notech_nand2 i_318648(.A(n_146988968), .B(n_146888967), .Z(write_data_31
		[2]));
	notech_nand2 i_418649(.A(n_147188970), .B(n_147088969), .Z(write_data_31
		[3]));
	notech_nand2 i_518650(.A(n_147388972), .B(n_147288971), .Z(write_data_31
		[4]));
	notech_nand2 i_618651(.A(n_147588974), .B(n_147488973), .Z(write_data_31
		[5]));
	notech_nand2 i_718652(.A(n_147788976), .B(n_147688975), .Z(write_data_31
		[6]));
	notech_nand2 i_818653(.A(n_147988978), .B(n_147888977), .Z(write_data_31
		[7]));
	notech_nand2 i_918654(.A(n_148188980), .B(n_148088979), .Z(write_data_31
		[8]));
	notech_nand2 i_1018655(.A(n_148388982), .B(n_148288981), .Z(write_data_31
		[9]));
	notech_nand2 i_1118656(.A(n_148588984), .B(n_148488983), .Z(write_data_31
		[10]));
	notech_nand2 i_1218657(.A(n_148788986), .B(n_148688985), .Z(write_data_31
		[11]));
	notech_nand2 i_1318658(.A(n_148988988), .B(n_148888987), .Z(write_data_31
		[12]));
	notech_nand2 i_1418659(.A(n_149188990), .B(n_149088989), .Z(write_data_31
		[13]));
	notech_nand2 i_1518660(.A(n_149388992), .B(n_149288991), .Z(write_data_31
		[14]));
	notech_nand2 i_1618661(.A(n_149588994), .B(n_149488993), .Z(write_data_31
		[15]));
	notech_nand2 i_1718662(.A(n_149788996), .B(n_149688995), .Z(write_data_31
		[16]));
	notech_nand2 i_1818663(.A(n_149988998), .B(n_149888997), .Z(write_data_31
		[17]));
	notech_nand2 i_1918664(.A(n_150189000), .B(n_150088999), .Z(write_data_31
		[18]));
	notech_nand2 i_2018665(.A(n_150389002), .B(n_150289001), .Z(write_data_31
		[19]));
	notech_nand2 i_2118666(.A(n_150589004), .B(n_150489003), .Z(write_data_31
		[20]));
	notech_nand2 i_2218667(.A(n_150789006), .B(n_150689005), .Z(write_data_31
		[21]));
	notech_nand2 i_2318668(.A(n_150989008), .B(n_150889007), .Z(write_data_31
		[22]));
	notech_nand2 i_2418669(.A(n_151189010), .B(n_151089009), .Z(write_data_31
		[23]));
	notech_nand2 i_2518670(.A(n_151389012), .B(n_151289011), .Z(write_data_31
		[24]));
	notech_nand2 i_2618671(.A(n_151589014), .B(n_151489013), .Z(write_data_31
		[25]));
	notech_nand2 i_2718672(.A(n_151789016), .B(n_151689015), .Z(write_data_31
		[26]));
	notech_nand2 i_2818673(.A(n_151989018), .B(n_151889017), .Z(write_data_31
		[27]));
	notech_nand2 i_3018675(.A(n_152189020), .B(n_152089019), .Z(write_data_31
		[29]));
	notech_nand2 i_3118676(.A(n_152389022), .B(n_152289021), .Z(write_data_31
		[30]));
	notech_nand2 i_3218677(.A(n_152589024), .B(n_152489023), .Z(write_data_31
		[31]));
	notech_nand2 i_52755(.A(n_60123), .B(n_58666), .Z(n_19986));
	notech_and4 i_111990(.A(n_256390062), .B(n_256190060), .C(n_255790056), 
		.D(n_254990048), .Z(to_acu100236[0]));
	notech_and4 i_211991(.A(n_256990068), .B(n_256890067), .C(n_256690065), 
		.D(n_256590064), .Z(to_acu100236[1]));
	notech_and4 i_311992(.A(n_257590074), .B(n_257490073), .C(n_257290071), 
		.D(n_257190070), .Z(to_acu100236[2]));
	notech_and4 i_411993(.A(n_258190080), .B(n_258090079), .C(n_257890077), 
		.D(n_257790076), .Z(to_acu100236[3]));
	notech_and4 i_511994(.A(n_258790086), .B(n_258690085), .C(n_258490083), 
		.D(n_258390082), .Z(to_acu100236[4]));
	notech_and4 i_611995(.A(n_259390092), .B(n_259290091), .C(n_259090089), 
		.D(n_258990088), .Z(to_acu100236[5]));
	notech_and4 i_711996(.A(n_259990098), .B(n_259890097), .C(n_259690095), 
		.D(n_259590094), .Z(to_acu100236[6]));
	notech_and4 i_811997(.A(n_260590104), .B(n_260490103), .C(n_260290101), 
		.D(n_260190100), .Z(to_acu100236[7]));
	notech_and4 i_911998(.A(n_261190110), .B(n_261090109), .C(n_260890107), 
		.D(n_260790106), .Z(to_acu100236[8]));
	notech_and4 i_1011999(.A(n_261790116), .B(n_261690115), .C(n_261490113),
		 .D(n_261390112), .Z(to_acu100236[9]));
	notech_and4 i_1112000(.A(n_262390122), .B(n_262290121), .C(n_262090119),
		 .D(n_261990118), .Z(to_acu100236[10]));
	notech_and4 i_1212001(.A(n_262990128), .B(n_262890127), .C(n_262690125),
		 .D(n_262590124), .Z(to_acu100236[11]));
	notech_and4 i_1312002(.A(n_263590134), .B(n_263490133), .C(n_263290131),
		 .D(n_263190130), .Z(to_acu100236[12]));
	notech_and4 i_1412003(.A(n_264190140), .B(n_264090139), .C(n_263890137),
		 .D(n_263790136), .Z(to_acu100236[13]));
	notech_and4 i_1512004(.A(n_264790146), .B(n_264690145), .C(n_264490143),
		 .D(n_264390142), .Z(to_acu100236[14]));
	notech_and4 i_1612005(.A(n_265390152), .B(n_265290151), .C(n_265090149),
		 .D(n_264990148), .Z(to_acu100236[15]));
	notech_and4 i_1712006(.A(n_265990158), .B(n_265890157), .C(n_265690155),
		 .D(n_265590154), .Z(to_acu100236[16]));
	notech_and4 i_1812007(.A(n_266590164), .B(n_266490163), .C(n_266290161),
		 .D(n_266190160), .Z(to_acu100236[17]));
	notech_and4 i_1912008(.A(n_267190170), .B(n_267090169), .C(n_266890167),
		 .D(n_266790166), .Z(to_acu100236[18]));
	notech_and4 i_2012009(.A(n_267790176), .B(n_267690175), .C(n_267490173),
		 .D(n_267390172), .Z(to_acu100236[19]));
	notech_and4 i_2112010(.A(n_268390182), .B(n_268290181), .C(n_268090179),
		 .D(n_267990178), .Z(to_acu100236[20]));
	notech_and4 i_2212011(.A(n_268990188), .B(n_268890187), .C(n_268690185),
		 .D(n_268590184), .Z(to_acu100236[21]));
	notech_and4 i_2312012(.A(n_269590194), .B(n_269490193), .C(n_269290191),
		 .D(n_269190190), .Z(to_acu100236[22]));
	notech_and4 i_2412013(.A(n_270190200), .B(n_270090199), .C(n_269890197),
		 .D(n_269790196), .Z(to_acu100236[23]));
	notech_and4 i_2512014(.A(n_270790206), .B(n_270690205), .C(n_270490203),
		 .D(n_270390202), .Z(to_acu100236[24]));
	notech_and4 i_2612015(.A(n_271390212), .B(n_271290211), .C(n_271090209),
		 .D(n_270990208), .Z(to_acu100236[25]));
	notech_and4 i_2712016(.A(n_271990218), .B(n_271890217), .C(n_271690215),
		 .D(n_271590214), .Z(to_acu100236[26]));
	notech_and4 i_2812017(.A(n_272590224), .B(n_272490223), .C(n_272290221),
		 .D(n_272190220), .Z(to_acu100236[27]));
	notech_and4 i_2912018(.A(n_273190230), .B(n_273090229), .C(n_272890227),
		 .D(n_272790226), .Z(to_acu100236[28]));
	notech_and4 i_3012019(.A(n_273790236), .B(n_273690235), .C(n_273490233),
		 .D(n_273390232), .Z(to_acu100236[29]));
	notech_and4 i_3112020(.A(n_274390242), .B(n_274290241), .C(n_274090239),
		 .D(n_273990238), .Z(to_acu100236[30]));
	notech_and4 i_3212021(.A(n_274990248), .B(n_274890247), .C(n_274690245),
		 .D(n_274590244), .Z(to_acu100236[31]));
	notech_and4 i_112246(.A(n_277090269), .B(n_276890267), .C(n_276190260), 
		.D(n_275790256), .Z(to_acu100236[32]));
	notech_and4 i_212247(.A(n_277690275), .B(n_277590274), .C(n_277390272), 
		.D(n_277290271), .Z(to_acu100236[33]));
	notech_and4 i_312248(.A(n_278290281), .B(n_278190280), .C(n_277990278), 
		.D(n_277890277), .Z(to_acu100236[34]));
	notech_and4 i_412249(.A(n_278890287), .B(n_278790286), .C(n_278590284), 
		.D(n_278490283), .Z(to_acu100236[35]));
	notech_and4 i_512250(.A(n_279490293), .B(n_279390292), .C(n_279190290), 
		.D(n_279090289), .Z(to_acu100236[36]));
	notech_and4 i_612251(.A(n_280090299), .B(n_279990298), .C(n_279790296), 
		.D(n_279690295), .Z(to_acu100236[37]));
	notech_and4 i_712252(.A(n_280690305), .B(n_280590304), .C(n_280390302), 
		.D(n_280290301), .Z(to_acu100236[38]));
	notech_and4 i_812253(.A(n_281290311), .B(n_281190310), .C(n_280990308), 
		.D(n_280890307), .Z(to_acu100236[39]));
	notech_and4 i_912254(.A(n_281890317), .B(n_281790316), .C(n_281590314), 
		.D(n_281490313), .Z(to_acu100236[40]));
	notech_and4 i_1012255(.A(n_282490323), .B(n_282390322), .C(n_282190320),
		 .D(n_282090319), .Z(to_acu100236[41]));
	notech_and4 i_1112256(.A(n_283090329), .B(n_282990328), .C(n_282790326),
		 .D(n_282690325), .Z(to_acu100236[42]));
	notech_and4 i_1212257(.A(n_283690335), .B(n_283590334), .C(n_283390332),
		 .D(n_283290331), .Z(to_acu100236[43]));
	notech_and4 i_1312258(.A(n_284290341), .B(n_284190340), .C(n_283990338),
		 .D(n_283890337), .Z(to_acu100236[44]));
	notech_and4 i_1412259(.A(n_284890347), .B(n_284790346), .C(n_284590344),
		 .D(n_284490343), .Z(to_acu100236[45]));
	notech_and4 i_1512260(.A(n_285490353), .B(n_285390352), .C(n_285190350),
		 .D(n_285090349), .Z(to_acu100236[46]));
	notech_and4 i_1612261(.A(n_286090359), .B(n_285990358), .C(n_285790356),
		 .D(n_285690355), .Z(to_acu100236[47]));
	notech_and4 i_1712262(.A(n_286690365), .B(n_286590364), .C(n_286390362),
		 .D(n_286290361), .Z(to_acu100236[48]));
	notech_and4 i_1812263(.A(n_287290371), .B(n_287190370), .C(n_286990368),
		 .D(n_286890367), .Z(to_acu100236[49]));
	notech_and4 i_1912264(.A(n_287890377), .B(n_287790376), .C(n_287590374),
		 .D(n_287490373), .Z(to_acu100236[50]));
	notech_and4 i_2012265(.A(n_288490383), .B(n_288390382), .C(n_288190380),
		 .D(n_288090379), .Z(to_acu100236[51]));
	notech_and4 i_2112266(.A(n_289090389), .B(n_288990388), .C(n_288790386),
		 .D(n_288690385), .Z(to_acu100236[52]));
	notech_and4 i_2212267(.A(n_289690395), .B(n_289590394), .C(n_289390392),
		 .D(n_289290391), .Z(to_acu100236[53]));
	notech_and4 i_2312268(.A(n_290290401), .B(n_290190400), .C(n_289990398),
		 .D(n_289890397), .Z(to_acu100236[54]));
	notech_and4 i_2412269(.A(n_290890407), .B(n_290790406), .C(n_290590404),
		 .D(n_290490403), .Z(to_acu100236[55]));
	notech_and4 i_2512270(.A(n_291490413), .B(n_291390412), .C(n_291190410),
		 .D(n_291090409), .Z(to_acu100236[56]));
	notech_and4 i_2612271(.A(n_292090419), .B(n_291990418), .C(n_291790416),
		 .D(n_291690415), .Z(to_acu100236[57]));
	notech_and4 i_2712272(.A(n_292690425), .B(n_292590424), .C(n_292390422),
		 .D(n_292290421), .Z(to_acu100236[58]));
	notech_and4 i_2812273(.A(n_293290431), .B(n_293190430), .C(n_292990428),
		 .D(n_292890427), .Z(to_acu100236[59]));
	notech_and4 i_2912274(.A(n_293890437), .B(n_293790436), .C(n_293590434),
		 .D(n_293490433), .Z(to_acu100236[60]));
	notech_and4 i_3012275(.A(n_294490443), .B(n_294390442), .C(n_294190440),
		 .D(n_294090439), .Z(to_acu100236[61]));
	notech_and4 i_3112276(.A(n_295090449), .B(n_294990448), .C(n_294790446),
		 .D(n_294690445), .Z(to_acu100236[62]));
	notech_and4 i_3212277(.A(n_295690455), .B(n_295590454), .C(n_295390452),
		 .D(n_295290451), .Z(to_acu100236[63]));
	notech_nand2 i_118006(.A(n_295990458), .B(n_295890457), .Z(write_data_26
		[0]));
	notech_nand2 i_218007(.A(n_296190460), .B(n_296090459), .Z(write_data_26
		[1]));
	notech_nand2 i_418009(.A(n_296390462), .B(n_296290461), .Z(write_data_26
		[3]));
	notech_nand2 i_518010(.A(n_296590464), .B(n_296490463), .Z(write_data_26
		[4]));
	notech_nand2 i_618011(.A(n_296790466), .B(n_296690465), .Z(write_data_26
		[5]));
	notech_nand2 i_718012(.A(n_296990468), .B(n_296890467), .Z(write_data_26
		[6]));
	notech_nand2 i_818013(.A(n_297190470), .B(n_297090469), .Z(write_data_26
		[7]));
	notech_nand2 i_918014(.A(n_297390472), .B(n_297290471), .Z(write_data_26
		[8]));
	notech_nand2 i_1018015(.A(n_297590474), .B(n_297490473), .Z(write_data_26
		[9]));
	notech_nand2 i_1118016(.A(n_297790476), .B(n_297690475), .Z(write_data_26
		[10]));
	notech_nand2 i_1218017(.A(n_297990478), .B(n_297890477), .Z(write_data_26
		[11]));
	notech_nand2 i_1418019(.A(n_298190480), .B(n_298090479), .Z(write_data_26
		[13]));
	notech_nand2 i_1518020(.A(n_298390482), .B(n_298290481), .Z(write_data_26
		[14]));
	notech_nand2 i_1618021(.A(n_298690484), .B(n_298490483), .Z(write_data_26
		[15]));
	notech_nand2 i_1718022(.A(n_298890486), .B(n_298790485), .Z(write_data_26
		[16]));
	notech_nand2 i_2318028(.A(n_299090488), .B(n_298990487), .Z(write_data_26
		[22]));
	notech_nand2 i_2418029(.A(n_299290490), .B(n_299190489), .Z(write_data_26
		[23]));
	notech_nand2 i_2518030(.A(n_299490492), .B(n_299390491), .Z(write_data_26
		[24]));
	notech_nand2 i_2718032(.A(n_299690494), .B(n_299590493), .Z(write_data_26
		[26]));
	notech_nand2 i_2818033(.A(n_299890496), .B(n_299790495), .Z(write_data_26
		[27]));
	notech_nand2 i_2918034(.A(n_300090498), .B(n_299990497), .Z(write_data_26
		[28]));
	notech_nand2 i_3018035(.A(n_300290500), .B(n_300190499), .Z(write_data_26
		[29]));
	notech_nand2 i_3118036(.A(n_300490502), .B(n_300390501), .Z(write_data_26
		[30]));
	notech_nand2 i_3218037(.A(n_300690504), .B(n_300590503), .Z(write_data_26
		[31]));
	notech_nand2 i_118134(.A(n_300890506), .B(n_300790505), .Z(write_data_27
		[0]));
	notech_nand2 i_218135(.A(n_301090508), .B(n_300990507), .Z(write_data_27
		[1]));
	notech_nand2 i_418137(.A(n_301290510), .B(n_301190509), .Z(write_data_27
		[3]));
	notech_nand2 i_518138(.A(n_301490512), .B(n_301390511), .Z(write_data_27
		[4]));
	notech_nand2 i_718140(.A(n_301690514), .B(n_301590513), .Z(write_data_27
		[6]));
	notech_nand2 i_818141(.A(n_301890516), .B(n_301790515), .Z(write_data_27
		[7]));
	notech_nand2 i_918142(.A(n_302090518), .B(n_301990517), .Z(write_data_27
		[8]));
	notech_nand2 i_1018143(.A(n_302290520), .B(n_302190519), .Z(write_data_27
		[9]));
	notech_nand2 i_1118144(.A(n_302490522), .B(n_302390521), .Z(write_data_27
		[10]));
	notech_nand2 i_1218145(.A(n_302690524), .B(n_302590523), .Z(write_data_27
		[11]));
	notech_nand2 i_1318146(.A(n_302890526), .B(n_302790525), .Z(write_data_27
		[12]));
	notech_nand2 i_1418147(.A(n_303090528), .B(n_302990527), .Z(write_data_27
		[13]));
	notech_nand2 i_1518148(.A(n_303290530), .B(n_303190529), .Z(write_data_27
		[14]));
	notech_nand2 i_1618149(.A(n_303490532), .B(n_303390531), .Z(write_data_27
		[15]));
	notech_nand2 i_1718150(.A(n_303690534), .B(n_303590533), .Z(write_data_27
		[16]));
	notech_nand2 i_1818151(.A(n_303890536), .B(n_303790535), .Z(write_data_27
		[17]));
	notech_nand2 i_1918152(.A(n_304090538), .B(n_303990537), .Z(write_data_27
		[18]));
	notech_nand2 i_2018153(.A(n_304290540), .B(n_304190539), .Z(write_data_27
		[19]));
	notech_nand2 i_2118154(.A(n_304490542), .B(n_304390541), .Z(write_data_27
		[20]));
	notech_nand2 i_2218155(.A(n_304690544), .B(n_304590543), .Z(write_data_27
		[21]));
	notech_nand2 i_2318156(.A(n_304890546), .B(n_304790545), .Z(write_data_27
		[22]));
	notech_nand2 i_2418157(.A(n_305090548), .B(n_304990547), .Z(write_data_27
		[23]));
	notech_nand2 i_2518158(.A(n_305290550), .B(n_305190549), .Z(write_data_27
		[24]));
	notech_nand2 i_2618159(.A(n_305490552), .B(n_305390551), .Z(write_data_27
		[25]));
	notech_nand2 i_2718160(.A(n_305690554), .B(n_305590553), .Z(write_data_27
		[26]));
	notech_nand2 i_2818161(.A(n_305890556), .B(n_305790555), .Z(write_data_27
		[27]));
	notech_nand2 i_2918162(.A(n_306090558), .B(n_305990557), .Z(write_data_27
		[28]));
	notech_nand2 i_3018163(.A(n_306290560), .B(n_306190559), .Z(write_data_27
		[29]));
	notech_nand2 i_3118164(.A(n_306490562), .B(n_306390561), .Z(write_data_27
		[30]));
	notech_nand2 i_3218165(.A(n_306690564), .B(n_306590563), .Z(write_data_27
		[31]));
	notech_nand2 i_318264(.A(n_306890566), .B(n_306790565), .Z(write_data_28
		[2]));
	notech_nand2 i_518266(.A(n_307090568), .B(n_306990567), .Z(write_data_28
		[4]));
	notech_nand2 i_618267(.A(n_307290570), .B(n_307190569), .Z(write_data_28
		[5]));
	notech_nand2 i_718268(.A(n_307490572), .B(n_307390571), .Z(write_data_28
		[6]));
	notech_nand2 i_818269(.A(n_307690574), .B(n_307590573), .Z(write_data_28
		[7]));
	notech_nand2 i_1018271(.A(n_307890576), .B(n_307790575), .Z(write_data_28
		[9]));
	notech_nand2 i_1118272(.A(n_308090578), .B(n_307990577), .Z(write_data_28
		[10]));
	notech_nand2 i_3218293(.A(n_308290580), .B(n_308190579), .Z(write_data_28
		[31]));
	notech_nand2 i_118390(.A(n_308790585), .B(n_308490582), .Z(write_data_29
		[0]));
	notech_nand2 i_218391(.A(n_308990587), .B(n_308890586), .Z(write_data_29
		[1]));
	notech_nand2 i_318392(.A(n_309190589), .B(n_309090588), .Z(write_data_29
		[2]));
	notech_nand2 i_418393(.A(n_309390591), .B(n_309290590), .Z(write_data_29
		[3]));
	notech_nand2 i_518394(.A(n_309590593), .B(n_309490592), .Z(write_data_29
		[4]));
	notech_nand2 i_618395(.A(n_309790595), .B(n_309690594), .Z(write_data_29
		[5]));
	notech_nand2 i_718396(.A(n_309990597), .B(n_309890596), .Z(write_data_29
		[6]));
	notech_nand2 i_818397(.A(n_310190599), .B(n_310090598), .Z(write_data_29
		[7]));
	notech_nand2 i_918398(.A(n_310390601), .B(n_310290600), .Z(write_data_29
		[8]));
	notech_nand2 i_1018399(.A(n_310590603), .B(n_310490602), .Z(write_data_29
		[9]));
	notech_nand2 i_1118400(.A(n_310790605), .B(n_310690604), .Z(write_data_29
		[10]));
	notech_nand2 i_1218401(.A(n_310990607), .B(n_310890606), .Z(write_data_29
		[11]));
	notech_nand2 i_1318402(.A(n_311190609), .B(n_311090608), .Z(write_data_29
		[12]));
	notech_nand2 i_1418403(.A(n_311390611), .B(n_311290610), .Z(write_data_29
		[13]));
	notech_nand2 i_1518404(.A(n_311590613), .B(n_311490612), .Z(write_data_29
		[14]));
	notech_nand2 i_1618405(.A(n_311790615), .B(n_311690614), .Z(write_data_29
		[15]));
	notech_nand2 i_1718406(.A(n_311990617), .B(n_311890616), .Z(write_data_29
		[16]));
	notech_nand2 i_1818407(.A(n_312190619), .B(n_312090618), .Z(write_data_29
		[17]));
	notech_nand2 i_1918408(.A(n_312390621), .B(n_312290620), .Z(write_data_29
		[18]));
	notech_nand2 i_2018409(.A(n_312590623), .B(n_312490622), .Z(write_data_29
		[19]));
	notech_nand2 i_2318412(.A(n_312790625), .B(n_312690624), .Z(write_data_29
		[22]));
	notech_nand2 i_2418413(.A(n_312990627), .B(n_312890626), .Z(write_data_29
		[23]));
	notech_nand2 i_2518414(.A(n_313190629), .B(n_313090628), .Z(write_data_29
		[24]));
	notech_nand2 i_2618415(.A(n_313390631), .B(n_313290630), .Z(write_data_29
		[25]));
	notech_nand2 i_2718416(.A(n_313590633), .B(n_313490632), .Z(write_data_29
		[26]));
	notech_nand2 i_2818417(.A(n_313790635), .B(n_313690634), .Z(write_data_29
		[27]));
	notech_nand2 i_2918418(.A(n_313990637), .B(n_313890636), .Z(write_data_29
		[28]));
	notech_nand2 i_3018419(.A(n_314190639), .B(n_314090638), .Z(write_data_29
		[29]));
	notech_nand2 i_3118420(.A(n_314390641), .B(n_314290640), .Z(write_data_29
		[30]));
	notech_nand2 i_3218421(.A(n_314590643), .B(n_314490642), .Z(write_data_29
		[31]));
	notech_nand2 i_118774(.A(n_315390651), .B(n_315090648), .Z(write_data_32
		[0]));
	notech_nand2 i_218775(.A(n_315590653), .B(n_315490652), .Z(write_data_32
		[1]));
	notech_nand2 i_318776(.A(n_315790655), .B(n_315690654), .Z(write_data_32
		[2]));
	notech_nand2 i_418777(.A(n_315990657), .B(n_315890656), .Z(write_data_32
		[3]));
	notech_nand2 i_518778(.A(n_316190659), .B(n_316090658), .Z(write_data_32
		[4]));
	notech_nand2 i_618779(.A(n_316390661), .B(n_316290660), .Z(write_data_32
		[5]));
	notech_nand2 i_718780(.A(n_316590663), .B(n_316490662), .Z(write_data_32
		[6]));
	notech_nand2 i_818781(.A(n_316790665), .B(n_316690664), .Z(write_data_32
		[7]));
	notech_nand2 i_918782(.A(n_316990667), .B(n_316890666), .Z(write_data_32
		[8]));
	notech_nand2 i_1018783(.A(n_317190669), .B(n_317090668), .Z(write_data_32
		[9]));
	notech_nand2 i_1118784(.A(n_317390671), .B(n_317290670), .Z(write_data_32
		[10]));
	notech_nand2 i_1218785(.A(n_317590673), .B(n_317490672), .Z(write_data_32
		[11]));
	notech_nand2 i_1318786(.A(n_317790675), .B(n_317690674), .Z(write_data_32
		[12]));
	notech_nand2 i_1418787(.A(n_317990677), .B(n_317890676), .Z(write_data_32
		[13]));
	notech_nand2 i_1518788(.A(n_318190679), .B(n_318090678), .Z(write_data_32
		[14]));
	notech_nand2 i_1618789(.A(n_318390681), .B(n_318290680), .Z(write_data_32
		[15]));
	notech_nand2 i_1718790(.A(n_318590683), .B(n_318490682), .Z(write_data_32
		[16]));
	notech_nand2 i_1818791(.A(n_318790685), .B(n_318690684), .Z(write_data_32
		[17]));
	notech_nand2 i_1918792(.A(n_318990687), .B(n_318890686), .Z(write_data_32
		[18]));
	notech_nand2 i_2018793(.A(n_319190689), .B(n_319090688), .Z(write_data_32
		[19]));
	notech_nand2 i_2118794(.A(n_319390691), .B(n_319290690), .Z(write_data_32
		[20]));
	notech_nand2 i_2218795(.A(n_319590693), .B(n_319490692), .Z(write_data_32
		[21]));
	notech_nand2 i_2318796(.A(n_319790695), .B(n_319690694), .Z(write_data_32
		[22]));
	notech_nand2 i_2418797(.A(n_319990697), .B(n_319890696), .Z(write_data_32
		[23]));
	notech_nand2 i_2518798(.A(n_320190699), .B(n_320090698), .Z(write_data_32
		[24]));
	notech_nand2 i_2618799(.A(n_320390701), .B(n_320290700), .Z(write_data_32
		[25]));
	notech_nand2 i_2718800(.A(n_320590703), .B(n_320490702), .Z(write_data_32
		[26]));
	notech_nand2 i_2818801(.A(n_320790705), .B(n_320690704), .Z(write_data_32
		[27]));
	notech_nand2 i_2918802(.A(n_320990707), .B(n_320890706), .Z(write_data_32
		[28]));
	notech_nand2 i_3018803(.A(n_321190709), .B(n_321090708), .Z(write_data_32
		[29]));
	notech_nand2 i_3118804(.A(n_321390711), .B(n_321290710), .Z(write_data_32
		[30]));
	notech_nand2 i_3218805(.A(n_321590713), .B(n_321490712), .Z(write_data_32
		[31]));
	notech_nand2 i_1529(.A(n_2825), .B(n_2838), .Z(n_2839));
	notech_and4 i_727966(.A(n_2826), .B(n_2835), .C(n_2645), .D(n_2632), .Z(n_2838
		));
	notech_or4 i_17836(.A(n_2896), .B(n_3790), .C(n_27069), .D(n_29655), .Z(n_327690774
		));
	notech_or4 i_17838(.A(n_60863), .B(n_61109), .C(n_69641311), .D(n_62870)
		, .Z(n_327790775));
	notech_or4 i_17839(.A(n_69641311), .B(n_61109), .C(n_62870), .D(n_59429)
		, .Z(n_327890776));
	notech_or4 i_17841(.A(n_69641311), .B(n_61109), .C(n_60874), .D(n_59429)
		, .Z(n_327990777));
	notech_or4 i_19238(.A(n_32443), .B(n_27994), .C(n_10157), .D(n_323190729
		), .Z(n_328090778));
	notech_nao3 i_19955(.A(n_60138), .B(n_60312), .C(n_57966), .Z(n_328190779
		));
	notech_or4 i_21347(.A(n_60863), .B(n_61109), .C(n_58220), .D(n_60845), .Z
		(n_328290780));
	notech_or4 i_26925(.A(n_61133), .B(n_60212), .C(n_29793), .D(n_268643294
		), .Z(n_328390781));
	notech_and4 i_17484(.A(n_62868), .B(n_32730), .C(n_55820), .D(n_2478), .Z
		(n_328490782));
	notech_ao3 i_18417(.A(tcmp_arithbox), .B(n_60312), .C(n_58072), .Z(n_328590783
		));
	notech_nand2 i_50248(.A(n_323590733), .B(n_58691), .Z(n_16532));
	notech_nand2 i_1417891(.A(n_325290750), .B(n_325190749), .Z(write_data_25
		[13]));
	notech_nand2 i_618139(.A(n_325490752), .B(n_325390751), .Z(write_data_27
		[5]));
	notech_nand2 i_2918674(.A(n_325990757), .B(n_325890756), .Z(write_data_31
		[28]));
	notech_ao3 i_18802(.A(n_2885), .B(n_326090758), .C(n_61151), .Z(n_328690784
		));
	notech_nand2 i_1918024(.A(n_327390771), .B(n_327290770), .Z(write_data_26
		[18]));
	notech_ao3 i_371(.A(n_2833), .B(n_2832), .C(n_2642), .Z(n_2835));
	notech_nand2 i_52786(.A(n_327590773), .B(n_58691), .Z(n_20021));
	notech_nand2 i_49752(.A(n_327490772), .B(n_58691), .Z(n_15633));
	notech_ao4 i_367(.A(n_275591872), .B(n_29133), .C(n_29648), .D(n_273591890
		), .Z(n_2833));
	notech_and4 i_368(.A(n_2829), .B(n_2828), .C(n_2827), .D(n_264191922), .Z
		(n_2832));
	notech_ao4 i_362(.A(n_275791870), .B(n_29124), .C(n_29173), .D(n_273791888
		), .Z(n_2829));
	notech_ao4 i_360(.A(n_274891879), .B(n_29157), .C(n_274491883), .D(n_29165
		), .Z(n_2828));
	notech_ao4 i_364(.A(n_275191876), .B(n_29141), .C(n_29666), .D(n_272791898
		), .Z(n_2827));
	notech_ao4 i_370(.A(n_29665), .B(n_273191894), .C(n_275291875), .D(n_29149
		), .Z(n_2826));
	notech_and4 i_527964(.A(n_2813), .B(n_2822), .C(n_2631), .D(n_2618), .Z(n_2825
		));
	notech_ao3 i_342(.A(n_2820), .B(n_2819), .C(n_2628), .Z(n_2822));
	notech_ao4 i_336(.A(n_275591872), .B(n_29131), .C(n_273591890), .D(n_29647
		), .Z(n_2820));
	notech_and4 i_338(.A(n_2816), .B(n_2815), .C(n_2814), .D(n_2627), .Z(n_2819
		));
	notech_ao4 i_332(.A(n_275791870), .B(n_29122), .C(n_29171), .D(n_273791888
		), .Z(n_2816));
	notech_ao4 i_330(.A(n_274891879), .B(n_29155), .C(n_274491883), .D(n_29163
		), .Z(n_2815));
	notech_ao4 i_333(.A(n_275191876), .B(n_29139), .C(n_272791898), .D(n_29634
		), .Z(n_2814));
	notech_ao4 i_341(.A(n_273191894), .B(n_29633), .C(n_275291875), .D(n_29147
		), .Z(n_2813));
	notech_ao3 i_255(.A(n_2808), .B(n_2807), .C(n_2586), .Z(n_2810));
	notech_ao4 i_250(.A(n_275591872), .B(n_29130), .C(n_273591890), .D(n_29646
		), .Z(n_2808));
	notech_and4 i_251(.A(n_2804), .B(n_2803), .C(n_2802), .D(n_2585), .Z(n_2807
		));
	notech_ao4 i_245(.A(n_275791870), .B(n_29121), .C(n_29170), .D(n_273791888
		), .Z(n_2804));
	notech_ao4 i_244(.A(n_274891879), .B(n_29154), .C(n_274491883), .D(n_29162
		), .Z(n_2803));
	notech_ao4 i_246(.A(n_275191876), .B(n_29138), .C(n_272791898), .D(n_29640
		), .Z(n_2802));
	notech_ao4 i_254(.A(n_273191894), .B(n_29639), .C(n_275291875), .D(n_29146
		), .Z(n_2801));
	notech_ao3 i_222(.A(n_2796), .B(n_2795), .C(n_2572), .Z(n_2798));
	notech_ao4 i_216(.A(n_275591872), .B(n_29127), .C(n_273591890), .D(n_29645
		), .Z(n_2796));
	notech_and4 i_217(.A(n_2792), .B(n_2791), .C(n_2790), .D(n_2571), .Z(n_2795
		));
	notech_ao4 i_212(.A(n_275791870), .B(n_29118), .C(n_29167), .D(n_273791888
		), .Z(n_2792));
	notech_ao4 i_211(.A(n_274891879), .B(n_29151), .C(n_274491883), .D(n_29159
		), .Z(n_2791));
	notech_ao4 i_213(.A(n_275191876), .B(n_29135), .C(n_29642), .D(n_272791898
		), .Z(n_2790));
	notech_ao4 i_221(.A(n_273191894), .B(n_29641), .C(n_275291875), .D(n_29143
		), .Z(n_2789));
	notech_nand3 i_194(.A(n_2777), .B(n_2786), .C(n_2560), .Z(n_2788));
	notech_ao3 i_192(.A(n_2784), .B(n_2783), .C(n_2557), .Z(n_2786));
	notech_ao4 i_188(.A(n_275591872), .B(n_29129), .C(n_273591890), .D(n_29644
		), .Z(n_2784));
	notech_and4 i_189(.A(n_2780), .B(n_2779), .C(n_2778), .D(n_2556), .Z(n_2783
		));
	notech_ao4 i_184(.A(n_275791870), .B(n_29120), .C(n_29169), .D(n_273791888
		), .Z(n_2780));
	notech_ao4 i_183(.A(n_274891879), .B(n_29153), .C(n_274491883), .D(n_29161
		), .Z(n_2779));
	notech_ao4 i_185(.A(n_275191876), .B(n_29137), .C(n_29668), .D(n_272791898
		), .Z(n_2778));
	notech_ao4 i_191(.A(n_273191894), .B(n_29667), .C(n_275291875), .D(n_29145
		), .Z(n_2777));
	notech_ao3 i_165(.A(n_2772), .B(n_2771), .C(n_2542), .Z(n_2774));
	notech_ao4 i_158(.A(n_275591872), .B(n_29128), .C(n_273591890), .D(n_29643
		), .Z(n_2772));
	notech_and4 i_159(.A(n_2768), .B(n_276791860), .C(n_276691861), .D(n_2541
		), .Z(n_2771));
	notech_and2 i_17941(.A(pt_fault), .B(n_30635), .Z(n_24991034));
	notech_and2 i_27104(.A(had_lgjmp), .B(\nbus_14522[31] ), .Z(pg_en));
	notech_ao4 i_91970130(.A(n_154379047), .B(n_27767), .C(n_27107), .D(n_27424
		), .Z(n_34391128));
	notech_ao4 i_91870131(.A(n_154179045), .B(n_56019), .C(n_154279046), .D(n_27729
		), .Z(n_34491129));
	notech_ao4 i_91770132(.A(n_154379047), .B(n_27768), .C(n_27107), .D(n_27426
		), .Z(n_34591130));
	notech_ao4 i_91670133(.A(n_154179045), .B(n_29733), .C(n_154279046), .D(n_27730
		), .Z(n_34691131));
	notech_ao4 i_91570134(.A(n_154379047), .B(n_27769), .C(n_27107), .D(n_27428
		), .Z(n_34791132));
	notech_ao4 i_91470135(.A(n_154179045), .B(n_29728), .C(n_154279046), .D(n_27731
		), .Z(n_34891133));
	notech_ao4 i_91370136(.A(n_154379047), .B(n_27770), .C(n_27107), .D(n_27430
		), .Z(n_34991134));
	notech_ao4 i_91270137(.A(n_154179045), .B(n_56055), .C(n_154279046), .D(n_27732
		), .Z(n_35091135));
	notech_ao4 i_91170138(.A(n_154379047), .B(n_27771), .C(n_27107), .D(n_27432
		), .Z(n_35191136));
	notech_ao4 i_91070139(.A(n_154179045), .B(n_29651), .C(n_154279046), .D(n_27733
		), .Z(n_35291137));
	notech_ao4 i_90970140(.A(n_154379047), .B(n_27773), .C(n_27107), .D(n_27434
		), .Z(n_35391138));
	notech_ao4 i_90870141(.A(n_154179045), .B(n_29723), .C(n_154279046), .D(n_27734
		), .Z(n_35491139));
	notech_ao4 i_90770142(.A(n_154379047), .B(n_27774), .C(n_27107), .D(n_27437
		), .Z(n_35591140));
	notech_ao4 i_90670143(.A(n_154179045), .B(n_29614), .C(n_154279046), .D(n_27735
		), .Z(n_35691141));
	notech_ao4 i_90570144(.A(n_54093), .B(n_27775), .C(n_54431), .D(n_27439)
		, .Z(n_35791142));
	notech_ao4 i_90470145(.A(n_54113), .B(n_29787), .C(n_54104), .D(n_27737)
		, .Z(n_35891143));
	notech_ao4 i_90370146(.A(n_54093), .B(n_27776), .C(n_54431), .D(n_27441)
		, .Z(n_35991144));
	notech_ao4 i_90270147(.A(n_54113), .B(n_56127), .C(n_54104), .D(n_27738)
		, .Z(n_36091145));
	notech_ao4 i_89370156(.A(n_54093), .B(n_27786), .C(n_54431), .D(n_27453)
		, .Z(n_36191146));
	notech_ao4 i_89270157(.A(n_54113), .B(n_56266), .C(n_54104), .D(n_27744)
		, .Z(n_36291147));
	notech_ao4 i_89170158(.A(n_54093), .B(n_27787), .C(n_54431), .D(n_27455)
		, .Z(n_36391148));
	notech_ao4 i_89070159(.A(n_54113), .B(n_29710), .C(n_54104), .D(n_27745)
		, .Z(n_36491149));
	notech_ao4 i_88970160(.A(n_54093), .B(n_27788), .C(n_54431), .D(n_27457)
		, .Z(n_36591150));
	notech_ao4 i_88870161(.A(n_54113), .B(n_29772), .C(n_54104), .D(n_27747)
		, .Z(n_36691151));
	notech_ao4 i_88770162(.A(n_54093), .B(n_27789), .C(n_54431), .D(n_27459)
		, .Z(n_36791152));
	notech_ao4 i_88670163(.A(n_54113), .B(n_29711), .C(n_54104), .D(n_27748)
		, .Z(n_36891153));
	notech_ao4 i_88570164(.A(n_54093), .B(n_27790), .C(n_54431), .D(n_27461)
		, .Z(n_36991154));
	notech_ao4 i_88470165(.A(n_54113), .B(n_29773), .C(n_54104), .D(n_27749)
		, .Z(n_37091155));
	notech_ao4 i_88370166(.A(n_54093), .B(n_27791), .C(n_54431), .D(n_27463)
		, .Z(n_37191156));
	notech_ao4 i_88270167(.A(n_54113), .B(n_29775), .C(n_54104), .D(n_27750)
		, .Z(n_37291157));
	notech_ao4 i_88170168(.A(n_54093), .B(n_27792), .C(n_54431), .D(n_27465)
		, .Z(n_37391158));
	notech_ao4 i_88070169(.A(n_54113), .B(n_29681), .C(n_54104), .D(n_27751)
		, .Z(n_37491159));
	notech_ao4 i_87970170(.A(n_54093), .B(n_27793), .C(n_54431), .D(n_27469)
		, .Z(n_37591160));
	notech_ao4 i_87870171(.A(n_54113), .B(n_29708), .C(n_54104), .D(n_27752)
		, .Z(n_37691161));
	notech_ao4 i_87770172(.A(n_54093), .B(n_27794), .C(n_27107), .D(n_27471)
		, .Z(n_37791162));
	notech_ao4 i_87670173(.A(n_54113), .B(n_29765), .C(n_154279046), .D(n_27755
		), .Z(n_37891163));
	notech_ao4 i_87570174(.A(n_54093), .B(n_27795), .C(n_54431), .D(n_27473)
		, .Z(n_37991164));
	notech_ao4 i_87470175(.A(n_54113), .B(n_29769), .C(n_54104), .D(n_27756)
		, .Z(n_38091165));
	notech_ao4 i_87370176(.A(n_54093), .B(n_27797), .C(n_54431), .D(n_27475)
		, .Z(n_38191166));
	notech_ao4 i_87270177(.A(n_54113), .B(n_29770), .C(n_54104), .D(n_27758)
		, .Z(n_38291167));
	notech_ao4 i_87170178(.A(n_54093), .B(n_27798), .C(n_54431), .D(n_27477)
		, .Z(n_38391168));
	notech_ao4 i_87070179(.A(n_54113), .B(n_29660), .C(n_54104), .D(n_27759)
		, .Z(n_38491169));
	notech_ao4 i_86970180(.A(n_54093), .B(n_27799), .C(n_54431), .D(n_27479)
		, .Z(n_38591170));
	notech_ao4 i_86870181(.A(n_54113), .B(n_29661), .C(n_54104), .D(n_27760)
		, .Z(n_38691171));
	notech_ao4 i_86770182(.A(n_54093), .B(n_27800), .C(n_54431), .D(n_27481)
		, .Z(n_38791172));
	notech_ao4 i_86670183(.A(n_54113), .B(n_29662), .C(n_54104), .D(n_27762)
		, .Z(n_38891173));
	notech_xor2 i_7767324(.A(n_32420), .B(all_cnt[2]), .Z(n_38991174));
	notech_xor2 i_7867323(.A(n_32421), .B(all_cnt[3]), .Z(n_39091175));
	notech_ao4 i_222479(.A(n_27853), .B(n_45891243), .C(n_60312), .D(n_3913)
		, .Z(n_12888));
	notech_ao4 i_6327542(.A(n_55514), .B(n_29537), .C(n_55498), .D(n_29535),
		 .Z(n_13681));
	notech_ao4 i_6227541(.A(n_55514), .B(n_29536), .C(n_55498), .D(n_29534),
		 .Z(n_13676));
	notech_ao4 i_6127540(.A(n_55519), .B(n_29535), .C(n_55498), .D(n_29533),
		 .Z(n_13671));
	notech_ao4 i_6027539(.A(n_55514), .B(n_29534), .C(n_55498), .D(n_29532),
		 .Z(n_13666));
	notech_ao4 i_5927538(.A(n_55514), .B(n_29533), .C(n_55498), .D(n_29531),
		 .Z(n_13661));
	notech_ao4 i_5827537(.A(n_55514), .B(n_29532), .C(n_55498), .D(n_29530),
		 .Z(n_13656));
	notech_ao4 i_5727536(.A(n_55514), .B(n_29531), .C(n_55498), .D(n_29529),
		 .Z(n_13651));
	notech_ao4 i_5627535(.A(n_55514), .B(n_29530), .C(n_55498), .D(n_29528),
		 .Z(n_13646));
	notech_ao4 i_5527534(.A(n_55514), .B(n_29529), .C(n_55498), .D(n_29527),
		 .Z(n_13641));
	notech_ao4 i_5427533(.A(n_55514), .B(n_29528), .C(n_55498), .D(n_29526),
		 .Z(n_13636));
	notech_ao4 i_5327532(.A(n_55514), .B(n_29527), .C(n_55498), .D(n_29525),
		 .Z(n_13631));
	notech_ao4 i_5227531(.A(n_55514), .B(n_29526), .C(n_55498), .D(n_29524),
		 .Z(n_13626));
	notech_ao4 i_5127530(.A(n_55514), .B(n_29525), .C(n_55503), .D(n_29523),
		 .Z(n_13621));
	notech_ao4 i_5027529(.A(n_55519), .B(n_29524), .C(n_55503), .D(n_29522),
		 .Z(n_13616));
	notech_ao4 i_4927528(.A(n_55519), .B(n_29523), .C(n_55503), .D(n_29521),
		 .Z(n_13611));
	notech_ao4 i_4827527(.A(n_55519), .B(n_29522), .C(n_55503), .D(n_29520),
		 .Z(n_13606));
	notech_ao4 i_4727526(.A(n_55519), .B(n_29521), .C(n_55503), .D(n_29519),
		 .Z(n_13601));
	notech_ao4 i_4627525(.A(n_55519), .B(n_29520), .C(n_55503), .D(n_29518),
		 .Z(n_13596));
	notech_ao4 i_4527524(.A(n_55524), .B(n_29519), .C(n_55503), .D(n_29517),
		 .Z(n_13591));
	notech_ao4 i_4427523(.A(n_55524), .B(n_29518), .C(n_55503), .D(n_29516),
		 .Z(n_13586));
	notech_ao4 i_4327522(.A(n_55519), .B(n_29517), .C(n_55503), .D(n_29515),
		 .Z(n_13581));
	notech_ao4 i_4227521(.A(n_55519), .B(n_29516), .C(n_55503), .D(n_29514),
		 .Z(n_13576));
	notech_ao4 i_4127520(.A(n_55519), .B(n_29515), .C(n_55503), .D(n_29513),
		 .Z(n_13571));
	notech_ao4 i_4027519(.A(n_55519), .B(n_29514), .C(n_55503), .D(n_29512),
		 .Z(n_13566));
	notech_ao4 i_3927518(.A(n_55519), .B(n_29513), .C(n_55503), .D(n_29511),
		 .Z(n_13561));
	notech_ao4 i_3827517(.A(n_55519), .B(n_29512), .C(n_55503), .D(n_29510),
		 .Z(n_13556));
	notech_ao4 i_3727516(.A(n_55519), .B(n_29511), .C(n_55503), .D(n_29509),
		 .Z(n_13551));
	notech_ao4 i_3627515(.A(n_55519), .B(n_29510), .C(n_55503), .D(n_29508),
		 .Z(n_13546));
	notech_ao4 i_3527514(.A(n_55519), .B(n_29509), .C(n_55503), .D(n_29507),
		 .Z(n_13541));
	notech_ao4 i_3427513(.A(n_55519), .B(n_29508), .C(n_55503), .D(n_29506),
		 .Z(n_13536));
	notech_ao3 i_24299(.A(n_60378), .B(opb[0]), .C(n_61151), .Z(n_45791242)
		);
	notech_ao4 i_154(.A(n_275791870), .B(n_29119), .C(n_29168), .D(n_273791888
		), .Z(n_2768));
	notech_ao4 i_153(.A(n_274891879), .B(n_29152), .C(n_274491883), .D(n_29160
		), .Z(n_276791860));
	notech_ao4 i_155(.A(n_275191876), .B(n_29136), .C(n_272791898), .D(n_29631
		), .Z(n_276691861));
	notech_ao4 i_164(.A(n_273191894), .B(n_29628), .C(n_275291875), .D(n_29144
		), .Z(n_276591862));
	notech_and4 i_64(.A(n_274191886), .B(n_2740), .C(n_276191866), .D(n_273891887
		), .Z(n_276391864));
	notech_and4 i_49(.A(n_275291875), .B(n_275191876), .C(n_274991878), .D(n_275991868
		), .Z(n_276191866));
	notech_and3 i_44(.A(n_275791870), .B(n_275591872), .C(n_275491873), .Z(n_275991868
		));
	notech_or4 i_50455(.A(vliw_pc[1]), .B(vliw_pc[3]), .C(n_272591900), .D(n_27722
		), .Z(n_275791870));
	notech_or4 i_50454(.A(vliw_pc[3]), .B(n_272591900), .C(n_27723), .D(vliw_pc
		[0]), .Z(n_275591872));
	notech_or4 i_50457(.A(vliw_pc[4]), .B(vliw_pc[2]), .C(vliw_pc[0]), .D(n_27493
		), .Z(n_275491873));
	notech_or4 i_1680219(.A(vliw_pc[4]), .B(vliw_pc[0]), .C(n_27724), .D(n_27493
		), .Z(n_275291875));
	notech_or4 i_50452(.A(vliw_pc[3]), .B(n_272591900), .C(n_27722), .D(n_27723
		), .Z(n_275191876));
	notech_and2 i_1380218(.A(n_274891879), .B(n_274491883), .Z(n_274991878)
		);
	notech_or4 i_50449(.A(vliw_pc[4]), .B(n_27722), .C(n_27724), .D(n_27493)
		, .Z(n_274891879));
	notech_nor2 i_2007(.A(vliw_pc[3]), .B(vliw_pc[1]), .Z(n_274591882));
	notech_or4 i_50448(.A(vliw_pc[3]), .B(n_27723), .C(n_27724), .D(n_272891897
		), .Z(n_274491883));
	notech_nao3 i_1780216(.A(n_273091895), .B(n_27722), .C(n_272591900), .Z(n_274191886
		));
	notech_nand3 i_50446(.A(n_32843), .B(n_2739), .C(vliw_pc[2]), .Z(n_2740)
		);
	notech_nor2 i_125(.A(vliw_pc[4]), .B(vliw_pc[3]), .Z(n_2739));
	notech_and2 i_1580215(.A(n_273591890), .B(n_273791888), .Z(n_273891887)
		);
	notech_nao3 i_50443(.A(n_273091895), .B(vliw_pc[0]), .C(n_272591900), .Z
		(n_273791888));
	notech_mux2 i_112278(.S(n_60537), .A(n_6053), .B(regs_14[0]), .Z(pc_out[
		0]));
	notech_mux2 i_212279(.S(n_60542), .A(n_6054), .B(regs_14[1]), .Z(pc_out[
		1]));
	notech_mux2 i_312280(.S(n_60537), .A(n_6055), .B(regs_14[2]), .Z(pc_out[
		2]));
	notech_mux2 i_412281(.S(n_60537), .A(n_6056), .B(regs_14[3]), .Z(pc_out[
		3]));
	notech_mux2 i_512282(.S(n_60537), .A(n_6057), .B(regs_14[4]), .Z(pc_out[
		4]));
	notech_mux2 i_612283(.S(n_60537), .A(n_6058), .B(regs_14[5]), .Z(pc_out[
		5]));
	notech_mux2 i_712284(.S(n_60537), .A(n_6059), .B(regs_14[6]), .Z(pc_out[
		6]));
	notech_mux2 i_812285(.S(n_60537), .A(n_6060), .B(regs_14[7]), .Z(pc_out[
		7]));
	notech_mux2 i_912286(.S(n_60537), .A(n_6061), .B(regs_14[8]), .Z(pc_out[
		8]));
	notech_mux2 i_1012287(.S(n_60537), .A(n_6062), .B(regs_14[9]), .Z(pc_out
		[9]));
	notech_mux2 i_1112288(.S(n_60537), .A(n_6063), .B(regs_14[10]), .Z(pc_out
		[10]));
	notech_mux2 i_1212289(.S(n_60542), .A(n_6064), .B(regs_14[11]), .Z(pc_out
		[11]));
	notech_mux2 i_1312290(.S(n_60542), .A(n_6065), .B(regs_14[12]), .Z(pc_out
		[12]));
	notech_mux2 i_1412291(.S(n_60542), .A(n_6066), .B(regs_14[13]), .Z(pc_out
		[13]));
	notech_mux2 i_1512292(.S(n_60542), .A(n_6067), .B(regs_14[14]), .Z(pc_out
		[14]));
	notech_mux2 i_1612293(.S(n_60542), .A(n_6068), .B(regs_14[15]), .Z(pc_out
		[15]));
	notech_mux2 i_1712294(.S(n_60542), .A(n_6069), .B(regs_14[16]), .Z(pc_out
		[16]));
	notech_mux2 i_1812295(.S(n_60548), .A(n_6070), .B(regs_14[17]), .Z(pc_out
		[17]));
	notech_mux2 i_1912296(.S(n_60542), .A(n_6071), .B(regs_14[18]), .Z(pc_out
		[18]));
	notech_mux2 i_2012297(.S(n_60542), .A(n_6072), .B(regs_14[19]), .Z(pc_out
		[19]));
	notech_mux2 i_2212299(.S(n_60542), .A(n_6074), .B(regs_14[21]), .Z(pc_out
		[21]));
	notech_mux2 i_2712304(.S(n_60542), .A(n_6079), .B(regs_14[26]), .Z(pc_out
		[26]));
	notech_mux2 i_2812305(.S(n_60542), .A(n_6080), .B(regs_14[27]), .Z(pc_out
		[27]));
	notech_mux2 i_2912306(.S(n_60542), .A(n_6081), .B(regs_14[28]), .Z(pc_out
		[28]));
	notech_mux2 i_3012307(.S(n_60542), .A(n_6082), .B(regs_14[29]), .Z(pc_out
		[29]));
	notech_mux2 i_3112308(.S(n_60542), .A(n_6083), .B(regs_14[30]), .Z(pc_out
		[30]));
	notech_nand2 i_217879(.A(n_34491129), .B(n_34391128), .Z(write_data_25[1
		]));
	notech_nand2 i_317880(.A(n_34691131), .B(n_34591130), .Z(write_data_25[2
		]));
	notech_nand2 i_417881(.A(n_34891133), .B(n_34791132), .Z(write_data_25[3
		]));
	notech_nand2 i_517882(.A(n_35091135), .B(n_34991134), .Z(write_data_25[4
		]));
	notech_nand2 i_617883(.A(n_35291137), .B(n_35191136), .Z(write_data_25[5
		]));
	notech_nand2 i_717884(.A(n_35491139), .B(n_35391138), .Z(write_data_25[6
		]));
	notech_nand2 i_817885(.A(n_35691141), .B(n_35591140), .Z(write_data_25[7
		]));
	notech_nand2 i_917886(.A(n_35891143), .B(n_35791142), .Z(write_data_25[8
		]));
	notech_nand2 i_1017887(.A(n_36091145), .B(n_35991144), .Z(write_data_25[
		9]));
	notech_nand2 i_1617893(.A(n_36291147), .B(n_36191146), .Z(write_data_25[
		15]));
	notech_nand2 i_1717894(.A(n_36491149), .B(n_36391148), .Z(write_data_25[
		16]));
	notech_nand2 i_1817895(.A(n_36691151), .B(n_36591150), .Z(write_data_25[
		17]));
	notech_nand2 i_1917896(.A(n_36891153), .B(n_36791152), .Z(write_data_25[
		18]));
	notech_nand2 i_2017897(.A(n_37091155), .B(n_36991154), .Z(write_data_25[
		19]));
	notech_nand2 i_2117898(.A(n_37291157), .B(n_37191156), .Z(write_data_25[
		20]));
	notech_nand2 i_2217899(.A(n_37491159), .B(n_37391158), .Z(write_data_25[
		21]));
	notech_nand2 i_2317900(.A(n_37691161), .B(n_37591160), .Z(write_data_25[
		22]));
	notech_nand2 i_2417901(.A(n_37891163), .B(n_37791162), .Z(write_data_25[
		23]));
	notech_nand2 i_2517902(.A(n_38091165), .B(n_37991164), .Z(write_data_25[
		24]));
	notech_nand2 i_2617903(.A(n_38291167), .B(n_38191166), .Z(write_data_25[
		25]));
	notech_nand2 i_2717904(.A(n_38491169), .B(n_38391168), .Z(write_data_25[
		26]));
	notech_nand2 i_2817905(.A(n_38691171), .B(n_38591170), .Z(write_data_25[
		27]));
	notech_nand2 i_2917906(.A(n_38891173), .B(n_38791172), .Z(write_data_25[
		28]));
	notech_xor2 i_11271051(.A(\eflags[7] ), .B(\eflags[11] ), .Z(\cond[12] )
		);
	notech_nand2 i_19571050(.A(n_30635), .B(n_60138), .Z(\nbus_11297[0] ));
	notech_or2 i_254471049(.A(\eflags[6] ), .B(\cond[12] ), .Z(\cond[14] )
		);
	notech_or2 i_233071048(.A(\eflags[6] ), .B(\eflags[0] ), .Z(\cond[6] )
		);
	notech_mux2 i_3211733(.S(n_60773), .A(cr2[31]), .B(icr2[31]), .Z(n_12629
		));
	notech_mux2 i_3111732(.S(n_60773), .A(cr2[30]), .B(icr2[30]), .Z(n_12623
		));
	notech_mux2 i_3011731(.S(n_60773), .A(cr2[29]), .B(icr2[29]), .Z(n_12617
		));
	notech_mux2 i_2911730(.S(n_60773), .A(cr2[28]), .B(icr2[28]), .Z(n_12611
		));
	notech_mux2 i_2811729(.S(n_60773), .A(cr2[27]), .B(icr2[27]), .Z(n_12605
		));
	notech_mux2 i_2711728(.S(n_60773), .A(cr2[26]), .B(icr2[26]), .Z(n_12599
		));
	notech_mux2 i_2611727(.S(n_60773), .A(cr2[25]), .B(icr2[25]), .Z(n_12593
		));
	notech_mux2 i_2511726(.S(n_60773), .A(cr2[24]), .B(icr2[24]), .Z(n_12587
		));
	notech_mux2 i_2411725(.S(n_60769), .A(cr2[23]), .B(icr2[23]), .Z(n_12581
		));
	notech_mux2 i_2311724(.S(n_60769), .A(cr2[22]), .B(icr2[22]), .Z(n_12575
		));
	notech_mux2 i_2211723(.S(n_60769), .A(cr2[21]), .B(icr2[21]), .Z(n_12569
		));
	notech_mux2 i_2111722(.S(n_60773), .A(cr2[20]), .B(icr2[20]), .Z(n_12563
		));
	notech_mux2 i_2011721(.S(n_60773), .A(cr2[19]), .B(icr2[19]), .Z(n_12557
		));
	notech_mux2 i_1911720(.S(n_60773), .A(cr2[18]), .B(icr2[18]), .Z(n_12551
		));
	notech_mux2 i_1811719(.S(n_60773), .A(cr2[17]), .B(icr2[17]), .Z(n_12545
		));
	notech_mux2 i_1711718(.S(n_60773), .A(cr2[16]), .B(icr2[16]), .Z(n_12539
		));
	notech_mux2 i_1611717(.S(n_60774), .A(cr2[15]), .B(icr2[15]), .Z(n_12533
		));
	notech_mux2 i_1511716(.S(n_60774), .A(cr2[14]), .B(icr2[14]), .Z(n_12527
		));
	notech_mux2 i_1411715(.S(n_60774), .A(cr2[13]), .B(icr2[13]), .Z(n_12521
		));
	notech_mux2 i_1311714(.S(n_60774), .A(cr2[12]), .B(icr2[12]), .Z(n_12515
		));
	notech_mux2 i_1211713(.S(n_60774), .A(cr2[11]), .B(icr2[11]), .Z(n_12509
		));
	notech_mux2 i_1111712(.S(n_60774), .A(cr2[10]), .B(icr2[10]), .Z(n_12503
		));
	notech_mux2 i_1011711(.S(n_60774), .A(cr2[9]), .B(icr2[9]), .Z(n_12497)
		);
	notech_mux2 i_911710(.S(n_60774), .A(cr2[8]), .B(icr2[8]), .Z(n_12491)
		);
	notech_mux2 i_811709(.S(n_60774), .A(cr2[7]), .B(icr2[7]), .Z(n_12485)
		);
	notech_mux2 i_711708(.S(n_60774), .A(cr2[6]), .B(icr2[6]), .Z(n_12479)
		);
	notech_mux2 i_611707(.S(n_60773), .A(cr2[5]), .B(icr2[5]), .Z(n_12473)
		);
	notech_mux2 i_511706(.S(n_60774), .A(cr2[4]), .B(icr2[4]), .Z(n_12467)
		);
	notech_mux2 i_411705(.S(n_60774), .A(cr2[3]), .B(icr2[3]), .Z(n_12461)
		);
	notech_mux2 i_311704(.S(n_60774), .A(cr2[2]), .B(icr2[2]), .Z(n_12455)
		);
	notech_mux2 i_211703(.S(n_60774), .A(cr2[1]), .B(icr2[1]), .Z(n_12449)
		);
	notech_mux2 i_111702(.S(n_60765), .A(cr2[0]), .B(icr2[0]), .Z(n_12443)
		);
	notech_mux2 i_3211765(.S(n_56006), .A(n_5490), .B(n_5489), .Z(n_23298)
		);
	notech_mux2 i_3111764(.S(n_56005), .A(n_5488), .B(n_5487), .Z(n_23291)
		);
	notech_mux2 i_3011763(.S(n_56006), .A(n_5486), .B(n_5485), .Z(n_23284)
		);
	notech_mux2 i_2911762(.S(n_56006), .A(n_5484), .B(n_5483), .Z(n_23277)
		);
	notech_mux2 i_2811761(.S(n_56006), .A(n_5482), .B(n_5481), .Z(n_23270)
		);
	notech_mux2 i_2711760(.S(n_56005), .A(n_5480), .B(n_5479), .Z(n_23263)
		);
	notech_mux2 i_2611759(.S(n_56005), .A(n_5478), .B(n_5477), .Z(n_23256)
		);
	notech_mux2 i_2511758(.S(n_56005), .A(n_5476), .B(n_5475), .Z(n_23249)
		);
	notech_mux2 i_2411757(.S(n_56005), .A(n_5474), .B(n_5473), .Z(n_23242)
		);
	notech_mux2 i_2311756(.S(n_56005), .A(n_5472), .B(n_5471), .Z(n_23235)
		);
	notech_mux2 i_2211755(.S(n_56006), .A(n_5470), .B(n_5469), .Z(n_23228)
		);
	notech_mux2 i_2111754(.S(n_56006), .A(n_5468), .B(n_5467), .Z(n_23221)
		);
	notech_mux2 i_2011753(.S(n_56006), .A(n_5466), .B(n_5465), .Z(n_23214)
		);
	notech_mux2 i_1911752(.S(n_56006), .A(n_5464), .B(n_5463), .Z(n_23207)
		);
	notech_mux2 i_1811751(.S(n_56006), .A(n_5462), .B(n_5461), .Z(n_23200)
		);
	notech_mux2 i_1711750(.S(n_56006), .A(n_5460), .B(n_5459), .Z(n_23193)
		);
	notech_mux2 i_1611749(.S(n_56006), .A(n_5458), .B(n_5457), .Z(n_23186)
		);
	notech_mux2 i_1511748(.S(n_56006), .A(n_5456), .B(n_5455), .Z(n_23179)
		);
	notech_mux2 i_1411747(.S(n_56006), .A(n_5454), .B(n_5453), .Z(n_23172)
		);
	notech_mux2 i_1311746(.S(n_56006), .A(n_5452), .B(n_5451), .Z(n_23165)
		);
	notech_mux2 i_1211745(.S(n_56005), .A(n_5450), .B(n_5449), .Z(n_23158)
		);
	notech_mux2 i_1111744(.S(n_56006), .A(n_5448), .B(n_5447), .Z(n_23151)
		);
	notech_mux2 i_1011743(.S(n_56006), .A(n_5446), .B(n_5445), .Z(n_23144)
		);
	notech_mux2 i_911742(.S(n_56006), .A(n_5444), .B(n_5443), .Z(n_23137));
	notech_mux2 i_811741(.S(n_56006), .A(n_5442), .B(n_5441), .Z(n_23130));
	notech_mux2 i_711740(.S(n_56006), .A(n_5440), .B(n_5439), .Z(n_23123));
	notech_mux2 i_611739(.S(n_56006), .A(n_5438), .B(n_5437), .Z(n_23116));
	notech_mux2 i_511738(.S(n_56005), .A(n_5436), .B(n_5435), .Z(n_23109));
	notech_mux2 i_411737(.S(n_56005), .A(n_5434), .B(n_5433), .Z(n_23102));
	notech_mux2 i_311736(.S(n_56005), .A(n_5432), .B(n_5431), .Z(n_23095));
	notech_mux2 i_211735(.S(n_56005), .A(n_5430), .B(n_5429), .Z(n_23088));
	notech_mux2 i_111734(.S(n_56005), .A(n_5428), .B(n_5427), .Z(n_23081));
	notech_nand3 i_50442(.A(vliw_pc[3]), .B(n_273391892), .C(vliw_pc[1]), .Z
		(n_273591890));
	notech_nand2 i_26920(.A(n_60212), .B(n_27852), .Z(n_45891243));
	notech_ao3 i_17464(.A(n_60378), .B(opb[2]), .C(n_61151), .Z(n_45991244)
		);
	notech_ao3 i_17467(.A(n_60378), .B(opb[5]), .C(n_61151), .Z(n_46091245)
		);
	notech_and2 i_26922(.A(n_38991174), .B(n_60212), .Z(n_46191246));
	notech_and2 i_26923(.A(n_39091175), .B(n_60212), .Z(n_46291247));
	notech_ao3 i_2004(.A(n_27724), .B(n_27722), .C(vliw_pc[4]), .Z(n_273391892
		));
	notech_and2 i_19(.A(n_273191894), .B(n_272791898), .Z(n_273291893));
	notech_reg_set fsmf_reg_0(.CP(n_62432), .D(fsm[0]), .SD(n_61560), .Q(fsmf
		[0]));
	notech_reg_set fsmf_reg_1(.CP(n_62432), .D(fsm[1]), .SD(n_61560), .Q(fsmf
		[1]));
	notech_reg_set fsmf_reg_2(.CP(n_62432), .D(n_61175), .SD(n_61559), .Q(fsmf
		[2]));
	notech_reg_set fsmf_reg_3(.CP(n_62432), .D(fsm[3]), .SD(n_61559), .Q(fsmf
		[3]));
	notech_reg fsmf_reg_4(.CP(n_62432), .D(n_61160), .CD(n_61559), .Q(fsmf[4
		]));
	notech_reg calc_sz_reg_0(.CP(n_62432), .D(n_16561), .CD(n_61555), .Q(calc_sz
		[0]));
	notech_mux2 i_629(.S(n_27114), .A(calc_sz[0]), .B(instrc[108]), .Z(n_16561
		));
	notech_nao3 i_1880214(.A(n_273091895), .B(vliw_pc[2]), .C(n_272891897), 
		.Z(n_273191894));
	notech_reg calc_sz_reg_1(.CP(n_62432), .D(n_16567), .CD(n_61559), .Q(calc_sz
		[1]));
	notech_mux2 i_662(.S(n_27114), .A(n_58101), .B(instrc[109]), .Z(n_16567)
		);
	notech_and2 i_2072(.A(vliw_pc[3]), .B(n_27723), .Z(n_273091895));
	notech_reg calc_sz_reg_2(.CP(n_62432), .D(n_16573), .CD(n_61559), .Q(calc_sz
		[2]));
	notech_mux2 i_1568(.S(n_27114), .A(calc_sz[2]), .B(instrc[110]), .Z(n_16573
		));
	notech_reg calc_sz_reg_3(.CP(n_62432), .D(n_16579), .CD(n_61559), .Q(calc_sz
		[3]));
	notech_mux2 i_198495651(.S(n_27114), .A(calc_sz[3]), .B(instrc[111]), .Z
		(n_16579));
	notech_or2 i_132(.A(vliw_pc[4]), .B(vliw_pc[0]), .Z(n_272891897));
	notech_reg tsc_reg_0(.CP(n_62432), .D(n_4970), .CD(n_61559), .Q(tsc[0])
		);
	notech_reg tsc_reg_1(.CP(n_62432), .D(n_4972), .CD(n_61559), .Q(tsc[1])
		);
	notech_reg tsc_reg_2(.CP(n_62432), .D(n_4974), .CD(n_61559), .Q(tsc[2])
		);
	notech_reg tsc_reg_3(.CP(n_62534), .D(n_4976), .CD(n_61561), .Q(tsc[3])
		);
	notech_reg tsc_reg_4(.CP(n_62534), .D(n_4978), .CD(n_61561), .Q(tsc[4])
		);
	notech_reg tsc_reg_5(.CP(n_62534), .D(n_4980), .CD(n_61561), .Q(tsc[5])
		);
	notech_reg tsc_reg_6(.CP(n_62534), .D(n_4982), .CD(n_61561), .Q(tsc[6])
		);
	notech_reg tsc_reg_7(.CP(n_62534), .D(n_4984), .CD(n_61561), .Q(tsc[7])
		);
	notech_reg tsc_reg_8(.CP(n_62534), .D(n_4986), .CD(n_61562), .Q(tsc[8])
		);
	notech_reg tsc_reg_9(.CP(n_62534), .D(n_4988), .CD(n_61562), .Q(tsc[9])
		);
	notech_reg tsc_reg_10(.CP(n_62534), .D(n_4990), .CD(n_61561), .Q(tsc[10]
		));
	notech_reg tsc_reg_11(.CP(n_62534), .D(n_4992), .CD(n_61562), .Q(tsc[11]
		));
	notech_reg tsc_reg_12(.CP(n_62534), .D(n_4994), .CD(n_61561), .Q(tsc[12]
		));
	notech_reg tsc_reg_13(.CP(n_62534), .D(n_4996), .CD(n_61560), .Q(tsc[13]
		));
	notech_reg tsc_reg_14(.CP(n_62534), .D(n_4998), .CD(n_61561), .Q(tsc[14]
		));
	notech_reg tsc_reg_15(.CP(n_62534), .D(n_5000), .CD(n_61560), .Q(tsc[15]
		));
	notech_reg tsc_reg_16(.CP(n_62534), .D(n_5002), .CD(n_61560), .Q(tsc[16]
		));
	notech_reg tsc_reg_17(.CP(n_62534), .D(n_5004), .CD(n_61561), .Q(tsc[17]
		));
	notech_reg tsc_reg_18(.CP(n_62534), .D(n_5006), .CD(n_61561), .Q(tsc[18]
		));
	notech_reg tsc_reg_19(.CP(n_62534), .D(n_5008), .CD(n_61561), .Q(tsc[19]
		));
	notech_reg tsc_reg_20(.CP(n_62534), .D(n_5010), .CD(n_61561), .Q(tsc[20]
		));
	notech_reg tsc_reg_21(.CP(n_62534), .D(n_5012), .CD(n_61561), .Q(tsc[21]
		));
	notech_reg tsc_reg_22(.CP(n_62532), .D(n_5014), .CD(n_61553), .Q(tsc[22]
		));
	notech_reg tsc_reg_23(.CP(n_62532), .D(n_5016), .CD(n_61554), .Q(tsc[23]
		));
	notech_reg tsc_reg_24(.CP(n_62594), .D(n_5018), .CD(n_61553), .Q(tsc[24]
		));
	notech_reg tsc_reg_25(.CP(n_62594), .D(n_5020), .CD(n_61553), .Q(tsc[25]
		));
	notech_reg tsc_reg_26(.CP(n_62594), .D(n_5022), .CD(n_61554), .Q(tsc[26]
		));
	notech_reg tsc_reg_27(.CP(n_62594), .D(n_5024), .CD(n_61554), .Q(tsc[27]
		));
	notech_reg tsc_reg_28(.CP(n_62594), .D(n_5026), .CD(n_61554), .Q(tsc[28]
		));
	notech_reg tsc_reg_29(.CP(n_62594), .D(n_5028), .CD(n_61554), .Q(tsc[29]
		));
	notech_reg tsc_reg_30(.CP(n_62594), .D(n_5030), .CD(n_61554), .Q(tsc[30]
		));
	notech_reg tsc_reg_31(.CP(n_62594), .D(n_5032), .CD(n_61553), .Q(tsc[31]
		));
	notech_reg tsc_reg_32(.CP(n_62594), .D(n_5034), .CD(n_61553), .Q(tsc[32]
		));
	notech_reg tsc_reg_33(.CP(n_62594), .D(n_5036), .CD(n_61553), .Q(tsc[33]
		));
	notech_reg tsc_reg_34(.CP(n_62594), .D(n_5038), .CD(n_61553), .Q(tsc[34]
		));
	notech_reg tsc_reg_35(.CP(n_62594), .D(n_5040), .CD(n_61553), .Q(tsc[35]
		));
	notech_reg tsc_reg_36(.CP(n_62594), .D(n_5042), .CD(n_61553), .Q(tsc[36]
		));
	notech_reg tsc_reg_37(.CP(n_62594), .D(n_5044), .CD(n_61553), .Q(tsc[37]
		));
	notech_reg tsc_reg_38(.CP(n_62594), .D(n_5046), .CD(n_61553), .Q(tsc[38]
		));
	notech_reg tsc_reg_39(.CP(n_62594), .D(n_5048), .CD(n_61553), .Q(tsc[39]
		));
	notech_reg tsc_reg_40(.CP(n_62594), .D(n_5050), .CD(n_61553), .Q(tsc[40]
		));
	notech_reg tsc_reg_41(.CP(n_62594), .D(n_5052), .CD(n_61555), .Q(tsc[41]
		));
	notech_reg tsc_reg_42(.CP(n_62532), .D(n_5054), .CD(n_61555), .Q(tsc[42]
		));
	notech_reg tsc_reg_43(.CP(n_62532), .D(n_5056), .CD(n_61555), .Q(tsc[43]
		));
	notech_reg tsc_reg_44(.CP(n_62532), .D(n_5058), .CD(n_61555), .Q(tsc[44]
		));
	notech_reg tsc_reg_45(.CP(n_62532), .D(n_5060), .CD(n_61555), .Q(tsc[45]
		));
	notech_reg tsc_reg_46(.CP(n_62532), .D(n_5062), .CD(n_61555), .Q(tsc[46]
		));
	notech_reg tsc_reg_47(.CP(n_62532), .D(n_5064), .CD(n_61555), .Q(tsc[47]
		));
	notech_reg tsc_reg_48(.CP(n_62532), .D(n_5066), .CD(n_61555), .Q(tsc[48]
		));
	notech_reg tsc_reg_49(.CP(n_62532), .D(n_5068), .CD(n_61555), .Q(tsc[49]
		));
	notech_reg tsc_reg_50(.CP(n_62532), .D(n_5070), .CD(n_61555), .Q(tsc[50]
		));
	notech_reg tsc_reg_51(.CP(n_62532), .D(n_5072), .CD(n_61554), .Q(tsc[51]
		));
	notech_reg tsc_reg_52(.CP(n_62594), .D(n_5074), .CD(n_61554), .Q(tsc[52]
		));
	notech_reg tsc_reg_53(.CP(n_62530), .D(n_5076), .CD(n_61554), .Q(tsc[53]
		));
	notech_reg tsc_reg_54(.CP(n_62530), .D(n_5078), .CD(n_61554), .Q(tsc[54]
		));
	notech_reg tsc_reg_55(.CP(n_62590), .D(n_5080), .CD(n_61554), .Q(tsc[55]
		));
	notech_reg tsc_reg_56(.CP(n_62590), .D(n_5082), .CD(n_61555), .Q(tsc[56]
		));
	notech_reg tsc_reg_57(.CP(n_62590), .D(n_5084), .CD(n_61555), .Q(tsc[57]
		));
	notech_reg tsc_reg_58(.CP(n_62590), .D(n_5086), .CD(n_61554), .Q(tsc[58]
		));
	notech_reg tsc_reg_59(.CP(n_62590), .D(n_5088), .CD(n_61554), .Q(tsc[59]
		));
	notech_reg tsc_reg_60(.CP(n_62590), .D(n_5090), .CD(n_61567), .Q(tsc[60]
		));
	notech_reg tsc_reg_61(.CP(n_62590), .D(n_5092), .CD(n_61567), .Q(tsc[61]
		));
	notech_reg tsc_reg_62(.CP(n_62590), .D(n_5094), .CD(n_61566), .Q(tsc[62]
		));
	notech_reg tsc_reg_63(.CP(n_62590), .D(n_5096), .CD(n_61567), .Q(tsc[63]
		));
	notech_reg_set first_rep_reg(.CP(n_62590), .D(n_16715), .SD(n_61567), .Q
		(first_rep));
	notech_mux2 i_2465(.S(n_19928), .A(first_rep), .B(n_26983), .Z(n_16715)
		);
	notech_nao3 i_50440(.A(vliw_pc[3]), .B(n_32843), .C(n_272591900), .Z(n_272791898
		));
	notech_reg_set fecx_reg(.CP(n_62674), .D(n_16722), .SD(1'b1), .Q(fecx)
		);
	notech_mux2 i_2473(.S(n_27115), .A(fecx), .B(n_322487498), .Z(n_16722)
		);
	notech_reg sav_ecx_reg_0(.CP(n_62674), .D(n_16729), .CD(n_61567), .Q(sav_ecx
		[0]));
	notech_mux2 i_2481(.S(n_59763), .A(ecx[0]), .B(sav_ecx[0]), .Z(n_16729)
		);
	notech_or2 i_1943(.A(vliw_pc[4]), .B(vliw_pc[2]), .Z(n_272591900));
	notech_reg sav_ecx_reg_1(.CP(n_62674), .D(n_16737), .CD(n_61567), .Q(sav_ecx
		[1]));
	notech_mux2 i_2489(.S(n_59763), .A(ecx[1]), .B(sav_ecx[1]), .Z(n_16737)
		);
	notech_ao3 i_1661(.A(n_27720), .B(n_27717), .C(fsm[0]), .Z(n_272491901)
		);
	notech_reg sav_ecx_reg_2(.CP(n_62674), .D(n_16744), .CD(n_61567), .Q(sav_ecx
		[2]));
	notech_mux2 i_2497(.S(n_59763), .A(ecx[2]), .B(sav_ecx[2]), .Z(n_16744)
		);
	notech_reg sav_ecx_reg_3(.CP(n_62674), .D(n_16751), .CD(n_61567), .Q(sav_ecx
		[3]));
	notech_mux2 i_2505(.S(n_59763), .A(ecx[3]), .B(sav_ecx[3]), .Z(n_16751)
		);
	notech_and4 i_617755(.A(n_2961), .B(n_298691832), .C(n_272191904), .D(n_2692
		), .Z(n_272291903));
	notech_reg sav_ecx_reg_4(.CP(n_62674), .D(n_16758), .CD(n_61566), .Q(sav_ecx
		[4]));
	notech_mux2 i_2513(.S(n_59763), .A(ecx[4]), .B(sav_ecx[4]), .Z(n_16758)
		);
	notech_nand2 i_977(.A(resa_shiftbox[5]), .B(n_26712), .Z(n_272191904));
	notech_reg sav_ecx_reg_5(.CP(n_62674), .D(n_16765), .CD(n_61566), .Q(sav_ecx
		[5]));
	notech_mux2 i_2521(.S(n_59764), .A(ecx[5]), .B(sav_ecx[5]), .Z(n_16765)
		);
	notech_or2 i_976(.A(n_57498), .B(n_29651), .Z(n_272091905));
	notech_reg sav_ecx_reg_6(.CP(n_62674), .D(n_16773), .CD(n_61566), .Q(sav_ecx
		[6]));
	notech_mux2 i_2529(.S(n_59764), .A(ecx[6]), .B(sav_ecx[6]), .Z(n_16773)
		);
	notech_reg sav_ecx_reg_7(.CP(n_62674), .D(n_16780), .CD(n_61566), .Q(sav_ecx
		[7]));
	notech_mux2 i_2537(.S(n_59764), .A(ecx[7]), .B(sav_ecx[7]), .Z(n_16780)
		);
	notech_reg sav_ecx_reg_8(.CP(n_62674), .D(n_16787), .CD(n_61566), .Q(sav_ecx
		[8]));
	notech_mux2 i_2545(.S(n_59763), .A(ecx[8]), .B(sav_ecx[8]), .Z(n_16787)
		);
	notech_nao3 i_985(.A(\nbus_14520[5] ), .B(n_2950), .C(n_57933), .Z(n_271791908
		));
	notech_reg sav_ecx_reg_9(.CP(n_62674), .D(n_16794), .CD(n_61566), .Q(sav_ecx
		[9]));
	notech_mux2 i_2553(.S(n_59763), .A(ecx[9]), .B(sav_ecx[9]), .Z(n_16794)
		);
	notech_reg sav_ecx_reg_10(.CP(n_62674), .D(n_16801), .CD(n_61566), .Q(sav_ecx
		[10]));
	notech_mux2 i_2562(.S(n_59764), .A(ecx[10]), .B(sav_ecx[10]), .Z(n_16801
		));
	notech_reg sav_ecx_reg_11(.CP(n_62674), .D(n_16809), .CD(n_61566), .Q(sav_ecx
		[11]));
	notech_mux2 i_2570(.S(n_59758), .A(ecx[11]), .B(sav_ecx[11]), .Z(n_16809
		));
	notech_nand2 i_975(.A(readio_data[5]), .B(n_26711), .Z(n_271491911));
	notech_reg sav_ecx_reg_12(.CP(n_62674), .D(n_16816), .CD(n_61566), .Q(sav_ecx
		[12]));
	notech_mux2 i_2579(.S(n_59758), .A(ecx[12]), .B(sav_ecx[12]), .Z(n_16816
		));
	notech_nand3 i_961(.A(n_1891), .B(mul64[5]), .C(n_60312), .Z(n_271391912
		));
	notech_reg sav_ecx_reg_13(.CP(n_62674), .D(n_16823), .CD(n_61566), .Q(sav_ecx
		[13]));
	notech_mux2 i_2587(.S(n_59758), .A(ecx[13]), .B(sav_ecx[13]), .Z(n_16823
		));
	notech_nao3 i_962(.A(resa_arithbox[5]), .B(n_60316), .C(n_58072), .Z(n_271291913
		));
	notech_reg sav_ecx_reg_14(.CP(n_62674), .D(n_16830), .CD(n_61570), .Q(sav_ecx
		[14]));
	notech_mux2 i_2595(.S(n_59758), .A(ecx[14]), .B(sav_ecx[14]), .Z(n_16830
		));
	notech_nao3 i_965(.A(n_32316), .B(nbus_14521[5]), .C(n_57933), .Z(n_271191914
		));
	notech_reg sav_ecx_reg_15(.CP(n_62674), .D(n_16837), .CD(n_61570), .Q(sav_ecx
		[15]));
	notech_mux2 i_2604(.S(n_59758), .A(ecx[15]), .B(sav_ecx[15]), .Z(n_16837
		));
	notech_or2 i_974(.A(n_22313), .B(n_59205), .Z(n_271091915));
	notech_reg sav_ecx_reg_16(.CP(n_62674), .D(n_16845), .CD(n_61570), .Q(sav_ecx
		[16]));
	notech_mux2 i_2612(.S(n_59758), .A(ecx[16]), .B(sav_ecx[16]), .Z(n_16845
		));
	notech_reg sav_ecx_reg_17(.CP(n_62590), .D(n_16852), .CD(n_61570), .Q(sav_ecx
		[17]));
	notech_mux2 i_2620(.S(n_59763), .A(ecx[17]), .B(sav_ecx[17]), .Z(n_16852
		));
	notech_reg sav_ecx_reg_18(.CP(n_62674), .D(n_16859), .CD(n_61570), .Q(sav_ecx
		[18]));
	notech_mux2 i_2628(.S(n_59763), .A(ecx[18]), .B(sav_ecx[18]), .Z(n_16859
		));
	notech_or2 i_980(.A(n_57165), .B(n_57653), .Z(n_2707));
	notech_reg sav_ecx_reg_19(.CP(n_62592), .D(n_16866), .CD(n_61570), .Q(sav_ecx
		[19]));
	notech_mux2 i_2636(.S(n_59763), .A(ecx[19]), .B(sav_ecx[19]), .Z(n_16866
		));
	notech_reg sav_ecx_reg_20(.CP(n_62592), .D(n_16873), .CD(n_61571), .Q(sav_ecx
		[20]));
	notech_mux2 i_2644(.S(n_59763), .A(ecx[20]), .B(sav_ecx[20]), .Z(n_16873
		));
	notech_reg sav_ecx_reg_21(.CP(n_62592), .D(n_16881), .CD(n_61570), .Q(sav_ecx
		[21]));
	notech_mux2 i_2652(.S(n_59763), .A(ecx[21]), .B(sav_ecx[21]), .Z(n_16881
		));
	notech_nand3 i_986(.A(n_25374), .B(\nbus_14522[5] ), .C(n_2952), .Z(n_270491919
		));
	notech_reg sav_ecx_reg_22(.CP(n_62592), .D(n_16888), .CD(n_61570), .Q(sav_ecx
		[22]));
	notech_mux2 i_2660(.S(n_59763), .A(ecx[22]), .B(sav_ecx[22]), .Z(n_16888
		));
	notech_reg sav_ecx_reg_23(.CP(n_62592), .D(n_16895), .CD(n_61570), .Q(sav_ecx
		[23]));
	notech_mux2 i_2668(.S(n_59766), .A(ecx[23]), .B(sav_ecx[23]), .Z(n_16895
		));
	notech_reg sav_ecx_reg_24(.CP(n_62592), .D(n_16901), .CD(n_61567), .Q(sav_ecx
		[24]));
	notech_mux2 i_2676(.S(n_59766), .A(ecx[24]), .B(sav_ecx[24]), .Z(n_16901
		));
	notech_reg sav_ecx_reg_25(.CP(n_62592), .D(n_16907), .CD(n_61567), .Q(sav_ecx
		[25]));
	notech_mux2 i_2684(.S(n_59766), .A(ecx[25]), .B(sav_ecx[25]), .Z(n_16907
		));
	notech_reg sav_ecx_reg_26(.CP(n_62592), .D(n_16913), .CD(n_61567), .Q(sav_ecx
		[26]));
	notech_mux2 i_2692(.S(n_59766), .A(ecx[26]), .B(sav_ecx[26]), .Z(n_16913
		));
	notech_reg sav_ecx_reg_27(.CP(n_62592), .D(n_16919), .CD(n_61567), .Q(sav_ecx
		[27]));
	notech_mux2 i_2700(.S(n_59766), .A(ecx[27]), .B(sav_ecx[27]), .Z(n_16919
		));
	notech_reg sav_ecx_reg_28(.CP(n_62592), .D(n_16925), .CD(n_61567), .Q(sav_ecx
		[28]));
	notech_mux2 i_2708(.S(n_59766), .A(ecx[28]), .B(sav_ecx[28]), .Z(n_16925
		));
	notech_or4 i_979(.A(n_59418), .B(n_315291671), .C(n_60207), .D(n_27905),
		 .Z(n_2697));
	notech_reg sav_ecx_reg_29(.CP(n_62592), .D(n_16931), .CD(n_61570), .Q(sav_ecx
		[29]));
	notech_mux2 i_2716(.S(n_59766), .A(ecx[29]), .B(sav_ecx[29]), .Z(n_16931
		));
	notech_nao3 i_982(.A(resa_shift4box[5]), .B(n_57899), .C(n_293591841), .Z
		(n_2696));
	notech_reg sav_ecx_reg_30(.CP(n_62592), .D(n_16937), .CD(n_61570), .Q(sav_ecx
		[30]));
	notech_mux2 i_2724(.S(n_59766), .A(ecx[30]), .B(sav_ecx[30]), .Z(n_16937
		));
	notech_reg sav_ecx_reg_31(.CP(n_62592), .D(n_16943), .CD(n_61570), .Q(sav_ecx
		[31]));
	notech_mux2 i_2732(.S(n_59766), .A(ecx[31]), .B(sav_ecx[31]), .Z(n_16943
		));
	notech_reg fesp_reg(.CP(n_62592), .D(n_16949), .CD(n_61570), .Q(fesp));
	notech_mux2 i_2740(.S(n_27152), .A(fesp), .B(n_322387497), .Z(n_16949)
		);
	notech_ao4 i_957(.A(n_57143), .B(nbus_11310[5]), .C(n_2653), .D(n_60207)
		, .Z(n_2693));
	notech_reg_set sav_esp_reg_0(.CP(n_62592), .D(n_16955), .SD(1'b1), .Q(sav_esp
		[0]));
	notech_mux2 i_2748(.S(n_328390781), .A(regs_4[0]), .B(sav_esp[0]), .Z(n_16955
		));
	notech_or2 i_991(.A(n_2693), .B(n_57583), .Z(n_2692));
	notech_reg_set sav_esp_reg_1(.CP(n_62592), .D(n_16961), .SD(1'b1), .Q(sav_esp
		[1]));
	notech_mux2 i_2756(.S(n_328390781), .A(regs_4[1]), .B(sav_esp[1]), .Z(n_16961
		));
	notech_xor2 i_954(.A(n_27885), .B(opa[5]), .Z(n_2691));
	notech_reg_set sav_esp_reg_2(.CP(n_62592), .D(n_16967), .SD(1'b1), .Q(sav_esp
		[2]));
	notech_mux2 i_2764(.S(n_328390781), .A(regs_4[2]), .B(sav_esp[2]), .Z(n_16967
		));
	notech_reg_set sav_esp_reg_3(.CP(n_62592), .D(n_16973), .SD(1'b1), .Q(sav_esp
		[3]));
	notech_mux2 i_2772(.S(n_328390781), .A(regs_4[3]), .B(sav_esp[3]), .Z(n_16973
		));
	notech_reg_set sav_esp_reg_4(.CP(n_62592), .D(n_16979), .SD(1'b1), .Q(sav_esp
		[4]));
	notech_mux2 i_2780(.S(n_328390781), .A(regs_4[4]), .B(sav_esp[4]), .Z(n_16979
		));
	notech_reg_set sav_esp_reg_5(.CP(n_62530), .D(n_16985), .SD(1'b1), .Q(sav_esp
		[5]));
	notech_mux2 i_2788(.S(n_328390781), .A(regs_4[5]), .B(sav_esp[5]), .Z(n_16985
		));
	notech_reg_set sav_esp_reg_6(.CP(n_62530), .D(n_16991), .SD(1'b1), .Q(sav_esp
		[6]));
	notech_mux2 i_2796(.S(n_328390781), .A(regs_4[6]), .B(sav_esp[6]), .Z(n_16991
		));
	notech_reg_set sav_esp_reg_7(.CP(n_62530), .D(n_16997), .SD(1'b1), .Q(sav_esp
		[7]));
	notech_mux2 i_2804(.S(n_328390781), .A(regs_4[7]), .B(sav_esp[7]), .Z(n_16997
		));
	notech_or4 i_572(.A(n_60969), .B(n_60958), .C(n_27924), .D(n_62836), .Z(n_2685
		));
	notech_reg_set sav_esp_reg_8(.CP(n_62530), .D(n_17003), .SD(1'b1), .Q(sav_esp
		[8]));
	notech_mux2 i_2812(.S(n_328390781), .A(regs_4[8]), .B(sav_esp[8]), .Z(n_17003
		));
	notech_or4 i_3150(.A(n_60969), .B(n_60958), .C(n_25619), .D(n_62836), .Z
		(n_2684));
	notech_reg_set sav_esp_reg_9(.CP(n_62530), .D(n_17009), .SD(1'b1), .Q(sav_esp
		[9]));
	notech_mux2 i_2820(.S(n_328390781), .A(regs_4[9]), .B(sav_esp[9]), .Z(n_17009
		));
	notech_nand2 i_1456(.A(n_23006), .B(n_2682), .Z(n_2683));
	notech_reg_set sav_esp_reg_10(.CP(n_62530), .D(n_17015), .SD(1'b1), .Q(sav_esp
		[10]));
	notech_mux2 i_2829(.S(n_328390781), .A(regs_4[10]), .B(sav_esp[10]), .Z(n_17015
		));
	notech_or4 i_565(.A(n_27925), .B(n_60863), .C(n_62870), .D(n_60986), .Z(n_2682
		));
	notech_reg_set sav_esp_reg_11(.CP(n_62530), .D(n_17021), .SD(1'b1), .Q(sav_esp
		[11]));
	notech_mux2 i_2838(.S(n_328390781), .A(regs_4[11]), .B(sav_esp[11]), .Z(n_17021
		));
	notech_reg_set sav_esp_reg_12(.CP(n_62530), .D(n_17027), .SD(1'b1), .Q(sav_esp
		[12]));
	notech_mux2 i_2847(.S(n_328390781), .A(regs_4[12]), .B(sav_esp[12]), .Z(n_17027
		));
	notech_reg_set sav_esp_reg_13(.CP(n_62530), .D(n_17033), .SD(1'b1), .Q(sav_esp
		[13]));
	notech_mux2 i_2856(.S(n_328390781), .A(regs_4[13]), .B(sav_esp[13]), .Z(n_17033
		));
	notech_reg_set sav_esp_reg_14(.CP(n_62530), .D(n_17039), .SD(1'b1), .Q(sav_esp
		[14]));
	notech_mux2 i_2865(.S(n_328390781), .A(regs_4[14]), .B(sav_esp[14]), .Z(n_17039
		));
	notech_or4 i_3132(.A(n_32729), .B(n_58086), .C(n_62836), .D(n_60933), .Z
		(n_2678));
	notech_reg_set sav_esp_reg_15(.CP(n_62590), .D(n_17045), .SD(1'b1), .Q(sav_esp
		[15]));
	notech_mux2 i_2874(.S(n_328390781), .A(regs_4[15]), .B(sav_esp[15]), .Z(n_17045
		));
	notech_or4 i_3183(.A(n_32643), .B(n_58086), .C(n_60933), .D(n_60904), .Z
		(n_2677));
	notech_reg_set sav_esp_reg_16(.CP(n_62584), .D(n_17051), .SD(1'b1), .Q(sav_esp
		[16]));
	notech_mux2 i_2882(.S(n_54389), .A(regs_4[16]), .B(sav_esp[16]), .Z(n_17051
		));
	notech_or4 i_551(.A(n_27925), .B(n_1868), .C(n_60933), .D(n_60904), .Z(n_2676
		));
	notech_reg_set sav_esp_reg_17(.CP(n_62528), .D(n_17057), .SD(1'b1), .Q(sav_esp
		[17]));
	notech_mux2 i_2890(.S(n_54389), .A(regs_4[17]), .B(sav_esp[17]), .Z(n_17057
		));
	notech_reg_set sav_esp_reg_18(.CP(n_62584), .D(n_17063), .SD(1'b1), .Q(sav_esp
		[18]));
	notech_mux2 i_2898(.S(n_54389), .A(regs_4[18]), .B(sav_esp[18]), .Z(n_17063
		));
	notech_reg_set sav_esp_reg_19(.CP(n_62584), .D(n_17069), .SD(1'b1), .Q(sav_esp
		[19]));
	notech_mux2 i_2906(.S(n_54389), .A(regs_4[19]), .B(sav_esp[19]), .Z(n_17069
		));
	notech_reg_set sav_esp_reg_20(.CP(n_62584), .D(n_17076), .SD(1'b1), .Q(sav_esp
		[20]));
	notech_mux2 i_2914(.S(n_54389), .A(regs_4[20]), .B(sav_esp[20]), .Z(n_17076
		));
	notech_reg_set sav_esp_reg_21(.CP(n_62584), .D(n_17083), .SD(1'b1), .Q(sav_esp
		[21]));
	notech_mux2 i_2922(.S(n_54389), .A(regs_4[21]), .B(sav_esp[21]), .Z(n_17083
		));
	notech_reg_set sav_esp_reg_22(.CP(n_62584), .D(n_17090), .SD(1'b1), .Q(sav_esp
		[22]));
	notech_mux2 i_2930(.S(n_54389), .A(regs_4[22]), .B(sav_esp[22]), .Z(n_17090
		));
	notech_reg_set sav_esp_reg_23(.CP(n_62584), .D(n_17097), .SD(1'b1), .Q(sav_esp
		[23]));
	notech_mux2 i_2939(.S(n_54389), .A(regs_4[23]), .B(sav_esp[23]), .Z(n_17097
		));
	notech_reg_set sav_esp_reg_24(.CP(n_62584), .D(n_17104), .SD(1'b1), .Q(sav_esp
		[24]));
	notech_mux2 i_2947(.S(n_54389), .A(regs_4[24]), .B(sav_esp[24]), .Z(n_17104
		));
	notech_ao4 i_275(.A(n_2896), .B(n_26757), .C(n_26983), .D(n_1874), .Z(n_266891921
		));
	notech_reg_set sav_esp_reg_25(.CP(n_62584), .D(n_17113), .SD(1'b1), .Q(sav_esp
		[25]));
	notech_mux2 i_2955(.S(n_54389), .A(regs_4[25]), .B(sav_esp[25]), .Z(n_17113
		));
	notech_reg_set sav_esp_reg_26(.CP(n_62584), .D(n_17120), .SD(1'b1), .Q(sav_esp
		[26]));
	notech_mux2 i_2963(.S(n_54389), .A(regs_4[26]), .B(sav_esp[26]), .Z(n_17120
		));
	notech_nao3 i_497(.A(reps[0]), .B(n_2665), .C(first_rep), .Z(n_2666));
	notech_reg_set sav_esp_reg_27(.CP(n_62584), .D(n_17127), .SD(1'b1), .Q(sav_esp
		[27]));
	notech_mux2 i_2971(.S(n_54389), .A(regs_4[27]), .B(sav_esp[27]), .Z(n_17127
		));
	notech_xor2 i_103(.A(nZF), .B(reps[1]), .Z(n_2665));
	notech_reg_set sav_esp_reg_28(.CP(n_62670), .D(n_17136), .SD(1'b1), .Q(sav_esp
		[28]));
	notech_mux2 i_2979(.S(n_54389), .A(regs_4[28]), .B(sav_esp[28]), .Z(n_17136
		));
	notech_nand2 i_495(.A(reps[0]), .B(first_rep), .Z(n_2664));
	notech_reg_set sav_esp_reg_29(.CP(n_62670), .D(n_17144), .SD(1'b1), .Q(sav_esp
		[29]));
	notech_mux2 i_2988(.S(n_54389), .A(regs_4[29]), .B(sav_esp[29]), .Z(n_17144
		));
	notech_nao3 i_496(.A(n_2659), .B(n_2664), .C(n_291691848), .Z(n_2663));
	notech_reg_set sav_esp_reg_30(.CP(n_62670), .D(n_17151), .SD(1'b1), .Q(sav_esp
		[30]));
	notech_mux2 i_2997(.S(n_54389), .A(regs_4[30]), .B(sav_esp[30]), .Z(n_17151
		));
	notech_reg_set sav_esp_reg_31(.CP(n_62670), .D(n_17158), .SD(1'b1), .Q(sav_esp
		[31]));
	notech_mux2 i_3005(.S(n_54389), .A(regs_4[31]), .B(sav_esp[31]), .Z(n_17158
		));
	notech_reg sav_esi_reg_0(.CP(n_62670), .D(n_17166), .CD(n_61564), .Q(sav_esi
		[0]));
	notech_mux2 i_3013(.S(n_59766), .A(regs_6[0]), .B(sav_esi[0]), .Z(n_17166
		));
	notech_or4 i_30(.A(n_291991845), .B(n_2929), .C(n_2926), .D(n_2922), .Z(n_2660
		));
	notech_reg sav_esi_reg_1(.CP(n_62670), .D(n_17173), .CD(n_61564), .Q(sav_esi
		[1]));
	notech_mux2 i_3021(.S(n_59766), .A(regs_6[1]), .B(sav_esi[1]), .Z(n_17173
		));
	notech_nand2 i_492(.A(n_2660), .B(n_60542), .Z(n_2659));
	notech_reg sav_esi_reg_2(.CP(n_62670), .D(n_17180), .CD(n_61564), .Q(sav_esi
		[2]));
	notech_mux2 i_3029(.S(n_59766), .A(regs_6[2]), .B(sav_esi[2]), .Z(n_17180
		));
	notech_or4 i_461(.A(n_27501), .B(n_62870), .C(n_60986), .D(n_2657), .Z(n_2658
		));
	notech_reg sav_esi_reg_3(.CP(n_62670), .D(n_17187), .CD(n_61564), .Q(sav_esi
		[3]));
	notech_mux2 i_3038(.S(n_59764), .A(regs_6[3]), .B(sav_esi[3]), .Z(n_17187
		));
	notech_and2 i_460(.A(n_60888), .B(n_59418), .Z(n_2657));
	notech_reg sav_esi_reg_4(.CP(n_62670), .D(n_17194), .CD(n_61564), .Q(sav_esi
		[4]));
	notech_mux2 i_3046(.S(n_59764), .A(regs_6[4]), .B(sav_esi[4]), .Z(n_17194
		));
	notech_reg sav_esi_reg_5(.CP(n_62670), .D(n_17202), .CD(n_61564), .Q(sav_esi
		[5]));
	notech_mux2 i_3055(.S(n_59764), .A(regs_6[5]), .B(sav_esi[5]), .Z(n_17202
		));
	notech_reg sav_esi_reg_6(.CP(n_62670), .D(n_17209), .CD(n_61564), .Q(sav_esi
		[6]));
	notech_mux2 i_3063(.S(n_59764), .A(regs_6[6]), .B(sav_esi[6]), .Z(n_17209
		));
	notech_or4 i_3082(.A(n_27994), .B(n_2877), .C(n_62836), .D(n_60931), .Z(n_2654
		));
	notech_reg sav_esi_reg_7(.CP(n_62670), .D(n_17216), .CD(n_61564), .Q(sav_esi
		[7]));
	notech_mux2 i_3072(.S(n_59764), .A(regs_6[7]), .B(sav_esi[7]), .Z(n_17216
		));
	notech_and4 i_441(.A(n_1870), .B(n_289791858), .C(n_58046), .D(n_25386),
		 .Z(n_2653));
	notech_reg sav_esi_reg_8(.CP(n_62670), .D(n_17223), .CD(n_61564), .Q(sav_esi
		[8]));
	notech_mux2 i_3081(.S(n_59764), .A(regs_6[8]), .B(sav_esi[8]), .Z(n_17223
		));
	notech_reg sav_esi_reg_9(.CP(n_62670), .D(n_17230), .CD(n_61562), .Q(sav_esi
		[9]));
	notech_mux2 i_3090(.S(n_59764), .A(regs_6[9]), .B(sav_esi[9]), .Z(n_17230
		));
	notech_reg sav_esi_reg_10(.CP(n_62670), .D(n_17238), .CD(n_61562), .Q(sav_esi
		[10]));
	notech_mux2 i_3100(.S(n_59766), .A(regs_6[10]), .B(sav_esi[10]), .Z(n_17238
		));
	notech_reg sav_esi_reg_11(.CP(n_62670), .D(n_17245), .CD(n_61562), .Q(sav_esi
		[11]));
	notech_mux2 i_3109(.S(n_59766), .A(regs_6[11]), .B(sav_esi[11]), .Z(n_17245
		));
	notech_nand2 i_419(.A(n_62892), .B(n_59429), .Z(n_2649));
	notech_reg sav_esi_reg_12(.CP(n_62670), .D(n_17252), .CD(n_61562), .Q(sav_esi
		[12]));
	notech_mux2 i_3118(.S(n_59764), .A(regs_6[12]), .B(sav_esi[12]), .Z(n_17252
		));
	notech_reg sav_esi_reg_13(.CP(n_62670), .D(n_17259), .CD(n_61562), .Q(sav_esi
		[13]));
	notech_mux2 i_3127(.S(n_59764), .A(regs_6[13]), .B(sav_esi[13]), .Z(n_17259
		));
	notech_and2 i_984(.A(n_1899), .B(n_1900), .Z(n_2647));
	notech_reg sav_esi_reg_14(.CP(n_62670), .D(n_17266), .CD(n_61562), .Q(sav_esi
		[14]));
	notech_mux2 i_3136(.S(n_59764), .A(regs_6[14]), .B(sav_esi[14]), .Z(n_17266
		));
	notech_reg sav_esi_reg_15(.CP(n_62734), .D(n_17272), .CD(n_61562), .Q(sav_esi
		[15]));
	notech_mux2 i_3144(.S(n_59758), .A(regs_6[15]), .B(sav_esi[15]), .Z(n_17272
		));
	notech_nand3 i_356(.A(n_273391892), .B(instrc[70]), .C(n_273091895), .Z(n_2645
		));
	notech_reg sav_esi_reg_16(.CP(n_62668), .D(n_17278), .CD(n_61562), .Q(sav_esi
		[16]));
	notech_mux2 i_3153(.S(n_59751), .A(regs_6[16]), .B(sav_esi[16]), .Z(n_17278
		));
	notech_reg sav_esi_reg_17(.CP(n_62734), .D(n_17284), .CD(n_61562), .Q(sav_esi
		[17]));
	notech_mux2 i_3161(.S(n_59751), .A(regs_6[17]), .B(sav_esi[17]), .Z(n_17284
		));
	notech_reg sav_esi_reg_18(.CP(n_62734), .D(n_17290), .CD(n_61562), .Q(sav_esi
		[18]));
	notech_mux2 i_3169(.S(n_59751), .A(regs_6[18]), .B(sav_esi[18]), .Z(n_17290
		));
	notech_and4 i_348(.A(vliw_pc[2]), .B(instrc[62]), .C(n_32843), .D(n_2739
		), .Z(n_2642));
	notech_reg sav_esi_reg_19(.CP(n_62734), .D(n_17296), .CD(n_61565), .Q(sav_esi
		[19]));
	notech_mux2 i_3177(.S(n_59751), .A(regs_6[19]), .B(sav_esi[19]), .Z(n_17296
		));
	notech_nand3 i_354(.A(instrc[6]), .B(n_273391892), .C(n_274591882), .Z(n_264191922
		));
	notech_reg sav_esi_reg_20(.CP(n_62734), .D(n_17302), .CD(n_61565), .Q(sav_esi
		[20]));
	notech_mux2 i_3186(.S(n_59751), .A(regs_6[20]), .B(sav_esi[20]), .Z(n_17302
		));
	notech_reg sav_esi_reg_21(.CP(n_62734), .D(n_17308), .CD(n_61565), .Q(sav_esi
		[21]));
	notech_mux2 i_3194(.S(n_59751), .A(regs_6[21]), .B(sav_esi[21]), .Z(n_17308
		));
	notech_reg sav_esi_reg_22(.CP(n_62734), .D(n_17314), .CD(n_61565), .Q(sav_esi
		[22]));
	notech_mux2 i_3202(.S(n_59764), .A(regs_6[22]), .B(sav_esi[22]), .Z(n_17314
		));
	notech_reg sav_esi_reg_23(.CP(n_62734), .D(n_17320), .CD(n_61565), .Q(sav_esi
		[23]));
	notech_mux2 i_3210(.S(n_59764), .A(regs_6[23]), .B(sav_esi[23]), .Z(n_17320
		));
	notech_reg sav_esi_reg_24(.CP(n_62734), .D(n_17326), .CD(n_61566), .Q(sav_esi
		[24]));
	notech_mux2 i_3218(.S(n_59764), .A(regs_6[24]), .B(sav_esi[24]), .Z(n_17326
		));
	notech_reg sav_esi_reg_25(.CP(n_62734), .D(n_17332), .CD(n_61566), .Q(sav_esi
		[25]));
	notech_mux2 i_3226(.S(n_59764), .A(regs_6[25]), .B(sav_esi[25]), .Z(n_17332
		));
	notech_reg sav_esi_reg_26(.CP(n_62734), .D(n_17338), .CD(n_61565), .Q(sav_esi
		[26]));
	notech_mux2 i_3234(.S(n_59764), .A(regs_6[26]), .B(sav_esi[26]), .Z(n_17338
		));
	notech_reg sav_esi_reg_27(.CP(n_62734), .D(n_17344), .CD(n_61565), .Q(sav_esi
		[27]));
	notech_mux2 i_3242(.S(n_59764), .A(regs_6[27]), .B(sav_esi[27]), .Z(n_17344
		));
	notech_reg sav_esi_reg_28(.CP(n_62734), .D(n_17350), .CD(n_61565), .Q(sav_esi
		[28]));
	notech_mux2 i_3250(.S(n_59751), .A(regs_6[28]), .B(sav_esi[28]), .Z(n_17350
		));
	notech_nand3 i_358(.A(n_276391864), .B(n_273291893), .C(instrc[126]), .Z
		(n_2632));
	notech_reg sav_esi_reg_29(.CP(n_62734), .D(n_17356), .CD(n_61564), .Q(sav_esi
		[29]));
	notech_mux2 i_3258(.S(n_59751), .A(regs_6[29]), .B(sav_esi[29]), .Z(n_17356
		));
	notech_nand3 i_326(.A(n_273391892), .B(n_273091895), .C(instrc[68]), .Z(n_2631
		));
	notech_reg sav_esi_reg_30(.CP(n_62734), .D(n_17362), .CD(n_61564), .Q(sav_esi
		[30]));
	notech_mux2 i_3266(.S(n_59751), .A(regs_6[30]), .B(sav_esi[30]), .Z(n_17362
		));
	notech_reg sav_esi_reg_31(.CP(n_62734), .D(n_17368), .CD(n_61564), .Q(sav_esi
		[31]));
	notech_mux2 i_3274(.S(n_59751), .A(regs_6[31]), .B(sav_esi[31]), .Z(n_17368
		));
	notech_reg sav_edi_reg_0(.CP(n_62734), .D(n_17374), .CD(n_61564), .Q(sav_edi
		[0]));
	notech_mux2 i_3282(.S(n_59751), .A(regs_7[0]), .B(sav_edi[0]), .Z(n_17374
		));
	notech_and4 i_317(.A(vliw_pc[2]), .B(n_32843), .C(n_2739), .D(instrc[60]
		), .Z(n_2628));
	notech_reg sav_edi_reg_1(.CP(n_62734), .D(n_17380), .CD(n_61565), .Q(sav_edi
		[1]));
	notech_mux2 i_3290(.S(n_59751), .A(regs_7[1]), .B(sav_edi[1]), .Z(n_17380
		));
	notech_nand3 i_324(.A(n_273391892), .B(n_274591882), .C(instrc[4]), .Z(n_2627
		));
	notech_reg sav_edi_reg_2(.CP(n_62734), .D(n_17386), .CD(n_61565), .Q(sav_edi
		[2]));
	notech_mux2 i_3298(.S(n_59751), .A(regs_7[2]), .B(sav_edi[2]), .Z(n_17386
		));
	notech_reg sav_edi_reg_3(.CP(n_62668), .D(n_17392), .CD(n_61565), .Q(sav_edi
		[3]));
	notech_mux2 i_3306(.S(n_59751), .A(regs_7[3]), .B(sav_edi[3]), .Z(n_17392
		));
	notech_reg sav_edi_reg_4(.CP(n_62668), .D(n_17398), .CD(n_61565), .Q(sav_edi
		[4]));
	notech_mux2 i_3314(.S(n_59751), .A(regs_7[4]), .B(sav_edi[4]), .Z(n_17398
		));
	notech_reg sav_edi_reg_5(.CP(n_62668), .D(n_17404), .CD(n_61565), .Q(sav_edi
		[5]));
	notech_mux2 i_3322(.S(n_59751), .A(regs_7[5]), .B(sav_edi[5]), .Z(n_17404
		));
	notech_reg sav_edi_reg_6(.CP(n_62668), .D(n_17410), .CD(n_61542), .Q(sav_edi
		[6]));
	notech_mux2 i_3332(.S(n_59751), .A(regs_7[6]), .B(sav_edi[6]), .Z(n_17410
		));
	notech_reg sav_edi_reg_7(.CP(n_62668), .D(n_17416), .CD(n_61542), .Q(sav_edi
		[7]));
	notech_mux2 i_3340(.S(n_59751), .A(regs_7[7]), .B(sav_edi[7]), .Z(n_17416
		));
	notech_reg sav_edi_reg_8(.CP(n_62668), .D(n_17422), .CD(n_61542), .Q(sav_edi
		[8]));
	notech_mux2 i_3348(.S(n_59758), .A(regs_7[8]), .B(sav_edi[8]), .Z(n_17422
		));
	notech_reg sav_edi_reg_9(.CP(n_62668), .D(n_17428), .CD(n_61542), .Q(sav_edi
		[9]));
	notech_mux2 i_3356(.S(n_59758), .A(regs_7[9]), .B(sav_edi[9]), .Z(n_17428
		));
	notech_reg sav_edi_reg_10(.CP(n_62668), .D(n_17435), .CD(n_61542), .Q(sav_edi
		[10]));
	notech_mux2 i_3364(.S(n_59758), .A(regs_7[10]), .B(sav_edi[10]), .Z(n_17435
		));
	notech_nand3 i_328(.A(n_276391864), .B(n_273291893), .C(instrc[124]), .Z
		(n_2618));
	notech_reg sav_edi_reg_11(.CP(n_62668), .D(n_17442), .CD(n_61542), .Q(sav_edi
		[11]));
	notech_mux2 i_3372(.S(n_59758), .A(regs_7[11]), .B(sav_edi[11]), .Z(n_17442
		));
	notech_nand3 i_298(.A(n_273391892), .B(n_273091895), .C(instrc[69]), .Z(n_2617
		));
	notech_reg sav_edi_reg_12(.CP(n_62668), .D(n_17449), .CD(n_61542), .Q(sav_edi
		[12]));
	notech_mux2 i_3380(.S(n_59758), .A(regs_7[12]), .B(sav_edi[12]), .Z(n_17449
		));
	notech_reg sav_edi_reg_13(.CP(n_62668), .D(n_17457), .CD(n_61542), .Q(sav_edi
		[13]));
	notech_mux2 i_3388(.S(n_59758), .A(regs_7[13]), .B(sav_edi[13]), .Z(n_17457
		));
	notech_reg sav_edi_reg_14(.CP(n_62584), .D(n_17464), .CD(n_61542), .Q(sav_edi
		[14]));
	notech_mux2 i_3397(.S(n_59758), .A(regs_7[14]), .B(sav_edi[14]), .Z(n_17464
		));
	notech_and4 i_290(.A(vliw_pc[2]), .B(n_32843), .C(n_2739), .D(instrc[61]
		), .Z(n_2614));
	notech_reg sav_edi_reg_15(.CP(n_62528), .D(n_17471), .CD(n_61541), .Q(sav_edi
		[15]));
	notech_mux2 i_3406(.S(n_59758), .A(regs_7[15]), .B(sav_edi[15]), .Z(n_17471
		));
	notech_nand3 i_296(.A(n_273391892), .B(n_274591882), .C(instrc[5]), .Z(n_2613
		));
	notech_reg sav_edi_reg_16(.CP(n_62672), .D(n_17481), .CD(n_61541), .Q(sav_edi
		[16]));
	notech_mux2 i_3414(.S(n_59758), .A(regs_7[16]), .B(sav_edi[16]), .Z(n_17481
		));
	notech_reg sav_edi_reg_17(.CP(n_62586), .D(n_17488), .CD(n_61541), .Q(sav_edi
		[17]));
	notech_mux2 i_3422(.S(n_59758), .A(regs_7[17]), .B(sav_edi[17]), .Z(n_17488
		));
	notech_reg sav_edi_reg_18(.CP(n_62586), .D(n_17495), .CD(n_61541), .Q(sav_edi
		[18]));
	notech_mux2 i_3432(.S(n_59758), .A(regs_7[18]), .B(sav_edi[18]), .Z(n_17495
		));
	notech_reg sav_edi_reg_19(.CP(n_62586), .D(n_17502), .CD(n_61541), .Q(sav_edi
		[19]));
	notech_mux2 i_3441(.S(n_59758), .A(regs_7[19]), .B(sav_edi[19]), .Z(n_17502
		));
	notech_reg sav_edi_reg_20(.CP(n_62586), .D(n_17509), .CD(n_61541), .Q(sav_edi
		[20]));
	notech_mux2 i_3449(.S(n_59763), .A(regs_7[20]), .B(sav_edi[20]), .Z(n_17509
		));
	notech_reg sav_edi_reg_21(.CP(n_62586), .D(n_17517), .CD(n_61541), .Q(sav_edi
		[21]));
	notech_mux2 i_3457(.S(n_59763), .A(regs_7[21]), .B(sav_edi[21]), .Z(n_17517
		));
	notech_reg sav_edi_reg_22(.CP(n_62586), .D(n_17524), .CD(n_61541), .Q(sav_edi
		[22]));
	notech_mux2 i_3466(.S(n_59763), .A(regs_7[22]), .B(sav_edi[22]), .Z(n_17524
		));
	notech_reg sav_edi_reg_23(.CP(n_62586), .D(n_17531), .CD(n_61541), .Q(sav_edi
		[23]));
	notech_mux2 i_3475(.S(n_59763), .A(regs_7[23]), .B(sav_edi[23]), .Z(n_17531
		));
	notech_reg sav_edi_reg_24(.CP(n_62586), .D(n_17538), .CD(n_61541), .Q(sav_edi
		[24]));
	notech_mux2 i_3483(.S(n_59763), .A(regs_7[24]), .B(sav_edi[24]), .Z(n_17538
		));
	notech_nand3 i_300(.A(n_276391864), .B(n_273291893), .C(instrc[125]), .Z
		(n_2604));
	notech_reg sav_edi_reg_25(.CP(n_62586), .D(n_17545), .CD(n_61543), .Q(sav_edi
		[25]));
	notech_mux2 i_3492(.S(n_59763), .A(regs_7[25]), .B(sav_edi[25]), .Z(n_17545
		));
	notech_nand3 i_270(.A(n_273391892), .B(n_273091895), .C(instrc[71]), .Z(n_2603
		));
	notech_reg sav_edi_reg_26(.CP(n_62586), .D(n_17553), .CD(n_61543), .Q(sav_edi
		[26]));
	notech_mux2 i_3502(.S(n_59766), .A(regs_7[26]), .B(sav_edi[26]), .Z(n_17553
		));
	notech_reg sav_edi_reg_27(.CP(n_62672), .D(n_17560), .CD(n_61543), .Q(sav_edi
		[27]));
	notech_mux2 i_3513(.S(n_59766), .A(regs_7[27]), .B(sav_edi[27]), .Z(n_17560
		));
	notech_reg sav_edi_reg_28(.CP(n_62672), .D(n_17567), .CD(n_61543), .Q(sav_edi
		[28]));
	notech_mux2 i_3522(.S(n_59766), .A(regs_7[28]), .B(sav_edi[28]), .Z(n_17567
		));
	notech_and4 i_262(.A(vliw_pc[2]), .B(n_32843), .C(n_2739), .D(instrc[63]
		), .Z(n_2600));
	notech_reg sav_edi_reg_29(.CP(n_62672), .D(n_17574), .CD(n_61543), .Q(sav_edi
		[29]));
	notech_mux2 i_3533(.S(n_59766), .A(regs_7[29]), .B(sav_edi[29]), .Z(n_17574
		));
	notech_nand3 i_268(.A(n_273391892), .B(n_274591882), .C(instrc[7]), .Z(n_2599
		));
	notech_reg sav_edi_reg_30(.CP(n_62672), .D(n_17581), .CD(n_61544), .Q(sav_edi
		[30]));
	notech_mux2 i_3541(.S(n_59766), .A(regs_7[30]), .B(sav_edi[30]), .Z(n_17581
		));
	notech_reg sav_edi_reg_31(.CP(n_62672), .D(n_17589), .CD(n_61544), .Q(sav_edi
		[31]));
	notech_mux2 i_3549(.S(n_59766), .A(regs_7[31]), .B(sav_edi[31]), .Z(n_17589
		));
	notech_reg fepc_reg(.CP(n_62672), .D(n_17596), .CD(n_61543), .Q(fepc));
	notech_mux2 i_3557(.S(n_13726), .A(fepc), .B(n_13729), .Z(n_17596));
	notech_reg_set sav_epc_reg_0(.CP(n_62672), .D(n_17603), .SD(1'b1), .Q(sav_epc
		[0]));
	notech_mux2 i_3565(.S(n_27270), .A(sav_epc[0]), .B(regs_14[0]), .Z(n_17603
		));
	notech_reg_set sav_epc_reg_1(.CP(n_62672), .D(n_17610), .SD(1'b1), .Q(sav_epc
		[1]));
	notech_mux2 i_3573(.S(n_27270), .A(sav_epc[1]), .B(regs_14[1]), .Z(n_17610
		));
	notech_reg_set sav_epc_reg_2(.CP(n_62672), .D(n_17617), .SD(1'b1), .Q(sav_epc
		[2]));
	notech_mux2 i_3582(.S(n_27270), .A(sav_epc[2]), .B(regs_14[2]), .Z(n_17617
		));
	notech_reg_set sav_epc_reg_3(.CP(n_62672), .D(n_17624), .SD(1'b1), .Q(sav_epc
		[3]));
	notech_mux2 i_3590(.S(n_27270), .A(sav_epc[3]), .B(regs_14[3]), .Z(n_17624
		));
	notech_reg_set sav_epc_reg_4(.CP(n_62672), .D(n_17630), .SD(1'b1), .Q(sav_epc
		[4]));
	notech_mux2 i_3598(.S(n_27270), .A(sav_epc[4]), .B(regs_14[4]), .Z(n_17630
		));
	notech_reg_set sav_epc_reg_5(.CP(n_62672), .D(n_17636), .SD(1'b1), .Q(sav_epc
		[5]));
	notech_mux2 i_3606(.S(n_27270), .A(sav_epc[5]), .B(regs_14[5]), .Z(n_17636
		));
	notech_nand3 i_272(.A(n_276391864), .B(n_273291893), .C(instrc[127]), .Z
		(n_2590));
	notech_reg_set sav_epc_reg_6(.CP(n_62672), .D(n_17642), .SD(1'b1), .Q(sav_epc
		[6]));
	notech_mux2 i_3614(.S(n_27270), .A(sav_epc[6]), .B(regs_14[6]), .Z(n_17642
		));
	notech_nand3 i_241(.A(n_273391892), .B(n_273091895), .C(instrc[67]), .Z(n_2589
		));
	notech_reg_set sav_epc_reg_7(.CP(n_62672), .D(n_17648), .SD(1'b1), .Q(sav_epc
		[7]));
	notech_mux2 i_3622(.S(n_27270), .A(sav_epc[7]), .B(regs_14[7]), .Z(n_17648
		));
	notech_reg_set sav_epc_reg_8(.CP(n_62672), .D(n_17654), .SD(1'b1), .Q(sav_epc
		[8]));
	notech_mux2 i_3630(.S(n_27270), .A(sav_epc[8]), .B(regs_14[8]), .Z(n_17654
		));
	notech_reg_set sav_epc_reg_9(.CP(n_62672), .D(n_17660), .SD(1'b1), .Q(sav_epc
		[9]));
	notech_mux2 i_3638(.S(n_27270), .A(sav_epc[9]), .B(regs_14[9]), .Z(n_17660
		));
	notech_and4 i_233(.A(vliw_pc[2]), .B(n_32843), .C(n_2739), .D(instrc[59]
		), .Z(n_2586));
	notech_reg_set sav_epc_reg_10(.CP(n_62672), .D(n_17666), .SD(1'b1), .Q(sav_epc
		[10]));
	notech_mux2 i_3646(.S(n_27270), .A(sav_epc[10]), .B(regs_14[10]), .Z(n_17666
		));
	notech_nand3 i_239(.A(n_273391892), .B(n_274591882), .C(instrc[3]), .Z(n_2585
		));
	notech_reg_set sav_epc_reg_11(.CP(n_62672), .D(n_17672), .SD(1'b1), .Q(sav_epc
		[11]));
	notech_mux2 i_3654(.S(n_27270), .A(sav_epc[11]), .B(regs_14[11]), .Z(n_17672
		));
	notech_reg_set sav_epc_reg_12(.CP(n_62586), .D(n_17678), .SD(1'b1), .Q(sav_epc
		[12]));
	notech_mux2 i_3662(.S(n_27270), .A(sav_epc[12]), .B(regs_14[12]), .Z(n_17678
		));
	notech_reg_set sav_epc_reg_13(.CP(n_62586), .D(n_17684), .SD(1'b1), .Q(sav_epc
		[13]));
	notech_mux2 i_3670(.S(n_27270), .A(sav_epc[13]), .B(regs_14[13]), .Z(n_17684
		));
	notech_reg_set sav_epc_reg_14(.CP(n_62588), .D(n_17690), .SD(1'b1), .Q(sav_epc
		[14]));
	notech_mux2 i_3678(.S(n_27270), .A(sav_epc[14]), .B(regs_14[14]), .Z(n_17690
		));
	notech_reg_set sav_epc_reg_15(.CP(n_62588), .D(n_17696), .SD(1'b1), .Q(sav_epc
		[15]));
	notech_mux2 i_3686(.S(n_27270), .A(sav_epc[15]), .B(regs_14[15]), .Z(n_17696
		));
	notech_reg_set sav_epc_reg_16(.CP(n_62588), .D(n_17702), .SD(1'b1), .Q(sav_epc
		[16]));
	notech_mux2 i_3694(.S(n_54618), .A(sav_epc[16]), .B(regs_14[16]), .Z(n_17702
		));
	notech_reg_set sav_epc_reg_17(.CP(n_62588), .D(n_17708), .SD(1'b1), .Q(sav_epc
		[17]));
	notech_mux2 i_3702(.S(n_54618), .A(sav_epc[17]), .B(regs_14[17]), .Z(n_17708
		));
	notech_reg_set sav_epc_reg_18(.CP(n_62588), .D(n_17714), .SD(1'b1), .Q(sav_epc
		[18]));
	notech_mux2 i_3710(.S(n_54618), .A(sav_epc[18]), .B(regs_14[18]), .Z(n_17714
		));
	notech_reg_set sav_epc_reg_19(.CP(n_62588), .D(n_17720), .SD(1'b1), .Q(sav_epc
		[19]));
	notech_mux2 i_3718(.S(n_54618), .A(sav_epc[19]), .B(regs_14[19]), .Z(n_17720
		));
	notech_nand3 i_243(.A(n_276391864), .B(n_273291893), .C(instrc[123]), .Z
		(n_2576));
	notech_reg_set sav_epc_reg_20(.CP(n_62588), .D(n_17726), .SD(1'b1), .Q(sav_epc
		[20]));
	notech_mux2 i_3726(.S(n_54618), .A(sav_epc[20]), .B(regs_14[20]), .Z(n_17726
		));
	notech_nand3 i_208(.A(n_273391892), .B(n_273091895), .C(instrc[64]), .Z(n_2575
		));
	notech_reg_set sav_epc_reg_21(.CP(n_62588), .D(n_17732), .SD(1'b1), .Q(sav_epc
		[21]));
	notech_mux2 i_3734(.S(n_54618), .A(sav_epc[21]), .B(regs_14[21]), .Z(n_17732
		));
	notech_reg_set sav_epc_reg_22(.CP(n_62588), .D(n_17738), .SD(1'b1), .Q(sav_epc
		[22]));
	notech_mux2 i_3742(.S(n_54618), .A(sav_epc[22]), .B(regs_14[22]), .Z(n_17738
		));
	notech_reg_set sav_epc_reg_23(.CP(n_62588), .D(n_17744), .SD(1'b1), .Q(sav_epc
		[23]));
	notech_mux2 i_3750(.S(n_54618), .A(sav_epc[23]), .B(regs_14[23]), .Z(n_17744
		));
	notech_and4 i_200(.A(vliw_pc[2]), .B(n_32843), .C(n_2739), .D(instrc[56]
		), .Z(n_2572));
	notech_reg_set sav_epc_reg_24(.CP(n_62588), .D(n_17750), .SD(1'b1), .Q(sav_epc
		[24]));
	notech_mux2 i_3758(.S(n_54618), .A(sav_epc[24]), .B(regs_14[24]), .Z(n_17750
		));
	notech_nand3 i_206(.A(n_273391892), .B(n_274591882), .C(instrc[0]), .Z(n_2571
		));
	notech_reg_set sav_epc_reg_25(.CP(n_62588), .D(n_17756), .SD(1'b1), .Q(sav_epc
		[25]));
	notech_mux2 i_3766(.S(n_54618), .A(sav_epc[25]), .B(regs_14[25]), .Z(n_17756
		));
	notech_reg_set sav_epc_reg_26(.CP(n_62588), .D(n_17762), .SD(1'b1), .Q(sav_epc
		[26]));
	notech_mux2 i_3774(.S(n_54618), .A(sav_epc[26]), .B(regs_14[26]), .Z(n_17762
		));
	notech_reg_set sav_epc_reg_27(.CP(n_62588), .D(n_17768), .SD(1'b1), .Q(sav_epc
		[27]));
	notech_mux2 i_3782(.S(n_54618), .A(sav_epc[27]), .B(regs_14[27]), .Z(n_17768
		));
	notech_reg_set sav_epc_reg_28(.CP(n_62588), .D(n_17774), .SD(1'b1), .Q(sav_epc
		[28]));
	notech_mux2 i_3790(.S(n_54618), .A(sav_epc[28]), .B(regs_14[28]), .Z(n_17774
		));
	notech_reg_set sav_epc_reg_29(.CP(n_62588), .D(n_17781), .SD(1'b1), .Q(sav_epc
		[29]));
	notech_mux2 i_3798(.S(n_54618), .A(sav_epc[29]), .B(regs_14[29]), .Z(n_17781
		));
	notech_reg_set sav_epc_reg_30(.CP(n_62588), .D(n_17788), .SD(1'b1), .Q(sav_epc
		[30]));
	notech_mux2 i_3806(.S(n_54618), .A(sav_epc[30]), .B(regs_14[30]), .Z(n_17788
		));
	notech_reg_set sav_epc_reg_31(.CP(n_62588), .D(n_17795), .SD(1'b1), .Q(sav_epc
		[31]));
	notech_mux2 i_3814(.S(n_54618), .A(sav_epc[31]), .B(regs_14[31]), .Z(n_17795
		));
	notech_reg_set all_cnt_reg_0(.CP(n_62588), .D(n_17802), .SD(1'b1), .Q(all_cnt
		[0]));
	notech_mux2 i_3822(.S(\nbus_11299[0] ), .A(all_cnt[0]), .B(n_27111), .Z(n_17802
		));
	notech_reg_set all_cnt_reg_1(.CP(n_62528), .D(n_17809), .SD(1'b1), .Q(all_cnt
		[1]));
	notech_mux2 i_3830(.S(\nbus_11299[0] ), .A(all_cnt[1]), .B(n_27271), .Z(n_17809
		));
	notech_nand3 i_210(.A(n_276391864), .B(n_273291893), .C(instrc[120]), .Z
		(n_2562));
	notech_reg_set all_cnt_reg_2(.CP(n_62528), .D(n_17817), .SD(1'b1), .Q(all_cnt
		[2]));
	notech_mux2 i_3838(.S(\nbus_11299[0] ), .A(all_cnt[2]), .B(n_46191246), 
		.Z(n_17817));
	notech_nor2 i_327962(.A(n_60969), .B(n_60958), .Z(n_2561));
	notech_reg_set all_cnt_reg_3(.CP(n_62528), .D(n_17824), .SD(1'b1), .Q(all_cnt
		[3]));
	notech_mux2 i_3846(.S(\nbus_11299[0] ), .A(all_cnt[3]), .B(n_46291247), 
		.Z(n_17824));
	notech_nand3 i_180(.A(n_273391892), .B(n_273091895), .C(instrc[66]), .Z(n_2560
		));
	notech_reg regs_reg_14_0(.CP(n_62528), .D(n_17831), .CD(n_61543), .Q(regs_14
		[0]));
	notech_mux2 i_3854(.S(n_3906), .A(n_24756), .B(regs_14[0]), .Z(n_17831)
		);
	notech_reg regs_reg_14_1(.CP(n_62528), .D(n_17838), .CD(n_61543), .Q(regs_14
		[1]));
	notech_mux2 i_3862(.S(n_3906), .A(n_24762), .B(regs_14[1]), .Z(n_17838)
		);
	notech_reg regs_reg_14_2(.CP(n_62528), .D(n_17845), .CD(n_61542), .Q(regs_14
		[2]));
	notech_mux2 i_3870(.S(n_3906), .A(n_24768), .B(regs_14[2]), .Z(n_17845)
		);
	notech_and4 i_172(.A(vliw_pc[2]), .B(n_32843), .C(n_2739), .D(instrc[58]
		), .Z(n_2557));
	notech_reg regs_reg_14_3(.CP(n_62528), .D(n_17853), .CD(n_61542), .Q(regs_14
		[3]));
	notech_mux2 i_3878(.S(n_3906), .A(n_24774), .B(regs_14[3]), .Z(n_17853)
		);
	notech_nand3 i_178(.A(n_273391892), .B(n_274591882), .C(instrc[2]), .Z(n_2556
		));
	notech_reg regs_reg_14_4(.CP(n_62528), .D(n_17860), .CD(n_61542), .Q(regs_14
		[4]));
	notech_mux2 i_3886(.S(n_3906), .A(n_24780), .B(regs_14[4]), .Z(n_17860)
		);
	notech_reg regs_reg_14_5(.CP(n_62528), .D(n_17867), .CD(n_61542), .Q(regs_14
		[5]));
	notech_mux2 i_3894(.S(n_3906), .A(n_24786), .B(regs_14[5]), .Z(n_17867)
		);
	notech_reg regs_reg_14_6(.CP(n_62528), .D(n_17874), .CD(n_61543), .Q(regs_14
		[6]));
	notech_mux2 i_3902(.S(n_3906), .A(n_24792), .B(regs_14[6]), .Z(n_17874)
		);
	notech_reg regs_reg_14_7(.CP(n_62668), .D(n_17881), .CD(n_61543), .Q(regs_14
		[7]));
	notech_mux2 i_3910(.S(n_3906), .A(n_24798), .B(regs_14[7]), .Z(n_17881)
		);
	notech_reg regs_reg_14_8(.CP(n_62526), .D(n_17889), .CD(n_61543), .Q(regs_14
		[8]));
	notech_mux2 i_3918(.S(n_3906), .A(n_24804), .B(regs_14[8]), .Z(n_17889)
		);
	notech_reg regs_reg_14_9(.CP(n_62526), .D(n_17896), .CD(n_61543), .Q(regs_14
		[9]));
	notech_mux2 i_3926(.S(n_3906), .A(n_24810), .B(regs_14[9]), .Z(n_17896)
		);
	notech_reg_set regs_reg_14_10(.CP(n_62576), .D(n_17903), .SD(n_61543), .Q
		(regs_14[10]));
	notech_mux2 i_3934(.S(n_3906), .A(n_24816), .B(regs_14[10]), .Z(n_17903)
		);
	notech_reg_set regs_reg_14_11(.CP(n_62576), .D(n_17910), .SD(n_61538), .Q
		(regs_14[11]));
	notech_mux2 i_3942(.S(n_3906), .A(n_24822), .B(regs_14[11]), .Z(n_17910)
		);
	notech_reg_set regs_reg_14_12(.CP(n_62576), .D(n_17917), .SD(n_61538), .Q
		(regs_14[12]));
	notech_mux2 i_3950(.S(n_3906), .A(n_24828), .B(regs_14[12]), .Z(n_17917)
		);
	notech_and3 i_182(.A(n_276391864), .B(n_273291893), .C(n_60975), .Z(n_2547
		));
	notech_reg_set regs_reg_14_13(.CP(n_62576), .D(n_17925), .SD(n_61538), .Q
		(regs_14[13]));
	notech_mux2 i_3958(.S(n_3906), .A(n_24834), .B(regs_14[13]), .Z(n_17925)
		);
	notech_and4 i_227961(.A(n_276591862), .B(n_2774), .C(n_2545), .D(n_2532)
		, .Z(n_2546));
	notech_reg_set regs_reg_14_14(.CP(n_62576), .D(n_17932), .SD(n_61538), .Q
		(regs_14[14]));
	notech_mux2 i_3966(.S(n_3906), .A(n_24840), .B(regs_14[14]), .Z(n_17932)
		);
	notech_nand3 i_150(.A(n_273391892), .B(n_273091895), .C(instrc[65]), .Z(n_2545
		));
	notech_reg_set regs_reg_14_15(.CP(n_62576), .D(n_17939), .SD(n_61538), .Q
		(regs_14[15]));
	notech_mux2 i_3974(.S(n_3906), .A(n_24846), .B(regs_14[15]), .Z(n_17939)
		);
	notech_reg_set regs_reg_14_16(.CP(n_62576), .D(n_17946), .SD(n_61538), .Q
		(regs_14[16]));
	notech_mux2 i_3982(.S(n_56210), .A(n_24852), .B(regs_14[16]), .Z(n_17946
		));
	notech_reg_set regs_reg_14_17(.CP(n_62576), .D(n_17953), .SD(n_61538), .Q
		(regs_14[17]));
	notech_mux2 i_3990(.S(n_56210), .A(n_24858), .B(regs_14[17]), .Z(n_17953
		));
	notech_and4 i_142(.A(vliw_pc[2]), .B(n_32843), .C(n_2739), .D(instrc[57]
		), .Z(n_2542));
	notech_reg_set regs_reg_14_18(.CP(n_62576), .D(n_17961), .SD(n_61538), .Q
		(regs_14[18]));
	notech_mux2 i_3998(.S(n_56210), .A(n_24864), .B(regs_14[18]), .Z(n_17961
		));
	notech_nand3 i_148(.A(n_273391892), .B(n_274591882), .C(instrc[1]), .Z(n_2541
		));
	notech_reg_set regs_reg_14_19(.CP(n_62576), .D(n_17968), .SD(n_61538), .Q
		(regs_14[19]));
	notech_mux2 i_4006(.S(n_56210), .A(n_24870), .B(regs_14[19]), .Z(n_17968
		));
	notech_reg regs_reg_14_20(.CP(n_62660), .D(n_17974), .CD(n_61538), .Q(regs_14
		[20]));
	notech_mux2 i_4014(.S(n_56210), .A(n_24876), .B(regs_14[20]), .Z(n_17974
		));
	notech_reg regs_reg_14_21(.CP(n_62660), .D(n_17980), .CD(n_61537), .Q(regs_14
		[21]));
	notech_mux2 i_4022(.S(n_56210), .A(n_24882), .B(regs_14[21]), .Z(n_17980
		));
	notech_reg regs_reg_14_22(.CP(n_62660), .D(n_17986), .CD(n_61537), .Q(regs_14
		[22]));
	notech_mux2 i_4030(.S(n_56210), .A(n_24888), .B(regs_14[22]), .Z(n_17986
		));
	notech_reg regs_reg_14_23(.CP(n_62660), .D(n_17992), .CD(n_61537), .Q(regs_14
		[23]));
	notech_mux2 i_4038(.S(n_56210), .A(n_24894), .B(regs_14[23]), .Z(n_17992
		));
	notech_reg regs_reg_14_24(.CP(n_62660), .D(n_17998), .CD(n_61537), .Q(regs_14
		[24]));
	notech_mux2 i_4046(.S(n_56210), .A(n_24900), .B(regs_14[24]), .Z(n_17998
		));
	notech_reg regs_reg_14_25(.CP(n_62660), .D(n_18004), .CD(n_61537), .Q(regs_14
		[25]));
	notech_mux2 i_4054(.S(n_56210), .A(n_24906), .B(regs_14[25]), .Z(n_18004
		));
	notech_reg regs_reg_14_26(.CP(n_62660), .D(n_18010), .CD(n_61537), .Q(regs_14
		[26]));
	notech_mux2 i_4062(.S(n_56210), .A(n_24912), .B(regs_14[26]), .Z(n_18010
		));
	notech_reg regs_reg_14_27(.CP(n_62660), .D(n_18016), .CD(n_61537), .Q(regs_14
		[27]));
	notech_mux2 i_4070(.S(n_56210), .A(n_24918), .B(regs_14[27]), .Z(n_18016
		));
	notech_nand3 i_152(.A(n_276391864), .B(n_273291893), .C(n_60915), .Z(n_2532
		));
	notech_reg regs_reg_14_28(.CP(n_62660), .D(n_18022), .CD(n_61537), .Q(regs_14
		[28]));
	notech_mux2 i_4078(.S(n_56210), .A(n_24924), .B(regs_14[28]), .Z(n_18022
		));
	notech_nao3 i_111(.A(n_29655), .B(n_18972), .C(n_3806), .Z(n_2531));
	notech_reg regs_reg_14_29(.CP(n_62660), .D(n_18028), .CD(n_61537), .Q(regs_14
		[29]));
	notech_mux2 i_4086(.S(n_56210), .A(n_1512), .B(regs_14[29]), .Z(n_18028)
		);
	notech_ao3 i_96(.A(n_1869), .B(n_23007), .C(n_2683), .Z(n_2530));
	notech_reg regs_reg_14_30(.CP(n_62660), .D(n_18034), .CD(n_61539), .Q(regs_14
		[30]));
	notech_mux2 i_4094(.S(n_56210), .A(n_24936), .B(regs_14[30]), .Z(n_18034
		));
	notech_mux2 i_65(.S(n_60316), .A(n_266891921), .B(n_1880), .Z(n_2529));
	notech_reg regs_reg_14_31(.CP(n_62660), .D(n_18040), .CD(n_61539), .Q(regs_14
		[31]));
	notech_mux2 i_4102(.S(n_56210), .A(n_24942), .B(regs_14[31]), .Z(n_18040
		));
	notech_or4 i_32071(.A(n_27125), .B(n_62870), .C(\opcode[3] ), .D(n_32695
		), .Z(n_27904));
	notech_reg regs_reg_13_0(.CP(n_62660), .D(n_18046), .CD(n_61539), .Q(gs[
		0]));
	notech_mux2 i_4110(.S(\nbus_11374[0] ), .A(gs[0]), .B(n_27275), .Z(n_18046
		));
	notech_reg regs_reg_13_1(.CP(n_62660), .D(n_18052), .CD(n_61539), .Q(gs[
		1]));
	notech_mux2 i_4118(.S(\nbus_11374[0] ), .A(gs[1]), .B(n_24436), .Z(n_18052
		));
	notech_reg regs_reg_13_2(.CP(n_62660), .D(n_18058), .CD(n_61539), .Q(gs[
		2]));
	notech_mux2 i_4126(.S(\nbus_11374[0] ), .A(n_56005), .B(n_24442), .Z(n_18058
		));
	notech_ao4 i_76532082(.A(write_ack), .B(n_318591638), .C(n_28533), .D(n_27084
		), .Z(n_2526));
	notech_reg regs_reg_13_3(.CP(n_62660), .D(n_18064), .CD(n_61541), .Q(gs[
		3]));
	notech_mux2 i_4134(.S(\nbus_11374[0] ), .A(gs[3]), .B(n_24448), .Z(n_18064
		));
	notech_and4 i_77032077(.A(n_242891974), .B(n_2524), .C(n_242991973), .D(n_243091972
		), .Z(n_2525));
	notech_reg regs_reg_13_4(.CP(n_62660), .D(n_18070), .CD(n_61541), .Q(gs[
		4]));
	notech_mux2 i_4142(.S(\nbus_11374[0] ), .A(gs[4]), .B(n_24454), .Z(n_18070
		));
	notech_ao4 i_76732080(.A(n_2359), .B(n_61133), .C(n_2358), .D(n_61109), 
		.Z(n_2524));
	notech_reg regs_reg_13_5(.CP(n_62660), .D(n_18076), .CD(n_61539), .Q(gs[
		5]));
	notech_mux2 i_4150(.S(\nbus_11374[0] ), .A(gs[5]), .B(n_24460), .Z(n_18076
		));
	notech_and4 i_77332074(.A(n_22015), .B(n_59115), .C(n_59106), .D(n_318491639
		), .Z(n_2523));
	notech_reg regs_reg_13_6(.CP(n_62660), .D(n_18082), .CD(n_61541), .Q(gs[
		6]));
	notech_mux2 i_4158(.S(\nbus_11374[0] ), .A(gs[6]), .B(n_24466), .Z(n_18082
		));
	notech_reg regs_reg_13_7(.CP(n_62658), .D(n_18088), .CD(n_61539), .Q(gs[
		7]));
	notech_mux2 i_4166(.S(\nbus_11374[0] ), .A(gs[7]), .B(n_24472), .Z(n_18088
		));
	notech_reg regs_reg_13_8(.CP(n_62658), .D(n_18094), .CD(n_61538), .Q(gs[
		8]));
	notech_mux2 i_4174(.S(\nbus_11374[0] ), .A(gs[8]), .B(n_27276), .Z(n_18094
		));
	notech_reg regs_reg_13_9(.CP(n_62730), .D(n_18100), .CD(n_61539), .Q(gs[
		9]));
	notech_mux2 i_4182(.S(\nbus_11374[0] ), .A(gs[9]), .B(n_27277), .Z(n_18100
		));
	notech_reg regs_reg_13_10(.CP(n_62730), .D(n_18106), .CD(n_61538), .Q(gs
		[10]));
	notech_mux2 i_4190(.S(\nbus_11374[0] ), .A(gs[10]), .B(n_27278), .Z(n_18106
		));
	notech_ao4 i_77532072(.A(n_2363), .B(n_60372), .C(n_2362), .D(n_25641), 
		.Z(n_2518));
	notech_reg regs_reg_13_11(.CP(n_62730), .D(n_18112), .CD(n_61538), .Q(gs
		[11]));
	notech_mux2 i_4198(.S(\nbus_11374[0] ), .A(gs[11]), .B(n_24496), .Z(n_18112
		));
	notech_reg regs_reg_13_12(.CP(n_62730), .D(n_18118), .CD(n_61539), .Q(gs
		[12]));
	notech_mux2 i_4206(.S(\nbus_11374[0] ), .A(gs[12]), .B(n_27279), .Z(n_18118
		));
	notech_reg regs_reg_13_13(.CP(n_62730), .D(n_18124), .CD(n_61539), .Q(gs
		[13]));
	notech_mux2 i_4214(.S(\nbus_11374[0] ), .A(gs[13]), .B(n_24508), .Z(n_18124
		));
	notech_reg regs_reg_13_14(.CP(n_62730), .D(n_18130), .CD(n_61539), .Q(gs
		[14]));
	notech_mux2 i_4222(.S(\nbus_11374[0] ), .A(gs[14]), .B(n_24514), .Z(n_18130
		));
	notech_reg regs_reg_13_15(.CP(n_62730), .D(n_18137), .CD(n_61539), .Q(gs
		[15]));
	notech_mux2 i_4231(.S(\nbus_11374[0] ), .A(gs[15]), .B(n_27281), .Z(n_18137
		));
	notech_reg regs_reg_13_16(.CP(n_62730), .D(n_18145), .CD(n_61539), .Q(gs
		[16]));
	notech_mux2 i_4240(.S(n_54687), .A(gs[16]), .B(n_27282), .Z(n_18145));
	notech_reg regs_reg_13_17(.CP(n_62730), .D(n_18152), .CD(n_61550), .Q(gs
		[17]));
	notech_mux2 i_4248(.S(n_54687), .A(gs[17]), .B(n_27283), .Z(n_18152));
	notech_reg regs_reg_13_18(.CP(n_62730), .D(n_18159), .CD(n_61550), .Q(gs
		[18]));
	notech_mux2 i_4256(.S(n_54687), .A(gs[18]), .B(n_27284), .Z(n_18159));
	notech_or4 i_102131846(.A(n_61175), .B(n_61160), .C(n_61151), .D(n_308891735
		), .Z(n_2510));
	notech_reg regs_reg_13_19(.CP(n_62730), .D(n_18166), .CD(n_61549), .Q(gs
		[19]));
	notech_mux2 i_4264(.S(n_54687), .A(gs[19]), .B(n_27285), .Z(n_18166));
	notech_reg regs_reg_13_20(.CP(n_62730), .D(n_18173), .CD(n_61549), .Q(gs
		[20]));
	notech_mux2 i_4272(.S(n_54687), .A(gs[20]), .B(n_27286), .Z(n_18173));
	notech_ao4 i_103731831(.A(n_59095), .B(n_19065), .C(n_2370), .D(n_61109)
		, .Z(n_2508));
	notech_reg regs_reg_13_21(.CP(n_62730), .D(n_18181), .CD(n_61550), .Q(gs
		[21]));
	notech_mux2 i_4280(.S(n_54687), .A(gs[21]), .B(n_27287), .Z(n_18181));
	notech_reg regs_reg_13_22(.CP(n_62730), .D(n_18188), .CD(n_61550), .Q(gs
		[22]));
	notech_mux2 i_4288(.S(n_54687), .A(gs[22]), .B(n_27288), .Z(n_18188));
	notech_reg regs_reg_13_23(.CP(n_62730), .D(n_18195), .CD(n_61550), .Q(gs
		[23]));
	notech_mux2 i_4296(.S(n_54687), .A(gs[23]), .B(n_27290), .Z(n_18195));
	notech_reg regs_reg_13_24(.CP(n_62730), .D(n_18202), .CD(n_61550), .Q(gs
		[24]));
	notech_mux2 i_4304(.S(n_54687), .A(gs[24]), .B(n_27291), .Z(n_18202));
	notech_ao4 i_103931829(.A(n_56570), .B(n_28558), .C(n_56666), .D(n_28255
		), .Z(n_2505));
	notech_reg regs_reg_13_25(.CP(n_62730), .D(n_18209), .CD(n_61550), .Q(gs
		[25]));
	notech_mux2 i_4312(.S(n_54687), .A(gs[25]), .B(n_27292), .Z(n_18209));
	notech_ao4 i_104031828(.A(n_56653), .B(n_28220), .C(n_56916), .D(n_29624
		), .Z(n_2504));
	notech_reg regs_reg_13_26(.CP(n_62730), .D(n_18217), .CD(n_61549), .Q(gs
		[26]));
	notech_mux2 i_4320(.S(n_54687), .A(gs[26]), .B(n_24586), .Z(n_18217));
	notech_and2 i_104431824(.A(n_2502), .B(n_2501), .Z(n_2503));
	notech_reg regs_reg_13_27(.CP(n_62658), .D(n_18224), .CD(n_61549), .Q(gs
		[27]));
	notech_mux2 i_4328(.S(n_54687), .A(gs[27]), .B(n_24592), .Z(n_18224));
	notech_ao4 i_104231826(.A(n_56640), .B(n_28287), .C(n_56532), .D(n_28320
		), .Z(n_2502));
	notech_reg regs_reg_13_28(.CP(n_62658), .D(n_18231), .CD(n_61549), .Q(gs
		[28]));
	notech_mux2 i_4336(.S(n_54687), .A(gs[28]), .B(n_24598), .Z(n_18231));
	notech_ao4 i_104331825(.A(n_56518), .B(n_29625), .C(n_56502), .D(n_28385
		), .Z(n_2501));
	notech_reg regs_reg_13_29(.CP(n_62658), .D(n_18238), .CD(n_61549), .Q(gs
		[29]));
	notech_mux2 i_4344(.S(n_54687), .A(gs[29]), .B(n_24604), .Z(n_18238));
	notech_and4 i_105231816(.A(n_2498), .B(n_2497), .C(n_2495), .D(n_2494), 
		.Z(n_2500));
	notech_reg regs_reg_13_30(.CP(n_62658), .D(n_18245), .CD(n_61549), .Q(gs
		[30]));
	notech_mux2 i_4352(.S(n_54687), .A(gs[30]), .B(n_27294), .Z(n_18245));
	notech_reg regs_reg_13_31(.CP(n_62658), .D(n_18253), .CD(n_61549), .Q(gs
		[31]));
	notech_mux2 i_4360(.S(n_54687), .A(gs[31]), .B(n_27295), .Z(n_18253));
	notech_ao4 i_104631822(.A(n_56489), .B(n_28353), .C(n_56627), .D(n_28449
		), .Z(n_2498));
	notech_reg regs_reg_12_0(.CP(n_62658), .D(n_18260), .CD(n_61549), .Q(regs_12
		[0]));
	notech_mux2 i_4368(.S(\nbus_11373[0] ), .A(regs_12[0]), .B(n_27296), .Z(n_18260
		));
	notech_ao4 i_104731821(.A(n_56605), .B(n_28481), .C(n_56553), .D(n_27892
		), .Z(n_2497));
	notech_reg regs_reg_12_1(.CP(n_62658), .D(n_18267), .CD(n_61549), .Q(regs_12
		[1]));
	notech_mux2 i_4376(.S(\nbus_11373[0] ), .A(regs_12[1]), .B(n_24088), .Z(n_18267
		));
	notech_reg regs_reg_12_2(.CP(n_62658), .D(n_18274), .CD(n_61549), .Q(regs_12
		[2]));
	notech_mux2 i_4384(.S(\nbus_11373[0] ), .A(regs_12[2]), .B(n_24094), .Z(n_18274
		));
	notech_ao4 i_104931819(.A(n_56547), .B(n_28591), .C(n_56592), .D(n_28188
		), .Z(n_2495));
	notech_reg regs_reg_12_3(.CP(n_62658), .D(n_18281), .CD(n_61549), .Q(regs_12
		[3]));
	notech_mux2 i_4392(.S(\nbus_11373[0] ), .A(regs_12[3]), .B(n_24100), .Z(n_18281
		));
	notech_ao4 i_105031818(.A(n_56614), .B(n_28417), .C(n_56583), .D(n_28514
		), .Z(n_2494));
	notech_reg regs_reg_12_4(.CP(n_62658), .D(n_18289), .CD(n_61552), .Q(regs_12
		[4]));
	notech_mux2 i_4400(.S(\nbus_11373[0] ), .A(regs_12[4]), .B(n_24106), .Z(n_18289
		));
	notech_reg regs_reg_12_5(.CP(n_62730), .D(n_18296), .CD(n_61552), .Q(regs_12
		[5]));
	notech_mux2 i_4408(.S(\nbus_11373[0] ), .A(regs_12[5]), .B(n_24112), .Z(n_18296
		));
	notech_ao3 i_31632471(.A(n_60139), .B(n_60207), .C(n_26580), .Z(n_2492)
		);
	notech_reg regs_reg_12_6(.CP(n_62726), .D(n_18303), .CD(n_61552), .Q(regs_12
		[6]));
	notech_mux2 i_4416(.S(\nbus_11373[0] ), .A(regs_12[6]), .B(n_27299), .Z(n_18303
		));
	notech_ao4 i_105531813(.A(n_2489), .B(all_cnt[3]), .C(n_246791942), .D(n_59364
		), .Z(n_2491));
	notech_reg regs_reg_12_7(.CP(n_62656), .D(n_18310), .CD(n_61552), .Q(regs_12
		[7]));
	notech_mux2 i_4424(.S(\nbus_11373[0] ), .A(regs_12[7]), .B(n_24124), .Z(n_18310
		));
	notech_ao4 i_105631812(.A(n_2379), .B(n_2380), .C(n_2378), .D(n_27192), 
		.Z(n_2490));
	notech_reg regs_reg_12_8(.CP(n_62726), .D(n_18317), .CD(n_61552), .Q(regs_12
		[8]));
	notech_mux2 i_4432(.S(\nbus_11373[0] ), .A(regs_12[8]), .B(n_24130), .Z(n_18317
		));
	notech_xor2 i_1030373(.A(n_59373), .B(n_246791942), .Z(n_2489));
	notech_reg regs_reg_12_9(.CP(n_62726), .D(n_18324), .CD(n_61552), .Q(regs_12
		[9]));
	notech_mux2 i_4440(.S(\nbus_11373[0] ), .A(regs_12[9]), .B(n_24136), .Z(n_18324
		));
	notech_nor2 i_530394(.A(n_2350), .B(n_2355), .Z(n_2488));
	notech_reg regs_reg_12_10(.CP(n_62726), .D(n_18330), .CD(n_61552), .Q(regs_12
		[10]));
	notech_mux2 i_4448(.S(\nbus_11373[0] ), .A(regs_12[10]), .B(n_24142), .Z
		(n_18330));
	notech_or4 i_2130206(.A(n_245991950), .B(n_245891951), .C(n_246091949), 
		.D(n_27558), .Z(n_3848598));
	notech_reg regs_reg_12_11(.CP(n_62726), .D(n_18336), .CD(n_61552), .Q(regs_12
		[11]));
	notech_mux2 i_4456(.S(\nbus_11373[0] ), .A(regs_12[11]), .B(n_24148), .Z
		(n_18336));
	notech_ao4 i_106731802(.A(n_27198), .B(n_27577), .C(n_59373), .D(n_27856
		), .Z(n_2487));
	notech_reg regs_reg_12_12(.CP(n_62726), .D(n_18342), .CD(n_61552), .Q(regs_12
		[12]));
	notech_mux2 i_4464(.S(\nbus_11373[0] ), .A(regs_12[12]), .B(n_24154), .Z
		(n_18342));
	notech_reg regs_reg_12_13(.CP(n_62726), .D(n_18348), .CD(n_61552), .Q(regs_12
		[13]));
	notech_mux2 i_4472(.S(\nbus_11373[0] ), .A(regs_12[13]), .B(n_24160), .Z
		(n_18348));
	notech_reg regs_reg_12_14(.CP(n_62726), .D(n_18354), .CD(n_61550), .Q(regs_12
		[14]));
	notech_mux2 i_4480(.S(\nbus_11373[0] ), .A(regs_12[14]), .B(n_24166), .Z
		(n_18354));
	notech_ao4 i_107031799(.A(n_59393), .B(n_27853), .C(n_59407), .D(n_27854
		), .Z(n_2484));
	notech_reg regs_reg_12_15(.CP(n_62726), .D(n_18360), .CD(n_61550), .Q(regs_12
		[15]));
	notech_mux2 i_4488(.S(\nbus_11373[0] ), .A(regs_12[15]), .B(n_24172), .Z
		(n_18360));
	notech_ao4 i_107131798(.A(n_27853), .B(n_27198), .C(n_59407), .D(n_27113
		), .Z(n_2483));
	notech_reg regs_reg_12_16(.CP(n_62726), .D(n_18366), .CD(n_61550), .Q(regs_12
		[16]));
	notech_mux2 i_4496(.S(n_54698), .A(regs_12[16]), .B(n_27303), .Z(n_18366
		));
	notech_ao4 i_10732632(.A(n_59373), .B(n_27852), .C(n_27856), .D(n_2481),
		 .Z(n_2482));
	notech_reg regs_reg_12_17(.CP(n_62726), .D(n_18372), .CD(n_61550), .Q(regs_12
		[17]));
	notech_mux2 i_4504(.S(n_54698), .A(regs_12[17]), .B(n_24184), .Z(n_18372
		));
	notech_and2 i_5332679(.A(n_59382), .B(n_27852), .Z(n_2481));
	notech_reg regs_reg_12_18(.CP(n_62726), .D(n_18378), .CD(n_61550), .Q(regs_12
		[18]));
	notech_mux2 i_4512(.S(n_54698), .A(regs_12[18]), .B(n_24190), .Z(n_18378
		));
	notech_or4 i_19032579(.A(n_61175), .B(n_61160), .C(n_61151), .D(n_32378)
		, .Z(n_2480));
	notech_reg regs_reg_12_19(.CP(n_62758), .D(n_18384), .CD(n_61552), .Q(regs_12
		[19]));
	notech_mux2 i_4520(.S(n_54698), .A(regs_12[19]), .B(n_24196), .Z(n_18384
		));
	notech_nand2 i_198932690(.A(n_59382), .B(n_59364), .Z(n_2479));
	notech_reg regs_reg_12_20(.CP(n_62758), .D(n_18390), .CD(n_61552), .Q(regs_12
		[20]));
	notech_mux2 i_4528(.S(n_54698), .A(regs_12[20]), .B(n_24202), .Z(n_18390
		));
	notech_or4 i_28932494(.A(n_32567), .B(n_26580), .C(n_19050), .D(n_19036)
		, .Z(n_4668680));
	notech_reg regs_reg_12_21(.CP(n_62758), .D(n_18396), .CD(n_61550), .Q(regs_12
		[21]));
	notech_mux2 i_4536(.S(n_54698), .A(regs_12[21]), .B(n_24208), .Z(n_18396
		));
	notech_and2 i_30532478(.A(n_27123), .B(n_32470), .Z(n_2478));
	notech_reg regs_reg_12_22(.CP(n_62758), .D(n_18402), .CD(n_61552), .Q(regs_12
		[22]));
	notech_mux2 i_4544(.S(n_54698), .A(regs_12[22]), .B(n_24214), .Z(n_18402
		));
	notech_reg regs_reg_12_23(.CP(n_62758), .D(n_18408), .CD(n_61547), .Q(regs_12
		[23]));
	notech_mux2 i_4552(.S(n_54698), .A(regs_12[23]), .B(n_24220), .Z(n_18408
		));
	notech_and4 i_30232481(.A(n_32432), .B(n_1897), .C(n_1898), .D(n_2354), 
		.Z(n_4758689));
	notech_reg regs_reg_12_24(.CP(n_62758), .D(n_18414), .CD(n_61547), .Q(regs_12
		[24]));
	notech_mux2 i_4560(.S(n_54698), .A(regs_12[24]), .B(n_24226), .Z(n_18414
		));
	notech_reg regs_reg_12_25(.CP(n_62758), .D(n_18420), .CD(n_61544), .Q(regs_12
		[25]));
	notech_mux2 i_4568(.S(n_54698), .A(regs_12[25]), .B(n_24232), .Z(n_18420
		));
	notech_reg regs_reg_12_26(.CP(n_62758), .D(n_18426), .CD(n_61547), .Q(regs_12
		[26]));
	notech_mux2 i_4576(.S(n_54698), .A(regs_12[26]), .B(n_24238), .Z(n_18426
		));
	notech_reg regs_reg_12_27(.CP(n_62758), .D(n_18432), .CD(n_61547), .Q(regs_12
		[27]));
	notech_mux2 i_4584(.S(n_54698), .A(regs_12[27]), .B(n_24244), .Z(n_18432
		));
	notech_reg regs_reg_12_28(.CP(n_62758), .D(n_18438), .CD(n_61547), .Q(regs_12
		[28]));
	notech_mux2 i_4592(.S(n_54698), .A(regs_12[28]), .B(n_24250), .Z(n_18438
		));
	notech_reg regs_reg_12_29(.CP(n_62758), .D(n_18444), .CD(n_61547), .Q(regs_12
		[29]));
	notech_mux2 i_4600(.S(n_54698), .A(regs_12[29]), .B(n_24256), .Z(n_18444
		));
	notech_or4 i_26132516(.A(n_4978711), .B(n_62836), .C(n_60931), .D(\opcode[3] 
		), .Z(n_4958709));
	notech_reg regs_reg_12_30(.CP(n_62758), .D(n_18450), .CD(n_61547), .Q(regs_12
		[30]));
	notech_mux2 i_4608(.S(n_54698), .A(regs_12[30]), .B(n_27307), .Z(n_18450
		));
	notech_reg regs_reg_12_31(.CP(n_62758), .D(n_18456), .CD(n_61547), .Q(regs_12
		[31]));
	notech_mux2 i_4616(.S(n_54698), .A(regs_12[31]), .B(n_24268), .Z(n_18456
		));
	notech_nand2 i_21032560(.A(n_2825), .B(n_2864), .Z(n_4978711));
	notech_reg regs_reg_11_0(.CP(n_62758), .D(n_18462), .CD(n_61544), .Q(regs_11
		[0]));
	notech_mux2 i_4624(.S(\nbus_11372[0] ), .A(regs_11[0]), .B(n_27308), .Z(n_18462
		));
	notech_nao3 i_26432513(.A(n_19117), .B(n_26761), .C(n_19109), .Z(n_5018715
		));
	notech_reg regs_reg_11_1(.CP(n_62758), .D(n_18468), .CD(n_61544), .Q(regs_11
		[1]));
	notech_mux2 i_4632(.S(\nbus_11372[0] ), .A(regs_11[1]), .B(n_23740), .Z(n_18468
		));
	notech_reg regs_reg_11_2(.CP(n_62758), .D(n_18474), .CD(n_61544), .Q(regs_11
		[2]));
	notech_mux2 i_4640(.S(\nbus_11372[0] ), .A(regs_11[2]), .B(n_23746), .Z(n_18474
		));
	notech_nor2 i_201332704(.A(n_59382), .B(n_59373), .Z(n_246991940));
	notech_reg regs_reg_11_3(.CP(n_62758), .D(n_18481), .CD(n_61544), .Q(regs_11
		[3]));
	notech_mux2 i_4648(.S(\nbus_11372[0] ), .A(regs_11[3]), .B(n_23752), .Z(n_18481
		));
	notech_or2 i_195232693(.A(n_59407), .B(n_29177), .Z(n_246891941));
	notech_reg regs_reg_11_4(.CP(n_62758), .D(n_18488), .CD(n_61544), .Q(regs_11
		[4]));
	notech_mux2 i_4656(.S(\nbus_11372[0] ), .A(regs_11[4]), .B(n_23758), .Z(n_18488
		));
	notech_nand2 i_194132695(.A(n_59407), .B(n_59393), .Z(n_246791942));
	notech_reg regs_reg_11_5(.CP(n_62726), .D(n_18495), .CD(n_61544), .Q(regs_11
		[5]));
	notech_mux2 i_4664(.S(\nbus_11372[0] ), .A(regs_11[5]), .B(n_23764), .Z(n_18495
		));
	notech_and2 i_193632696(.A(all_cnt[1]), .B(all_cnt[2]), .Z(n_6858899));
	notech_reg regs_reg_11_6(.CP(n_62758), .D(n_18502), .CD(n_61544), .Q(regs_11
		[6]));
	notech_mux2 i_4672(.S(\nbus_11372[0] ), .A(regs_11[6]), .B(n_27309), .Z(n_18502
		));
	notech_nao3 i_138331506(.A(calc_sz[0]), .B(n_27895), .C(calc_sz[3]), .Z(n_246691943
		));
	notech_reg regs_reg_11_7(.CP(n_62728), .D(n_18509), .CD(n_61544), .Q(regs_11
		[7]));
	notech_mux2 i_4680(.S(\nbus_11372[0] ), .A(regs_11[7]), .B(n_23776), .Z(n_18509
		));
	notech_reg regs_reg_11_8(.CP(n_62728), .D(n_18517), .CD(n_61544), .Q(regs_11
		[8]));
	notech_mux2 i_4688(.S(\nbus_11372[0] ), .A(regs_11[8]), .B(n_27310), .Z(n_18517
		));
	notech_and3 i_27581(.A(n_57020), .B(n_57042), .C(n_57078), .Z(n_246591944
		));
	notech_reg regs_reg_11_9(.CP(n_62728), .D(n_18524), .CD(n_61544), .Q(regs_11
		[9]));
	notech_mux2 i_4696(.S(\nbus_11372[0] ), .A(regs_11[9]), .B(n_27311), .Z(n_18524
		));
	notech_or4 i_27718(.A(n_62844), .B(n_32729), .C(n_32259), .D(n_60931), .Z
		(n_32257));
	notech_reg regs_reg_11_10(.CP(n_62728), .D(n_18531), .CD(n_61548), .Q(regs_11
		[10]));
	notech_mux2 i_4704(.S(\nbus_11372[0] ), .A(regs_11[10]), .B(n_27312), .Z
		(n_18531));
	notech_reg regs_reg_11_11(.CP(n_62728), .D(n_18538), .CD(n_61548), .Q(regs_11
		[11]));
	notech_mux2 i_4712(.S(\nbus_11372[0] ), .A(regs_11[11]), .B(n_23800), .Z
		(n_18538));
	notech_ao4 i_26632511(.A(n_32351), .B(n_32373), .C(n_56843), .D(n_61133)
		, .Z(n_32350));
	notech_reg regs_reg_11_12(.CP(n_62728), .D(n_18545), .CD(n_61548), .Q(regs_11
		[12]));
	notech_mux2 i_4720(.S(\nbus_11372[0] ), .A(regs_11[12]), .B(n_27313), .Z
		(n_18545));
	notech_reg regs_reg_11_13(.CP(n_62728), .D(n_18553), .CD(n_61548), .Q(regs_11
		[13]));
	notech_mux2 i_4728(.S(\nbus_11372[0] ), .A(regs_11[13]), .B(n_23812), .Z
		(n_18553));
	notech_reg regs_reg_11_14(.CP(n_62728), .D(n_18561), .CD(n_61548), .Q(regs_11
		[14]));
	notech_mux2 i_4736(.S(\nbus_11372[0] ), .A(regs_11[14]), .B(n_23818), .Z
		(n_18561));
	notech_reg regs_reg_11_15(.CP(n_62728), .D(n_18568), .CD(n_61548), .Q(regs_11
		[15]));
	notech_mux2 i_4744(.S(\nbus_11372[0] ), .A(regs_11[15]), .B(n_27314), .Z
		(n_18568));
	notech_reg regs_reg_11_16(.CP(n_62728), .D(n_18575), .CD(n_61549), .Q(regs_11
		[16]));
	notech_mux2 i_4752(.S(n_54745), .A(regs_11[16]), .B(n_27315), .Z(n_18575
		));
	notech_reg regs_reg_11_17(.CP(n_62728), .D(n_18583), .CD(n_61548), .Q(regs_11
		[17]));
	notech_mux2 i_4760(.S(n_54745), .A(regs_11[17]), .B(n_27316), .Z(n_18583
		));
	notech_and2 i_59832235(.A(n_318791636), .B(n_27571), .Z(n_246091949));
	notech_reg regs_reg_11_18(.CP(n_62728), .D(n_18591), .CD(n_61548), .Q(regs_11
		[18]));
	notech_mux2 i_4768(.S(n_54745), .A(regs_11[18]), .B(n_27317), .Z(n_18591
		));
	notech_ao4 i_59732236(.A(n_6858899), .B(n_27563), .C(n_59286), .D(n_27571
		), .Z(n_245991950));
	notech_reg regs_reg_11_19(.CP(n_62728), .D(n_18599), .CD(n_61548), .Q(regs_11
		[19]));
	notech_mux2 i_4776(.S(n_54745), .A(regs_11[19]), .B(n_27318), .Z(n_18599
		));
	notech_ao4 i_59632237(.A(n_2406), .B(n_27566), .C(all_cnt[3]), .D(n_59364
		), .Z(n_245891951));
	notech_reg regs_reg_11_20(.CP(n_62728), .D(n_18607), .CD(n_61547), .Q(regs_11
		[20]));
	notech_mux2 i_4784(.S(n_54745), .A(regs_11[20]), .B(n_27320), .Z(n_18607
		));
	notech_reg regs_reg_11_21(.CP(n_62728), .D(n_18614), .CD(n_61547), .Q(regs_11
		[21]));
	notech_mux2 i_4792(.S(n_54745), .A(regs_11[21]), .B(n_27321), .Z(n_18614
		));
	notech_reg regs_reg_11_22(.CP(n_62728), .D(n_18621), .CD(n_61547), .Q(regs_11
		[22]));
	notech_mux2 i_4800(.S(n_54745), .A(regs_11[22]), .B(n_23866), .Z(n_18621
		));
	notech_reg regs_reg_11_23(.CP(n_62728), .D(n_18628), .CD(n_61547), .Q(regs_11
		[23]));
	notech_mux2 i_4808(.S(n_54745), .A(regs_11[23]), .B(n_23872), .Z(n_18628
		));
	notech_reg regs_reg_11_24(.CP(n_62728), .D(n_18635), .CD(n_61547), .Q(regs_11
		[24]));
	notech_mux2 i_4816(.S(n_54745), .A(regs_11[24]), .B(n_23878), .Z(n_18635
		));
	notech_reg regs_reg_11_25(.CP(n_62728), .D(n_18643), .CD(n_61548), .Q(regs_11
		[25]));
	notech_mux2 i_4824(.S(n_54745), .A(regs_11[25]), .B(n_23884), .Z(n_18643
		));
	notech_reg regs_reg_11_26(.CP(n_62656), .D(n_18650), .CD(n_61548), .Q(regs_11
		[26]));
	notech_mux2 i_4832(.S(n_54745), .A(regs_11[26]), .B(n_23890), .Z(n_18650
		));
	notech_reg regs_reg_11_27(.CP(n_62656), .D(n_18657), .CD(n_61548), .Q(regs_11
		[27]));
	notech_mux2 i_4840(.S(n_54745), .A(regs_11[27]), .B(n_23896), .Z(n_18657
		));
	notech_reg regs_reg_11_28(.CP(n_62656), .D(n_18664), .CD(n_61548), .Q(regs_11
		[28]));
	notech_mux2 i_4848(.S(n_54745), .A(regs_11[28]), .B(n_23902), .Z(n_18664
		));
	notech_reg regs_reg_11_29(.CP(n_62656), .D(n_18671), .CD(n_61592), .Q(regs_11
		[29]));
	notech_mux2 i_4856(.S(n_54745), .A(regs_11[29]), .B(n_23908), .Z(n_18671
		));
	notech_reg regs_reg_11_30(.CP(n_62656), .D(n_18677), .CD(n_61592), .Q(regs_11
		[30]));
	notech_mux2 i_4864(.S(n_54745), .A(regs_11[30]), .B(n_23914), .Z(n_18677
		));
	notech_reg regs_reg_11_31(.CP(n_62656), .D(n_18683), .CD(n_61592), .Q(regs_11
		[31]));
	notech_mux2 i_4872(.S(n_54745), .A(regs_11[31]), .B(n_23920), .Z(n_18683
		));
	notech_reg regs_reg_10_0(.CP(n_62656), .D(n_18689), .CD(n_61592), .Q(regs_10
		[0]));
	notech_mux2 i_4880(.S(\nbus_11302[0] ), .A(regs_10[0]), .B(n_27322), .Z(n_18689
		));
	notech_reg regs_reg_10_1(.CP(n_62656), .D(n_18695), .CD(n_61592), .Q(regs_10
		[1]));
	notech_mux2 i_4889(.S(\nbus_11302[0] ), .A(regs_10[1]), .B(n_13980), .Z(n_18695
		));
	notech_reg regs_reg_10_2(.CP(n_62656), .D(n_18701), .CD(n_61593), .Q(regs_10
		[2]));
	notech_mux2 i_4897(.S(\nbus_11302[0] ), .A(regs_10[2]), .B(n_13986), .Z(n_18701
		));
	notech_reg regs_reg_10_3(.CP(n_62656), .D(n_18707), .CD(n_61593), .Q(regs_10
		[3]));
	notech_mux2 i_4905(.S(\nbus_11302[0] ), .A(regs_10[3]), .B(n_13992), .Z(n_18707
		));
	notech_reg regs_reg_10_4(.CP(n_62576), .D(n_18713), .CD(n_61592), .Q(regs_10
		[4]));
	notech_mux2 i_4913(.S(\nbus_11302[0] ), .A(regs_10[4]), .B(n_13998), .Z(n_18713
		));
	notech_reg regs_reg_10_5(.CP(n_62656), .D(n_18719), .CD(n_61592), .Q(regs_10
		[5]));
	notech_mux2 i_4921(.S(\nbus_11302[0] ), .A(regs_10[5]), .B(n_14004), .Z(n_18719
		));
	notech_reg regs_reg_10_6(.CP(n_62662), .D(n_18725), .CD(n_61592), .Q(regs_10
		[6]));
	notech_mux2 i_4929(.S(\nbus_11302[0] ), .A(regs_10[6]), .B(n_14010), .Z(n_18725
		));
	notech_reg regs_reg_10_7(.CP(n_62578), .D(n_18731), .CD(n_61589), .Q(regs_10
		[7]));
	notech_mux2 i_4937(.S(\nbus_11302[0] ), .A(regs_10[7]), .B(n_14016), .Z(n_18731
		));
	notech_reg regs_reg_10_8(.CP(n_62578), .D(n_18737), .CD(n_61589), .Q(regs_10
		[8]));
	notech_mux2 i_4945(.S(\nbus_11302[0] ), .A(regs_10[8]), .B(n_27323), .Z(n_18737
		));
	notech_reg regs_reg_10_9(.CP(n_62578), .D(n_18743), .CD(n_61589), .Q(regs_10
		[9]));
	notech_mux2 i_4953(.S(\nbus_11302[0] ), .A(regs_10[9]), .B(n_27324), .Z(n_18743
		));
	notech_reg regs_reg_10_10(.CP(n_62578), .D(n_18749), .CD(n_61589), .Q(regs_10
		[10]));
	notech_mux2 i_4961(.S(\nbus_11302[0] ), .A(regs_10[10]), .B(n_27325), .Z
		(n_18749));
	notech_reg regs_reg_10_11(.CP(n_62578), .D(n_18755), .CD(n_61592), .Q(regs_10
		[11]));
	notech_mux2 i_4969(.S(\nbus_11302[0] ), .A(regs_10[11]), .B(n_14040), .Z
		(n_18755));
	notech_reg regs_reg_10_12(.CP(n_62578), .D(n_18761), .CD(n_61592), .Q(regs_10
		[12]));
	notech_mux2 i_4977(.S(\nbus_11302[0] ), .A(regs_10[12]), .B(n_27326), .Z
		(n_18761));
	notech_or4 i_55032281(.A(n_61109), .B(n_2893), .C(n_62836), .D(n_60933),
		 .Z(n_243491968));
	notech_reg regs_reg_10_13(.CP(n_62578), .D(n_18767), .CD(n_61592), .Q(regs_10
		[13]));
	notech_mux2 i_4985(.S(\nbus_11302[0] ), .A(regs_10[13]), .B(n_14052), .Z
		(n_18767));
	notech_nand2 i_27723(.A(n_62776), .B(opc[30]), .Z(n_32252));
	notech_reg regs_reg_10_14(.CP(n_62578), .D(n_18773), .CD(n_61592), .Q(regs_10
		[14]));
	notech_mux2 i_4993(.S(\nbus_11302[0] ), .A(regs_10[14]), .B(n_14058), .Z
		(n_18773));
	notech_nand2 i_34264(.A(n_19137), .B(n_60207), .Z(n_25641));
	notech_reg regs_reg_10_15(.CP(n_62578), .D(n_18779), .CD(n_61592), .Q(regs_10
		[15]));
	notech_mux2 i_5001(.S(\nbus_11302[0] ), .A(regs_10[15]), .B(n_27327), .Z
		(n_18779));
	notech_nand3 i_34265(.A(n_60378), .B(n_3794), .C(n_61151), .Z(n_25640)
		);
	notech_reg regs_reg_10_16(.CP(n_62578), .D(n_18785), .CD(n_61594), .Q(regs_10
		[16]));
	notech_mux2 i_5009(.S(n_54783), .A(regs_10[16]), .B(n_27328), .Z(n_18785
		));
	notech_reg regs_reg_10_17(.CP(n_62664), .D(n_18791), .CD(n_61594), .Q(regs_10
		[17]));
	notech_mux2 i_5017(.S(n_54783), .A(regs_10[17]), .B(n_27330), .Z(n_18791
		));
	notech_reg regs_reg_10_18(.CP(n_62664), .D(n_18797), .CD(n_61593), .Q(regs_10
		[18]));
	notech_mux2 i_5025(.S(n_54783), .A(regs_10[18]), .B(n_27331), .Z(n_18797
		));
	notech_nao3 i_39832403(.A(n_60207), .B(n_29655), .C(n_19137), .Z(n_243191971
		));
	notech_reg regs_reg_10_19(.CP(n_62664), .D(n_18803), .CD(n_61594), .Q(regs_10
		[19]));
	notech_mux2 i_5033(.S(n_54783), .A(regs_10[19]), .B(n_27332), .Z(n_18803
		));
	notech_or4 i_38932412(.A(n_32581), .B(n_2357), .C(n_26900), .D(n_61133),
		 .Z(n_243091972));
	notech_reg regs_reg_10_20(.CP(n_62664), .D(n_18809), .CD(n_61594), .Q(regs_10
		[20]));
	notech_mux2 i_5041(.S(n_54783), .A(regs_10[20]), .B(n_14094), .Z(n_18809
		));
	notech_or4 i_38732413(.A(n_3806), .B(n_32579), .C(n_1878), .D(n_29655), 
		.Z(n_242991973));
	notech_reg regs_reg_10_21(.CP(n_62664), .D(n_18815), .CD(n_61594), .Q(regs_10
		[21]));
	notech_mux2 i_5049(.S(n_54783), .A(regs_10[21]), .B(n_27333), .Z(n_18815
		));
	notech_or4 i_38632414(.A(n_32403), .B(n_26999), .C(read_ack), .D(n_32567
		), .Z(n_242891974));
	notech_reg regs_reg_10_22(.CP(n_62664), .D(n_18821), .CD(n_61594), .Q(regs_10
		[22]));
	notech_mux2 i_5057(.S(n_54783), .A(regs_10[22]), .B(n_14106), .Z(n_18821
		));
	notech_reg regs_reg_10_23(.CP(n_62664), .D(n_18827), .CD(n_61594), .Q(regs_10
		[23]));
	notech_mux2 i_5065(.S(n_54783), .A(regs_10[23]), .B(n_14112), .Z(n_18827
		));
	notech_reg regs_reg_10_24(.CP(n_62664), .D(n_18834), .CD(n_61594), .Q(regs_10
		[24]));
	notech_mux2 i_5073(.S(n_54783), .A(regs_10[24]), .B(n_14118), .Z(n_18834
		));
	notech_reg regs_reg_10_25(.CP(n_62664), .D(n_18842), .CD(n_61593), .Q(regs_10
		[25]));
	notech_mux2 i_5081(.S(n_54783), .A(regs_10[25]), .B(n_14124), .Z(n_18842
		));
	notech_reg regs_reg_10_26(.CP(n_62664), .D(n_18849), .CD(n_61593), .Q(regs_10
		[26]));
	notech_mux2 i_5089(.S(n_54783), .A(regs_10[26]), .B(n_216059241), .Z(n_18849
		));
	notech_reg regs_reg_10_27(.CP(n_62664), .D(n_18856), .CD(n_61593), .Q(regs_10
		[27]));
	notech_mux2 i_5097(.S(n_54783), .A(regs_10[27]), .B(n_14136), .Z(n_18856
		));
	notech_reg regs_reg_10_28(.CP(n_62664), .D(n_18863), .CD(n_61593), .Q(regs_10
		[28]));
	notech_mux2 i_5105(.S(n_54783), .A(regs_10[28]), .B(n_215159232), .Z(n_18863
		));
	notech_reg regs_reg_10_29(.CP(n_62664), .D(n_18870), .CD(n_61593), .Q(regs_10
		[29]));
	notech_mux2 i_5113(.S(n_54783), .A(regs_10[29]), .B(n_14148), .Z(n_18870
		));
	notech_reg regs_reg_10_30(.CP(n_62664), .D(n_18878), .CD(n_61593), .Q(regs_10
		[30]));
	notech_mux2 i_5121(.S(n_54783), .A(regs_10[30]), .B(n_14154), .Z(n_18878
		));
	notech_or4 i_64232193(.A(n_59478), .B(n_62794), .C(n_60904), .D(n_27573)
		, .Z(n_2419));
	notech_reg regs_reg_10_31(.CP(n_62664), .D(n_18885), .CD(n_61593), .Q(regs_10
		[31]));
	notech_mux2 i_5129(.S(n_54783), .A(regs_10[31]), .B(n_14160), .Z(n_18885
		));
	notech_reg regs_reg_9_0(.CP(n_62664), .D(n_18892), .CD(n_61593), .Q(cs[0
		]));
	notech_mux2 i_5137(.S(\nbus_11335[0] ), .A(cs[0]), .B(n_27336), .Z(n_18892
		));
	notech_nand2 i_61632218(.A(n_317091653), .B(n_32350), .Z(n_2417));
	notech_reg regs_reg_9_1(.CP(n_62664), .D(n_18899), .CD(n_61593), .Q(cs[1
		]));
	notech_mux2 i_5145(.S(\nbus_11335[0] ), .A(cs[1]), .B(n_18835), .Z(n_18899
		));
	notech_reg regs_reg_9_2(.CP(n_62664), .D(n_18906), .CD(n_61593), .Q(\nbus_14523[2] 
		));
	notech_mux2 i_5153(.S(\nbus_11335[0] ), .A(\nbus_14523[2] ), .B(n_27337)
		, .Z(n_18906));
	notech_reg regs_reg_9_3(.CP(n_62664), .D(n_18914), .CD(n_61587), .Q(\nbus_14523[3] 
		));
	notech_mux2 i_5161(.S(\nbus_11335[0] ), .A(\nbus_14523[3] ), .B(n_18847)
		, .Z(n_18914));
	notech_nand2 i_61232222(.A(n_23513), .B(n_23514), .Z(n_2414));
	notech_reg regs_reg_9_4(.CP(n_62732), .D(n_18921), .CD(n_61587), .Q(\nbus_14523[4] 
		));
	notech_mux2 i_5169(.S(\nbus_11335[0] ), .A(\nbus_14523[4] ), .B(n_18853)
		, .Z(n_18921));
	notech_reg regs_reg_9_5(.CP(n_62662), .D(n_18928), .CD(n_61587), .Q(\nbus_14523[5] 
		));
	notech_mux2 i_5177(.S(\nbus_11335[0] ), .A(\nbus_14523[5] ), .B(n_18859)
		, .Z(n_18928));
	notech_reg regs_reg_9_6(.CP(n_62732), .D(n_18935), .CD(n_61587), .Q(\nbus_14523[6] 
		));
	notech_mux2 i_5185(.S(\nbus_11335[0] ), .A(\nbus_14523[6] ), .B(n_18865)
		, .Z(n_18935));
	notech_reg regs_reg_9_7(.CP(n_62732), .D(n_18942), .CD(n_61587), .Q(\nbus_14523[7] 
		));
	notech_mux2 i_5193(.S(\nbus_11335[0] ), .A(\nbus_14523[7] ), .B(n_18871)
		, .Z(n_18942));
	notech_reg regs_reg_9_8(.CP(n_62732), .D(n_18950), .CD(n_61588), .Q(\nbus_14523[8] 
		));
	notech_mux2 i_5201(.S(\nbus_11335[0] ), .A(\nbus_14523[8] ), .B(n_18877)
		, .Z(n_18950));
	notech_reg regs_reg_9_9(.CP(n_62732), .D(n_18957), .CD(n_61588), .Q(\nbus_14523[9] 
		));
	notech_mux2 i_5209(.S(\nbus_11335[0] ), .A(\nbus_14523[9] ), .B(n_27338)
		, .Z(n_18957));
	notech_reg regs_reg_9_10(.CP(n_62732), .D(n_18965), .CD(n_61587), .Q(\nbus_14523[10] 
		));
	notech_mux2 i_5217(.S(\nbus_11335[0] ), .A(\nbus_14523[10] ), .B(n_18889
		), .Z(n_18965));
	notech_reg regs_reg_9_11(.CP(n_62732), .D(n_18974), .CD(n_61588), .Q(\nbus_14523[11] 
		));
	notech_mux2 i_5225(.S(\nbus_11335[0] ), .A(\nbus_14523[11] ), .B(n_18895
		), .Z(n_18974));
	notech_nor2 i_60232232(.A(n_59397), .B(n_27854), .Z(n_2406));
	notech_reg regs_reg_9_12(.CP(n_62732), .D(n_18982), .CD(n_61587), .Q(\nbus_14523[12] 
		));
	notech_mux2 i_5233(.S(\nbus_11335[0] ), .A(\nbus_14523[12] ), .B(n_18901
		), .Z(n_18982));
	notech_reg regs_reg_9_13(.CP(n_62732), .D(n_18990), .CD(n_61586), .Q(\nbus_14523[13] 
		));
	notech_mux2 i_5241(.S(\nbus_11335[0] ), .A(\nbus_14523[13] ), .B(n_18907
		), .Z(n_18990));
	notech_reg regs_reg_9_14(.CP(n_62732), .D(n_18999), .CD(n_61587), .Q(\nbus_14523[14] 
		));
	notech_mux2 i_5249(.S(\nbus_11335[0] ), .A(\nbus_14523[14] ), .B(n_18913
		), .Z(n_18999));
	notech_reg regs_reg_9_15(.CP(n_62732), .D(n_19007), .CD(n_61586), .Q(\nbus_14523[15] 
		));
	notech_mux2 i_5258(.S(\nbus_11335[0] ), .A(\nbus_14523[15] ), .B(n_18919
		), .Z(n_19007));
	notech_reg regs_reg_9_16(.CP(n_62732), .D(n_19016), .CD(n_61586), .Q(\nbus_14523[16] 
		));
	notech_mux2 i_5266(.S(n_56872), .A(\nbus_14523[16] ), .B(n_18925), .Z(n_19016
		));
	notech_reg regs_reg_9_17(.CP(n_62732), .D(n_19023), .CD(n_61587), .Q(\nbus_14523[17] 
		));
	notech_mux2 i_5274(.S(n_56872), .A(\nbus_14523[17] ), .B(n_18931), .Z(n_19023
		));
	notech_reg regs_reg_9_18(.CP(n_62732), .D(n_19030), .CD(n_61587), .Q(\nbus_14523[18] 
		));
	notech_mux2 i_5282(.S(n_56872), .A(\nbus_14523[18] ), .B(n_18937), .Z(n_19030
		));
	notech_reg regs_reg_9_19(.CP(n_62732), .D(n_19037), .CD(n_61587), .Q(\nbus_14523[19] 
		));
	notech_mux2 i_5290(.S(n_56872), .A(\nbus_14523[19] ), .B(n_18943), .Z(n_19037
		));
	notech_reg regs_reg_9_20(.CP(n_62732), .D(n_19044), .CD(n_61587), .Q(\nbus_14523[20] 
		));
	notech_mux2 i_5298(.S(n_56872), .A(\nbus_14523[20] ), .B(n_27339), .Z(n_19044
		));
	notech_reg regs_reg_9_21(.CP(n_62732), .D(n_19051), .CD(n_61587), .Q(\nbus_14523[21] 
		));
	notech_mux2 i_5306(.S(n_56872), .A(\nbus_14523[21] ), .B(n_18955), .Z(n_19051
		));
	notech_reg regs_reg_9_22(.CP(n_62732), .D(n_19058), .CD(n_61589), .Q(\nbus_14523[22] 
		));
	notech_mux2 i_5315(.S(n_56872), .A(\nbus_14523[22] ), .B(n_27341), .Z(n_19058
		));
	notech_reg regs_reg_9_23(.CP(n_62732), .D(n_19064), .CD(n_61589), .Q(\nbus_14523[23] 
		));
	notech_mux2 i_5326(.S(n_56872), .A(\nbus_14523[23] ), .B(n_27342), .Z(n_19064
		));
	notech_reg regs_reg_9_24(.CP(n_62662), .D(n_19071), .CD(n_61589), .Q(\nbus_14523[24] 
		));
	notech_mux2 i_5337(.S(n_56872), .A(\nbus_14523[24] ), .B(n_27343), .Z(n_19071
		));
	notech_reg regs_reg_9_25(.CP(n_62662), .D(n_19078), .CD(n_61589), .Q(\nbus_14523[25] 
		));
	notech_mux2 i_5345(.S(n_56872), .A(\nbus_14523[25] ), .B(n_27345), .Z(n_19078
		));
	notech_reg regs_reg_9_26(.CP(n_62662), .D(n_19085), .CD(n_61589), .Q(\nbus_14523[26] 
		));
	notech_mux2 i_5353(.S(n_56872), .A(\nbus_14523[26] ), .B(n_18985), .Z(n_19085
		));
	notech_reg regs_reg_9_27(.CP(n_62662), .D(n_19092), .CD(n_61589), .Q(\nbus_14523[27] 
		));
	notech_mux2 i_5361(.S(n_56872), .A(\nbus_14523[27] ), .B(n_18991), .Z(n_19092
		));
	notech_reg regs_reg_9_28(.CP(n_62662), .D(n_19099), .CD(n_61589), .Q(\nbus_14523[28] 
		));
	notech_mux2 i_5369(.S(n_56872), .A(\nbus_14523[28] ), .B(n_18997), .Z(n_19099
		));
	notech_and2 i_28432497(.A(all_cnt[1]), .B(n_27572), .Z(n_2389));
	notech_reg regs_reg_9_29(.CP(n_62662), .D(n_19107), .CD(n_61589), .Q(\nbus_14523[29] 
		));
	notech_mux2 i_5377(.S(n_56872), .A(\nbus_14523[29] ), .B(n_19003), .Z(n_19107
		));
	notech_reg regs_reg_9_30(.CP(n_62662), .D(n_19115), .CD(n_61589), .Q(\nbus_14523[30] 
		));
	notech_mux2 i_5385(.S(n_56872), .A(\nbus_14523[30] ), .B(n_27347), .Z(n_19115
		));
	notech_ao4 i_37832422(.A(n_59407), .B(n_2389), .C(all_cnt[1]), .D(n_27572
		), .Z(n_2387));
	notech_reg regs_reg_9_31(.CP(n_62662), .D(n_19123), .CD(n_61588), .Q(\nbus_14523[31] 
		));
	notech_mux2 i_5393(.S(n_56872), .A(\nbus_14523[31] ), .B(n_27350), .Z(n_19123
		));
	notech_and2 i_13832603(.A(n_27192), .B(all_cnt[2]), .Z(n_2386));
	notech_reg regs_reg_8_0(.CP(n_62662), .D(n_19132), .CD(n_61588), .Q(regs_8
		[0]));
	notech_mux2 i_5401(.S(n_27365), .A(regs_8[0]), .B(n_27351), .Z(n_19132)
		);
	notech_reg regs_reg_8_1(.CP(n_62662), .D(n_19140), .CD(n_61588), .Q(regs_8
		[1]));
	notech_mux2 i_5409(.S(n_27365), .A(regs_8[1]), .B(n_18486), .Z(n_19140)
		);
	notech_ao3 i_37732423(.A(all_cnt[1]), .B(all_cnt[2]), .C(n_2481), .Z(n_2384
		));
	notech_reg regs_reg_8_2(.CP(n_62578), .D(n_19147), .CD(n_61588), .Q(regs_8
		[2]));
	notech_mux2 i_5417(.S(n_27365), .A(regs_8[2]), .B(n_18492), .Z(n_19147)
		);
	notech_reg regs_reg_8_3(.CP(n_62578), .D(n_19155), .CD(n_61588), .Q(regs_8
		[3]));
	notech_mux2 i_5425(.S(n_27365), .A(regs_8[3]), .B(n_18498), .Z(n_19155)
		);
	notech_reg regs_reg_8_4(.CP(n_62666), .D(n_19162), .CD(n_61588), .Q(regs_8
		[4]));
	notech_mux2 i_5433(.S(n_27365), .A(regs_8[4]), .B(n_18504), .Z(n_19162)
		);
	notech_or2 i_57732256(.A(n_2489), .B(all_cnt[2]), .Z(n_2381));
	notech_reg regs_reg_8_5(.CP(n_62580), .D(n_19169), .CD(n_61588), .Q(regs_8
		[5]));
	notech_mux2 i_5441(.S(n_27365), .A(regs_8[5]), .B(n_18510), .Z(n_19169)
		);
	notech_and2 i_24132533(.A(n_2489), .B(all_cnt[3]), .Z(n_2380));
	notech_reg regs_reg_8_6(.CP(n_62580), .D(n_19176), .CD(n_61588), .Q(regs_8
		[6]));
	notech_mux2 i_5449(.S(n_27365), .A(regs_8[6]), .B(n_27354), .Z(n_19176)
		);
	notech_ao4 i_6432675(.A(n_2387), .B(n_2386), .C(n_59275), .D(n_2384), .Z
		(n_2379));
	notech_reg regs_reg_8_7(.CP(n_62580), .D(n_19183), .CD(n_61588), .Q(regs_8
		[7]));
	notech_mux2 i_5457(.S(n_27365), .A(regs_8[7]), .B(n_18522), .Z(n_19183)
		);
	notech_and2 i_27532504(.A(n_27070), .B(n_2381), .Z(n_2378));
	notech_reg regs_reg_8_8(.CP(n_62580), .D(n_19191), .CD(n_61588), .Q(regs_8
		[8]));
	notech_mux2 i_5465(.S(n_27365), .A(regs_8[8]), .B(n_27355), .Z(n_19191)
		);
	notech_reg regs_reg_8_9(.CP(n_62580), .D(n_19198), .CD(n_61599), .Q(regs_8
		[9]));
	notech_mux2 i_5473(.S(n_27365), .A(regs_8[9]), .B(n_27356), .Z(n_19198)
		);
	notech_and2 i_35832441(.A(n_2491), .B(n_2490), .Z(n_2376));
	notech_reg regs_reg_8_10(.CP(n_62580), .D(n_19205), .CD(n_61599), .Q(regs_8
		[10]));
	notech_mux2 i_5481(.S(n_27365), .A(regs_8[10]), .B(n_27357), .Z(n_19205)
		);
	notech_reg regs_reg_8_11(.CP(n_62580), .D(n_19212), .CD(n_61599), .Q(regs_8
		[11]));
	notech_mux2 i_5489(.S(n_27365), .A(regs_8[11]), .B(n_18546), .Z(n_19212)
		);
	notech_reg regs_reg_8_12(.CP(n_62580), .D(n_19219), .CD(n_61599), .Q(regs_8
		[12]));
	notech_mux2 i_5497(.S(n_27365), .A(regs_8[12]), .B(n_27358), .Z(n_19219)
		);
	notech_reg regs_reg_8_13(.CP(n_62580), .D(n_19227), .CD(n_61599), .Q(regs_8
		[13]));
	notech_mux2 i_5505(.S(n_27365), .A(regs_8[13]), .B(n_18558), .Z(n_19227)
		);
	notech_nand3 i_56932263(.A(n_32393), .B(n_62794), .C(n_26818), .Z(n_2372
		));
	notech_reg regs_reg_8_14(.CP(n_62580), .D(n_19234), .CD(n_61599), .Q(regs_8
		[14]));
	notech_mux2 i_5513(.S(n_27365), .A(regs_8[14]), .B(n_18564), .Z(n_19234)
		);
	notech_reg regs_reg_8_15(.CP(n_62666), .D(n_19241), .CD(n_61599), .Q(regs_8
		[15]));
	notech_mux2 i_5521(.S(n_27365), .A(regs_8[15]), .B(n_27359), .Z(n_19241)
		);
	notech_and4 i_34032453(.A(n_32446), .B(n_27085), .C(n_1869), .D(n_2939),
		 .Z(n_2370));
	notech_reg regs_reg_8_16(.CP(n_62666), .D(n_19248), .CD(n_61599), .Q(regs_8
		[16]));
	notech_mux2 i_5529(.S(n_54803), .A(regs_8[16]), .B(n_27360), .Z(n_19248)
		);
	notech_reg regs_reg_8_17(.CP(n_62666), .D(n_19255), .CD(n_61599), .Q(regs_8
		[17]));
	notech_mux2 i_5537(.S(n_54803), .A(regs_8[17]), .B(n_27361), .Z(n_19255)
		);
	notech_and3 i_54032287(.A(n_32434), .B(n_2419), .C(n_1881), .Z(n_2368)
		);
	notech_reg regs_reg_8_18(.CP(n_62666), .D(n_19263), .CD(n_61598), .Q(regs_8
		[18]));
	notech_mux2 i_5545(.S(n_54803), .A(regs_8[18]), .B(n_27362), .Z(n_19263)
		);
	notech_reg regs_reg_8_19(.CP(n_62666), .D(n_19270), .CD(n_61598), .Q(regs_8
		[19]));
	notech_mux2 i_5553(.S(n_54803), .A(regs_8[19]), .B(n_27363), .Z(n_19270)
		);
	notech_ao4 i_52932298(.A(n_32405), .B(n_3848598), .C(n_319391630), .D(n_4668680
		), .Z(n_2366));
	notech_reg regs_reg_8_20(.CP(n_62666), .D(n_19277), .CD(n_61598), .Q(regs_8
		[20]));
	notech_mux2 i_5561(.S(n_54803), .A(regs_8[20]), .B(n_18600), .Z(n_19277)
		);
	notech_reg regs_reg_8_21(.CP(n_62666), .D(n_19284), .CD(n_61598), .Q(regs_8
		[21]));
	notech_mux2 i_5569(.S(n_54803), .A(regs_8[21]), .B(n_27364), .Z(n_19284)
		);
	notech_reg regs_reg_8_22(.CP(n_62666), .D(n_19291), .CD(n_61598), .Q(regs_8
		[22]));
	notech_mux2 i_5577(.S(n_54803), .A(regs_8[22]), .B(n_18612), .Z(n_19291)
		);
	notech_and2 i_27832502(.A(n_1862), .B(n_29656), .Z(n_2363));
	notech_reg regs_reg_8_23(.CP(n_62666), .D(n_19298), .CD(n_61598), .Q(regs_8
		[23]));
	notech_mux2 i_5585(.S(n_54803), .A(regs_8[23]), .B(n_18618), .Z(n_19298)
		);
	notech_ao4 i_28132500(.A(write_ack), .B(n_26761), .C(n_5219), .D(n_5018715
		), .Z(n_2362));
	notech_reg regs_reg_8_24(.CP(n_62666), .D(n_19304), .CD(n_61598), .Q(regs_8
		[24]));
	notech_mux2 i_5593(.S(n_54803), .A(regs_8[24]), .B(n_18624), .Z(n_19304)
		);
	notech_reg regs_reg_8_25(.CP(n_62666), .D(n_19310), .CD(n_61598), .Q(regs_8
		[25]));
	notech_mux2 i_5601(.S(n_54803), .A(regs_8[25]), .B(n_18630), .Z(n_19310)
		);
	notech_reg regs_reg_8_26(.CP(n_62666), .D(n_19317), .CD(n_61598), .Q(regs_8
		[26]));
	notech_mux2 i_5609(.S(n_54803), .A(regs_8[26]), .B(n_18636), .Z(n_19317)
		);
	notech_and4 i_36532435(.A(n_59124), .B(n_2518), .C(n_2523), .D(n_243191971
		), .Z(n_2359));
	notech_reg regs_reg_8_27(.CP(n_62666), .D(n_19323), .CD(n_61598), .Q(regs_8
		[27]));
	notech_mux2 i_5617(.S(n_54803), .A(regs_8[27]), .B(n_18642), .Z(n_19323)
		);
	notech_and4 i_36432436(.A(n_2685), .B(n_22024), .C(n_4758689), .D(n_23625
		), .Z(n_2358));
	notech_reg regs_reg_8_28(.CP(n_62666), .D(n_19329), .CD(n_61600), .Q(regs_8
		[28]));
	notech_mux2 i_5625(.S(n_54803), .A(regs_8[28]), .B(n_18648), .Z(n_19329)
		);
	notech_ao4 i_36332437(.A(n_319791626), .B(n_23755), .C(n_319991624), .D(read_ack
		), .Z(n_2357));
	notech_reg regs_reg_8_29(.CP(n_62666), .D(n_19335), .CD(n_61600), .Q(regs_8
		[29]));
	notech_mux2 i_5633(.S(n_54803), .A(regs_8[29]), .B(n_18654), .Z(n_19335)
		);
	notech_reg regs_reg_8_30(.CP(n_62666), .D(n_19341), .CD(n_61600), .Q(regs_8
		[30]));
	notech_mux2 i_5641(.S(n_54803), .A(regs_8[30]), .B(n_18660), .Z(n_19341)
		);
	notech_xor2 i_37232428(.A(cs[0]), .B(sav_cs[0]), .Z(n_2355));
	notech_reg regs_reg_8_31(.CP(n_62666), .D(n_19347), .CD(n_61600), .Q(regs_8
		[31]));
	notech_mux2 i_5649(.S(n_54803), .A(regs_8[31]), .B(n_18666), .Z(n_19347)
		);
	notech_nao3 i_9632643(.A(n_62798), .B(n_62836), .C(n_59451), .Z(n_2354)
		);
	notech_reg regs_reg_7_0(.CP(n_62666), .D(n_19353), .CD(n_61600), .Q(regs_7
		[0]));
	notech_mux2 i_5657(.S(\nbus_11350[0] ), .A(regs_7[0]), .B(n_27366), .Z(n_19353
		));
	notech_reg regs_reg_7_1(.CP(n_62580), .D(n_19359), .CD(n_61600), .Q(regs_7
		[1]));
	notech_mux2 i_5665(.S(\nbus_11350[0] ), .A(regs_7[1]), .B(n_21342), .Z(n_19359
		));
	notech_reg regs_reg_7_2(.CP(n_62580), .D(n_19365), .CD(n_61600), .Q(regs_7
		[2]));
	notech_mux2 i_5673(.S(\nbus_11350[0] ), .A(regs_7[2]), .B(n_27367), .Z(n_19365
		));
	notech_ao4 i_83232706(.A(n_62776), .B(n_60904), .C(n_60888), .D(n_17107)
		, .Z(n_2351));
	notech_reg regs_reg_7_3(.CP(n_62582), .D(n_19371), .CD(n_61600), .Q(regs_7
		[3]));
	notech_mux2 i_5681(.S(\nbus_11350[0] ), .A(regs_7[3]), .B(n_21354), .Z(n_19371
		));
	notech_or2 i_15232589(.A(n_19029), .B(n_19043), .Z(n_26580));
	notech_reg regs_reg_7_4(.CP(n_62582), .D(n_19377), .CD(n_61600), .Q(regs_7
		[4]));
	notech_mux2 i_5689(.S(\nbus_11350[0] ), .A(regs_7[4]), .B(n_21360), .Z(n_19377
		));
	notech_xor2 i_14232599(.A(cs[1]), .B(sav_cs[1]), .Z(n_2350));
	notech_reg regs_reg_7_5(.CP(n_62582), .D(n_19383), .CD(n_61600), .Q(regs_7
		[5]));
	notech_mux2 i_5697(.S(\nbus_11350[0] ), .A(regs_7[5]), .B(n_21366), .Z(n_19383
		));
	notech_nao3 i_12832613(.A(n_62868), .B(\opcode[3] ), .C(n_27925), .Z(n_24989
		));
	notech_reg regs_reg_7_6(.CP(n_62582), .D(n_19389), .CD(n_61599), .Q(regs_7
		[6]));
	notech_mux2 i_5705(.S(\nbus_11350[0] ), .A(regs_7[6]), .B(n_27368), .Z(n_19389
		));
	notech_nand2 i_11532626(.A(n_62868), .B(\opcode[3] ), .Z(n_25617));
	notech_reg regs_reg_7_7(.CP(n_62582), .D(n_19395), .CD(n_61599), .Q(regs_7
		[7]));
	notech_mux2 i_5713(.S(\nbus_11350[0] ), .A(regs_7[7]), .B(n_27300), .Z(n_19395
		));
	notech_nao3 i_3507(.A(n_27170), .B(n_27123), .C(n_32443), .Z(n_32378));
	notech_reg regs_reg_7_8(.CP(n_62582), .D(n_19403), .CD(n_61599), .Q(regs_7
		[8]));
	notech_mux2 i_5721(.S(\nbus_11350[0] ), .A(regs_7[8]), .B(n_21384), .Z(n_19403
		));
	notech_ao3 i_165232918(.A(n_56950), .B(n_60139), .C(n_56858), .Z(n_2349)
		);
	notech_reg regs_reg_7_9(.CP(n_62582), .D(n_19409), .CD(n_61599), .Q(regs_7
		[9]));
	notech_mux2 i_5729(.S(\nbus_11350[0] ), .A(regs_7[9]), .B(n_27369), .Z(n_19409
		));
	notech_reg regs_reg_7_10(.CP(n_62582), .D(n_19415), .CD(n_61599), .Q(regs_7
		[10]));
	notech_mux2 i_5737(.S(\nbus_11350[0] ), .A(regs_7[10]), .B(n_21396), .Z(n_19415
		));
	notech_or4 i_72232793(.A(n_58101), .B(n_56970), .C(n_56827), .D(n_61133)
		, .Z(n_32347));
	notech_reg regs_reg_7_11(.CP(n_62582), .D(n_19421), .CD(n_61600), .Q(regs_7
		[11]));
	notech_mux2 i_5745(.S(\nbus_11350[0] ), .A(regs_7[11]), .B(n_27370), .Z(n_19421
		));
	notech_or4 i_72132796(.A(n_58062), .B(n_2937), .C(n_56827), .D(n_61133),
		 .Z(n_32351));
	notech_reg regs_reg_7_12(.CP(n_62582), .D(n_19427), .CD(n_61600), .Q(regs_7
		[12]));
	notech_mux2 i_5753(.S(\nbus_11350[0] ), .A(regs_7[12]), .B(n_21408), .Z(n_19427
		));
	notech_nao3 i_72032800(.A(n_32386), .B(n_60139), .C(n_56829), .Z(n_32355
		));
	notech_reg regs_reg_7_13(.CP(n_62582), .D(n_19433), .CD(n_61600), .Q(regs_7
		[13]));
	notech_mux2 i_5761(.S(\nbus_11350[0] ), .A(regs_7[13]), .B(n_27371), .Z(n_19433
		));
	notech_or4 i_33232801(.A(n_32378), .B(n_60207), .C(n_60986), .D(n_56983)
		, .Z(n_32356));
	notech_reg regs_reg_7_14(.CP(n_62582), .D(n_19439), .CD(n_61600), .Q(regs_7
		[14]));
	notech_mux2 i_5769(.S(\nbus_11350[0] ), .A(regs_7[14]), .B(n_27372), .Z(n_19439
		));
	notech_nor2 i_162132921(.A(n_305391770), .B(n_61136), .Z(n_234791985));
	notech_reg regs_reg_7_15(.CP(n_62582), .D(n_19445), .CD(n_61595), .Q(regs_7
		[15]));
	notech_mux2 i_5777(.S(\nbus_11350[0] ), .A(regs_7[15]), .B(n_27373), .Z(n_19445
		));
	notech_reg regs_reg_7_16(.CP(n_62582), .D(n_19451), .CD(n_61595), .Q(regs_7
		[16]));
	notech_mux2 i_5785(.S(n_54823), .A(regs_7[16]), .B(n_27374), .Z(n_19451)
		);
	notech_or4 i_58455618(.A(n_61171), .B(n_61160), .C(n_61151), .D(n_26634)
		, .Z(n_27753));
	notech_reg regs_reg_7_17(.CP(n_62582), .D(n_19457), .CD(n_61595), .Q(regs_7
		[17]));
	notech_mux2 i_5793(.S(n_54823), .A(regs_7[17]), .B(n_21438), .Z(n_19457)
		);
	notech_nand3 i_194755555(.A(n_56983), .B(n_314291681), .C(n_27273), .Z(n_30822
		));
	notech_reg regs_reg_7_18(.CP(n_62582), .D(n_19463), .CD(n_61595), .Q(regs_7
		[18]));
	notech_mux2 i_5801(.S(n_54823), .A(regs_7[18]), .B(n_21444), .Z(n_19463)
		);
	notech_reg regs_reg_7_19(.CP(n_62582), .D(n_19469), .CD(n_61595), .Q(regs_7
		[19]));
	notech_mux2 i_5809(.S(n_54823), .A(regs_7[19]), .B(n_21450), .Z(n_19469)
		);
	notech_reg regs_reg_7_20(.CP(n_62582), .D(n_19475), .CD(n_61595), .Q(regs_7
		[20]));
	notech_mux2 i_5817(.S(n_54823), .A(regs_7[20]), .B(n_21456), .Z(n_19475)
		);
	notech_ao4 i_170736599(.A(n_57976), .B(n_28321), .C(n_60845), .D(n_28515
		), .Z(n_2343));
	notech_reg regs_reg_7_21(.CP(n_62582), .D(n_19481), .CD(n_61595), .Q(regs_7
		[21]));
	notech_mux2 i_5825(.S(n_54823), .A(regs_7[21]), .B(n_21462), .Z(n_19481)
		);
	notech_ao4 i_170836598(.A(n_58009), .B(n_27893), .C(n_56463), .D(n_29618
		), .Z(n_2342));
	notech_reg regs_reg_7_22(.CP(n_62526), .D(n_19487), .CD(n_61595), .Q(regs_7
		[22]));
	notech_mux2 i_5833(.S(n_54823), .A(regs_7[22]), .B(n_21468), .Z(n_19487)
		);
	notech_and2 i_171236594(.A(n_2340), .B(n_2339), .Z(n_2341));
	notech_reg regs_reg_7_23(.CP(n_62526), .D(n_19493), .CD(n_61595), .Q(regs_7
		[23]));
	notech_mux2 i_5841(.S(n_54823), .A(regs_7[23]), .B(n_21474), .Z(n_19493)
		);
	notech_ao4 i_171036596(.A(n_56400), .B(n_28189), .C(n_56385), .D(n_28418
		), .Z(n_2340));
	notech_reg regs_reg_7_24(.CP(n_62526), .D(n_19499), .CD(n_61595), .Q(regs_7
		[24]));
	notech_mux2 i_5849(.S(n_54823), .A(regs_7[24]), .B(n_21480), .Z(n_19499)
		);
	notech_ao4 i_171136595(.A(n_59344), .B(n_28559), .C(n_56371), .D(n_28354
		), .Z(n_2339));
	notech_reg regs_reg_7_25(.CP(n_62526), .D(n_19505), .CD(n_61594), .Q(regs_7
		[25]));
	notech_mux2 i_5857(.S(n_54823), .A(regs_7[25]), .B(n_21486), .Z(n_19505)
		);
	notech_and4 i_172036586(.A(n_2336), .B(n_2335), .C(n_2333), .D(n_2332), 
		.Z(n_2338));
	notech_reg regs_reg_7_26(.CP(n_62526), .D(n_19511), .CD(n_61594), .Q(regs_7
		[26]));
	notech_mux2 i_5865(.S(n_54823), .A(regs_7[26]), .B(n_1561), .Z(n_19511)
		);
	notech_reg regs_reg_7_27(.CP(n_62526), .D(n_19517), .CD(n_61594), .Q(regs_7
		[27]));
	notech_mux2 i_5873(.S(n_54823), .A(regs_7[27]), .B(n_21498), .Z(n_19517)
		);
	notech_ao4 i_171436592(.A(n_56452), .B(n_28288), .C(n_58024), .D(n_28482
		), .Z(n_2336));
	notech_reg regs_reg_7_28(.CP(n_62526), .D(n_19524), .CD(n_61594), .Q(regs_7
		[28]));
	notech_mux2 i_5881(.S(n_54823), .A(regs_7[28]), .B(n_218659267), .Z(n_19524
		));
	notech_ao4 i_171536591(.A(n_56447), .B(n_28256), .C(n_56432), .D(n_28221
		), .Z(n_2335));
	notech_reg regs_reg_7_29(.CP(n_62526), .D(n_19530), .CD(n_61594), .Q(regs_7
		[29]));
	notech_mux2 i_5890(.S(n_54823), .A(regs_7[29]), .B(n_217359254), .Z(n_19530
		));
	notech_reg regs_reg_7_30(.CP(n_62526), .D(n_19536), .CD(n_61595), .Q(regs_7
		[30]));
	notech_mux2 i_5898(.S(n_54823), .A(regs_7[30]), .B(n_21516), .Z(n_19536)
		);
	notech_ao4 i_171736589(.A(n_56908), .B(n_29617), .C(n_56427), .D(n_28386
		), .Z(n_2333));
	notech_reg regs_reg_7_31(.CP(n_62526), .D(n_19542), .CD(n_61595), .Q(regs_7
		[31]));
	notech_mux2 i_5906(.S(n_54823), .A(regs_7[31]), .B(n_27375), .Z(n_19542)
		);
	notech_ao4 i_171836588(.A(n_56414), .B(n_28450), .C(n_56405), .D(n_28592
		), .Z(n_2332));
	notech_reg pipe_mul_reg_0(.CP(n_62576), .D(n_19548), .CD(n_61594), .Q(pipe_mul
		[0]));
	notech_mux2 i_5914(.S(\nbus_11306[0] ), .A(pipe_mul[0]), .B(n_194086214)
		, .Z(n_19548));
	notech_reg pipe_mul_reg_1(.CP(n_62566), .D(n_19554), .CD(n_61595), .Q(pipe_mul
		[1]));
	notech_mux2 i_5922(.S(\nbus_11306[0] ), .A(pipe_mul[1]), .B(n_194186215)
		, .Z(n_19554));
	notech_reg CFOF_mul_reg(.CP(n_62566), .D(n_19560), .CD(n_61597), .Q(CFOF_mul
		));
	notech_mux2 i_5931(.S(n_114468161), .A(n_12393), .B(CFOF_mul), .Z(n_19560
		));
	notech_ao4 i_172136585(.A(n_57976), .B(n_28319), .C(n_60845), .D(n_28513
		), .Z(n_2329));
	notech_reg eval_flag_reg(.CP(n_62566), .D(n_19566), .CD(n_61597), .Q(eval_flag
		));
	notech_mux2 i_5941(.S(n_15683), .A(eval_flag), .B(n_328690784), .Z(n_19566
		));
	notech_ao4 i_172236584(.A(n_58009), .B(n_27891), .C(n_56463), .D(n_29613
		), .Z(n_2328));
	notech_reg rep_en1_reg(.CP(n_62566), .D(n_19572), .CD(n_61597), .Q(rep_en1
		));
	notech_mux2 i_5950(.S(n_14570), .A(rep_en1), .B(n_60316), .Z(n_19572));
	notech_and2 i_172636580(.A(n_2326), .B(n_2325), .Z(n_2327));
	notech_reg rep_en2_reg(.CP(n_62566), .D(n_19578), .CD(n_61597), .Q(rep_en2
		));
	notech_mux2 i_5958(.S(n_14425), .A(rep_en2), .B(n_60316), .Z(n_19578));
	notech_ao4 i_172436582(.A(n_56400), .B(n_28187), .C(n_28416), .D(n_56385
		), .Z(n_2326));
	notech_reg rep_en3_reg(.CP(n_62566), .D(n_19584), .CD(n_61597), .Q(rep_en3
		));
	notech_mux2 i_5967(.S(n_16532), .A(rep_en3), .B(n_60321), .Z(n_19584));
	notech_ao4 i_172536581(.A(n_59344), .B(n_28557), .C(n_56371), .D(n_28352
		), .Z(n_2325));
	notech_reg rep_en4_reg(.CP(n_62566), .D(n_19590), .CD(n_61598), .Q(rep_en4
		));
	notech_mux2 i_5976(.S(n_20021), .A(rep_en4), .B(n_60321), .Z(n_19590));
	notech_and4 i_173436572(.A(n_2322), .B(n_232191987), .C(n_2319), .D(n_2318
		), .Z(n_2324));
	notech_reg rep_en5_reg(.CP(n_62566), .D(n_19596), .CD(n_61598), .Q(rep_en5
		));
	notech_mux2 i_5984(.S(n_15633), .A(rep_en5), .B(n_60318), .Z(n_19596));
	notech_reg nCF_reg(.CP(n_62566), .D(n_19602), .CD(n_61598), .Q(nCF));
	notech_mux2 i_5993(.S(n_12057), .A(nCF), .B(n_27022), .Z(n_19602));
	notech_ao4 i_172836578(.A(n_56452), .B(n_28286), .C(n_58024), .D(n_28480
		), .Z(n_2322));
	notech_reg nPF_reg(.CP(n_62566), .D(n_19608), .CD(n_61598), .Q(nPF));
	notech_mux2 i_6003(.S(n_15649), .A(nPF), .B(n_309787371), .Z(n_19608));
	notech_ao4 i_172936577(.A(n_56447), .B(n_28254), .C(n_56432), .D(n_28219
		), .Z(n_232191987));
	notech_reg nAF_reg(.CP(n_62566), .D(n_19614), .CD(n_61597), .Q(nAF));
	notech_mux2 i_6011(.S(n_328484275), .A(nAF_arithbox), .B(nAF), .Z(n_19614
		));
	notech_reg nSF_reg(.CP(n_62566), .D(n_19620), .CD(n_61597), .Q(nSF));
	notech_mux2 i_6019(.S(n_58219), .A(n_26608), .B(nSF), .Z(n_19620));
	notech_ao4 i_173136575(.A(n_56908), .B(n_29612), .C(n_56427), .D(n_28384
		), .Z(n_2319));
	notech_reg opas_reg(.CP(n_62642), .D(n_19629), .CD(n_61597), .Q(opas));
	notech_mux2 i_6027(.S(n_328484275), .A(opas_arithbox), .B(opas), .Z(n_19629
		));
	notech_ao4 i_173236574(.A(n_56414), .B(n_28448), .C(n_56405), .D(n_28590
		), .Z(n_2318));
	notech_reg opbs_reg(.CP(n_62642), .D(n_19635), .CD(n_61595), .Q(opbs));
	notech_mux2 i_6035(.S(n_328484275), .A(opbs_arithbox), .B(opbs), .Z(n_19635
		));
	notech_reg nOF_reg(.CP(n_62642), .D(n_19641), .CD(n_61597), .Q(nOF));
	notech_mux2 i_6043(.S(n_27386), .A(nOF), .B(n_27384), .Z(n_19641));
	notech_reg regs_reg_15_0(.CP(n_62642), .D(n_19648), .CD(n_61597), .Q(\eflags[0] 
		));
	notech_mux2 i_6051(.S(\nbus_11376[0] ), .A(\eflags[0] ), .B(n_27387), .Z
		(n_19648));
	notech_ao4 i_173536571(.A(n_57976), .B(n_28318), .C(n_60845), .D(n_28512
		), .Z(n_231591988));
	notech_reg regs_reg_15_1(.CP(n_62642), .D(n_19655), .CD(n_61597), .Q(\eflags[1] 
		));
	notech_mux2 i_6059(.S(n_3907), .A(n_25252), .B(\eflags[1] ), .Z(n_19655)
		);
	notech_ao4 i_173636570(.A(n_58009), .B(n_27890), .C(n_56468), .D(n_29611
		), .Z(n_2314));
	notech_reg regs_reg_15_2(.CP(n_62642), .D(n_19662), .CD(n_61597), .Q(\eflags[2] 
		));
	notech_mux2 i_6067(.S(\nbus_11376[2] ), .A(\eflags[2] ), .B(n_3895), .Z(n_19662
		));
	notech_and2 i_174036566(.A(n_2312), .B(n_2311), .Z(n_2313));
	notech_reg regs_reg_15_3(.CP(n_62642), .D(n_19669), .CD(n_61597), .Q(\eflags[3] 
		));
	notech_mux2 i_6075(.S(n_3907), .A(n_25264), .B(\eflags[3] ), .Z(n_19669)
		);
	notech_ao4 i_173836568(.A(n_56400), .B(n_28186), .C(n_56385), .D(n_28415
		), .Z(n_2312));
	notech_reg regs_reg_15_4(.CP(n_62642), .D(n_19676), .CD(n_61597), .Q(\eflags[4] 
		));
	notech_mux2 i_6083(.S(\nbus_11376[0] ), .A(\eflags[4] ), .B(n_25270), .Z
		(n_19676));
	notech_ao4 i_173936567(.A(n_59349), .B(n_28556), .C(n_56371), .D(n_28351
		), .Z(n_2311));
	notech_reg regs_reg_15_5(.CP(n_62642), .D(n_19682), .CD(n_61575), .Q(\eflags[5] 
		));
	notech_mux2 i_6091(.S(n_3907), .A(n_25276), .B(\eflags[5] ), .Z(n_19682)
		);
	notech_and4 i_174836558(.A(n_2308), .B(n_2307), .C(n_2305), .D(n_2304), 
		.Z(n_2310));
	notech_reg regs_reg_15_6(.CP(n_62642), .D(n_19688), .CD(n_61576), .Q(\eflags[6] 
		));
	notech_mux2 i_6099(.S(n_27393), .A(\eflags[6] ), .B(n_3869), .Z(n_19688)
		);
	notech_reg regs_reg_15_7(.CP(n_62642), .D(n_19694), .CD(n_61575), .Q(\eflags[7] 
		));
	notech_mux2 i_6107(.S(n_27393), .A(\eflags[7] ), .B(n_25288), .Z(n_19694
		));
	notech_ao4 i_174236564(.A(n_56452), .B(n_28285), .C(n_58024), .D(n_28479
		), .Z(n_2308));
	notech_reg regs_reg_15_8(.CP(n_62642), .D(n_19700), .CD(n_61575), .Q(\eflags[8] 
		));
	notech_mux2 i_6115(.S(\nbus_11376[8] ), .A(\eflags[8] ), .B(n_27388), .Z
		(n_19700));
	notech_ao4 i_174336563(.A(n_56447), .B(n_28253), .C(n_56432), .D(n_28218
		), .Z(n_2307));
	notech_reg regs_reg_15_9(.CP(n_62642), .D(n_19706), .CD(n_61576), .Q(ie)
		);
	notech_mux2 i_6123(.S(n_27390), .A(ie), .B(n_27389), .Z(n_19706));
	notech_reg regs_reg_15_10(.CP(n_62642), .D(n_19712), .CD(n_61576), .Q(\eflags[10] 
		));
	notech_mux2 i_6131(.S(n_27392), .A(n_56172), .B(n_27391), .Z(n_19712));
	notech_ao4 i_174536561(.A(n_56908), .B(n_29610), .C(n_56427), .D(n_28383
		), .Z(n_2305));
	notech_reg regs_reg_15_11(.CP(n_62642), .D(n_19718), .CD(n_61576), .Q(\eflags[11] 
		));
	notech_mux2 i_6139(.S(n_27393), .A(\eflags[11] ), .B(n_1598), .Z(n_19718
		));
	notech_ao4 i_174636560(.A(n_56414), .B(n_28447), .C(n_56405), .D(n_28589
		), .Z(n_2304));
	notech_reg regs_reg_15_12(.CP(n_62642), .D(n_19724), .CD(n_61576), .Q(\eflags[12] 
		));
	notech_mux2 i_6147(.S(\nbus_11376[12] ), .A(\eflags[12] ), .B(n_27394), 
		.Z(n_19724));
	notech_reg regs_reg_15_13(.CP(n_62642), .D(n_19730), .CD(n_61576), .Q(\eflags[13] 
		));
	notech_mux2 i_6155(.S(\nbus_11376[12] ), .A(\eflags[13] ), .B(n_27395), 
		.Z(n_19730));
	notech_reg regs_reg_15_14(.CP(n_62642), .D(n_19736), .CD(n_61575), .Q(\eflags[14] 
		));
	notech_mux2 i_6163(.S(\nbus_11376[12] ), .A(\eflags[14] ), .B(n_27396), 
		.Z(n_19736));
	notech_ao4 i_174936557(.A(n_57976), .B(n_28316), .C(n_60845), .D(n_28510
		), .Z(n_2301));
	notech_reg regs_reg_15_15(.CP(n_62642), .D(n_19742), .CD(n_61575), .Q(\eflags[15] 
		));
	notech_mux2 i_6171(.S(n_3907), .A(n_27397), .B(\eflags[15] ), .Z(n_19742
		));
	notech_ao4 i_175036556(.A(n_58009), .B(n_27888), .C(n_56463), .D(n_29607
		), .Z(n_2300));
	notech_reg regs_reg_15_16(.CP(n_62640), .D(n_19748), .CD(n_61575), .Q(\eflags[16] 
		));
	notech_mux2 i_6179(.S(\nbus_11376[12] ), .A(\eflags[16] ), .B(n_25342), 
		.Z(n_19748));
	notech_and2 i_175436552(.A(n_2298), .B(n_2297), .Z(n_2299));
	notech_reg regs_reg_15_17(.CP(n_62640), .D(n_19754), .CD(n_61575), .Q(\eflags[17] 
		));
	notech_mux2 i_6187(.S(\nbus_11376[12] ), .A(\eflags[17] ), .B(n_27398), 
		.Z(n_19754));
	notech_ao4 i_175236554(.A(n_56400), .B(n_28184), .C(n_28413), .D(n_56385
		), .Z(n_2298));
	notech_reg regs_reg_15_18(.CP(n_62716), .D(n_19760), .CD(n_61575), .Q(\eflags[18] 
		));
	notech_mux2 i_6195(.S(\nbus_11376[12] ), .A(\eflags[18] ), .B(n_27399), 
		.Z(n_19760));
	notech_ao4 i_175336553(.A(n_59344), .B(n_28554), .C(n_56371), .D(n_28349
		), .Z(n_2297));
	notech_reg regs_reg_15_19(.CP(n_62716), .D(n_19766), .CD(n_61575), .Q(\eflags[19] 
		));
	notech_mux2 i_6203(.S(\nbus_11376[12] ), .A(\eflags[19] ), .B(n_27400), 
		.Z(n_19766));
	notech_and4 i_176236544(.A(n_2294), .B(n_2293), .C(n_2291), .D(n_2290), 
		.Z(n_2296));
	notech_reg regs_reg_15_20(.CP(n_62716), .D(n_19772), .CD(n_61575), .Q(\eflags[20] 
		));
	notech_mux2 i_6211(.S(\nbus_11376[12] ), .A(\eflags[20] ), .B(n_25366), 
		.Z(n_19772));
	notech_reg regs_reg_15_21(.CP(n_62716), .D(n_19778), .CD(n_61575), .Q(\eflags[21] 
		));
	notech_mux2 i_6219(.S(\nbus_11376[12] ), .A(\eflags[21] ), .B(n_27401), 
		.Z(n_19778));
	notech_ao4 i_175636550(.A(n_56452), .B(n_28283), .C(n_58024), .D(n_28477
		), .Z(n_2294));
	notech_reg regs_reg_15_22(.CP(n_62716), .D(n_19784), .CD(n_61575), .Q(\eflags[22] 
		));
	notech_mux2 i_6227(.S(\nbus_11376[12] ), .A(\eflags[22] ), .B(n_25378), 
		.Z(n_19784));
	notech_ao4 i_175736549(.A(n_56447), .B(n_28251), .C(n_56432), .D(n_28216
		), .Z(n_2293));
	notech_reg regs_reg_15_23(.CP(n_62716), .D(n_19790), .CD(n_61575), .Q(\eflags[23] 
		));
	notech_mux2 i_6235(.S(\nbus_11376[12] ), .A(\eflags[23] ), .B(n_25384), 
		.Z(n_19790));
	notech_reg regs_reg_15_24(.CP(n_62716), .D(n_19796), .CD(n_61577), .Q(\eflags[24] 
		));
	notech_mux2 i_6243(.S(\nbus_11376[12] ), .A(\eflags[24] ), .B(n_25390), 
		.Z(n_19796));
	notech_ao4 i_175936547(.A(n_56908), .B(n_29606), .C(n_56427), .D(n_28381
		), .Z(n_2291));
	notech_reg regs_reg_15_25(.CP(n_62716), .D(n_19802), .CD(n_61577), .Q(\eflags[25] 
		));
	notech_mux2 i_6251(.S(\nbus_11376[12] ), .A(\eflags[25] ), .B(n_25396), 
		.Z(n_19802));
	notech_ao4 i_176036546(.A(n_56414), .B(n_28445), .C(n_56405), .D(n_28587
		), .Z(n_2290));
	notech_reg regs_reg_15_26(.CP(n_62716), .D(n_19809), .CD(n_61577), .Q(\eflags[26] 
		));
	notech_mux2 i_6259(.S(\nbus_11376[12] ), .A(\eflags[26] ), .B(n_25402), 
		.Z(n_19809));
	notech_reg regs_reg_15_27(.CP(n_62716), .D(n_19815), .CD(n_61577), .Q(\eflags[27] 
		));
	notech_mux2 i_6267(.S(\nbus_11376[12] ), .A(\eflags[27] ), .B(n_25408), 
		.Z(n_19815));
	notech_reg regs_reg_15_28(.CP(n_62716), .D(n_19821), .CD(n_61577), .Q(\eflags[28] 
		));
	notech_mux2 i_6275(.S(\nbus_11376[12] ), .A(\eflags[28] ), .B(n_25414), 
		.Z(n_19821));
	notech_ao4 i_193336375(.A(n_57976), .B(n_28301), .C(n_60845), .D(n_28494
		), .Z(n_2287));
	notech_reg regs_reg_15_29(.CP(n_62716), .D(n_19827), .CD(n_61577), .Q(\eflags[29] 
		));
	notech_mux2 i_6283(.S(\nbus_11376[12] ), .A(\eflags[29] ), .B(n_1577), .Z
		(n_19827));
	notech_ao4 i_193436374(.A(n_58009), .B(n_27869), .C(n_56463), .D(n_29620
		), .Z(n_2286));
	notech_reg regs_reg_15_30(.CP(n_62716), .D(n_19833), .CD(n_61577), .Q(\eflags[30] 
		));
	notech_mux2 i_6291(.S(\nbus_11376[12] ), .A(\eflags[30] ), .B(n_25426), 
		.Z(n_19833));
	notech_and2 i_193836370(.A(n_2284), .B(n_2283), .Z(n_2285));
	notech_reg regs_reg_15_31(.CP(n_62716), .D(n_19839), .CD(n_61577), .Q(\eflags[31] 
		));
	notech_mux2 i_6299(.S(\nbus_11376[12] ), .A(\eflags[31] ), .B(n_27402), 
		.Z(n_19839));
	notech_ao4 i_193636372(.A(n_56396), .B(n_28169), .C(n_56385), .D(n_28398
		), .Z(n_2284));
	notech_reg regs_reg_6_0(.CP(n_62716), .D(n_19845), .CD(n_61577), .Q(regs_6
		[0]));
	notech_mux2 i_6307(.S(n_3815), .A(n_27403), .B(regs_6[0]), .Z(n_19845)
		);
	notech_ao4 i_193736371(.A(n_59344), .B(n_28529), .C(n_56371), .D(n_28334
		), .Z(n_2283));
	notech_reg regs_reg_6_1(.CP(n_62716), .D(n_19851), .CD(n_61577), .Q(regs_6
		[1]));
	notech_mux2 i_6315(.S(n_3815), .A(n_18138), .B(regs_6[1]), .Z(n_19851)
		);
	notech_and4 i_194636362(.A(n_2280), .B(n_2279), .C(n_2277), .D(n_2276), 
		.Z(n_2282));
	notech_reg regs_reg_6_2(.CP(n_62716), .D(n_19857), .CD(n_61576), .Q(regs_6
		[2]));
	notech_mux2 i_6323(.S(n_3815), .A(n_27404), .B(regs_6[2]), .Z(n_19857)
		);
	notech_reg regs_reg_6_3(.CP(n_62716), .D(n_19863), .CD(n_61576), .Q(regs_6
		[3]));
	notech_mux2 i_6331(.S(n_3815), .A(n_18150), .B(regs_6[3]), .Z(n_19863)
		);
	notech_ao4 i_194036368(.A(n_56452), .B(n_28268), .C(n_58024), .D(n_28462
		), .Z(n_2280));
	notech_reg regs_reg_6_4(.CP(n_62640), .D(n_19869), .CD(n_61576), .Q(regs_6
		[4]));
	notech_mux2 i_6339(.S(n_3815), .A(n_18156), .B(regs_6[4]), .Z(n_19869)
		);
	notech_ao4 i_194136367(.A(n_56443), .B(n_28235), .C(n_56432), .D(n_28201
		), .Z(n_2279));
	notech_reg regs_reg_6_5(.CP(n_62640), .D(n_19875), .CD(n_61576), .Q(regs_6
		[5]));
	notech_mux2 i_6347(.S(n_3815), .A(n_18162), .B(regs_6[5]), .Z(n_19875)
		);
	notech_reg regs_reg_6_6(.CP(n_62640), .D(n_19881), .CD(n_61576), .Q(regs_6
		[6]));
	notech_mux2 i_6355(.S(n_3815), .A(n_18168), .B(regs_6[6]), .Z(n_19881)
		);
	notech_ao4 i_194336365(.A(n_56908), .B(n_29621), .C(n_56423), .D(n_28366
		), .Z(n_2277));
	notech_reg regs_reg_6_7(.CP(n_62640), .D(n_19887), .CD(n_61577), .Q(regs_6
		[7]));
	notech_mux2 i_6363(.S(n_3815), .A(n_27405), .B(regs_6[7]), .Z(n_19887)
		);
	notech_ao4 i_194436364(.A(n_56414), .B(n_28430), .C(n_56405), .D(n_28572
		), .Z(n_2276));
	notech_reg regs_reg_6_8(.CP(n_62640), .D(n_19893), .CD(n_61577), .Q(regs_6
		[8]));
	notech_mux2 i_6371(.S(n_3815), .A(n_18180), .B(regs_6[8]), .Z(n_19893)
		);
	notech_reg regs_reg_6_9(.CP(n_62640), .D(n_19900), .CD(n_61576), .Q(regs_6
		[9]));
	notech_mux2 i_6379(.S(n_3815), .A(n_18186), .B(regs_6[9]), .Z(n_19900)
		);
	notech_reg regs_reg_6_10(.CP(n_62640), .D(n_19906), .CD(n_61576), .Q(regs_6
		[10]));
	notech_mux2 i_6387(.S(n_3815), .A(n_18192), .B(regs_6[10]), .Z(n_19906)
		);
	notech_ao4 i_198936319(.A(n_57976), .B(n_28296), .C(n_60845), .D(n_28490
		), .Z(n_2273));
	notech_reg regs_reg_6_11(.CP(n_62640), .D(n_19912), .CD(n_61572), .Q(regs_6
		[11]));
	notech_mux2 i_6395(.S(n_3815), .A(n_27298), .B(regs_6[11]), .Z(n_19912)
		);
	notech_ao4 i_199036318(.A(n_58009), .B(n_27865), .C(n_56463), .D(n_29615
		), .Z(n_2272));
	notech_reg regs_reg_6_12(.CP(n_62640), .D(n_19918), .CD(n_61572), .Q(regs_6
		[12]));
	notech_mux2 i_6403(.S(n_3815), .A(n_18204), .B(regs_6[12]), .Z(n_19918)
		);
	notech_and2 i_199436314(.A(n_2270), .B(n_2269), .Z(n_2271));
	notech_reg regs_reg_6_13(.CP(n_62640), .D(n_19924), .CD(n_61571), .Q(regs_6
		[13]));
	notech_mux2 i_6411(.S(n_3815), .A(n_27406), .B(regs_6[13]), .Z(n_19924)
		);
	notech_ao4 i_199236316(.A(n_56396), .B(n_28165), .C(n_56385), .D(n_28394
		), .Z(n_2270));
	notech_reg regs_reg_6_14(.CP(n_62716), .D(n_19932), .CD(n_61571), .Q(regs_6
		[14]));
	notech_mux2 i_6419(.S(n_3815), .A(n_27407), .B(regs_6[14]), .Z(n_19932)
		);
	notech_ao4 i_199336315(.A(n_59344), .B(n_28523), .C(n_56371), .D(n_28329
		), .Z(n_2269));
	notech_reg regs_reg_6_15(.CP(n_62638), .D(n_19938), .CD(n_61572), .Q(regs_6
		[15]));
	notech_mux2 i_6427(.S(n_3815), .A(n_18222), .B(regs_6[15]), .Z(n_19938)
		);
	notech_and4 i_200236306(.A(n_2266), .B(n_2265), .C(n_2263), .D(n_2262), 
		.Z(n_2268));
	notech_reg regs_reg_6_16(.CP(n_62638), .D(n_19944), .CD(n_61572), .Q(regs_6
		[16]));
	notech_mux2 i_6435(.S(n_54843), .A(n_18228), .B(regs_6[16]), .Z(n_19944)
		);
	notech_reg regs_reg_6_17(.CP(n_62712), .D(n_19950), .CD(n_61572), .Q(regs_6
		[17]));
	notech_mux2 i_6443(.S(n_54843), .A(n_18234), .B(regs_6[17]), .Z(n_19950)
		);
	notech_ao4 i_199636312(.A(n_56452), .B(n_28264), .C(n_58024), .D(n_28458
		), .Z(n_2266));
	notech_reg regs_reg_6_18(.CP(n_62712), .D(n_19956), .CD(n_61572), .Q(regs_6
		[18]));
	notech_mux2 i_6451(.S(n_54843), .A(n_18240), .B(regs_6[18]), .Z(n_19956)
		);
	notech_ao4 i_199736311(.A(n_56443), .B(n_28230), .C(n_56432), .D(n_28197
		), .Z(n_2265));
	notech_reg regs_reg_6_19(.CP(n_62712), .D(n_19962), .CD(n_61572), .Q(regs_6
		[19]));
	notech_mux2 i_6459(.S(n_54843), .A(n_18246), .B(regs_6[19]), .Z(n_19962)
		);
	notech_reg regs_reg_6_20(.CP(n_62712), .D(n_19970), .CD(n_61571), .Q(regs_6
		[20]));
	notech_mux2 i_6467(.S(n_54843), .A(n_18252), .B(regs_6[20]), .Z(n_19970)
		);
	notech_ao4 i_199936309(.A(n_56908), .B(n_29616), .C(n_56423), .D(n_28362
		), .Z(n_2263));
	notech_reg regs_reg_6_21(.CP(n_62712), .D(n_19976), .CD(n_61571), .Q(regs_6
		[21]));
	notech_mux2 i_6475(.S(n_54843), .A(n_18258), .B(regs_6[21]), .Z(n_19976)
		);
	notech_ao4 i_200036308(.A(n_56414), .B(n_28426), .C(n_56405), .D(n_28567
		), .Z(n_2262));
	notech_reg regs_reg_6_22(.CP(n_62712), .D(n_19982), .CD(n_61571), .Q(regs_6
		[22]));
	notech_mux2 i_6483(.S(n_54843), .A(n_18264), .B(regs_6[22]), .Z(n_19982)
		);
	notech_reg regs_reg_6_23(.CP(n_62712), .D(n_19989), .CD(n_61571), .Q(regs_6
		[23]));
	notech_mux2 i_6491(.S(n_54843), .A(n_18270), .B(regs_6[23]), .Z(n_19989)
		);
	notech_reg regs_reg_6_24(.CP(n_62712), .D(n_19995), .CD(n_61571), .Q(regs_6
		[24]));
	notech_mux2 i_6499(.S(n_54843), .A(n_18276), .B(regs_6[24]), .Z(n_19995)
		);
	notech_ao4 i_208736221(.A(n_57976), .B(n_28320), .C(n_60845), .D(n_28514
		), .Z(n_2259));
	notech_reg regs_reg_6_25(.CP(n_62712), .D(n_20001), .CD(n_61571), .Q(regs_6
		[25]));
	notech_mux2 i_6507(.S(n_54843), .A(n_18282), .B(regs_6[25]), .Z(n_20001)
		);
	notech_ao4 i_208836220(.A(n_58009), .B(n_27892), .C(n_56463), .D(n_29625
		), .Z(n_2258));
	notech_reg regs_reg_6_26(.CP(n_62712), .D(n_20007), .CD(n_61571), .Q(regs_6
		[26]));
	notech_mux2 i_6515(.S(n_54843), .A(n_1623), .B(regs_6[26]), .Z(n_20007)
		);
	notech_and2 i_209236216(.A(n_2256), .B(n_2255), .Z(n_2257));
	notech_reg regs_reg_6_27(.CP(n_62754), .D(n_20013), .CD(n_61571), .Q(regs_6
		[27]));
	notech_mux2 i_6523(.S(n_54843), .A(n_1611), .B(regs_6[27]), .Z(n_20013)
		);
	notech_ao4 i_209036218(.A(n_56396), .B(n_28188), .C(n_56385), .D(n_28417
		), .Z(n_2256));
	notech_reg regs_reg_6_28(.CP(n_62754), .D(n_20019), .CD(n_61571), .Q(regs_6
		[28]));
	notech_mux2 i_6531(.S(n_54843), .A(n_227859359), .B(regs_6[28]), .Z(n_20019
		));
	notech_ao4 i_209136217(.A(n_59344), .B(n_28558), .C(n_56371), .D(n_28353
		), .Z(n_2255));
	notech_reg regs_reg_6_29(.CP(n_62754), .D(n_20026), .CD(n_61571), .Q(regs_6
		[29]));
	notech_mux2 i_6539(.S(n_54843), .A(n_226659347), .B(regs_6[29]), .Z(n_20026
		));
	notech_and4 i_210036208(.A(n_2252), .B(n_2251), .C(n_2249), .D(n_2248), 
		.Z(n_2254));
	notech_reg regs_reg_6_30(.CP(n_62754), .D(n_20032), .CD(n_61573), .Q(regs_6
		[30]));
	notech_mux2 i_6547(.S(n_54843), .A(n_301391810), .B(regs_6[30]), .Z(n_20032
		));
	notech_reg regs_reg_6_31(.CP(n_62754), .D(n_20038), .CD(n_61573), .Q(regs_6
		[31]));
	notech_mux2 i_6555(.S(n_54843), .A(n_27408), .B(regs_6[31]), .Z(n_20038)
		);
	notech_ao4 i_209436214(.A(n_56452), .B(n_28287), .C(n_58024), .D(n_28481
		), .Z(n_2252));
	notech_reg regs_reg_5_0(.CP(n_62754), .D(n_20044), .CD(n_61573), .Q(regs_5
		[0]));
	notech_mux2 i_6563(.S(\nbus_11332[0] ), .A(regs_5[0]), .B(n_27409), .Z(n_20044
		));
	notech_ao4 i_209536213(.A(n_56443), .B(n_28255), .C(n_56432), .D(n_28220
		), .Z(n_2251));
	notech_reg regs_reg_5_1(.CP(n_62754), .D(n_20050), .CD(n_61573), .Q(regs_5
		[1]));
	notech_mux2 i_6571(.S(\nbus_11332[0] ), .A(regs_5[1]), .B(n_17786), .Z(n_20050
		));
	notech_reg regs_reg_5_2(.CP(n_62754), .D(n_20056), .CD(n_61573), .Q(regs_5
		[2]));
	notech_mux2 i_6579(.S(\nbus_11332[0] ), .A(regs_5[2]), .B(n_27410), .Z(n_20056
		));
	notech_ao4 i_209736211(.A(n_56908), .B(n_29624), .C(n_56423), .D(n_28385
		), .Z(n_2249));
	notech_reg regs_reg_5_3(.CP(n_62754), .D(n_20062), .CD(n_61573), .Q(regs_5
		[3]));
	notech_mux2 i_6587(.S(\nbus_11332[0] ), .A(regs_5[3]), .B(n_17798), .Z(n_20062
		));
	notech_ao4 i_209836210(.A(n_56414), .B(n_28449), .C(n_56405), .D(n_28591
		), .Z(n_2248));
	notech_reg regs_reg_5_4(.CP(n_62754), .D(n_20068), .CD(n_61573), .Q(regs_5
		[4]));
	notech_mux2 i_6595(.S(\nbus_11332[0] ), .A(regs_5[4]), .B(n_17804), .Z(n_20068
		));
	notech_reg regs_reg_5_5(.CP(n_62754), .D(n_20074), .CD(n_61573), .Q(regs_5
		[5]));
	notech_mux2 i_6603(.S(\nbus_11332[0] ), .A(regs_5[5]), .B(n_17810), .Z(n_20074
		));
	notech_reg regs_reg_5_6(.CP(n_62754), .D(n_20080), .CD(n_61573), .Q(regs_5
		[6]));
	notech_mux2 i_6611(.S(\nbus_11332[0] ), .A(regs_5[6]), .B(n_17816), .Z(n_20080
		));
	notech_ao4 i_210136207(.A(n_57976), .B(n_28317), .C(n_60845), .D(n_28511
		), .Z(n_2245));
	notech_reg regs_reg_5_7(.CP(n_62754), .D(n_20086), .CD(n_61573), .Q(regs_5
		[7]));
	notech_mux2 i_6619(.S(\nbus_11332[0] ), .A(regs_5[7]), .B(n_17822), .Z(n_20086
		));
	notech_ao4 i_210236206(.A(n_58009), .B(n_27889), .C(n_56463), .D(n_29609
		), .Z(n_2244));
	notech_reg regs_reg_5_8(.CP(n_62754), .D(n_20092), .CD(n_61572), .Q(regs_5
		[8]));
	notech_mux2 i_6627(.S(\nbus_11332[0] ), .A(regs_5[8]), .B(n_27411), .Z(n_20092
		));
	notech_and2 i_210636202(.A(n_2242), .B(n_2241), .Z(n_2243));
	notech_reg regs_reg_5_9(.CP(n_62754), .D(n_20099), .CD(n_61572), .Q(regs_5
		[9]));
	notech_mux2 i_6635(.S(\nbus_11332[0] ), .A(regs_5[9]), .B(n_27412), .Z(n_20099
		));
	notech_ao4 i_210436204(.A(n_56400), .B(n_28185), .C(n_28414), .D(n_56385
		), .Z(n_2242));
	notech_reg regs_reg_5_10(.CP(n_62754), .D(n_20107), .CD(n_61572), .Q(regs_5
		[10]));
	notech_mux2 i_6643(.S(\nbus_11332[0] ), .A(regs_5[10]), .B(n_27413), .Z(n_20107
		));
	notech_ao4 i_210536203(.A(n_59344), .B(n_28555), .C(n_56371), .D(n_28350
		), .Z(n_2241));
	notech_reg regs_reg_5_11(.CP(n_62754), .D(n_20114), .CD(n_61572), .Q(regs_5
		[11]));
	notech_mux2 i_6651(.S(\nbus_11332[0] ), .A(regs_5[11]), .B(n_17846), .Z(n_20114
		));
	notech_and4 i_211436194(.A(n_2238), .B(n_2237), .C(n_2235), .D(n_2234), 
		.Z(n_2240));
	notech_reg regs_reg_5_12(.CP(n_62754), .D(n_20122), .CD(n_61572), .Q(regs_5
		[12]));
	notech_mux2 i_6659(.S(\nbus_11332[0] ), .A(regs_5[12]), .B(n_27414), .Z(n_20122
		));
	notech_reg regs_reg_5_13(.CP(n_62712), .D(n_20129), .CD(n_61573), .Q(regs_5
		[13]));
	notech_mux2 i_6667(.S(\nbus_11332[0] ), .A(regs_5[13]), .B(n_17858), .Z(n_20129
		));
	notech_ao4 i_210836200(.A(n_56452), .B(n_28284), .C(n_58024), .D(n_28478
		), .Z(n_2238));
	notech_reg regs_reg_5_14(.CP(n_62754), .D(n_20137), .CD(n_61573), .Q(regs_5
		[14]));
	notech_mux2 i_6675(.S(\nbus_11332[0] ), .A(regs_5[14]), .B(n_17864), .Z(n_20137
		));
	notech_ao4 i_210936199(.A(n_56447), .B(n_28252), .C(n_56432), .D(n_28217
		), .Z(n_2237));
	notech_reg regs_reg_5_15(.CP(n_62714), .D(n_20144), .CD(n_61572), .Q(regs_5
		[15]));
	notech_mux2 i_6683(.S(\nbus_11332[0] ), .A(regs_5[15]), .B(n_27415), .Z(n_20144
		));
	notech_reg regs_reg_5_16(.CP(n_62714), .D(n_20152), .CD(n_61573), .Q(regs_5
		[16]));
	notech_mux2 i_6691(.S(n_54854), .A(regs_5[16]), .B(n_27416), .Z(n_20152)
		);
	notech_ao4 i_211136197(.A(n_56908), .B(n_29608), .C(n_56427), .D(n_28382
		), .Z(n_2235));
	notech_reg regs_reg_5_17(.CP(n_62714), .D(n_20159), .CD(n_61583), .Q(regs_5
		[17]));
	notech_mux2 i_6699(.S(n_54854), .A(regs_5[17]), .B(n_27417), .Z(n_20159)
		);
	notech_ao4 i_211236196(.A(n_56414), .B(n_28446), .C(n_56405), .D(n_28588
		), .Z(n_2234));
	notech_reg regs_reg_5_18(.CP(n_62714), .D(n_20167), .CD(n_61583), .Q(regs_5
		[18]));
	notech_mux2 i_6707(.S(n_54854), .A(regs_5[18]), .B(n_27418), .Z(n_20167)
		);
	notech_reg regs_reg_5_19(.CP(n_62714), .D(n_20174), .CD(n_61583), .Q(regs_5
		[19]));
	notech_mux2 i_6715(.S(n_54854), .A(regs_5[19]), .B(n_27419), .Z(n_20174)
		);
	notech_reg regs_reg_5_20(.CP(n_62714), .D(n_20182), .CD(n_61583), .Q(regs_5
		[20]));
	notech_mux2 i_6723(.S(n_54854), .A(regs_5[20]), .B(n_17900), .Z(n_20182)
		);
	notech_ao4 i_211536193(.A(n_57976), .B(n_28303), .C(n_60845), .D(n_28496
		), .Z(n_2231));
	notech_reg regs_reg_5_21(.CP(n_62714), .D(n_20189), .CD(n_61583), .Q(regs_5
		[21]));
	notech_mux2 i_6731(.S(n_54854), .A(regs_5[21]), .B(n_27420), .Z(n_20189)
		);
	notech_ao4 i_211636192(.A(n_58009), .B(n_27871), .C(n_56463), .D(n_29622
		), .Z(n_2230));
	notech_reg regs_reg_5_22(.CP(n_62714), .D(n_20197), .CD(n_61584), .Q(regs_5
		[22]));
	notech_mux2 i_6739(.S(n_54854), .A(regs_5[22]), .B(n_17912), .Z(n_20197)
		);
	notech_and2 i_212036188(.A(n_2228), .B(n_2227), .Z(n_2229));
	notech_reg regs_reg_5_23(.CP(n_62714), .D(n_20204), .CD(n_61584), .Q(regs_5
		[23]));
	notech_mux2 i_6747(.S(n_54854), .A(regs_5[23]), .B(n_17918), .Z(n_20204)
		);
	notech_ao4 i_211836190(.A(n_56400), .B(n_28171), .C(n_56385), .D(n_28400
		), .Z(n_2228));
	notech_reg regs_reg_5_24(.CP(n_62714), .D(n_20212), .CD(n_61584), .Q(regs_5
		[24]));
	notech_mux2 i_6755(.S(n_54854), .A(regs_5[24]), .B(n_17924), .Z(n_20212)
		);
	notech_ao4 i_211936189(.A(n_59344), .B(n_28534), .C(n_56371), .D(n_28336
		), .Z(n_2227));
	notech_reg regs_reg_5_25(.CP(n_62714), .D(n_20219), .CD(n_61584), .Q(regs_5
		[25]));
	notech_mux2 i_6763(.S(n_54854), .A(regs_5[25]), .B(n_17930), .Z(n_20219)
		);
	notech_and4 i_212836180(.A(n_2224), .B(n_2223), .C(n_2221), .D(n_2220), 
		.Z(n_2226));
	notech_reg regs_reg_5_26(.CP(n_62714), .D(n_20229), .CD(n_61583), .Q(regs_5
		[26]));
	notech_mux2 i_6771(.S(n_54854), .A(regs_5[26]), .B(n_17936), .Z(n_20229)
		);
	notech_reg regs_reg_5_27(.CP(n_62714), .D(n_20238), .CD(n_61583), .Q(regs_5
		[27]));
	notech_mux2 i_6779(.S(n_54854), .A(regs_5[27]), .B(n_17942), .Z(n_20238)
		);
	notech_ao4 i_212236186(.A(n_56452), .B(n_28270), .C(n_58024), .D(n_28464
		), .Z(n_2224));
	notech_reg regs_reg_5_28(.CP(n_62714), .D(n_20246), .CD(n_61583), .Q(regs_5
		[28]));
	notech_mux2 i_6787(.S(n_54854), .A(regs_5[28]), .B(n_17948), .Z(n_20246)
		);
	notech_ao4 i_212336185(.A(n_56447), .B(n_28238), .C(n_56432), .D(n_28203
		), .Z(n_2223));
	notech_reg regs_reg_5_29(.CP(n_62714), .D(n_20253), .CD(n_61582), .Q(regs_5
		[29]));
	notech_mux2 i_6795(.S(n_54854), .A(regs_5[29]), .B(n_17954), .Z(n_20253)
		);
	notech_reg regs_reg_5_30(.CP(n_62714), .D(n_20259), .CD(n_61582), .Q(regs_5
		[30]));
	notech_mux2 i_6803(.S(n_54854), .A(regs_5[30]), .B(n_17960), .Z(n_20259)
		);
	notech_ao4 i_212536183(.A(n_56908), .B(n_29623), .C(n_56427), .D(n_28368
		), .Z(n_2221));
	notech_reg regs_reg_5_31(.CP(n_62714), .D(n_20265), .CD(n_61583), .Q(regs_5
		[31]));
	notech_mux2 i_6811(.S(n_54854), .A(regs_5[31]), .B(n_17966), .Z(n_20265)
		);
	notech_ao4 i_212636182(.A(n_56414), .B(n_28432), .C(n_56405), .D(n_28574
		), .Z(n_2220));
	notech_reg sav_cs_reg_0(.CP(n_62714), .D(n_20271), .CD(n_61583), .Q(sav_cs
		[0]));
	notech_mux2 i_6819(.S(n_60136), .A(cs[0]), .B(sav_cs[0]), .Z(n_20271));
	notech_reg sav_cs_reg_1(.CP(n_62714), .D(n_20277), .CD(n_61583), .Q(sav_cs
		[1]));
	notech_mux2 i_6827(.S(n_60136), .A(cs[1]), .B(sav_cs[1]), .Z(n_20277));
	notech_nao3 i_2838206(.A(instrc[123]), .B(n_60975), .C(instrc[120]), .Z(n_101413114
		));
	notech_reg tss_esp0_reg(.CP(n_62638), .D(n_20283), .CD(n_61583), .Q(tss_esp0
		));
	notech_mux2 i_6835(.S(n_19896), .A(tss_esp0), .B(n_60318), .Z(n_20283)
		);
	notech_reg_set temp_sp_reg_0(.CP(n_62638), .D(n_20289), .SD(1'b1), .Q(temp_sp
		[0]));
	notech_mux2 i_6843(.S(\nbus_11363[0] ), .A(temp_sp[0]), .B(n_27421), .Z(n_20289
		));
	notech_reg_set temp_sp_reg_1(.CP(n_62638), .D(n_20295), .SD(1'b1), .Q(temp_sp
		[1]));
	notech_mux2 i_6851(.S(\nbus_11363[0] ), .A(temp_sp[1]), .B(n_27423), .Z(n_20295
		));
	notech_reg_set temp_sp_reg_2(.CP(n_62638), .D(n_20301), .SD(1'b1), .Q(temp_sp
		[2]));
	notech_mux2 i_6859(.S(\nbus_11363[0] ), .A(temp_sp[2]), .B(n_27425), .Z(n_20301
		));
	notech_reg_set temp_sp_reg_3(.CP(n_62638), .D(n_20307), .SD(1'b1), .Q(temp_sp
		[3]));
	notech_mux2 i_6867(.S(\nbus_11363[0] ), .A(temp_sp[3]), .B(n_27427), .Z(n_20307
		));
	notech_reg_set temp_sp_reg_4(.CP(n_62638), .D(n_20316), .SD(1'b1), .Q(temp_sp
		[4]));
	notech_mux2 i_6875(.S(\nbus_11363[0] ), .A(temp_sp[4]), .B(n_27429), .Z(n_20316
		));
	notech_reg_set temp_sp_reg_5(.CP(n_62638), .D(n_20322), .SD(1'b1), .Q(temp_sp
		[5]));
	notech_mux2 i_6883(.S(\nbus_11363[0] ), .A(temp_sp[5]), .B(n_27431), .Z(n_20322
		));
	notech_reg_set temp_sp_reg_6(.CP(n_62638), .D(n_20328), .SD(1'b1), .Q(temp_sp
		[6]));
	notech_mux2 i_6891(.S(\nbus_11363[0] ), .A(temp_sp[6]), .B(n_27433), .Z(n_20328
		));
	notech_reg_set temp_sp_reg_7(.CP(n_62638), .D(n_20334), .SD(1'b1), .Q(temp_sp
		[7]));
	notech_mux2 i_6899(.S(\nbus_11363[0] ), .A(temp_sp[7]), .B(n_27435), .Z(n_20334
		));
	notech_reg_set temp_sp_reg_8(.CP(n_62638), .D(n_20340), .SD(1'b1), .Q(temp_sp
		[8]));
	notech_mux2 i_6907(.S(\nbus_11363[0] ), .A(temp_sp[8]), .B(n_27438), .Z(n_20340
		));
	notech_reg_set temp_sp_reg_9(.CP(n_62712), .D(n_20346), .SD(1'b1), .Q(temp_sp
		[9]));
	notech_mux2 i_6915(.S(\nbus_11363[0] ), .A(temp_sp[9]), .B(n_27440), .Z(n_20346
		));
	notech_reg_set temp_sp_reg_10(.CP(n_62706), .D(n_20352), .SD(1'b1), .Q(temp_sp
		[10]));
	notech_mux2 i_6923(.S(\nbus_11363[0] ), .A(temp_sp[10]), .B(n_27442), .Z
		(n_20352));
	notech_reg_set temp_sp_reg_11(.CP(n_62706), .D(n_20358), .SD(1'b1), .Q(temp_sp
		[11]));
	notech_mux2 i_6931(.S(\nbus_11363[0] ), .A(temp_sp[11]), .B(n_27444), .Z
		(n_20358));
	notech_reg_set temp_sp_reg_12(.CP(n_62706), .D(n_20364), .SD(1'b1), .Q(temp_sp
		[12]));
	notech_mux2 i_6939(.S(\nbus_11363[0] ), .A(temp_sp[12]), .B(n_27446), .Z
		(n_20364));
	notech_reg_set temp_sp_reg_13(.CP(n_62706), .D(n_20370), .SD(1'b1), .Q(temp_sp
		[13]));
	notech_mux2 i_6947(.S(\nbus_11363[0] ), .A(temp_sp[13]), .B(n_27448), .Z
		(n_20370));
	notech_reg_set temp_sp_reg_14(.CP(n_62706), .D(n_20376), .SD(1'b1), .Q(temp_sp
		[14]));
	notech_mux2 i_6955(.S(\nbus_11363[0] ), .A(temp_sp[14]), .B(n_27450), .Z
		(n_20376));
	notech_reg_set temp_sp_reg_15(.CP(n_62706), .D(n_20382), .SD(1'b1), .Q(temp_sp
		[15]));
	notech_mux2 i_6963(.S(\nbus_11363[0] ), .A(temp_sp[15]), .B(n_27452), .Z
		(n_20382));
	notech_reg_set temp_sp_reg_16(.CP(n_62706), .D(n_20388), .SD(1'b1), .Q(temp_sp
		[16]));
	notech_mux2 i_6971(.S(n_54420), .A(temp_sp[16]), .B(n_27454), .Z(n_20388
		));
	notech_reg_set temp_sp_reg_17(.CP(n_62706), .D(n_20395), .SD(1'b1), .Q(temp_sp
		[17]));
	notech_mux2 i_6979(.S(n_54420), .A(temp_sp[17]), .B(n_27456), .Z(n_20395
		));
	notech_reg_set temp_sp_reg_18(.CP(n_62706), .D(n_20403), .SD(1'b1), .Q(temp_sp
		[18]));
	notech_mux2 i_6987(.S(n_54420), .A(temp_sp[18]), .B(n_27458), .Z(n_20403
		));
	notech_reg_set temp_sp_reg_19(.CP(n_62706), .D(n_20409), .SD(1'b1), .Q(temp_sp
		[19]));
	notech_mux2 i_6995(.S(n_54420), .A(temp_sp[19]), .B(n_27460), .Z(n_20409
		));
	notech_reg_set temp_sp_reg_20(.CP(n_62706), .D(n_20415), .SD(1'b1), .Q(temp_sp
		[20]));
	notech_mux2 i_7003(.S(n_54420), .A(temp_sp[20]), .B(n_27462), .Z(n_20415
		));
	notech_reg_set temp_sp_reg_21(.CP(n_62706), .D(n_20421), .SD(1'b1), .Q(temp_sp
		[21]));
	notech_mux2 i_7011(.S(n_54420), .A(temp_sp[21]), .B(n_27464), .Z(n_20421
		));
	notech_reg_set temp_sp_reg_22(.CP(n_62750), .D(n_20427), .SD(1'b1), .Q(temp_sp
		[22]));
	notech_mux2 i_7019(.S(n_54420), .A(temp_sp[22]), .B(n_27466), .Z(n_20427
		));
	notech_reg_set temp_sp_reg_23(.CP(n_62750), .D(n_20433), .SD(1'b1), .Q(temp_sp
		[23]));
	notech_mux2 i_7027(.S(n_54420), .A(temp_sp[23]), .B(n_27470), .Z(n_20433
		));
	notech_reg_set temp_sp_reg_24(.CP(n_62750), .D(n_20439), .SD(1'b1), .Q(temp_sp
		[24]));
	notech_mux2 i_7035(.S(n_54420), .A(temp_sp[24]), .B(n_27472), .Z(n_20439
		));
	notech_reg_set temp_sp_reg_25(.CP(n_62750), .D(n_20445), .SD(1'b1), .Q(temp_sp
		[25]));
	notech_mux2 i_7043(.S(n_54420), .A(temp_sp[25]), .B(n_27474), .Z(n_20445
		));
	notech_reg_set temp_sp_reg_26(.CP(n_62750), .D(n_20451), .SD(1'b1), .Q(temp_sp
		[26]));
	notech_mux2 i_7051(.S(n_54420), .A(temp_sp[26]), .B(n_27476), .Z(n_20451
		));
	notech_reg_set temp_sp_reg_27(.CP(n_62750), .D(n_20457), .SD(1'b1), .Q(temp_sp
		[27]));
	notech_mux2 i_7059(.S(n_54420), .A(temp_sp[27]), .B(n_27478), .Z(n_20457
		));
	notech_reg_set temp_sp_reg_28(.CP(n_62750), .D(n_20463), .SD(1'b1), .Q(temp_sp
		[28]));
	notech_mux2 i_7067(.S(n_54420), .A(temp_sp[28]), .B(n_27480), .Z(n_20463
		));
	notech_reg_set temp_sp_reg_29(.CP(n_62750), .D(n_20469), .SD(1'b1), .Q(temp_sp
		[29]));
	notech_mux2 i_7075(.S(n_54420), .A(temp_sp[29]), .B(n_27482), .Z(n_20469
		));
	notech_reg_set temp_sp_reg_30(.CP(n_62750), .D(n_20476), .SD(1'b1), .Q(temp_sp
		[30]));
	notech_mux2 i_7083(.S(n_54420), .A(temp_sp[30]), .B(n_27484), .Z(n_20476
		));
	notech_reg_set temp_sp_reg_31(.CP(n_62750), .D(n_20484), .SD(1'b1), .Q(temp_sp
		[31]));
	notech_mux2 i_7091(.S(n_54420), .A(temp_sp[31]), .B(n_27486), .Z(n_20484
		));
	notech_reg regs_reg_4_0(.CP(n_62750), .D(n_20490), .CD(n_61583), .Q(regs_4
		[0]));
	notech_mux2 i_7099(.S(n_177458870), .A(n_27488), .B(regs_4[0]), .Z(n_20490
		));
	notech_reg regs_reg_4_1(.CP(n_62750), .D(n_20496), .CD(n_61586), .Q(regs_4
		[1]));
	notech_mux2 i_7107(.S(n_177458870), .A(n_20990), .B(regs_4[1]), .Z(n_20496
		));
	notech_reg regs_reg_4_2(.CP(n_62750), .D(n_20502), .CD(n_61586), .Q(regs_4
		[2]));
	notech_mux2 i_7115(.S(n_177458870), .A(n_20996), .B(regs_4[2]), .Z(n_20502
		));
	notech_reg regs_reg_4_3(.CP(n_62750), .D(n_20508), .CD(n_61586), .Q(regs_4
		[3]));
	notech_mux2 i_7123(.S(n_177458870), .A(n_21002), .B(regs_4[3]), .Z(n_20508
		));
	notech_reg regs_reg_4_4(.CP(n_62750), .D(n_20514), .CD(n_61586), .Q(regs_4
		[4]));
	notech_mux2 i_7131(.S(n_177458870), .A(n_21008), .B(regs_4[4]), .Z(n_20514
		));
	notech_reg regs_reg_4_5(.CP(n_62750), .D(n_20520), .CD(n_61586), .Q(regs_4
		[5]));
	notech_mux2 i_7139(.S(n_177458870), .A(n_21014), .B(regs_4[5]), .Z(n_20520
		));
	notech_reg regs_reg_4_6(.CP(n_62750), .D(n_20526), .CD(n_61586), .Q(regs_4
		[6]));
	notech_mux2 i_7147(.S(n_177458870), .A(n_21020), .B(regs_4[6]), .Z(n_20526
		));
	notech_reg regs_reg_4_7(.CP(n_62750), .D(n_20532), .CD(n_61586), .Q(regs_4
		[7]));
	notech_mux2 i_7155(.S(n_177458870), .A(n_21026), .B(regs_4[7]), .Z(n_20532
		));
	notech_reg regs_reg_4_8(.CP(n_62750), .D(n_20538), .CD(n_61586), .Q(regs_4
		[8]));
	notech_mux2 i_7163(.S(n_177458870), .A(n_21032), .B(regs_4[8]), .Z(n_20538
		));
	notech_reg regs_reg_4_9(.CP(n_62762), .D(n_20544), .CD(n_61586), .Q(regs_4
		[9]));
	notech_mux2 i_7171(.S(n_177458870), .A(n_21038), .B(regs_4[9]), .Z(n_20544
		));
	notech_reg regs_reg_4_10(.CP(n_62762), .D(n_20550), .CD(n_61586), .Q(regs_4
		[10]));
	notech_mux2 i_7179(.S(n_177458870), .A(n_21044), .B(regs_4[10]), .Z(n_20550
		));
	notech_reg regs_reg_4_11(.CP(n_62762), .D(n_20556), .CD(n_61584), .Q(regs_4
		[11]));
	notech_mux2 i_7187(.S(n_177458870), .A(n_27489), .B(regs_4[11]), .Z(n_20556
		));
	notech_reg regs_reg_4_12(.CP(n_62762), .D(n_20562), .CD(n_61584), .Q(regs_4
		[12]));
	notech_mux2 i_7195(.S(n_177458870), .A(n_21056), .B(regs_4[12]), .Z(n_20562
		));
	notech_reg regs_reg_4_13(.CP(n_62762), .D(n_20568), .CD(n_61584), .Q(regs_4
		[13]));
	notech_mux2 i_7203(.S(n_177458870), .A(n_27490), .B(regs_4[13]), .Z(n_20568
		));
	notech_reg regs_reg_4_14(.CP(n_62762), .D(n_20574), .CD(n_61584), .Q(regs_4
		[14]));
	notech_mux2 i_7211(.S(n_177458870), .A(n_27491), .B(regs_4[14]), .Z(n_20574
		));
	notech_reg regs_reg_4_15(.CP(n_62762), .D(n_20580), .CD(n_61584), .Q(regs_4
		[15]));
	notech_mux2 i_7219(.S(n_177458870), .A(n_21074), .B(regs_4[15]), .Z(n_20580
		));
	notech_reg regs_reg_4_16(.CP(n_62762), .D(n_20586), .CD(n_61584), .Q(regs_4
		[16]));
	notech_mux2 i_7227(.S(n_54905), .A(n_21080), .B(regs_4[16]), .Z(n_20586)
		);
	notech_reg regs_reg_4_17(.CP(n_62762), .D(n_20592), .CD(n_61584), .Q(regs_4
		[17]));
	notech_mux2 i_7235(.S(n_54905), .A(n_21086), .B(regs_4[17]), .Z(n_20592)
		);
	notech_reg regs_reg_4_18(.CP(n_62762), .D(n_20598), .CD(n_61584), .Q(regs_4
		[18]));
	notech_mux2 i_7243(.S(n_54905), .A(n_21092), .B(regs_4[18]), .Z(n_20598)
		);
	notech_reg regs_reg_4_19(.CP(n_62762), .D(n_20604), .CD(n_61584), .Q(regs_4
		[19]));
	notech_mux2 i_7251(.S(n_54905), .A(n_21098), .B(regs_4[19]), .Z(n_20604)
		);
	notech_reg regs_reg_4_20(.CP(n_62762), .D(n_20610), .CD(n_61578), .Q(regs_4
		[20]));
	notech_mux2 i_7259(.S(n_54905), .A(n_21104), .B(regs_4[20]), .Z(n_20610)
		);
	notech_reg regs_reg_4_21(.CP(n_62762), .D(n_20616), .CD(n_61578), .Q(regs_4
		[21]));
	notech_mux2 i_7267(.S(n_54905), .A(n_21110), .B(regs_4[21]), .Z(n_20616)
		);
	notech_reg regs_reg_4_22(.CP(n_62762), .D(n_20623), .CD(n_61578), .Q(regs_4
		[22]));
	notech_mux2 i_7275(.S(n_54905), .A(n_21116), .B(regs_4[22]), .Z(n_20623)
		);
	notech_reg regs_reg_4_23(.CP(n_62762), .D(n_20631), .CD(n_61578), .Q(regs_4
		[23]));
	notech_mux2 i_7283(.S(n_54905), .A(n_21122), .B(regs_4[23]), .Z(n_20631)
		);
	notech_reg regs_reg_4_24(.CP(n_62762), .D(n_20638), .CD(n_61581), .Q(regs_4
		[24]));
	notech_mux2 i_7291(.S(n_54905), .A(n_21128), .B(regs_4[24]), .Z(n_20638)
		);
	notech_reg regs_reg_4_25(.CP(n_62762), .D(n_20645), .CD(n_61581), .Q(regs_4
		[25]));
	notech_mux2 i_7299(.S(n_54905), .A(n_21134), .B(regs_4[25]), .Z(n_20645)
		);
	notech_reg regs_reg_4_26(.CP(n_62762), .D(n_20652), .CD(n_61581), .Q(regs_4
		[26]));
	notech_mux2 i_7307(.S(n_54905), .A(n_1637), .B(regs_4[26]), .Z(n_20652)
		);
	notech_reg regs_reg_4_27(.CP(n_62762), .D(n_20659), .CD(n_61581), .Q(regs_4
		[27]));
	notech_mux2 i_7315(.S(n_54905), .A(n_21146), .B(regs_4[27]), .Z(n_20659)
		);
	notech_reg regs_reg_4_28(.CP(n_62762), .D(n_20667), .CD(n_61581), .Q(regs_4
		[28]));
	notech_mux2 i_7323(.S(n_54905), .A(n_230659387), .B(regs_4[28]), .Z(n_20667
		));
	notech_reg regs_reg_4_29(.CP(n_62748), .D(n_20674), .CD(n_61578), .Q(regs_4
		[29]));
	notech_mux2 i_7331(.S(n_54905), .A(n_229259373), .B(regs_4[29]), .Z(n_20674
		));
	notech_reg regs_reg_4_30(.CP(n_62748), .D(n_20681), .CD(n_61578), .Q(regs_4
		[30]));
	notech_mux2 i_7339(.S(n_54905), .A(n_21164), .B(regs_4[30]), .Z(n_20681)
		);
	notech_reg regs_reg_4_31(.CP(n_62748), .D(n_20688), .CD(n_61578), .Q(regs_4
		[31]));
	notech_mux2 i_7347(.S(n_54905), .A(n_21170), .B(regs_4[31]), .Z(n_20688)
		);
	notech_reg regs_reg_3_0(.CP(n_62748), .D(n_20695), .CD(n_61577), .Q(regs_3
		[0]));
	notech_mux2 i_7355(.S(n_3816), .A(n_20618), .B(regs_3[0]), .Z(n_20695)
		);
	notech_reg regs_reg_3_1(.CP(n_62748), .D(n_20703), .CD(n_61578), .Q(regs_3
		[1]));
	notech_mux2 i_7363(.S(n_3816), .A(n_27492), .B(regs_3[1]), .Z(n_20703)
		);
	notech_reg regs_reg_3_2(.CP(n_62748), .D(n_20710), .CD(n_61578), .Q(regs_3
		[2]));
	notech_mux2 i_7371(.S(n_3816), .A(n_27494), .B(regs_3[2]), .Z(n_20710)
		);
	notech_reg regs_reg_3_3(.CP(n_62748), .D(n_20717), .CD(n_61578), .Q(regs_3
		[3]));
	notech_mux2 i_7379(.S(n_3816), .A(n_20636), .B(regs_3[3]), .Z(n_20717)
		);
	notech_reg regs_reg_3_4(.CP(n_62748), .D(n_20724), .CD(n_61578), .Q(regs_3
		[4]));
	notech_mux2 i_7387(.S(n_3816), .A(n_20642), .B(regs_3[4]), .Z(n_20724)
		);
	notech_reg regs_reg_3_5(.CP(n_62748), .D(n_20731), .CD(n_61578), .Q(regs_3
		[5]));
	notech_mux2 i_7395(.S(n_3816), .A(n_20648), .B(regs_3[5]), .Z(n_20731)
		);
	notech_reg regs_reg_3_6(.CP(n_62748), .D(n_20739), .CD(n_61578), .Q(regs_3
		[6]));
	notech_mux2 i_7403(.S(n_3816), .A(n_27495), .B(regs_3[6]), .Z(n_20739)
		);
	notech_reg regs_reg_3_7(.CP(n_62748), .D(n_20746), .CD(n_61582), .Q(regs_3
		[7]));
	notech_mux2 i_7411(.S(n_3816), .A(n_27496), .B(regs_3[7]), .Z(n_20746)
		);
	notech_reg regs_reg_3_8(.CP(n_62748), .D(n_20753), .CD(n_61582), .Q(regs_3
		[8]));
	notech_mux2 i_7419(.S(n_3816), .A(n_20666), .B(regs_3[8]), .Z(n_20753)
		);
	notech_reg regs_reg_3_9(.CP(n_62748), .D(n_20760), .CD(n_61582), .Q(regs_3
		[9]));
	notech_mux2 i_7427(.S(n_3816), .A(n_27497), .B(regs_3[9]), .Z(n_20760)
		);
	notech_reg regs_reg_3_10(.CP(n_62752), .D(n_20767), .CD(n_61582), .Q(regs_3
		[10]));
	notech_mux2 i_7435(.S(n_3816), .A(n_20678), .B(regs_3[10]), .Z(n_20767)
		);
	notech_reg regs_reg_3_11(.CP(n_62708), .D(n_20775), .CD(n_61582), .Q(regs_3
		[11]));
	notech_mux2 i_7443(.S(n_3816), .A(n_20684), .B(regs_3[11]), .Z(n_20775)
		);
	notech_reg regs_reg_3_12(.CP(n_62708), .D(n_20782), .CD(n_61582), .Q(regs_3
		[12]));
	notech_mux2 i_7451(.S(n_3816), .A(n_27498), .B(regs_3[12]), .Z(n_20782)
		);
	notech_reg regs_reg_3_13(.CP(n_62708), .D(n_20789), .CD(n_61582), .Q(regs_3
		[13]));
	notech_mux2 i_7459(.S(n_3816), .A(n_27297), .B(regs_3[13]), .Z(n_20789)
		);
	notech_reg regs_reg_3_14(.CP(n_62708), .D(n_20796), .CD(n_61582), .Q(regs_3
		[14]));
	notech_mux2 i_7467(.S(n_3816), .A(n_27499), .B(regs_3[14]), .Z(n_20796)
		);
	notech_reg regs_reg_3_15(.CP(n_62708), .D(n_20803), .CD(n_61582), .Q(regs_3
		[15]));
	notech_mux2 i_7475(.S(n_3816), .A(n_27502), .B(regs_3[15]), .Z(n_20803)
		);
	notech_reg regs_reg_3_16(.CP(n_62708), .D(n_20810), .CD(n_61582), .Q(regs_3
		[16]));
	notech_mux2 i_7483(.S(n_54943), .A(n_27503), .B(regs_3[16]), .Z(n_20810)
		);
	notech_reg regs_reg_3_17(.CP(n_62708), .D(n_20816), .CD(n_61581), .Q(regs_3
		[17]));
	notech_mux2 i_7491(.S(n_54943), .A(n_20720), .B(regs_3[17]), .Z(n_20816)
		);
	notech_reg regs_reg_3_18(.CP(n_62708), .D(n_20822), .CD(n_61581), .Q(regs_3
		[18]));
	notech_mux2 i_7499(.S(n_54943), .A(n_20726), .B(regs_3[18]), .Z(n_20822)
		);
	notech_reg regs_reg_3_19(.CP(n_62708), .D(n_20828), .CD(n_61581), .Q(regs_3
		[19]));
	notech_mux2 i_7507(.S(n_54943), .A(n_20732), .B(regs_3[19]), .Z(n_20828)
		);
	notech_reg regs_reg_3_20(.CP(n_62708), .D(n_20834), .CD(n_61581), .Q(regs_3
		[20]));
	notech_mux2 i_7515(.S(n_54943), .A(n_20738), .B(regs_3[20]), .Z(n_20834)
		);
	notech_reg regs_reg_3_21(.CP(n_62752), .D(n_20840), .CD(n_61581), .Q(regs_3
		[21]));
	notech_mux2 i_7524(.S(n_54943), .A(n_20744), .B(regs_3[21]), .Z(n_20840)
		);
	notech_reg regs_reg_3_22(.CP(n_62752), .D(n_20846), .CD(n_61581), .Q(regs_3
		[22]));
	notech_mux2 i_7532(.S(n_54943), .A(n_27504), .B(regs_3[22]), .Z(n_20846)
		);
	notech_reg regs_reg_3_23(.CP(n_62752), .D(n_20852), .CD(n_61582), .Q(regs_3
		[23]));
	notech_mux2 i_7540(.S(n_54943), .A(n_20756), .B(regs_3[23]), .Z(n_20852)
		);
	notech_reg regs_reg_3_24(.CP(n_62752), .D(n_20858), .CD(n_61581), .Q(regs_3
		[24]));
	notech_mux2 i_7548(.S(n_54943), .A(n_27506), .B(regs_3[24]), .Z(n_20858)
		);
	notech_reg regs_reg_3_25(.CP(n_62752), .D(n_20864), .CD(n_61581), .Q(regs_3
		[25]));
	notech_mux2 i_7556(.S(n_54943), .A(n_20768), .B(regs_3[25]), .Z(n_20864)
		);
	notech_reg regs_reg_3_26(.CP(n_62752), .D(n_20870), .CD(n_61491), .Q(regs_3
		[26]));
	notech_mux2 i_7564(.S(n_54943), .A(n_27507), .B(regs_3[26]), .Z(n_20870)
		);
	notech_reg regs_reg_3_27(.CP(n_62752), .D(n_20876), .CD(n_61491), .Q(regs_3
		[27]));
	notech_mux2 i_7572(.S(n_54943), .A(n_20780), .B(regs_3[27]), .Z(n_20876)
		);
	notech_reg regs_reg_3_28(.CP(n_62752), .D(n_20882), .CD(n_61491), .Q(regs_3
		[28]));
	notech_mux2 i_7580(.S(n_54943), .A(n_27020), .B(regs_3[28]), .Z(n_20882)
		);
	notech_reg regs_reg_3_29(.CP(n_62752), .D(n_20888), .CD(n_61491), .Q(regs_3
		[29]));
	notech_mux2 i_7588(.S(n_54943), .A(n_27508), .B(regs_3[29]), .Z(n_20888)
		);
	notech_reg regs_reg_3_30(.CP(n_62752), .D(n_20894), .CD(n_61492), .Q(regs_3
		[30]));
	notech_mux2 i_7596(.S(n_54943), .A(n_27510), .B(regs_3[30]), .Z(n_20894)
		);
	notech_reg regs_reg_3_31(.CP(n_62752), .D(n_20900), .CD(n_61492), .Q(regs_3
		[31]));
	notech_mux2 i_7604(.S(n_54943), .A(n_27511), .B(regs_3[31]), .Z(n_20900)
		);
	notech_reg_set cr0_reg_0(.CP(n_62752), .D(n_20906), .SD(n_61492), .Q(\nbus_14526[0] 
		));
	notech_mux2 i_7612(.S(n_328290780), .A(opa[0]), .B(n_60542), .Z(n_20906)
		);
	notech_reg cr0_reg_1(.CP(n_62752), .D(n_20912), .CD(n_61492), .Q(\nbus_14522[1] 
		));
	notech_mux2 i_7620(.S(n_328290780), .A(opa[1]), .B(\nbus_14522[1] ), .Z(n_20912
		));
	notech_reg cr0_reg_2(.CP(n_62752), .D(n_20918), .CD(n_61492), .Q(cr0[2])
		);
	notech_mux2 i_7628(.S(n_328290780), .A(opa[2]), .B(cr0[2]), .Z(n_20918)
		);
	notech_reg cr0_reg_3(.CP(n_62752), .D(n_20924), .CD(n_61491), .Q(\nbus_14522[3] 
		));
	notech_mux2 i_7636(.S(n_328290780), .A(opa[3]), .B(\nbus_14522[3] ), .Z(n_20924
		));
	notech_reg cr0_reg_4(.CP(n_62752), .D(n_20930), .CD(n_61491), .Q(\nbus_14522[4] 
		));
	notech_mux2 i_7644(.S(n_328290780), .A(opa[4]), .B(\nbus_14522[4] ), .Z(n_20930
		));
	notech_reg cr0_reg_5(.CP(n_62752), .D(n_20936), .CD(n_61491), .Q(\nbus_14522[5] 
		));
	notech_mux2 i_7652(.S(n_328290780), .A(opa[5]), .B(\nbus_14522[5] ), .Z(n_20936
		));
	notech_reg cr0_reg_6(.CP(n_62752), .D(n_20942), .CD(n_61488), .Q(\nbus_14522[6] 
		));
	notech_mux2 i_7662(.S(n_328290780), .A(opa[6]), .B(\nbus_14522[6] ), .Z(n_20942
		));
	notech_reg cr0_reg_7(.CP(n_62708), .D(n_20948), .CD(n_61488), .Q(\nbus_14522[7] 
		));
	notech_mux2 i_7670(.S(n_328290780), .A(opa[7]), .B(\nbus_14522[7] ), .Z(n_20948
		));
	notech_reg cr0_reg_8(.CP(n_62708), .D(n_20954), .CD(n_61491), .Q(\nbus_14522[8] 
		));
	notech_mux2 i_7678(.S(n_328290780), .A(opa[8]), .B(\nbus_14522[8] ), .Z(n_20954
		));
	notech_reg cr0_reg_9(.CP(n_62710), .D(n_20960), .CD(n_61491), .Q(\nbus_14522[9] 
		));
	notech_mux2 i_7686(.S(n_328290780), .A(opa[9]), .B(\nbus_14522[9] ), .Z(n_20960
		));
	notech_reg cr0_reg_10(.CP(n_62710), .D(n_20966), .CD(n_61491), .Q(\nbus_14522[10] 
		));
	notech_mux2 i_7694(.S(n_328290780), .A(opa[10]), .B(\nbus_14522[10] ), .Z
		(n_20966));
	notech_reg cr0_reg_11(.CP(n_62710), .D(n_20972), .CD(n_61491), .Q(\nbus_14522[11] 
		));
	notech_mux2 i_7702(.S(n_328290780), .A(opa[11]), .B(\nbus_14522[11] ), .Z
		(n_20972));
	notech_reg cr0_reg_12(.CP(n_62710), .D(n_20978), .CD(n_61491), .Q(\nbus_14522[12] 
		));
	notech_mux2 i_7710(.S(n_328290780), .A(opa[12]), .B(\nbus_14522[12] ), .Z
		(n_20978));
	notech_reg cr0_reg_13(.CP(n_62710), .D(n_20985), .CD(n_61493), .Q(\nbus_14522[13] 
		));
	notech_mux2 i_7718(.S(n_328290780), .A(opa[13]), .B(\nbus_14522[13] ), .Z
		(n_20985));
	notech_reg cr0_reg_14(.CP(n_62710), .D(n_20992), .CD(n_61493), .Q(\nbus_14522[14] 
		));
	notech_mux2 i_7727(.S(n_328290780), .A(opa[14]), .B(\nbus_14522[14] ), .Z
		(n_20992));
	notech_reg cr0_reg_15(.CP(n_62710), .D(n_20999), .CD(n_61493), .Q(\nbus_14522[15] 
		));
	notech_mux2 i_7735(.S(n_328290780), .A(opa[15]), .B(\nbus_14522[15] ), .Z
		(n_20999));
	notech_reg cr0_reg_16(.CP(n_62710), .D(n_21006), .CD(n_61493), .Q(cr0[16
		]));
	notech_mux2 i_7743(.S(n_60830), .A(opa[16]), .B(cr0[16]), .Z(n_21006));
	notech_reg cr0_reg_17(.CP(n_62710), .D(n_21013), .CD(n_61493), .Q(\nbus_14522[17] 
		));
	notech_mux2 i_7751(.S(n_60830), .A(opa[17]), .B(\nbus_14522[17] ), .Z(n_21013
		));
	notech_reg cr0_reg_18(.CP(n_62710), .D(n_21021), .CD(n_61493), .Q(\nbus_14522[18] 
		));
	notech_mux2 i_7759(.S(n_60830), .A(opa[18]), .B(\nbus_14522[18] ), .Z(n_21021
		));
	notech_reg cr0_reg_19(.CP(n_62710), .D(n_21028), .CD(n_61493), .Q(\nbus_14522[19] 
		));
	notech_mux2 i_7767(.S(n_60830), .A(opa[19]), .B(\nbus_14522[19] ), .Z(n_21028
		));
	notech_reg cr0_reg_20(.CP(n_62710), .D(n_21035), .CD(n_61493), .Q(\nbus_14522[20] 
		));
	notech_mux2 i_7776(.S(n_60830), .A(opa[20]), .B(\nbus_14522[20] ), .Z(n_21035
		));
	notech_reg cr0_reg_21(.CP(n_62710), .D(n_21042), .CD(n_61493), .Q(\nbus_14522[21] 
		));
	notech_mux2 i_7785(.S(n_60830), .A(opa[21]), .B(\nbus_14522[21] ), .Z(n_21042
		));
	notech_reg cr0_reg_22(.CP(n_62710), .D(n_21049), .CD(n_61493), .Q(\nbus_14522[22] 
		));
	notech_mux2 i_7793(.S(n_60830), .A(opa[22]), .B(\nbus_14522[22] ), .Z(n_21049
		));
	notech_reg cr0_reg_23(.CP(n_62710), .D(n_21057), .CD(n_61492), .Q(\nbus_14522[23] 
		));
	notech_mux2 i_7801(.S(n_60830), .A(opa[23]), .B(\nbus_14522[23] ), .Z(n_21057
		));
	notech_reg cr0_reg_24(.CP(n_62710), .D(n_21064), .CD(n_61492), .Q(\nbus_14522[24] 
		));
	notech_mux2 i_7809(.S(n_60830), .A(opa[24]), .B(\nbus_14522[24] ), .Z(n_21064
		));
	notech_reg cr0_reg_25(.CP(n_62710), .D(n_21071), .CD(n_61492), .Q(\nbus_14522[25] 
		));
	notech_mux2 i_7817(.S(n_60830), .A(opa[25]), .B(\nbus_14522[25] ), .Z(n_21071
		));
	notech_reg cr0_reg_26(.CP(n_62710), .D(n_21078), .CD(n_61492), .Q(\nbus_14522[26] 
		));
	notech_mux2 i_7825(.S(n_60830), .A(opa[26]), .B(\nbus_14522[26] ), .Z(n_21078
		));
	notech_reg cr0_reg_27(.CP(n_62710), .D(n_21085), .CD(n_61492), .Q(\nbus_14522[27] 
		));
	notech_mux2 i_7833(.S(n_60830), .A(opa[27]), .B(\nbus_14522[27] ), .Z(n_21085
		));
	notech_reg cr0_reg_28(.CP(n_62636), .D(n_21093), .CD(n_61493), .Q(\nbus_14522[28] 
		));
	notech_mux2 i_7841(.S(n_60830), .A(opa[28]), .B(\nbus_14522[28] ), .Z(n_21093
		));
	notech_reg cr0_reg_29(.CP(n_62636), .D(n_21100), .CD(n_61493), .Q(\nbus_14522[29] 
		));
	notech_mux2 i_7849(.S(n_60830), .A(opa[29]), .B(\nbus_14522[29] ), .Z(n_21100
		));
	notech_reg cr0_reg_30(.CP(n_62636), .D(n_21107), .CD(n_61492), .Q(\nbus_14522[30] 
		));
	notech_mux2 i_7857(.S(n_60830), .A(opa[30]), .B(\nbus_14522[30] ), .Z(n_21107
		));
	notech_reg cr0_reg_31(.CP(n_62636), .D(n_21114), .CD(n_61492), .Q(\nbus_14522[31] 
		));
	notech_mux2 i_7865(.S(n_60830), .A(opa[31]), .B(\nbus_14522[31] ), .Z(n_21114
		));
	notech_reg mask8b_reg_0(.CP(n_62636), .D(n_21121), .CD(n_61486), .Q(mask8b
		[0]));
	notech_mux2 i_7873(.S(\nbus_11326[0] ), .A(mask8b[0]), .B(n_27540), .Z(n_21121
		));
	notech_reg mask8b_reg_1(.CP(n_62636), .D(n_21129), .CD(n_61486), .Q(mask8b
		[1]));
	notech_mux2 i_7881(.S(\nbus_11326[0] ), .A(mask8b[1]), .B(n_27542), .Z(n_21129
		));
	notech_reg mask8b_reg_2(.CP(n_62636), .D(n_21136), .CD(n_61486), .Q(mask8b
		[2]));
	notech_mux2 i_7889(.S(\nbus_11326[0] ), .A(mask8b[2]), .B(n_16501), .Z(n_21136
		));
	notech_reg opb_reg_0(.CP(n_62636), .D(n_21143), .CD(n_61486), .Q(opb[0])
		);
	notech_mux2 i_7897(.S(n_3817), .A(n_19106), .B(opb[0]), .Z(n_21143));
	notech_reg opb_reg_1(.CP(n_62636), .D(n_21150), .CD(n_61486), .Q(opb[1])
		);
	notech_mux2 i_7905(.S(n_3817), .A(n_19112), .B(opb[1]), .Z(n_21150));
	notech_reg opb_reg_2(.CP(n_62636), .D(n_21157), .CD(n_61487), .Q(opb[2])
		);
	notech_mux2 i_7913(.S(n_3817), .A(n_3881), .B(opb[2]), .Z(n_21157));
	notech_reg opb_reg_3(.CP(n_62636), .D(n_21165), .CD(n_61487), .Q(opb[3])
		);
	notech_mux2 i_7921(.S(n_3817), .A(n_19124), .B(opb[3]), .Z(n_21165));
	notech_reg opb_reg_4(.CP(n_62636), .D(n_21172), .CD(n_61486), .Q(opb[4])
		);
	notech_mux2 i_7929(.S(n_3817), .A(n_19130), .B(opb[4]), .Z(n_21172));
	notech_reg opb_reg_5(.CP(n_62718), .D(n_21178), .CD(n_61487), .Q(opb[5])
		);
	notech_mux2 i_7937(.S(n_3817), .A(n_19136), .B(opb[5]), .Z(n_21178));
	notech_reg opb_reg_6(.CP(n_62568), .D(n_21184), .CD(n_61486), .Q(opb[6])
		);
	notech_mux2 i_7945(.S(n_3817), .A(n_19142), .B(opb[6]), .Z(n_21184));
	notech_reg opb_reg_7(.CP(n_62568), .D(n_21190), .CD(n_61485), .Q(opb[7])
		);
	notech_mux2 i_7953(.S(n_3817), .A(n_19148), .B(opb[7]), .Z(n_21190));
	notech_reg opb_reg_8(.CP(n_62568), .D(n_21196), .CD(n_61485), .Q(opb[8])
		);
	notech_mux2 i_7961(.S(n_3817), .A(n_27543), .B(opb[8]), .Z(n_21196));
	notech_reg opb_reg_9(.CP(n_62568), .D(n_21202), .CD(n_61485), .Q(opb[9])
		);
	notech_mux2 i_7969(.S(n_3817), .A(n_27544), .B(opb[9]), .Z(n_21202));
	notech_reg opb_reg_10(.CP(n_62568), .D(n_21208), .CD(n_61485), .Q(opb[10
		]));
	notech_mux2 i_7977(.S(n_3817), .A(n_27545), .B(opb[10]), .Z(n_21208));
	notech_reg opb_reg_11(.CP(n_62568), .D(n_21214), .CD(n_61486), .Q(opb[11
		]));
	notech_mux2 i_7985(.S(n_3817), .A(n_27546), .B(opb[11]), .Z(n_21214));
	notech_reg opb_reg_12(.CP(n_62568), .D(n_21220), .CD(n_61486), .Q(opb[12
		]));
	notech_mux2 i_7993(.S(n_3817), .A(n_27547), .B(opb[12]), .Z(n_21220));
	notech_reg opb_reg_13(.CP(n_62568), .D(n_21226), .CD(n_61486), .Q(opb[13
		]));
	notech_mux2 i_8001(.S(n_3817), .A(n_27548), .B(opb[13]), .Z(n_21226));
	notech_nand2 i_2638208(.A(instrc[120]), .B(instrc[123]), .Z(n_32339));
	notech_reg opb_reg_14(.CP(n_62568), .D(n_21232), .CD(n_61486), .Q(opb[14
		]));
	notech_mux2 i_8009(.S(n_3817), .A(n_27549), .B(opb[14]), .Z(n_21232));
	notech_nor2 i_1838216(.A(instrc[120]), .B(n_29180), .Z(n_32367));
	notech_reg opb_reg_15(.CP(n_62568), .D(n_21238), .CD(n_61486), .Q(opb[15
		]));
	notech_mux2 i_8017(.S(n_3817), .A(n_19196), .B(opb[15]), .Z(n_21238));
	notech_reg opb_reg_16(.CP(n_62648), .D(n_21244), .CD(n_61488), .Q(opb[16
		]));
	notech_mux2 i_8025(.S(n_27550), .A(opb[16]), .B(n_19202), .Z(n_21244));
	notech_reg opb_reg_17(.CP(n_62648), .D(n_21250), .CD(n_61488), .Q(opb[17
		]));
	notech_mux2 i_8033(.S(n_27550), .A(opb[17]), .B(n_19208), .Z(n_21250));
	notech_ao4 i_192039479(.A(n_56666), .B(n_28235), .C(n_56653), .D(n_28201
		), .Z(n_2071));
	notech_reg opb_reg_18(.CP(n_62648), .D(n_21256), .CD(n_61488), .Q(opb[18
		]));
	notech_mux2 i_8041(.S(n_27550), .A(opb[18]), .B(n_19214), .Z(n_21256));
	notech_ao4 i_192139478(.A(n_56916), .B(n_29621), .C(n_56640), .D(n_28268
		), .Z(n_2070));
	notech_reg opb_reg_19(.CP(n_62648), .D(n_21262), .CD(n_61488), .Q(opb[19
		]));
	notech_mux2 i_8049(.S(n_27550), .A(opb[19]), .B(n_19220), .Z(n_21262));
	notech_and2 i_192539474(.A(n_2068), .B(n_2067), .Z(n_2069));
	notech_reg opb_reg_20(.CP(n_62648), .D(n_21268), .CD(n_61488), .Q(opb[20
		]));
	notech_mux2 i_8057(.S(n_27550), .A(opb[20]), .B(n_19226), .Z(n_21268));
	notech_ao4 i_192339476(.A(n_56532), .B(n_28301), .C(n_56518), .D(n_29620
		), .Z(n_2068));
	notech_reg opb_reg_21(.CP(n_62648), .D(n_21274), .CD(n_61488), .Q(opb[21
		]));
	notech_mux2 i_8065(.S(n_27550), .A(opb[21]), .B(n_19232), .Z(n_21274));
	notech_ao4 i_192439475(.A(n_56502), .B(n_28366), .C(n_56489), .D(n_28334
		), .Z(n_2067));
	notech_reg opb_reg_22(.CP(n_62648), .D(n_21280), .CD(n_61488), .Q(opb[22
		]));
	notech_mux2 i_8073(.S(n_27550), .A(opb[22]), .B(n_19238), .Z(n_21280));
	notech_and4 i_193339466(.A(n_2064), .B(n_2063), .C(n_2061), .D(n_2060), 
		.Z(n_2066));
	notech_reg opb_reg_23(.CP(n_62648), .D(n_21286), .CD(n_61488), .Q(opb[23
		]));
	notech_mux2 i_8081(.S(n_27550), .A(opb[23]), .B(n_19244), .Z(n_21286));
	notech_reg opb_reg_24(.CP(n_62648), .D(n_21292), .CD(n_61488), .Q(opb[24
		]));
	notech_mux2 i_8089(.S(n_27550), .A(opb[24]), .B(n_19250), .Z(n_21292));
	notech_ao4 i_192739472(.A(n_56627), .B(n_28430), .C(n_56614), .D(n_28398
		), .Z(n_2064));
	notech_reg opb_reg_25(.CP(n_62648), .D(n_21298), .CD(n_61488), .Q(opb[25
		]));
	notech_mux2 i_8097(.S(n_27550), .A(opb[25]), .B(n_19256), .Z(n_21298));
	notech_ao4 i_192839471(.A(n_56605), .B(n_28462), .C(n_56592), .D(n_28169
		), .Z(n_2063));
	notech_reg opb_reg_26(.CP(n_62648), .D(n_21304), .CD(n_61487), .Q(opb[26
		]));
	notech_mux2 i_8105(.S(n_27550), .A(opb[26]), .B(n_19262), .Z(n_21304));
	notech_reg opb_reg_27(.CP(n_62648), .D(n_21310), .CD(n_61487), .Q(opb[27
		]));
	notech_mux2 i_8113(.S(n_27550), .A(opb[27]), .B(n_19268), .Z(n_21310));
	notech_ao4 i_193039469(.A(n_56583), .B(n_28494), .C(n_56570), .D(n_28529
		), .Z(n_2061));
	notech_reg opb_reg_28(.CP(n_62648), .D(n_21316), .CD(n_61487), .Q(opb[28
		]));
	notech_mux2 i_8121(.S(n_27550), .A(opb[28]), .B(n_19274), .Z(n_21316));
	notech_ao4 i_193139468(.A(n_56557), .B(n_27869), .C(n_56547), .D(n_28572
		), .Z(n_2060));
	notech_reg opb_reg_29(.CP(n_62648), .D(n_21322), .CD(n_61487), .Q(opb[29
		]));
	notech_mux2 i_8129(.S(n_27550), .A(opb[29]), .B(n_19280), .Z(n_21322));
	notech_reg opb_reg_30(.CP(n_62648), .D(n_21328), .CD(n_61487), .Q(opb[30
		]));
	notech_mux2 i_8137(.S(n_27550), .A(opb[30]), .B(n_19286), .Z(n_21328));
	notech_reg opb_reg_31(.CP(n_62648), .D(n_21334), .CD(n_61487), .Q(opb[31
		]));
	notech_mux2 i_8145(.S(n_27550), .A(opb[31]), .B(n_19292), .Z(n_21334));
	notech_reg regs_reg_2_0(.CP(n_62648), .D(n_21341), .CD(n_61487), .Q(regs_2
		[0]));
	notech_mux2 i_8153(.S(n_27575), .A(regs_2[0]), .B(n_27551), .Z(n_21341)
		);
	notech_reg regs_reg_2_1(.CP(n_62648), .D(n_21352), .CD(n_61487), .Q(regs_2
		[1]));
	notech_mux2 i_8162(.S(n_27575), .A(regs_2[1]), .B(n_17438), .Z(n_21352)
		);
	notech_reg regs_reg_2_2(.CP(n_62648), .D(n_21359), .CD(n_61487), .Q(regs_2
		[2]));
	notech_mux2 i_8170(.S(n_27575), .A(regs_2[2]), .B(n_27553), .Z(n_21359)
		);
	notech_ao4 i_202739374(.A(n_56666), .B(n_28238), .C(n_56653), .D(n_28203
		), .Z(n_2054));
	notech_reg regs_reg_2_3(.CP(n_62646), .D(n_21367), .CD(n_61499), .Q(regs_2
		[3]));
	notech_mux2 i_8178(.S(n_27575), .A(regs_2[3]), .B(n_17450), .Z(n_21367)
		);
	notech_ao4 i_202839373(.A(n_56916), .B(n_29623), .C(n_56640), .D(n_28270
		), .Z(n_2053));
	notech_reg regs_reg_2_4(.CP(n_62646), .D(n_21374), .CD(n_61499), .Q(regs_2
		[4]));
	notech_mux2 i_8186(.S(n_27575), .A(regs_2[4]), .B(n_27026), .Z(n_21374)
		);
	notech_and2 i_203239369(.A(n_2051), .B(n_2050), .Z(n_2052));
	notech_reg regs_reg_2_5(.CP(n_62722), .D(n_21381), .CD(n_61499), .Q(regs_2
		[5]));
	notech_mux2 i_8194(.S(n_27575), .A(regs_2[5]), .B(n_17462), .Z(n_21381)
		);
	notech_ao4 i_203039371(.A(n_56532), .B(n_28303), .C(n_56518), .D(n_29622
		), .Z(n_2051));
	notech_reg regs_reg_2_6(.CP(n_62722), .D(n_21388), .CD(n_61499), .Q(regs_2
		[6]));
	notech_mux2 i_8202(.S(n_27575), .A(regs_2[6]), .B(n_27554), .Z(n_21388)
		);
	notech_ao4 i_203139370(.A(n_56502), .B(n_28368), .C(n_56489), .D(n_28336
		), .Z(n_2050));
	notech_reg regs_reg_2_7(.CP(n_62722), .D(n_21395), .CD(n_61499), .Q(regs_2
		[7]));
	notech_mux2 i_8210(.S(n_27575), .A(regs_2[7]), .B(n_27555), .Z(n_21395)
		);
	notech_and4 i_204039361(.A(n_2047), .B(n_2046), .C(n_2044), .D(n_204392003
		), .Z(n_2049));
	notech_reg regs_reg_2_8(.CP(n_62722), .D(n_21403), .CD(n_61499), .Q(regs_2
		[8]));
	notech_mux2 i_8218(.S(n_27575), .A(regs_2[8]), .B(n_17480), .Z(n_21403)
		);
	notech_reg regs_reg_2_9(.CP(n_62722), .D(n_21410), .CD(n_61499), .Q(regs_2
		[9]));
	notech_mux2 i_8226(.S(n_27575), .A(regs_2[9]), .B(n_17486), .Z(n_21410)
		);
	notech_ao4 i_203439367(.A(n_56627), .B(n_28432), .C(n_56614), .D(n_28400
		), .Z(n_2047));
	notech_reg regs_reg_2_10(.CP(n_62722), .D(n_21417), .CD(n_61499), .Q(regs_2
		[10]));
	notech_mux2 i_8234(.S(n_27575), .A(regs_2[10]), .B(n_27556), .Z(n_21417)
		);
	notech_ao4 i_203539366(.A(n_56605), .B(n_28464), .C(n_56592), .D(n_28171
		), .Z(n_2046));
	notech_reg regs_reg_2_11(.CP(n_62722), .D(n_21424), .CD(n_61499), .Q(regs_2
		[11]));
	notech_mux2 i_8242(.S(n_27575), .A(regs_2[11]), .B(n_27557), .Z(n_21424)
		);
	notech_reg regs_reg_2_12(.CP(n_62722), .D(n_21431), .CD(n_61498), .Q(regs_2
		[12]));
	notech_mux2 i_8250(.S(n_27575), .A(regs_2[12]), .B(n_17504), .Z(n_21431)
		);
	notech_ao4 i_203739364(.A(n_56583), .B(n_28496), .C(n_56570), .D(n_28534
		), .Z(n_2044));
	notech_reg regs_reg_2_13(.CP(n_62722), .D(n_21439), .CD(n_61498), .Q(regs_2
		[13]));
	notech_mux2 i_8258(.S(n_27575), .A(regs_2[13]), .B(n_27559), .Z(n_21439)
		);
	notech_ao4 i_203839363(.A(n_56557), .B(n_27871), .C(n_56547), .D(n_28574
		), .Z(n_204392003));
	notech_reg regs_reg_2_14(.CP(n_62722), .D(n_21446), .CD(n_61498), .Q(regs_2
		[14]));
	notech_mux2 i_8266(.S(n_27575), .A(regs_2[14]), .B(n_27560), .Z(n_21446)
		);
	notech_reg regs_reg_2_15(.CP(n_62722), .D(n_21453), .CD(n_61498), .Q(regs_2
		[15]));
	notech_mux2 i_8274(.S(n_27575), .A(regs_2[15]), .B(n_17522), .Z(n_21453)
		);
	notech_reg regs_reg_2_16(.CP(n_62722), .D(n_21460), .CD(n_61498), .Q(regs_2
		[16]));
	notech_mux2 i_8282(.S(n_54963), .A(regs_2[16]), .B(n_17528), .Z(n_21460)
		);
	notech_reg regs_reg_2_17(.CP(n_62722), .D(n_21467), .CD(n_61498), .Q(regs_2
		[17]));
	notech_mux2 i_8290(.S(n_54963), .A(regs_2[17]), .B(n_27561), .Z(n_21467)
		);
	notech_reg regs_reg_2_18(.CP(n_62722), .D(n_21475), .CD(n_61498), .Q(regs_2
		[18]));
	notech_mux2 i_8298(.S(n_54963), .A(regs_2[18]), .B(n_17540), .Z(n_21475)
		);
	notech_reg regs_reg_2_19(.CP(n_62722), .D(n_21482), .CD(n_61498), .Q(regs_2
		[19]));
	notech_mux2 i_8306(.S(n_54963), .A(regs_2[19]), .B(n_27562), .Z(n_21482)
		);
	notech_reg regs_reg_2_20(.CP(n_62722), .D(n_21489), .CD(n_61498), .Q(regs_2
		[20]));
	notech_mux2 i_8314(.S(n_54963), .A(regs_2[20]), .B(n_27564), .Z(n_21489)
		);
	notech_reg regs_reg_2_21(.CP(n_62722), .D(n_21496), .CD(n_61498), .Q(regs_2
		[21]));
	notech_mux2 i_8322(.S(n_54963), .A(regs_2[21]), .B(n_17558), .Z(n_21496)
		);
	notech_reg regs_reg_2_22(.CP(n_62722), .D(n_21503), .CD(n_61502), .Q(regs_2
		[22]));
	notech_mux2 i_8330(.S(n_54963), .A(regs_2[22]), .B(n_27565), .Z(n_21503)
		);
	notech_reg regs_reg_2_23(.CP(n_62646), .D(n_21511), .CD(n_61502), .Q(regs_2
		[23]));
	notech_mux2 i_8338(.S(n_54963), .A(regs_2[23]), .B(n_27567), .Z(n_21511)
		);
	notech_reg regs_reg_2_24(.CP(n_62646), .D(n_21518), .CD(n_61502), .Q(regs_2
		[24]));
	notech_mux2 i_8346(.S(n_54963), .A(regs_2[24]), .B(n_27568), .Z(n_21518)
		);
	notech_reg regs_reg_2_25(.CP(n_62646), .D(n_21525), .CD(n_61502), .Q(regs_2
		[25]));
	notech_mux2 i_8354(.S(n_54963), .A(regs_2[25]), .B(n_27569), .Z(n_21525)
		);
	notech_reg regs_reg_2_26(.CP(n_62646), .D(n_21531), .CD(n_61502), .Q(regs_2
		[26]));
	notech_mux2 i_8362(.S(n_54963), .A(regs_2[26]), .B(n_233659417), .Z(n_21531
		));
	notech_reg regs_reg_2_27(.CP(n_62646), .D(n_21537), .CD(n_61503), .Q(regs_2
		[27]));
	notech_mux2 i_8370(.S(n_54963), .A(regs_2[27]), .B(n_17594), .Z(n_21537)
		);
	notech_reg regs_reg_2_28(.CP(n_62646), .D(n_21543), .CD(n_61503), .Q(regs_2
		[28]));
	notech_mux2 i_8378(.S(n_54963), .A(regs_2[28]), .B(n_232659407), .Z(n_21543
		));
	notech_reg regs_reg_2_29(.CP(n_62646), .D(n_21549), .CD(n_61503), .Q(regs_2
		[29]));
	notech_mux2 i_8386(.S(n_54963), .A(regs_2[29]), .B(n_1647), .Z(n_21549)
		);
	notech_reg regs_reg_2_30(.CP(n_62646), .D(n_21555), .CD(n_61503), .Q(regs_2
		[30]));
	notech_mux2 i_8394(.S(n_54963), .A(regs_2[30]), .B(n_27574), .Z(n_21555)
		);
	notech_or2 i_33904(.A(n_57020), .B(n_57042), .Z(n_26062));
	notech_reg regs_reg_2_31(.CP(n_62646), .D(n_21561), .CD(n_61502), .Q(regs_2
		[31]));
	notech_mux2 i_8403(.S(n_54963), .A(regs_2[31]), .B(n_17618), .Z(n_21561)
		);
	notech_and2 i_32621(.A(n_57055), .B(n_57082), .Z(n_2026));
	notech_reg regs_reg_1_0(.CP(n_62646), .D(n_21567), .CD(n_61499), .Q(ecx[
		0]));
	notech_mux2 i_8411(.S(\nbus_11330[0] ), .A(ecx[0]), .B(n_27576), .Z(n_21567
		));
	notech_or4 i_100040328(.A(n_59382), .B(n_246791942), .C(n_32351), .D(n_59373
		), .Z(n_2025));
	notech_reg regs_reg_1_1(.CP(n_62722), .D(n_21573), .CD(n_61502), .Q(ecx[
		1]));
	notech_mux2 i_8419(.S(\nbus_11330[0] ), .A(ecx[1]), .B(n_3842), .Z(n_21573
		));
	notech_reg regs_reg_1_2(.CP(n_62568), .D(n_21579), .CD(n_61499), .Q(ecx[
		2]));
	notech_mux2 i_8427(.S(\nbus_11330[0] ), .A(ecx[2]), .B(n_27015), .Z(n_21579
		));
	notech_reg regs_reg_1_3(.CP(n_62644), .D(n_21587), .CD(n_61499), .Q(ecx[
		3]));
	notech_mux2 i_8435(.S(\nbus_11330[0] ), .A(ecx[3]), .B(n_27005), .Z(n_21587
		));
	notech_reg regs_reg_1_4(.CP(n_62718), .D(n_21593), .CD(n_61502), .Q(ecx[
		4]));
	notech_mux2 i_8443(.S(\nbus_11330[0] ), .A(ecx[4]), .B(n_17099), .Z(n_21593
		));
	notech_reg regs_reg_1_5(.CP(n_62718), .D(n_21599), .CD(n_61502), .Q(ecx[
		5]));
	notech_mux2 i_8451(.S(\nbus_11330[0] ), .A(ecx[5]), .B(n_27006), .Z(n_21599
		));
	notech_reg regs_reg_1_6(.CP(n_62718), .D(n_21605), .CD(n_61502), .Q(ecx[
		6]));
	notech_mux2 i_8459(.S(\nbus_11330[0] ), .A(ecx[6]), .B(n_3870), .Z(n_21605
		));
	notech_reg regs_reg_1_7(.CP(n_62718), .D(n_21611), .CD(n_61502), .Q(ecx[
		7]));
	notech_mux2 i_8467(.S(\nbus_11330[0] ), .A(ecx[7]), .B(n_17117), .Z(n_21611
		));
	notech_reg regs_reg_1_8(.CP(n_62718), .D(n_21617), .CD(n_61502), .Q(ecx[
		8]));
	notech_mux2 i_8475(.S(\nbus_11330[0] ), .A(ecx[8]), .B(n_17123), .Z(n_21617
		));
	notech_reg regs_reg_1_9(.CP(n_62718), .D(n_21623), .CD(n_61496), .Q(ecx[
		9]));
	notech_mux2 i_8483(.S(\nbus_11330[0] ), .A(ecx[9]), .B(n_17129), .Z(n_21623
		));
	notech_reg regs_reg_1_10(.CP(n_62718), .D(n_21629), .CD(n_61496), .Q(ecx
		[10]));
	notech_mux2 i_8491(.S(\nbus_11330[0] ), .A(ecx[10]), .B(n_3848), .Z(n_21629
		));
	notech_reg regs_reg_1_11(.CP(n_62718), .D(n_21635), .CD(n_61494), .Q(ecx
		[11]));
	notech_mux2 i_8499(.S(\nbus_11330[0] ), .A(ecx[11]), .B(n_17141), .Z(n_21635
		));
	notech_reg regs_reg_1_12(.CP(n_62718), .D(n_21641), .CD(n_61494), .Q(ecx
		[12]));
	notech_mux2 i_8507(.S(\nbus_11330[0] ), .A(ecx[12]), .B(n_3841), .Z(n_21641
		));
	notech_reg regs_reg_1_13(.CP(n_62718), .D(n_21647), .CD(n_61496), .Q(ecx
		[13]));
	notech_mux2 i_8515(.S(\nbus_11330[0] ), .A(ecx[13]), .B(n_27027), .Z(n_21647
		));
	notech_reg regs_reg_1_14(.CP(n_62718), .D(n_21655), .CD(n_61496), .Q(ecx
		[14]));
	notech_mux2 i_8523(.S(\nbus_11330[0] ), .A(ecx[14]), .B(n_27028), .Z(n_21655
		));
	notech_reg regs_reg_1_15(.CP(n_62756), .D(n_21661), .CD(n_61496), .Q(ecx
		[15]));
	notech_mux2 i_8531(.S(\nbus_11330[0] ), .A(ecx[15]), .B(n_17165), .Z(n_21661
		));
	notech_reg regs_reg_1_16(.CP(n_62756), .D(n_21667), .CD(n_61496), .Q(ecx
		[16]));
	notech_mux2 i_8539(.S(\nbus_11330[16] ), .A(ecx[16]), .B(n_27011), .Z(n_21667
		));
	notech_reg regs_reg_1_17(.CP(n_62756), .D(n_21674), .CD(n_61496), .Q(ecx
		[17]));
	notech_mux2 i_8547(.S(\nbus_11330[16] ), .A(ecx[17]), .B(n_17177), .Z(n_21674
		));
	notech_nand3 i_28399(.A(n_60904), .B(n_62794), .C(\opa_12[13] ), .Z(n_31576
		));
	notech_reg regs_reg_1_18(.CP(n_62756), .D(n_21684), .CD(n_61494), .Q(ecx
		[18]));
	notech_mux2 i_8555(.S(\nbus_11330[16] ), .A(ecx[18]), .B(n_3862), .Z(n_21684
		));
	notech_nand2 i_28415(.A(n_62776), .B(opc_10[13]), .Z(n_31560));
	notech_reg regs_reg_1_19(.CP(n_62756), .D(n_21692), .CD(n_61494), .Q(ecx
		[19]));
	notech_mux2 i_8563(.S(\nbus_11330[16] ), .A(ecx[19]), .B(n_17189), .Z(n_21692
		));
	notech_or4 i_28435(.A(n_60969), .B(n_60958), .C(\opcode[1] ), .D(n_56239
		), .Z(n_31540));
	notech_reg regs_reg_1_20(.CP(n_62756), .D(n_21701), .CD(n_61494), .Q(ecx
		[20]));
	notech_mux2 i_8571(.S(\nbus_11330[16] ), .A(ecx[20]), .B(n_27578), .Z(n_21701
		));
	notech_nand3 i_28483(.A(n_60904), .B(n_62794), .C(\opa_12[11] ), .Z(n_31492
		));
	notech_reg regs_reg_1_21(.CP(n_62756), .D(n_21708), .CD(n_61494), .Q(ecx
		[21]));
	notech_mux2 i_8579(.S(\nbus_11330[16] ), .A(ecx[21]), .B(n_3838), .Z(n_21708
		));
	notech_nand2 i_28499(.A(n_62798), .B(opc_10[11]), .Z(n_31476));
	notech_reg regs_reg_1_22(.CP(n_62756), .D(n_21716), .CD(n_61494), .Q(ecx
		[22]));
	notech_mux2 i_8587(.S(\nbus_11330[16] ), .A(ecx[22]), .B(n_3859), .Z(n_21716
		));
	notech_or2 i_29381(.A(n_308891735), .B(n_56959), .Z(n_30594));
	notech_reg regs_reg_1_23(.CP(n_62756), .D(n_21723), .CD(n_61494), .Q(ecx
		[23]));
	notech_mux2 i_8595(.S(\nbus_11330[16] ), .A(ecx[23]), .B(n_27579), .Z(n_21723
		));
	notech_nao3 i_29406(.A(n_60378), .B(n_1476), .C(n_61151), .Z(n_30569));
	notech_reg regs_reg_1_24(.CP(n_62756), .D(n_21731), .CD(n_61494), .Q(ecx
		[24]));
	notech_mux2 i_8603(.S(\nbus_11330[16] ), .A(ecx[24]), .B(n_27581), .Z(n_21731
		));
	notech_or4 i_29407(.A(n_61171), .B(n_61160), .C(n_61151), .D(n_27305), .Z
		(n_30568));
	notech_reg regs_reg_1_25(.CP(n_62756), .D(n_21738), .CD(n_61494), .Q(ecx
		[25]));
	notech_mux2 i_8611(.S(\nbus_11330[16] ), .A(ecx[25]), .B(n_27582), .Z(n_21738
		));
	notech_or4 i_32833(.A(n_59382), .B(n_246791942), .C(n_32347), .D(n_59373
		), .Z(n_27142));
	notech_reg regs_reg_1_26(.CP(n_62756), .D(n_21746), .CD(n_61494), .Q(ecx
		[26]));
	notech_mux2 i_8619(.S(\nbus_11330[16] ), .A(ecx[26]), .B(n_237259453), .Z
		(n_21746));
	notech_reg regs_reg_1_27(.CP(n_62756), .D(n_21753), .CD(n_61494), .Q(ecx
		[27]));
	notech_mux2 i_8627(.S(\nbus_11330[16] ), .A(ecx[27]), .B(n_236059441), .Z
		(n_21753));
	notech_reg regs_reg_1_28(.CP(n_62756), .D(n_21761), .CD(n_61497), .Q(ecx
		[28]));
	notech_mux2 i_8635(.S(\nbus_11330[16] ), .A(ecx[28]), .B(n_1659), .Z(n_21761
		));
	notech_reg regs_reg_1_29(.CP(n_62756), .D(n_21768), .CD(n_61497), .Q(ecx
		[29]));
	notech_mux2 i_8643(.S(\nbus_11330[16] ), .A(ecx[29]), .B(n_234859429), .Z
		(n_21768));
	notech_reg regs_reg_1_30(.CP(n_62756), .D(n_21776), .CD(n_61497), .Q(ecx
		[30]));
	notech_mux2 i_8651(.S(\nbus_11330[16] ), .A(ecx[30]), .B(n_3856), .Z(n_21776
		));
	notech_or4 i_101540317(.A(n_58062), .B(n_2937), .C(n_56829), .D(n_32295)
		, .Z(n_2004));
	notech_reg regs_reg_1_31(.CP(n_62756), .D(n_21783), .CD(n_61497), .Q(ecx
		[31]));
	notech_mux2 i_8659(.S(\nbus_11330[16] ), .A(ecx[31]), .B(n_27233), .Z(n_21783
		));
	notech_reg_set divq_reg_0(.CP(n_62756), .D(n_21791), .SD(1'b1), .Q(divq[
		0]));
	notech_mux2 i_8667(.S(n_55535), .A(divq[0]), .B(n_13371), .Z(n_21791));
	notech_reg_set divq_reg_1(.CP(n_62718), .D(n_21798), .SD(1'b1), .Q(divq[
		1]));
	notech_mux2 i_8675(.S(n_55535), .A(divq[1]), .B(n_13376), .Z(n_21798));
	notech_nao3 i_100540323(.A(n_3879), .B(n_28552), .C(n_55581), .Z(n_2001)
		);
	notech_reg_set divq_reg_2(.CP(n_62756), .D(n_21806), .SD(1'b1), .Q(divq[
		2]));
	notech_mux2 i_8683(.S(n_55535), .A(divq[2]), .B(n_13381), .Z(n_21806));
	notech_or2 i_100440324(.A(n_4011), .B(n_56605), .Z(n_2000));
	notech_reg_set divq_reg_3(.CP(n_62720), .D(n_21813), .SD(1'b1), .Q(divq[
		3]));
	notech_mux2 i_8691(.S(n_55535), .A(divq[3]), .B(n_13386), .Z(n_21813));
	notech_and3 i_79240512(.A(n_303791786), .B(n_27346), .C(n_300891815), .Z
		(n_1999));
	notech_reg_set divq_reg_4(.CP(n_62720), .D(n_21821), .SD(1'b1), .Q(divq[
		4]));
	notech_mux2 i_8699(.S(n_55535), .A(divq[4]), .B(n_13391), .Z(n_21821));
	notech_or4 i_135541259(.A(n_57064), .B(n_57011), .C(n_54916), .D(n_1999)
		, .Z(n_27157));
	notech_reg_set divq_reg_5(.CP(n_62720), .D(n_21828), .SD(1'b1), .Q(divq[
		5]));
	notech_mux2 i_8707(.S(n_55535), .A(divq[5]), .B(n_13396), .Z(n_21828));
	notech_reg_set divq_reg_6(.CP(n_62720), .D(n_21838), .SD(1'b1), .Q(divq[
		6]));
	notech_mux2 i_8715(.S(n_55535), .A(divq[6]), .B(n_13401), .Z(n_21838));
	notech_and4 i_136343204(.A(n_38618568), .B(n_1995), .C(n_1918), .D(n_1915
		), .Z(n_1998));
	notech_reg_set divq_reg_7(.CP(n_62720), .D(n_21852), .SD(1'b1), .Q(divq[
		7]));
	notech_mux2 i_8723(.S(n_55535), .A(divq[7]), .B(n_13406), .Z(n_21852));
	notech_reg_set divq_reg_8(.CP(n_62720), .D(n_21859), .SD(1'b1), .Q(divq[
		8]));
	notech_mux2 i_8731(.S(n_55535), .A(divq[8]), .B(n_13411), .Z(n_21859));
	notech_reg_set divq_reg_9(.CP(n_62720), .D(n_21867), .SD(1'b1), .Q(divq[
		9]));
	notech_mux2 i_8739(.S(n_55535), .A(divq[9]), .B(n_13416), .Z(n_21867));
	notech_ao4 i_136143206(.A(n_60139), .B(n_27151), .C(n_83019012), .D(n_308791736
		), .Z(n_1995));
	notech_reg_set divq_reg_10(.CP(n_62720), .D(n_21874), .SD(1'b1), .Q(divq
		[10]));
	notech_mux2 i_8747(.S(n_55535), .A(divq[10]), .B(n_13421), .Z(n_21874)
		);
	notech_reg_set divq_reg_11(.CP(n_62720), .D(n_21882), .SD(1'b1), .Q(divq
		[11]));
	notech_mux2 i_8755(.S(n_55535), .A(divq[11]), .B(n_13426), .Z(n_21882)
		);
	notech_ao4 i_136443203(.A(n_96519147), .B(n_307891745), .C(n_314591678),
		 .D(n_56557), .Z(n_1992));
	notech_reg_set divq_reg_12(.CP(n_62720), .D(n_21889), .SD(1'b1), .Q(divq
		[12]));
	notech_mux2 i_8763(.S(n_55535), .A(divq[12]), .B(n_13431), .Z(n_21889)
		);
	notech_reg_set divq_reg_13(.CP(n_62720), .D(n_21897), .SD(1'b1), .Q(divq
		[13]));
	notech_mux2 i_8771(.S(n_55535), .A(divq[13]), .B(n_13436), .Z(n_21897)
		);
	notech_ao4 i_136543202(.A(n_29619), .B(n_187357098), .C(n_306791756), .D
		(n_1867), .Z(n_1990));
	notech_reg_set divq_reg_14(.CP(n_62720), .D(n_21904), .SD(1'b1), .Q(divq
		[14]));
	notech_mux2 i_8779(.S(n_55535), .A(divq[14]), .B(n_13441), .Z(n_21904)
		);
	notech_ao4 i_80744477(.A(n_61109), .B(n_1908), .C(n_314791676), .D(n_1988
		), .Z(n_38618568));
	notech_reg_set divq_reg_15(.CP(n_62720), .D(n_21912), .SD(1'b1), .Q(divq
		[15]));
	notech_mux2 i_8787(.S(n_55535), .A(divq[15]), .B(n_13446), .Z(n_21912)
		);
	notech_or4 i_168142907(.A(n_61136), .B(n_60207), .C(n_59708), .D(n_32380
		), .Z(n_1988));
	notech_reg_set divq_reg_16(.CP(n_62720), .D(n_21919), .SD(1'b1), .Q(divq
		[16]));
	notech_mux2 i_8796(.S(n_55537), .A(divq[16]), .B(n_13451), .Z(n_21919)
		);
	notech_nand2 i_3044497(.A(n_62776), .B(opc_10[31]), .Z(n_83019012));
	notech_reg_set divq_reg_17(.CP(n_62720), .D(n_21927), .SD(1'b1), .Q(divq
		[17]));
	notech_mux2 i_8804(.S(n_55537), .A(divq[17]), .B(n_13456), .Z(n_21927)
		);
	notech_reg_set divq_reg_18(.CP(n_62720), .D(n_21934), .SD(1'b1), .Q(divq
		[18]));
	notech_mux2 i_8812(.S(n_55537), .A(divq[18]), .B(n_13461), .Z(n_21934)
		);
	notech_reg_set divq_reg_19(.CP(n_62720), .D(n_21942), .SD(1'b1), .Q(divq
		[19]));
	notech_mux2 i_8820(.S(n_55537), .A(divq[19]), .B(n_13466), .Z(n_21942)
		);
	notech_ao4 i_211942471(.A(n_56666), .B(n_28256), .C(n_56653), .D(n_28221
		), .Z(n_1983));
	notech_reg_set divq_reg_20(.CP(n_62720), .D(n_21949), .SD(1'b1), .Q(divq
		[20]));
	notech_mux2 i_8828(.S(n_55537), .A(divq[20]), .B(n_13471), .Z(n_21949)
		);
	notech_ao4 i_212042470(.A(n_56916), .B(n_29617), .C(n_56636), .D(n_28288
		), .Z(n_1982));
	notech_reg_set divq_reg_21(.CP(n_62720), .D(n_21957), .SD(1'b1), .Q(divq
		[21]));
	notech_mux2 i_8836(.S(n_55537), .A(divq[21]), .B(n_13476), .Z(n_21957)
		);
	notech_and2 i_212442466(.A(n_197857105), .B(n_1977), .Z(n_1981));
	notech_reg_set divq_reg_22(.CP(n_62644), .D(n_21964), .SD(1'b1), .Q(divq
		[22]));
	notech_mux2 i_8844(.S(n_55537), .A(divq[22]), .B(n_13481), .Z(n_21964)
		);
	notech_ao4 i_212242468(.A(n_56527), .B(n_28321), .C(n_56502), .D(n_28386
		), .Z(n_197857105));
	notech_reg_set divq_reg_23(.CP(n_62644), .D(n_21972), .SD(1'b1), .Q(divq
		[23]));
	notech_mux2 i_8852(.S(n_55537), .A(divq[23]), .B(n_13486), .Z(n_21972)
		);
	notech_ao4 i_212342467(.A(n_56489), .B(n_28354), .C(n_56627), .D(n_28450
		), .Z(n_1977));
	notech_reg_set divq_reg_24(.CP(n_62644), .D(n_21979), .SD(1'b1), .Q(divq
		[24]));
	notech_mux2 i_8860(.S(n_55537), .A(divq[24]), .B(n_13491), .Z(n_21979)
		);
	notech_and4 i_213242458(.A(n_1974), .B(n_1973), .C(n_1971), .D(n_1970), 
		.Z(n_1976));
	notech_reg_set divq_reg_25(.CP(n_62644), .D(n_21987), .SD(1'b1), .Q(divq
		[25]));
	notech_mux2 i_8868(.S(n_55537), .A(divq[25]), .B(n_13496), .Z(n_21987)
		);
	notech_reg_set divq_reg_26(.CP(n_62644), .D(n_21995), .SD(1'b1), .Q(divq
		[26]));
	notech_mux2 i_8876(.S(n_55537), .A(divq[26]), .B(n_13501), .Z(n_21995)
		);
	notech_ao4 i_212642464(.A(n_56614), .B(n_28418), .C(n_56605), .D(n_28482
		), .Z(n_1974));
	notech_reg_set divq_reg_27(.CP(n_62644), .D(n_22005), .SD(1'b1), .Q(divq
		[27]));
	notech_mux2 i_8884(.S(n_55537), .A(divq[27]), .B(n_13506), .Z(n_22005)
		);
	notech_ao4 i_212742463(.A(n_56583), .B(n_28515), .C(n_56570), .D(n_28559
		), .Z(n_1973));
	notech_reg_set divq_reg_28(.CP(n_62644), .D(n_22011), .SD(1'b1), .Q(divq
		[28]));
	notech_mux2 i_8892(.S(n_55537), .A(divq[28]), .B(n_13511), .Z(n_22011)
		);
	notech_reg_set divq_reg_29(.CP(n_62644), .D(n_22018), .SD(1'b1), .Q(divq
		[29]));
	notech_mux2 i_8900(.S(n_55537), .A(divq[29]), .B(n_13516), .Z(n_22018)
		);
	notech_ao4 i_212942461(.A(n_56557), .B(n_27893), .C(n_56547), .D(n_28592
		), .Z(n_1971));
	notech_reg_set divq_reg_30(.CP(n_62644), .D(n_22025), .SD(1'b1), .Q(divq
		[30]));
	notech_mux2 i_8908(.S(n_55537), .A(divq[30]), .B(n_13521), .Z(n_22025)
		);
	notech_ao4 i_213042460(.A(n_56592), .B(n_28189), .C(n_56518), .D(n_29618
		), .Z(n_1970));
	notech_reg_set divq_reg_31(.CP(n_62644), .D(n_22034), .SD(1'b1), .Q(divq
		[31]));
	notech_mux2 i_8916(.S(n_55537), .A(divq[31]), .B(n_13526), .Z(n_22034)
		);
	notech_nand2 i_41544495(.A(n_62776), .B(opc[31]), .Z(n_96519147));
	notech_reg_set divq_reg_32(.CP(n_62568), .D(n_22042), .SD(1'b1), .Q(divq
		[32]));
	notech_mux2 i_8924(.S(n_55530), .A(divq[32]), .B(n_13531), .Z(n_22042)
		);
	notech_reg_set divq_reg_33(.CP(n_62644), .D(n_22048), .SD(1'b1), .Q(divq
		[33]));
	notech_mux2 i_8932(.S(n_55530), .A(divq[33]), .B(n_27583), .Z(n_22048)
		);
	notech_reg_set divq_reg_34(.CP(n_62650), .D(n_22055), .SD(1'b1), .Q(divq
		[34]));
	notech_mux2 i_8940(.S(n_55530), .A(divq[34]), .B(n_27584), .Z(n_22055)
		);
	notech_ao4 i_216042430(.A(n_56662), .B(n_28230), .C(n_56649), .D(n_28197
		), .Z(n_1967));
	notech_reg_set divq_reg_35(.CP(n_62570), .D(n_22061), .SD(1'b1), .Q(divq
		[35]));
	notech_mux2 i_8948(.S(n_55530), .A(divq[35]), .B(n_27585), .Z(n_22061)
		);
	notech_ao4 i_216142429(.A(n_56916), .B(n_29616), .C(n_56636), .D(n_28264
		), .Z(n_1966));
	notech_reg_set divq_reg_36(.CP(n_62570), .D(n_22067), .SD(1'b1), .Q(divq
		[36]));
	notech_mux2 i_8956(.S(n_55530), .A(divq[36]), .B(n_27586), .Z(n_22067)
		);
	notech_and2 i_216542425(.A(n_1964), .B(n_1963), .Z(n_1965));
	notech_reg_set divq_reg_37(.CP(n_62570), .D(n_22073), .SD(1'b1), .Q(divq
		[37]));
	notech_mux2 i_8964(.S(n_55530), .A(divq[37]), .B(n_27587), .Z(n_22073)
		);
	notech_ao4 i_216342427(.A(n_56527), .B(n_28296), .C(n_56498), .D(n_28362
		), .Z(n_1964));
	notech_reg_set divq_reg_38(.CP(n_62570), .D(n_22079), .SD(1'b1), .Q(divq
		[38]));
	notech_mux2 i_8972(.S(n_55530), .A(divq[38]), .B(n_27588), .Z(n_22079)
		);
	notech_ao4 i_216442426(.A(n_56485), .B(n_28329), .C(n_56627), .D(n_28426
		), .Z(n_1963));
	notech_reg_set divq_reg_39(.CP(n_62570), .D(n_22085), .SD(1'b1), .Q(divq
		[39]));
	notech_mux2 i_8980(.S(n_55530), .A(divq[39]), .B(n_27589), .Z(n_22085)
		);
	notech_and4 i_217342417(.A(n_1960), .B(n_1959), .C(n_1957), .D(n_1956), 
		.Z(n_196257103));
	notech_reg_set divq_reg_40(.CP(n_62570), .D(n_22091), .SD(1'b1), .Q(divq
		[40]));
	notech_mux2 i_8988(.S(n_55530), .A(divq[40]), .B(n_27590), .Z(n_22091)
		);
	notech_reg_set divq_reg_41(.CP(n_62570), .D(n_22097), .SD(1'b1), .Q(divq
		[41]));
	notech_mux2 i_8996(.S(n_55530), .A(divq[41]), .B(n_27591), .Z(n_22097)
		);
	notech_ao4 i_216742423(.A(n_56614), .B(n_28394), .C(n_56601), .D(n_28458
		), .Z(n_1960));
	notech_reg_set divq_reg_42(.CP(n_62570), .D(n_22103), .SD(1'b1), .Q(divq
		[42]));
	notech_mux2 i_9004(.S(n_55530), .A(divq[42]), .B(n_27592), .Z(n_22103)
		);
	notech_ao4 i_216842422(.A(n_56592), .B(n_28165), .C(n_56583), .D(n_28490
		), .Z(n_1959));
	notech_reg_set divq_reg_43(.CP(n_62570), .D(n_22109), .SD(1'b1), .Q(divq
		[43]));
	notech_mux2 i_9012(.S(n_55530), .A(divq[43]), .B(n_27593), .Z(n_22109)
		);
	notech_reg_set divq_reg_44(.CP(n_62570), .D(n_22115), .SD(1'b1), .Q(divq
		[44]));
	notech_mux2 i_9020(.S(n_55530), .A(divq[44]), .B(n_27594), .Z(n_22115)
		);
	notech_ao4 i_217042420(.A(n_56570), .B(n_28523), .C(n_56557), .D(n_27865
		), .Z(n_1957));
	notech_reg_set divq_reg_45(.CP(n_62652), .D(n_22121), .SD(1'b1), .Q(divq
		[45]));
	notech_mux2 i_9028(.S(n_55530), .A(divq[45]), .B(n_27595), .Z(n_22121)
		);
	notech_ao4 i_217142419(.A(n_56547), .B(n_28567), .C(n_56518), .D(n_29615
		), .Z(n_1956));
	notech_reg_set divq_reg_46(.CP(n_62652), .D(n_22127), .SD(1'b1), .Q(divq
		[46]));
	notech_mux2 i_9037(.S(n_55530), .A(divq[46]), .B(n_27596), .Z(n_22127)
		);
	notech_reg_set divq_reg_47(.CP(n_62652), .D(n_22133), .SD(1'b1), .Q(divq
		[47]));
	notech_mux2 i_9045(.S(n_55530), .A(divq[47]), .B(n_27597), .Z(n_22133)
		);
	notech_reg_set divq_reg_48(.CP(n_62652), .D(n_22139), .SD(1'b1), .Q(divq
		[48]));
	notech_mux2 i_9053(.S(n_55532), .A(divq[48]), .B(n_27598), .Z(n_22139)
		);
	notech_reg_set divq_reg_49(.CP(n_62652), .D(n_22145), .SD(1'b1), .Q(divq
		[49]));
	notech_mux2 i_9061(.S(n_55532), .A(divq[49]), .B(n_27599), .Z(n_22145)
		);
	notech_reg_set divq_reg_50(.CP(n_62652), .D(n_22151), .SD(1'b1), .Q(divq
		[50]));
	notech_mux2 i_9069(.S(n_55532), .A(divq[50]), .B(n_27600), .Z(n_22151)
		);
	notech_reg_set divq_reg_51(.CP(n_62652), .D(n_22157), .SD(1'b1), .Q(divq
		[51]));
	notech_mux2 i_9077(.S(n_55532), .A(divq[51]), .B(n_27602), .Z(n_22157)
		);
	notech_reg_set divq_reg_52(.CP(n_62652), .D(n_22163), .SD(1'b1), .Q(divq
		[52]));
	notech_mux2 i_9085(.S(n_55532), .A(divq[52]), .B(n_27603), .Z(n_22163)
		);
	notech_reg_set divq_reg_53(.CP(n_62652), .D(n_22169), .SD(1'b1), .Q(divq
		[53]));
	notech_mux2 i_9093(.S(n_55532), .A(divq[53]), .B(n_27605), .Z(n_22169)
		);
	notech_reg_set divq_reg_54(.CP(n_62652), .D(n_22175), .SD(1'b1), .Q(divq
		[54]));
	notech_mux2 i_9101(.S(n_55532), .A(divq[54]), .B(n_27606), .Z(n_22175)
		);
	notech_reg_set divq_reg_55(.CP(n_62652), .D(n_22181), .SD(1'b1), .Q(divq
		[55]));
	notech_mux2 i_9109(.S(n_55532), .A(divq[55]), .B(n_27607), .Z(n_22181)
		);
	notech_reg_set divq_reg_56(.CP(n_62652), .D(n_22187), .SD(1'b1), .Q(divq
		[56]));
	notech_mux2 i_9117(.S(n_55532), .A(divq[56]), .B(n_27608), .Z(n_22187)
		);
	notech_reg_set divq_reg_57(.CP(n_62652), .D(n_22193), .SD(1'b1), .Q(divq
		[57]));
	notech_mux2 i_9125(.S(n_55532), .A(divq[57]), .B(n_27609), .Z(n_22193)
		);
	notech_reg_set divq_reg_58(.CP(n_62652), .D(n_22199), .SD(1'b1), .Q(divq
		[58]));
	notech_mux2 i_9133(.S(n_55532), .A(divq[58]), .B(n_27610), .Z(n_22199)
		);
	notech_reg_set divq_reg_59(.CP(n_62652), .D(n_22205), .SD(1'b1), .Q(divq
		[59]));
	notech_mux2 i_9141(.S(n_55532), .A(divq[59]), .B(n_27611), .Z(n_22205)
		);
	notech_reg_set divq_reg_60(.CP(n_62652), .D(n_22211), .SD(1'b1), .Q(divq
		[60]));
	notech_mux2 i_9149(.S(n_55532), .A(divq[60]), .B(n_27613), .Z(n_22211)
		);
	notech_reg_set divq_reg_61(.CP(n_62652), .D(n_22218), .SD(1'b1), .Q(divq
		[61]));
	notech_mux2 i_9157(.S(n_55532), .A(divq[61]), .B(n_27614), .Z(n_22218)
		);
	notech_reg_set divq_reg_62(.CP(n_62652), .D(n_22225), .SD(1'b1), .Q(divq
		[62]));
	notech_mux2 i_9165(.S(n_55532), .A(divq[62]), .B(n_27615), .Z(n_22225)
		);
	notech_nand2 i_6144433(.A(n_62776), .B(opc_10[7]), .Z(n_31309));
	notech_reg_set divq_reg_63(.CP(n_62652), .D(n_22232), .SD(1'b1), .Q(divq
		[63]));
	notech_mux2 i_9173(.S(n_55532), .A(divq[63]), .B(n_101485291), .Z(n_22232
		));
	notech_nand2 i_4444450(.A(n_62776), .B(opc[7]), .Z(n_31307));
	notech_reg_set divr_reg_0(.CP(n_62724), .D(n_22240), .SD(1'b1), .Q(divr[
		0]));
	notech_mux2 i_9182(.S(n_55575), .A(divr[0]), .B(n_21670), .Z(n_22240));
	notech_reg_set divr_reg_1(.CP(n_62650), .D(n_22247), .SD(1'b1), .Q(divr[
		1]));
	notech_mux2 i_9190(.S(n_55575), .A(divr[1]), .B(n_21675), .Z(n_22247));
	notech_reg_set divr_reg_2(.CP(n_62724), .D(n_22254), .SD(1'b1), .Q(divr[
		2]));
	notech_mux2 i_9198(.S(n_55575), .A(divr[2]), .B(n_21680), .Z(n_22254));
	notech_reg_set divr_reg_3(.CP(n_62724), .D(n_22261), .SD(1'b1), .Q(divr[
		3]));
	notech_mux2 i_9206(.S(n_55575), .A(divr[3]), .B(n_21685), .Z(n_22261));
	notech_reg_set divr_reg_4(.CP(n_62724), .D(n_22268), .SD(1'b1), .Q(divr[
		4]));
	notech_mux2 i_9214(.S(n_55575), .A(divr[4]), .B(n_21690), .Z(n_22268));
	notech_reg_set divr_reg_5(.CP(n_62724), .D(n_22276), .SD(1'b1), .Q(divr[
		5]));
	notech_mux2 i_9222(.S(n_55575), .A(divr[5]), .B(n_21695), .Z(n_22276));
	notech_reg_set divr_reg_6(.CP(n_62724), .D(n_22283), .SD(1'b1), .Q(divr[
		6]));
	notech_mux2 i_9230(.S(n_55575), .A(divr[6]), .B(n_21700), .Z(n_22283));
	notech_reg_set divr_reg_7(.CP(n_62724), .D(n_22290), .SD(1'b1), .Q(divr[
		7]));
	notech_mux2 i_9238(.S(n_55575), .A(divr[7]), .B(n_21705), .Z(n_22290));
	notech_reg_set divr_reg_8(.CP(n_62724), .D(n_22297), .SD(1'b1), .Q(divr[
		8]));
	notech_mux2 i_9246(.S(n_55575), .A(divr[8]), .B(n_21710), .Z(n_22297));
	notech_reg_set divr_reg_9(.CP(n_62724), .D(n_22304), .SD(1'b1), .Q(divr[
		9]));
	notech_mux2 i_9254(.S(n_55575), .A(divr[9]), .B(n_21715), .Z(n_22304));
	notech_reg_set divr_reg_10(.CP(n_62724), .D(n_22314), .SD(1'b1), .Q(divr
		[10]));
	notech_mux2 i_9262(.S(n_55575), .A(divr[10]), .B(n_21720), .Z(n_22314)
		);
	notech_reg_set divr_reg_11(.CP(n_62724), .D(n_22321), .SD(1'b1), .Q(divr
		[11]));
	notech_mux2 i_9270(.S(n_55575), .A(divr[11]), .B(n_21725), .Z(n_22321)
		);
	notech_reg_set divr_reg_12(.CP(n_62724), .D(n_22330), .SD(1'b1), .Q(divr
		[12]));
	notech_mux2 i_9279(.S(n_55575), .A(divr[12]), .B(n_21730), .Z(n_22330)
		);
	notech_reg_set divr_reg_13(.CP(n_62724), .D(n_22337), .SD(1'b1), .Q(divr
		[13]));
	notech_mux2 i_9287(.S(n_55575), .A(divr[13]), .B(n_21735), .Z(n_22337)
		);
	notech_reg_set divr_reg_14(.CP(n_62724), .D(n_22344), .SD(1'b1), .Q(divr
		[14]));
	notech_mux2 i_9295(.S(n_55575), .A(divr[14]), .B(n_21740), .Z(n_22344)
		);
	notech_reg_set divr_reg_15(.CP(n_62724), .D(n_22351), .SD(1'b1), .Q(divr
		[15]));
	notech_mux2 i_9303(.S(n_55575), .A(divr[15]), .B(n_21745), .Z(n_22351)
		);
	notech_reg_set divr_reg_16(.CP(n_62724), .D(n_22358), .SD(1'b1), .Q(divr
		[16]));
	notech_mux2 i_9311(.S(n_55577), .A(divr[16]), .B(n_21750), .Z(n_22358)
		);
	notech_or2 i_26844228(.A(n_314791676), .B(n_187592028), .Z(n_1923));
	notech_reg_set divr_reg_17(.CP(n_62724), .D(n_22366), .SD(1'b1), .Q(divr
		[17]));
	notech_mux2 i_9319(.S(n_55577), .A(divr[17]), .B(n_21755), .Z(n_22366)
		);
	notech_reg_set divr_reg_18(.CP(n_62724), .D(n_22373), .SD(1'b1), .Q(divr
		[18]));
	notech_mux2 i_9327(.S(n_55577), .A(divr[18]), .B(n_21760), .Z(n_22373)
		);
	notech_reg_set divr_reg_19(.CP(n_62724), .D(n_22380), .SD(1'b1), .Q(divr
		[19]));
	notech_mux2 i_9335(.S(n_55577), .A(divr[19]), .B(n_21765), .Z(n_22380)
		);
	notech_reg_set divr_reg_20(.CP(n_62650), .D(n_22387), .SD(1'b1), .Q(divr
		[20]));
	notech_mux2 i_9343(.S(n_55577), .A(divr[20]), .B(n_21770), .Z(n_22387)
		);
	notech_reg_set divr_reg_21(.CP(n_62650), .D(n_22394), .SD(1'b1), .Q(divr
		[21]));
	notech_mux2 i_9351(.S(n_55577), .A(divr[21]), .B(n_21775), .Z(n_22394)
		);
	notech_or4 i_27344223(.A(n_61136), .B(n_60321), .C(n_60283), .D(n_28123)
		, .Z(n_1918));
	notech_reg_set divr_reg_22(.CP(n_62650), .D(n_22402), .SD(1'b1), .Q(divr
		[22]));
	notech_mux2 i_9359(.S(n_55577), .A(divr[22]), .B(n_21780), .Z(n_22402)
		);
	notech_reg_set divr_reg_23(.CP(n_62650), .D(n_22408), .SD(1'b1), .Q(divr
		[23]));
	notech_mux2 i_9367(.S(n_55577), .A(divr[23]), .B(n_21785), .Z(n_22408)
		);
	notech_reg_set divr_reg_24(.CP(n_62650), .D(n_22414), .SD(1'b1), .Q(divr
		[24]));
	notech_mux2 i_9375(.S(n_55577), .A(divr[24]), .B(n_21790), .Z(n_22414)
		);
	notech_nao3 i_27444222(.A(\regs_1_0[31] ), .B(n_60283), .C(n_59322), .Z(n_1915
		));
	notech_reg_set divr_reg_25(.CP(n_62650), .D(n_22420), .SD(1'b1), .Q(divr
		[25]));
	notech_mux2 i_9384(.S(n_55577), .A(divr[25]), .B(n_21795), .Z(n_22420)
		);
	notech_reg_set divr_reg_26(.CP(n_62650), .D(n_22426), .SD(1'b1), .Q(divr
		[26]));
	notech_mux2 i_9392(.S(n_55577), .A(divr[26]), .B(n_21800), .Z(n_22426)
		);
	notech_reg_set divr_reg_27(.CP(n_62650), .D(n_22432), .SD(1'b1), .Q(divr
		[27]));
	notech_mux2 i_9400(.S(n_55577), .A(divr[27]), .B(n_21805), .Z(n_22432)
		);
	notech_reg_set divr_reg_28(.CP(n_62650), .D(n_22438), .SD(1'b1), .Q(divr
		[28]));
	notech_mux2 i_9408(.S(n_55577), .A(divr[28]), .B(n_21810), .Z(n_22438)
		);
	notech_reg_set divr_reg_29(.CP(n_62650), .D(n_22444), .SD(1'b1), .Q(divr
		[29]));
	notech_mux2 i_9416(.S(n_55577), .A(divr[29]), .B(n_21815), .Z(n_22444)
		);
	notech_reg_set divr_reg_30(.CP(n_62570), .D(n_22452), .SD(1'b1), .Q(divr
		[30]));
	notech_mux2 i_9424(.S(n_55577), .A(divr[30]), .B(n_21820), .Z(n_22452)
		);
	notech_nand2 i_66643850(.A(n_313991684), .B(\regs_13_14[31] ), .Z(n_1909
		));
	notech_reg_set divr_reg_31(.CP(n_62570), .D(n_22458), .SD(1'b1), .Q(divr
		[31]));
	notech_mux2 i_9432(.S(n_55577), .A(divr[31]), .B(n_21825), .Z(n_22458)
		);
	notech_and2 i_16944327(.A(n_314691677), .B(n_1909), .Z(n_1908));
	notech_reg_set divr_reg_32(.CP(n_62654), .D(n_22464), .SD(1'b1), .Q(divr
		[32]));
	notech_mux2 i_9440(.S(n_55570), .A(divr[32]), .B(n_21830), .Z(n_22464)
		);
	notech_reg_set divr_reg_33(.CP(n_62572), .D(n_22470), .SD(1'b1), .Q(divr
		[33]));
	notech_mux2 i_9448(.S(n_55570), .A(divr[33]), .B(n_21835), .Z(n_22470)
		);
	notech_reg_set divr_reg_34(.CP(n_62572), .D(n_22476), .SD(1'b1), .Q(divr
		[34]));
	notech_mux2 i_9456(.S(n_55570), .A(divr[34]), .B(n_21840), .Z(n_22476)
		);
	notech_or4 i_27844218(.A(n_60854), .B(n_32614), .C(n_307691747), .D(n_24589
		), .Z(n_188857101));
	notech_reg_set divr_reg_35(.CP(n_62572), .D(n_22482), .SD(1'b1), .Q(divr
		[35]));
	notech_mux2 i_9464(.S(n_55570), .A(divr[35]), .B(n_21845), .Z(n_22482)
		);
	notech_or2 i_27744219(.A(n_307391750), .B(n_24589), .Z(n_188357100));
	notech_reg_set divr_reg_36(.CP(n_62572), .D(n_22488), .SD(1'b1), .Q(divr
		[36]));
	notech_mux2 i_9472(.S(n_55570), .A(divr[36]), .B(n_21850), .Z(n_22488)
		);
	notech_reg_set divr_reg_37(.CP(n_62572), .D(n_22494), .SD(1'b1), .Q(divr
		[37]));
	notech_mux2 i_9480(.S(n_55570), .A(divr[37]), .B(n_21855), .Z(n_22494)
		);
	notech_reg_set divr_reg_38(.CP(n_62572), .D(n_22500), .SD(1'b1), .Q(divr
		[38]));
	notech_mux2 i_9488(.S(n_55570), .A(divr[38]), .B(n_21860), .Z(n_22500)
		);
	notech_and2 i_16344333(.A(n_307591748), .B(n_188857101), .Z(n_187592028)
		);
	notech_reg_set divr_reg_39(.CP(n_62572), .D(n_22506), .SD(1'b1), .Q(divr
		[39]));
	notech_mux2 i_9496(.S(n_55570), .A(divr[39]), .B(n_21865), .Z(n_22506)
		);
	notech_and2 i_16244334(.A(n_307291751), .B(n_188357100), .Z(n_187357098)
		);
	notech_reg_set divr_reg_40(.CP(n_62572), .D(n_22512), .SD(1'b1), .Q(divr
		[40]));
	notech_mux2 i_9504(.S(n_55570), .A(divr[40]), .B(n_21870), .Z(n_22512)
		);
	notech_ao4 i_16144335(.A(n_24590), .B(n_57837), .C(n_59726), .D(n_307391750
		), .Z(n_1867));
	notech_reg_set divr_reg_41(.CP(n_62572), .D(n_22518), .SD(1'b1), .Q(divr
		[41]));
	notech_mux2 i_9512(.S(n_55570), .A(divr[41]), .B(n_21875), .Z(n_22518)
		);
	notech_or2 i_8244412(.A(n_308891735), .B(n_56983), .Z(n_30825));
	notech_reg_set divr_reg_42(.CP(n_62572), .D(n_22524), .SD(1'b1), .Q(divr
		[42]));
	notech_mux2 i_9520(.S(n_55570), .A(divr[42]), .B(n_21880), .Z(n_22524)
		);
	notech_reg_set divr_reg_43(.CP(n_62654), .D(n_22530), .SD(1'b1), .Q(divr
		[43]));
	notech_mux2 i_9528(.S(n_55570), .A(divr[43]), .B(n_21885), .Z(n_22530)
		);
	notech_ao4 i_215645627(.A(n_55735), .B(n_27746), .C(n_30803), .D(eval_flag
		), .Z(n_1865));
	notech_reg_set divr_reg_44(.CP(n_62654), .D(n_22536), .SD(1'b1), .Q(divr
		[44]));
	notech_mux2 i_9536(.S(n_55570), .A(divr[44]), .B(n_21890), .Z(n_22536)
		);
	notech_reg_set divr_reg_45(.CP(n_62654), .D(n_22542), .SD(1'b1), .Q(divr
		[45]));
	notech_mux2 i_9545(.S(n_55570), .A(divr[45]), .B(n_21895), .Z(n_22542)
		);
	notech_reg_set divr_reg_46(.CP(n_62654), .D(n_22548), .SD(1'b1), .Q(divr
		[46]));
	notech_mux2 i_9553(.S(n_55570), .A(divr[46]), .B(n_21900), .Z(n_22548)
		);
	notech_reg_set divr_reg_47(.CP(n_62654), .D(n_22554), .SD(1'b1), .Q(divr
		[47]));
	notech_mux2 i_9561(.S(n_55570), .A(divr[47]), .B(n_21905), .Z(n_22554)
		);
	notech_reg_set divr_reg_48(.CP(n_62654), .D(n_22560), .SD(1'b1), .Q(divr
		[48]));
	notech_mux2 i_9569(.S(n_55572), .A(divr[48]), .B(n_21910), .Z(n_22560)
		);
	notech_ao4 i_5847641(.A(n_306291761), .B(n_306391760), .C(n_27761), .D(n_304591778
		), .Z(n_104722311));
	notech_reg_set divr_reg_49(.CP(n_62654), .D(n_22566), .SD(1'b1), .Q(divr
		[49]));
	notech_mux2 i_9577(.S(n_55572), .A(divr[49]), .B(n_21915), .Z(n_22566)
		);
	notech_or2 i_115846579(.A(n_312191702), .B(n_26611), .Z(n_1857));
	notech_reg_set divr_reg_50(.CP(n_62654), .D(n_22574), .SD(1'b1), .Q(divr
		[50]));
	notech_mux2 i_9585(.S(n_55572), .A(divr[50]), .B(n_21920), .Z(n_22574)
		);
	notech_reg_set divr_reg_51(.CP(n_62654), .D(n_22581), .SD(1'b1), .Q(divr
		[51]));
	notech_mux2 i_9593(.S(n_55572), .A(divr[51]), .B(n_21925), .Z(n_22581)
		);
	notech_reg_set divr_reg_52(.CP(n_62654), .D(n_22589), .SD(1'b1), .Q(divr
		[52]));
	notech_mux2 i_9601(.S(n_55572), .A(divr[52]), .B(n_21930), .Z(n_22589)
		);
	notech_reg_set divr_reg_53(.CP(n_62654), .D(n_22598), .SD(1'b1), .Q(divr
		[53]));
	notech_mux2 i_9609(.S(n_55572), .A(divr[53]), .B(n_21935), .Z(n_22598)
		);
	notech_reg_set divr_reg_54(.CP(n_62654), .D(n_22604), .SD(1'b1), .Q(divr
		[54]));
	notech_mux2 i_9617(.S(n_55572), .A(divr[54]), .B(n_21940), .Z(n_22604)
		);
	notech_reg_set divr_reg_55(.CP(n_62654), .D(n_22610), .SD(1'b1), .Q(divr
		[55]));
	notech_mux2 i_9625(.S(n_55572), .A(divr[55]), .B(n_21945), .Z(n_22610)
		);
	notech_reg_set divr_reg_56(.CP(n_62654), .D(n_22616), .SD(1'b1), .Q(divr
		[56]));
	notech_mux2 i_9633(.S(n_55572), .A(divr[56]), .B(n_21950), .Z(n_22616)
		);
	notech_reg_set divr_reg_57(.CP(n_62654), .D(n_22622), .SD(1'b1), .Q(divr
		[57]));
	notech_mux2 i_9641(.S(n_55572), .A(divr[57]), .B(n_21955), .Z(n_22622)
		);
	notech_and3 i_115046587(.A(n_28544), .B(n_28543), .C(n_28545), .Z(n_184992034
		));
	notech_reg_set divr_reg_58(.CP(n_62654), .D(n_22628), .SD(1'b1), .Q(divr
		[58]));
	notech_mux2 i_9649(.S(n_55572), .A(divr[58]), .B(n_21960), .Z(n_22628)
		);
	notech_and3 i_3347666(.A(n_300891815), .B(n_27346), .C(n_27349), .Z(n_184892035
		));
	notech_reg_set divr_reg_59(.CP(n_62654), .D(n_22634), .SD(1'b1), .Q(divr
		[59]));
	notech_mux2 i_9657(.S(n_55572), .A(divr[59]), .B(n_21965), .Z(n_22634)
		);
	notech_and4 i_3247667(.A(n_56843), .B(n_1441), .C(n_55735), .D(n_305191772
		), .Z(n_184792036));
	notech_reg_set divr_reg_60(.CP(n_62654), .D(n_22640), .SD(1'b1), .Q(divr
		[60]));
	notech_mux2 i_9665(.S(n_55572), .A(divr[60]), .B(n_21970), .Z(n_22640)
		);
	notech_nand2 i_12544(.A(n_304491779), .B(n_32616), .Z(n_184692037));
	notech_reg_set divr_reg_61(.CP(n_62572), .D(n_22646), .SD(1'b1), .Q(divr
		[61]));
	notech_mux2 i_9673(.S(n_55572), .A(divr[61]), .B(n_21975), .Z(n_22646)
		);
	notech_reg_set divr_reg_62(.CP(n_62572), .D(n_22652), .SD(1'b1), .Q(divr
		[62]));
	notech_mux2 i_9681(.S(n_55572), .A(divr[62]), .B(n_21980), .Z(n_22652)
		);
	notech_reg_set divr_reg_63(.CP(n_62574), .D(n_22658), .SD(1'b1), .Q(divr
		[63]));
	notech_mux2 i_9689(.S(n_55572), .A(divr[63]), .B(n_21985), .Z(n_22658)
		);
	notech_or4 i_103949654(.A(n_32343), .B(n_32342), .C(n_314891675), .D(n_184192042
		), .Z(n_184392040));
	notech_reg sign_div_reg(.CP(n_62574), .D(n_22664), .CD(n_61497), .Q(sign_div
		));
	notech_mux2 i_9697(.S(n_328190779), .A(n_26990), .B(sign_div), .Z(n_22664
		));
	notech_nao3 i_103649657(.A(n_57992), .B(n_27221), .C(n_311991704), .Z(n_184292041
		));
	notech_reg_set opc_reg_0(.CP(n_62574), .D(n_22672), .SD(1'b1), .Q(opc[0]
		));
	notech_mux2 i_9705(.S(n_27622), .A(opc[0]), .B(n_27619), .Z(n_22672));
	notech_and3 i_1050639(.A(n_56843), .B(n_2004), .C(n_24994), .Z(n_184192042
		));
	notech_reg_set opc_reg_1(.CP(n_62574), .D(n_22678), .SD(1'b1), .Q(opc[1]
		));
	notech_mux2 i_9713(.S(n_27622), .A(opc[1]), .B(n_27620), .Z(n_22678));
	notech_reg_set opc_reg_2(.CP(n_62574), .D(n_22684), .SD(1'b1), .Q(opc[2]
		));
	notech_mux2 i_9721(.S(n_27622), .A(opc[2]), .B(n_15031), .Z(n_22684));
	notech_reg_set opc_reg_3(.CP(n_62574), .D(n_22690), .SD(1'b1), .Q(opc[3]
		));
	notech_mux2 i_9729(.S(n_27622), .A(opc[3]), .B(n_27621), .Z(n_22690));
	notech_reg_set opc_reg_4(.CP(n_62574), .D(n_22696), .SD(1'b1), .Q(opc[4]
		));
	notech_mux2 i_9737(.S(n_27622), .A(opc[4]), .B(n_15041), .Z(n_22696));
	notech_reg_set opc_reg_5(.CP(n_62574), .D(n_22702), .SD(1'b1), .Q(opc[5]
		));
	notech_mux2 i_9745(.S(n_27623), .A(opc[5]), .B(n_15046), .Z(n_22702));
	notech_ao4 i_170452272(.A(n_174292094), .B(n_311491709), .C(n_174992087)
		, .D(n_311391710), .Z(n_1836));
	notech_reg_set opc_reg_6(.CP(n_62574), .D(n_22708), .SD(1'b1), .Q(opc[6]
		));
	notech_mux2 i_9753(.S(n_27623), .A(opc[6]), .B(n_15051), .Z(n_22708));
	notech_reg_set opc_reg_7(.CP(n_62574), .D(n_22714), .SD(1'b1), .Q(opc[7]
		));
	notech_mux2 i_9761(.S(n_27623), .A(opc[7]), .B(n_15056), .Z(n_22714));
	notech_and4 i_170252274(.A(n_1832), .B(n_1831), .C(n_1829), .D(n_1667), 
		.Z(n_1834));
	notech_reg_set opc_reg_8(.CP(n_62574), .D(n_22721), .SD(1'b1), .Q(opc[8]
		));
	notech_mux2 i_9769(.S(n_138582386), .A(n_15061), .B(opc[8]), .Z(n_22721)
		);
	notech_reg_set opc_reg_9(.CP(n_62574), .D(n_22728), .SD(1'b1), .Q(opc[9]
		));
	notech_mux2 i_9777(.S(n_138582386), .A(n_15066), .B(opc[9]), .Z(n_22728)
		);
	notech_ao4 i_169952277(.A(n_26696), .B(n_29660), .C(n_133728614), .D(n_151428791
		), .Z(n_1832));
	notech_reg_set opc_reg_10(.CP(n_62574), .D(n_22736), .SD(1'b1), .Q(opc[
		10]));
	notech_mux2 i_9785(.S(n_138582386), .A(n_15071), .B(opc[10]), .Z(n_22736
		));
	notech_ao4 i_169852278(.A(n_311191712), .B(n_55947), .C(n_311091713), .D
		(n_57783), .Z(n_1831));
	notech_reg_set opc_reg_11(.CP(n_62574), .D(n_22743), .SD(1'b1), .Q(opc[
		11]));
	notech_mux2 i_9793(.S(n_138582386), .A(n_15076), .B(opc[11]), .Z(n_22743
		));
	notech_reg_set opc_reg_12(.CP(n_62574), .D(n_22751), .SD(1'b1), .Q(opc[
		12]));
	notech_mux2 i_9801(.S(n_138582386), .A(n_15081), .B(opc[12]), .Z(n_22751
		));
	notech_ao4 i_169752279(.A(n_59124), .B(nbus_11295[26]), .C(n_54638), .D(n_28958
		), .Z(n_1829));
	notech_reg_set opc_reg_13(.CP(n_62574), .D(n_22758), .SD(1'b1), .Q(opc[
		13]));
	notech_mux2 i_9809(.S(n_138582386), .A(n_15086), .B(opc[13]), .Z(n_22758
		));
	notech_reg_set opc_reg_14(.CP(n_62574), .D(n_22766), .SD(1'b1), .Q(opc[
		14]));
	notech_mux2 i_9817(.S(n_138582386), .A(n_15091), .B(opc[14]), .Z(n_22766
		));
	notech_reg_set opc_reg_15(.CP(n_62574), .D(n_22773), .SD(1'b1), .Q(opc[
		15]));
	notech_mux2 i_9825(.S(n_138582386), .A(n_15096), .B(opc[15]), .Z(n_22773
		));
	notech_and4 i_159952377(.A(n_1824), .B(n_1823), .C(n_1821), .D(n_1820), 
		.Z(n_1826));
	notech_reg_set opc_reg_16(.CP(n_62574), .D(n_22781), .SD(1'b1), .Q(opc[
		16]));
	notech_mux2 i_9833(.S(n_27640), .A(opc[16]), .B(n_27624), .Z(n_22781));
	notech_reg_set opc_reg_17(.CP(n_62524), .D(n_22788), .SD(1'b1), .Q(opc[
		17]));
	notech_mux2 i_9842(.S(n_27640), .A(opc[17]), .B(n_27625), .Z(n_22788));
	notech_ao4 i_159652380(.A(n_60139), .B(n_27150), .C(n_308591738), .D(n_28013
		), .Z(n_1824));
	notech_reg_set opc_reg_18(.CP(n_62524), .D(n_22796), .SD(1'b1), .Q(opc[
		18]));
	notech_mux2 i_9851(.S(n_27640), .A(opc[18]), .B(n_27626), .Z(n_22796));
	notech_ao4 i_159552381(.A(n_59095), .B(n_28117), .C(n_150628783), .D(n_29662
		), .Z(n_1823));
	notech_reg_set opc_reg_19(.CP(n_62524), .D(n_22803), .SD(1'b1), .Q(opc[
		19]));
	notech_mux2 i_9860(.S(n_27640), .A(opc[19]), .B(n_27627), .Z(n_22803));
	notech_reg_set opc_reg_20(.CP(n_62524), .D(n_22811), .SD(1'b1), .Q(opc[
		20]));
	notech_mux2 i_9868(.S(n_27640), .A(opc[20]), .B(n_27628), .Z(n_22811));
	notech_ao4 i_159452382(.A(n_130528582), .B(n_150728784), .C(n_150528782)
		, .D(n_55974), .Z(n_1821));
	notech_reg_set opc_reg_21(.CP(n_62524), .D(n_22818), .SD(1'b1), .Q(opc[
		21]));
	notech_mux2 i_9876(.S(n_27640), .A(opc[21]), .B(n_27629), .Z(n_22818));
	notech_ao4 i_159352383(.A(n_150428781), .B(n_57802), .C(n_26648), .D(n_29605
		), .Z(n_1820));
	notech_reg_set opc_reg_22(.CP(n_62524), .D(n_22826), .SD(1'b1), .Q(opc[
		22]));
	notech_mux2 i_9884(.S(n_27640), .A(opc[22]), .B(n_27630), .Z(n_22826));
	notech_reg_set opc_reg_23(.CP(n_62524), .D(n_22833), .SD(1'b1), .Q(opc[
		23]));
	notech_mux2 i_9892(.S(n_27640), .A(opc[23]), .B(n_27631), .Z(n_22833));
	notech_reg_set opc_reg_24(.CP(n_62524), .D(n_22841), .SD(1'b1), .Q(opc[
		24]));
	notech_mux2 i_9900(.S(n_27640), .A(opc[24]), .B(n_27632), .Z(n_22841));
	notech_and4 i_150152475(.A(n_1814), .B(n_1813), .C(n_1812), .D(n_3883), 
		.Z(n_1817));
	notech_reg_set opc_reg_25(.CP(n_62524), .D(n_22848), .SD(1'b1), .Q(opc[
		25]));
	notech_mux2 i_9908(.S(n_27640), .A(opc[25]), .B(n_27633), .Z(n_22848));
	notech_reg_set opc_reg_26(.CP(n_62524), .D(n_22856), .SD(1'b1), .Q(opc[
		26]));
	notech_mux2 i_9916(.S(n_27640), .A(opc[26]), .B(n_27634), .Z(n_22856));
	notech_reg_set opc_reg_27(.CP(n_62524), .D(n_22863), .SD(1'b1), .Q(opc[
		27]));
	notech_mux2 i_9924(.S(n_27640), .A(opc[27]), .B(n_27635), .Z(n_22863));
	notech_ao4 i_149752479(.A(n_128228559), .B(n_149128768), .C(n_149428771)
		, .D(n_55956), .Z(n_1814));
	notech_reg_set opc_reg_28(.CP(n_62524), .D(n_22871), .SD(1'b1), .Q(opc[
		28]));
	notech_mux2 i_9932(.S(n_27640), .A(opc[28]), .B(n_27636), .Z(n_22871));
	notech_ao4 i_149652480(.A(n_149328770), .B(n_57815), .C(n_54638), .D(n_28984
		), .Z(n_1813));
	notech_reg_set opc_reg_29(.CP(n_62740), .D(n_22878), .SD(1'b1), .Q(opc[
		29]));
	notech_mux2 i_9940(.S(n_27640), .A(opc[29]), .B(n_27637), .Z(n_22878));
	notech_ao4 i_149852478(.A(n_310691717), .B(n_28014), .C(n_149228769), .D
		(n_29659), .Z(n_1812));
	notech_reg_set opc_reg_30(.CP(n_62448), .D(n_22884), .SD(1'b1), .Q(opc[
		30]));
	notech_mux2 i_9948(.S(n_27640), .A(opc[30]), .B(n_27638), .Z(n_22884));
	notech_reg_set opc_reg_31(.CP(n_62448), .D(n_22890), .SD(1'b1), .Q(opc[
		31]));
	notech_mux2 i_9956(.S(n_27640), .A(opc[31]), .B(n_27639), .Z(n_22890));
	notech_reg nZF_reg(.CP(n_62448), .D(n_22896), .CD(n_61498), .Q(nZF));
	notech_mux2 i_9964(.S(n_21998), .A(nZF), .B(n_22001), .Z(n_22896));
	notech_nand3 i_141052560(.A(n_1802), .B(n_180192047), .C(n_1808), .Z(n_1809
		));
	notech_reg regs_reg_0_0(.CP(n_62448), .D(n_22902), .CD(n_61498), .Q(regs_0
		[0]));
	notech_mux2 i_9972(.S(n_27652), .A(regs_0[0]), .B(n_27642), .Z(n_22902)
		);
	notech_and3 i_140952561(.A(n_1806), .B(n_1805), .C(n_1804), .Z(n_1808)
		);
	notech_reg regs_reg_0_1(.CP(n_62448), .D(n_22908), .CD(n_61497), .Q(regs_0
		[1]));
	notech_mux2 i_9980(.S(n_27652), .A(regs_0[1]), .B(n_16712), .Z(n_22908)
		);
	notech_reg regs_reg_0_2(.CP(n_62448), .D(n_22914), .CD(n_61497), .Q(regs_0
		[2]));
	notech_mux2 i_9988(.S(n_27652), .A(regs_0[2]), .B(n_27643), .Z(n_22914)
		);
	notech_ao4 i_140352567(.A(n_146928746), .B(\nbus_11365[26] ), .C(n_54865
		), .D(n_29604), .Z(n_1806));
	notech_reg regs_reg_0_3(.CP(n_62448), .D(n_22920), .CD(n_61497), .Q(regs_0
		[3]));
	notech_mux2 i_9996(.S(n_27652), .A(regs_0[3]), .B(n_16724), .Z(n_22920)
		);
	notech_ao4 i_140252568(.A(n_54883), .B(n_28619), .C(n_54894), .D(n_27477
		), .Z(n_1805));
	notech_reg regs_reg_0_4(.CP(n_62448), .D(n_22926), .CD(n_61496), .Q(regs_0
		[4]));
	notech_mux2 i_10004(.S(n_27652), .A(regs_0[4]), .B(n_27644), .Z(n_22926)
		);
	notech_ao4 i_140652564(.A(n_60144), .B(n_27184), .C(n_310391720), .D(n_28011
		), .Z(n_1804));
	notech_reg regs_reg_0_5(.CP(n_62448), .D(n_22932), .CD(n_61496), .Q(regs_0
		[5]));
	notech_mux2 i_10012(.S(n_27652), .A(regs_0[5]), .B(n_16736), .Z(n_22932)
		);
	notech_reg regs_reg_0_6(.CP(n_62544), .D(n_22938), .CD(n_61496), .Q(regs_0
		[6]));
	notech_mux2 i_10020(.S(n_27652), .A(regs_0[6]), .B(n_16742), .Z(n_22938)
		);
	notech_ao4 i_140552565(.A(n_54874), .B(n_28115), .C(n_147128748), .D(n_29660
		), .Z(n_1802));
	notech_reg regs_reg_0_7(.CP(n_62544), .D(n_22944), .CD(n_61496), .Q(regs_0
		[7]));
	notech_mux2 i_10028(.S(n_27652), .A(regs_0[7]), .B(n_27645), .Z(n_22944)
		);
	notech_ao4 i_140452566(.A(n_133728614), .B(n_147228749), .C(n_147028747)
		, .D(\nbus_11358[26] ), .Z(n_180192047));
	notech_reg regs_reg_0_8(.CP(n_62544), .D(n_22950), .CD(n_61496), .Q(regs_0
		[8]));
	notech_mux2 i_10036(.S(n_27652), .A(regs_0[8]), .B(n_16754), .Z(n_22950)
		);
	notech_reg regs_reg_0_9(.CP(n_62544), .D(n_22956), .CD(n_61497), .Q(regs_0
		[9]));
	notech_mux2 i_10044(.S(n_27652), .A(regs_0[9]), .B(n_27646), .Z(n_22956)
		);
	notech_reg regs_reg_0_10(.CP(n_62544), .D(n_22962), .CD(n_61497), .Q(regs_0
		[10]));
	notech_mux2 i_10052(.S(n_27652), .A(regs_0[10]), .B(n_27647), .Z(n_22962
		));
	notech_nand3 i_124452724(.A(n_179292055), .B(n_179192056), .C(n_179792050
		), .Z(n_179892049));
	notech_reg regs_reg_0_11(.CP(n_62544), .D(n_22968), .CD(n_61497), .Q(regs_0
		[11]));
	notech_mux2 i_10060(.S(n_27652), .A(regs_0[11]), .B(n_27648), .Z(n_22968
		));
	notech_and3 i_124352725(.A(n_179592052), .B(n_179492053), .C(n_1620), .Z
		(n_179792050));
	notech_reg regs_reg_0_12(.CP(n_62544), .D(n_22974), .CD(n_61497), .Q(regs_0
		[12]));
	notech_mux2 i_10068(.S(n_27652), .A(regs_0[12]), .B(n_16778), .Z(n_22974
		));
	notech_reg regs_reg_0_13(.CP(n_62544), .D(n_22980), .CD(n_61474), .Q(regs_0
		[13]));
	notech_mux2 i_10076(.S(n_27652), .A(regs_0[13]), .B(n_16784), .Z(n_22980
		));
	notech_ao4 i_123752731(.A(n_54658), .B(n_29602), .C(n_27334), .D(n_29600
		), .Z(n_179592052));
	notech_reg regs_reg_0_14(.CP(n_62544), .D(n_22986), .CD(n_61474), .Q(regs_0
		[14]));
	notech_mux2 i_10084(.S(n_27652), .A(regs_0[14]), .B(n_27649), .Z(n_22986
		));
	notech_ao4 i_124052728(.A(n_27319), .B(n_28011), .C(n_59322), .D(n_28115
		), .Z(n_179492053));
	notech_reg regs_reg_0_15(.CP(n_62544), .D(n_22992), .CD(n_61474), .Q(regs_0
		[15]));
	notech_mux2 i_10092(.S(n_27652), .A(regs_0[15]), .B(n_27650), .Z(n_22992
		));
	notech_reg regs_reg_0_16(.CP(n_62544), .D(n_22999), .CD(n_61474), .Q(regs_0
		[16]));
	notech_mux2 i_10100(.S(n_54983), .A(regs_0[16]), .B(n_16802), .Z(n_22999
		));
	notech_ao4 i_123952729(.A(n_145028727), .B(n_29660), .C(n_133728614), .D
		(n_145128728), .Z(n_179292055));
	notech_reg regs_reg_0_17(.CP(n_62544), .D(n_23008), .CD(n_61474), .Q(regs_0
		[17]));
	notech_mux2 i_10108(.S(n_54983), .A(regs_0[17]), .B(n_16808), .Z(n_23008
		));
	notech_ao4 i_123852730(.A(n_144928726), .B(n_55947), .C(n_144828725), .D
		(n_57783), .Z(n_179192056));
	notech_reg regs_reg_0_18(.CP(n_62544), .D(n_23015), .CD(n_61474), .Q(regs_0
		[18]));
	notech_mux2 i_10116(.S(n_54983), .A(regs_0[18]), .B(n_16814), .Z(n_23015
		));
	notech_reg regs_reg_0_19(.CP(n_62544), .D(n_23022), .CD(n_61474), .Q(regs_0
		[19]));
	notech_mux2 i_10124(.S(n_54983), .A(regs_0[19]), .B(n_16820), .Z(n_23022
		));
	notech_reg regs_reg_0_20(.CP(n_62544), .D(n_23030), .CD(n_61474), .Q(regs_0
		[20]));
	notech_mux2 i_10132(.S(n_54983), .A(regs_0[20]), .B(n_16826), .Z(n_23030
		));
	notech_nand3 i_122152747(.A(n_178692061), .B(n_178592062), .C(n_178492063
		), .Z(n_178892059));
	notech_reg regs_reg_0_21(.CP(n_62544), .D(n_23038), .CD(n_61474), .Q(regs_0
		[21]));
	notech_mux2 i_10140(.S(n_54983), .A(regs_0[21]), .B(n_16832), .Z(n_23038
		));
	notech_reg regs_reg_0_22(.CP(n_62544), .D(n_23046), .CD(n_61472), .Q(regs_0
		[22]));
	notech_mux2 i_10148(.S(n_54983), .A(regs_0[22]), .B(n_16838), .Z(n_23046
		));
	notech_ao4 i_121552753(.A(n_144828725), .B(n_57792), .C(n_27329), .D(n_310091723
		), .Z(n_178692061));
	notech_reg regs_reg_0_23(.CP(n_62544), .D(n_23054), .CD(n_61472), .Q(regs_0
		[23]));
	notech_mux2 i_10156(.S(n_54983), .A(regs_0[23]), .B(n_16844), .Z(n_23054
		));
	notech_ao4 i_121452754(.A(n_54658), .B(n_29598), .C(n_27334), .D(n_29597
		), .Z(n_178592062));
	notech_reg regs_reg_0_24(.CP(n_62544), .D(n_23061), .CD(n_61472), .Q(regs_0
		[24]));
	notech_mux2 i_10164(.S(n_54983), .A(regs_0[24]), .B(n_16850), .Z(n_23061
		));
	notech_ao4 i_121852750(.A(n_60144), .B(n_27215), .C(n_27319), .D(n_28012
		), .Z(n_178492063));
	notech_reg regs_reg_0_25(.CP(n_62542), .D(n_23067), .CD(n_61472), .Q(regs_0
		[25]));
	notech_mux2 i_10172(.S(n_54983), .A(regs_0[25]), .B(n_16856), .Z(n_23067
		));
	notech_nand2 i_122052748(.A(n_178292065), .B(n_178192066), .Z(n_178392064
		));
	notech_reg regs_reg_0_26(.CP(n_62542), .D(n_23073), .CD(n_61472), .Q(regs_0
		[26]));
	notech_mux2 i_10180(.S(n_54983), .A(regs_0[26]), .B(n_27268), .Z(n_23073
		));
	notech_ao4 i_121752751(.A(n_59326), .B(n_28116), .C(n_145028727), .D(n_29661
		), .Z(n_178292065));
	notech_reg regs_reg_0_27(.CP(n_62614), .D(n_23079), .CD(n_61472), .Q(regs_0
		[27]));
	notech_mux2 i_10188(.S(n_54983), .A(regs_0[27]), .B(n_16868), .Z(n_23079
		));
	notech_ao4 i_121652752(.A(n_131228589), .B(n_145128728), .C(n_144928726)
		, .D(n_55938), .Z(n_178192066));
	notech_reg regs_reg_0_28(.CP(n_62614), .D(n_23086), .CD(n_61472), .Q(regs_0
		[28]));
	notech_mux2 i_10196(.S(n_54983), .A(regs_0[28]), .B(n_27019), .Z(n_23086
		));
	notech_reg regs_reg_0_29(.CP(n_62614), .D(n_23093), .CD(n_61472), .Q(regs_0
		[29]));
	notech_mux2 i_10204(.S(n_54983), .A(regs_0[29]), .B(n_27651), .Z(n_23093
		));
	notech_ao4 i_115252816(.A(n_1583), .B(n_56190), .C(n_3885), .D(n_3997), 
		.Z(n_177992068));
	notech_reg regs_reg_0_30(.CP(n_62614), .D(n_23100), .CD(n_61472), .Q(regs_0
		[30]));
	notech_mux2 i_10212(.S(n_54983), .A(regs_0[30]), .B(n_16886), .Z(n_23100
		));
	notech_and4 i_115352815(.A(n_177592072), .B(n_1592), .C(n_1593), .D(n_1596
		), .Z(n_177892069));
	notech_reg regs_reg_0_31(.CP(n_62614), .D(n_23107), .CD(n_61472), .Q(regs_0
		[31]));
	notech_mux2 i_10220(.S(n_54983), .A(regs_0[31]), .B(n_16892), .Z(n_23107
		));
	notech_reg cr1_reg_0(.CP(n_62614), .D(n_23114), .CD(n_61475), .Q(nbus_14521
		[0]));
	notech_mux2 i_10228(.S(n_328084271), .A(opa[0]), .B(nbus_14521[0]), .Z(n_23114
		));
	notech_reg cr1_reg_1(.CP(n_62614), .D(n_23121), .CD(n_61475), .Q(nbus_14521
		[1]));
	notech_mux2 i_10236(.S(n_328084271), .A(opa[1]), .B(nbus_14521[1]), .Z(n_23121
		));
	notech_and4 i_114852819(.A(n_1771), .B(n_177092073), .C(n_1773), .D(n_1591
		), .Z(n_177592072));
	notech_reg cr1_reg_2(.CP(n_62614), .D(n_23128), .CD(n_61475), .Q(nbus_14521
		[2]));
	notech_mux2 i_10244(.S(n_328084271), .A(opa[2]), .B(nbus_14521[2]), .Z(n_23128
		));
	notech_reg cr1_reg_3(.CP(n_62614), .D(n_23135), .CD(n_61475), .Q(nbus_14521
		[3]));
	notech_mux2 i_10252(.S(n_328084271), .A(opa[3]), .B(nbus_14521[3]), .Z(n_23135
		));
	notech_ao4 i_114652821(.A(n_31492), .B(n_27604), .C(n_56518), .D(n_30528
		), .Z(n_1773));
	notech_reg cr1_reg_4(.CP(n_62614), .D(n_23142), .CD(n_61475), .Q(nbus_14521
		[4]));
	notech_mux2 i_10260(.S(n_328084271), .A(opa[4]), .B(nbus_14521[4]), .Z(n_23142
		));
	notech_reg cr1_reg_5(.CP(n_62614), .D(n_23149), .CD(n_61476), .Q(nbus_14521
		[5]));
	notech_mux2 i_10268(.S(n_328084271), .A(opa[5]), .B(nbus_14521[5]), .Z(n_23149
		));
	notech_ao4 i_114452823(.A(n_55726), .B(n_28100), .C(n_307091753), .D(n_27385
		), .Z(n_1771));
	notech_reg cr1_reg_6(.CP(n_62614), .D(n_23156), .CD(n_61476), .Q(nbus_14521
		[6]));
	notech_mux2 i_10276(.S(n_328084271), .A(opa[6]), .B(nbus_14521[6]), .Z(n_23156
		));
	notech_ao4 i_114352824(.A(n_307991744), .B(n_31476), .C(n_55735), .D(n_31456
		), .Z(n_177092073));
	notech_reg cr1_reg_7(.CP(n_62614), .D(n_23163), .CD(n_61476), .Q(nbus_14521
		[7]));
	notech_mux2 i_10284(.S(n_328084271), .A(opa[7]), .B(nbus_14521[7]), .Z(n_23163
		));
	notech_reg cr1_reg_8(.CP(n_62614), .D(n_23170), .CD(n_61476), .Q(nbus_14521
		[8]));
	notech_mux2 i_10292(.S(n_328084271), .A(opa[8]), .B(nbus_14521[8]), .Z(n_23170
		));
	notech_reg cr1_reg_9(.CP(n_62614), .D(n_23177), .CD(n_61475), .Q(nbus_14521
		[9]));
	notech_mux2 i_10300(.S(n_328084271), .A(opa[9]), .B(nbus_14521[9]), .Z(n_23177
		));
	notech_nand3 i_105552911(.A(n_176592074), .B(n_176492075), .C(n_176392076
		), .Z(n_1767));
	notech_reg cr1_reg_10(.CP(n_62614), .D(n_23185), .CD(n_61474), .Q(nbus_14521
		[10]));
	notech_mux2 i_10308(.S(n_328084271), .A(opa[10]), .B(nbus_14521[10]), .Z
		(n_23185));
	notech_reg cr1_reg_11(.CP(n_62614), .D(n_23192), .CD(n_61475), .Q(nbus_14521
		[11]));
	notech_mux2 i_10316(.S(n_328084271), .A(opa[11]), .B(nbus_14521[11]), .Z
		(n_23192));
	notech_ao4 i_105252914(.A(n_142928706), .B(n_29659), .C(n_128228559), .D
		(n_143028707), .Z(n_176592074));
	notech_reg cr1_reg_12(.CP(n_62614), .D(n_23201), .CD(n_61474), .Q(nbus_14521
		[12]));
	notech_mux2 i_10324(.S(n_328084271), .A(opa[12]), .B(nbus_14521[12]), .Z
		(n_23201));
	notech_ao4 i_105152915(.A(n_142828705), .B(n_55956), .C(n_142728704), .D
		(n_57815), .Z(n_176492075));
	notech_reg cr1_reg_13(.CP(n_62542), .D(n_23210), .CD(n_61474), .Q(nbus_14521
		[13]));
	notech_mux2 i_10332(.S(n_328084271), .A(opa[13]), .B(nbus_14521[13]), .Z
		(n_23210));
	notech_ao4 i_105352913(.A(n_4014), .B(n_28014), .C(n_55726), .D(n_28118)
		, .Z(n_176392076));
	notech_reg cr1_reg_14(.CP(n_62542), .D(n_23217), .CD(n_61475), .Q(nbus_14521
		[14]));
	notech_mux2 i_10340(.S(n_328084271), .A(opa[14]), .B(nbus_14521[14]), .Z
		(n_23217));
	notech_nand2 i_103852928(.A(opbs), .B(opas), .Z(n_176292077));
	notech_reg cr1_reg_15(.CP(n_62542), .D(n_23224), .CD(n_61475), .Q(nbus_14521
		[15]));
	notech_mux2 i_10348(.S(n_328084271), .A(opa[15]), .B(nbus_14521[15]), .Z
		(n_23224));
	notech_ao4 i_103452932(.A(opa[15]), .B(n_306391760), .C(opa[31]), .D(n_57967
		), .Z(n_176192078));
	notech_reg cr1_reg_16(.CP(n_62542), .D(n_23231), .CD(n_61475), .Q(nbus_14521
		[16]));
	notech_mux2 i_10356(.S(n_55005), .A(opa[16]), .B(nbus_14521[16]), .Z(n_23231
		));
	notech_or2 i_103752929(.A(opbs), .B(opas), .Z(n_176092079));
	notech_reg cr1_reg_17(.CP(n_62542), .D(n_23238), .CD(n_61475), .Q(nbus_14521
		[17]));
	notech_mux2 i_10364(.S(n_55005), .A(opa[17]), .B(nbus_14521[17]), .Z(n_23238
		));
	notech_reg cr1_reg_18(.CP(n_62542), .D(n_23245), .CD(n_61475), .Q(nbus_14521
		[18]));
	notech_mux2 i_10372(.S(n_55005), .A(opa[18]), .B(nbus_14521[18]), .Z(n_23245
		));
	notech_reg cr1_reg_19(.CP(n_62542), .D(n_23252), .CD(n_61470), .Q(nbus_14521
		[19]));
	notech_mux2 i_10380(.S(n_55005), .A(opa[19]), .B(nbus_14521[19]), .Z(n_23252
		));
	notech_nand3 i_91953044(.A(n_175192085), .B(n_175092086), .C(n_175692082
		), .Z(n_175792081));
	notech_reg cr1_reg_20(.CP(n_62542), .D(n_23259), .CD(n_61470), .Q(nbus_14521
		[20]));
	notech_mux2 i_10390(.S(n_55005), .A(opa[20]), .B(nbus_14521[20]), .Z(n_23259
		));
	notech_and3 i_91853045(.A(n_1754), .B(n_175392083), .C(n_1558), .Z(n_175692082
		));
	notech_reg cr1_reg_21(.CP(n_62542), .D(n_23266), .CD(n_61469), .Q(nbus_14521
		[21]));
	notech_mux2 i_10398(.S(n_55005), .A(opa[21]), .B(nbus_14521[21]), .Z(n_23266
		));
	notech_reg cr1_reg_22(.CP(n_62614), .D(n_23273), .CD(n_61469), .Q(nbus_14521
		[22]));
	notech_mux2 i_10406(.S(n_55005), .A(opa[22]), .B(nbus_14521[22]), .Z(n_23273
		));
	notech_ao4 i_91253051(.A(n_54649), .B(n_29595), .C(n_28527), .D(n_29594)
		, .Z(n_1754));
	notech_reg cr1_reg_23(.CP(n_62540), .D(n_23280), .CD(n_61470), .Q(nbus_14521
		[23]));
	notech_mux2 i_10414(.S(n_55005), .A(opa[23]), .B(nbus_14521[23]), .Z(n_23280
		));
	notech_ao4 i_91553048(.A(n_303591788), .B(n_28011), .C(n_59326), .D(n_28115
		), .Z(n_175392083));
	notech_reg cr1_reg_24(.CP(n_62540), .D(n_23287), .CD(n_61470), .Q(nbus_14521
		[24]));
	notech_mux2 i_10422(.S(n_55005), .A(opa[24]), .B(nbus_14521[24]), .Z(n_23287
		));
	notech_reg cr1_reg_25(.CP(n_62610), .D(n_23294), .CD(n_61470), .Q(nbus_14521
		[25]));
	notech_mux2 i_10430(.S(n_55005), .A(opa[25]), .B(nbus_14521[25]), .Z(n_23294
		));
	notech_ao4 i_91453049(.A(n_140328680), .B(n_29660), .C(n_133728614), .D(n_140428681
		), .Z(n_175192085));
	notech_reg cr1_reg_26(.CP(n_62610), .D(n_23301), .CD(n_61470), .Q(nbus_14521
		[26]));
	notech_mux2 i_10438(.S(n_55005), .A(opa[26]), .B(nbus_14521[26]), .Z(n_23301
		));
	notech_ao4 i_91353050(.A(n_140228679), .B(n_55947), .C(n_140128678), .D(n_57783
		), .Z(n_175092086));
	notech_reg cr1_reg_27(.CP(n_62610), .D(n_23308), .CD(n_61470), .Q(nbus_14521
		[27]));
	notech_mux2 i_10446(.S(n_55005), .A(opa[27]), .B(nbus_14521[27]), .Z(n_23308
		));
	notech_nand2 i_2653928(.A(opc_10[26]), .B(n_62794), .Z(n_174992087));
	notech_reg cr1_reg_28(.CP(n_62610), .D(n_23316), .CD(n_61469), .Q(nbus_14521
		[28]));
	notech_mux2 i_10454(.S(n_55005), .A(opa[28]), .B(nbus_14521[28]), .Z(n_23316
		));
	notech_and3 i_68253918(.A(n_174692090), .B(n_174592091), .C(n_3884), .Z(n_174892088
		));
	notech_reg cr1_reg_29(.CP(n_62610), .D(n_23322), .CD(n_61469), .Q(nbus_14521
		[29]));
	notech_mux2 i_10462(.S(n_55005), .A(opa[29]), .B(nbus_14521[29]), .Z(n_23322
		));
	notech_reg cr1_reg_30(.CP(n_62610), .D(n_23328), .CD(n_61469), .Q(nbus_14521
		[30]));
	notech_mux2 i_10470(.S(n_55005), .A(opa[30]), .B(nbus_14521[30]), .Z(n_23328
		));
	notech_ao4 i_47153480(.A(n_309591728), .B(n_29660), .C(n_133728614), .D(n_30803
		), .Z(n_174692090));
	notech_reg cr1_reg_31(.CP(n_62610), .D(n_23334), .CD(n_61469), .Q(nbus_14521
		[31]));
	notech_mux2 i_10478(.S(n_55005), .A(opa[31]), .B(nbus_14521[31]), .Z(n_23334
		));
	notech_ao4 i_47053481(.A(n_304691777), .B(n_55947), .C(n_309491729), .D(n_57783
		), .Z(n_174592091));
	notech_reg cr2_reg_reg_0(.CP(n_62610), .D(n_23340), .CD(n_61469), .Q(cr2_reg
		[0]));
	notech_mux2 i_10486(.S(\nbus_11297[0] ), .A(cr2_reg[0]), .B(n_12443), .Z
		(n_23340));
	notech_nand2 i_2753927(.A(opc_10[28]), .B(n_62794), .Z(n_174492092));
	notech_reg cr2_reg_reg_1(.CP(n_62610), .D(n_23346), .CD(n_61469), .Q(cr2_reg
		[1]));
	notech_mux2 i_10494(.S(\nbus_11297[0] ), .A(cr2_reg[1]), .B(n_12449), .Z
		(n_23346));
	notech_nand2 i_2853926(.A(opc_10[29]), .B(n_62794), .Z(n_174392093));
	notech_reg cr2_reg_reg_2(.CP(n_62694), .D(n_23352), .CD(n_61469), .Q(cr2_reg
		[2]));
	notech_mux2 i_10502(.S(\nbus_11297[0] ), .A(cr2_reg[2]), .B(n_12455), .Z
		(n_23352));
	notech_nand2 i_42353919(.A(opc[26]), .B(n_62794), .Z(n_174292094));
	notech_reg cr2_reg_reg_3(.CP(n_62694), .D(n_23358), .CD(n_61469), .Q(cr2_reg
		[3]));
	notech_mux2 i_10510(.S(\nbus_11297[0] ), .A(cr2_reg[3]), .B(n_12461), .Z
		(n_23358));
	notech_reg cr2_reg_reg_4(.CP(n_62694), .D(n_23364), .CD(n_61469), .Q(cr2_reg
		[4]));
	notech_mux2 i_10518(.S(\nbus_11297[0] ), .A(cr2_reg[4]), .B(n_12467), .Z
		(n_23364));
	notech_reg cr2_reg_reg_5(.CP(n_62694), .D(n_23370), .CD(n_61469), .Q(cr2_reg
		[5]));
	notech_mux2 i_10526(.S(\nbus_11297[0] ), .A(cr2_reg[5]), .B(n_12473), .Z
		(n_23370));
	notech_ao4 i_36353583(.A(n_56547), .B(n_28587), .C(n_56557), .D(n_27888)
		, .Z(n_173992096));
	notech_reg cr2_reg_reg_6(.CP(n_62694), .D(n_23376), .CD(n_61471), .Q(cr2_reg
		[6]));
	notech_mux2 i_10534(.S(\nbus_11297[0] ), .A(cr2_reg[6]), .B(n_12479), .Z
		(n_23376));
	notech_ao4 i_36253584(.A(n_56566), .B(n_28554), .C(n_56579), .D(n_28510)
		, .Z(n_173892097));
	notech_reg cr2_reg_reg_7(.CP(n_62694), .D(n_23382), .CD(n_61471), .Q(cr2_reg
		[7]));
	notech_mux2 i_10542(.S(\nbus_11297[0] ), .A(cr2_reg[7]), .B(n_12485), .Z
		(n_23382));
	notech_and2 i_36653580(.A(n_173692098), .B(n_1735), .Z(n_1737));
	notech_reg cr2_reg_reg_8(.CP(n_62694), .D(n_23389), .CD(n_61471), .Q(cr2_reg
		[8]));
	notech_mux2 i_10550(.S(\nbus_11297[0] ), .A(cr2_reg[8]), .B(n_12491), .Z
		(n_23389));
	notech_ao4 i_36153585(.A(n_56592), .B(n_28184), .C(n_56601), .D(n_28477)
		, .Z(n_173692098));
	notech_reg cr2_reg_reg_9(.CP(n_62694), .D(n_23395), .CD(n_61471), .Q(cr2_reg
		[9]));
	notech_mux2 i_10558(.S(\nbus_11297[0] ), .A(cr2_reg[9]), .B(n_12497), .Z
		(n_23395));
	notech_ao4 i_36053586(.A(n_56614), .B(n_28413), .C(n_56627), .D(n_28445)
		, .Z(n_1735));
	notech_reg cr2_reg_reg_10(.CP(n_62694), .D(n_23401), .CD(n_61471), .Q(cr2_reg
		[10]));
	notech_mux2 i_10566(.S(\nbus_11297[0] ), .A(cr2_reg[10]), .B(n_12503), .Z
		(n_23401));
	notech_and4 i_36853578(.A(n_173292101), .B(n_173192102), .C(n_172992104)
		, .D(n_172892105), .Z(n_173492099));
	notech_reg cr2_reg_reg_11(.CP(n_62694), .D(n_23407), .CD(n_61472), .Q(cr2_reg
		[11]));
	notech_mux2 i_10574(.S(\nbus_11297[0] ), .A(cr2_reg[11]), .B(n_12509), .Z
		(n_23407));
	notech_reg cr2_reg_reg_12(.CP(n_62694), .D(n_23413), .CD(n_61472), .Q(cr2_reg
		[12]));
	notech_mux2 i_10582(.S(\nbus_11297[0] ), .A(cr2_reg[12]), .B(n_12515), .Z
		(n_23413));
	notech_ao4 i_35953587(.A(n_56485), .B(n_28349), .C(n_56498), .D(n_28381)
		, .Z(n_173292101));
	notech_reg cr2_reg_reg_13(.CP(n_62694), .D(n_23419), .CD(n_61471), .Q(cr2_reg
		[13]));
	notech_mux2 i_10593(.S(\nbus_11297[0] ), .A(cr2_reg[13]), .B(n_12521), .Z
		(n_23419));
	notech_ao4 i_35853588(.A(n_56513), .B(n_29607), .C(n_56527), .D(n_28316)
		, .Z(n_173192102));
	notech_reg cr2_reg_reg_14(.CP(n_62694), .D(n_23425), .CD(n_61471), .Q(cr2_reg
		[14]));
	notech_mux2 i_10601(.S(\nbus_11297[0] ), .A(cr2_reg[14]), .B(n_12527), .Z
		(n_23425));
	notech_reg cr2_reg_reg_15(.CP(n_62694), .D(n_23431), .CD(n_61471), .Q(cr2_reg
		[15]));
	notech_mux2 i_10609(.S(\nbus_11297[0] ), .A(cr2_reg[15]), .B(n_12533), .Z
		(n_23431));
	notech_ao4 i_35753589(.A(n_56636), .B(n_28283), .C(n_56916), .D(n_29606)
		, .Z(n_172992104));
	notech_reg cr2_reg_reg_16(.CP(n_62694), .D(n_23437), .CD(n_61470), .Q(cr2_reg
		[16]));
	notech_mux2 i_10617(.S(\nbus_11297[0] ), .A(cr2_reg[16]), .B(n_12539), .Z
		(n_23437));
	notech_ao4 i_35653590(.A(n_56649), .B(n_28216), .C(n_56662), .D(n_28251)
		, .Z(n_172892105));
	notech_reg cr2_reg_reg_17(.CP(n_62694), .D(n_23443), .CD(n_61470), .Q(cr2_reg
		[17]));
	notech_mux2 i_10625(.S(\nbus_11297[0] ), .A(cr2_reg[17]), .B(n_12545), .Z
		(n_23443));
	notech_nand2 i_40153921(.A(opc[28]), .B(n_62794), .Z(n_172792106));
	notech_reg cr2_reg_reg_18(.CP(n_62694), .D(n_23449), .CD(n_61470), .Q(cr2_reg
		[18]));
	notech_mux2 i_10633(.S(n_55016), .A(cr2_reg[18]), .B(n_12551), .Z(n_23449
		));
	notech_reg cr2_reg_reg_19(.CP(n_62694), .D(n_23455), .CD(n_61470), .Q(cr2_reg
		[19]));
	notech_mux2 i_10642(.S(n_55016), .A(cr2_reg[19]), .B(n_12557), .Z(n_23455
		));
	notech_reg cr2_reg_reg_20(.CP(n_62610), .D(n_23461), .CD(n_61470), .Q(cr2_reg
		[20]));
	notech_mux2 i_10650(.S(n_55016), .A(cr2_reg[20]), .B(n_12563), .Z(n_23461
		));
	notech_ao4 i_28653659(.A(n_56547), .B(n_28589), .C(n_56557), .D(n_27890)
		, .Z(n_172492109));
	notech_reg cr2_reg_reg_21(.CP(n_62694), .D(n_23467), .CD(n_61471), .Q(cr2_reg
		[21]));
	notech_mux2 i_10658(.S(n_55016), .A(cr2_reg[21]), .B(n_12569), .Z(n_23467
		));
	notech_ao4 i_28553660(.A(n_56566), .B(n_28556), .C(n_56579), .D(n_28512)
		, .Z(n_1723));
	notech_reg cr2_reg_reg_22(.CP(n_62612), .D(n_23473), .CD(n_61471), .Q(cr2_reg
		[22]));
	notech_mux2 i_10666(.S(n_55016), .A(cr2_reg[22]), .B(n_12575), .Z(n_23473
		));
	notech_and2 i_28953656(.A(n_172192110), .B(n_172092111), .Z(n_1722));
	notech_reg cr2_reg_reg_23(.CP(n_62612), .D(n_23479), .CD(n_61471), .Q(cr2_reg
		[23]));
	notech_mux2 i_10674(.S(n_55016), .A(cr2_reg[23]), .B(n_12581), .Z(n_23479
		));
	notech_ao4 i_28453661(.A(n_56592), .B(n_28186), .C(n_56601), .D(n_28479)
		, .Z(n_172192110));
	notech_reg cr2_reg_reg_24(.CP(n_62612), .D(n_23485), .CD(n_61471), .Q(cr2_reg
		[24]));
	notech_mux2 i_10682(.S(n_55016), .A(cr2_reg[24]), .B(n_12587), .Z(n_23485
		));
	notech_ao4 i_28353662(.A(n_56614), .B(n_28415), .C(n_56627), .D(n_28447)
		, .Z(n_172092111));
	notech_reg cr2_reg_reg_25(.CP(n_62612), .D(n_23491), .CD(n_61482), .Q(cr2_reg
		[25]));
	notech_mux2 i_10690(.S(n_55016), .A(cr2_reg[25]), .B(n_12593), .Z(n_23491
		));
	notech_and4 i_29153654(.A(n_171792114), .B(n_171692115), .C(n_171492117)
		, .D(n_171392118), .Z(n_171992112));
	notech_reg cr2_reg_reg_26(.CP(n_62612), .D(n_23497), .CD(n_61482), .Q(cr2_reg
		[26]));
	notech_mux2 i_10698(.S(n_55016), .A(cr2_reg[26]), .B(n_12599), .Z(n_23497
		));
	notech_reg cr2_reg_reg_27(.CP(n_62612), .D(n_23503), .CD(n_61482), .Q(cr2_reg
		[27]));
	notech_mux2 i_10706(.S(n_55016), .A(cr2_reg[27]), .B(n_12605), .Z(n_23503
		));
	notech_ao4 i_28253663(.A(n_56489), .B(n_28351), .C(n_56502), .D(n_28383)
		, .Z(n_171792114));
	notech_reg cr2_reg_reg_28(.CP(n_62612), .D(n_23515), .CD(n_61482), .Q(cr2_reg
		[28]));
	notech_mux2 i_10714(.S(n_55016), .A(cr2_reg[28]), .B(n_12611), .Z(n_23515
		));
	notech_ao4 i_28153664(.A(n_56513), .B(n_29611), .C(n_56532), .D(n_28318)
		, .Z(n_171692115));
	notech_reg cr2_reg_reg_29(.CP(n_62612), .D(n_23521), .CD(n_61482), .Q(cr2_reg
		[29]));
	notech_mux2 i_10723(.S(n_55016), .A(cr2_reg[29]), .B(n_12617), .Z(n_23521
		));
	notech_reg cr2_reg_reg_30(.CP(n_62612), .D(n_23527), .CD(n_61482), .Q(cr2_reg
		[30]));
	notech_mux2 i_10731(.S(n_55016), .A(cr2_reg[30]), .B(n_12623), .Z(n_23527
		));
	notech_ao4 i_28053665(.A(n_56640), .B(n_28285), .C(n_56916), .D(n_29610)
		, .Z(n_171492117));
	notech_reg cr2_reg_reg_31(.CP(n_62612), .D(n_23533), .CD(n_61483), .Q(cr2_reg
		[31]));
	notech_mux2 i_10739(.S(n_55016), .A(cr2_reg[31]), .B(n_12629), .Z(n_23533
		));
	notech_ao4 i_27953666(.A(n_56653), .B(n_28218), .C(n_56666), .D(n_28253)
		, .Z(n_171392118));
	notech_reg cr3_reg_0(.CP(n_62612), .D(n_23539), .CD(n_61482), .Q(\nbus_14520[0] 
		));
	notech_mux2 i_10747(.S(n_328090778), .A(opa[0]), .B(\nbus_14520[0] ), .Z
		(n_23539));
	notech_reg cr3_reg_1(.CP(n_62612), .D(n_23545), .CD(n_61482), .Q(\nbus_14520[1] 
		));
	notech_mux2 i_10755(.S(n_328090778), .A(opa[1]), .B(\nbus_14520[1] ), .Z
		(n_23545));
	notech_reg cr3_reg_2(.CP(n_62612), .D(n_23551), .CD(n_61482), .Q(\nbus_14520[2] 
		));
	notech_mux2 i_10763(.S(n_328090778), .A(opa[2]), .B(\nbus_14520[2] ), .Z
		(n_23551));
	notech_nand3 i_25853686(.A(n_170492127), .B(n_170392128), .C(n_170992122
		), .Z(n_171092121));
	notech_reg cr3_reg_3(.CP(n_62612), .D(n_23557), .CD(n_61481), .Q(\nbus_14520[3] 
		));
	notech_mux2 i_10771(.S(n_328090778), .A(opa[3]), .B(\nbus_14520[3] ), .Z
		(n_23557));
	notech_and3 i_25753687(.A(n_170792124), .B(n_170692125), .C(n_1509), .Z(n_170992122
		));
	notech_reg cr3_reg_4(.CP(n_62612), .D(n_23563), .CD(n_61481), .Q(\nbus_14520[4] 
		));
	notech_mux2 i_10779(.S(n_328090778), .A(opa[4]), .B(\nbus_14520[4] ), .Z
		(n_23563));
	notech_reg cr3_reg_5(.CP(n_62612), .D(n_23570), .CD(n_61481), .Q(\nbus_14520[5] 
		));
	notech_mux2 i_10787(.S(n_328090778), .A(opa[5]), .B(\nbus_14520[5] ), .Z
		(n_23570));
	notech_ao4 i_24853693(.A(n_309091733), .B(n_55956), .C(n_308991734), .D(n_57815
		), .Z(n_170792124));
	notech_reg cr3_reg_6(.CP(n_62612), .D(n_23576), .CD(n_61481), .Q(\nbus_14520[6] 
		));
	notech_mux2 i_10795(.S(n_328090778), .A(opa[6]), .B(\nbus_14520[6] ), .Z
		(n_23576));
	notech_ao4 i_25153690(.A(n_121628493), .B(n_28014), .C(n_309291731), .D(n_28118
		), .Z(n_170692125));
	notech_reg cr3_reg_7(.CP(n_62612), .D(n_23582), .CD(n_61481), .Q(\nbus_14520[7] 
		));
	notech_mux2 i_10803(.S(n_328090778), .A(opa[7]), .B(\nbus_14520[7] ), .Z
		(n_23582));
	notech_reg cr3_reg_8(.CP(n_62612), .D(n_23588), .CD(n_61482), .Q(\nbus_14520[8] 
		));
	notech_mux2 i_10811(.S(n_328090778), .A(opa[8]), .B(\nbus_14520[8] ), .Z
		(n_23588));
	notech_ao4 i_25053691(.A(n_56091), .B(n_29593), .C(n_29659), .D(n_26765)
		, .Z(n_170492127));
	notech_reg cr3_reg_9(.CP(n_62540), .D(n_23594), .CD(n_61482), .Q(\nbus_14520[9] 
		));
	notech_mux2 i_10819(.S(n_328090778), .A(opa[9]), .B(\nbus_14520[9] ), .Z
		(n_23594));
	notech_ao4 i_24953692(.A(n_122428501), .B(n_28155), .C(n_122528502), .D(n_128228559
		), .Z(n_170392128));
	notech_reg cr3_reg_10(.CP(n_62540), .D(n_23600), .CD(n_61481), .Q(\nbus_14520[10] 
		));
	notech_mux2 i_10827(.S(n_328090778), .A(opa[10]), .B(\nbus_14520[10] ), 
		.Z(n_23600));
	notech_nand2 i_42253920(.A(opc[29]), .B(n_62794), .Z(n_170292129));
	notech_reg cr3_reg_11(.CP(n_62540), .D(n_23606), .CD(n_61482), .Q(\nbus_14520[11] 
		));
	notech_mux2 i_10835(.S(n_328090778), .A(opa[11]), .B(\nbus_14520[11] ), 
		.Z(n_23606));
	notech_reg cr3_reg_12(.CP(n_62540), .D(n_23612), .CD(n_61485), .Q(cr3[12
		]));
	notech_mux2 i_10843(.S(n_328090778), .A(opa[12]), .B(cr3[12]), .Z(n_23612
		));
	notech_reg cr3_reg_13(.CP(n_62540), .D(n_23618), .CD(n_61485), .Q(cr3[13
		]));
	notech_mux2 i_10851(.S(n_328090778), .A(opa[13]), .B(cr3[13]), .Z(n_23618
		));
	notech_ao4 i_22653712(.A(n_56592), .B(n_28187), .C(n_56547), .D(n_28590)
		, .Z(n_169992130));
	notech_reg cr3_reg_14(.CP(n_62540), .D(n_23624), .CD(n_61483), .Q(cr3[14
		]));
	notech_mux2 i_10859(.S(n_328090778), .A(opa[14]), .B(cr3[14]), .Z(n_23624
		));
	notech_ao4 i_22553713(.A(n_56557), .B(n_27891), .C(n_56566), .D(n_28557)
		, .Z(n_1698));
	notech_reg cr3_reg_15(.CP(n_62540), .D(n_23632), .CD(n_61485), .Q(cr3[15
		]));
	notech_mux2 i_10867(.S(n_328090778), .A(n_60102), .B(cr3[15]), .Z(n_23632
		));
	notech_and2 i_22953709(.A(n_169692132), .B(n_1695), .Z(n_169792131));
	notech_reg cr3_reg_16(.CP(n_62540), .D(n_23638), .CD(n_61485), .Q(cr3[16
		]));
	notech_mux2 i_10875(.S(n_55918), .A(opa[16]), .B(cr3[16]), .Z(n_23638)
		);
	notech_ao4 i_22453714(.A(n_56583), .B(n_28513), .C(n_56605), .D(n_28480)
		, .Z(n_169692132));
	notech_reg cr3_reg_17(.CP(n_62540), .D(n_23644), .CD(n_61485), .Q(cr3[17
		]));
	notech_mux2 i_10883(.S(n_55918), .A(opa[17]), .B(cr3[17]), .Z(n_23644)
		);
	notech_ao4 i_22353715(.A(n_56614), .B(n_28416), .C(n_56627), .D(n_28448)
		, .Z(n_1695));
	notech_reg cr3_reg_18(.CP(n_62610), .D(n_23650), .CD(n_61485), .Q(cr3[18
		]));
	notech_mux2 i_10891(.S(n_55918), .A(opa[18]), .B(cr3[18]), .Z(n_23650)
		);
	notech_and4 i_23153707(.A(n_1692), .B(n_169192135), .C(n_1689), .D(n_168892137
		), .Z(n_169492133));
	notech_reg cr3_reg_19(.CP(n_62604), .D(n_23656), .CD(n_61485), .Q(cr3[19
		]));
	notech_mux2 i_10899(.S(n_55918), .A(opa[19]), .B(cr3[19]), .Z(n_23656)
		);
	notech_reg cr3_reg_20(.CP(n_62538), .D(n_23662), .CD(n_61485), .Q(cr3[20
		]));
	notech_mux2 i_10907(.S(n_55918), .A(opa[20]), .B(cr3[20]), .Z(n_23662)
		);
	notech_ao4 i_22253716(.A(n_56489), .B(n_28352), .C(n_56502), .D(n_28384)
		, .Z(n_1692));
	notech_reg cr3_reg_21(.CP(n_62604), .D(n_23668), .CD(n_61483), .Q(cr3[21
		]));
	notech_mux2 i_10915(.S(n_55918), .A(opa[21]), .B(cr3[21]), .Z(n_23668)
		);
	notech_ao4 i_22053717(.A(n_56513), .B(n_29613), .C(n_56532), .D(n_28319)
		, .Z(n_169192135));
	notech_reg cr3_reg_22(.CP(n_62604), .D(n_23674), .CD(n_61483), .Q(cr3[22
		]));
	notech_mux2 i_10923(.S(n_55918), .A(opa[22]), .B(cr3[22]), .Z(n_23674)
		);
	notech_reg cr3_reg_23(.CP(n_62604), .D(n_23680), .CD(n_61483), .Q(cr3[23
		]));
	notech_mux2 i_10931(.S(n_55918), .A(opa[23]), .B(cr3[23]), .Z(n_23680)
		);
	notech_ao4 i_21953718(.A(n_56640), .B(n_28286), .C(n_56916), .D(n_29612)
		, .Z(n_1689));
	notech_reg cr3_reg_24(.CP(n_62604), .D(n_23686), .CD(n_61483), .Q(cr3[24
		]));
	notech_mux2 i_10939(.S(n_55918), .A(opa[24]), .B(cr3[24]), .Z(n_23686)
		);
	notech_ao4 i_21853719(.A(n_56653), .B(n_28219), .C(n_56666), .D(n_28254)
		, .Z(n_168892137));
	notech_reg cr3_reg_25(.CP(n_62604), .D(n_23692), .CD(n_61483), .Q(cr3[25
		]));
	notech_mux2 i_10947(.S(n_55918), .A(opa[25]), .B(cr3[25]), .Z(n_23692)
		);
	notech_ao4 i_18553750(.A(n_57671), .B(n_306391760), .C(n_57967), .D(n_59726
		), .Z(n_168792138));
	notech_reg cr3_reg_26(.CP(n_62604), .D(n_23698), .CD(n_61483), .Q(cr3[26
		]));
	notech_mux2 i_10955(.S(n_55918), .A(opa[26]), .B(cr3[26]), .Z(n_23698)
		);
	notech_nao3 i_167755569(.A(n_27377), .B(n_60321), .C(n_26702), .Z(n_1686
		));
	notech_reg cr3_reg_27(.CP(n_62604), .D(n_23704), .CD(n_61483), .Q(cr3[27
		]));
	notech_mux2 i_10963(.S(n_55918), .A(opa[27]), .B(cr3[27]), .Z(n_23704)
		);
	notech_reg cr3_reg_28(.CP(n_62604), .D(n_23710), .CD(n_61483), .Q(cr3[28
		]));
	notech_mux2 i_10971(.S(n_55918), .A(opa[28]), .B(cr3[28]), .Z(n_23710)
		);
	notech_reg cr3_reg_29(.CP(n_62604), .D(n_23716), .CD(n_61483), .Q(cr3[29
		]));
	notech_mux2 i_10979(.S(n_55918), .A(opa[29]), .B(cr3[29]), .Z(n_23716)
		);
	notech_reg cr3_reg_30(.CP(n_62690), .D(n_23722), .CD(n_61483), .Q(cr3[30
		]));
	notech_mux2 i_10987(.S(n_55918), .A(opa[30]), .B(cr3[30]), .Z(n_23722)
		);
	notech_ao4 i_8953823(.A(n_56547), .B(n_28588), .C(n_56557), .D(n_27889),
		 .Z(n_168292141));
	notech_reg cr3_reg_31(.CP(n_62690), .D(n_23729), .CD(n_61477), .Q(cr3[31
		]));
	notech_mux2 i_10995(.S(n_55918), .A(opa[31]), .B(cr3[31]), .Z(n_23729)
		);
	notech_ao4 i_8853824(.A(n_56570), .B(n_28555), .C(n_56583), .D(n_28511),
		 .Z(n_168192142));
	notech_reg opa_reg_0(.CP(n_62690), .D(n_23737), .CD(n_61477), .Q(opa[0])
		);
	notech_mux2 i_11003(.S(n_27702), .A(opa[0]), .B(n_27700), .Z(n_23737));
	notech_and2 i_9253820(.A(n_167992143), .B(n_167892144), .Z(n_1680));
	notech_reg opa_reg_1(.CP(n_62690), .D(n_23744), .CD(n_61477), .Q(opa[1])
		);
	notech_mux2 i_11011(.S(n_27702), .A(opa[1]), .B(n_27701), .Z(n_23744));
	notech_ao4 i_8753825(.A(n_56592), .B(n_28185), .C(n_56605), .D(n_28478),
		 .Z(n_167992143));
	notech_reg opa_reg_2(.CP(n_62690), .D(n_23751), .CD(n_61477), .Q(opa[2])
		);
	notech_mux2 i_11019(.S(n_27702), .A(opa[2]), .B(n_26995), .Z(n_23751));
	notech_ao4 i_8653826(.A(n_56614), .B(n_28414), .C(n_56627), .D(n_28446),
		 .Z(n_167892144));
	notech_reg opa_reg_3(.CP(n_62690), .D(n_23762), .CD(n_61477), .Q(opa[3])
		);
	notech_mux2 i_11027(.S(n_27702), .A(opa[3]), .B(n_26996), .Z(n_23762));
	notech_and4 i_9453818(.A(n_167592147), .B(n_1674), .C(n_1672), .D(n_1671
		), .Z(n_167792145));
	notech_reg opa_reg_4(.CP(n_62690), .D(n_23769), .CD(n_61477), .Q(opa[4])
		);
	notech_mux2 i_11035(.S(n_27702), .A(opa[4]), .B(n_26997), .Z(n_23769));
	notech_reg opa_reg_5(.CP(n_62690), .D(n_23778), .CD(n_61477), .Q(opa[5])
		);
	notech_mux2 i_11043(.S(n_27702), .A(opa[5]), .B(n_27128), .Z(n_23778));
	notech_ao4 i_8553827(.A(n_56489), .B(n_28350), .C(n_56502), .D(n_28382),
		 .Z(n_167592147));
	notech_reg opa_reg_6(.CP(n_62690), .D(n_23786), .CD(n_61477), .Q(opa[6])
		);
	notech_mux2 i_11051(.S(n_27702), .A(opa[6]), .B(n_26998), .Z(n_23786));
	notech_ao4 i_8453828(.A(n_56518), .B(n_29609), .C(n_56532), .D(n_28317),
		 .Z(n_1674));
	notech_reg opa_reg_7(.CP(n_62690), .D(n_23793), .CD(n_61477), .Q(opa[7])
		);
	notech_mux2 i_11059(.S(n_27702), .A(opa[7]), .B(n_27000), .Z(n_23793));
	notech_reg opa_reg_8(.CP(n_62690), .D(n_23801), .CD(n_61477), .Q(opa[8])
		);
	notech_mux2 i_11067(.S(n_27711), .A(opa[8]), .B(n_27703), .Z(n_23801));
	notech_ao4 i_8353829(.A(n_56636), .B(n_28284), .C(n_56916), .D(n_29608),
		 .Z(n_1672));
	notech_reg opa_reg_9(.CP(n_62690), .D(n_23808), .CD(n_61476), .Q(opa[9])
		);
	notech_mux2 i_11075(.S(n_27711), .A(opa[9]), .B(n_27704), .Z(n_23808));
	notech_ao4 i_8253830(.A(n_56653), .B(n_28217), .C(n_56666), .D(n_28252),
		 .Z(n_1671));
	notech_reg opa_reg_10(.CP(n_62690), .D(n_23815), .CD(n_61476), .Q(opa[10
		]));
	notech_mux2 i_11083(.S(n_27711), .A(opa[10]), .B(n_27705), .Z(n_23815)
		);
	notech_and4 i_2717616(.A(n_174892088), .B(n_1834), .C(n_1836), .D(n_1660
		), .Z(n_1670));
	notech_reg opa_reg_11(.CP(n_62690), .D(n_23822), .CD(n_61476), .Q(opa[11
		]));
	notech_mux2 i_11091(.S(n_27711), .A(opa[11]), .B(n_27706), .Z(n_23822)
		);
	notech_reg opa_reg_12(.CP(n_62690), .D(n_23829), .CD(n_61476), .Q(opa[12
		]));
	notech_mux2 i_11099(.S(n_27711), .A(opa[12]), .B(n_27707), .Z(n_23829)
		);
	notech_reg opa_reg_13(.CP(n_62690), .D(n_23837), .CD(n_61476), .Q(opa[13
		]));
	notech_mux2 i_11107(.S(n_27711), .A(opa[13]), .B(n_27708), .Z(n_23837)
		);
	notech_or4 i_169352283(.A(n_56827), .B(n_56944), .C(n_56583), .D(n_28011
		), .Z(n_1667));
	notech_reg opa_reg_14(.CP(n_62690), .D(n_23844), .CD(n_61476), .Q(opa[14
		]));
	notech_mux2 i_11115(.S(n_27711), .A(opa[14]), .B(n_27709), .Z(n_23844)
		);
	notech_reg opa_reg_15(.CP(n_62690), .D(n_23851), .CD(n_61477), .Q(opa[15
		]));
	notech_mux2 i_11123(.S(n_27711), .A(n_60102), .B(n_27710), .Z(n_23851)
		);
	notech_reg opa_reg_16(.CP(n_62690), .D(n_23858), .CD(n_61476), .Q(opa[16
		]));
	notech_mux2 i_11131(.S(n_27713), .A(opa[16]), .B(n_22311), .Z(n_23858)
		);
	notech_reg opa_reg_17(.CP(n_62744), .D(n_23865), .CD(n_61476), .Q(opa[17
		]));
	notech_mux2 i_11139(.S(n_27713), .A(opa[17]), .B(n_22317), .Z(n_23865)
		);
	notech_reg opa_reg_18(.CP(n_62688), .D(n_23873), .CD(n_61480), .Q(opa[18
		]));
	notech_mux2 i_11147(.S(n_27713), .A(opa[18]), .B(n_22323), .Z(n_23873)
		);
	notech_reg opa_reg_19(.CP(n_62744), .D(n_23880), .CD(n_61481), .Q(opa[19
		]));
	notech_mux2 i_11155(.S(n_27713), .A(opa[19]), .B(n_22329), .Z(n_23880)
		);
	notech_reg opa_reg_20(.CP(n_62744), .D(n_23887), .CD(n_61480), .Q(opa[20
		]));
	notech_mux2 i_11163(.S(n_27713), .A(opa[20]), .B(n_22335), .Z(n_23887)
		);
	notech_or2 i_169452282(.A(n_151128788), .B(n_3983), .Z(n_1660));
	notech_reg opa_reg_21(.CP(n_62744), .D(n_23894), .CD(n_61480), .Q(opa[21
		]));
	notech_mux2 i_11171(.S(n_27713), .A(opa[21]), .B(n_22341), .Z(n_23894)
		);
	notech_or4 i_2917042(.A(n_1657), .B(n_1658), .C(n_1648), .D(n_27772), .Z
		(n_1659));
	notech_reg opa_reg_22(.CP(n_62744), .D(n_23901), .CD(n_61481), .Q(opa[22
		]));
	notech_mux2 i_11179(.S(n_27713), .A(opa[22]), .B(n_22347), .Z(n_23901)
		);
	notech_ao3 i_159252384(.A(opc[28]), .B(n_62772), .C(n_307891745), .Z(n_1658
		));
	notech_reg opa_reg_23(.CP(n_62744), .D(n_23909), .CD(n_61481), .Q(opa[23
		]));
	notech_mux2 i_11187(.S(n_27713), .A(opa[23]), .B(n_22353), .Z(n_23909)
		);
	notech_ao3 i_159152385(.A(opc_10[28]), .B(n_62794), .C(n_308791736), .Z(n_1657
		));
	notech_reg opa_reg_24(.CP(n_62744), .D(n_23916), .CD(n_61481), .Q(opa[24
		]));
	notech_mux2 i_11195(.S(n_27713), .A(opa[24]), .B(n_22359), .Z(n_23916)
		);
	notech_reg opa_reg_25(.CP(n_62744), .D(n_23923), .CD(n_61481), .Q(opa[25
		]));
	notech_mux2 i_11203(.S(n_27713), .A(opa[25]), .B(n_22365), .Z(n_23923)
		);
	notech_reg opa_reg_26(.CP(n_62744), .D(n_23930), .CD(n_61481), .Q(opa[26
		]));
	notech_mux2 i_11211(.S(n_27713), .A(opa[26]), .B(n_22371), .Z(n_23930)
		);
	notech_reg opa_reg_27(.CP(n_62744), .D(n_23938), .CD(n_61480), .Q(opa[27
		]));
	notech_mux2 i_11219(.S(n_27713), .A(opa[27]), .B(n_22377), .Z(n_23938)
		);
	notech_reg opa_reg_28(.CP(n_62744), .D(n_23949), .CD(n_61480), .Q(opa[28
		]));
	notech_mux2 i_11227(.S(n_27713), .A(opa[28]), .B(n_22383), .Z(n_23949)
		);
	notech_reg opa_reg_29(.CP(n_62744), .D(n_23955), .CD(n_61480), .Q(opa[29
		]));
	notech_mux2 i_11235(.S(n_27713), .A(opa[29]), .B(n_22389), .Z(n_23955)
		);
	notech_reg opa_reg_30(.CP(n_62744), .D(n_23961), .CD(n_61477), .Q(opa[30
		]));
	notech_mux2 i_11243(.S(n_27713), .A(opa[30]), .B(n_22395), .Z(n_23961)
		);
	notech_reg opa_reg_31(.CP(n_62744), .D(n_23967), .CD(n_61480), .Q(opa[31
		]));
	notech_mux2 i_11251(.S(n_27713), .A(opa[31]), .B(n_22401), .Z(n_23967)
		);
	notech_reg tcmp_reg(.CP(n_62744), .D(n_23973), .CD(n_61480), .Q(tcmp));
	notech_mux2 i_11259(.S(n_3818), .A(n_328590783), .B(tcmp), .Z(n_23973)
		);
	notech_nor2 i_159052386(.A(n_3982), .B(n_150228779), .Z(n_1648));
	notech_reg sema_rw_reg(.CP(n_62744), .D(n_23979), .CD(n_61480), .Q(sema_rw
		));
	notech_mux2 i_11267(.S(n_23569), .A(sema_rw), .B(n_27715), .Z(n_23979)
		);
	notech_or4 i_3021939(.A(n_1645), .B(n_1646), .C(n_1638), .D(n_27796), .Z
		(n_1647));
	notech_reg_set fsm_reg_0(.CP(n_62744), .D(n_23985), .SD(n_61480), .Q(fsm
		[0]));
	notech_mux2 i_11275(.S(\nbus_11340[0] ), .A(fsm[0]), .B(n_27174), .Z(n_23985
		));
	notech_ao3 i_149552481(.A(opc[29]), .B(\opcode[2] ), .C(n_310891715), .Z
		(n_1646));
	notech_reg_set fsm_reg_1(.CP(n_62744), .D(n_23991), .SD(n_61480), .Q(fsm
		[1]));
	notech_mux2 i_11283(.S(\nbus_11340[0] ), .A(fsm[1]), .B(n_27716), .Z(n_23991
		));
	notech_ao3 i_149452482(.A(opc_10[29]), .B(\opcode[2] ), .C(n_310791716),
		 .Z(n_1645));
	notech_reg_set fsm_reg_2(.CP(n_62744), .D(n_23997), .SD(n_61480), .Q(fsm
		[2]));
	notech_mux2 i_11293(.S(\nbus_11340[0] ), .A(n_61171), .B(n_27718), .Z(n_23997
		));
	notech_reg_set fsm_reg_3(.CP(n_62688), .D(n_24003), .SD(n_61526), .Q(fsm
		[3]));
	notech_mux2 i_11301(.S(\nbus_11340[0] ), .A(fsm[3]), .B(n_19665), .Z(n_24003
		));
	notech_reg fsm_reg_4(.CP(n_62688), .D(n_24009), .CD(n_61526), .Q(fsm[4])
		);
	notech_mux2 i_11309(.S(\nbus_11340[0] ), .A(n_61160), .B(n_27721), .Z(n_24009
		));
	notech_reg vliw_pc_reg_0(.CP(n_62688), .D(n_24015), .CD(n_61526), .Q(vliw_pc
		[0]));
	notech_mux2 i_11317(.S(\nbus_11308[0] ), .A(vliw_pc[0]), .B(n_14515), .Z
		(n_24015));
	notech_reg vliw_pc_reg_1(.CP(n_62688), .D(n_24023), .CD(n_61526), .Q(vliw_pc
		[1]));
	notech_mux2 i_11325(.S(\nbus_11308[0] ), .A(vliw_pc[1]), .B(n_214286416)
		, .Z(n_24023));
	notech_reg vliw_pc_reg_2(.CP(n_62688), .D(n_24030), .CD(n_61526), .Q(vliw_pc
		[2]));
	notech_mux2 i_11333(.S(\nbus_11308[0] ), .A(vliw_pc[2]), .B(n_214386417)
		, .Z(n_24030));
	notech_reg vliw_pc_reg_3(.CP(n_62688), .D(n_24036), .CD(n_61526), .Q(vliw_pc
		[3]));
	notech_mux2 i_11341(.S(\nbus_11308[0] ), .A(vliw_pc[3]), .B(n_214486418)
		, .Z(n_24036));
	notech_nor2 i_149352483(.A(n_148728764), .B(n_3981), .Z(n_1638));
	notech_reg vliw_pc_reg_4(.CP(n_62688), .D(n_24042), .CD(n_61526), .Q(vliw_pc
		[4]));
	notech_mux2 i_11349(.S(\nbus_11308[0] ), .A(vliw_pc[4]), .B(n_214586419)
		, .Z(n_24042));
	notech_or4 i_2721808(.A(n_1635), .B(n_1809), .C(n_1636), .D(n_1624), .Z(n_1637
		));
	notech_reg_set opd_reg_0(.CP(n_62688), .D(n_24048), .SD(1'b1), .Q(opd[0]
		));
	notech_mux2 i_11357(.S(\nbus_11380[0] ), .A(opd[0]), .B(n_25948), .Z(n_24048
		));
	notech_ao3 i_140152569(.A(opc[26]), .B(\opcode[2] ), .C(n_310491719), .Z
		(n_1636));
	notech_reg_set opd_reg_1(.CP(n_62688), .D(n_24054), .SD(1'b1), .Q(opd[1]
		));
	notech_mux2 i_11365(.S(\nbus_11380[0] ), .A(opd[1]), .B(n_27725), .Z(n_24054
		));
	notech_ao3 i_140052570(.A(opc_10[26]), .B(\opcode[2] ), .C(n_301791806),
		 .Z(n_1635));
	notech_reg_set opd_reg_2(.CP(n_62688), .D(n_24060), .SD(1'b1), .Q(opd[2]
		));
	notech_mux2 i_11373(.S(\nbus_11380[0] ), .A(opd[2]), .B(n_25958), .Z(n_24060
		));
	notech_reg_set opd_reg_3(.CP(n_62604), .D(n_24066), .SD(1'b1), .Q(opd[3]
		));
	notech_mux2 i_11381(.S(\nbus_11380[0] ), .A(opd[3]), .B(n_27726), .Z(n_24066
		));
	notech_reg_set opd_reg_4(.CP(n_62538), .D(n_24072), .SD(1'b1), .Q(opd[4]
		));
	notech_mux2 i_11389(.S(\nbus_11380[0] ), .A(opd[4]), .B(n_25968), .Z(n_24072
		));
	notech_reg_set opd_reg_5(.CP(n_62692), .D(n_24078), .SD(1'b1), .Q(opd[5]
		));
	notech_mux2 i_11397(.S(\nbus_11380[0] ), .A(opd[5]), .B(n_25973), .Z(n_24078
		));
	notech_reg_set opd_reg_6(.CP(n_62606), .D(n_24085), .SD(1'b1), .Q(opd[6]
		));
	notech_mux2 i_11405(.S(n_60129), .A(n_25978), .B(opd[6]), .Z(n_24085));
	notech_reg_set opd_reg_7(.CP(n_62606), .D(n_24092), .SD(1'b1), .Q(opd[7]
		));
	notech_mux2 i_11413(.S(n_60129), .A(n_25983), .B(opd[7]), .Z(n_24092));
	notech_reg_set opd_reg_8(.CP(n_62606), .D(n_24099), .SD(1'b1), .Q(opd[8]
		));
	notech_mux2 i_11421(.S(n_60129), .A(n_25988), .B(opd[8]), .Z(n_24099));
	notech_reg_set opd_reg_9(.CP(n_62606), .D(n_24108), .SD(1'b1), .Q(opd[9]
		));
	notech_mux2 i_11429(.S(n_60129), .A(n_25993), .B(opd[9]), .Z(n_24108));
	notech_reg_set opd_reg_10(.CP(n_62606), .D(n_24115), .SD(1'b1), .Q(opd[
		10]));
	notech_mux2 i_11437(.S(n_60129), .A(n_25998), .B(opd[10]), .Z(n_24115)
		);
	notech_reg_set opd_reg_11(.CP(n_62606), .D(n_24122), .SD(1'b1), .Q(opd[
		11]));
	notech_mux2 i_11445(.S(n_60129), .A(n_26003), .B(opd[11]), .Z(n_24122)
		);
	notech_reg_set opd_reg_12(.CP(n_62606), .D(n_24129), .SD(1'b1), .Q(opd[
		12]));
	notech_mux2 i_11453(.S(n_60129), .A(n_26008), .B(opd[12]), .Z(n_24129)
		);
	notech_nor2 i_139952571(.A(n_146428741), .B(n_3983), .Z(n_1624));
	notech_reg_set opd_reg_13(.CP(n_62606), .D(n_24137), .SD(1'b1), .Q(opd[
		13]));
	notech_mux2 i_11461(.S(n_60129), .A(n_26013), .B(opd[13]), .Z(n_24137)
		);
	notech_or4 i_2721552(.A(n_1621), .B(n_179892049), .C(n_1622), .D(n_161292148
		), .Z(n_1623));
	notech_reg_set opd_reg_14(.CP(n_62606), .D(n_24144), .SD(1'b1), .Q(opd[
		14]));
	notech_mux2 i_11469(.S(n_60129), .A(n_26018), .B(opd[14]), .Z(n_24144)
		);
	notech_and3 i_123652732(.A(opc[26]), .B(\opcode[2] ), .C(n_27340), .Z(n_1622
		));
	notech_reg_set opd_reg_15(.CP(n_62692), .D(n_24151), .SD(1'b1), .Q(opd[
		15]));
	notech_mux2 i_11478(.S(n_60129), .A(n_26023), .B(opd[15]), .Z(n_24151)
		);
	notech_ao3 i_123552733(.A(opc_10[26]), .B(\opcode[2] ), .C(n_27329), .Z(n_1621
		));
	notech_reg_set opd_reg_16(.CP(n_62692), .D(n_24158), .SD(1'b1), .Q(opd[
		16]));
	notech_mux2 i_11486(.S(\nbus_11380[16] ), .A(opd[16]), .B(n_26028), .Z(n_24158
		));
	notech_nand2 i_123352735(.A(sav_esi[26]), .B(n_61136), .Z(n_1620));
	notech_reg_set opd_reg_17(.CP(n_62692), .D(n_24165), .SD(1'b1), .Q(opd[
		17]));
	notech_mux2 i_11494(.S(\nbus_11380[16] ), .A(opd[17]), .B(n_26033), .Z(n_24165
		));
	notech_reg_set opd_reg_18(.CP(n_62692), .D(n_24173), .SD(1'b1), .Q(opd[
		18]));
	notech_mux2 i_11502(.S(\nbus_11380[16] ), .A(opd[18]), .B(n_26038), .Z(n_24173
		));
	notech_reg_set opd_reg_19(.CP(n_62692), .D(n_24180), .SD(1'b1), .Q(opd[
		19]));
	notech_mux2 i_11510(.S(\nbus_11380[16] ), .A(opd[19]), .B(n_26043), .Z(n_24180
		));
	notech_reg_set opd_reg_20(.CP(n_62692), .D(n_24187), .SD(1'b1), .Q(opd[
		20]));
	notech_mux2 i_11518(.S(\nbus_11380[16] ), .A(opd[20]), .B(n_26048), .Z(n_24187
		));
	notech_reg_set opd_reg_21(.CP(n_62692), .D(n_24194), .SD(1'b1), .Q(opd[
		21]));
	notech_mux2 i_11526(.S(\nbus_11380[16] ), .A(opd[21]), .B(n_26053), .Z(n_24194
		));
	notech_reg_set opd_reg_22(.CP(n_62692), .D(n_24201), .SD(1'b1), .Q(opd[
		22]));
	notech_mux2 i_11534(.S(\nbus_11380[16] ), .A(opd[22]), .B(n_26058), .Z(n_24201
		));
	notech_reg_set opd_reg_23(.CP(n_62692), .D(n_24210), .SD(1'b1), .Q(opd[
		23]));
	notech_mux2 i_11542(.S(\nbus_11380[16] ), .A(opd[23]), .B(n_26063), .Z(n_24210
		));
	notech_reg_set opd_reg_24(.CP(n_62692), .D(n_24217), .SD(1'b1), .Q(opd[
		24]));
	notech_mux2 i_11550(.S(\nbus_11380[16] ), .A(opd[24]), .B(n_26068), .Z(n_24217
		));
	notech_nor2 i_123452734(.A(n_3983), .B(n_144428721), .Z(n_161292148));
	notech_reg_set opd_reg_25(.CP(n_62692), .D(n_24225), .SD(1'b1), .Q(opd[
		25]));
	notech_mux2 i_11558(.S(\nbus_11380[16] ), .A(opd[25]), .B(n_26073), .Z(n_24225
		));
	notech_or4 i_2821553(.A(n_178892059), .B(n_178392064), .C(n_1610), .D(n_1599
		), .Z(n_1611));
	notech_reg_set opd_reg_26(.CP(n_62692), .D(n_24233), .SD(1'b1), .Q(opd[
		26]));
	notech_mux2 i_11566(.S(\nbus_11380[16] ), .A(opd[26]), .B(n_26078), .Z(n_24233
		));
	notech_and3 i_121352755(.A(opc[27]), .B(\opcode[2] ), .C(n_27340), .Z(n_1610
		));
	notech_reg_set opd_reg_27(.CP(n_62692), .D(n_24241), .SD(1'b1), .Q(opd[
		27]));
	notech_mux2 i_11574(.S(\nbus_11380[16] ), .A(opd[27]), .B(n_26083), .Z(n_24241
		));
	notech_reg_set opd_reg_28(.CP(n_62692), .D(n_24248), .SD(1'b1), .Q(opd[
		28]));
	notech_mux2 i_11582(.S(\nbus_11380[16] ), .A(opd[28]), .B(n_26088), .Z(n_24248
		));
	notech_reg_set opd_reg_29(.CP(n_62692), .D(n_24255), .SD(1'b1), .Q(opd[
		29]));
	notech_mux2 i_11590(.S(\nbus_11380[16] ), .A(opd[29]), .B(n_26093), .Z(n_24255
		));
	notech_reg_set opd_reg_30(.CP(n_62692), .D(n_24263), .SD(1'b1), .Q(opd[
		30]));
	notech_mux2 i_11598(.S(\nbus_11380[16] ), .A(opd[30]), .B(n_26098), .Z(n_24263
		));
	notech_reg_set opd_reg_31(.CP(n_62692), .D(n_24270), .SD(1'b1), .Q(opd[
		31]));
	notech_mux2 i_11606(.S(\nbus_11380[16] ), .A(opd[31]), .B(n_27727), .Z(n_24270
		));
	notech_reg_set temp_ss_reg_0(.CP(n_62692), .D(n_24276), .SD(1'b1), .Q(temp_ss
		[0]));
	notech_mux2 i_11614(.S(\nbus_11346[0] ), .A(temp_ss[0]), .B(n_319287466)
		, .Z(n_24276));
	notech_reg_set temp_ss_reg_1(.CP(n_62606), .D(n_24282), .SD(1'b1), .Q(temp_ss
		[1]));
	notech_mux2 i_11622(.S(\nbus_11346[0] ), .A(temp_ss[1]), .B(n_319387467)
		, .Z(n_24282));
	notech_reg_set temp_ss_reg_2(.CP(n_62606), .D(n_24288), .SD(1'b1), .Q(temp_ss
		[2]));
	notech_mux2 i_11630(.S(\nbus_11346[0] ), .A(temp_ss[2]), .B(n_319487468)
		, .Z(n_24288));
	notech_reg_set temp_ss_reg_3(.CP(n_62608), .D(n_24294), .SD(1'b1), .Q(temp_ss
		[3]));
	notech_mux2 i_11638(.S(\nbus_11346[0] ), .A(temp_ss[3]), .B(n_319587469)
		, .Z(n_24294));
	notech_reg_set temp_ss_reg_4(.CP(n_62608), .D(n_24300), .SD(1'b1), .Q(temp_ss
		[4]));
	notech_mux2 i_11646(.S(\nbus_11346[0] ), .A(temp_ss[4]), .B(n_319687470)
		, .Z(n_24300));
	notech_reg_set temp_ss_reg_5(.CP(n_62608), .D(n_24306), .SD(1'b1), .Q(temp_ss
		[5]));
	notech_mux2 i_11654(.S(\nbus_11346[0] ), .A(temp_ss[5]), .B(n_319787471)
		, .Z(n_24306));
	notech_nor2 i_121252756(.A(n_4016), .B(n_144428721), .Z(n_1599));
	notech_reg_set temp_ss_reg_6(.CP(n_62608), .D(n_24312), .SD(1'b1), .Q(temp_ss
		[6]));
	notech_mux2 i_11662(.S(\nbus_11346[0] ), .A(temp_ss[6]), .B(n_319887472)
		, .Z(n_24312));
	notech_nand3 i_1221377(.A(n_177992068), .B(n_177892069), .C(n_1597), .Z(n_1598
		));
	notech_reg_set temp_ss_reg_7(.CP(n_62608), .D(n_24318), .SD(1'b1), .Q(temp_ss
		[7]));
	notech_mux2 i_11670(.S(\nbus_11346[0] ), .A(temp_ss[7]), .B(n_319987473)
		, .Z(n_24318));
	notech_or2 i_113552832(.A(n_4008), .B(n_56181), .Z(n_1597));
	notech_reg_set temp_ss_reg_8(.CP(n_62608), .D(n_24324), .SD(1'b1), .Q(temp_ss
		[8]));
	notech_mux2 i_11678(.S(\nbus_11346[0] ), .A(temp_ss[8]), .B(n_320087474)
		, .Z(n_24324));
	notech_nand2 i_113452833(.A(n_26640), .B(opd[11]), .Z(n_1596));
	notech_reg_set temp_ss_reg_9(.CP(n_62608), .D(n_24332), .SD(1'b1), .Q(temp_ss
		[9]));
	notech_mux2 i_11686(.S(\nbus_11346[0] ), .A(temp_ss[9]), .B(n_320187475)
		, .Z(n_24332));
	notech_reg_set temp_ss_reg_10(.CP(n_62608), .D(n_24338), .SD(1'b1), .Q(temp_ss
		[10]));
	notech_mux2 i_11694(.S(\nbus_11346[0] ), .A(temp_ss[10]), .B(n_320287476
		), .Z(n_24338));
	notech_reg_set temp_ss_reg_11(.CP(n_62608), .D(n_24345), .SD(1'b1), .Q(temp_ss
		[11]));
	notech_mux2 i_11702(.S(\nbus_11346[0] ), .A(temp_ss[11]), .B(n_320387477
		), .Z(n_24345));
	notech_nao3 i_113852829(.A(n_62776), .B(opc[11]), .C(n_4009), .Z(n_1593)
		);
	notech_reg_set temp_ss_reg_12(.CP(n_62608), .D(n_24351), .SD(1'b1), .Q(temp_ss
		[12]));
	notech_mux2 i_11710(.S(\nbus_11346[0] ), .A(temp_ss[12]), .B(n_320487478
		), .Z(n_24351));
	notech_nand2 i_114252825(.A(opa[11]), .B(n_1584), .Z(n_1592));
	notech_reg_set temp_ss_reg_13(.CP(n_62608), .D(n_24357), .SD(1'b1), .Q(temp_ss
		[13]));
	notech_mux2 i_11720(.S(\nbus_11346[0] ), .A(temp_ss[13]), .B(n_320587479
		), .Z(n_24357));
	notech_or2 i_113652831(.A(n_4007), .B(n_302491799), .Z(n_1591));
	notech_reg_set temp_ss_reg_14(.CP(n_62608), .D(n_24363), .SD(1'b1), .Q(temp_ss
		[14]));
	notech_mux2 i_11728(.S(\nbus_11346[0] ), .A(temp_ss[14]), .B(n_320687480
		), .Z(n_24363));
	notech_reg_set temp_ss_reg_15(.CP(n_62608), .D(n_24369), .SD(1'b1), .Q(temp_ss
		[15]));
	notech_mux2 i_11736(.S(\nbus_11346[0] ), .A(temp_ss[15]), .B(n_320787481
		), .Z(n_24369));
	notech_reg_set temp_ss_reg_16(.CP(n_62608), .D(n_24377), .SD(1'b1), .Q(temp_ss
		[16]));
	notech_mux2 i_11744(.S(n_53270), .A(temp_ss[16]), .B(n_320887482), .Z(n_24377
		));
	notech_reg_set temp_ss_reg_17(.CP(n_62608), .D(n_24383), .SD(1'b1), .Q(temp_ss
		[17]));
	notech_mux2 i_11752(.S(n_53270), .A(temp_ss[17]), .B(n_168285959), .Z(n_24383
		));
	notech_reg_set temp_ss_reg_18(.CP(n_62608), .D(n_24389), .SD(1'b1), .Q(temp_ss
		[18]));
	notech_mux2 i_11760(.S(n_53270), .A(temp_ss[18]), .B(n_320987483), .Z(n_24389
		));
	notech_reg_set temp_ss_reg_19(.CP(n_62608), .D(n_24395), .SD(1'b1), .Q(temp_ss
		[19]));
	notech_mux2 i_11768(.S(n_53270), .A(temp_ss[19]), .B(n_321087484), .Z(n_24395
		));
	notech_reg_set temp_ss_reg_20(.CP(n_62608), .D(n_24401), .SD(1'b1), .Q(temp_ss
		[20]));
	notech_mux2 i_11778(.S(n_53270), .A(temp_ss[20]), .B(n_321187485), .Z(n_24401
		));
	notech_nao3 i_3353879(.A(n_27257), .B(n_27272), .C(n_1580), .Z(n_1584)
		);
	notech_reg_set temp_ss_reg_21(.CP(n_62608), .D(n_24407), .SD(1'b1), .Q(temp_ss
		[21]));
	notech_mux2 i_11786(.S(n_53270), .A(temp_ss[21]), .B(n_321287486), .Z(n_24407
		));
	notech_ao4 i_3453878(.A(n_56959), .B(n_4005), .C(n_55735), .D(n_306991754
		), .Z(n_1583));
	notech_reg_set temp_ss_reg_22(.CP(n_62538), .D(n_24413), .SD(1'b1), .Q(temp_ss
		[22]));
	notech_mux2 i_11794(.S(n_53270), .A(temp_ss[22]), .B(n_321387487), .Z(n_24413
		));
	notech_reg_set temp_ss_reg_23(.CP(n_62538), .D(n_24419), .SD(1'b1), .Q(temp_ss
		[23]));
	notech_mux2 i_11802(.S(n_53270), .A(temp_ss[23]), .B(n_321487488), .Z(n_24419
		));
	notech_reg_set temp_ss_reg_24(.CP(n_62538), .D(n_24425), .SD(1'b1), .Q(temp_ss
		[24]));
	notech_mux2 i_11810(.S(n_53270), .A(temp_ss[24]), .B(n_321587489), .Z(n_24425
		));
	notech_ao4 i_112952838(.A(n_56950), .B(n_26626), .C(n_311591708), .D(n_306191762
		), .Z(n_1580));
	notech_reg_set temp_ss_reg_25(.CP(n_62538), .D(n_24432), .SD(1'b1), .Q(temp_ss
		[25]));
	notech_mux2 i_11818(.S(n_53270), .A(temp_ss[25]), .B(n_321687490), .Z(n_24432
		));
	notech_reg_set temp_ss_reg_26(.CP(n_62538), .D(n_24439), .SD(1'b1), .Q(temp_ss
		[26]));
	notech_mux2 i_11826(.S(n_53270), .A(temp_ss[26]), .B(n_321787491), .Z(n_24439
		));
	notech_reg_set temp_ss_reg_27(.CP(n_62538), .D(n_24446), .SD(1'b1), .Q(temp_ss
		[27]));
	notech_mux2 i_11834(.S(n_53270), .A(temp_ss[27]), .B(n_321887492), .Z(n_24446
		));
	notech_or4 i_3021395(.A(n_1575), .B(n_1767), .C(n_1576), .D(n_1568), .Z(n_1577
		));
	notech_reg_set temp_ss_reg_28(.CP(n_62538), .D(n_24453), .SD(1'b1), .Q(temp_ss
		[28]));
	notech_mux2 i_11842(.S(n_53270), .A(temp_ss[28]), .B(n_321987493), .Z(n_24453
		));
	notech_and3 i_105052916(.A(opc[29]), .B(\opcode[2] ), .C(n_4010), .Z(n_1576
		));
	notech_reg_set temp_ss_reg_29(.CP(n_62538), .D(n_24461), .SD(1'b1), .Q(temp_ss
		[29]));
	notech_mux2 i_11850(.S(n_53270), .A(temp_ss[29]), .B(n_322087494), .Z(n_24461
		));
	notech_ao3 i_104952917(.A(opc_10[29]), .B(\opcode[2] ), .C(n_295269964),
		 .Z(n_1575));
	notech_reg_set temp_ss_reg_30(.CP(n_62538), .D(n_24468), .SD(1'b1), .Q(temp_ss
		[30]));
	notech_mux2 i_11858(.S(n_53270), .A(temp_ss[30]), .B(n_322187495), .Z(n_24468
		));
	notech_reg_set temp_ss_reg_31(.CP(n_62688), .D(n_24475), .SD(1'b1), .Q(temp_ss
		[31]));
	notech_mux2 i_11866(.S(n_53270), .A(temp_ss[31]), .B(n_322287496), .Z(n_24475
		));
	notech_reg errco_reg_0(.CP(n_62596), .D(n_24482), .CD(n_61526), .Q(errco
		[0]));
	notech_mux2 i_11874(.S(n_55016), .A(errco[0]), .B(n_24991034), .Z(n_24482
		));
	notech_reg errco_reg_1(.CP(n_62536), .D(n_24489), .CD(n_61526), .Q(errco
		[1]));
	notech_mux2 i_11882(.S(n_55016), .A(errco[1]), .B(wr_fault), .Z(n_24489)
		);
	notech_reg errco_reg_2(.CP(n_62596), .D(n_24497), .CD(n_61526), .Q(errco
		[2]));
	notech_mux2 i_11890(.S(n_55016), .A(errco[2]), .B(cs[1]), .Z(n_24497));
	notech_reg errco_reg_3(.CP(n_62596), .D(n_24507), .CD(n_61525), .Q(errco
		[3]));
	notech_ao3 i_11900(.A(n_60139), .B(errco[3]), .C(n_60765), .Z(n_24507)
		);
	notech_reg errco_reg_4(.CP(n_62596), .D(n_24511), .CD(n_61525), .Q(errco
		[4]));
	notech_mux2 i_11906(.S(n_55016), .A(errco[4]), .B(n_60765), .Z(n_24511)
		);
	notech_nor2 i_104852918(.A(n_3981), .B(n_309891725), .Z(n_1568));
	notech_reg errco_reg_5(.CP(n_62596), .D(n_24522), .CD(n_61525), .Q(errco
		[5]));
	notech_ao3 i_11916(.A(n_60139), .B(errco[5]), .C(n_60765), .Z(n_24522)
		);
	notech_and2 i_3753875(.A(n_176192078), .B(n_1562), .Z(n_1567));
	notech_reg errco_reg_6(.CP(n_62596), .D(n_24529), .CD(n_61525), .Q(errco
		[6]));
	notech_ao3 i_11924(.A(n_60139), .B(errco[6]), .C(n_60773), .Z(n_24529)
		);
	notech_reg errco_reg_7(.CP(n_62596), .D(n_24536), .CD(n_61525), .Q(errco
		[7]));
	notech_ao3 i_11933(.A(n_60139), .B(errco[7]), .C(n_60765), .Z(n_24536)
		);
	notech_reg errco_reg_8(.CP(n_62596), .D(n_24543), .CD(n_61526), .Q(errco
		[8]));
	notech_ao3 i_11943(.A(n_60139), .B(errco[8]), .C(n_60765), .Z(n_24543)
		);
	notech_reg errco_reg_9(.CP(n_62596), .D(n_24551), .CD(n_61526), .Q(errco
		[9]));
	notech_ao3 i_11951(.A(n_60139), .B(errco[9]), .C(n_60765), .Z(n_24551)
		);
	notech_reg errco_reg_10(.CP(n_62596), .D(n_24558), .CD(n_61525), .Q(errco
		[10]));
	notech_ao3 i_11959(.A(n_60139), .B(errco[10]), .C(n_60765), .Z(n_24558)
		);
	notech_or2 i_103352933(.A(n_56959), .B(opa[7]), .Z(n_1562));
	notech_reg errco_reg_11(.CP(n_62680), .D(n_24565), .CD(n_61526), .Q(errco
		[11]));
	notech_ao3 i_11967(.A(n_60139), .B(errco[11]), .C(n_60765), .Z(n_24565)
		);
	notech_or4 i_2721360(.A(n_1559), .B(n_175792081), .C(n_1560), .D(n_1549)
		, .Z(n_1561));
	notech_reg errco_reg_12(.CP(n_62680), .D(n_24572), .CD(n_61527), .Q(errco
		[12]));
	notech_ao3 i_11975(.A(n_60139), .B(errco[12]), .C(n_60765), .Z(n_24572)
		);
	notech_and3 i_91153052(.A(opc[26]), .B(\opcode[2] ), .C(n_309791726), .Z
		(n_1560));
	notech_reg errco_reg_13(.CP(n_62680), .D(n_24579), .CD(n_61528), .Q(errco
		[13]));
	notech_ao3 i_11983(.A(n_60128), .B(errco[13]), .C(n_60765), .Z(n_24579)
		);
	notech_ao3 i_91053053(.A(opc_10[26]), .B(\opcode[2] ), .C(n_309691727), 
		.Z(n_1559));
	notech_reg errco_reg_14(.CP(n_62680), .D(n_24591), .CD(n_61527), .Q(errco
		[14]));
	notech_ao3 i_11991(.A(n_60128), .B(errco[14]), .C(n_60765), .Z(n_24591)
		);
	notech_nand2 i_90853055(.A(sav_edi[26]), .B(n_61136), .Z(n_1558));
	notech_reg errco_reg_15(.CP(n_62680), .D(n_24600), .CD(n_61527), .Q(errco
		[15]));
	notech_ao3 i_11999(.A(n_60128), .B(errco[15]), .C(n_60765), .Z(n_24600)
		);
	notech_reg errco_reg_16(.CP(n_62680), .D(n_24607), .CD(n_61528), .Q(errco
		[16]));
	notech_ao3 i_12007(.A(n_60128), .B(errco[16]), .C(n_60765), .Z(n_24607)
		);
	notech_reg errco_reg_17(.CP(n_62680), .D(n_24615), .CD(n_61528), .Q(errco
		[17]));
	notech_ao3 i_12015(.A(n_60128), .B(errco[17]), .C(n_60773), .Z(n_24615)
		);
	notech_reg errco_reg_18(.CP(n_62680), .D(n_24622), .CD(n_61528), .Q(errco
		[18]));
	notech_ao3 i_12023(.A(n_60128), .B(errco[18]), .C(n_60769), .Z(n_24622)
		);
	notech_reg errco_reg_19(.CP(n_62680), .D(n_24628), .CD(n_61528), .Q(errco
		[19]));
	notech_ao3 i_12032(.A(n_60128), .B(errco[19]), .C(n_60769), .Z(n_24628)
		);
	notech_reg errco_reg_20(.CP(n_62680), .D(n_24635), .CD(n_61528), .Q(errco
		[20]));
	notech_ao3 i_12040(.A(n_60128), .B(errco[20]), .C(n_60769), .Z(n_24635)
		);
	notech_reg errco_reg_21(.CP(n_62680), .D(n_24641), .CD(n_61527), .Q(errco
		[21]));
	notech_ao3 i_12048(.A(n_60127), .B(errco[21]), .C(n_60769), .Z(n_24641)
		);
	notech_reg errco_reg_22(.CP(n_62680), .D(n_24647), .CD(n_61527), .Q(errco
		[22]));
	notech_ao3 i_12056(.A(n_60127), .B(errco[22]), .C(n_60769), .Z(n_24647)
		);
	notech_reg errco_reg_23(.CP(n_62680), .D(n_24653), .CD(n_61527), .Q(errco
		[23]));
	notech_ao3 i_12064(.A(n_60127), .B(errco[23]), .C(n_60769), .Z(n_24653)
		);
	notech_nor2 i_90953054(.A(n_139728674), .B(n_3983), .Z(n_1549));
	notech_reg errco_reg_24(.CP(n_62680), .D(n_24659), .CD(n_61527), .Q(errco
		[24]));
	notech_ao3 i_12072(.A(n_60127), .B(errco[24]), .C(n_60769), .Z(n_24659)
		);
	notech_reg errco_reg_25(.CP(n_62680), .D(n_24665), .CD(n_61527), .Q(errco
		[25]));
	notech_ao3 i_12080(.A(n_60128), .B(errco[25]), .C(n_60769), .Z(n_24665)
		);
	notech_reg errco_reg_26(.CP(n_62680), .D(n_24671), .CD(n_61527), .Q(errco
		[26]));
	notech_ao3 i_12088(.A(n_60128), .B(errco[26]), .C(n_60773), .Z(n_24671)
		);
	notech_reg errco_reg_27(.CP(n_62680), .D(n_24677), .CD(n_61527), .Q(errco
		[27]));
	notech_ao3 i_12096(.A(n_60128), .B(errco[27]), .C(n_60773), .Z(n_24677)
		);
	notech_reg errco_reg_28(.CP(n_62680), .D(n_24683), .CD(n_61527), .Q(errco
		[28]));
	notech_ao3 i_12104(.A(n_60128), .B(errco[28]), .C(n_60773), .Z(n_24683)
		);
	notech_reg errco_reg_29(.CP(n_62680), .D(n_24690), .CD(n_61527), .Q(errco
		[29]));
	notech_ao3 i_12112(.A(n_60133), .B(errco[29]), .C(n_60773), .Z(n_24690)
		);
	notech_reg errco_reg_30(.CP(n_62678), .D(n_24696), .CD(n_61527), .Q(errco
		[30]));
	notech_ao3 i_12120(.A(n_60133), .B(errco[30]), .C(n_60769), .Z(n_24696)
		);
	notech_reg errco_reg_31(.CP(n_62678), .D(n_24702), .CD(n_61521), .Q(errco
		[31]));
	notech_ao3 i_12128(.A(n_60133), .B(errco[31]), .C(n_60769), .Z(n_24702)
		);
	notech_reg_set write_data_reg_0(.CP(n_62740), .D(n_24706), .SD(1'b1), .Q
		(write_data[0]));
	notech_mux2 i_12134(.S(\nbus_11378[0] ), .A(write_data[0]), .B(n_25704),
		 .Z(n_24706));
	notech_reg_set write_data_reg_1(.CP(n_62740), .D(n_24715), .SD(1'b1), .Q
		(write_data[1]));
	notech_mux2 i_12142(.S(\nbus_11378[0] ), .A(write_data[1]), .B(n_25709),
		 .Z(n_24715));
	notech_reg_set write_data_reg_2(.CP(n_62740), .D(n_24721), .SD(1'b1), .Q
		(write_data[2]));
	notech_mux2 i_12150(.S(\nbus_11378[0] ), .A(write_data[2]), .B(n_25714),
		 .Z(n_24721));
	notech_reg_set write_data_reg_3(.CP(n_62740), .D(n_24727), .SD(1'b1), .Q
		(write_data[3]));
	notech_mux2 i_12158(.S(\nbus_11378[0] ), .A(write_data[3]), .B(n_25719),
		 .Z(n_24727));
	notech_reg_set write_data_reg_4(.CP(n_62740), .D(n_24733), .SD(1'b1), .Q
		(write_data[4]));
	notech_mux2 i_12166(.S(\nbus_11378[0] ), .A(write_data[4]), .B(n_25724),
		 .Z(n_24733));
	notech_reg_set write_data_reg_5(.CP(n_62740), .D(n_24739), .SD(1'b1), .Q
		(write_data[5]));
	notech_mux2 i_12174(.S(\nbus_11378[0] ), .A(write_data[5]), .B(n_25729),
		 .Z(n_24739));
	notech_reg_set write_data_reg_6(.CP(n_62740), .D(n_24745), .SD(1'b1), .Q
		(write_data[6]));
	notech_mux2 i_12182(.S(\nbus_11378[0] ), .A(write_data[6]), .B(n_25734),
		 .Z(n_24745));
	notech_reg_set write_data_reg_7(.CP(n_62740), .D(n_24751), .SD(1'b1), .Q
		(write_data[7]));
	notech_mux2 i_12190(.S(\nbus_11378[0] ), .A(write_data[7]), .B(n_25739),
		 .Z(n_24751));
	notech_reg_set write_data_reg_8(.CP(n_62740), .D(n_24758), .SD(1'b1), .Q
		(write_data[8]));
	notech_mux2 i_12198(.S(\nbus_11378[0] ), .A(write_data[8]), .B(n_25744),
		 .Z(n_24758));
	notech_reg_set write_data_reg_9(.CP(n_62740), .D(n_24765), .SD(1'b1), .Q
		(write_data[9]));
	notech_mux2 i_12207(.S(\nbus_11378[0] ), .A(write_data[9]), .B(n_25749),
		 .Z(n_24765));
	notech_reg_set write_data_reg_10(.CP(n_62740), .D(n_24772), .SD(1'b1), .Q
		(write_data[10]));
	notech_mux2 i_12215(.S(\nbus_11378[0] ), .A(write_data[10]), .B(n_25754)
		, .Z(n_24772));
	notech_reg_set write_data_reg_11(.CP(n_62448), .D(n_24779), .SD(1'b1), .Q
		(write_data[11]));
	notech_mux2 i_12223(.S(\nbus_11378[0] ), .A(write_data[11]), .B(n_25759)
		, .Z(n_24779));
	notech_reg_set write_data_reg_12(.CP(n_62740), .D(n_24787), .SD(1'b1), .Q
		(write_data[12]));
	notech_mux2 i_12231(.S(\nbus_11378[0] ), .A(write_data[12]), .B(n_25764)
		, .Z(n_24787));
	notech_reg_set write_data_reg_13(.CP(n_62740), .D(n_24794), .SD(1'b1), .Q
		(write_data[13]));
	notech_mux2 i_12239(.S(\nbus_11378[0] ), .A(write_data[13]), .B(n_25769)
		, .Z(n_24794));
	notech_reg_set write_data_reg_14(.CP(n_62740), .D(n_24801), .SD(1'b1), .Q
		(write_data[14]));
	notech_mux2 i_12247(.S(\nbus_11378[0] ), .A(write_data[14]), .B(n_25774)
		, .Z(n_24801));
	notech_reg_set write_data_reg_15(.CP(n_62740), .D(n_24811), .SD(1'b1), .Q
		(write_data[15]));
	notech_mux2 i_12256(.S(\nbus_11378[0] ), .A(write_data[15]), .B(n_25779)
		, .Z(n_24811));
	notech_reg_set write_data_reg_16(.CP(n_62740), .D(n_24818), .SD(1'b1), .Q
		(write_data[16]));
	notech_mux2 i_12264(.S(n_54146), .A(write_data[16]), .B(n_25784), .Z(n_24818
		));
	notech_reg_set write_data_reg_17(.CP(n_62740), .D(n_24825), .SD(1'b1), .Q
		(write_data[17]));
	notech_mux2 i_12272(.S(n_54146), .A(write_data[17]), .B(n_25789), .Z(n_24825
		));
	notech_reg_set write_data_reg_18(.CP(n_62678), .D(n_24832), .SD(1'b1), .Q
		(write_data[18]));
	notech_mux2 i_12280(.S(n_54146), .A(write_data[18]), .B(n_25794), .Z(n_24832
		));
	notech_reg_set write_data_reg_19(.CP(n_62678), .D(n_24839), .SD(1'b1), .Q
		(write_data[19]));
	notech_mux2 i_12289(.S(n_54146), .A(write_data[19]), .B(n_25799), .Z(n_24839
		));
	notech_reg_set write_data_reg_20(.CP(n_62678), .D(n_24847), .SD(1'b1), .Q
		(write_data[20]));
	notech_mux2 i_12297(.S(n_54146), .A(write_data[20]), .B(n_25804), .Z(n_24847
		));
	notech_reg_set write_data_reg_21(.CP(n_62678), .D(n_24854), .SD(1'b1), .Q
		(write_data[21]));
	notech_mux2 i_12305(.S(n_54146), .A(write_data[21]), .B(n_25809), .Z(n_24854
		));
	notech_reg_set write_data_reg_22(.CP(n_62678), .D(n_24861), .SD(1'b1), .Q
		(write_data[22]));
	notech_mux2 i_12313(.S(n_54146), .A(write_data[22]), .B(n_25814), .Z(n_24861
		));
	notech_reg_set write_data_reg_23(.CP(n_62678), .D(n_24868), .SD(1'b1), .Q
		(write_data[23]));
	notech_mux2 i_12321(.S(n_54146), .A(write_data[23]), .B(n_25819), .Z(n_24868
		));
	notech_reg_set write_data_reg_24(.CP(n_62678), .D(n_24875), .SD(1'b1), .Q
		(write_data[24]));
	notech_mux2 i_12329(.S(n_54146), .A(write_data[24]), .B(n_25824), .Z(n_24875
		));
	notech_reg_set write_data_reg_25(.CP(n_62678), .D(n_24883), .SD(1'b1), .Q
		(write_data[25]));
	notech_mux2 i_12338(.S(n_54146), .A(write_data[25]), .B(n_25829), .Z(n_24883
		));
	notech_reg_set write_data_reg_26(.CP(n_62678), .D(n_24890), .SD(1'b1), .Q
		(write_data[26]));
	notech_mux2 i_12346(.S(n_54146), .A(write_data[26]), .B(n_25834), .Z(n_24890
		));
	notech_reg_set write_data_reg_27(.CP(n_62740), .D(n_24897), .SD(1'b1), .Q
		(write_data[27]));
	notech_mux2 i_12354(.S(n_54146), .A(write_data[27]), .B(n_25839), .Z(n_24897
		));
	notech_reg_set write_data_reg_28(.CP(n_62736), .D(n_24904), .SD(1'b1), .Q
		(write_data[28]));
	notech_mux2 i_12362(.S(n_54146), .A(write_data[28]), .B(n_25844), .Z(n_24904
		));
	notech_or4 i_3020723(.A(n_1510), .B(n_171092121), .C(n_1511), .D(n_1500)
		, .Z(n_1512));
	notech_reg_set write_data_reg_29(.CP(n_62676), .D(n_24911), .SD(1'b1), .Q
		(write_data[29]));
	notech_mux2 i_12370(.S(n_54146), .A(write_data[29]), .B(n_25849), .Z(n_24911
		));
	notech_ao3 i_24753694(.A(opc[29]), .B(\opcode[2] ), .C(n_309391730), .Z(n_1511
		));
	notech_reg_set write_data_reg_30(.CP(n_62736), .D(n_24919), .SD(1'b1), .Q
		(write_data[30]));
	notech_mux2 i_12378(.S(n_54146), .A(write_data[30]), .B(n_25854), .Z(n_24919
		));
	notech_and2 i_24353696(.A(add_len_pc[29]), .B(n_26766), .Z(n_1510));
	notech_reg_set write_data_reg_31(.CP(n_62736), .D(n_24926), .SD(1'b1), .Q
		(write_data[31]));
	notech_mux2 i_12386(.S(n_54146), .A(write_data[31]), .B(n_25859), .Z(n_24926
		));
	notech_nand2 i_24253697(.A(sav_epc[29]), .B(n_61136), .Z(n_1509));
	notech_reg ldtr_reg_0(.CP(n_62736), .D(n_24933), .CD(n_61521), .Q(ldtr[0
		]));
	notech_mux2 i_12394(.S(n_327990777), .A(opb[0]), .B(ldtr[0]), .Z(n_24933
		));
	notech_reg ldtr_reg_1(.CP(n_62736), .D(n_24940), .CD(n_61521), .Q(ldtr[1
		]));
	notech_mux2 i_12402(.S(n_327990777), .A(opb[1]), .B(ldtr[1]), .Z(n_24940
		));
	notech_reg ldtr_reg_2(.CP(n_62736), .D(n_24947), .CD(n_61521), .Q(ldtr[2
		]));
	notech_mux2 i_12410(.S(n_327990777), .A(opb[2]), .B(ldtr[2]), .Z(n_24947
		));
	notech_reg ldtr_reg_3(.CP(n_62736), .D(n_24953), .CD(n_61521), .Q(ldtr[3
		]));
	notech_mux2 i_12418(.S(n_327990777), .A(opb[3]), .B(ldtr[3]), .Z(n_24953
		));
	notech_reg ldtr_reg_4(.CP(n_62736), .D(n_24959), .CD(n_61521), .Q(ldtr[4
		]));
	notech_mux2 i_12426(.S(n_327990777), .A(opb[4]), .B(ldtr[4]), .Z(n_24959
		));
	notech_reg ldtr_reg_5(.CP(n_62736), .D(n_24965), .CD(n_61522), .Q(ldtr[5
		]));
	notech_mux2 i_12434(.S(n_327990777), .A(opb[5]), .B(ldtr[5]), .Z(n_24965
		));
	notech_reg ldtr_reg_6(.CP(n_62736), .D(n_24971), .CD(n_61521), .Q(ldtr[6
		]));
	notech_mux2 i_12442(.S(n_327990777), .A(opb[6]), .B(ldtr[6]), .Z(n_24971
		));
	notech_reg ldtr_reg_7(.CP(n_62736), .D(n_24977), .CD(n_61521), .Q(ldtr[7
		]));
	notech_mux2 i_12450(.S(n_327990777), .A(opb[7]), .B(ldtr[7]), .Z(n_24977
		));
	notech_reg ldtr_reg_8(.CP(n_62760), .D(n_24983), .CD(n_61521), .Q(ldtr[8
		]));
	notech_mux2 i_12458(.S(n_327990777), .A(opb[8]), .B(ldtr[8]), .Z(n_24983
		));
	notech_nor2 i_24553695(.A(n_124328520), .B(n_3981), .Z(n_1500));
	notech_reg ldtr_reg_9(.CP(n_62760), .D(n_24990), .CD(n_61520), .Q(ldtr[9
		]));
	notech_mux2 i_12466(.S(n_327990777), .A(opb[9]), .B(ldtr[9]), .Z(n_24990
		));
	notech_reg ldtr_reg_10(.CP(n_62760), .D(n_24999), .CD(n_61520), .Q(ldtr[
		10]));
	notech_mux2 i_12474(.S(n_327990777), .A(opb[10]), .B(ldtr[10]), .Z(n_24999
		));
	notech_reg ldtr_reg_11(.CP(n_62760), .D(n_25006), .CD(n_61520), .Q(ldtr[
		11]));
	notech_mux2 i_12482(.S(n_327990777), .A(opb[11]), .B(ldtr[11]), .Z(n_25006
		));
	notech_reg ldtr_reg_12(.CP(n_62760), .D(n_25014), .CD(n_61520), .Q(ldtr[
		12]));
	notech_mux2 i_12490(.S(n_327990777), .A(opb[12]), .B(ldtr[12]), .Z(n_25014
		));
	notech_reg ldtr_reg_13(.CP(n_62760), .D(n_25020), .CD(n_61520), .Q(ldtr[
		13]));
	notech_mux2 i_12498(.S(n_327990777), .A(opb[13]), .B(ldtr[13]), .Z(n_25020
		));
	notech_reg ldtr_reg_14(.CP(n_62760), .D(n_25026), .CD(n_61521), .Q(ldtr[
		14]));
	notech_mux2 i_12506(.S(n_327990777), .A(opb[14]), .B(ldtr[14]), .Z(n_25026
		));
	notech_reg ldtr_reg_15(.CP(n_62760), .D(n_25032), .CD(n_61521), .Q(ldtr[
		15]));
	notech_mux2 i_12514(.S(n_327990777), .A(opb[15]), .B(ldtr[15]), .Z(n_25032
		));
	notech_reg ldtr_reg_16(.CP(n_62760), .D(n_25038), .CD(n_61521), .Q(ldtr[
		16]));
	notech_mux2 i_12522(.S(n_54378), .A(opb[16]), .B(ldtr[16]), .Z(n_25038)
		);
	notech_reg ldtr_reg_17(.CP(n_62760), .D(n_25044), .CD(n_61521), .Q(ldtr[
		17]));
	notech_mux2 i_12530(.S(n_54378), .A(opb[17]), .B(ldtr[17]), .Z(n_25044)
		);
	notech_reg ldtr_reg_18(.CP(n_62760), .D(n_25050), .CD(n_61525), .Q(ldtr[
		18]));
	notech_mux2 i_12538(.S(n_54378), .A(opb[18]), .B(ldtr[18]), .Z(n_25050)
		);
	notech_reg ldtr_reg_19(.CP(n_62760), .D(n_25056), .CD(n_61525), .Q(ldtr[
		19]));
	notech_mux2 i_12549(.S(n_54378), .A(opb[19]), .B(ldtr[19]), .Z(n_25056)
		);
	notech_reg ldtr_reg_20(.CP(n_62760), .D(n_25062), .CD(n_61522), .Q(ldtr[
		20]));
	notech_mux2 i_12557(.S(n_54378), .A(opb[20]), .B(ldtr[20]), .Z(n_25062)
		);
	notech_reg ldtr_reg_21(.CP(n_62760), .D(n_25068), .CD(n_61522), .Q(ldtr[
		21]));
	notech_mux2 i_12565(.S(n_54378), .A(opb[21]), .B(ldtr[21]), .Z(n_25068)
		);
	notech_reg ldtr_reg_22(.CP(n_62760), .D(n_25074), .CD(n_61525), .Q(ldtr[
		22]));
	notech_mux2 i_12573(.S(n_54378), .A(opb[22]), .B(ldtr[22]), .Z(n_25074)
		);
	notech_reg ldtr_reg_23(.CP(n_62760), .D(n_25080), .CD(n_61525), .Q(ldtr[
		23]));
	notech_mux2 i_12581(.S(n_54378), .A(opb[23]), .B(ldtr[23]), .Z(n_25080)
		);
	notech_reg ldtr_reg_24(.CP(n_62760), .D(n_25086), .CD(n_61525), .Q(ldtr[
		24]));
	notech_mux2 i_12589(.S(n_54378), .A(opb[24]), .B(ldtr[24]), .Z(n_25086)
		);
	notech_reg ldtr_reg_25(.CP(n_62760), .D(n_25092), .CD(n_61525), .Q(ldtr[
		25]));
	notech_mux2 i_12597(.S(n_54378), .A(opb[25]), .B(ldtr[25]), .Z(n_25092)
		);
	notech_reg ldtr_reg_26(.CP(n_62736), .D(n_25098), .CD(n_61525), .Q(ldtr[
		26]));
	notech_mux2 i_12605(.S(n_54378), .A(opb[26]), .B(ldtr[26]), .Z(n_25098)
		);
	notech_reg ldtr_reg_27(.CP(n_62760), .D(n_25104), .CD(n_61522), .Q(ldtr[
		27]));
	notech_mux2 i_12613(.S(n_54378), .A(opb[27]), .B(ldtr[27]), .Z(n_25104)
		);
	notech_reg ldtr_reg_28(.CP(n_62738), .D(n_25110), .CD(n_61522), .Q(ldtr[
		28]));
	notech_mux2 i_12621(.S(n_54378), .A(opb[28]), .B(ldtr[28]), .Z(n_25110)
		);
	notech_reg ldtr_reg_29(.CP(n_62738), .D(n_25116), .CD(n_61522), .Q(ldtr[
		29]));
	notech_mux2 i_12629(.S(n_54378), .A(opb[29]), .B(ldtr[29]), .Z(n_25116)
		);
	notech_or2 i_18453751(.A(n_56959), .B(n_57957), .Z(n_1479));
	notech_reg ldtr_reg_30(.CP(n_62738), .D(n_25122), .CD(n_61522), .Q(ldtr[
		30]));
	notech_mux2 i_12637(.S(n_54378), .A(opb[30]), .B(ldtr[30]), .Z(n_25122)
		);
	notech_or4 i_18053755(.A(n_2868), .B(\opcode[2] ), .C(n_60904), .D(n_60207
		), .Z(n_1478));
	notech_reg ldtr_reg_31(.CP(n_62738), .D(n_25128), .CD(n_61522), .Q(ldtr[
		31]));
	notech_mux2 i_12645(.S(n_54378), .A(opb[31]), .B(ldtr[31]), .Z(n_25128)
		);
	notech_reg gdtr_reg_0(.CP(n_62738), .D(n_25134), .CD(n_61522), .Q(gdtr[0
		]));
	notech_mux2 i_12653(.S(n_327890776), .A(opb[0]), .B(gdtr[0]), .Z(n_25134
		));
	notech_or4 i_108755516(.A(n_61175), .B(n_61160), .C(n_61151), .D(eval_flag
		), .Z(n_27754));
	notech_reg gdtr_reg_1(.CP(n_62738), .D(n_25140), .CD(n_61522), .Q(gdtr[1
		]));
	notech_mux2 i_12661(.S(n_327890776), .A(opb[1]), .B(gdtr[1]), .Z(n_25140
		));
	notech_ao4 i_46853981(.A(n_1903), .B(n_1901), .C(n_56950), .D(n_26626), 
		.Z(n_1476));
	notech_reg gdtr_reg_2(.CP(n_62738), .D(n_25146), .CD(n_61522), .Q(gdtr[2
		]));
	notech_mux2 i_12669(.S(n_327890776), .A(opb[2]), .B(gdtr[2]), .Z(n_25146
		));
	notech_nand3 i_12653787(.A(n_1476), .B(n_27377), .C(n_60321), .Z(n_1475)
		);
	notech_reg gdtr_reg_3(.CP(n_62738), .D(n_25152), .CD(n_61522), .Q(gdtr[3
		]));
	notech_mux2 i_12677(.S(n_327890776), .A(opb[3]), .B(gdtr[3]), .Z(n_25152
		));
	notech_nao3 i_12453789(.A(n_246591944), .B(n_57068), .C(n_306591758), .Z
		(n_1474));
	notech_reg gdtr_reg_4(.CP(n_62738), .D(n_25158), .CD(n_61522), .Q(gdtr[4
		]));
	notech_mux2 i_12685(.S(n_327890776), .A(opb[4]), .B(gdtr[4]), .Z(n_25158
		));
	notech_or2 i_10553807(.A(n_4011), .B(n_56518), .Z(n_1473));
	notech_reg gdtr_reg_5(.CP(n_62738), .D(n_25164), .CD(n_61533), .Q(gdtr[5
		]));
	notech_mux2 i_12693(.S(n_327890776), .A(opb[5]), .B(gdtr[5]), .Z(n_25164
		));
	notech_reg gdtr_reg_6(.CP(n_62738), .D(n_25170), .CD(n_61533), .Q(gdtr[6
		]));
	notech_mux2 i_12701(.S(n_327890776), .A(opb[6]), .B(gdtr[6]), .Z(n_25170
		));
	notech_reg gdtr_reg_7(.CP(n_62738), .D(n_25176), .CD(n_61533), .Q(gdtr[7
		]));
	notech_mux2 i_12709(.S(n_327890776), .A(opb[7]), .B(gdtr[7]), .Z(n_25176
		));
	notech_reg gdtr_reg_8(.CP(n_62738), .D(n_25182), .CD(n_61533), .Q(gdtr[8
		]));
	notech_mux2 i_12717(.S(n_327890776), .A(opb[8]), .B(gdtr[8]), .Z(n_25182
		));
	notech_reg gdtr_reg_9(.CP(n_62738), .D(n_25188), .CD(n_61533), .Q(gdtr[9
		]));
	notech_mux2 i_12725(.S(n_327890776), .A(opb[9]), .B(gdtr[9]), .Z(n_25188
		));
	notech_reg gdtr_reg_10(.CP(n_62738), .D(n_25194), .CD(n_61533), .Q(gdtr[
		10]));
	notech_mux2 i_12733(.S(n_327890776), .A(opb[10]), .B(gdtr[10]), .Z(n_25194
		));
	notech_reg gdtr_reg_11(.CP(n_62738), .D(n_25200), .CD(n_61533), .Q(gdtr[
		11]));
	notech_mux2 i_12741(.S(n_327890776), .A(opb[11]), .B(gdtr[11]), .Z(n_25200
		));
	notech_reg gdtr_reg_12(.CP(n_62738), .D(n_25206), .CD(n_61533), .Q(gdtr[
		12]));
	notech_mux2 i_12749(.S(n_327890776), .A(opb[12]), .B(gdtr[12]), .Z(n_25206
		));
	notech_reg gdtr_reg_13(.CP(n_62738), .D(n_25212), .CD(n_61533), .Q(gdtr[
		13]));
	notech_mux2 i_12757(.S(n_327890776), .A(opb[13]), .B(gdtr[13]), .Z(n_25212
		));
	notech_reg gdtr_reg_14(.CP(n_62738), .D(n_25218), .CD(n_61533), .Q(gdtr[
		14]));
	notech_mux2 i_12765(.S(n_327890776), .A(opb[14]), .B(gdtr[14]), .Z(n_25218
		));
	notech_reg gdtr_reg_15(.CP(n_62676), .D(n_25224), .CD(n_61532), .Q(gdtr[
		15]));
	notech_mux2 i_12773(.S(n_327890776), .A(opb[15]), .B(gdtr[15]), .Z(n_25224
		));
	notech_reg gdtr_reg_16(.CP(n_62676), .D(n_25230), .CD(n_61532), .Q(gdtr[
		16]));
	notech_mux2 i_12781(.S(n_54535), .A(opb[16]), .B(gdtr[16]), .Z(n_25230)
		);
	notech_reg gdtr_reg_17(.CP(n_62676), .D(n_25236), .CD(n_61532), .Q(gdtr[
		17]));
	notech_mux2 i_12789(.S(n_54535), .A(opb[17]), .B(gdtr[17]), .Z(n_25236)
		);
	notech_reg gdtr_reg_18(.CP(n_62676), .D(n_25242), .CD(n_61532), .Q(gdtr[
		18]));
	notech_mux2 i_12797(.S(n_54535), .A(opb[18]), .B(gdtr[18]), .Z(n_25242)
		);
	notech_reg gdtr_reg_19(.CP(n_62676), .D(n_25249), .CD(n_61532), .Q(gdtr[
		19]));
	notech_mux2 i_12805(.S(n_54535), .A(opb[19]), .B(gdtr[19]), .Z(n_25249)
		);
	notech_reg gdtr_reg_20(.CP(n_62676), .D(n_25256), .CD(n_61532), .Q(gdtr[
		20]));
	notech_mux2 i_12813(.S(n_54535), .A(opb[20]), .B(gdtr[20]), .Z(n_25256)
		);
	notech_reg gdtr_reg_21(.CP(n_62676), .D(n_25263), .CD(n_61533), .Q(gdtr[
		21]));
	notech_mux2 i_12821(.S(n_54535), .A(opb[21]), .B(gdtr[21]), .Z(n_25263)
		);
	notech_reg gdtr_reg_22(.CP(n_62676), .D(n_25271), .CD(n_61532), .Q(gdtr[
		22]));
	notech_mux2 i_12829(.S(n_54535), .A(opb[22]), .B(gdtr[22]), .Z(n_25271)
		);
	notech_or4 i_29157(.A(n_61175), .B(n_61160), .C(n_61151), .D(n_59708), .Z
		(n_30818));
	notech_reg gdtr_reg_23(.CP(n_62676), .D(n_25278), .CD(n_61532), .Q(gdtr[
		23]));
	notech_mux2 i_12837(.S(n_54535), .A(opb[23]), .B(gdtr[23]), .Z(n_25278)
		);
	notech_reg gdtr_reg_24(.CP(n_62596), .D(n_25285), .CD(n_61536), .Q(gdtr[
		24]));
	notech_mux2 i_12845(.S(n_54535), .A(opb[24]), .B(gdtr[24]), .Z(n_25285)
		);
	notech_reg gdtr_reg_25(.CP(n_62676), .D(n_25292), .CD(n_61536), .Q(gdtr[
		25]));
	notech_mux2 i_12853(.S(n_54535), .A(opb[25]), .B(gdtr[25]), .Z(n_25292)
		);
	notech_reg gdtr_reg_26(.CP(n_62682), .D(n_25299), .CD(n_61536), .Q(gdtr[
		26]));
	notech_mux2 i_12861(.S(n_54535), .A(opb[26]), .B(gdtr[26]), .Z(n_25299)
		);
	notech_nao3 i_98254606(.A(n_60133), .B(n_60321), .C(n_308891735), .Z(n_1452
		));
	notech_reg gdtr_reg_27(.CP(n_62598), .D(n_25307), .CD(n_61536), .Q(gdtr[
		27]));
	notech_mux2 i_12869(.S(n_54535), .A(opb[27]), .B(gdtr[27]), .Z(n_25307)
		);
	notech_reg gdtr_reg_28(.CP(n_62598), .D(n_25314), .CD(n_61536), .Q(gdtr[
		28]));
	notech_mux2 i_12877(.S(n_54535), .A(opb[28]), .B(gdtr[28]), .Z(n_25314)
		);
	notech_and2 i_31423(.A(n_57068), .B(n_57082), .Z(n_28552));
	notech_reg gdtr_reg_29(.CP(n_62598), .D(n_25321), .CD(n_61537), .Q(gdtr[
		29]));
	notech_mux2 i_12885(.S(n_54535), .A(opb[29]), .B(gdtr[29]), .Z(n_25321)
		);
	notech_reg gdtr_reg_30(.CP(n_62598), .D(n_25328), .CD(n_61537), .Q(gdtr[
		30]));
	notech_mux2 i_12893(.S(n_54535), .A(opb[30]), .B(gdtr[30]), .Z(n_25328)
		);
	notech_reg gdtr_reg_31(.CP(n_62598), .D(n_25337), .CD(n_61537), .Q(gdtr[
		31]));
	notech_mux2 i_12901(.S(n_54535), .A(opb[31]), .B(gdtr[31]), .Z(n_25337)
		);
	notech_reg Daddrgs_reg_0(.CP(n_62598), .D(n_23081), .CD(n_61537), .Q(Daddrgs
		[0]));
	notech_reg Daddrgs_reg_1(.CP(n_62598), .D(n_23088), .CD(n_61536), .Q(Daddrgs
		[1]));
	notech_reg Daddrgs_reg_2(.CP(n_62598), .D(n_23095), .CD(n_61536), .Q(Daddrgs
		[2]));
	notech_reg Daddrgs_reg_3(.CP(n_62598), .D(n_23102), .CD(n_61536), .Q(Daddrgs
		[3]));
	notech_reg Daddrgs_reg_4(.CP(n_62684), .D(n_23109), .CD(n_61533), .Q(Daddrgs
		[4]));
	notech_reg Daddrgs_reg_5(.CP(n_62684), .D(n_23116), .CD(n_61533), .Q(Daddrgs
		[5]));
	notech_reg Daddrgs_reg_6(.CP(n_62684), .D(n_23123), .CD(n_61536), .Q(Daddrgs
		[6]));
	notech_reg Daddrgs_reg_7(.CP(n_62684), .D(n_23130), .CD(n_61536), .Q(Daddrgs
		[7]));
	notech_reg Daddrgs_reg_8(.CP(n_62684), .D(n_23137), .CD(n_61536), .Q(Daddrgs
		[8]));
	notech_reg Daddrgs_reg_9(.CP(n_62684), .D(n_23144), .CD(n_61536), .Q(Daddrgs
		[9]));
	notech_reg Daddrgs_reg_10(.CP(n_62684), .D(n_23151), .CD(n_61536), .Q(Daddrgs
		[10]));
	notech_reg Daddrgs_reg_11(.CP(n_62684), .D(n_23158), .CD(n_61530), .Q(Daddrgs
		[11]));
	notech_reg Daddrgs_reg_12(.CP(n_62684), .D(n_23165), .CD(n_61530), .Q(Daddrgs
		[12]));
	notech_reg Daddrgs_reg_13(.CP(n_62684), .D(n_23172), .CD(n_61530), .Q(Daddrgs
		[13]));
	notech_reg Daddrgs_reg_14(.CP(n_62684), .D(n_23179), .CD(n_61530), .Q(Daddrgs
		[14]));
	notech_reg Daddrgs_reg_15(.CP(n_62684), .D(n_23186), .CD(n_61530), .Q(Daddrgs
		[15]));
	notech_reg Daddrgs_reg_16(.CP(n_62684), .D(n_23193), .CD(n_61530), .Q(Daddrgs
		[16]));
	notech_reg Daddrgs_reg_17(.CP(n_62684), .D(n_23200), .CD(n_61530), .Q(Daddrgs
		[17]));
	notech_reg Daddrgs_reg_18(.CP(n_62684), .D(n_23207), .CD(n_61530), .Q(Daddrgs
		[18]));
	notech_reg Daddrgs_reg_19(.CP(n_62684), .D(n_23214), .CD(n_61530), .Q(Daddrgs
		[19]));
	notech_reg Daddrgs_reg_20(.CP(n_62684), .D(n_23221), .CD(n_61530), .Q(Daddrgs
		[20]));
	notech_reg Daddrgs_reg_21(.CP(n_62684), .D(n_23228), .CD(n_61528), .Q(Daddrgs
		[21]));
	notech_reg Daddrgs_reg_22(.CP(n_62684), .D(n_23235), .CD(n_61528), .Q(Daddrgs
		[22]));
	notech_reg Daddrgs_reg_23(.CP(n_62742), .D(n_23242), .CD(n_61528), .Q(Daddrgs
		[23]));
	notech_reg Daddrgs_reg_24(.CP(n_62682), .D(n_23249), .CD(n_61528), .Q(Daddrgs
		[24]));
	notech_reg Daddrgs_reg_25(.CP(n_62742), .D(n_23256), .CD(n_61528), .Q(Daddrgs
		[25]));
	notech_reg Daddrgs_reg_26(.CP(n_62742), .D(n_23263), .CD(n_61530), .Q(Daddrgs
		[26]));
	notech_reg Daddrgs_reg_27(.CP(n_62742), .D(n_23270), .CD(n_61530), .Q(Daddrgs
		[27]));
	notech_reg Daddrgs_reg_28(.CP(n_62742), .D(n_23277), .CD(n_61528), .Q(Daddrgs
		[28]));
	notech_reg Daddrgs_reg_29(.CP(n_62742), .D(n_23284), .CD(n_61528), .Q(Daddrgs
		[29]));
	notech_reg Daddrgs_reg_30(.CP(n_62742), .D(n_23291), .CD(n_61531), .Q(Daddrgs
		[30]));
	notech_reg Daddrgs_reg_31(.CP(n_62742), .D(n_23298), .CD(n_61531), .Q(Daddrgs
		[31]));
	notech_reg idtr_reg_0(.CP(n_62742), .D(n_25434), .CD(n_61531), .Q(idtr[0
		]));
	notech_mux2 i_13037(.S(n_327790775), .A(opb[0]), .B(idtr[0]), .Z(n_25434
		));
	notech_ao3 i_50355029(.A(n_32386), .B(n_56513), .C(n_56827), .Z(n_1448)
		);
	notech_reg idtr_reg_1(.CP(n_62742), .D(n_25440), .CD(n_61531), .Q(idtr[1
		]));
	notech_mux2 i_13045(.S(n_327790775), .A(opb[1]), .B(idtr[1]), .Z(n_25440
		));
	notech_reg idtr_reg_2(.CP(n_62742), .D(n_25446), .CD(n_61532), .Q(idtr[2
		]));
	notech_mux2 i_13053(.S(n_327790775), .A(opb[2]), .B(idtr[2]), .Z(n_25446
		));
	notech_reg idtr_reg_3(.CP(n_62742), .D(n_25452), .CD(n_61532), .Q(idtr[3
		]));
	notech_mux2 i_13061(.S(n_327790775), .A(opb[3]), .B(idtr[3]), .Z(n_25452
		));
	notech_reg idtr_reg_4(.CP(n_62742), .D(n_25458), .CD(n_61532), .Q(idtr[4
		]));
	notech_mux2 i_13069(.S(n_327790775), .A(opb[4]), .B(idtr[4]), .Z(n_25458
		));
	notech_reg idtr_reg_5(.CP(n_62742), .D(n_25464), .CD(n_61532), .Q(idtr[5
		]));
	notech_mux2 i_13077(.S(n_327790775), .A(opb[5]), .B(idtr[5]), .Z(n_25464
		));
	notech_reg idtr_reg_6(.CP(n_62742), .D(n_25470), .CD(n_61532), .Q(idtr[6
		]));
	notech_mux2 i_13085(.S(n_327790775), .A(opb[6]), .B(idtr[6]), .Z(n_25470
		));
	notech_ao3 i_48055047(.A(n_60133), .B(n_56557), .C(n_56813), .Z(n_1442)
		);
	notech_reg idtr_reg_7(.CP(n_62742), .D(n_25476), .CD(n_61531), .Q(idtr[7
		]));
	notech_mux2 i_13093(.S(n_327790775), .A(opb[7]), .B(idtr[7]), .Z(n_25476
		));
	notech_or4 i_47855048(.A(n_58062), .B(n_2937), .C(n_56827), .D(n_32294),
		 .Z(n_1441));
	notech_reg idtr_reg_8(.CP(n_62742), .D(n_25482), .CD(n_61531), .Q(idtr[8
		]));
	notech_mux2 i_13101(.S(n_327790775), .A(opb[8]), .B(idtr[8]), .Z(n_25482
		));
	notech_ao3 i_47355052(.A(n_56557), .B(n_60133), .C(n_56688), .Z(n_1440)
		);
	notech_reg idtr_reg_9(.CP(n_62742), .D(n_25489), .CD(n_61531), .Q(idtr[9
		]));
	notech_mux2 i_13109(.S(n_327790775), .A(opb[9]), .B(idtr[9]), .Z(n_25489
		));
	notech_reg idtr_reg_10(.CP(n_62742), .D(n_25496), .CD(n_61530), .Q(idtr[
		10]));
	notech_mux2 i_13117(.S(n_327790775), .A(opb[10]), .B(idtr[10]), .Z(n_25496
		));
	notech_ao4 i_7155446(.A(n_60888), .B(n_2893), .C(n_32458), .D(n_27377), 
		.Z(n_1438));
	notech_reg idtr_reg_11(.CP(n_62682), .D(n_25503), .CD(n_61531), .Q(idtr[
		11]));
	notech_mux2 i_13125(.S(n_327790775), .A(opb[11]), .B(idtr[11]), .Z(n_25503
		));
	notech_reg idtr_reg_12(.CP(n_62682), .D(n_25510), .CD(n_61531), .Q(idtr[
		12]));
	notech_mux2 i_13133(.S(n_327790775), .A(opb[12]), .B(idtr[12]), .Z(n_25510
		));
	notech_reg idtr_reg_13(.CP(n_62682), .D(n_25517), .CD(n_61531), .Q(idtr[
		13]));
	notech_mux2 i_13141(.S(n_327790775), .A(opb[13]), .B(idtr[13]), .Z(n_25517
		));
	notech_reg idtr_reg_14(.CP(n_62682), .D(n_25525), .CD(n_61531), .Q(idtr[
		14]));
	notech_mux2 i_13149(.S(n_327790775), .A(opb[14]), .B(idtr[14]), .Z(n_25525
		));
	notech_and3 i_46355062(.A(n_24582), .B(n_24583), .C(n_24589), .Z(n_1434)
		);
	notech_reg idtr_reg_15(.CP(n_62682), .D(n_25532), .CD(n_61531), .Q(idtr[
		15]));
	notech_mux2 i_13157(.S(n_327790775), .A(opb[15]), .B(idtr[15]), .Z(n_25532
		));
	notech_ao4 i_84255518(.A(n_62776), .B(n_60904), .C(n_60888), .D(n_27757)
		, .Z(n_1433));
	notech_reg idtr_reg_16(.CP(n_62682), .D(n_25539), .CD(n_61531), .Q(idtr[
		16]));
	notech_mux2 i_13165(.S(n_54546), .A(opb[16]), .B(idtr[16]), .Z(n_25539)
		);
	notech_reg idtr_reg_17(.CP(n_62682), .D(n_25546), .CD(n_61508), .Q(idtr[
		17]));
	notech_mux2 i_13173(.S(n_54546), .A(opb[17]), .B(idtr[17]), .Z(n_25546)
		);
	notech_nand2 i_2955521(.A(n_62776), .B(opc_10[30]), .Z(n_30809));
	notech_reg idtr_reg_18(.CP(n_62682), .D(n_25553), .CD(n_61508), .Q(idtr[
		18]));
	notech_mux2 i_13181(.S(n_54546), .A(opb[18]), .B(idtr[18]), .Z(n_25553)
		);
	notech_reg idtr_reg_19(.CP(n_62682), .D(n_25561), .CD(n_61508), .Q(idtr[
		19]));
	notech_mux2 i_13189(.S(n_54546), .A(opb[19]), .B(idtr[19]), .Z(n_25561)
		);
	notech_ao3 i_7458417(.A(n_60133), .B(n_60318), .C(n_28532), .Z(n_1430)
		);
	notech_reg idtr_reg_20(.CP(n_62598), .D(n_25568), .CD(n_61508), .Q(idtr[
		20]));
	notech_mux2 i_13197(.S(n_54546), .A(opb[20]), .B(idtr[20]), .Z(n_25568)
		);
	notech_ao3 i_8958402(.A(n_60133), .B(n_60316), .C(n_304091783), .Z(n_1429
		));
	notech_reg idtr_reg_21(.CP(n_62598), .D(n_25575), .CD(n_61508), .Q(idtr[
		21]));
	notech_mux2 i_13205(.S(n_54546), .A(opb[21]), .B(idtr[21]), .Z(n_25575)
		);
	notech_ao4 i_31432(.A(n_56843), .B(n_61133), .C(n_32351), .D(n_32616), .Z
		(n_28543));
	notech_reg idtr_reg_22(.CP(n_62686), .D(n_25582), .CD(n_61508), .Q(idtr[
		22]));
	notech_mux2 i_13213(.S(n_54546), .A(opb[22]), .B(idtr[22]), .Z(n_25582)
		);
	notech_reg idtr_reg_23(.CP(n_62600), .D(n_25589), .CD(n_61509), .Q(idtr[
		23]));
	notech_mux2 i_13221(.S(n_54546), .A(opb[23]), .B(idtr[23]), .Z(n_25589)
		);
	notech_or4 i_31739(.A(n_28544), .B(n_57055), .C(n_57011), .D(n_54916), .Z
		(n_28236));
	notech_reg idtr_reg_24(.CP(n_62600), .D(n_25597), .CD(n_61508), .Q(idtr[
		24]));
	notech_mux2 i_13229(.S(n_54546), .A(opb[24]), .B(idtr[24]), .Z(n_25597)
		);
	notech_or4 i_31741(.A(n_303891785), .B(n_57055), .C(n_57011), .D(n_54916
		), .Z(n_28234));
	notech_reg idtr_reg_25(.CP(n_62600), .D(n_25604), .CD(n_61508), .Q(idtr[
		25]));
	notech_mux2 i_13237(.S(n_54546), .A(opb[25]), .B(idtr[25]), .Z(n_25604)
		);
	notech_or4 i_7058421(.A(n_60274), .B(n_59478), .C(n_2839), .D(n_303991784
		), .Z(n_28532));
	notech_reg idtr_reg_26(.CP(n_62600), .D(n_25611), .CD(n_61508), .Q(idtr[
		26]));
	notech_mux2 i_13245(.S(n_54546), .A(opb[26]), .B(idtr[26]), .Z(n_25611)
		);
	notech_reg idtr_reg_27(.CP(n_62600), .D(n_25627), .CD(n_61507), .Q(idtr[
		27]));
	notech_mux2 i_13253(.S(n_54546), .A(opb[27]), .B(idtr[27]), .Z(n_25627)
		);
	notech_or4 i_34068(.A(n_32614), .B(n_32342), .C(n_54954), .D(n_26054), .Z
		(n_25875));
	notech_reg idtr_reg_28(.CP(n_62600), .D(n_25635), .CD(n_61507), .Q(idtr[
		28]));
	notech_mux2 i_13261(.S(n_54546), .A(opb[28]), .B(idtr[28]), .Z(n_25635)
		);
	notech_nand2 i_34069(.A(n_26767), .B(n_26669), .Z(n_25874));
	notech_reg idtr_reg_29(.CP(n_62600), .D(n_25645), .CD(n_61507), .Q(idtr[
		29]));
	notech_mux2 i_13269(.S(n_54546), .A(opb[29]), .B(idtr[29]), .Z(n_25645)
		);
	notech_reg idtr_reg_30(.CP(n_62600), .D(n_25654), .CD(n_61507), .Q(idtr[
		30]));
	notech_mux2 i_13277(.S(n_54546), .A(opb[30]), .B(idtr[30]), .Z(n_25654)
		);
	notech_ao3 i_105257475(.A(n_60133), .B(n_56570), .C(n_56813), .Z(n_1427)
		);
	notech_reg idtr_reg_31(.CP(n_62600), .D(n_25661), .CD(n_61507), .Q(idtr[
		31]));
	notech_mux2 i_13285(.S(n_54546), .A(opb[31]), .B(idtr[31]), .Z(n_25661)
		);
	notech_reg tr_reg_3(.CP(n_62686), .D(n_25671), .CD(n_61508), .Q(\tr[3] )
		);
	notech_mux2 i_13293(.S(n_317787451), .A(opb[3]), .B(\tr[3] ), .Z(n_25671
		));
	notech_reg tr_reg_4(.CP(n_62686), .D(n_25678), .CD(n_61508), .Q(\tr[4] )
		);
	notech_mux2 i_13301(.S(n_317787451), .A(opb[4]), .B(\tr[4] ), .Z(n_25678
		));
	notech_reg tr_reg_5(.CP(n_62686), .D(n_25684), .CD(n_61507), .Q(\tr[5] )
		);
	notech_mux2 i_13310(.S(n_317787451), .A(opb[5]), .B(\tr[5] ), .Z(n_25684
		));
	notech_reg tr_reg_6(.CP(n_62686), .D(n_25690), .CD(n_61508), .Q(\tr[6] )
		);
	notech_mux2 i_13318(.S(n_317787451), .A(opb[6]), .B(\tr[6] ), .Z(n_25690
		));
	notech_reg tr_reg_7(.CP(n_62686), .D(n_25696), .CD(n_61510), .Q(\tr[7] )
		);
	notech_mux2 i_13326(.S(n_317787451), .A(opb[7]), .B(\tr[7] ), .Z(n_25696
		));
	notech_reg tr_reg_8(.CP(n_62686), .D(n_25702), .CD(n_61510), .Q(\tr[8] )
		);
	notech_mux2 i_13334(.S(n_317787451), .A(opb[8]), .B(\tr[8] ), .Z(n_25702
		));
	notech_reg tr_reg_9(.CP(n_62686), .D(n_25710), .CD(n_61509), .Q(\tr[9] )
		);
	notech_mux2 i_13342(.S(n_317787451), .A(opb[9]), .B(\tr[9] ), .Z(n_25710
		));
	notech_reg tr_reg_10(.CP(n_62686), .D(n_25717), .CD(n_61510), .Q(\tr[10] 
		));
	notech_mux2 i_13350(.S(n_317787451), .A(opb[10]), .B(\tr[10] ), .Z(n_25717
		));
	notech_reg tr_reg_11(.CP(n_62686), .D(n_25725), .CD(n_61510), .Q(\tr[11] 
		));
	notech_mux2 i_13358(.S(n_317787451), .A(opb[11]), .B(\tr[11] ), .Z(n_25725
		));
	notech_reg tr_reg_12(.CP(n_62686), .D(n_25732), .CD(n_61510), .Q(\tr[12] 
		));
	notech_mux2 i_13366(.S(n_317787451), .A(opb[12]), .B(\tr[12] ), .Z(n_25732
		));
	notech_ao4 i_83858517(.A(n_62776), .B(n_60904), .C(n_60888), .D(n_27353)
		, .Z(n_1416));
	notech_reg tr_reg_13(.CP(n_62686), .D(n_25740), .CD(n_61510), .Q(\tr[13] 
		));
	notech_mux2 i_13374(.S(n_317787451), .A(opb[13]), .B(\tr[13] ), .Z(n_25740
		));
	notech_reg tr_reg_14(.CP(n_62686), .D(n_25747), .CD(n_61510), .Q(\tr[14] 
		));
	notech_mux2 i_13382(.S(n_317787451), .A(opb[14]), .B(\tr[14] ), .Z(n_25747
		));
	notech_and3 i_147460329(.A(n_93835734), .B(n_54667), .C(n_131792187), .Z
		(n_1414));
	notech_reg tr_reg_15(.CP(n_62686), .D(n_25755), .CD(n_61510), .Q(\tr[15] 
		));
	notech_mux2 i_13390(.S(n_317787451), .A(opb[15]), .B(\tr[15] ), .Z(n_25755
		));
	notech_reg desc_reg_0(.CP(n_62686), .D(n_25762), .CD(n_61509), .Q(desc[0
		]));
	notech_mux2 i_13398(.S(n_58662), .A(read_data[0]), .B(desc[0]), .Z(n_25762
		));
	notech_reg desc_reg_1(.CP(n_62686), .D(n_25772), .CD(n_61509), .Q(desc[1
		]));
	notech_mux2 i_13406(.S(n_58662), .A(read_data[1]), .B(desc[1]), .Z(n_25772
		));
	notech_ao4 i_147560328(.A(n_302391800), .B(n_27998), .C(n_54934), .D(n_31540
		), .Z(n_1411));
	notech_reg desc_reg_2(.CP(n_62686), .D(n_25783), .CD(n_61509), .Q(desc[2
		]));
	notech_mux2 i_13414(.S(n_58662), .A(read_data[2]), .B(desc[2]), .Z(n_25783
		));
	notech_and4 i_148260321(.A(n_1408), .B(n_132692178), .C(n_1406), .D(n_132392181
		), .Z(n_1410));
	notech_reg desc_reg_3(.CP(n_62686), .D(n_25791), .CD(n_61509), .Q(desc[3
		]));
	notech_mux2 i_13422(.S(n_58662), .A(read_data[3]), .B(desc[3]), .Z(n_25791
		));
	notech_reg desc_reg_4(.CP(n_62686), .D(n_25798), .CD(n_61509), .Q(desc[4
		]));
	notech_mux2 i_13430(.S(n_58662), .A(read_data[4]), .B(desc[4]), .Z(n_25798
		));
	notech_ao4 i_147860325(.A(n_27293), .B(n_57653), .C(n_302091803), .D(n_25875
		), .Z(n_1408));
	notech_reg desc_reg_5(.CP(n_62600), .D(n_25806), .CD(n_61509), .Q(desc[5
		]));
	notech_mux2 i_13438(.S(n_58662), .A(read_data[5]), .B(desc[5]), .Z(n_25806
		));
	notech_reg desc_reg_6(.CP(n_62600), .D(n_25813), .CD(n_61509), .Q(desc[6
		]));
	notech_mux2 i_13446(.S(n_58662), .A(read_data[6]), .B(desc[6]), .Z(n_25813
		));
	notech_ao4 i_148060323(.A(n_301991804), .B(n_30109), .C(n_56605), .D(n_94935745
		), .Z(n_1406));
	notech_reg desc_reg_7(.CP(n_62602), .D(n_25821), .CD(n_61509), .Q(desc[7
		]));
	notech_mux2 i_13454(.S(n_58662), .A(read_data[7]), .B(desc[7]), .Z(n_25821
		));
	notech_reg desc_reg_8(.CP(n_62602), .D(n_25828), .CD(n_61509), .Q(desc[8
		]));
	notech_mux2 i_13462(.S(n_58662), .A(read_data[8]), .B(desc[8]), .Z(n_25828
		));
	notech_and3 i_173060086(.A(n_130992195), .B(n_65435450), .C(n_1403), .Z(n_1404
		));
	notech_reg desc_reg_9(.CP(n_62602), .D(n_25836), .CD(n_61509), .Q(desc[9
		]));
	notech_mux2 i_13470(.S(n_58662), .A(read_data[9]), .B(desc[9]), .Z(n_25836
		));
	notech_ao4 i_172960087(.A(n_27334), .B(n_29590), .C(n_54658), .D(n_29589
		), .Z(n_1403));
	notech_reg desc_reg_10(.CP(n_62602), .D(n_25843), .CD(n_61504), .Q(desc[
		10]));
	notech_mux2 i_13478(.S(n_58662), .A(read_data[10]), .B(desc[10]), .Z(n_25843
		));
	notech_reg desc_reg_11(.CP(n_62602), .D(n_25851), .CD(n_61504), .Q(desc[
		11]));
	notech_mux2 i_13486(.S(n_59158), .A(read_data[11]), .B(desc[11]), .Z(n_25851
		));
	notech_ao4 i_173160085(.A(n_27157), .B(n_30088), .C(n_27142), .D(n_302891795
		), .Z(n_1401));
	notech_reg desc_reg_12(.CP(n_62602), .D(n_25858), .CD(n_61504), .Q(desc[
		12]));
	notech_mux2 i_13494(.S(n_59158), .A(read_data[12]), .B(desc[12]), .Z(n_25858
		));
	notech_ao4 i_173260084(.A(n_27348), .B(n_31476), .C(n_302791796), .D(n_56181
		), .Z(n_1400));
	notech_reg desc_reg_13(.CP(n_62602), .D(n_25865), .CD(n_61504), .Q(desc[
		13]));
	notech_mux2 i_13502(.S(n_59158), .A(read_data[13]), .B(desc[13]), .Z(n_25865
		));
	notech_and4 i_174560076(.A(n_1397), .B(n_1395), .C(n_1394), .D(n_133592169
		), .Z(n_1399));
	notech_reg desc_reg_14(.CP(n_62602), .D(n_25871), .CD(n_61504), .Q(desc[
		14]));
	notech_mux2 i_13510(.S(n_59158), .A(read_data[14]), .B(desc[14]), .Z(n_25871
		));
	notech_reg desc_reg_15(.CP(n_62602), .D(n_25880), .CD(n_61504), .Q(desc[
		15]));
	notech_mux2 i_13518(.S(n_59158), .A(read_data[15]), .B(desc[15]), .Z(n_25880
		));
	notech_ao4 i_173560081(.A(n_27349), .B(n_31456), .C(n_302591798), .D(n_27996
		), .Z(n_1397));
	notech_reg desc_reg_16(.CP(n_62602), .D(n_25888), .CD(n_61504), .Q(desc[
		16]));
	notech_mux2 i_13526(.S(n_59158), .A(read_data[16]), .B(desc[16]), .Z(n_25888
		));
	notech_reg desc_reg_17(.CP(n_62602), .D(n_25894), .CD(n_61504), .Q(desc[
		17]));
	notech_mux2 i_13534(.S(n_59158), .A(read_data[17]), .B(desc[17]), .Z(n_25894
		));
	notech_ao4 i_174060079(.A(n_31492), .B(n_51735313), .C(n_60128), .D(n_27200
		), .Z(n_1395));
	notech_reg desc_reg_18(.CP(n_62602), .D(n_25900), .CD(n_61504), .Q(desc[
		18]));
	notech_mux2 i_13542(.S(n_59158), .A(read_data[18]), .B(desc[18]), .Z(n_25900
		));
	notech_ao4 i_174360078(.A(n_52135317), .B(n_56190), .C(n_302491799), .D(n_52335319
		), .Z(n_1394));
	notech_reg desc_reg_19(.CP(n_62602), .D(n_25906), .CD(n_61504), .Q(desc[
		19]));
	notech_mux2 i_13550(.S(n_59158), .A(read_data[19]), .B(desc[19]), .Z(n_25906
		));
	notech_or2 i_174961734(.A(n_1393), .B(n_27349), .Z(n_52135317));
	notech_reg desc_reg_20(.CP(n_62602), .D(n_25912), .CD(n_61503), .Q(desc[
		20]));
	notech_mux2 i_13558(.S(n_58662), .A(read_data[20]), .B(desc[20]), .Z(n_25912
		));
	notech_or2 i_178360040(.A(n_1416), .B(n_32318), .Z(n_1393));
	notech_reg desc_reg_21(.CP(n_62602), .D(n_25918), .CD(n_61503), .Q(desc[
		21]));
	notech_mux2 i_13566(.S(n_59158), .A(read_data[21]), .B(desc[21]), .Z(n_25918
		));
	notech_nand2 i_184561728(.A(n_26591), .B(n_27344), .Z(n_52335319));
	notech_reg desc_reg_22(.CP(n_62602), .D(n_25924), .CD(n_61503), .Q(desc[
		22]));
	notech_mux2 i_13574(.S(n_59158), .A(read_data[22]), .B(desc[22]), .Z(n_25924
		));
	notech_nor2 i_178460039(.A(n_1416), .B(n_56405), .Z(n_27344));
	notech_reg desc_reg_23(.CP(n_62602), .D(n_25930), .CD(n_61503), .Q(desc[
		23]));
	notech_mux2 i_13582(.S(n_59158), .A(read_data[23]), .B(desc[23]), .Z(n_25930
		));
	notech_and4 i_181360014(.A(n_1390), .B(n_134592159), .C(n_1388), .D(n_134292162
		), .Z(n_1392));
	notech_reg desc_reg_24(.CP(n_62602), .D(n_25936), .CD(n_61503), .Q(desc[
		24]));
	notech_mux2 i_13590(.S(n_327690774), .A(read_data[24]), .B(desc[24]), .Z
		(n_25936));
	notech_reg desc_reg_25(.CP(n_62602), .D(n_25942), .CD(n_61503), .Q(desc[
		25]));
	notech_mux2 i_13598(.S(n_327690774), .A(read_data[25]), .B(desc[25]), .Z
		(n_25942));
	notech_ao4 i_180860018(.A(n_54658), .B(n_29588), .C(n_59326), .D(n_28121
		), .Z(n_1390));
	notech_reg desc_reg_26(.CP(n_62536), .D(n_25949), .CD(n_61504), .Q(desc[
		26]));
	notech_mux2 i_13606(.S(n_327690774), .A(read_data[26]), .B(desc[26]), .Z
		(n_25949));
	notech_reg desc_reg_27(.CP(n_62536), .D(n_25956), .CD(n_61503), .Q(desc[
		27]));
	notech_mux2 i_13615(.S(n_327690774), .A(read_data[27]), .B(desc[27]), .Z
		(n_25956));
	notech_ao4 i_181160016(.A(n_32252), .B(n_26803), .C(n_27319), .D(n_28015
		), .Z(n_1388));
	notech_reg desc_reg_28(.CP(n_62536), .D(n_25964), .CD(n_61503), .Q(desc[
		28]));
	notech_mux2 i_13624(.S(n_327690774), .A(read_data[28]), .B(desc[28]), .Z
		(n_25964));
	notech_and4 i_181860009(.A(n_1385), .B(n_1383), .C(n_134892156), .D(n_135192153
		), .Z(n_1387));
	notech_reg desc_reg_29(.CP(n_62536), .D(n_25971), .CD(n_61505), .Q(desc[
		29]));
	notech_mux2 i_13633(.S(n_327690774), .A(read_data[29]), .B(desc[29]), .Z
		(n_25971));
	notech_reg desc_reg_30(.CP(n_62536), .D(n_25979), .CD(n_61507), .Q(desc[
		30]));
	notech_mux2 i_13641(.S(n_327690774), .A(read_data[30]), .B(desc[30]), .Z
		(n_25979));
	notech_ao4 i_181460013(.A(n_145028727), .B(n_29591), .C(n_144928726), .D
		(n_55929), .Z(n_1385));
	notech_reg desc_reg_31(.CP(n_62536), .D(n_25986), .CD(n_61505), .Q(desc[
		31]));
	notech_mux2 i_13649(.S(n_327690774), .A(read_data[31]), .B(desc[31]), .Z
		(n_25986));
	notech_reg Daddrs_reg_0(.CP(n_62536), .D(n_25994), .CD(n_61505), .Q(Daddr
		[0]));
	notech_mux2 i_13657(.S(\nbus_11377[0] ), .A(Daddr[0]), .B(n_27835), .Z(n_25994
		));
	notech_ao4 i_181660011(.A(n_144828725), .B(n_57828), .C(n_60128), .D(n_27216
		), .Z(n_1383));
	notech_reg Daddrs_reg_1(.CP(n_62536), .D(n_26001), .CD(n_61507), .Q(Daddr
		[1]));
	notech_mux2 i_13665(.S(\nbus_11377[0] ), .A(Daddr[1]), .B(n_27836), .Z(n_26001
		));
	notech_reg Daddrs_reg_2(.CP(n_62536), .D(n_26009), .CD(n_61507), .Q(Daddr
		[2]));
	notech_mux2 i_13673(.S(\nbus_11377[0] ), .A(Daddr[2]), .B(n_27837), .Z(n_26009
		));
	notech_and3 i_189259939(.A(n_62935425), .B(n_1380), .C(n_130692198), .Z(n_1381
		));
	notech_reg Daddrs_reg_3(.CP(n_62448), .D(n_26016), .CD(n_61507), .Q(Daddr
		[3]));
	notech_mux2 i_13681(.S(\nbus_11377[0] ), .A(Daddr[3]), .B(n_27838), .Z(n_26016
		));
	notech_ao4 i_188959940(.A(n_31309), .B(n_28236), .C(n_31307), .D(n_28234
		), .Z(n_1380));
	notech_reg Daddrs_reg_4(.CP(n_62536), .D(n_26025), .CD(n_61507), .Q(Daddr
		[4]));
	notech_mux2 i_13689(.S(\nbus_11377[0] ), .A(Daddr[4]), .B(n_27839), .Z(n_26025
		));
	notech_reg Daddrs_reg_5(.CP(n_62634), .D(n_26032), .CD(n_61507), .Q(Daddr
		[5]));
	notech_mux2 i_13697(.S(\nbus_11377[0] ), .A(Daddr[5]), .B(n_27840), .Z(n_26032
		));
	notech_ao4 i_127361754(.A(n_28222), .B(n_56109), .C(n_57957), .D(n_298991830
		), .Z(n_62935425));
	notech_reg Daddrs_reg_6(.CP(n_62490), .D(n_26041), .CD(n_61505), .Q(Daddr
		[6]));
	notech_mux2 i_13705(.S(\nbus_11377[0] ), .A(Daddr[6]), .B(n_27841), .Z(n_26041
		));
	notech_reg Daddrs_reg_7(.CP(n_62490), .D(n_26049), .CD(n_61505), .Q(Daddr
		[7]));
	notech_mux2 i_13713(.S(\nbus_11377[0] ), .A(Daddr[7]), .B(n_27842), .Z(n_26049
		));
	notech_ao4 i_189359938(.A(n_303291791), .B(n_56100), .C(n_28544), .D(n_31279
		), .Z(n_1378));
	notech_reg Daddrs_reg_8(.CP(n_62490), .D(n_26064), .CD(n_61505), .Q(Daddr
		[8]));
	notech_mux2 i_13721(.S(\nbus_11377[0] ), .A(Daddr[8]), .B(n_27843), .Z(n_26064
		));
	notech_and4 i_190359930(.A(n_1375), .B(n_1373), .C(n_1372), .D(n_1359), 
		.Z(n_1377));
	notech_reg Daddrs_reg_9(.CP(n_62562), .D(n_26071), .CD(n_61504), .Q(Daddr
		[9]));
	notech_mux2 i_13729(.S(\nbus_11377[0] ), .A(Daddr[9]), .B(n_27844), .Z(n_26071
		));
	notech_reg Daddrs_reg_10(.CP(n_62562), .D(n_26079), .CD(n_61505), .Q(Daddr
		[10]));
	notech_mux2 i_13737(.S(\nbus_11377[0] ), .A(Daddr[10]), .B(n_25548), .Z(n_26079
		));
	notech_ao4 i_189659935(.A(n_54649), .B(n_29587), .C(n_60133), .D(n_27224
		), .Z(n_1375));
	notech_reg Daddrs_reg_11(.CP(n_62562), .D(n_26086), .CD(n_61505), .Q(Daddr
		[11]));
	notech_mux2 i_13745(.S(\nbus_11377[0] ), .A(Daddr[11]), .B(n_25554), .Z(n_26086
		));
	notech_reg Daddrs_reg_12(.CP(n_62562), .D(n_26094), .CD(n_61505), .Q(Daddr
		[12]));
	notech_mux2 i_13753(.S(\nbus_11377[0] ), .A(Daddr[12]), .B(n_25560), .Z(n_26094
		));
	notech_ao4 i_189859933(.A(n_303191792), .B(n_300091823), .C(n_300291821)
		, .D(n_29614), .Z(n_1373));
	notech_reg Daddrs_reg_13(.CP(n_62562), .D(n_26101), .CD(n_61505), .Q(Daddr
		[13]));
	notech_mux2 i_13761(.S(\nbus_11377[0] ), .A(Daddr[13]), .B(n_25566), .Z(n_26101
		));
	notech_ao4 i_189959932(.A(n_130492200), .B(n_56109), .C(n_57957), .D(n_30233
		), .Z(n_1372));
	notech_reg Daddrs_reg_14(.CP(n_62562), .D(n_26108), .CD(n_61505), .Q(Daddr
		[14]));
	notech_mux2 i_13769(.S(\nbus_11377[0] ), .A(Daddr[14]), .B(n_25572), .Z(n_26108
		));
	notech_reg Daddrs_reg_15(.CP(n_62562), .D(n_26114), .CD(n_61505), .Q(Daddr
		[15]));
	notech_mux2 i_13777(.S(\nbus_11377[0] ), .A(Daddr[15]), .B(n_25578), .Z(n_26114
		));
	notech_ao4 i_114361759(.A(n_302491799), .B(n_102135817), .C(n_102035816)
		, .D(n_56190), .Z(n_65435450));
	notech_reg Daddrs_reg_16(.CP(n_62562), .D(n_26120), .CD(n_61517), .Q(Daddr
		[16]));
	notech_mux2 i_13785(.S(n_55438), .A(Daddr[16]), .B(n_25584), .Z(n_26120)
		);
	notech_and3 i_66361770(.A(n_1369), .B(n_1371), .C(n_1368), .Z(n_93835734
		));
	notech_reg Daddrs_reg_17(.CP(n_62562), .D(n_26126), .CD(n_61517), .Q(Daddr
		[17]));
	notech_mux2 i_13793(.S(n_55438), .A(Daddr[17]), .B(n_25590), .Z(n_26126)
		);
	notech_ao4 i_220259636(.A(n_56230), .B(n_30569), .C(n_30568), .D(n_57653
		), .Z(n_1371));
	notech_reg Daddrs_reg_18(.CP(n_62562), .D(n_26132), .CD(n_61517), .Q(Daddr
		[18]));
	notech_mux2 i_13801(.S(n_55438), .A(Daddr[18]), .B(n_25596), .Z(n_26132)
		);
	notech_reg Daddrs_reg_19(.CP(n_62562), .D(n_26138), .CD(n_61517), .Q(Daddr
		[19]));
	notech_mux2 i_13809(.S(n_55438), .A(Daddr[19]), .B(n_25602), .Z(n_26138)
		);
	notech_ao4 i_220359635(.A(n_60316), .B(n_28102), .C(n_30570), .D(n_56239
		), .Z(n_1369));
	notech_reg Daddrs_reg_20(.CP(n_62562), .D(n_26144), .CD(n_61517), .Q(Daddr
		[20]));
	notech_mux2 i_13817(.S(n_55438), .A(Daddr[20]), .B(n_25608), .Z(n_26144)
		);
	notech_or4 i_65761771(.A(n_58101), .B(n_56970), .C(n_56827), .D(n_301691807
		), .Z(n_94935745));
	notech_reg Daddrs_reg_21(.CP(n_62562), .D(n_26150), .CD(n_61519), .Q(Daddr
		[21]));
	notech_mux2 i_13825(.S(n_55438), .A(Daddr[21]), .B(n_25614), .Z(n_26150)
		);
	notech_or4 i_114060643(.A(n_59708), .B(n_56959), .C(n_302091803), .D(n_60207
		), .Z(n_1368));
	notech_reg Daddrs_reg_22(.CP(n_62562), .D(n_26156), .CD(n_61519), .Q(Daddr
		[22]));
	notech_mux2 i_13833(.S(n_55438), .A(Daddr[22]), .B(n_25620), .Z(n_26156)
		);
	notech_reg Daddrs_reg_23(.CP(n_62562), .D(n_26162), .CD(n_61517), .Q(Daddr
		[23]));
	notech_mux2 i_13841(.S(n_55438), .A(Daddr[23]), .B(n_25626), .Z(n_26162)
		);
	notech_reg Daddrs_reg_24(.CP(n_62562), .D(n_26168), .CD(n_61517), .Q(Daddr
		[24]));
	notech_mux2 i_13849(.S(n_55438), .A(Daddr[24]), .B(n_25632), .Z(n_26168)
		);
	notech_reg Daddrs_reg_25(.CP(n_62562), .D(n_26174), .CD(n_61517), .Q(Daddr
		[25]));
	notech_mux2 i_13857(.S(n_55438), .A(Daddr[25]), .B(n_25638), .Z(n_26174)
		);
	notech_reg Daddrs_reg_26(.CP(n_62562), .D(n_26180), .CD(n_61516), .Q(Daddr
		[26]));
	notech_mux2 i_13865(.S(n_55438), .A(Daddr[26]), .B(n_25644), .Z(n_26180)
		);
	notech_reg Daddrs_reg_27(.CP(n_62562), .D(n_26186), .CD(n_61516), .Q(Daddr
		[27]));
	notech_mux2 i_13873(.S(n_55438), .A(Daddr[27]), .B(n_25650), .Z(n_26186)
		);
	notech_reg Daddrs_reg_28(.CP(n_62634), .D(n_26192), .CD(n_61516), .Q(Daddr
		[28]));
	notech_mux2 i_13881(.S(n_55438), .A(Daddr[28]), .B(n_25656), .Z(n_26192)
		);
	notech_reg Daddrs_reg_29(.CP(n_62560), .D(n_26198), .CD(n_61516), .Q(Daddr
		[29]));
	notech_mux2 i_13889(.S(n_55438), .A(Daddr[29]), .B(n_239659477), .Z(n_26198
		));
	notech_reg Daddrs_reg_30(.CP(n_62634), .D(n_26204), .CD(n_61517), .Q(Daddr
		[30]));
	notech_mux2 i_13897(.S(n_55438), .A(Daddr[30]), .B(n_25668), .Z(n_26204)
		);
	notech_nand3 i_75760995(.A(n_1430), .B(n_6363), .C(n_56163), .Z(n_1359)
		);
	notech_reg Daddrs_reg_31(.CP(n_62634), .D(n_26210), .CD(n_61517), .Q(Daddr
		[31]));
	notech_mux2 i_13905(.S(n_55438), .A(Daddr[31]), .B(n_25674), .Z(n_26210)
		);
	notech_reg write_sz_reg_0(.CP(n_62634), .D(n_26216), .CD(n_61517), .Q(write_sz
		[0]));
	notech_mux2 i_13913(.S(n_27846), .A(write_sz[0]), .B(n_307084061), .Z(n_26216
		));
	notech_reg_set write_sz_reg_1(.CP(n_62634), .D(n_26222), .SD(n_61517), .Q
		(write_sz[1]));
	notech_mux2 i_13921(.S(n_27846), .A(write_sz[1]), .B(n_27845), .Z(n_26222
		));
	notech_or4 i_76060992(.A(n_56675), .B(n_56566), .C(n_303391790), .D(n_61136
		), .Z(n_1356));
	notech_reg flush_tlb_reg(.CP(n_62634), .D(n_26229), .CD(n_61517), .Q(flush_tlb
		));
	notech_mux2 i_13929(.S(n_22030), .A(flush_tlb), .B(n_60316), .Z(n_26229)
		);
	notech_reg read_req_reg(.CP(n_62634), .D(n_26235), .CD(n_61520), .Q(read_reqs
		));
	notech_mux2 i_13937(.S(n_21582), .A(read_reqs), .B(n_21585), .Z(n_26235)
		);
	notech_reg writeio_req_reg(.CP(n_62634), .D(n_26241), .CD(n_61520), .Q(writeio_req
		));
	notech_mux2 i_13945(.S(n_19986), .A(writeio_req), .B(n_60316), .Z(n_26241
		));
	notech_reg flush_Dtlb_reg(.CP(n_62634), .D(n_26247), .CD(n_61519), .Q(flush_Dtlb
		));
	notech_mux2 i_13953(.S(n_19963), .A(flush_Dtlb), .B(n_328490782), .Z(n_26247
		));
	notech_reg write_req_reg(.CP(n_62634), .D(n_26254), .CD(n_61520), .Q(write_reqs
		));
	notech_mux2 i_13961(.S(n_14840), .A(write_reqs), .B(n_14843), .Z(n_26254
		));
	notech_or2 i_65361093(.A(n_302991794), .B(n_145128728), .Z(n_135192153)
		);
	notech_reg_set terms_reg(.CP(n_62634), .D(n_26261), .SD(n_61520), .Q(terminate
		));
	notech_mux2 i_13969(.S(n_14789), .A(terminate), .B(n_14792), .Z(n_26261)
		);
	notech_reg writeio_data_reg_0(.CP(n_62634), .D(n_26267), .CD(n_61520), .Q
		(writeio_data[0]));
	notech_mux2 i_13977(.S(n_60123), .A(n_60072), .B(writeio_data[0]), .Z(n_26267
		));
	notech_reg writeio_data_reg_1(.CP(n_62634), .D(n_26273), .CD(n_61520), .Q
		(writeio_data[1]));
	notech_mux2 i_13985(.S(n_60123), .A(opa[1]), .B(writeio_data[1]), .Z(n_26273
		));
	notech_or2 i_65861090(.A(n_303091793), .B(n_144428721), .Z(n_134892156)
		);
	notech_reg writeio_data_reg_2(.CP(n_62634), .D(n_26279), .CD(n_61520), .Q
		(writeio_data[2]));
	notech_mux2 i_13993(.S(n_60123), .A(opa[2]), .B(writeio_data[2]), .Z(n_26279
		));
	notech_reg writeio_data_reg_3(.CP(n_62634), .D(n_26285), .CD(n_61520), .Q
		(writeio_data[3]));
	notech_mux2 i_14001(.S(n_60123), .A(opa[3]), .B(writeio_data[3]), .Z(n_26285
		));
	notech_reg writeio_data_reg_4(.CP(n_62634), .D(n_26291), .CD(n_61519), .Q
		(writeio_data[4]));
	notech_mux2 i_14009(.S(n_60123), .A(opa[4]), .B(writeio_data[4]), .Z(n_26291
		));
	notech_or4 i_66161087(.A(n_184892035), .B(n_30809), .C(n_54916), .D(n_27712
		), .Z(n_134592159));
	notech_reg writeio_data_reg_5(.CP(n_62634), .D(n_26297), .CD(n_61519), .Q
		(writeio_data[5]));
	notech_mux2 i_14017(.S(n_60123), .A(opa[5]), .B(writeio_data[5]), .Z(n_26297
		));
	notech_reg writeio_data_reg_6(.CP(n_62634), .D(n_26303), .CD(n_61519), .Q
		(writeio_data[6]));
	notech_mux2 i_14025(.S(n_60123), .A(n_60082), .B(writeio_data[6]), .Z(n_26303
		));
	notech_reg writeio_data_reg_7(.CP(n_62490), .D(n_26309), .CD(n_61519), .Q
		(writeio_data[7]));
	notech_mux2 i_14033(.S(n_60123), .A(n_60091), .B(writeio_data[7]), .Z(n_26309
		));
	notech_nand3 i_66661084(.A(n_54834), .B(n_7342), .C(n_56172), .Z(n_134292162
		));
	notech_reg writeio_data_reg_8(.CP(n_62560), .D(n_26315), .CD(n_61519), .Q
		(writeio_data[8]));
	notech_mux2 i_14041(.S(n_60123), .A(opa[8]), .B(writeio_data[8]), .Z(n_26315
		));
	notech_reg writeio_data_reg_9(.CP(n_62560), .D(n_26321), .CD(n_61519), .Q
		(writeio_data[9]));
	notech_mux2 i_14049(.S(n_60123), .A(opa[9]), .B(writeio_data[9]), .Z(n_26321
		));
	notech_reg writeio_data_reg_10(.CP(n_62560), .D(n_26327), .CD(n_61519), 
		.Q(writeio_data[10]));
	notech_mux2 i_14057(.S(n_60123), .A(opa[10]), .B(writeio_data[10]), .Z(n_26327
		));
	notech_reg writeio_data_reg_11(.CP(n_62490), .D(n_26333), .CD(n_61519), 
		.Q(writeio_data[11]));
	notech_mux2 i_14065(.S(n_60123), .A(opa[11]), .B(writeio_data[11]), .Z(n_26333
		));
	notech_reg writeio_data_reg_12(.CP(n_62560), .D(n_26339), .CD(n_61519), 
		.Q(writeio_data[12]));
	notech_mux2 i_14073(.S(n_60123), .A(opa[12]), .B(writeio_data[12]), .Z(n_26339
		));
	notech_reg writeio_data_reg_13(.CP(n_62564), .D(n_26345), .CD(n_61519), 
		.Q(writeio_data[13]));
	notech_mux2 i_14081(.S(n_60123), .A(opa[13]), .B(writeio_data[13]), .Z(n_26345
		));
	notech_reg writeio_data_reg_14(.CP(n_62518), .D(n_26351), .CD(n_61514), 
		.Q(writeio_data[14]));
	notech_mux2 i_14089(.S(n_60123), .A(opa[14]), .B(writeio_data[14]), .Z(n_26351
		));
	notech_or2 i_57061164(.A(n_302691797), .B(n_57635), .Z(n_133592169));
	notech_reg writeio_data_reg_15(.CP(n_62518), .D(n_26357), .CD(n_61514), 
		.Q(writeio_data[15]));
	notech_mux2 i_14097(.S(n_60387), .A(n_60102), .B(writeio_data[15]), .Z(n_26357
		));
	notech_reg writeio_data_reg_16(.CP(n_62518), .D(n_26363), .CD(n_61514), 
		.Q(writeio_data[16]));
	notech_mux2 i_14105(.S(n_60387), .A(opa[16]), .B(writeio_data[16]), .Z(n_26363
		));
	notech_reg writeio_data_reg_17(.CP(n_62564), .D(n_26369), .CD(n_61514), 
		.Q(writeio_data[17]));
	notech_mux2 i_14113(.S(n_60387), .A(opa[17]), .B(writeio_data[17]), .Z(n_26369
		));
	notech_reg writeio_data_reg_18(.CP(n_62564), .D(n_26375), .CD(n_61514), 
		.Q(writeio_data[18]));
	notech_mux2 i_14121(.S(n_60387), .A(opa[18]), .B(writeio_data[18]), .Z(n_26375
		));
	notech_reg writeio_data_reg_19(.CP(n_62564), .D(n_26381), .CD(n_61515), 
		.Q(writeio_data[19]));
	notech_mux2 i_14129(.S(n_60387), .A(opa[19]), .B(writeio_data[19]), .Z(n_26381
		));
	notech_reg writeio_data_reg_20(.CP(n_62564), .D(n_26387), .CD(n_61515), 
		.Q(writeio_data[20]));
	notech_mux2 i_14137(.S(n_60387), .A(opa[20]), .B(writeio_data[20]), .Z(n_26387
		));
	notech_reg writeio_data_reg_21(.CP(n_62564), .D(n_26394), .CD(n_61514), 
		.Q(writeio_data[21]));
	notech_mux2 i_14145(.S(n_60387), .A(opa[21]), .B(writeio_data[21]), .Z(n_26394
		));
	notech_reg writeio_data_reg_22(.CP(n_62564), .D(n_26400), .CD(n_61514), 
		.Q(writeio_data[22]));
	notech_mux2 i_14153(.S(n_60387), .A(opa[22]), .B(writeio_data[22]), .Z(n_26400
		));
	notech_reg writeio_data_reg_23(.CP(n_62564), .D(n_26406), .CD(n_61514), 
		.Q(writeio_data[23]));
	notech_mux2 i_14161(.S(n_60387), .A(opa[23]), .B(writeio_data[23]), .Z(n_26406
		));
	notech_or4 i_28861440(.A(n_54954), .B(n_54934), .C(n_32335), .D(n_56239)
		, .Z(n_132692178));
	notech_reg writeio_data_reg_24(.CP(n_62564), .D(n_26412), .CD(n_61510), 
		.Q(writeio_data[24]));
	notech_mux2 i_14170(.S(n_60387), .A(opa[24]), .B(writeio_data[24]), .Z(n_26412
		));
	notech_reg writeio_data_reg_25(.CP(n_62564), .D(n_26418), .CD(n_61510), 
		.Q(writeio_data[25]));
	notech_mux2 i_14178(.S(n_60387), .A(opa[25]), .B(writeio_data[25]), .Z(n_26418
		));
	notech_reg writeio_data_reg_26(.CP(n_62564), .D(n_26424), .CD(n_61510), 
		.Q(writeio_data[26]));
	notech_mux2 i_14186(.S(n_60123), .A(opa[26]), .B(writeio_data[26]), .Z(n_26424
		));
	notech_or2 i_29161437(.A(n_302291801), .B(n_56230), .Z(n_132392181));
	notech_reg writeio_data_reg_27(.CP(n_62564), .D(n_26430), .CD(n_61510), 
		.Q(writeio_data[27]));
	notech_mux2 i_14194(.S(n_60387), .A(opa[27]), .B(writeio_data[27]), .Z(n_26430
		));
	notech_reg writeio_data_reg_28(.CP(n_62564), .D(n_26436), .CD(n_61514), 
		.Q(writeio_data[28]));
	notech_mux2 i_14202(.S(n_60387), .A(opa[28]), .B(writeio_data[28]), .Z(n_26436
		));
	notech_reg writeio_data_reg_29(.CP(n_62564), .D(n_26442), .CD(n_61514), 
		.Q(writeio_data[29]));
	notech_mux2 i_14210(.S(n_60387), .A(opa[29]), .B(writeio_data[29]), .Z(n_26442
		));
	notech_or4 i_29461434(.A(n_55581), .B(n_31560), .C(n_27119), .D(n_54934)
		, .Z(n_132092184));
	notech_reg writeio_data_reg_30(.CP(n_62564), .D(n_26448), .CD(n_61514), 
		.Q(writeio_data[30]));
	notech_mux2 i_14218(.S(n_60387), .A(opa[30]), .B(writeio_data[30]), .Z(n_26448
		));
	notech_reg writeio_data_reg_31(.CP(n_62518), .D(n_26454), .CD(n_61514), 
		.Q(writeio_data[31]));
	notech_mux2 i_14226(.S(n_60387), .A(opa[31]), .B(writeio_data[31]), .Z(n_26454
		));
	notech_reg io_add_reg_0(.CP(n_62564), .D(n_26460), .CD(n_61514), .Q(io_add
		[0]));
	notech_mux2 i_14234(.S(\nbus_11298[0] ), .A(io_add[0]), .B(n_45791242), 
		.Z(n_26460));
	notech_or4 i_29561433(.A(n_62830), .B(n_25874), .C(n_60933), .D(n_56239)
		, .Z(n_131792187));
	notech_reg io_add_reg_1(.CP(n_62564), .D(n_26466), .CD(n_61516), .Q(io_add
		[1]));
	notech_mux2 i_14242(.S(\nbus_11298[0] ), .A(io_add[1]), .B(n_317987453),
		 .Z(n_26466));
	notech_nao3 i_123460559(.A(n_60133), .B(n_60318), .C(n_30470), .Z(n_131692188
		));
	notech_reg io_add_reg_2(.CP(n_62564), .D(n_26472), .CD(n_61516), .Q(io_add
		[2]));
	notech_mux2 i_14250(.S(\nbus_11298[0] ), .A(io_add[2]), .B(n_45991244), 
		.Z(n_26472));
	notech_reg io_add_reg_3(.CP(n_62518), .D(n_26478), .CD(n_61516), .Q(io_add
		[3]));
	notech_mux2 i_14258(.S(\nbus_11298[0] ), .A(io_add[3]), .B(n_318087454),
		 .Z(n_26478));
	notech_reg io_add_reg_4(.CP(n_62564), .D(n_26484), .CD(n_61516), .Q(io_add
		[4]));
	notech_mux2 i_14266(.S(\nbus_11298[0] ), .A(io_add[4]), .B(n_318187455),
		 .Z(n_26484));
	notech_reg io_add_reg_5(.CP(n_62518), .D(n_26490), .CD(n_61516), .Q(io_add
		[5]));
	notech_mux2 i_14274(.S(\nbus_11298[0] ), .A(io_add[5]), .B(n_46091245), 
		.Z(n_26490));
	notech_and3 i_119060601(.A(n_26613), .B(n_26614), .C(n_26616), .Z(n_131292192
		));
	notech_reg io_add_reg_6(.CP(n_62518), .D(n_26496), .CD(n_61516), .Q(io_add
		[6]));
	notech_mux2 i_14282(.S(\nbus_11298[0] ), .A(io_add[6]), .B(n_318287456),
		 .Z(n_26496));
	notech_reg io_add_reg_7(.CP(n_62518), .D(n_26502), .CD(n_61516), .Q(io_add
		[7]));
	notech_mux2 i_14290(.S(\nbus_11298[0] ), .A(io_add[7]), .B(n_318387457),
		 .Z(n_26502));
	notech_reg io_add_reg_8(.CP(n_62518), .D(n_26508), .CD(n_61516), .Q(io_add
		[8]));
	notech_mux2 i_14298(.S(\nbus_11298[0] ), .A(io_add[8]), .B(n_318487458),
		 .Z(n_26508));
	notech_nand3 i_79760957(.A(n_60133), .B(n_60207), .C(read_data[11]), .Z(n_130992195
		));
	notech_reg io_add_reg_9(.CP(n_62518), .D(n_26514), .CD(n_61516), .Q(io_add
		[9]));
	notech_mux2 i_14306(.S(\nbus_11298[0] ), .A(io_add[9]), .B(n_318587459),
		 .Z(n_26514));
	notech_reg io_add_reg_10(.CP(n_62518), .D(n_26520), .CD(n_61515), .Q(io_add
		[10]));
	notech_mux2 i_14314(.S(\nbus_11298[0] ), .A(io_add[10]), .B(n_318687460)
		, .Z(n_26520));
	notech_reg io_add_reg_11(.CP(n_62518), .D(n_26526), .CD(n_61515), .Q(io_add
		[11]));
	notech_mux2 i_14322(.S(\nbus_11298[0] ), .A(io_add[11]), .B(n_318787461)
		, .Z(n_26526));
	notech_nand3 i_76560988(.A(n_60133), .B(n_60207), .C(read_data[7]), .Z(n_130692198
		));
	notech_reg io_add_reg_12(.CP(n_62518), .D(n_26532), .CD(n_61515), .Q(io_add
		[12]));
	notech_mux2 i_14330(.S(\nbus_11298[0] ), .A(io_add[12]), .B(n_318887462)
		, .Z(n_26532));
	notech_reg io_add_reg_13(.CP(n_62518), .D(n_26538), .CD(n_61515), .Q(io_add
		[13]));
	notech_mux2 i_14338(.S(\nbus_11298[0] ), .A(io_add[13]), .B(n_318987463)
		, .Z(n_26538));
	notech_and2 i_1661708(.A(n_301891805), .B(n_299991824), .Z(n_130492200)
		);
	notech_reg io_add_reg_14(.CP(n_62518), .D(n_26544), .CD(n_61515), .Q(io_add
		[14]));
	notech_mux2 i_14346(.S(\nbus_11298[0] ), .A(io_add[14]), .B(n_319087464)
		, .Z(n_26544));
	notech_ao4 i_1561709(.A(n_59441), .B(n_27302), .C(n_28332), .D(n_26683),
		 .Z(n_130392201));
	notech_reg io_add_reg_15(.CP(n_62518), .D(n_26550), .CD(n_61515), .Q(io_add
		[15]));
	notech_mux2 i_14354(.S(\nbus_11298[0] ), .A(io_add[15]), .B(n_319187465)
		, .Z(n_26550));
	notech_nand2 i_108961763(.A(n_28544), .B(n_28543), .Z(n_28542));
	notech_reg pc_req_reg(.CP(n_62518), .D(n_26556), .CD(n_61515), .Q(pc_req
		));
	notech_mux2 i_14362(.S(n_12360), .A(pc_req), .B(n_60318), .Z(n_26556));
	notech_nand2 i_3761780(.A(n_62776), .B(opc[13]), .Z(n_30109));
	notech_reg had_lgjmp_reg(.CP(n_62518), .D(n_26562), .CD(n_61515), .Q(had_lgjmp
		));
	notech_mux2 i_14370(.S(n_317687450), .A(\nbus_14522[31] ), .B(had_lgjmp)
		, .Z(n_26562));
	notech_reg readio_req_reg(.CP(n_62518), .D(n_26568), .CD(n_61515), .Q(readio_req
		));
	notech_mux2 i_14378(.S(n_12080), .A(readio_req), .B(n_60316), .Z(n_26568
		));
	notech_inv i_30623(.A(n_212669138), .Z(n_26574));
	notech_inv i_30624(.A(n_257069582), .Z(n_26575));
	notech_inv i_30626(.A(n_207269084), .Z(n_26576));
	notech_inv i_30627(.A(n_207169083), .Z(n_26577));
	notech_inv i_30628(.A(n_258969601), .Z(n_26578));
	notech_inv i_30629(.A(n_259669608), .Z(n_26579));
	notech_inv i_30630(.A(n_261169623), .Z(n_26581));
	notech_inv i_30631(.A(n_204069052), .Z(n_26582));
	notech_inv i_30632(.A(n_266969681), .Z(n_26583));
	notech_inv i_30633(.A(n_267669688), .Z(n_26584));
	notech_inv i_30634(.A(n_203169043), .Z(n_26585));
	notech_inv i_30636(.A(n_203069042), .Z(n_26586));
	notech_inv i_30637(.A(n_272069732), .Z(n_26587));
	notech_inv i_30638(.A(n_272969741), .Z(n_26588));
	notech_inv i_30639(.A(n_273869750), .Z(n_26589));
	notech_inv i_30640(.A(n_289369905), .Z(n_26590));
	notech_inv i_30641(.A(n_27349), .Z(n_26591));
	notech_inv i_30642(.A(n_197268985), .Z(n_26592));
	notech_inv i_30643(.A(n_307091753), .Z(n_26593));
	notech_inv i_30644(.A(n_112564654), .Z(n_26594));
	notech_inv i_30645(.A(n_4010), .Z(n_26595));
	notech_inv i_30646(.A(n_24994), .Z(n_26596));
	notech_inv i_30647(.A(n_313470145), .Z(n_26597));
	notech_inv i_30648(.A(n_313870149), .Z(n_26598));
	notech_inv i_30649(.A(n_58504), .Z(n_26599));
	notech_inv i_30650(.A(n_322670237), .Z(n_26600));
	notech_inv i_30651(.A(n_27757), .Z(n_26601));
	notech_inv i_30652(.A(n_1901), .Z(n_26602));
	notech_inv i_30653(.A(n_346170472), .Z(n_26603));
	notech_inv i_30654(.A(n_117868195), .Z(n_26604));
	notech_inv i_30655(.A(n_157368590), .Z(n_26605));
	notech_inv i_30656(.A(n_311591708), .Z(n_26606));
	notech_inv i_30657(.A(n_313170142), .Z(n_26607));
	notech_inv i_30658(.A(n_3996), .Z(n_26608));
	notech_inv i_30659(.A(n_186768883), .Z(n_26609));
	notech_inv i_30660(.A(n_32386), .Z(n_26610));
	notech_inv i_30661(.A(n_213069142), .Z(n_26612));
	notech_inv i_30662(.A(n_287027252), .Z(n_26615));
	notech_inv i_30663(.A(n_258469596), .Z(n_26617));
	notech_inv i_30664(.A(n_258069592), .Z(n_26618));
	notech_inv i_30665(.A(n_257669588), .Z(n_26619));
	notech_inv i_30666(.A(n_288369895), .Z(n_26621));
	notech_inv i_30667(.A(n_287969891), .Z(n_26622));
	notech_inv i_30668(.A(n_287569887), .Z(n_26623));
	notech_inv i_30669(.A(n_288769899), .Z(n_26624));
	notech_inv i_30670(.A(n_306191762), .Z(n_26625));
	notech_inv i_30671(.A(n_306391760), .Z(n_26626));
	notech_inv i_30672(.A(n_314291681), .Z(n_26627));
	notech_inv i_30673(.A(n_124871728), .Z(n_26628));
	notech_inv i_30674(.A(n_122071700), .Z(n_26629));
	notech_inv i_30675(.A(n_127871758), .Z(n_26630));
	notech_inv i_30676(.A(n_153372013), .Z(n_26631));
	notech_inv i_30677(.A(n_183772317), .Z(n_26632));
	notech_inv i_30678(.A(n_184272322), .Z(n_26633));
	notech_inv i_30679(.A(n_1904), .Z(n_26634));
	notech_inv i_30680(.A(n_184472324), .Z(n_26635));
	notech_inv i_30681(.A(n_184772327), .Z(n_26636));
	notech_inv i_30682(.A(n_185372333), .Z(n_26637));
	notech_inv i_30683(.A(n_27906), .Z(n_26638));
	notech_inv i_30684(.A(n_4013), .Z(n_26640));
	notech_inv i_30685(.A(n_58496), .Z(n_26641));
	notech_inv i_30686(.A(n_148128758), .Z(n_26642));
	notech_inv i_30687(.A(n_1902), .Z(n_26643));
	notech_inv i_30688(.A(n_344466973), .Z(n_26644));
	notech_inv i_30689(.A(n_312147737), .Z(n_26645));
	notech_inv i_30690(.A(n_58622), .Z(n_26646));
	notech_inv i_30691(.A(n_58714), .Z(n_26647));
	notech_inv i_30692(.A(n_310991714), .Z(n_26648));
	notech_inv i_30694(.A(n_32294), .Z(n_26649));
	notech_inv i_30699(.A(n_32373), .Z(n_26651));
	notech_inv i_30700(.A(n_250972989), .Z(n_26652));
	notech_inv i_30701(.A(n_251672996), .Z(n_26653));
	notech_inv i_30702(.A(n_252373003), .Z(n_26654));
	notech_inv i_30703(.A(n_255573035), .Z(n_26655));
	notech_inv i_30704(.A(n_256473044), .Z(n_26656));
	notech_inv i_30705(.A(n_263073110), .Z(n_26657));
	notech_inv i_30706(.A(n_266173141), .Z(n_26658));
	notech_inv i_30707(.A(n_275173231), .Z(n_26659));
	notech_inv i_30708(.A(n_312073600), .Z(n_26660));
	notech_inv i_30709(.A(n_317673656), .Z(n_26661));
	notech_inv i_30710(.A(n_58482), .Z(n_26662));
	notech_inv i_30712(.A(n_32344), .Z(n_26664));
	notech_inv i_30720(.A(n_292666455), .Z(n_26667));
	notech_inv i_30721(.A(n_28544), .Z(n_26668));
	notech_inv i_30722(.A(n_54934), .Z(n_26669));
	notech_inv i_30723(.A(n_3845), .Z(n_26670));
	notech_inv i_30725(.A(n_58316), .Z(n_26671));
	notech_inv i_30726(.A(n_152672006), .Z(n_26672));
	notech_inv i_30727(.A(n_278566314), .Z(n_26673));
	notech_inv i_30728(.A(n_284566374), .Z(n_26674));
	notech_inv i_30729(.A(n_307324337), .Z(n_26675));
	notech_inv i_30730(.A(n_306073540), .Z(n_26676));
	notech_inv i_30731(.A(n_306273542), .Z(n_26677));
	notech_inv i_30732(.A(n_309791726), .Z(n_26678));
	notech_inv i_30733(.A(n_58055), .Z(n_26679));
	notech_inv i_30734(.A(n_58378), .Z(n_26680));
	notech_inv i_30736(.A(n_28546), .Z(n_26681));
	notech_inv i_30737(.A(n_119175135), .Z(n_26682));
	notech_inv i_30738(.A(n_28545), .Z(n_26683));
	notech_inv i_30739(.A(n_155075494), .Z(n_26684));
	notech_inv i_30740(.A(n_155175495), .Z(n_26685));
	notech_inv i_30741(.A(n_178175725), .Z(n_26686));
	notech_inv i_30742(.A(n_178875732), .Z(n_26687));
	notech_inv i_30743(.A(n_179575739), .Z(n_26688));
	notech_inv i_30744(.A(n_180275746), .Z(n_26689));
	notech_inv i_30746(.A(n_183375777), .Z(n_26690));
	notech_inv i_30747(.A(n_184075784), .Z(n_26691));
	notech_inv i_30748(.A(n_184775791), .Z(n_26692));
	notech_inv i_30753(.A(n_185475798), .Z(n_26693));
	notech_inv i_30757(.A(n_186175805), .Z(n_26694));
	notech_inv i_30758(.A(n_186875812), .Z(n_26695));
	notech_inv i_30759(.A(n_151328790), .Z(n_26696));
	notech_inv i_30761(.A(n_122175165), .Z(n_26697));
	notech_inv i_30762(.A(n_58163), .Z(n_26698));
	notech_inv i_30764(.A(n_215276091), .Z(n_26699));
	notech_inv i_30765(.A(n_105022314), .Z(n_26700));
	notech_inv i_30767(.A(n_217176110), .Z(n_26701));
	notech_inv i_30769(.A(n_1903), .Z(n_26702));
	notech_inv i_30770(.A(n_193865467), .Z(n_26704));
	notech_inv i_30772(.A(n_192365452), .Z(n_26705));
	notech_inv i_30773(.A(n_54974), .Z(n_26707));
	notech_inv i_30774(.A(n_121375157), .Z(n_26708));
	notech_inv i_30775(.A(n_215876097), .Z(n_26710));
	notech_inv i_30776(.A(n_57512), .Z(n_26711));
	notech_inv i_30777(.A(n_57121), .Z(n_26712));
	notech_inv i_30782(.A(n_24594), .Z(n_26718));
	notech_inv i_30783(.A(n_115978663), .Z(n_26719));
	notech_inv i_30784(.A(n_318891635), .Z(n_26720));
	notech_inv i_30785(.A(n_32280), .Z(n_26721));
	notech_inv i_30786(.A(n_329463511), .Z(n_26723));
	notech_inv i_30787(.A(n_3810), .Z(n_26724));
	notech_inv i_30788(.A(n_30366), .Z(n_26725));
	notech_inv i_30789(.A(n_3811), .Z(n_26727));
	notech_inv i_30790(.A(n_30301), .Z(n_26728));
	notech_inv i_30791(.A(n_130878812), .Z(n_26729));
	notech_inv i_30792(.A(n_131178815), .Z(n_26730));
	notech_inv i_30793(.A(n_58087), .Z(n_26731));
	notech_inv i_30795(.A(n_58325), .Z(n_26733));
	notech_inv i_30796(.A(n_135778861), .Z(n_26734));
	notech_inv i_30797(.A(n_32367), .Z(n_26735));
	notech_inv i_30798(.A(n_160979113), .Z(n_26736));
	notech_inv i_30799(.A(n_57249), .Z(n_26737));
	notech_inv i_30800(.A(n_161279116), .Z(n_26738));
	notech_inv i_30801(.A(n_158379087), .Z(n_26739));
	notech_inv i_30802(.A(n_161579119), .Z(n_26740));
	notech_inv i_30803(.A(n_162779131), .Z(n_26741));
	notech_inv i_30804(.A(n_163479138), .Z(n_26742));
	notech_inv i_30805(.A(n_164279146), .Z(n_26743));
	notech_inv i_30806(.A(n_164979153), .Z(n_26744));
	notech_inv i_30807(.A(n_154679050), .Z(n_26745));
	notech_inv i_30808(.A(n_158465113), .Z(n_26746));
	notech_inv i_30809(.A(n_156865097), .Z(n_26747));
	notech_inv i_30810(.A(n_301091813), .Z(n_26748));
	notech_inv i_30811(.A(n_113564664), .Z(n_26749));
	notech_inv i_30812(.A(n_112964658), .Z(n_26750));
	notech_inv i_30813(.A(n_113064659), .Z(n_26751));
	notech_inv i_30815(.A(n_54814), .Z(n_26753));
	notech_inv i_30816(.A(n_111264641), .Z(n_26754));
	notech_inv i_30817(.A(n_19022), .Z(n_26755));
	notech_inv i_30818(.A(n_19036), .Z(n_26756));
	notech_inv i_30819(.A(n_32605), .Z(n_26757));
	notech_inv i_30820(.A(n_32562), .Z(n_26758));
	notech_inv i_30821(.A(n_314863415), .Z(n_26759));
	notech_inv i_30822(.A(n_314663413), .Z(n_26760));
	notech_inv i_30823(.A(n_19127), .Z(n_26761));
	notech_inv i_30824(.A(n_309721261), .Z(n_26762));
	notech_inv i_30825(.A(n_281263079), .Z(n_26763));
	notech_inv i_30826(.A(n_209379594), .Z(n_26764));
	notech_inv i_30827(.A(n_122228499), .Z(n_26765));
	notech_inv i_30828(.A(n_122628503), .Z(n_26766));
	notech_inv i_30829(.A(n_26061), .Z(n_26767));
	notech_inv i_30831(.A(n_54718), .Z(n_26769));
	notech_inv i_30832(.A(n_30946), .Z(n_26770));
	notech_inv i_30833(.A(n_233679837), .Z(n_26771));
	notech_inv i_30834(.A(n_223979740), .Z(n_26772));
	notech_inv i_30835(.A(n_57616), .Z(n_26773));
	notech_inv i_30836(.A(n_58169), .Z(n_26774));
	notech_inv i_30837(.A(n_24589), .Z(n_26775));
	notech_inv i_30838(.A(n_125361536), .Z(n_26776));
	notech_inv i_30839(.A(n_215879659), .Z(n_26777));
	notech_inv i_30840(.A(n_144861731), .Z(n_26778));
	notech_inv i_30841(.A(n_57839), .Z(n_26779));
	notech_inv i_30842(.A(n_3812), .Z(n_26780));
	notech_inv i_30843(.A(n_330263519), .Z(n_26781));
	notech_inv i_30844(.A(n_57967), .Z(n_26782));
	notech_inv i_30845(.A(n_190262174), .Z(n_26783));
	notech_inv i_30846(.A(n_58806), .Z(n_26784));
	notech_inv i_30847(.A(n_329563512), .Z(n_26785));
	notech_inv i_30848(.A(n_56809), .Z(n_26789));
	notech_inv i_30849(.A(n_58132), .Z(n_26790));
	notech_inv i_30850(.A(n_54765), .Z(n_26791));
	notech_inv i_30851(.A(n_57926), .Z(n_26792));
	notech_inv i_30852(.A(n_249179992), .Z(n_26793));
	notech_inv i_30853(.A(n_255380054), .Z(n_26794));
	notech_inv i_30854(.A(n_256080061), .Z(n_26795));
	notech_inv i_30855(.A(n_256780068), .Z(n_26797));
	notech_inv i_30856(.A(n_257480075), .Z(n_26798));
	notech_inv i_30857(.A(n_58493), .Z(n_26800));
	notech_inv i_30858(.A(n_261780118), .Z(n_26801));
	notech_inv i_30859(.A(n_91719099), .Z(n_26802));
	notech_inv i_30860(.A(n_27340), .Z(n_26803));
	notech_inv i_30861(.A(n_58485), .Z(n_26804));
	notech_inv i_30862(.A(n_58486), .Z(n_26805));
	notech_inv i_30863(.A(n_266380164), .Z(n_26806));
	notech_inv i_30864(.A(n_56482), .Z(n_26807));
	notech_inv i_30865(.A(n_58488), .Z(n_26808));
	notech_inv i_30866(.A(n_58802), .Z(n_26809));
	notech_inv i_30867(.A(n_58078), .Z(n_26810));
	notech_inv i_30868(.A(n_58419), .Z(n_26811));
	notech_inv i_30869(.A(n_58490), .Z(n_26812));
	notech_inv i_30870(.A(n_58421), .Z(n_26813));
	notech_inv i_30871(.A(n_290580406), .Z(n_26814));
	notech_inv i_30872(.A(n_27344), .Z(n_26815));
	notech_inv i_30873(.A(n_58487), .Z(n_26816));
	notech_inv i_30874(.A(n_32350), .Z(n_26817));
	notech_inv i_30875(.A(n_316891655), .Z(n_26818));
	notech_inv i_30876(.A(n_58098), .Z(n_26819));
	notech_inv i_30877(.A(n_58097), .Z(n_26820));
	notech_inv i_30878(.A(n_58481), .Z(n_26821));
	notech_inv i_30880(.A(n_57808), .Z(n_26823));
	notech_inv i_30881(.A(n_58422), .Z(n_26824));
	notech_inv i_30882(.A(n_56803), .Z(n_26825));
	notech_inv i_30883(.A(n_58495), .Z(n_26826));
	notech_inv i_30884(.A(n_57927), .Z(n_26827));
	notech_inv i_30885(.A(n_58479), .Z(n_26828));
	notech_inv i_30886(.A(n_57505), .Z(n_26829));
	notech_inv i_30887(.A(n_332380824), .Z(n_26830));
	notech_inv i_30888(.A(n_312580626), .Z(n_26831));
	notech_inv i_30889(.A(n_316591658), .Z(n_26832));
	notech_inv i_30890(.A(n_297363240), .Z(n_26833));
	notech_inv i_30891(.A(n_54774), .Z(n_26834));
	notech_inv i_30892(.A(n_286663133), .Z(n_26835));
	notech_inv i_30893(.A(n_3829), .Z(n_26836));
	notech_inv i_30894(.A(n_3827), .Z(n_26837));
	notech_inv i_30895(.A(n_3813), .Z(n_26838));
	notech_inv i_30896(.A(n_341380914), .Z(n_26839));
	notech_inv i_30897(.A(n_30905), .Z(n_26840));
	notech_inv i_30898(.A(n_30359), .Z(n_26841));
	notech_inv i_30899(.A(n_282063087), .Z(n_26842));
	notech_inv i_30900(.A(n_58162), .Z(n_26843));
	notech_inv i_30901(.A(n_131578819), .Z(n_26844));
	notech_inv i_30902(.A(n_275063017), .Z(n_26845));
	notech_inv i_30903(.A(n_250140519), .Z(n_26846));
	notech_inv i_30905(.A(n_346280963), .Z(n_26847));
	notech_inv i_30906(.A(n_160079104), .Z(n_26849));
	notech_inv i_30908(.A(n_58377), .Z(n_26850));
	notech_inv i_30909(.A(n_58053), .Z(n_26851));
	notech_inv i_30910(.A(n_58164), .Z(n_26852));
	notech_inv i_30911(.A(n_58050), .Z(n_26853));
	notech_inv i_30912(.A(n_58051), .Z(n_26854));
	notech_inv i_30913(.A(n_57179), .Z(n_26855));
	notech_inv i_30914(.A(n_57180), .Z(n_26856));
	notech_inv i_30915(.A(n_290918108), .Z(n_26857));
	notech_inv i_30919(.A(n_340580906), .Z(n_26858));
	notech_inv i_30920(.A(n_345480955), .Z(n_26859));
	notech_inv i_30921(.A(n_320391620), .Z(n_26860));
	notech_inv i_30922(.A(n_110982110), .Z(n_26861));
	notech_inv i_30923(.A(n_123182232), .Z(n_26862));
	notech_inv i_30924(.A(n_123282233), .Z(n_26863));
	notech_inv i_30925(.A(n_123982240), .Z(n_26864));
	notech_inv i_30926(.A(n_124082241), .Z(n_26865));
	notech_inv i_30927(.A(n_124782248), .Z(n_26866));
	notech_inv i_30928(.A(n_124882249), .Z(n_26867));
	notech_inv i_30929(.A(n_125582256), .Z(n_26868));
	notech_inv i_30930(.A(n_125682257), .Z(n_26869));
	notech_inv i_30931(.A(n_126382264), .Z(n_26870));
	notech_inv i_30932(.A(n_126482265), .Z(n_26871));
	notech_inv i_30933(.A(n_127182272), .Z(n_26872));
	notech_inv i_30934(.A(n_127282273), .Z(n_26873));
	notech_inv i_30935(.A(n_127982280), .Z(n_26874));
	notech_inv i_30936(.A(n_128082281), .Z(n_26875));
	notech_inv i_30937(.A(n_128782288), .Z(n_26876));
	notech_inv i_30938(.A(n_128882289), .Z(n_26877));
	notech_inv i_30939(.A(n_129582296), .Z(n_26878));
	notech_inv i_30940(.A(n_129682297), .Z(n_26879));
	notech_inv i_30941(.A(n_315191672), .Z(n_26880));
	notech_inv i_30942(.A(n_132182322), .Z(n_26881));
	notech_inv i_30943(.A(n_57758), .Z(n_26882));
	notech_inv i_30944(.A(n_74438764), .Z(n_26883));
	notech_inv i_30945(.A(n_54736), .Z(n_26884));
	notech_inv i_30946(.A(n_76638786), .Z(n_26885));
	notech_inv i_30947(.A(n_76238782), .Z(n_26886));
	notech_inv i_30948(.A(n_30961), .Z(n_26887));
	notech_inv i_30949(.A(n_30937), .Z(n_26888));
	notech_inv i_30950(.A(n_30966), .Z(n_26889));
	notech_inv i_30951(.A(n_28551), .Z(n_26890));
	notech_inv i_30952(.A(n_28120), .Z(n_26891));
	notech_inv i_30953(.A(n_28132), .Z(n_26892));
	notech_inv i_30954(.A(n_143682437), .Z(n_26893));
	notech_inv i_30955(.A(n_30352), .Z(n_26894));
	notech_inv i_30956(.A(n_57602), .Z(n_26895));
	notech_inv i_30957(.A(n_145182452), .Z(n_26896));
	notech_inv i_30958(.A(n_145382454), .Z(n_26897));
	notech_inv i_30959(.A(n_30930), .Z(n_26898));
	notech_inv i_30960(.A(n_29967), .Z(n_26899));
	notech_inv i_30961(.A(n_32586), .Z(n_26900));
	notech_inv i_30962(.A(n_137382374), .Z(n_26901));
	notech_inv i_30963(.A(n_58144), .Z(n_26902));
	notech_inv i_30964(.A(n_155282553), .Z(n_26903));
	notech_inv i_30965(.A(n_58646), .Z(n_26904));
	notech_inv i_30966(.A(n_58610), .Z(n_26905));
	notech_inv i_30967(.A(n_58167), .Z(n_26906));
	notech_inv i_30968(.A(n_58489), .Z(n_26908));
	notech_inv i_30969(.A(n_180682807), .Z(n_26910));
	notech_inv i_30970(.A(n_226362530), .Z(n_26911));
	notech_inv i_30971(.A(n_206683057), .Z(n_26912));
	notech_inv i_30972(.A(n_206783058), .Z(n_26913));
	notech_inv i_30973(.A(n_206883059), .Z(n_26915));
	notech_inv i_30974(.A(n_58498), .Z(n_26916));
	notech_inv i_30975(.A(n_58146), .Z(n_26918));
	notech_inv i_30976(.A(n_32292), .Z(n_26920));
	notech_inv i_30977(.A(n_58497), .Z(n_26921));
	notech_inv i_30978(.A(n_32301), .Z(n_26922));
	notech_inv i_30979(.A(n_32304), .Z(n_26924));
	notech_inv i_30980(.A(n_32408), .Z(n_26925));
	notech_inv i_30981(.A(n_32295), .Z(n_26927));
	notech_inv i_30982(.A(n_32284), .Z(n_26928));
	notech_inv i_30983(.A(n_58148), .Z(n_26929));
	notech_inv i_30984(.A(n_32291), .Z(n_26933));
	notech_inv i_30985(.A(n_57569), .Z(n_26937));
	notech_inv i_30986(.A(n_25010), .Z(n_26938));
	notech_inv i_30987(.A(n_25007), .Z(n_26939));
	notech_inv i_30988(.A(n_242983420), .Z(n_26940));
	notech_inv i_30989(.A(n_23512), .Z(n_26941));
	notech_inv i_30990(.A(n_23510), .Z(n_26942));
	notech_inv i_30991(.A(n_243883429), .Z(n_26943));
	notech_inv i_30992(.A(n_243983430), .Z(n_26944));
	notech_inv i_30993(.A(n_54794), .Z(n_26945));
	notech_inv i_30995(.A(n_175362036), .Z(n_26947));
	notech_inv i_30996(.A(n_18912289), .Z(n_26948));
	notech_inv i_30997(.A(n_19512295), .Z(n_26949));
	notech_inv i_30998(.A(n_32318), .Z(n_26950));
	notech_inv i_30999(.A(n_169561978), .Z(n_26951));
	notech_inv i_31000(.A(n_168861971), .Z(n_26952));
	notech_inv i_31001(.A(n_160061883), .Z(n_26953));
	notech_inv i_31003(.A(n_168561968), .Z(n_26954));
	notech_inv i_31004(.A(n_168361966), .Z(n_26955));
	notech_inv i_31006(.A(n_152561808), .Z(n_26958));
	notech_inv i_31007(.A(n_24583), .Z(n_26960));
	notech_inv i_31008(.A(n_131461597), .Z(n_26961));
	notech_inv i_31009(.A(n_32384), .Z(n_26962));
	notech_inv i_31010(.A(n_19043), .Z(n_26963));
	notech_inv i_31011(.A(n_19057), .Z(n_26964));
	notech_inv i_31013(.A(n_25374), .Z(n_26965));
	notech_inv i_31014(.A(n_148261765), .Z(n_26966));
	notech_inv i_31015(.A(n_17409952), .Z(n_26967));
	notech_inv i_31016(.A(n_30931), .Z(n_26968));
	notech_inv i_31017(.A(n_32298), .Z(n_26969));
	notech_inv i_31018(.A(n_30350), .Z(n_26970));
	notech_inv i_31019(.A(n_30342), .Z(n_26971));
	notech_inv i_31020(.A(n_30357), .Z(n_26972));
	notech_inv i_31021(.A(n_30322), .Z(n_26973));
	notech_inv i_31022(.A(n_317784168), .Z(n_26974));
	notech_inv i_31023(.A(n_143861721), .Z(n_26975));
	notech_inv i_31024(.A(n_142761710), .Z(n_26976));
	notech_inv i_31025(.A(n_142461707), .Z(n_26977));
	notech_inv i_31026(.A(n_323984230), .Z(n_26978));
	notech_inv i_31027(.A(n_141161694), .Z(n_26979));
	notech_inv i_31028(.A(n_138561668), .Z(n_26980));
	notech_inv i_31029(.A(n_129561578), .Z(n_26981));
	notech_inv i_31030(.A(n_130361586), .Z(n_26982));
	notech_inv i_31031(.A(n_60283), .Z(n_26983));
	notech_inv i_31032(.A(n_58088), .Z(n_26984));
	notech_inv i_31033(.A(n_19079), .Z(n_26985));
	notech_inv i_31034(.A(n_54865), .Z(n_26986));
	notech_inv i_31036(.A(n_109682097), .Z(n_26988));
	notech_inv i_31037(.A(n_18989), .Z(n_26989));
	notech_inv i_31038(.A(n_60074), .Z(n_26990));
	notech_inv i_31039(.A(n_3915), .Z(n_26991));
	notech_inv i_31040(.A(n_3819), .Z(n_26992));
	notech_inv i_31041(.A(n_346670477), .Z(n_26993));
	notech_inv i_31042(.A(n_46630), .Z(n_26994));
	notech_inv i_31043(.A(n_3900), .Z(n_26995));
	notech_inv i_31044(.A(n_3899), .Z(n_26996));
	notech_inv i_31045(.A(n_3898), .Z(n_26997));
	notech_inv i_31046(.A(n_3897), .Z(n_26998));
	notech_inv i_31047(.A(n_19050), .Z(n_26999));
	notech_inv i_31048(.A(n_3896), .Z(n_27000));
	notech_inv i_31049(.A(n_55800), .Z(n_27001));
	notech_inv i_31050(.A(n_3886), .Z(n_27002));
	notech_inv i_31051(.A(n_55891), .Z(n_27003));
	notech_inv i_31053(.A(n_3872), .Z(n_27005));
	notech_inv i_31054(.A(n_3871), .Z(n_27006));
	notech_inv i_31055(.A(n_106985346), .Z(n_27007));
	notech_inv i_31056(.A(n_114785424), .Z(n_27008));
	notech_inv i_31057(.A(n_115685433), .Z(n_27009));
	notech_inv i_31058(.A(n_116585442), .Z(n_27010));
	notech_inv i_31059(.A(n_3863), .Z(n_27011));
	notech_inv i_31060(.A(n_117485451), .Z(n_27012));
	notech_inv i_31061(.A(n_118385460), .Z(n_27013));
	notech_inv i_31062(.A(n_119285469), .Z(n_27014));
	notech_inv i_31063(.A(n_3860), .Z(n_27015));
	notech_inv i_31064(.A(n_120185478), .Z(n_27016));
	notech_inv i_31065(.A(n_121085487), .Z(n_27017));
	notech_inv i_31066(.A(n_121985496), .Z(n_27018));
	notech_inv i_31067(.A(n_238359464), .Z(n_27019));
	notech_inv i_31068(.A(n_231559396), .Z(n_27020));
	notech_inv i_31069(.A(n_122885505), .Z(n_27021));
	notech_inv i_31070(.A(n_225459335), .Z(n_27022));
	notech_inv i_31071(.A(n_3853), .Z(n_27023));
	notech_inv i_31072(.A(n_305291771), .Z(n_27024));
	notech_inv i_31073(.A(n_3596), .Z(n_27025));
	notech_inv i_31074(.A(n_3847), .Z(n_27026));
	notech_inv i_31075(.A(n_3840), .Z(n_27027));
	notech_inv i_31076(.A(n_3839), .Z(n_27028));
	notech_inv i_31077(.A(n_3834), .Z(n_27029));
	notech_inv i_31078(.A(n_60933), .Z(\opcode[2] ));
	notech_inv i_31079(.A(n_3832), .Z(n_27031));
	notech_inv i_31082(.A(n_3824), .Z(n_27033));
	notech_inv i_31083(.A(n_3823), .Z(n_27034));
	notech_inv i_31084(.A(n_3822), .Z(n_27035));
	notech_inv i_31085(.A(n_32616), .Z(n_27036));
	notech_inv i_31086(.A(n_3796), .Z(n_27037));
	notech_inv i_31087(.A(n_3787), .Z(n_27038));
	notech_inv i_31090(.A(n_3776), .Z(n_27039));
	notech_inv i_31091(.A(n_144385720), .Z(n_27040));
	notech_inv i_31092(.A(n_3628), .Z(n_27041));
	notech_inv i_31093(.A(n_3724), .Z(n_27042));
	notech_inv i_31094(.A(n_3714), .Z(n_27043));
	notech_inv i_31095(.A(n_315891665), .Z(n_27044));
	notech_inv i_31096(.A(n_3672), .Z(n_27045));
	notech_inv i_31097(.A(n_3632), .Z(n_27046));
	notech_inv i_31098(.A(n_209886372), .Z(n_27047));
	notech_inv i_31099(.A(n_213886412), .Z(n_27048));
	notech_inv i_31100(.A(n_212886402), .Z(n_27049));
	notech_inv i_31101(.A(n_58697), .Z(n_27050));
	notech_inv i_31102(.A(n_290618105), .Z(n_27051));
	notech_inv i_31103(.A(n_18964), .Z(n_27052));
	notech_inv i_31108(.A(n_58675), .Z(n_27053));
	notech_inv i_31112(.A(n_57406), .Z(n_27054));
	notech_inv i_31113(.A(n_269686970), .Z(n_27055));
	notech_inv i_31114(.A(n_57899), .Z(n_27056));
	notech_inv i_31116(.A(n_342991444), .Z(n_27057));
	notech_inv i_31117(.A(n_342591448), .Z(n_27058));
	notech_inv i_31119(.A(n_342491449), .Z(n_27059));
	notech_inv i_31120(.A(n_341191462), .Z(n_27060));
	notech_inv i_31121(.A(n_305191772), .Z(n_27061));
	notech_inv i_31123(.A(n_312960210), .Z(n_27062));
	notech_inv i_31125(.A(n_58812), .Z(n_27063));
	notech_inv i_31126(.A(n_19006), .Z(n_27065));
	notech_inv i_31128(.A(n_55378), .Z(n_27066));
	notech_inv i_31130(.A(n_18972), .Z(n_27068));
	notech_inv i_31131(.A(n_32551), .Z(n_27069));
	notech_inv i_31133(.A(n_320191622), .Z(n_27070));
	notech_inv i_31135(.A(n_296760048), .Z(n_27071));
	notech_inv i_31136(.A(n_287959960), .Z(n_27072));
	notech_inv i_31139(.A(n_4005), .Z(n_27075));
	notech_inv i_31140(.A(n_277959860), .Z(n_27076));
	notech_inv i_31141(.A(n_53174), .Z(n_27077));
	notech_inv i_31142(.A(n_256290061), .Z(n_27078));
	notech_inv i_31143(.A(n_305891765), .Z(n_27079));
	notech_inv i_31144(.A(n_267459755), .Z(n_27080));
	notech_inv i_31145(.A(n_53252), .Z(n_27081));
	notech_inv i_31146(.A(n_256459645), .Z(n_27082));
	notech_inv i_31147(.A(n_255659637), .Z(n_27083));
	notech_inv i_31148(.A(n_32272), .Z(n_27084));
	notech_inv i_31149(.A(n_317291651), .Z(n_27085));
	notech_inv i_31150(.A(n_60986), .Z(\opcode[3] ));
	notech_inv i_31151(.A(n_60874), .Z(\opcode[0] ));
	notech_inv i_31153(.A(n_32335), .Z(n_27089));
	notech_inv i_31154(.A(n_3919), .Z(n_27090));
	notech_inv i_31156(.A(n_40675), .Z(n_27092));
	notech_inv i_31158(.A(n_32319), .Z(n_27094));
	notech_inv i_31159(.A(n_27922), .Z(n_27095));
	notech_inv i_31160(.A(n_27880), .Z(n_27096));
	notech_inv i_31161(.A(n_58666), .Z(n_27097));
	notech_inv i_31162(.A(n_243459515), .Z(n_27098));
	notech_inv i_31163(.A(n_242759508), .Z(n_27099));
	notech_inv i_31164(.A(n_224759328), .Z(n_27100));
	notech_inv i_31165(.A(n_186058956), .Z(n_27101));
	notech_inv i_31166(.A(n_313491689), .Z(n_27102));
	notech_inv i_31167(.A(n_183958935), .Z(n_27103));
	notech_inv i_31168(.A(n_32323), .Z(n_27104));
	notech_inv i_31169(.A(n_55820), .Z(n_27105));
	notech_inv i_31170(.A(n_58691), .Z(n_27106));
	notech_inv i_31171(.A(n_3922), .Z(n_27107));
	notech_inv i_31172(.A(n_177558871), .Z(n_27108));
	notech_inv i_31173(.A(n_312091703), .Z(n_27109));
	notech_inv i_31174(.A(n_319291631), .Z(n_27110));
	notech_inv i_31175(.A(n_45891243), .Z(n_27111));
	notech_inv i_31176(.A(fsmf[4]), .Z(n_27112));
	notech_inv i_31177(.A(n_6858899), .Z(n_27113));
	notech_inv i_31178(.A(\nbus_11351[0] ), .Z(n_27114));
	notech_inv i_31179(.A(n_13782), .Z(n_27115));
	notech_inv i_31180(.A(sav_ecx[0]), .Z(n_27116));
	notech_inv i_31181(.A(sav_ecx[1]), .Z(n_27117));
	notech_inv i_31182(.A(sav_ecx[2]), .Z(n_27118));
	notech_inv i_31183(.A(n_28552), .Z(n_27119));
	notech_inv i_31184(.A(sav_ecx[3]), .Z(n_27120));
	notech_inv i_31185(.A(sav_ecx[4]), .Z(n_27121));
	notech_inv i_31186(.A(sav_ecx[5]), .Z(n_27122));
	notech_inv i_31187(.A(n_32695), .Z(n_27123));
	notech_inv i_31188(.A(sav_ecx[6]), .Z(n_27124));
	notech_inv i_31189(.A(n_32470), .Z(n_27125));
	notech_inv i_31190(.A(sav_ecx[7]), .Z(n_27126));
	notech_inv i_31191(.A(sav_ecx[8]), .Z(n_27127));
	notech_inv i_31192(.A(n_272291903), .Z(n_27128));
	notech_inv i_31194(.A(sav_ecx[9]), .Z(n_27129));
	notech_inv i_31195(.A(sav_ecx[10]), .Z(n_27130));
	notech_inv i_31196(.A(sav_ecx[11]), .Z(n_27131));
	notech_inv i_31197(.A(n_2838), .Z(n_27132));
	notech_inv i_31198(.A(sav_ecx[12]), .Z(n_27133));
	notech_inv i_31199(.A(sav_ecx[13]), .Z(n_27134));
	notech_inv i_31200(.A(sav_ecx[14]), .Z(n_27135));
	notech_inv i_31201(.A(sav_ecx[15]), .Z(n_27136));
	notech_inv i_31202(.A(sav_ecx[17]), .Z(n_27137));
	notech_inv i_31203(.A(sav_ecx[18]), .Z(n_27138));
	notech_inv i_31204(.A(sav_ecx[19]), .Z(n_27139));
	notech_inv i_31205(.A(sav_ecx[20]), .Z(n_27140));
	notech_inv i_31206(.A(sav_ecx[21]), .Z(n_27141));
	notech_inv i_31208(.A(sav_ecx[22]), .Z(n_27144));
	notech_inv i_31209(.A(n_2880), .Z(n_27145));
	notech_inv i_31210(.A(sav_ecx[23]), .Z(n_27146));
	notech_inv i_31211(.A(sav_ecx[24]), .Z(n_27147));
	notech_inv i_31212(.A(sav_ecx[25]), .Z(n_27148));
	notech_inv i_31213(.A(sav_ecx[27]), .Z(n_27149));
	notech_inv i_31214(.A(sav_ecx[28]), .Z(n_27150));
	notech_inv i_31215(.A(sav_ecx[31]), .Z(n_27151));
	notech_inv i_31216(.A(n_14391), .Z(n_27152));
	notech_inv i_31217(.A(sav_esp[0]), .Z(n_27153));
	notech_inv i_31218(.A(sav_esp[1]), .Z(n_27154));
	notech_inv i_31219(.A(n_60904), .Z(\opcode[1] ));
	notech_inv i_31220(.A(sav_esp[2]), .Z(n_27156));
	notech_inv i_31221(.A(sav_esp[3]), .Z(n_27158));
	notech_inv i_31222(.A(sav_esp[4]), .Z(n_27159));
	notech_inv i_31223(.A(sav_esp[5]), .Z(n_27160));
	notech_inv i_31224(.A(sav_esp[6]), .Z(n_27161));
	notech_inv i_31225(.A(sav_esp[7]), .Z(n_27162));
	notech_inv i_31226(.A(sav_esp[8]), .Z(n_27164));
	notech_inv i_31227(.A(sav_esp[9]), .Z(n_27165));
	notech_inv i_31228(.A(sav_esp[10]), .Z(n_27166));
	notech_inv i_31229(.A(sav_esp[11]), .Z(n_27167));
	notech_inv i_31230(.A(sav_esp[12]), .Z(n_27168));
	notech_inv i_31231(.A(sav_esp[14]), .Z(n_27169));
	notech_inv i_31232(.A(n_2864), .Z(n_27170));
	notech_inv i_31233(.A(sav_esp[16]), .Z(n_27171));
	notech_inv i_31234(.A(sav_esp[17]), .Z(n_27172));
	notech_inv i_31235(.A(sav_esp[18]), .Z(n_27173));
	notech_inv i_31236(.A(n_320091623), .Z(n_27174));
	notech_inv i_31237(.A(sav_esp[19]), .Z(n_27175));
	notech_inv i_31238(.A(sav_esp[21]), .Z(n_27176));
	notech_inv i_31239(.A(n_317591648), .Z(n_27177));
	notech_inv i_31240(.A(sav_esp[22]), .Z(n_27178));
	notech_inv i_31242(.A(n_319891625), .Z(n_27179));
	notech_inv i_31243(.A(sav_esp[23]), .Z(n_27181));
	notech_inv i_31245(.A(sav_esp[24]), .Z(n_27182));
	notech_inv i_31246(.A(sav_esp[25]), .Z(n_27183));
	notech_inv i_31247(.A(sav_esp[26]), .Z(n_27184));
	notech_inv i_31248(.A(sav_esp[28]), .Z(n_27185));
	notech_inv i_31249(.A(sav_esp[29]), .Z(n_27186));
	notech_inv i_31250(.A(sav_esp[30]), .Z(n_27187));
	notech_inv i_31252(.A(sav_esp[31]), .Z(n_27188));
	notech_inv i_31255(.A(sav_esi[1]), .Z(n_27189));
	notech_inv i_31256(.A(sav_esi[3]), .Z(n_27190));
	notech_inv i_31257(.A(sav_esi[4]), .Z(n_27191));
	notech_inv i_31258(.A(n_319091633), .Z(n_27192));
	notech_inv i_31259(.A(sav_esi[5]), .Z(n_27193));
	notech_inv i_31260(.A(n_317391650), .Z(n_27194));
	notech_inv i_31261(.A(sav_esi[6]), .Z(n_27195));
	notech_inv i_31262(.A(n_318991634), .Z(n_27196));
	notech_inv i_31263(.A(sav_esi[7]), .Z(n_27197));
	notech_inv i_31264(.A(n_318791636), .Z(n_27198));
	notech_inv i_31265(.A(sav_esi[10]), .Z(n_27199));
	notech_inv i_31266(.A(sav_esi[11]), .Z(n_27200));
	notech_inv i_31267(.A(sav_esi[12]), .Z(n_27201));
	notech_inv i_31268(.A(sav_esi[13]), .Z(n_27202));
	notech_inv i_31269(.A(sav_esi[14]), .Z(n_27203));
	notech_inv i_31270(.A(sav_esi[15]), .Z(n_27204));
	notech_inv i_31271(.A(sav_esi[16]), .Z(n_27205));
	notech_inv i_31272(.A(sav_esi[17]), .Z(n_27206));
	notech_inv i_31273(.A(sav_esi[18]), .Z(n_27207));
	notech_inv i_31274(.A(sav_esi[19]), .Z(n_27208));
	notech_inv i_31275(.A(sav_esi[20]), .Z(n_27209));
	notech_inv i_31276(.A(sav_esi[21]), .Z(n_27210));
	notech_inv i_31277(.A(sav_esi[22]), .Z(n_27211));
	notech_inv i_31278(.A(sav_esi[23]), .Z(n_27212));
	notech_inv i_31279(.A(sav_esi[24]), .Z(n_27213));
	notech_inv i_31280(.A(sav_esi[25]), .Z(n_27214));
	notech_inv i_31281(.A(sav_esi[27]), .Z(n_27215));
	notech_inv i_31282(.A(sav_esi[30]), .Z(n_27216));
	notech_inv i_31283(.A(sav_esi[31]), .Z(n_27217));
	notech_inv i_31284(.A(sav_edi[1]), .Z(n_27218));
	notech_inv i_31285(.A(sav_edi[3]), .Z(n_27219));
	notech_inv i_31286(.A(sav_edi[4]), .Z(n_27220));
	notech_inv i_31287(.A(n_314891675), .Z(n_27221));
	notech_inv i_31288(.A(sav_edi[5]), .Z(n_27222));
	notech_inv i_31289(.A(sav_edi[6]), .Z(n_27223));
	notech_inv i_31290(.A(sav_edi[7]), .Z(n_27224));
	notech_inv i_31291(.A(sav_edi[9]), .Z(n_27225));
	notech_inv i_31292(.A(sav_edi[10]), .Z(n_27226));
	notech_inv i_31293(.A(sav_edi[11]), .Z(n_27227));
	notech_inv i_31294(.A(sav_edi[12]), .Z(n_27228));
	notech_inv i_31295(.A(sav_edi[13]), .Z(n_27229));
	notech_inv i_31296(.A(sav_edi[14]), .Z(n_27230));
	notech_inv i_31297(.A(sav_edi[15]), .Z(n_27231));
	notech_inv i_31298(.A(sav_edi[16]), .Z(n_27232));
	notech_inv i_31299(.A(n_314491679), .Z(n_27233));
	notech_inv i_31300(.A(sav_edi[17]), .Z(n_27234));
	notech_inv i_31301(.A(sav_edi[18]), .Z(n_27235));
	notech_inv i_31302(.A(sav_edi[19]), .Z(n_27236));
	notech_inv i_31303(.A(sav_edi[20]), .Z(n_27237));
	notech_inv i_31304(.A(sav_edi[21]), .Z(n_27238));
	notech_inv i_31305(.A(sav_edi[22]), .Z(n_27239));
	notech_inv i_31306(.A(sav_edi[23]), .Z(n_27240));
	notech_inv i_31307(.A(sav_edi[24]), .Z(n_27241));
	notech_inv i_31308(.A(sav_edi[25]), .Z(n_27242));
	notech_inv i_31309(.A(sav_edi[27]), .Z(n_27243));
	notech_inv i_31310(.A(sav_edi[30]), .Z(n_27244));
	notech_inv i_31311(.A(sav_edi[31]), .Z(n_27245));
	notech_inv i_31312(.A(fepc), .Z(n_27246));
	notech_inv i_31313(.A(sav_epc[1]), .Z(n_27247));
	notech_inv i_31314(.A(sav_epc[3]), .Z(n_27248));
	notech_inv i_31315(.A(sav_epc[4]), .Z(n_27249));
	notech_inv i_31316(.A(sav_epc[5]), .Z(n_27250));
	notech_inv i_31317(.A(sav_epc[6]), .Z(n_27251));
	notech_inv i_31318(.A(sav_epc[7]), .Z(n_27252));
	notech_inv i_31319(.A(sav_epc[11]), .Z(n_27253));
	notech_inv i_31320(.A(sav_epc[13]), .Z(n_27254));
	notech_inv i_31321(.A(sav_epc[14]), .Z(n_27255));
	notech_inv i_31322(.A(sav_epc[16]), .Z(n_27256));
	notech_inv i_31323(.A(n_308391740), .Z(n_27257));
	notech_inv i_31324(.A(sav_epc[17]), .Z(n_27258));
	notech_inv i_31325(.A(n_304791776), .Z(n_27259));
	notech_inv i_31326(.A(sav_epc[18]), .Z(n_27260));
	notech_inv i_31327(.A(sav_epc[19]), .Z(n_27261));
	notech_inv i_31328(.A(sav_epc[20]), .Z(n_27262));
	notech_inv i_31330(.A(sav_epc[21]), .Z(n_27263));
	notech_inv i_31331(.A(sav_epc[22]), .Z(n_27264));
	notech_inv i_31332(.A(sav_epc[23]), .Z(n_27265));
	notech_inv i_31333(.A(sav_epc[24]), .Z(n_27266));
	notech_inv i_31334(.A(sav_epc[25]), .Z(n_27267));
	notech_inv i_31335(.A(n_1670), .Z(n_27268));
	notech_inv i_31336(.A(sav_epc[31]), .Z(n_27269));
	notech_inv i_31337(.A(\nbus_11311[0] ), .Z(n_27270));
	notech_inv i_31338(.A(n_12888), .Z(n_27271));
	notech_inv i_31340(.A(n_306491759), .Z(n_27272));
	notech_inv i_31341(.A(n_307791746), .Z(n_27273));
	notech_inv i_31342(.A(n_307491749), .Z(n_27274));
	notech_inv i_31343(.A(n_24430), .Z(n_27275));
	notech_inv i_31344(.A(n_24478), .Z(n_27276));
	notech_inv i_31345(.A(n_24484), .Z(n_27277));
	notech_inv i_31346(.A(n_24490), .Z(n_27278));
	notech_inv i_31347(.A(n_24502), .Z(n_27279));
	notech_inv i_31348(.A(n_303891785), .Z(n_27280));
	notech_inv i_31349(.A(n_24520), .Z(n_27281));
	notech_inv i_31350(.A(n_24526), .Z(n_27282));
	notech_inv i_31351(.A(n_24532), .Z(n_27283));
	notech_inv i_31352(.A(n_24538), .Z(n_27284));
	notech_inv i_31353(.A(n_24544), .Z(n_27285));
	notech_inv i_31354(.A(n_24550), .Z(n_27286));
	notech_inv i_31355(.A(n_24556), .Z(n_27287));
	notech_inv i_31356(.A(n_24562), .Z(n_27288));
	notech_inv i_31357(.A(n_302791796), .Z(n_27289));
	notech_inv i_31358(.A(n_24568), .Z(n_27290));
	notech_inv i_31359(.A(n_24574), .Z(n_27291));
	notech_inv i_31360(.A(n_24580), .Z(n_27292));
	notech_inv i_31361(.A(n_302191802), .Z(n_27293));
	notech_inv i_31362(.A(n_24610), .Z(n_27294));
	notech_inv i_31363(.A(n_24616), .Z(n_27295));
	notech_inv i_31364(.A(n_24082), .Z(n_27296));
	notech_inv i_31365(.A(n_301591808), .Z(n_27297));
	notech_inv i_31366(.A(n_301491809), .Z(n_27298));
	notech_inv i_31367(.A(n_24118), .Z(n_27299));
	notech_inv i_31368(.A(n_301291811), .Z(n_27300));
	notech_inv i_31369(.A(n_299891825), .Z(n_27301));
	notech_inv i_31370(.A(n_300491819), .Z(n_27302));
	notech_inv i_31371(.A(n_24178), .Z(n_27303));
	notech_inv i_31372(.A(n_299691827), .Z(n_27304));
	notech_inv i_31373(.A(n_299491829), .Z(n_27305));
	notech_inv i_31374(.A(n_2988), .Z(n_27306));
	notech_inv i_31375(.A(n_24262), .Z(n_27307));
	notech_inv i_31376(.A(n_23734), .Z(n_27308));
	notech_inv i_31377(.A(n_23770), .Z(n_27309));
	notech_inv i_31378(.A(n_23782), .Z(n_27310));
	notech_inv i_31379(.A(n_23788), .Z(n_27311));
	notech_inv i_31380(.A(n_23794), .Z(n_27312));
	notech_inv i_31381(.A(n_23806), .Z(n_27313));
	notech_inv i_31382(.A(n_23824), .Z(n_27314));
	notech_inv i_31383(.A(n_23830), .Z(n_27315));
	notech_inv i_31384(.A(n_23836), .Z(n_27316));
	notech_inv i_31385(.A(n_23842), .Z(n_27317));
	notech_inv i_31386(.A(n_23848), .Z(n_27318));
	notech_inv i_31387(.A(n_23854), .Z(n_27320));
	notech_inv i_31388(.A(n_23860), .Z(n_27321));
	notech_inv i_31389(.A(n_13974), .Z(n_27322));
	notech_inv i_31390(.A(n_14022), .Z(n_27323));
	notech_inv i_31391(.A(n_14028), .Z(n_27324));
	notech_inv i_31392(.A(n_14034), .Z(n_27325));
	notech_inv i_31393(.A(n_14046), .Z(n_27326));
	notech_inv i_31394(.A(n_14064), .Z(n_27327));
	notech_inv i_31395(.A(n_14070), .Z(n_27328));
	notech_inv i_31396(.A(n_14076), .Z(n_27330));
	notech_inv i_31397(.A(n_14082), .Z(n_27331));
	notech_inv i_31398(.A(n_14088), .Z(n_27332));
	notech_inv i_31399(.A(n_14100), .Z(n_27333));
	notech_inv i_31400(.A(n_18829), .Z(n_27336));
	notech_inv i_31401(.A(n_18841), .Z(n_27337));
	notech_inv i_31402(.A(n_18883), .Z(n_27338));
	notech_inv i_31403(.A(n_18949), .Z(n_27339));
	notech_inv i_31404(.A(n_18961), .Z(n_27341));
	notech_inv i_31405(.A(n_18967), .Z(n_27342));
	notech_inv i_31407(.A(n_18973), .Z(n_27343));
	notech_inv i_31408(.A(n_18979), .Z(n_27345));
	notech_inv i_31409(.A(n_19009), .Z(n_27347));
	notech_inv i_31410(.A(n_19015), .Z(n_27350));
	notech_inv i_31411(.A(n_18480), .Z(n_27351));
	notech_inv i_31412(.A(n_291691848), .Z(n_27352));
	notech_inv i_31413(.A(n_18516), .Z(n_27354));
	notech_inv i_31414(.A(n_18528), .Z(n_27355));
	notech_inv i_31415(.A(n_18534), .Z(n_27356));
	notech_inv i_31416(.A(n_18540), .Z(n_27357));
	notech_inv i_31417(.A(n_18552), .Z(n_27358));
	notech_inv i_31418(.A(n_18570), .Z(n_27359));
	notech_inv i_31419(.A(n_18576), .Z(n_27360));
	notech_inv i_31420(.A(n_18582), .Z(n_27361));
	notech_inv i_31421(.A(n_18588), .Z(n_27362));
	notech_inv i_31422(.A(n_18594), .Z(n_27363));
	notech_inv i_31424(.A(n_18606), .Z(n_27364));
	notech_inv i_31425(.A(\nbus_11334[0] ), .Z(n_27365));
	notech_inv i_31426(.A(n_21336), .Z(n_27366));
	notech_inv i_31427(.A(n_21348), .Z(n_27367));
	notech_inv i_31428(.A(n_21372), .Z(n_27368));
	notech_inv i_31429(.A(n_21390), .Z(n_27369));
	notech_inv i_31430(.A(n_21402), .Z(n_27370));
	notech_inv i_31431(.A(n_21414), .Z(n_27371));
	notech_inv i_31433(.A(n_21420), .Z(n_27372));
	notech_inv i_31434(.A(n_21426), .Z(n_27373));
	notech_inv i_31435(.A(n_21432), .Z(n_27374));
	notech_inv i_31436(.A(n_21522), .Z(n_27375));
	notech_inv i_31437(.A(pipe_mul[0]), .Z(n_27376));
	notech_inv i_31438(.A(eval_flag), .Z(n_27377));
	notech_inv i_31439(.A(rep_en1), .Z(n_27378));
	notech_inv i_31440(.A(n_14570), .Z(n_27379));
	notech_inv i_31441(.A(rep_en4), .Z(n_27380));
	notech_inv i_31442(.A(nCF), .Z(n_27381));
	notech_inv i_31443(.A(nAF), .Z(n_27382));
	notech_inv i_31444(.A(nSF), .Z(n_27383));
	notech_inv i_31445(.A(n_21654), .Z(n_27384));
	notech_inv i_31446(.A(nOF), .Z(n_27385));
	notech_inv i_31447(.A(n_21651), .Z(n_27386));
	notech_inv i_31448(.A(n_25246), .Z(n_27387));
	notech_inv i_31449(.A(n_25294), .Z(n_27388));
	notech_inv i_31450(.A(n_25300), .Z(n_27389));
	notech_inv i_31452(.A(\nbus_11376[9] ), .Z(n_27390));
	notech_inv i_31453(.A(n_25306), .Z(n_27391));
	notech_inv i_31454(.A(\nbus_11376[10] ), .Z(n_27392));
	notech_inv i_31455(.A(\nbus_11376[6] ), .Z(n_27393));
	notech_inv i_31456(.A(n_25318), .Z(n_27394));
	notech_inv i_31457(.A(n_25324), .Z(n_27395));
	notech_inv i_31458(.A(n_25330), .Z(n_27396));
	notech_inv i_31459(.A(n_25336), .Z(n_27397));
	notech_inv i_31460(.A(n_25348), .Z(n_27398));
	notech_inv i_31461(.A(n_25354), .Z(n_27399));
	notech_inv i_31462(.A(n_25360), .Z(n_27400));
	notech_inv i_31463(.A(n_25372), .Z(n_27401));
	notech_inv i_31464(.A(n_25432), .Z(n_27402));
	notech_inv i_31465(.A(n_18132), .Z(n_27403));
	notech_inv i_31466(.A(n_18144), .Z(n_27404));
	notech_inv i_31467(.A(n_18174), .Z(n_27405));
	notech_inv i_31468(.A(n_18210), .Z(n_27406));
	notech_inv i_31469(.A(n_18216), .Z(n_27407));
	notech_inv i_31470(.A(n_18318), .Z(n_27408));
	notech_inv i_31471(.A(n_17780), .Z(n_27409));
	notech_inv i_31472(.A(n_17792), .Z(n_27410));
	notech_inv i_31473(.A(n_17828), .Z(n_27411));
	notech_inv i_31474(.A(n_17834), .Z(n_27412));
	notech_inv i_31475(.A(n_17840), .Z(n_27413));
	notech_inv i_31476(.A(n_17852), .Z(n_27414));
	notech_inv i_31477(.A(n_17870), .Z(n_27415));
	notech_inv i_31478(.A(n_17876), .Z(n_27416));
	notech_inv i_31479(.A(n_17882), .Z(n_27417));
	notech_inv i_31480(.A(n_17888), .Z(n_27418));
	notech_inv i_31481(.A(n_17894), .Z(n_27419));
	notech_inv i_31482(.A(n_17906), .Z(n_27420));
	notech_inv i_31483(.A(n_22720), .Z(n_27421));
	notech_inv i_31484(.A(temp_sp[0]), .Z(n_27422));
	notech_inv i_31485(.A(n_22725), .Z(n_27423));
	notech_inv i_31486(.A(temp_sp[1]), .Z(n_27424));
	notech_inv i_31487(.A(n_22730), .Z(n_27425));
	notech_inv i_31488(.A(temp_sp[2]), .Z(n_27426));
	notech_inv i_31489(.A(n_22735), .Z(n_27427));
	notech_inv i_31490(.A(temp_sp[3]), .Z(n_27428));
	notech_inv i_31491(.A(n_22740), .Z(n_27429));
	notech_inv i_31492(.A(temp_sp[4]), .Z(n_27430));
	notech_inv i_31493(.A(n_22745), .Z(n_27431));
	notech_inv i_31494(.A(temp_sp[5]), .Z(n_27432));
	notech_inv i_31495(.A(n_22750), .Z(n_27433));
	notech_inv i_31496(.A(temp_sp[6]), .Z(n_27434));
	notech_inv i_31497(.A(n_22755), .Z(n_27435));
	notech_inv i_31498(.A(temp_sp[7]), .Z(n_27437));
	notech_inv i_31499(.A(n_22760), .Z(n_27438));
	notech_inv i_31500(.A(temp_sp[8]), .Z(n_27439));
	notech_inv i_31501(.A(n_22765), .Z(n_27440));
	notech_inv i_31502(.A(temp_sp[9]), .Z(n_27441));
	notech_inv i_31503(.A(n_22770), .Z(n_27442));
	notech_inv i_31504(.A(temp_sp[10]), .Z(n_27443));
	notech_inv i_31505(.A(n_22775), .Z(n_27444));
	notech_inv i_31506(.A(temp_sp[11]), .Z(n_27445));
	notech_inv i_31507(.A(n_22780), .Z(n_27446));
	notech_inv i_31508(.A(temp_sp[12]), .Z(n_27447));
	notech_inv i_31509(.A(n_22785), .Z(n_27448));
	notech_inv i_31510(.A(temp_sp[13]), .Z(n_27449));
	notech_inv i_31511(.A(n_22790), .Z(n_27450));
	notech_inv i_31512(.A(temp_sp[14]), .Z(n_27451));
	notech_inv i_31513(.A(n_22795), .Z(n_27452));
	notech_inv i_31514(.A(temp_sp[15]), .Z(n_27453));
	notech_inv i_31515(.A(n_22800), .Z(n_27454));
	notech_inv i_31516(.A(temp_sp[16]), .Z(n_27455));
	notech_inv i_31517(.A(n_22805), .Z(n_27456));
	notech_inv i_31518(.A(temp_sp[17]), .Z(n_27457));
	notech_inv i_31519(.A(n_22810), .Z(n_27458));
	notech_inv i_31520(.A(temp_sp[18]), .Z(n_27459));
	notech_inv i_31521(.A(n_22815), .Z(n_27460));
	notech_inv i_31522(.A(temp_sp[19]), .Z(n_27461));
	notech_inv i_31523(.A(n_22820), .Z(n_27462));
	notech_inv i_31524(.A(temp_sp[20]), .Z(n_27463));
	notech_inv i_31525(.A(n_22825), .Z(n_27464));
	notech_inv i_31526(.A(temp_sp[21]), .Z(n_27465));
	notech_inv i_31527(.A(n_22830), .Z(n_27466));
	notech_inv i_31528(.A(temp_sp[22]), .Z(n_27469));
	notech_inv i_31529(.A(n_22835), .Z(n_27470));
	notech_inv i_31530(.A(temp_sp[23]), .Z(n_27471));
	notech_inv i_31531(.A(n_22840), .Z(n_27472));
	notech_inv i_31532(.A(temp_sp[24]), .Z(n_27473));
	notech_inv i_31533(.A(n_22845), .Z(n_27474));
	notech_inv i_31534(.A(temp_sp[25]), .Z(n_27475));
	notech_inv i_31535(.A(n_22850), .Z(n_27476));
	notech_inv i_31536(.A(temp_sp[26]), .Z(n_27477));
	notech_inv i_31537(.A(n_22855), .Z(n_27478));
	notech_inv i_31538(.A(temp_sp[27]), .Z(n_27479));
	notech_inv i_31539(.A(n_22860), .Z(n_27480));
	notech_inv i_31540(.A(temp_sp[28]), .Z(n_27481));
	notech_inv i_31541(.A(n_22865), .Z(n_27482));
	notech_inv i_31542(.A(temp_sp[29]), .Z(n_27483));
	notech_inv i_31543(.A(n_22870), .Z(n_27484));
	notech_inv i_31544(.A(temp_sp[30]), .Z(n_27485));
	notech_inv i_31545(.A(n_22875), .Z(n_27486));
	notech_inv i_31546(.A(temp_sp[31]), .Z(n_27487));
	notech_inv i_31547(.A(n_20984), .Z(n_27488));
	notech_inv i_31548(.A(n_21050), .Z(n_27489));
	notech_inv i_31549(.A(n_21062), .Z(n_27490));
	notech_inv i_31550(.A(n_21068), .Z(n_27491));
	notech_inv i_31551(.A(n_20624), .Z(n_27492));
	notech_inv i_31552(.A(n_274591882), .Z(n_27493));
	notech_inv i_31553(.A(n_20630), .Z(n_27494));
	notech_inv i_31554(.A(n_20654), .Z(n_27495));
	notech_inv i_31555(.A(n_20660), .Z(n_27496));
	notech_inv i_31556(.A(n_20672), .Z(n_27497));
	notech_inv i_31557(.A(n_20690), .Z(n_27498));
	notech_inv i_31558(.A(n_20702), .Z(n_27499));
	notech_inv i_31559(.A(n_20708), .Z(n_27502));
	notech_inv i_31560(.A(n_20714), .Z(n_27503));
	notech_inv i_31561(.A(n_20750), .Z(n_27504));
	notech_inv i_31562(.A(n_20762), .Z(n_27506));
	notech_inv i_31563(.A(n_20774), .Z(n_27507));
	notech_inv i_31564(.A(n_20792), .Z(n_27508));
	notech_inv i_31565(.A(n_20798), .Z(n_27510));
	notech_inv i_31566(.A(n_20804), .Z(n_27511));
	notech_inv i_31567(.A(\nbus_14522[1] ), .Z(n_27512));
	notech_inv i_31568(.A(\nbus_14522[3] ), .Z(n_27513));
	notech_inv i_31569(.A(\nbus_14522[4] ), .Z(n_27514));
	notech_inv i_31570(.A(\nbus_14522[6] ), .Z(n_27515));
	notech_inv i_31571(.A(\nbus_14522[7] ), .Z(n_27516));
	notech_inv i_31572(.A(\nbus_14522[8] ), .Z(n_27517));
	notech_inv i_31573(.A(\nbus_14522[9] ), .Z(n_27518));
	notech_inv i_31574(.A(\nbus_14522[10] ), .Z(n_27519));
	notech_inv i_31575(.A(\nbus_14522[11] ), .Z(n_27520));
	notech_inv i_31576(.A(\nbus_14522[12] ), .Z(n_27521));
	notech_inv i_31577(.A(\nbus_14522[13] ), .Z(n_27522));
	notech_inv i_31578(.A(\nbus_14522[14] ), .Z(n_27523));
	notech_inv i_31579(.A(\nbus_14522[15] ), .Z(n_27524));
	notech_inv i_31580(.A(\nbus_14522[17] ), .Z(n_27525));
	notech_inv i_31581(.A(\nbus_14522[18] ), .Z(n_27526));
	notech_inv i_31582(.A(\nbus_14522[19] ), .Z(n_27527));
	notech_inv i_31583(.A(\nbus_14522[20] ), .Z(n_27528));
	notech_inv i_31584(.A(\nbus_14522[21] ), .Z(n_27529));
	notech_inv i_31585(.A(\nbus_14522[22] ), .Z(n_27530));
	notech_inv i_31586(.A(\nbus_14522[23] ), .Z(n_27531));
	notech_inv i_31587(.A(\nbus_14522[24] ), .Z(n_27532));
	notech_inv i_31588(.A(\nbus_14522[25] ), .Z(n_27533));
	notech_inv i_31589(.A(\nbus_14522[26] ), .Z(n_27534));
	notech_inv i_31590(.A(\nbus_14522[27] ), .Z(n_27536));
	notech_inv i_31591(.A(\nbus_14522[28] ), .Z(n_27537));
	notech_inv i_31592(.A(\nbus_14522[29] ), .Z(n_27538));
	notech_inv i_31593(.A(\nbus_14522[30] ), .Z(n_27539));
	notech_inv i_31594(.A(n_16489), .Z(n_27540));
	notech_inv i_31595(.A(mask8b[0]), .Z(n_27541));
	notech_inv i_31596(.A(n_16495), .Z(n_27542));
	notech_inv i_31597(.A(n_19154), .Z(n_27543));
	notech_inv i_31598(.A(n_19160), .Z(n_27544));
	notech_inv i_31599(.A(n_19166), .Z(n_27545));
	notech_inv i_31600(.A(n_19172), .Z(n_27546));
	notech_inv i_31601(.A(n_19178), .Z(n_27547));
	notech_inv i_31602(.A(n_19184), .Z(n_27548));
	notech_inv i_31603(.A(n_19190), .Z(n_27549));
	notech_inv i_31604(.A(\nbus_11337[16] ), .Z(n_27550));
	notech_inv i_31605(.A(n_17432), .Z(n_27551));
	notech_inv i_31606(.A(n_2492), .Z(n_27552));
	notech_inv i_31607(.A(n_17444), .Z(n_27553));
	notech_inv i_31608(.A(n_17468), .Z(n_27554));
	notech_inv i_31609(.A(n_17474), .Z(n_27555));
	notech_inv i_31610(.A(n_17492), .Z(n_27556));
	notech_inv i_31611(.A(n_17498), .Z(n_27557));
	notech_inv i_31612(.A(n_2487), .Z(n_27558));
	notech_inv i_31613(.A(n_17510), .Z(n_27559));
	notech_inv i_31614(.A(n_17516), .Z(n_27560));
	notech_inv i_31615(.A(n_17534), .Z(n_27561));
	notech_inv i_31616(.A(n_17546), .Z(n_27562));
	notech_inv i_31617(.A(n_2484), .Z(n_27563));
	notech_inv i_31618(.A(n_17552), .Z(n_27564));
	notech_inv i_31619(.A(n_17564), .Z(n_27565));
	notech_inv i_31620(.A(n_2483), .Z(n_27566));
	notech_inv i_31621(.A(n_17570), .Z(n_27567));
	notech_inv i_31622(.A(n_17576), .Z(n_27568));
	notech_inv i_31623(.A(n_17582), .Z(n_27569));
	notech_inv i_31624(.A(n_2482), .Z(n_27571));
	notech_inv i_31625(.A(n_2481), .Z(n_27572));
	notech_inv i_31626(.A(n_2478), .Z(n_27573));
	notech_inv i_31627(.A(n_17612), .Z(n_27574));
	notech_inv i_31629(.A(\nbus_11331[0] ), .Z(n_27575));
	notech_inv i_31630(.A(n_17075), .Z(n_27576));
	notech_inv i_31631(.A(n_59286), .Z(n_27577));
	notech_inv i_31632(.A(n_17195), .Z(n_27578));
	notech_inv i_31633(.A(n_17213), .Z(n_27579));
	notech_inv i_31634(.A(n_17219), .Z(n_27581));
	notech_inv i_31635(.A(n_17225), .Z(n_27582));
	notech_inv i_31636(.A(n_13536), .Z(n_27583));
	notech_inv i_31637(.A(n_13541), .Z(n_27584));
	notech_inv i_31638(.A(n_13546), .Z(n_27585));
	notech_inv i_31639(.A(n_13551), .Z(n_27586));
	notech_inv i_31640(.A(n_13556), .Z(n_27587));
	notech_inv i_31641(.A(n_13561), .Z(n_27588));
	notech_inv i_31642(.A(n_13566), .Z(n_27589));
	notech_inv i_31643(.A(n_13571), .Z(n_27590));
	notech_inv i_31644(.A(n_13576), .Z(n_27591));
	notech_inv i_31645(.A(n_13581), .Z(n_27592));
	notech_inv i_31646(.A(n_13586), .Z(n_27593));
	notech_inv i_31647(.A(n_13591), .Z(n_27594));
	notech_inv i_31648(.A(n_13596), .Z(n_27595));
	notech_inv i_31650(.A(n_13601), .Z(n_27596));
	notech_inv i_31651(.A(n_13606), .Z(n_27597));
	notech_inv i_31652(.A(n_13611), .Z(n_27598));
	notech_inv i_31653(.A(n_13616), .Z(n_27599));
	notech_inv i_31654(.A(n_13621), .Z(n_27600));
	notech_inv i_31655(.A(n_13626), .Z(n_27602));
	notech_inv i_31656(.A(n_13631), .Z(n_27603));
	notech_inv i_31657(.A(n_13636), .Z(n_27605));
	notech_inv i_31658(.A(n_13641), .Z(n_27606));
	notech_inv i_31659(.A(n_13646), .Z(n_27607));
	notech_inv i_31660(.A(n_13651), .Z(n_27608));
	notech_inv i_31661(.A(n_13656), .Z(n_27609));
	notech_inv i_31662(.A(n_13661), .Z(n_27610));
	notech_inv i_31663(.A(n_13666), .Z(n_27611));
	notech_inv i_31664(.A(n_13671), .Z(n_27613));
	notech_inv i_31665(.A(n_13676), .Z(n_27614));
	notech_inv i_31666(.A(n_13681), .Z(n_27615));
	notech_inv i_31669(.A(n_15021), .Z(n_27619));
	notech_inv i_31670(.A(n_15026), .Z(n_27620));
	notech_inv i_31671(.A(n_15036), .Z(n_27621));
	notech_inv i_31672(.A(\nbus_11313[0] ), .Z(n_27622));
	notech_inv i_31673(.A(\nbus_11313[5] ), .Z(n_27623));
	notech_inv i_31674(.A(n_15101), .Z(n_27624));
	notech_inv i_31676(.A(n_15106), .Z(n_27625));
	notech_inv i_31677(.A(n_15111), .Z(n_27626));
	notech_inv i_31678(.A(n_15116), .Z(n_27627));
	notech_inv i_31679(.A(n_15121), .Z(n_27628));
	notech_inv i_31680(.A(n_15126), .Z(n_27629));
	notech_inv i_31681(.A(n_15131), .Z(n_27630));
	notech_inv i_31682(.A(n_15136), .Z(n_27631));
	notech_inv i_31683(.A(n_15141), .Z(n_27632));
	notech_inv i_31684(.A(n_15146), .Z(n_27633));
	notech_inv i_31685(.A(n_15151), .Z(n_27634));
	notech_inv i_31686(.A(n_15156), .Z(n_27635));
	notech_inv i_31687(.A(n_15161), .Z(n_27636));
	notech_inv i_31688(.A(n_15166), .Z(n_27637));
	notech_inv i_31689(.A(n_15171), .Z(n_27638));
	notech_inv i_31690(.A(n_15176), .Z(n_27639));
	notech_inv i_31691(.A(\nbus_11313[16] ), .Z(n_27640));
	notech_inv i_31692(.A(nZF), .Z(n_27641));
	notech_inv i_31693(.A(n_16706), .Z(n_27642));
	notech_inv i_31694(.A(n_16718), .Z(n_27643));
	notech_inv i_31695(.A(n_16730), .Z(n_27644));
	notech_inv i_31696(.A(n_16748), .Z(n_27645));
	notech_inv i_31697(.A(n_16760), .Z(n_27646));
	notech_inv i_31698(.A(n_16766), .Z(n_27647));
	notech_inv i_31699(.A(n_16772), .Z(n_27648));
	notech_inv i_31700(.A(n_16790), .Z(n_27649));
	notech_inv i_31701(.A(n_16796), .Z(n_27650));
	notech_inv i_31702(.A(n_16880), .Z(n_27651));
	notech_inv i_31703(.A(\nbus_11329[0] ), .Z(n_27652));
	notech_inv i_31704(.A(nbus_14521[0]), .Z(n_27653));
	notech_inv i_31705(.A(nbus_14521[1]), .Z(n_27654));
	notech_inv i_31706(.A(nbus_14521[2]), .Z(n_27655));
	notech_inv i_31707(.A(nbus_14521[3]), .Z(n_27656));
	notech_inv i_31708(.A(nbus_14521[4]), .Z(n_27657));
	notech_inv i_31709(.A(nbus_14521[6]), .Z(n_27658));
	notech_inv i_31710(.A(nbus_14521[7]), .Z(n_27659));
	notech_inv i_31711(.A(nbus_14521[15]), .Z(n_27660));
	notech_inv i_31712(.A(nbus_14521[16]), .Z(n_27661));
	notech_inv i_31713(.A(nbus_14521[17]), .Z(n_27662));
	notech_inv i_31714(.A(nbus_14521[18]), .Z(n_27663));
	notech_inv i_31715(.A(nbus_14521[19]), .Z(n_27664));
	notech_inv i_31716(.A(nbus_14521[20]), .Z(n_27665));
	notech_inv i_31717(.A(nbus_14521[21]), .Z(n_27666));
	notech_inv i_31718(.A(nbus_14521[22]), .Z(n_27667));
	notech_inv i_31719(.A(nbus_14521[23]), .Z(n_27668));
	notech_inv i_31720(.A(nbus_14521[24]), .Z(n_27669));
	notech_inv i_31721(.A(nbus_14521[25]), .Z(n_27670));
	notech_inv i_31722(.A(nbus_14521[26]), .Z(n_27671));
	notech_inv i_31723(.A(nbus_14521[27]), .Z(n_27672));
	notech_inv i_31724(.A(nbus_14521[28]), .Z(n_27673));
	notech_inv i_31725(.A(nbus_14521[29]), .Z(n_27674));
	notech_inv i_31726(.A(nbus_14521[30]), .Z(n_27675));
	notech_inv i_31727(.A(cr2_reg[0]), .Z(n_27676));
	notech_inv i_31728(.A(cr2_reg[1]), .Z(n_27677));
	notech_inv i_31729(.A(cr2_reg[3]), .Z(n_27678));
	notech_inv i_31730(.A(cr2_reg[4]), .Z(n_27679));
	notech_inv i_31731(.A(cr2_reg[5]), .Z(n_27680));
	notech_inv i_31732(.A(cr2_reg[6]), .Z(n_27681));
	notech_inv i_31733(.A(cr2_reg[7]), .Z(n_27682));
	notech_inv i_31734(.A(cr2_reg[8]), .Z(n_27683));
	notech_inv i_31735(.A(cr2_reg[9]), .Z(n_27684));
	notech_inv i_31736(.A(cr2_reg[10]), .Z(n_27685));
	notech_inv i_31737(.A(cr2_reg[11]), .Z(n_27686));
	notech_inv i_31738(.A(cr2_reg[12]), .Z(n_27687));
	notech_inv i_31740(.A(cr2_reg[13]), .Z(n_27688));
	notech_inv i_31742(.A(cr2_reg[14]), .Z(n_27689));
	notech_inv i_31743(.A(cr2_reg[15]), .Z(n_27690));
	notech_inv i_31744(.A(cr2_reg[31]), .Z(n_27691));
	notech_inv i_31745(.A(\nbus_14520[0] ), .Z(n_27692));
	notech_inv i_31746(.A(\nbus_14520[1] ), .Z(n_27693));
	notech_inv i_31747(.A(\nbus_14520[2] ), .Z(n_27694));
	notech_inv i_31748(.A(\nbus_14520[6] ), .Z(n_27695));
	notech_inv i_31749(.A(\nbus_14520[8] ), .Z(n_27696));
	notech_inv i_31750(.A(\nbus_14520[9] ), .Z(n_27697));
	notech_inv i_31751(.A(\nbus_14520[10] ), .Z(n_27698));
	notech_inv i_31752(.A(\nbus_14520[11] ), .Z(n_27699));
	notech_inv i_31753(.A(n_22215), .Z(n_27700));
	notech_inv i_31754(.A(n_22221), .Z(n_27701));
	notech_inv i_31755(.A(\nbus_11356[0] ), .Z(n_27702));
	notech_inv i_31756(.A(n_22263), .Z(n_27703));
	notech_inv i_31757(.A(n_22269), .Z(n_27704));
	notech_inv i_31758(.A(n_22275), .Z(n_27705));
	notech_inv i_31759(.A(n_22281), .Z(n_27706));
	notech_inv i_31760(.A(n_22287), .Z(n_27707));
	notech_inv i_31762(.A(n_22293), .Z(n_27708));
	notech_inv i_31763(.A(n_22299), .Z(n_27709));
	notech_inv i_31764(.A(n_22305), .Z(n_27710));
	notech_inv i_31765(.A(\nbus_11356[8] ), .Z(n_27711));
	notech_inv i_31766(.A(n_2026), .Z(n_27712));
	notech_inv i_31767(.A(\nbus_11356[16] ), .Z(n_27713));
	notech_inv i_31768(.A(tcmp), .Z(n_27714));
	notech_inv i_31769(.A(n_1881), .Z(n_27715));
	notech_inv i_31770(.A(n_19653), .Z(n_27716));
	notech_inv i_31771(.A(fsm[1]), .Z(n_27717));
	notech_inv i_31772(.A(n_19659), .Z(n_27718));
	notech_inv i_31773(.A(n_61171), .Z(n_27719));
	notech_inv i_31774(.A(fsm[3]), .Z(n_27720));
	notech_inv i_31775(.A(n_19671), .Z(n_27721));
	notech_inv i_31776(.A(vliw_pc[0]), .Z(n_27722));
	notech_inv i_31777(.A(vliw_pc[1]), .Z(n_27723));
	notech_inv i_31778(.A(vliw_pc[2]), .Z(n_27724));
	notech_inv i_31779(.A(n_25953), .Z(n_27725));
	notech_inv i_31780(.A(n_25963), .Z(n_27726));
	notech_inv i_31781(.A(n_26103), .Z(n_27727));
	notech_inv i_31782(.A(temp_ss[0]), .Z(n_27728));
	notech_inv i_31783(.A(temp_ss[1]), .Z(n_27729));
	notech_inv i_31784(.A(temp_ss[2]), .Z(n_27730));
	notech_inv i_31785(.A(temp_ss[3]), .Z(n_27731));
	notech_inv i_31786(.A(temp_ss[4]), .Z(n_27732));
	notech_inv i_31787(.A(temp_ss[5]), .Z(n_27733));
	notech_inv i_31788(.A(temp_ss[6]), .Z(n_27734));
	notech_inv i_31789(.A(temp_ss[7]), .Z(n_27735));
	notech_inv i_31790(.A(temp_ss[8]), .Z(n_27737));
	notech_inv i_31791(.A(temp_ss[9]), .Z(n_27738));
	notech_inv i_31792(.A(temp_ss[10]), .Z(n_27739));
	notech_inv i_31793(.A(temp_ss[11]), .Z(n_27740));
	notech_inv i_31794(.A(temp_ss[12]), .Z(n_27741));
	notech_inv i_31795(.A(temp_ss[13]), .Z(n_27742));
	notech_inv i_31796(.A(temp_ss[14]), .Z(n_27743));
	notech_inv i_31797(.A(temp_ss[15]), .Z(n_27744));
	notech_inv i_31798(.A(temp_ss[16]), .Z(n_27745));
	notech_inv i_31799(.A(temp_ss[17]), .Z(n_27747));
	notech_inv i_31800(.A(temp_ss[18]), .Z(n_27748));
	notech_inv i_31801(.A(temp_ss[19]), .Z(n_27749));
	notech_inv i_31802(.A(temp_ss[20]), .Z(n_27750));
	notech_inv i_31803(.A(temp_ss[21]), .Z(n_27751));
	notech_inv i_31804(.A(temp_ss[22]), .Z(n_27752));
	notech_inv i_31805(.A(temp_ss[23]), .Z(n_27755));
	notech_inv i_31806(.A(temp_ss[24]), .Z(n_27756));
	notech_inv i_31807(.A(temp_ss[25]), .Z(n_27758));
	notech_inv i_31808(.A(temp_ss[26]), .Z(n_27759));
	notech_inv i_31809(.A(temp_ss[27]), .Z(n_27760));
	notech_inv i_31810(.A(temp_ss[28]), .Z(n_27762));
	notech_inv i_31811(.A(temp_ss[29]), .Z(n_27763));
	notech_inv i_31812(.A(temp_ss[30]), .Z(n_27764));
	notech_inv i_31813(.A(temp_ss[31]), .Z(n_27765));
	notech_inv i_31814(.A(errco[0]), .Z(n_27766));
	notech_inv i_31815(.A(errco[1]), .Z(n_27767));
	notech_inv i_31816(.A(errco[2]), .Z(n_27768));
	notech_inv i_31817(.A(errco[3]), .Z(n_27769));
	notech_inv i_31818(.A(errco[4]), .Z(n_27770));
	notech_inv i_31819(.A(errco[5]), .Z(n_27771));
	notech_inv i_31820(.A(n_1826), .Z(n_27772));
	notech_inv i_31821(.A(errco[6]), .Z(n_27773));
	notech_inv i_31822(.A(errco[7]), .Z(n_27774));
	notech_inv i_31823(.A(errco[8]), .Z(n_27775));
	notech_inv i_31824(.A(errco[9]), .Z(n_27776));
	notech_inv i_31825(.A(errco[10]), .Z(n_27777));
	notech_inv i_31826(.A(errco[11]), .Z(n_27779));
	notech_inv i_31827(.A(errco[12]), .Z(n_27780));
	notech_inv i_31828(.A(errco[13]), .Z(n_27783));
	notech_inv i_31829(.A(errco[14]), .Z(n_27785));
	notech_inv i_31830(.A(errco[15]), .Z(n_27786));
	notech_inv i_31831(.A(errco[16]), .Z(n_27787));
	notech_inv i_31832(.A(errco[17]), .Z(n_27788));
	notech_inv i_31833(.A(errco[18]), .Z(n_27789));
	notech_inv i_31834(.A(errco[19]), .Z(n_27790));
	notech_inv i_31835(.A(errco[20]), .Z(n_27791));
	notech_inv i_31836(.A(errco[21]), .Z(n_27792));
	notech_inv i_31837(.A(errco[22]), .Z(n_27793));
	notech_inv i_31838(.A(errco[23]), .Z(n_27794));
	notech_inv i_31839(.A(errco[24]), .Z(n_27795));
	notech_inv i_31840(.A(n_1817), .Z(n_27796));
	notech_inv i_31841(.A(errco[25]), .Z(n_27797));
	notech_inv i_31842(.A(errco[26]), .Z(n_27798));
	notech_inv i_31843(.A(errco[27]), .Z(n_27799));
	notech_inv i_31844(.A(errco[28]), .Z(n_27800));
	notech_inv i_31845(.A(errco[29]), .Z(n_27801));
	notech_inv i_31846(.A(errco[30]), .Z(n_27802));
	notech_inv i_31847(.A(errco[31]), .Z(n_27803));
	notech_inv i_31848(.A(Daddrgs[0]), .Z(n_27804));
	notech_inv i_31849(.A(Daddrgs[2]), .Z(n_27805));
	notech_inv i_31850(.A(Daddrgs[3]), .Z(n_27806));
	notech_inv i_31851(.A(Daddrgs[4]), .Z(n_27807));
	notech_inv i_31852(.A(Daddrgs[5]), .Z(n_27808));
	notech_inv i_31853(.A(Daddrgs[6]), .Z(n_27809));
	notech_inv i_31854(.A(Daddrgs[7]), .Z(n_27810));
	notech_inv i_31855(.A(Daddrgs[8]), .Z(n_27811));
	notech_inv i_31857(.A(Daddrgs[9]), .Z(n_27812));
	notech_inv i_31858(.A(Daddrgs[10]), .Z(n_27813));
	notech_inv i_31859(.A(Daddrgs[11]), .Z(n_27814));
	notech_inv i_31860(.A(Daddrgs[12]), .Z(n_27815));
	notech_inv i_31861(.A(Daddrgs[13]), .Z(n_27816));
	notech_inv i_31862(.A(Daddrgs[14]), .Z(n_27817));
	notech_inv i_31863(.A(Daddrgs[15]), .Z(n_27818));
	notech_inv i_31864(.A(Daddrgs[16]), .Z(n_27819));
	notech_inv i_31865(.A(Daddrgs[17]), .Z(n_27820));
	notech_inv i_31867(.A(Daddrgs[18]), .Z(n_27821));
	notech_inv i_31868(.A(Daddrgs[19]), .Z(n_27822));
	notech_inv i_31869(.A(Daddrgs[20]), .Z(n_27823));
	notech_inv i_31870(.A(Daddrgs[21]), .Z(n_27824));
	notech_inv i_31871(.A(Daddrgs[22]), .Z(n_27825));
	notech_inv i_31872(.A(Daddrgs[23]), .Z(n_27826));
	notech_inv i_31873(.A(Daddrgs[24]), .Z(n_27827));
	notech_inv i_31874(.A(Daddrgs[25]), .Z(n_27828));
	notech_inv i_31875(.A(Daddrgs[26]), .Z(n_27829));
	notech_inv i_31876(.A(Daddrgs[27]), .Z(n_27830));
	notech_inv i_31877(.A(Daddrgs[28]), .Z(n_27831));
	notech_inv i_31878(.A(Daddrgs[29]), .Z(n_27832));
	notech_inv i_31879(.A(Daddrgs[30]), .Z(n_27833));
	notech_inv i_31880(.A(Daddrgs[31]), .Z(n_27834));
	notech_inv i_31881(.A(n_25488), .Z(n_27835));
	notech_inv i_31882(.A(n_25494), .Z(n_27836));
	notech_inv i_31883(.A(n_25500), .Z(n_27837));
	notech_inv i_31884(.A(n_25506), .Z(n_27838));
	notech_inv i_31885(.A(n_25512), .Z(n_27839));
	notech_inv i_31886(.A(n_25518), .Z(n_27840));
	notech_inv i_31887(.A(n_25524), .Z(n_27841));
	notech_inv i_31888(.A(n_25530), .Z(n_27842));
	notech_inv i_31889(.A(n_25536), .Z(n_27843));
	notech_inv i_31890(.A(n_25542), .Z(n_27844));
	notech_inv i_31891(.A(n_22451), .Z(n_27845));
	notech_inv i_31892(.A(\nbus_11357[0] ), .Z(n_27846));
	notech_inv i_31893(.A(\nbus_14522[31] ), .Z(n_27847));
	notech_inv i_31895(.A(cs[0]), .Z(n_27849));
	notech_inv i_31897(.A(cs[1]), .Z(n_27851));
	notech_inv i_31898(.A(all_cnt[0]), .Z(n_27852));
	notech_inv i_31900(.A(all_cnt[1]), .Z(n_27853));
	notech_inv i_31901(.A(all_cnt[2]), .Z(n_27854));
	notech_inv i_31903(.A(all_cnt[3]), .Z(n_27856));
	notech_inv i_31905(.A(ecx[0]), .Z(n_27858));
	notech_inv i_31906(.A(ecx[1]), .Z(n_27859));
	notech_inv i_31907(.A(ecx[2]), .Z(n_27860));
	notech_inv i_31908(.A(ecx[3]), .Z(n_27861));
	notech_inv i_31909(.A(ecx[4]), .Z(n_27862));
	notech_inv i_31910(.A(ecx[5]), .Z(n_27863));
	notech_inv i_31911(.A(ecx[6]), .Z(n_27864));
	notech_inv i_31912(.A(ecx[7]), .Z(n_27865));
	notech_inv i_31913(.A(ecx[8]), .Z(n_27866));
	notech_inv i_31914(.A(ecx[9]), .Z(n_27867));
	notech_inv i_31915(.A(ecx[10]), .Z(n_27868));
	notech_inv i_31916(.A(ecx[11]), .Z(n_27869));
	notech_inv i_31917(.A(ecx[12]), .Z(n_27870));
	notech_inv i_31918(.A(ecx[13]), .Z(n_27871));
	notech_inv i_31919(.A(ecx[14]), .Z(n_27872));
	notech_inv i_31920(.A(ecx[15]), .Z(n_27873));
	notech_inv i_31921(.A(ecx[16]), .Z(n_27874));
	notech_inv i_31922(.A(ecx[17]), .Z(n_27875));
	notech_inv i_31923(.A(ecx[18]), .Z(n_27876));
	notech_inv i_31924(.A(ecx[19]), .Z(n_27878));
	notech_inv i_31925(.A(ecx[20]), .Z(n_27881));
	notech_inv i_31926(.A(ecx[21]), .Z(n_27882));
	notech_inv i_31927(.A(ecx[22]), .Z(n_27883));
	notech_inv i_31928(.A(ecx[23]), .Z(n_27884));
	notech_inv i_31929(.A(ecx[24]), .Z(n_27886));
	notech_inv i_31930(.A(ecx[25]), .Z(n_27887));
	notech_inv i_31931(.A(ecx[26]), .Z(n_27888));
	notech_inv i_31932(.A(ecx[27]), .Z(n_27889));
	notech_inv i_31933(.A(ecx[28]), .Z(n_27890));
	notech_inv i_31934(.A(ecx[29]), .Z(n_27891));
	notech_inv i_31935(.A(ecx[30]), .Z(n_27892));
	notech_inv i_31936(.A(ecx[31]), .Z(n_27893));
	notech_inv i_31937(.A(calc_sz[0]), .Z(n_27894));
	notech_inv i_31938(.A(calc_sz[2]), .Z(n_27895));
	notech_inv i_31939(.A(nbus_11310[0]), .Z(n_27897));
	notech_inv i_31940(.A(nbus_11310[1]), .Z(n_27898));
	notech_inv i_31941(.A(nbus_11310[2]), .Z(n_27899));
	notech_inv i_31942(.A(nbus_11310[3]), .Z(n_27901));
	notech_inv i_31943(.A(nbus_11310[4]), .Z(n_27902));
	notech_inv i_31944(.A(nbus_11310[5]), .Z(n_27905));
	notech_inv i_31945(.A(nbus_11310[6]), .Z(n_27909));
	notech_inv i_31946(.A(nbus_11310[7]), .Z(n_27910));
	notech_inv i_31947(.A(nbus_11310[8]), .Z(n_27911));
	notech_inv i_31948(.A(nbus_11310[9]), .Z(n_27912));
	notech_inv i_31949(.A(nbus_11310[10]), .Z(n_27913));
	notech_inv i_31950(.A(nbus_11310[11]), .Z(n_27914));
	notech_inv i_31951(.A(nbus_11310[12]), .Z(n_27915));
	notech_inv i_31952(.A(nbus_11310[13]), .Z(n_27916));
	notech_inv i_31953(.A(nbus_11310[14]), .Z(n_27918));
	notech_inv i_31954(.A(nbus_11310[15]), .Z(n_27923));
	notech_inv i_31955(.A(nbus_11310[16]), .Z(n_27926));
	notech_inv i_31956(.A(nbus_11310[17]), .Z(n_27927));
	notech_inv i_31957(.A(nbus_11310[18]), .Z(n_27928));
	notech_inv i_31958(.A(nbus_11310[19]), .Z(n_27929));
	notech_inv i_31959(.A(nbus_11310[20]), .Z(n_27930));
	notech_inv i_31960(.A(nbus_11310[21]), .Z(n_27931));
	notech_inv i_31961(.A(nbus_11310[22]), .Z(n_27932));
	notech_inv i_31962(.A(nbus_11310[23]), .Z(n_27933));
	notech_inv i_31963(.A(nbus_11310[24]), .Z(n_27934));
	notech_inv i_31964(.A(nbus_11310[25]), .Z(n_27935));
	notech_inv i_31965(.A(nbus_11310[26]), .Z(n_27936));
	notech_inv i_31966(.A(nbus_11310[27]), .Z(n_27937));
	notech_inv i_31967(.A(nbus_11310[28]), .Z(n_27938));
	notech_inv i_31968(.A(nbus_11310[29]), .Z(n_27939));
	notech_inv i_31969(.A(nbus_11310[30]), .Z(n_27940));
	notech_inv i_31970(.A(nbus_11310[31]), .Z(n_27941));
	notech_inv i_31971(.A(n_60072), .Z(\nbus_11307[0] ));
	notech_inv i_31972(.A(opa[1]), .Z(\nbus_11307[1] ));
	notech_inv i_31974(.A(opa[3]), .Z(\nbus_11307[3] ));
	notech_inv i_31975(.A(opa[4]), .Z(\nbus_11307[4] ));
	notech_inv i_31976(.A(opa[5]), .Z(\nbus_11307[5] ));
	notech_inv i_31977(.A(n_60082), .Z(\nbus_11307[6] ));
	notech_inv i_31978(.A(n_60091), .Z(\nbus_11307[7] ));
	notech_inv i_31979(.A(opa[8]), .Z(\nbus_11307[8] ));
	notech_inv i_31983(.A(opa[9]), .Z(\nbus_11307[9] ));
	notech_inv i_31984(.A(opa[10]), .Z(\nbus_11307[10] ));
	notech_inv i_31985(.A(opa[11]), .Z(\nbus_11307[11] ));
	notech_inv i_31986(.A(opa[12]), .Z(\nbus_11307[12] ));
	notech_inv i_31987(.A(opa[13]), .Z(\nbus_11307[13] ));
	notech_inv i_31988(.A(opa[14]), .Z(\nbus_11307[14] ));
	notech_inv i_31989(.A(n_60102), .Z(\nbus_11307[15] ));
	notech_inv i_31990(.A(opa[16]), .Z(\nbus_11365[16] ));
	notech_inv i_31991(.A(opa[17]), .Z(\nbus_11365[17] ));
	notech_inv i_31992(.A(opa[18]), .Z(\nbus_11365[18] ));
	notech_inv i_31994(.A(opa[19]), .Z(\nbus_11365[19] ));
	notech_inv i_31995(.A(opa[20]), .Z(\nbus_11365[20] ));
	notech_inv i_31996(.A(opa[21]), .Z(\nbus_11365[21] ));
	notech_inv i_31997(.A(opa[22]), .Z(\nbus_11365[22] ));
	notech_inv i_31999(.A(opa[23]), .Z(\nbus_11365[23] ));
	notech_inv i_32000(.A(opa[24]), .Z(\nbus_11365[24] ));
	notech_inv i_32001(.A(opa[25]), .Z(\nbus_11365[25] ));
	notech_inv i_32002(.A(opa[26]), .Z(\nbus_11365[26] ));
	notech_inv i_32003(.A(opa[27]), .Z(\nbus_11365[27] ));
	notech_inv i_32004(.A(opa[28]), .Z(\nbus_11365[28] ));
	notech_inv i_32006(.A(opa[29]), .Z(\nbus_11365[29] ));
	notech_inv i_32007(.A(opa[30]), .Z(\nbus_11365[30] ));
	notech_inv i_32008(.A(opa[31]), .Z(\nbus_11365[31] ));
	notech_inv i_32009(.A(reps[2]), .Z(n_27980));
	notech_inv i_32011(.A(opd[0]), .Z(n_27981));
	notech_inv i_32012(.A(opd[1]), .Z(n_27983));
	notech_inv i_32014(.A(opd[2]), .Z(n_27984));
	notech_inv i_32015(.A(opd[3]), .Z(n_27985));
	notech_inv i_32016(.A(opd[4]), .Z(n_27986));
	notech_inv i_32017(.A(opd[5]), .Z(n_27987));
	notech_inv i_32018(.A(opd[6]), .Z(n_27989));
	notech_inv i_32019(.A(opd[7]), .Z(n_27990));
	notech_inv i_32020(.A(opd[8]), .Z(n_27991));
	notech_inv i_32021(.A(opd[9]), .Z(n_27992));
	notech_inv i_32023(.A(opd[10]), .Z(n_27993));
	notech_inv i_32024(.A(opd[11]), .Z(n_27996));
	notech_inv i_32025(.A(opd[12]), .Z(n_27997));
	notech_inv i_32026(.A(opd[13]), .Z(n_27998));
	notech_inv i_32027(.A(opd[14]), .Z(n_27999));
	notech_inv i_32028(.A(opd[15]), .Z(n_28000));
	notech_inv i_32029(.A(opd[16]), .Z(n_28001));
	notech_inv i_32030(.A(opd[17]), .Z(n_28002));
	notech_inv i_32031(.A(opd[18]), .Z(n_28003));
	notech_inv i_32032(.A(opd[19]), .Z(n_28004));
	notech_inv i_32033(.A(opd[20]), .Z(n_28005));
	notech_inv i_32034(.A(opd[21]), .Z(n_28006));
	notech_inv i_32035(.A(opd[22]), .Z(n_28007));
	notech_inv i_32036(.A(opd[23]), .Z(n_28008));
	notech_inv i_32037(.A(opd[24]), .Z(n_28009));
	notech_inv i_32038(.A(opd[25]), .Z(n_28010));
	notech_inv i_32039(.A(opd[26]), .Z(n_28011));
	notech_inv i_32040(.A(opd[27]), .Z(n_28012));
	notech_inv i_32041(.A(opd[28]), .Z(n_28013));
	notech_inv i_32042(.A(opd[29]), .Z(n_28014));
	notech_inv i_32043(.A(opd[30]), .Z(n_28015));
	notech_inv i_32044(.A(opd[31]), .Z(n_28016));
	notech_inv i_32045(.A(opb[0]), .Z(\nbus_11358[0] ));
	notech_inv i_32046(.A(opb[1]), .Z(\nbus_11358[1] ));
	notech_inv i_32047(.A(opb[2]), .Z(\nbus_11358[2] ));
	notech_inv i_32048(.A(opb[3]), .Z(\nbus_11358[3] ));
	notech_inv i_32049(.A(opb[4]), .Z(\nbus_11358[4] ));
	notech_inv i_32050(.A(opb[5]), .Z(\nbus_11358[5] ));
	notech_inv i_32051(.A(opb[6]), .Z(\nbus_11358[6] ));
	notech_inv i_32052(.A(opb[7]), .Z(\nbus_11358[7] ));
	notech_inv i_32057(.A(opb[8]), .Z(\nbus_11358[8] ));
	notech_inv i_32058(.A(opb[9]), .Z(\nbus_11358[9] ));
	notech_inv i_32059(.A(opb[10]), .Z(\nbus_11358[10] ));
	notech_inv i_32060(.A(opb[11]), .Z(\nbus_11358[11] ));
	notech_inv i_32061(.A(opb[12]), .Z(\nbus_11358[12] ));
	notech_inv i_32062(.A(opb[13]), .Z(\nbus_11358[13] ));
	notech_inv i_32063(.A(opb[14]), .Z(\nbus_11358[14] ));
	notech_inv i_32064(.A(opb[15]), .Z(\nbus_11358[15] ));
	notech_inv i_32065(.A(opb[16]), .Z(\nbus_11358[16] ));
	notech_inv i_32066(.A(opb[17]), .Z(\nbus_11358[17] ));
	notech_inv i_32067(.A(opb[18]), .Z(\nbus_11358[18] ));
	notech_inv i_32068(.A(opb[19]), .Z(\nbus_11358[19] ));
	notech_inv i_32069(.A(opb[20]), .Z(\nbus_11358[20] ));
	notech_inv i_32070(.A(opb[21]), .Z(\nbus_11358[21] ));
	notech_inv i_32072(.A(opb[22]), .Z(\nbus_11358[22] ));
	notech_inv i_32073(.A(opb[23]), .Z(\nbus_11358[23] ));
	notech_inv i_32074(.A(opb[24]), .Z(\nbus_11358[24] ));
	notech_inv i_32076(.A(opb[25]), .Z(\nbus_11358[25] ));
	notech_inv i_32077(.A(opb[26]), .Z(\nbus_11358[26] ));
	notech_inv i_32078(.A(opb[27]), .Z(\nbus_11358[27] ));
	notech_inv i_32079(.A(opb[28]), .Z(\nbus_11358[28] ));
	notech_inv i_32080(.A(opb[29]), .Z(\nbus_11358[29] ));
	notech_inv i_32081(.A(opb[30]), .Z(\nbus_11358[30] ));
	notech_inv i_32082(.A(opb[31]), .Z(\nbus_11358[31] ));
	notech_inv i_32083(.A(opz[0]), .Z(n_28049));
	notech_inv i_32084(.A(opz[1]), .Z(n_28050));
	notech_inv i_32085(.A(opz[2]), .Z(n_28051));
	notech_inv i_32086(.A(opc[0]), .Z(nbus_11295[0]));
	notech_inv i_32087(.A(opc[1]), .Z(nbus_11295[1]));
	notech_inv i_32088(.A(opc[2]), .Z(nbus_11295[2]));
	notech_inv i_32089(.A(opc[3]), .Z(nbus_11295[3]));
	notech_inv i_32090(.A(opc[4]), .Z(nbus_11295[4]));
	notech_inv i_32091(.A(opc[5]), .Z(nbus_11295[5]));
	notech_inv i_32092(.A(opc[6]), .Z(nbus_11295[6]));
	notech_inv i_32093(.A(opc[7]), .Z(nbus_11295[7]));
	notech_inv i_32094(.A(opc[8]), .Z(nbus_11295[8]));
	notech_inv i_32095(.A(opc[9]), .Z(nbus_11295[9]));
	notech_inv i_32096(.A(opc[10]), .Z(nbus_11295[10]));
	notech_inv i_32097(.A(opc[11]), .Z(nbus_11295[11]));
	notech_inv i_32098(.A(opc[12]), .Z(nbus_11295[12]));
	notech_inv i_32099(.A(opc[13]), .Z(nbus_11295[13]));
	notech_inv i_32100(.A(opc[14]), .Z(nbus_11295[14]));
	notech_inv i_32101(.A(opc[15]), .Z(nbus_11295[15]));
	notech_inv i_32102(.A(opc[16]), .Z(nbus_11295[16]));
	notech_inv i_32103(.A(opc[17]), .Z(nbus_11295[17]));
	notech_inv i_32104(.A(opc[18]), .Z(nbus_11295[18]));
	notech_inv i_32105(.A(opc[19]), .Z(nbus_11295[19]));
	notech_inv i_32106(.A(opc[20]), .Z(nbus_11295[20]));
	notech_inv i_32107(.A(opc[21]), .Z(nbus_11295[21]));
	notech_inv i_32108(.A(opc[22]), .Z(nbus_11295[22]));
	notech_inv i_32109(.A(opc[23]), .Z(nbus_11295[23]));
	notech_inv i_32110(.A(opc[24]), .Z(nbus_11295[24]));
	notech_inv i_32111(.A(opc[25]), .Z(nbus_11295[25]));
	notech_inv i_32112(.A(opc[26]), .Z(nbus_11295[26]));
	notech_inv i_32113(.A(opc[27]), .Z(nbus_11295[27]));
	notech_inv i_32114(.A(opc[28]), .Z(nbus_11295[28]));
	notech_inv i_32115(.A(opc[29]), .Z(nbus_11295[29]));
	notech_inv i_32116(.A(opc[30]), .Z(nbus_11295[30]));
	notech_inv i_32117(.A(opc[31]), .Z(nbus_11295[31]));
	notech_inv i_32118(.A(read_data[0]), .Z(n_28089));
	notech_inv i_32121(.A(read_data[1]), .Z(n_28090));
	notech_inv i_32122(.A(read_data[2]), .Z(n_28091));
	notech_inv i_32123(.A(read_data[3]), .Z(n_28092));
	notech_inv i_32124(.A(read_data[4]), .Z(n_28093));
	notech_inv i_32126(.A(read_data[5]), .Z(n_28094));
	notech_inv i_32127(.A(read_data[6]), .Z(n_28095));
	notech_inv i_32128(.A(read_data[7]), .Z(n_28096));
	notech_inv i_32129(.A(read_data[8]), .Z(n_28097));
	notech_inv i_32130(.A(read_data[9]), .Z(n_28098));
	notech_inv i_32131(.A(read_data[10]), .Z(n_28099));
	notech_inv i_32132(.A(read_data[11]), .Z(n_28100));
	notech_inv i_32133(.A(read_data[12]), .Z(n_28101));
	notech_inv i_32134(.A(read_data[13]), .Z(n_28102));
	notech_inv i_32135(.A(read_data[14]), .Z(n_28103));
	notech_inv i_32136(.A(read_data[15]), .Z(n_28104));
	notech_inv i_32137(.A(read_data[16]), .Z(n_28105));
	notech_inv i_32138(.A(read_data[17]), .Z(n_28106));
	notech_inv i_32139(.A(read_data[18]), .Z(n_28107));
	notech_inv i_32140(.A(read_data[19]), .Z(n_28108));
	notech_inv i_32141(.A(read_data[20]), .Z(n_28109));
	notech_inv i_32142(.A(read_data[21]), .Z(n_28110));
	notech_inv i_32143(.A(read_data[22]), .Z(n_28111));
	notech_inv i_32144(.A(read_data[23]), .Z(n_28112));
	notech_inv i_32145(.A(read_data[24]), .Z(n_28113));
	notech_inv i_32146(.A(read_data[25]), .Z(n_28114));
	notech_inv i_32147(.A(read_data[26]), .Z(n_28115));
	notech_inv i_32148(.A(read_data[27]), .Z(n_28116));
	notech_inv i_32149(.A(read_data[28]), .Z(n_28117));
	notech_inv i_32150(.A(read_data[29]), .Z(n_28118));
	notech_inv i_32151(.A(read_data[30]), .Z(n_28121));
	notech_inv i_32152(.A(read_data[31]), .Z(n_28123));
	notech_inv i_32153(.A(opc_10[0]), .Z(n_28124));
	notech_inv i_32154(.A(opc_10[1]), .Z(n_28125));
	notech_inv i_32155(.A(opc_10[2]), .Z(n_28126));
	notech_inv i_32156(.A(opc_10[3]), .Z(n_28127));
	notech_inv i_32157(.A(opc_10[4]), .Z(n_28128));
	notech_inv i_32158(.A(opc_10[5]), .Z(n_28129));
	notech_inv i_32159(.A(opc_10[6]), .Z(n_28131));
	notech_inv i_32160(.A(opc_10[7]), .Z(n_28133));
	notech_inv i_32161(.A(opc_10[8]), .Z(n_28134));
	notech_inv i_32162(.A(opc_10[9]), .Z(n_28135));
	notech_inv i_32163(.A(opc_10[10]), .Z(n_28136));
	notech_inv i_32164(.A(opc_10[11]), .Z(n_28137));
	notech_inv i_32165(.A(opc_10[12]), .Z(n_28138));
	notech_inv i_32166(.A(opc_10[13]), .Z(n_28139));
	notech_inv i_32167(.A(opc_10[14]), .Z(n_28140));
	notech_inv i_32168(.A(opc_10[15]), .Z(n_28141));
	notech_inv i_32169(.A(opc_10[16]), .Z(n_28142));
	notech_inv i_32170(.A(opc_10[17]), .Z(n_28143));
	notech_inv i_32171(.A(opc_10[18]), .Z(n_28144));
	notech_inv i_32172(.A(opc_10[19]), .Z(n_28145));
	notech_inv i_32173(.A(opc_10[20]), .Z(n_28146));
	notech_inv i_32174(.A(opc_10[21]), .Z(n_28147));
	notech_inv i_32175(.A(opc_10[22]), .Z(n_28148));
	notech_inv i_32176(.A(opc_10[23]), .Z(n_28149));
	notech_inv i_32177(.A(opc_10[24]), .Z(n_28150));
	notech_inv i_32178(.A(opc_10[25]), .Z(n_28151));
	notech_inv i_32179(.A(opc_10[26]), .Z(n_28152));
	notech_inv i_32180(.A(opc_10[27]), .Z(n_28153));
	notech_inv i_32181(.A(opc_10[28]), .Z(n_28154));
	notech_inv i_32182(.A(opc_10[29]), .Z(n_28155));
	notech_inv i_32183(.A(opc_10[30]), .Z(n_28156));
	notech_inv i_32184(.A(opc_10[31]), .Z(n_28157));
	notech_inv i_32185(.A(regs_14[0]), .Z(n_28158));
	notech_inv i_32186(.A(regs_14[1]), .Z(n_28159));
	notech_inv i_32187(.A(regs_14[2]), .Z(n_28160));
	notech_inv i_32188(.A(regs_14[3]), .Z(n_28161));
	notech_inv i_32189(.A(regs_14[4]), .Z(n_28162));
	notech_inv i_32190(.A(regs_14[5]), .Z(n_28163));
	notech_inv i_32191(.A(regs_14[6]), .Z(n_28164));
	notech_inv i_32192(.A(regs_14[7]), .Z(n_28165));
	notech_inv i_32193(.A(regs_14[8]), .Z(n_28166));
	notech_inv i_32195(.A(regs_14[9]), .Z(n_28167));
	notech_inv i_32196(.A(regs_14[10]), .Z(n_28168));
	notech_inv i_32197(.A(regs_14[11]), .Z(n_28169));
	notech_inv i_32198(.A(regs_14[12]), .Z(n_28170));
	notech_inv i_32199(.A(regs_14[13]), .Z(n_28171));
	notech_inv i_32200(.A(regs_14[14]), .Z(n_28172));
	notech_inv i_32201(.A(regs_14[15]), .Z(n_28173));
	notech_inv i_32202(.A(regs_14[16]), .Z(n_28174));
	notech_inv i_32203(.A(regs_14[17]), .Z(n_28175));
	notech_inv i_32204(.A(regs_14[18]), .Z(n_28176));
	notech_inv i_32205(.A(regs_14[19]), .Z(n_28177));
	notech_inv i_32206(.A(regs_14[20]), .Z(n_28178));
	notech_inv i_32207(.A(regs_14[21]), .Z(n_28179));
	notech_inv i_32208(.A(regs_14[22]), .Z(n_28180));
	notech_inv i_32209(.A(regs_14[23]), .Z(n_28181));
	notech_inv i_32210(.A(regs_14[24]), .Z(n_28182));
	notech_inv i_32211(.A(regs_14[25]), .Z(n_28183));
	notech_inv i_32212(.A(regs_14[26]), .Z(n_28184));
	notech_inv i_32213(.A(regs_14[27]), .Z(n_28185));
	notech_inv i_32214(.A(regs_14[28]), .Z(n_28186));
	notech_inv i_32215(.A(regs_14[29]), .Z(n_28187));
	notech_inv i_32216(.A(regs_14[30]), .Z(n_28188));
	notech_inv i_32217(.A(regs_14[31]), .Z(n_28189));
	notech_inv i_32218(.A(regs_11[0]), .Z(n_28190));
	notech_inv i_32219(.A(regs_11[1]), .Z(n_28191));
	notech_inv i_32220(.A(regs_11[2]), .Z(n_28192));
	notech_inv i_32221(.A(regs_11[3]), .Z(n_28193));
	notech_inv i_32222(.A(regs_11[4]), .Z(n_28194));
	notech_inv i_32223(.A(regs_11[5]), .Z(n_28195));
	notech_inv i_32224(.A(regs_11[6]), .Z(n_28196));
	notech_inv i_32225(.A(regs_11[7]), .Z(n_28197));
	notech_inv i_32226(.A(regs_11[8]), .Z(n_28198));
	notech_inv i_32227(.A(regs_11[9]), .Z(n_28199));
	notech_inv i_32228(.A(regs_11[10]), .Z(n_28200));
	notech_inv i_32229(.A(regs_11[11]), .Z(n_28201));
	notech_inv i_32230(.A(regs_11[12]), .Z(n_28202));
	notech_inv i_32231(.A(regs_11[13]), .Z(n_28203));
	notech_inv i_32232(.A(regs_11[14]), .Z(n_28204));
	notech_inv i_32234(.A(regs_11[15]), .Z(n_28205));
	notech_inv i_32235(.A(regs_11[16]), .Z(n_28206));
	notech_inv i_32236(.A(regs_11[17]), .Z(n_28207));
	notech_inv i_32237(.A(regs_11[18]), .Z(n_28208));
	notech_inv i_32238(.A(regs_11[19]), .Z(n_28209));
	notech_inv i_32240(.A(regs_11[20]), .Z(n_28210));
	notech_inv i_32241(.A(regs_11[21]), .Z(n_28211));
	notech_inv i_32242(.A(regs_11[22]), .Z(n_28212));
	notech_inv i_32243(.A(regs_11[23]), .Z(n_28213));
	notech_inv i_32244(.A(regs_11[24]), .Z(n_28214));
	notech_inv i_32245(.A(regs_11[25]), .Z(n_28215));
	notech_inv i_32246(.A(regs_11[26]), .Z(n_28216));
	notech_inv i_32247(.A(regs_11[27]), .Z(n_28217));
	notech_inv i_32248(.A(regs_11[28]), .Z(n_28218));
	notech_inv i_32249(.A(regs_11[29]), .Z(n_28219));
	notech_inv i_32250(.A(regs_11[30]), .Z(n_28220));
	notech_inv i_32251(.A(regs_11[31]), .Z(n_28221));
	notech_inv i_32252(.A(regs_12[0]), .Z(n_28223));
	notech_inv i_32253(.A(regs_12[1]), .Z(n_28224));
	notech_inv i_32254(.A(regs_12[2]), .Z(n_28225));
	notech_inv i_32255(.A(regs_12[3]), .Z(n_28226));
	notech_inv i_32256(.A(regs_12[4]), .Z(n_28227));
	notech_inv i_32257(.A(regs_12[5]), .Z(n_28228));
	notech_inv i_32258(.A(regs_12[6]), .Z(n_28229));
	notech_inv i_32259(.A(regs_12[7]), .Z(n_28230));
	notech_inv i_32260(.A(regs_12[8]), .Z(n_28231));
	notech_inv i_32261(.A(regs_12[9]), .Z(n_28232));
	notech_inv i_32262(.A(regs_12[10]), .Z(n_28233));
	notech_inv i_32263(.A(regs_12[11]), .Z(n_28235));
	notech_inv i_32264(.A(regs_12[12]), .Z(n_28237));
	notech_inv i_32265(.A(regs_12[13]), .Z(n_28238));
	notech_inv i_32266(.A(regs_12[14]), .Z(n_28239));
	notech_inv i_32267(.A(regs_12[15]), .Z(n_28240));
	notech_inv i_32268(.A(regs_12[16]), .Z(n_28241));
	notech_inv i_32269(.A(regs_12[17]), .Z(n_28242));
	notech_inv i_32270(.A(regs_12[18]), .Z(n_28243));
	notech_inv i_32271(.A(regs_12[19]), .Z(n_28244));
	notech_inv i_32272(.A(regs_12[20]), .Z(n_28245));
	notech_inv i_32273(.A(regs_12[21]), .Z(n_28246));
	notech_inv i_32274(.A(regs_12[22]), .Z(n_28247));
	notech_inv i_32275(.A(regs_12[23]), .Z(n_28248));
	notech_inv i_32276(.A(regs_12[24]), .Z(n_28249));
	notech_inv i_32277(.A(regs_12[25]), .Z(n_28250));
	notech_inv i_32278(.A(regs_12[26]), .Z(n_28251));
	notech_inv i_32279(.A(regs_12[27]), .Z(n_28252));
	notech_inv i_32280(.A(regs_12[28]), .Z(n_28253));
	notech_inv i_32281(.A(regs_12[29]), .Z(n_28254));
	notech_inv i_32282(.A(regs_12[30]), .Z(n_28255));
	notech_inv i_32283(.A(regs_12[31]), .Z(n_28256));
	notech_inv i_32284(.A(gs[0]), .Z(n_28257));
	notech_inv i_32285(.A(gs[1]), .Z(n_28258));
	notech_inv i_32286(.A(n_56005), .Z(n_28259));
	notech_inv i_32287(.A(gs[3]), .Z(n_28260));
	notech_inv i_32288(.A(gs[4]), .Z(n_28261));
	notech_inv i_32289(.A(gs[5]), .Z(n_28262));
	notech_inv i_32290(.A(gs[6]), .Z(n_28263));
	notech_inv i_32291(.A(gs[7]), .Z(n_28264));
	notech_inv i_32292(.A(gs[8]), .Z(n_28265));
	notech_inv i_32293(.A(gs[9]), .Z(n_28266));
	notech_inv i_32294(.A(gs[10]), .Z(n_28267));
	notech_inv i_32295(.A(gs[11]), .Z(n_28268));
	notech_inv i_32296(.A(gs[12]), .Z(n_28269));
	notech_inv i_32297(.A(gs[13]), .Z(n_28270));
	notech_inv i_32298(.A(gs[14]), .Z(n_28271));
	notech_inv i_32299(.A(gs[15]), .Z(n_28272));
	notech_inv i_32300(.A(gs[16]), .Z(n_28273));
	notech_inv i_32301(.A(gs[17]), .Z(n_28274));
	notech_inv i_32302(.A(gs[18]), .Z(n_28275));
	notech_inv i_32303(.A(gs[19]), .Z(n_28276));
	notech_inv i_32304(.A(gs[20]), .Z(n_28277));
	notech_inv i_32305(.A(gs[21]), .Z(n_28278));
	notech_inv i_32306(.A(gs[22]), .Z(n_28279));
	notech_inv i_32307(.A(gs[23]), .Z(n_28280));
	notech_inv i_32308(.A(gs[24]), .Z(n_28281));
	notech_inv i_32309(.A(gs[25]), .Z(n_28282));
	notech_inv i_32310(.A(gs[26]), .Z(n_28283));
	notech_inv i_32311(.A(gs[27]), .Z(n_28284));
	notech_inv i_32312(.A(gs[28]), .Z(n_28285));
	notech_inv i_32313(.A(gs[29]), .Z(n_28286));
	notech_inv i_32314(.A(gs[30]), .Z(n_28287));
	notech_inv i_32315(.A(gs[31]), .Z(n_28288));
	notech_inv i_32316(.A(regs_2[0]), .Z(n_28289));
	notech_inv i_32317(.A(regs_2[1]), .Z(n_28290));
	notech_inv i_32318(.A(regs_2[2]), .Z(n_28291));
	notech_inv i_32319(.A(regs_2[3]), .Z(n_28292));
	notech_inv i_32320(.A(regs_2[4]), .Z(n_28293));
	notech_inv i_32321(.A(regs_2[5]), .Z(n_28294));
	notech_inv i_32322(.A(regs_2[6]), .Z(n_28295));
	notech_inv i_32323(.A(regs_2[7]), .Z(n_28296));
	notech_inv i_32324(.A(regs_2[8]), .Z(n_28297));
	notech_inv i_32325(.A(regs_2[9]), .Z(n_28298));
	notech_inv i_32326(.A(regs_2[10]), .Z(n_28299));
	notech_inv i_32327(.A(regs_2[11]), .Z(n_28301));
	notech_inv i_32328(.A(regs_2[12]), .Z(n_28302));
	notech_inv i_32329(.A(regs_2[13]), .Z(n_28303));
	notech_inv i_32330(.A(regs_2[14]), .Z(n_28304));
	notech_inv i_32331(.A(regs_2[15]), .Z(n_28305));
	notech_inv i_32332(.A(regs_2[16]), .Z(n_28306));
	notech_inv i_32333(.A(regs_2[17]), .Z(n_28307));
	notech_inv i_32334(.A(regs_2[18]), .Z(n_28308));
	notech_inv i_32335(.A(regs_2[19]), .Z(n_28309));
	notech_inv i_32336(.A(regs_2[20]), .Z(n_28310));
	notech_inv i_32337(.A(regs_2[21]), .Z(n_28311));
	notech_inv i_32338(.A(regs_2[22]), .Z(n_28312));
	notech_inv i_32339(.A(regs_2[23]), .Z(n_28313));
	notech_inv i_32340(.A(regs_2[24]), .Z(n_28314));
	notech_inv i_32341(.A(regs_2[25]), .Z(n_28315));
	notech_inv i_32342(.A(regs_2[26]), .Z(n_28316));
	notech_inv i_32343(.A(regs_2[27]), .Z(n_28317));
	notech_inv i_32344(.A(regs_2[28]), .Z(n_28318));
	notech_inv i_32345(.A(regs_2[29]), .Z(n_28319));
	notech_inv i_32346(.A(regs_2[30]), .Z(n_28320));
	notech_inv i_32347(.A(regs_2[31]), .Z(n_28321));
	notech_inv i_32348(.A(regs_5[0]), .Z(n_28322));
	notech_inv i_32349(.A(regs_5[1]), .Z(n_28323));
	notech_inv i_32350(.A(regs_5[2]), .Z(n_28324));
	notech_inv i_32351(.A(regs_5[3]), .Z(n_28325));
	notech_inv i_32352(.A(regs_5[4]), .Z(n_28326));
	notech_inv i_32353(.A(regs_5[5]), .Z(n_28327));
	notech_inv i_32354(.A(regs_5[6]), .Z(n_28328));
	notech_inv i_32355(.A(regs_5[7]), .Z(n_28329));
	notech_inv i_32356(.A(regs_5[8]), .Z(n_28330));
	notech_inv i_32357(.A(regs_5[9]), .Z(n_28331));
	notech_inv i_32358(.A(regs_5[10]), .Z(n_28333));
	notech_inv i_32360(.A(regs_5[11]), .Z(n_28334));
	notech_inv i_32361(.A(regs_5[12]), .Z(n_28335));
	notech_inv i_32362(.A(regs_5[13]), .Z(n_28336));
	notech_inv i_32364(.A(regs_5[14]), .Z(n_28337));
	notech_inv i_32365(.A(regs_5[15]), .Z(n_28338));
	notech_inv i_32367(.A(regs_5[16]), .Z(n_28339));
	notech_inv i_32368(.A(regs_5[17]), .Z(n_28340));
	notech_inv i_32369(.A(regs_5[18]), .Z(n_28341));
	notech_inv i_32370(.A(regs_5[19]), .Z(n_28342));
	notech_inv i_32372(.A(regs_5[20]), .Z(n_28343));
	notech_inv i_32373(.A(regs_5[21]), .Z(n_28344));
	notech_inv i_32375(.A(regs_5[22]), .Z(n_28345));
	notech_inv i_32376(.A(regs_5[23]), .Z(n_28346));
	notech_inv i_32377(.A(regs_5[24]), .Z(n_28347));
	notech_inv i_32378(.A(regs_5[25]), .Z(n_28348));
	notech_inv i_32379(.A(regs_5[26]), .Z(n_28349));
	notech_inv i_32380(.A(regs_5[27]), .Z(n_28350));
	notech_inv i_32381(.A(regs_5[28]), .Z(n_28351));
	notech_inv i_32382(.A(regs_5[29]), .Z(n_28352));
	notech_inv i_32383(.A(regs_5[30]), .Z(n_28353));
	notech_inv i_32384(.A(regs_5[31]), .Z(n_28354));
	notech_inv i_32385(.A(regs_8[0]), .Z(n_28355));
	notech_inv i_32386(.A(regs_8[1]), .Z(n_28356));
	notech_inv i_32387(.A(regs_8[2]), .Z(n_28357));
	notech_inv i_32388(.A(regs_8[3]), .Z(n_28358));
	notech_inv i_32389(.A(regs_8[4]), .Z(n_28359));
	notech_inv i_32390(.A(regs_8[5]), .Z(n_28360));
	notech_inv i_32391(.A(regs_8[6]), .Z(n_28361));
	notech_inv i_32392(.A(regs_8[7]), .Z(n_28362));
	notech_inv i_32393(.A(regs_8[8]), .Z(n_28363));
	notech_inv i_32394(.A(regs_8[9]), .Z(n_28364));
	notech_inv i_32395(.A(regs_8[10]), .Z(n_28365));
	notech_inv i_32397(.A(regs_8[11]), .Z(n_28366));
	notech_inv i_32398(.A(regs_8[12]), .Z(n_28367));
	notech_inv i_32400(.A(regs_8[13]), .Z(n_28368));
	notech_inv i_32401(.A(regs_8[14]), .Z(n_28369));
	notech_inv i_32403(.A(regs_8[15]), .Z(n_28370));
	notech_inv i_32404(.A(regs_8[16]), .Z(n_28371));
	notech_inv i_32406(.A(regs_8[17]), .Z(n_28372));
	notech_inv i_32407(.A(regs_8[18]), .Z(n_28373));
	notech_inv i_32408(.A(regs_8[19]), .Z(n_28374));
	notech_inv i_32409(.A(regs_8[20]), .Z(n_28375));
	notech_inv i_32410(.A(regs_8[21]), .Z(n_28376));
	notech_inv i_32411(.A(regs_8[22]), .Z(n_28377));
	notech_inv i_32412(.A(regs_8[23]), .Z(n_28378));
	notech_inv i_32413(.A(regs_8[24]), .Z(n_28379));
	notech_inv i_32414(.A(regs_8[25]), .Z(n_28380));
	notech_inv i_32415(.A(regs_8[26]), .Z(n_28381));
	notech_inv i_32416(.A(regs_8[27]), .Z(n_28382));
	notech_inv i_32417(.A(regs_8[28]), .Z(n_28383));
	notech_inv i_32418(.A(regs_8[29]), .Z(n_28384));
	notech_inv i_32419(.A(regs_8[30]), .Z(n_28385));
	notech_inv i_32420(.A(regs_8[31]), .Z(n_28386));
	notech_inv i_32421(.A(regs_4[0]), .Z(n_28387));
	notech_inv i_32422(.A(regs_4[1]), .Z(n_28388));
	notech_inv i_32423(.A(regs_4[2]), .Z(n_28389));
	notech_inv i_32424(.A(regs_4[3]), .Z(n_28390));
	notech_inv i_32425(.A(regs_4[4]), .Z(n_28391));
	notech_inv i_32426(.A(regs_4[5]), .Z(n_28392));
	notech_inv i_32428(.A(regs_4[6]), .Z(n_28393));
	notech_inv i_32429(.A(regs_4[7]), .Z(n_28394));
	notech_inv i_32430(.A(regs_4[8]), .Z(n_28395));
	notech_inv i_32431(.A(regs_4[9]), .Z(n_28396));
	notech_inv i_32432(.A(regs_4[10]), .Z(n_28397));
	notech_inv i_32433(.A(regs_4[11]), .Z(n_28398));
	notech_inv i_32434(.A(regs_4[12]), .Z(n_28399));
	notech_inv i_32435(.A(regs_4[13]), .Z(n_28400));
	notech_inv i_32436(.A(regs_4[14]), .Z(n_28401));
	notech_inv i_32437(.A(regs_4[15]), .Z(n_28402));
	notech_inv i_32438(.A(regs_4[16]), .Z(n_28403));
	notech_inv i_32439(.A(regs_4[17]), .Z(n_28404));
	notech_inv i_32440(.A(regs_4[18]), .Z(n_28405));
	notech_inv i_32441(.A(regs_4[19]), .Z(n_28406));
	notech_inv i_32442(.A(regs_4[20]), .Z(n_28407));
	notech_inv i_32443(.A(regs_4[21]), .Z(n_28408));
	notech_inv i_32444(.A(regs_4[22]), .Z(n_28409));
	notech_inv i_32445(.A(regs_4[23]), .Z(n_28410));
	notech_inv i_32446(.A(regs_4[24]), .Z(n_28411));
	notech_inv i_32447(.A(regs_4[25]), .Z(n_28412));
	notech_inv i_32448(.A(regs_4[26]), .Z(n_28413));
	notech_inv i_32449(.A(regs_4[27]), .Z(n_28414));
	notech_inv i_32450(.A(regs_4[28]), .Z(n_28415));
	notech_inv i_32451(.A(regs_4[29]), .Z(n_28416));
	notech_inv i_32452(.A(regs_4[30]), .Z(n_28417));
	notech_inv i_32453(.A(regs_4[31]), .Z(n_28418));
	notech_inv i_32454(.A(regs_10[0]), .Z(n_28419));
	notech_inv i_32455(.A(regs_10[1]), .Z(n_28420));
	notech_inv i_32456(.A(regs_10[2]), .Z(n_28421));
	notech_inv i_32457(.A(regs_10[3]), .Z(n_28422));
	notech_inv i_32458(.A(regs_10[4]), .Z(n_28423));
	notech_inv i_32459(.A(regs_10[5]), .Z(n_28424));
	notech_inv i_32460(.A(regs_10[6]), .Z(n_28425));
	notech_inv i_32461(.A(regs_10[7]), .Z(n_28426));
	notech_inv i_32462(.A(regs_10[8]), .Z(n_28427));
	notech_inv i_32463(.A(regs_10[9]), .Z(n_28428));
	notech_inv i_32464(.A(regs_10[10]), .Z(n_28429));
	notech_inv i_32467(.A(regs_10[11]), .Z(n_28430));
	notech_inv i_32468(.A(regs_10[12]), .Z(n_28431));
	notech_inv i_32469(.A(regs_10[13]), .Z(n_28432));
	notech_inv i_32470(.A(regs_10[14]), .Z(n_28433));
	notech_inv i_32471(.A(regs_10[15]), .Z(n_28434));
	notech_inv i_32473(.A(regs_10[16]), .Z(n_28435));
	notech_inv i_32474(.A(regs_10[17]), .Z(n_28436));
	notech_inv i_32475(.A(regs_10[18]), .Z(n_28437));
	notech_inv i_32477(.A(regs_10[19]), .Z(n_28438));
	notech_inv i_32478(.A(regs_10[20]), .Z(n_28439));
	notech_inv i_32479(.A(regs_10[21]), .Z(n_28440));
	notech_inv i_32480(.A(regs_10[22]), .Z(n_28441));
	notech_inv i_32481(.A(regs_10[23]), .Z(n_28442));
	notech_inv i_32482(.A(regs_10[24]), .Z(n_28443));
	notech_inv i_32483(.A(regs_10[25]), .Z(n_28444));
	notech_inv i_32484(.A(regs_10[26]), .Z(n_28445));
	notech_inv i_32485(.A(regs_10[27]), .Z(n_28446));
	notech_inv i_32486(.A(regs_10[28]), .Z(n_28447));
	notech_inv i_32487(.A(regs_10[29]), .Z(n_28448));
	notech_inv i_32489(.A(regs_10[30]), .Z(n_28449));
	notech_inv i_32490(.A(regs_10[31]), .Z(n_28450));
	notech_inv i_32491(.A(regs_3[0]), .Z(n_28451));
	notech_inv i_32492(.A(regs_3[1]), .Z(n_28452));
	notech_inv i_32493(.A(regs_3[2]), .Z(n_28453));
	notech_inv i_32494(.A(regs_3[3]), .Z(n_28454));
	notech_inv i_32495(.A(regs_3[4]), .Z(n_28455));
	notech_inv i_32496(.A(regs_3[5]), .Z(n_28456));
	notech_inv i_32497(.A(regs_3[6]), .Z(n_28457));
	notech_inv i_32498(.A(regs_3[7]), .Z(n_28458));
	notech_inv i_32499(.A(regs_3[8]), .Z(n_28459));
	notech_inv i_32500(.A(regs_3[9]), .Z(n_28460));
	notech_inv i_32501(.A(regs_3[10]), .Z(n_28461));
	notech_inv i_32502(.A(regs_3[11]), .Z(n_28462));
	notech_inv i_32503(.A(regs_3[12]), .Z(n_28463));
	notech_inv i_32504(.A(regs_3[13]), .Z(n_28464));
	notech_inv i_32505(.A(regs_3[14]), .Z(n_28465));
	notech_inv i_32506(.A(regs_3[15]), .Z(n_28466));
	notech_inv i_32508(.A(regs_3[16]), .Z(n_28467));
	notech_inv i_32509(.A(regs_3[17]), .Z(n_28468));
	notech_inv i_32510(.A(regs_3[18]), .Z(n_28469));
	notech_inv i_32511(.A(regs_3[19]), .Z(n_28470));
	notech_inv i_32512(.A(regs_3[20]), .Z(n_28471));
	notech_inv i_32513(.A(regs_3[21]), .Z(n_28472));
	notech_inv i_32514(.A(regs_3[22]), .Z(n_28473));
	notech_inv i_32515(.A(regs_3[23]), .Z(n_28474));
	notech_inv i_32516(.A(regs_3[24]), .Z(n_28475));
	notech_inv i_32517(.A(regs_3[25]), .Z(n_28476));
	notech_inv i_32518(.A(regs_3[26]), .Z(n_28477));
	notech_inv i_32519(.A(regs_3[27]), .Z(n_28478));
	notech_inv i_32520(.A(regs_3[28]), .Z(n_28479));
	notech_inv i_32521(.A(regs_3[29]), .Z(n_28480));
	notech_inv i_32522(.A(regs_3[30]), .Z(n_28481));
	notech_inv i_32523(.A(regs_3[31]), .Z(n_28482));
	notech_inv i_32524(.A(regs_0[0]), .Z(n_28483));
	notech_inv i_32525(.A(regs_0[1]), .Z(n_28484));
	notech_inv i_32526(.A(regs_0[2]), .Z(n_28485));
	notech_inv i_32527(.A(regs_0[3]), .Z(n_28486));
	notech_inv i_32528(.A(regs_0[4]), .Z(n_28487));
	notech_inv i_32529(.A(regs_0[5]), .Z(n_28488));
	notech_inv i_32530(.A(regs_0[6]), .Z(n_28489));
	notech_inv i_32531(.A(regs_0[7]), .Z(n_28490));
	notech_inv i_32532(.A(regs_0[8]), .Z(n_28491));
	notech_inv i_32533(.A(regs_0[9]), .Z(n_28492));
	notech_inv i_32534(.A(regs_0[10]), .Z(n_28493));
	notech_inv i_32535(.A(regs_0[11]), .Z(n_28494));
	notech_inv i_32536(.A(regs_0[12]), .Z(n_28495));
	notech_inv i_32537(.A(regs_0[13]), .Z(n_28496));
	notech_inv i_32538(.A(regs_0[14]), .Z(n_28497));
	notech_inv i_32539(.A(regs_0[15]), .Z(n_28498));
	notech_inv i_32540(.A(regs_0[16]), .Z(n_28499));
	notech_inv i_32541(.A(regs_0[17]), .Z(n_28500));
	notech_inv i_32542(.A(regs_0[18]), .Z(n_28501));
	notech_inv i_32543(.A(regs_0[19]), .Z(n_28503));
	notech_inv i_32544(.A(regs_0[20]), .Z(n_28504));
	notech_inv i_32545(.A(regs_0[21]), .Z(n_28505));
	notech_inv i_32546(.A(regs_0[22]), .Z(n_28506));
	notech_inv i_32547(.A(regs_0[23]), .Z(n_28507));
	notech_inv i_32548(.A(regs_0[24]), .Z(n_28508));
	notech_inv i_32549(.A(regs_0[25]), .Z(n_28509));
	notech_inv i_32550(.A(regs_0[26]), .Z(n_28510));
	notech_inv i_32551(.A(regs_0[27]), .Z(n_28511));
	notech_inv i_32552(.A(regs_0[28]), .Z(n_28512));
	notech_inv i_32553(.A(regs_0[29]), .Z(n_28513));
	notech_inv i_32554(.A(regs_0[30]), .Z(n_28514));
	notech_inv i_32555(.A(regs_0[31]), .Z(n_28515));
	notech_inv i_32556(.A(regs_7[0]), .Z(n_28516));
	notech_inv i_32557(.A(regs_7[1]), .Z(n_28517));
	notech_inv i_32558(.A(regs_7[2]), .Z(n_28518));
	notech_inv i_32559(.A(regs_7[3]), .Z(n_28519));
	notech_inv i_32560(.A(regs_7[4]), .Z(n_28520));
	notech_inv i_32561(.A(regs_7[5]), .Z(n_28521));
	notech_inv i_32562(.A(regs_7[6]), .Z(n_28522));
	notech_inv i_32563(.A(regs_7[7]), .Z(n_28523));
	notech_inv i_32564(.A(regs_7[8]), .Z(n_28525));
	notech_inv i_32565(.A(regs_7[9]), .Z(n_28526));
	notech_inv i_32566(.A(regs_7[10]), .Z(n_28528));
	notech_inv i_32567(.A(regs_7[11]), .Z(n_28529));
	notech_inv i_32568(.A(regs_7[12]), .Z(n_28531));
	notech_inv i_32569(.A(regs_7[13]), .Z(n_28534));
	notech_inv i_32570(.A(regs_7[14]), .Z(n_28535));
	notech_inv i_32571(.A(regs_7[15]), .Z(n_28536));
	notech_inv i_32572(.A(regs_7[16]), .Z(n_28537));
	notech_inv i_32573(.A(regs_7[17]), .Z(n_28538));
	notech_inv i_32574(.A(regs_7[18]), .Z(n_28539));
	notech_inv i_32575(.A(regs_7[19]), .Z(n_28540));
	notech_inv i_32576(.A(regs_7[20]), .Z(n_28541));
	notech_inv i_32577(.A(regs_7[21]), .Z(n_28547));
	notech_inv i_32578(.A(regs_7[22]), .Z(n_28548));
	notech_inv i_32579(.A(regs_7[23]), .Z(n_28549));
	notech_inv i_32580(.A(regs_7[24]), .Z(n_28550));
	notech_inv i_32581(.A(regs_7[25]), .Z(n_28553));
	notech_inv i_32582(.A(regs_7[26]), .Z(n_28554));
	notech_inv i_32583(.A(regs_7[27]), .Z(n_28555));
	notech_inv i_32584(.A(regs_7[28]), .Z(n_28556));
	notech_inv i_32585(.A(regs_7[29]), .Z(n_28557));
	notech_inv i_32586(.A(regs_7[30]), .Z(n_28558));
	notech_inv i_32587(.A(regs_7[31]), .Z(n_28559));
	notech_inv i_32588(.A(regs_6[0]), .Z(n_28560));
	notech_inv i_32589(.A(regs_6[1]), .Z(n_28561));
	notech_inv i_32590(.A(regs_6[2]), .Z(n_28562));
	notech_inv i_32591(.A(regs_6[3]), .Z(n_28563));
	notech_inv i_32592(.A(regs_6[4]), .Z(n_28564));
	notech_inv i_32593(.A(regs_6[5]), .Z(n_28565));
	notech_inv i_32594(.A(regs_6[6]), .Z(n_28566));
	notech_inv i_32595(.A(regs_6[7]), .Z(n_28567));
	notech_inv i_32596(.A(regs_6[8]), .Z(n_28568));
	notech_inv i_32597(.A(regs_6[9]), .Z(n_28570));
	notech_inv i_32598(.A(regs_6[10]), .Z(n_28571));
	notech_inv i_32599(.A(regs_6[11]), .Z(n_28572));
	notech_inv i_32600(.A(regs_6[12]), .Z(n_28573));
	notech_inv i_32601(.A(regs_6[13]), .Z(n_28574));
	notech_inv i_32602(.A(regs_6[14]), .Z(n_28575));
	notech_inv i_32603(.A(regs_6[15]), .Z(n_28576));
	notech_inv i_32604(.A(regs_6[16]), .Z(n_28577));
	notech_inv i_32605(.A(regs_6[17]), .Z(n_28578));
	notech_inv i_32606(.A(regs_6[18]), .Z(n_28579));
	notech_inv i_32607(.A(regs_6[19]), .Z(n_28580));
	notech_inv i_32608(.A(regs_6[20]), .Z(n_28581));
	notech_inv i_32609(.A(regs_6[21]), .Z(n_28582));
	notech_inv i_32610(.A(regs_6[22]), .Z(n_28583));
	notech_inv i_32611(.A(regs_6[23]), .Z(n_28584));
	notech_inv i_32612(.A(regs_6[24]), .Z(n_28585));
	notech_inv i_32613(.A(regs_6[25]), .Z(n_28586));
	notech_inv i_32614(.A(regs_6[26]), .Z(n_28587));
	notech_inv i_32615(.A(regs_6[27]), .Z(n_28588));
	notech_inv i_32616(.A(regs_6[28]), .Z(n_28589));
	notech_inv i_32617(.A(regs_6[29]), .Z(n_28590));
	notech_inv i_32618(.A(regs_6[30]), .Z(n_28591));
	notech_inv i_32619(.A(regs_6[31]), .Z(n_28592));
	notech_inv i_32620(.A(regs_4_2[0]), .Z(n_28593));
	notech_inv i_32622(.A(regs_4_2[1]), .Z(n_28594));
	notech_inv i_32623(.A(regs_4_2[2]), .Z(n_28595));
	notech_inv i_32624(.A(regs_4_2[3]), .Z(n_28596));
	notech_inv i_32625(.A(regs_4_2[4]), .Z(n_28597));
	notech_inv i_32626(.A(regs_4_2[5]), .Z(n_28598));
	notech_inv i_32627(.A(regs_4_2[6]), .Z(n_28599));
	notech_inv i_32628(.A(regs_4_2[7]), .Z(n_28600));
	notech_inv i_32629(.A(regs_4_2[8]), .Z(n_28601));
	notech_inv i_32630(.A(regs_4_2[9]), .Z(n_28602));
	notech_inv i_32631(.A(regs_4_2[10]), .Z(n_28603));
	notech_inv i_32632(.A(regs_4_2[11]), .Z(n_28604));
	notech_inv i_32633(.A(regs_4_2[12]), .Z(n_28605));
	notech_inv i_32635(.A(regs_4_2[13]), .Z(n_28606));
	notech_inv i_32637(.A(regs_4_2[14]), .Z(n_28607));
	notech_inv i_32638(.A(regs_4_2[15]), .Z(n_28608));
	notech_inv i_32639(.A(regs_4_2[16]), .Z(n_28609));
	notech_inv i_32640(.A(regs_4_2[17]), .Z(n_28610));
	notech_inv i_32641(.A(regs_4_2[18]), .Z(n_28611));
	notech_inv i_32642(.A(regs_4_2[19]), .Z(n_28612));
	notech_inv i_32643(.A(regs_4_2[20]), .Z(n_28613));
	notech_inv i_32644(.A(regs_4_2[21]), .Z(n_28614));
	notech_inv i_32645(.A(regs_4_2[22]), .Z(n_28615));
	notech_inv i_32646(.A(regs_4_2[23]), .Z(n_28616));
	notech_inv i_32647(.A(regs_4_2[24]), .Z(n_28617));
	notech_inv i_32648(.A(regs_4_2[25]), .Z(n_28618));
	notech_inv i_32649(.A(regs_4_2[26]), .Z(n_28619));
	notech_inv i_32650(.A(regs_4_2[27]), .Z(n_28620));
	notech_inv i_32651(.A(regs_4_2[28]), .Z(n_28621));
	notech_inv i_32652(.A(regs_4_2[29]), .Z(n_28622));
	notech_inv i_32653(.A(regs_4_2[30]), .Z(n_28623));
	notech_inv i_32654(.A(regs_4_2[31]), .Z(n_28624));
	notech_inv i_32655(.A(nbus_159[0]), .Z(n_28625));
	notech_inv i_32656(.A(nbus_159[1]), .Z(n_28626));
	notech_inv i_32657(.A(nbus_159[2]), .Z(n_28627));
	notech_inv i_32658(.A(nbus_159[3]), .Z(n_28628));
	notech_inv i_32659(.A(nbus_159[4]), .Z(n_28629));
	notech_inv i_32660(.A(nbus_159[5]), .Z(n_28631));
	notech_inv i_32661(.A(nbus_159[6]), .Z(n_28632));
	notech_inv i_32662(.A(nbus_159[7]), .Z(n_28634));
	notech_inv i_32663(.A(nbus_159[8]), .Z(n_28635));
	notech_inv i_32664(.A(nbus_163[2]), .Z(n_28637));
	notech_inv i_32665(.A(nbus_163[5]), .Z(n_28638));
	notech_inv i_32666(.A(nbus_163[7]), .Z(n_28639));
	notech_inv i_32667(.A(nbus_163[8]), .Z(n_28640));
	notech_inv i_32668(.A(nbus_163[9]), .Z(n_28641));
	notech_inv i_32669(.A(nbus_163[10]), .Z(n_28642));
	notech_inv i_32670(.A(nbus_163[11]), .Z(n_28643));
	notech_inv i_32671(.A(nbus_163[12]), .Z(n_28644));
	notech_inv i_32672(.A(nbus_163[13]), .Z(n_28645));
	notech_inv i_32673(.A(nbus_163[14]), .Z(n_28647));
	notech_inv i_32674(.A(nbus_163[15]), .Z(n_28648));
	notech_inv i_32675(.A(nbus_165[0]), .Z(n_28649));
	notech_inv i_32676(.A(nbus_165[1]), .Z(n_28650));
	notech_inv i_32677(.A(nbus_165[2]), .Z(n_28652));
	notech_inv i_32678(.A(nbus_165[3]), .Z(n_28653));
	notech_inv i_32679(.A(nbus_165[4]), .Z(n_28654));
	notech_inv i_32680(.A(nbus_165[5]), .Z(n_28657));
	notech_inv i_32681(.A(nbus_165[6]), .Z(n_28658));
	notech_inv i_32682(.A(nbus_165[7]), .Z(n_28659));
	notech_inv i_32683(.A(nbus_165[8]), .Z(n_28660));
	notech_inv i_32684(.A(nbus_165[9]), .Z(n_28661));
	notech_inv i_32685(.A(nbus_165[10]), .Z(n_28662));
	notech_inv i_32686(.A(nbus_165[11]), .Z(n_28663));
	notech_inv i_32687(.A(nbus_165[12]), .Z(n_28664));
	notech_inv i_32688(.A(nbus_165[13]), .Z(n_28665));
	notech_inv i_32689(.A(nbus_165[14]), .Z(n_28666));
	notech_inv i_32690(.A(nbus_165[15]), .Z(n_28667));
	notech_inv i_32691(.A(nbus_165[16]), .Z(n_28668));
	notech_inv i_32692(.A(nbus_158[5]), .Z(n_28669));
	notech_inv i_32693(.A(nbus_158[7]), .Z(n_28670));
	notech_inv i_32694(.A(nbus_158[8]), .Z(n_28671));
	notech_inv i_32695(.A(nbus_158[9]), .Z(n_28672));
	notech_inv i_32696(.A(nbus_158[10]), .Z(n_28673));
	notech_inv i_32697(.A(nbus_158[11]), .Z(n_28674));
	notech_inv i_32698(.A(nbus_158[12]), .Z(n_28675));
	notech_inv i_32699(.A(nbus_158[13]), .Z(n_28676));
	notech_inv i_32700(.A(nbus_158[14]), .Z(n_28677));
	notech_inv i_32701(.A(nbus_158[15]), .Z(n_28678));
	notech_inv i_32702(.A(nbus_158[16]), .Z(n_28679));
	notech_inv i_32703(.A(n_60542), .Z(n_28680));
	notech_inv i_32704(.A(cr0[2]), .Z(n_28681));
	notech_inv i_32705(.A(cr0[16]), .Z(n_28682));
	notech_inv i_32706(.A(resa_shift4box[0]), .Z(n_28683));
	notech_inv i_32707(.A(resa_shift4box[1]), .Z(n_28684));
	notech_inv i_32708(.A(resa_shift4box[2]), .Z(n_28685));
	notech_inv i_32709(.A(resa_shift4box[3]), .Z(n_28686));
	notech_inv i_32710(.A(resa_shift4box[4]), .Z(n_28687));
	notech_inv i_32711(.A(resa_shift4box[6]), .Z(n_28688));
	notech_inv i_32712(.A(resa_shift4box[7]), .Z(n_28689));
	notech_inv i_32713(.A(resa_shift4box[8]), .Z(n_28690));
	notech_inv i_32714(.A(resa_shift4box[9]), .Z(n_28691));
	notech_inv i_32715(.A(resa_shift4box[10]), .Z(n_28692));
	notech_inv i_32716(.A(resa_shift4box[11]), .Z(n_28693));
	notech_inv i_32717(.A(resa_shift4box[12]), .Z(n_28694));
	notech_inv i_32718(.A(resa_shift4box[13]), .Z(n_28695));
	notech_inv i_32719(.A(resa_shift4box[14]), .Z(n_28696));
	notech_inv i_32720(.A(resa_shift4box[15]), .Z(n_28697));
	notech_inv i_32721(.A(cr3[12]), .Z(n_28698));
	notech_inv i_32722(.A(cr3[13]), .Z(n_28699));
	notech_inv i_32723(.A(cr3[14]), .Z(n_28700));
	notech_inv i_32724(.A(cr3[15]), .Z(n_28701));
	notech_inv i_32725(.A(cr3[16]), .Z(n_28702));
	notech_inv i_32726(.A(cr3[17]), .Z(n_28703));
	notech_inv i_32727(.A(cr3[18]), .Z(n_28704));
	notech_inv i_32728(.A(cr3[19]), .Z(n_28705));
	notech_inv i_32729(.A(cr3[20]), .Z(n_28706));
	notech_inv i_32730(.A(cr3[21]), .Z(n_28707));
	notech_inv i_32731(.A(cr3[22]), .Z(n_28708));
	notech_inv i_32732(.A(cr3[23]), .Z(n_28709));
	notech_inv i_32733(.A(cr3[24]), .Z(n_28710));
	notech_inv i_32734(.A(cr3[25]), .Z(n_28711));
	notech_inv i_32735(.A(cr3[26]), .Z(n_28712));
	notech_inv i_32736(.A(cr3[27]), .Z(n_28713));
	notech_inv i_32737(.A(cr3[28]), .Z(n_28714));
	notech_inv i_32738(.A(cr3[29]), .Z(n_28715));
	notech_inv i_32739(.A(cr3[30]), .Z(n_28716));
	notech_inv i_32740(.A(cr3[31]), .Z(n_28717));
	notech_inv i_32741(.A(resa_arithbox[0]), .Z(n_28718));
	notech_inv i_32742(.A(resa_arithbox[1]), .Z(n_28719));
	notech_inv i_32743(.A(resa_arithbox[2]), .Z(n_28720));
	notech_inv i_32744(.A(resa_arithbox[3]), .Z(n_28723));
	notech_inv i_32745(.A(resa_arithbox[4]), .Z(n_28725));
	notech_inv i_32746(.A(resa_arithbox[6]), .Z(n_28726));
	notech_inv i_32747(.A(resa_arithbox[7]), .Z(n_28727));
	notech_inv i_32748(.A(resa_arithbox[8]), .Z(n_28728));
	notech_inv i_32749(.A(resa_arithbox[9]), .Z(n_28729));
	notech_inv i_32750(.A(resa_arithbox[10]), .Z(n_28730));
	notech_inv i_32751(.A(resa_arithbox[11]), .Z(n_28732));
	notech_inv i_32752(.A(resa_arithbox[12]), .Z(n_28733));
	notech_inv i_32753(.A(resa_arithbox[13]), .Z(n_28735));
	notech_inv i_32754(.A(resa_arithbox[14]), .Z(n_28736));
	notech_inv i_32755(.A(resa_arithbox[31]), .Z(n_28737));
	notech_inv i_32756(.A(opa_0[0]), .Z(n_28738));
	notech_inv i_32757(.A(opa_0[1]), .Z(n_28739));
	notech_inv i_32758(.A(opa_0[2]), .Z(n_28740));
	notech_inv i_32759(.A(opa_0[3]), .Z(n_28741));
	notech_inv i_32760(.A(opa_0[4]), .Z(n_28742));
	notech_inv i_32761(.A(opa_0[5]), .Z(n_28743));
	notech_inv i_32762(.A(opa_0[6]), .Z(n_28744));
	notech_inv i_32763(.A(opa_0[7]), .Z(n_28745));
	notech_inv i_32764(.A(opa_0[8]), .Z(n_28746));
	notech_inv i_32765(.A(opa_0[9]), .Z(n_28747));
	notech_inv i_32766(.A(opa_0[10]), .Z(n_28748));
	notech_inv i_32767(.A(opa_0[11]), .Z(n_28749));
	notech_inv i_32768(.A(opa_0[12]), .Z(n_28750));
	notech_inv i_32769(.A(opa_0[13]), .Z(n_28751));
	notech_inv i_32770(.A(opa_0[14]), .Z(n_28752));
	notech_inv i_32771(.A(opa_0[15]), .Z(n_28753));
	notech_inv i_32772(.A(opa_0[16]), .Z(n_28754));
	notech_inv i_32773(.A(opa_0[17]), .Z(n_28755));
	notech_inv i_32774(.A(opa_0[18]), .Z(n_28756));
	notech_inv i_32775(.A(opa_0[19]), .Z(n_28757));
	notech_inv i_32776(.A(opa_0[20]), .Z(n_28758));
	notech_inv i_32777(.A(opa_0[21]), .Z(n_28759));
	notech_inv i_32778(.A(opa_0[22]), .Z(n_28760));
	notech_inv i_32779(.A(opa_0[23]), .Z(n_28761));
	notech_inv i_32780(.A(opa_0[24]), .Z(n_28762));
	notech_inv i_32781(.A(opa_0[25]), .Z(n_28763));
	notech_inv i_32782(.A(opa_0[26]), .Z(n_28764));
	notech_inv i_32783(.A(opa_0[27]), .Z(n_28765));
	notech_inv i_32784(.A(opa_0[28]), .Z(n_28766));
	notech_inv i_32785(.A(opa_0[29]), .Z(n_28767));
	notech_inv i_32786(.A(opa_0[30]), .Z(n_28768));
	notech_inv i_32787(.A(opa_0[31]), .Z(n_28769));
	notech_inv i_32788(.A(nbus_157[0]), .Z(n_28770));
	notech_inv i_32789(.A(nbus_157[1]), .Z(n_28771));
	notech_inv i_32790(.A(nbus_157[2]), .Z(n_28772));
	notech_inv i_32791(.A(nbus_157[3]), .Z(n_28773));
	notech_inv i_32792(.A(nbus_157[4]), .Z(n_28774));
	notech_inv i_32793(.A(nbus_157[5]), .Z(n_28775));
	notech_inv i_32794(.A(nbus_157[6]), .Z(n_28776));
	notech_inv i_32796(.A(nbus_157[7]), .Z(n_28777));
	notech_inv i_32797(.A(nbus_157[8]), .Z(n_28778));
	notech_inv i_32798(.A(nbus_157[9]), .Z(n_28779));
	notech_inv i_32799(.A(nbus_157[10]), .Z(n_28780));
	notech_inv i_32800(.A(nbus_157[11]), .Z(n_28781));
	notech_inv i_32801(.A(nbus_157[12]), .Z(n_28783));
	notech_inv i_32802(.A(nbus_157[13]), .Z(n_28784));
	notech_inv i_32803(.A(nbus_157[14]), .Z(n_28785));
	notech_inv i_32804(.A(nbus_157[15]), .Z(n_28786));
	notech_inv i_32805(.A(nbus_157[16]), .Z(n_28787));
	notech_inv i_32806(.A(nbus_157[17]), .Z(n_28788));
	notech_inv i_32807(.A(nbus_157[18]), .Z(n_28789));
	notech_inv i_32808(.A(nbus_157[19]), .Z(n_28790));
	notech_inv i_32809(.A(nbus_157[20]), .Z(n_28791));
	notech_inv i_32810(.A(nbus_157[21]), .Z(n_28792));
	notech_inv i_32811(.A(nbus_157[22]), .Z(n_28793));
	notech_inv i_32812(.A(nbus_157[23]), .Z(n_28794));
	notech_inv i_32813(.A(nbus_157[24]), .Z(n_28795));
	notech_inv i_32814(.A(nbus_157[25]), .Z(n_28796));
	notech_inv i_32815(.A(nbus_157[26]), .Z(n_28797));
	notech_inv i_32816(.A(nbus_157[27]), .Z(n_28798));
	notech_inv i_32817(.A(nbus_157[28]), .Z(n_28799));
	notech_inv i_32818(.A(nbus_157[29]), .Z(n_28800));
	notech_inv i_32819(.A(nbus_157[30]), .Z(n_28801));
	notech_inv i_32820(.A(nbus_157[32]), .Z(n_28802));
	notech_inv i_32821(.A(readio_data[1]), .Z(n_28803));
	notech_inv i_32822(.A(readio_data[2]), .Z(n_28804));
	notech_inv i_32823(.A(readio_data[3]), .Z(n_28805));
	notech_inv i_32824(.A(readio_data[4]), .Z(n_28806));
	notech_inv i_32825(.A(readio_data[6]), .Z(n_28807));
	notech_inv i_32826(.A(readio_data[7]), .Z(n_28808));
	notech_inv i_32827(.A(readio_data[8]), .Z(n_28809));
	notech_inv i_32828(.A(readio_data[9]), .Z(n_28810));
	notech_inv i_32829(.A(readio_data[10]), .Z(n_28811));
	notech_inv i_32830(.A(readio_data[11]), .Z(n_28812));
	notech_inv i_32831(.A(readio_data[12]), .Z(n_28813));
	notech_inv i_32832(.A(readio_data[13]), .Z(n_28814));
	notech_inv i_32834(.A(readio_data[14]), .Z(n_28815));
	notech_inv i_32835(.A(readio_data[15]), .Z(n_28816));
	notech_inv i_32836(.A(readio_data[16]), .Z(n_28817));
	notech_inv i_32837(.A(readio_data[17]), .Z(n_28818));
	notech_inv i_32838(.A(readio_data[18]), .Z(n_28819));
	notech_inv i_32839(.A(readio_data[19]), .Z(n_28820));
	notech_inv i_32840(.A(readio_data[20]), .Z(n_28821));
	notech_inv i_32841(.A(readio_data[21]), .Z(n_28822));
	notech_inv i_32842(.A(readio_data[22]), .Z(n_28823));
	notech_inv i_32843(.A(readio_data[23]), .Z(n_28824));
	notech_inv i_32844(.A(readio_data[24]), .Z(n_28825));
	notech_inv i_32845(.A(readio_data[25]), .Z(n_28826));
	notech_inv i_32846(.A(readio_data[26]), .Z(n_28827));
	notech_inv i_32847(.A(readio_data[27]), .Z(n_28828));
	notech_inv i_32848(.A(readio_data[28]), .Z(n_28829));
	notech_inv i_32849(.A(readio_data[29]), .Z(n_28830));
	notech_inv i_32850(.A(readio_data[30]), .Z(n_28831));
	notech_inv i_32851(.A(readio_data[31]), .Z(n_28832));
	notech_inv i_32852(.A(resa_shiftbox[0]), .Z(n_28833));
	notech_inv i_32853(.A(resa_shiftbox[1]), .Z(n_28834));
	notech_inv i_32854(.A(resa_shiftbox[2]), .Z(n_28835));
	notech_inv i_32855(.A(resa_shiftbox[3]), .Z(n_28836));
	notech_inv i_32856(.A(resa_shiftbox[4]), .Z(n_28837));
	notech_inv i_32857(.A(resa_shiftbox[6]), .Z(n_28838));
	notech_inv i_32858(.A(resa_shiftbox[7]), .Z(n_28839));
	notech_inv i_32859(.A(resa_shiftbox[8]), .Z(n_28840));
	notech_inv i_32860(.A(resa_shiftbox[9]), .Z(n_28842));
	notech_inv i_32861(.A(resa_shiftbox[10]), .Z(n_28844));
	notech_inv i_32862(.A(resa_shiftbox[11]), .Z(n_28845));
	notech_inv i_32863(.A(resa_shiftbox[12]), .Z(n_28846));
	notech_inv i_32864(.A(resa_shiftbox[13]), .Z(n_28847));
	notech_inv i_32865(.A(resa_shiftbox[14]), .Z(n_28849));
	notech_inv i_32866(.A(resa_shiftbox[15]), .Z(n_28850));
	notech_inv i_32867(.A(resa_shiftbox[16]), .Z(n_28852));
	notech_inv i_32868(.A(resa_shiftbox[17]), .Z(n_28854));
	notech_inv i_32869(.A(resa_shiftbox[18]), .Z(n_28855));
	notech_inv i_32870(.A(resa_shiftbox[19]), .Z(n_28856));
	notech_inv i_32871(.A(resa_shiftbox[20]), .Z(n_28858));
	notech_inv i_32872(.A(resa_shiftbox[21]), .Z(n_28859));
	notech_inv i_32873(.A(resa_shiftbox[22]), .Z(n_28861));
	notech_inv i_32874(.A(resa_shiftbox[23]), .Z(n_28863));
	notech_inv i_32875(.A(resa_shiftbox[24]), .Z(n_28867));
	notech_inv i_32876(.A(resa_shiftbox[25]), .Z(n_28872));
	notech_inv i_32877(.A(resa_shiftbox[26]), .Z(n_28873));
	notech_inv i_32878(.A(resa_shiftbox[27]), .Z(n_28874));
	notech_inv i_32879(.A(resa_shiftbox[28]), .Z(n_28875));
	notech_inv i_32880(.A(resa_shiftbox[29]), .Z(n_28876));
	notech_inv i_32881(.A(resa_shiftbox[30]), .Z(n_28877));
	notech_inv i_32882(.A(nbus_162[0]), .Z(n_28878));
	notech_inv i_32883(.A(nbus_162[1]), .Z(n_28879));
	notech_inv i_32884(.A(nbus_162[3]), .Z(n_28880));
	notech_inv i_32885(.A(nbus_162[4]), .Z(n_28881));
	notech_inv i_32886(.A(nbus_162[5]), .Z(n_28882));
	notech_inv i_32887(.A(nbus_162[6]), .Z(n_28883));
	notech_inv i_32888(.A(nbus_162[7]), .Z(n_28884));
	notech_inv i_32889(.A(nbus_162[8]), .Z(n_28885));
	notech_inv i_32890(.A(nbus_162[9]), .Z(n_28886));
	notech_inv i_32891(.A(nbus_162[10]), .Z(n_28887));
	notech_inv i_32892(.A(nbus_162[11]), .Z(n_28888));
	notech_inv i_32893(.A(nbus_162[12]), .Z(n_28889));
	notech_inv i_32894(.A(nbus_162[13]), .Z(n_28890));
	notech_inv i_32895(.A(nbus_162[14]), .Z(n_28891));
	notech_inv i_32896(.A(nbus_162[15]), .Z(n_28892));
	notech_inv i_32897(.A(nbus_162[16]), .Z(n_28893));
	notech_inv i_32898(.A(nbus_162[17]), .Z(n_28894));
	notech_inv i_32899(.A(nbus_162[18]), .Z(n_28895));
	notech_inv i_32900(.A(nbus_162[19]), .Z(n_28896));
	notech_inv i_32901(.A(nbus_162[20]), .Z(n_28897));
	notech_inv i_32902(.A(nbus_162[21]), .Z(n_28898));
	notech_inv i_32903(.A(nbus_162[22]), .Z(n_28899));
	notech_inv i_32904(.A(nbus_162[23]), .Z(n_28900));
	notech_inv i_32905(.A(nbus_162[24]), .Z(n_28901));
	notech_inv i_32906(.A(nbus_162[25]), .Z(n_28902));
	notech_inv i_32907(.A(nbus_162[26]), .Z(n_28903));
	notech_inv i_32908(.A(nbus_162[27]), .Z(n_28904));
	notech_inv i_32909(.A(nbus_162[28]), .Z(n_28905));
	notech_inv i_32910(.A(nbus_162[29]), .Z(n_28906));
	notech_inv i_32912(.A(nbus_162[30]), .Z(n_28907));
	notech_inv i_32913(.A(nbus_162[31]), .Z(n_28908));
	notech_inv i_32914(.A(nbus_164[0]), .Z(n_28909));
	notech_inv i_32915(.A(nbus_164[1]), .Z(n_28910));
	notech_inv i_32916(.A(nbus_164[2]), .Z(n_28911));
	notech_inv i_32917(.A(nbus_164[3]), .Z(n_28912));
	notech_inv i_32918(.A(nbus_164[4]), .Z(n_28913));
	notech_inv i_32919(.A(nbus_164[5]), .Z(n_28914));
	notech_inv i_32920(.A(nbus_164[6]), .Z(n_28915));
	notech_inv i_32921(.A(nbus_164[7]), .Z(n_28916));
	notech_inv i_32922(.A(nbus_164[8]), .Z(n_28917));
	notech_inv i_32923(.A(nbus_164[9]), .Z(n_28918));
	notech_inv i_32924(.A(nbus_164[10]), .Z(n_28919));
	notech_inv i_32925(.A(nbus_164[11]), .Z(n_28920));
	notech_inv i_32926(.A(nbus_164[12]), .Z(n_28921));
	notech_inv i_32928(.A(nbus_164[13]), .Z(n_28922));
	notech_inv i_32929(.A(nbus_164[14]), .Z(n_28923));
	notech_inv i_32930(.A(nbus_164[15]), .Z(n_28924));
	notech_inv i_32931(.A(nbus_164[32]), .Z(n_28925));
	notech_inv i_32932(.A(nbus_167[0]), .Z(n_28926));
	notech_inv i_32933(.A(nbus_167[1]), .Z(n_28927));
	notech_inv i_32934(.A(nbus_167[2]), .Z(n_28928));
	notech_inv i_32935(.A(nbus_167[3]), .Z(n_28929));
	notech_inv i_32936(.A(nbus_167[4]), .Z(n_28930));
	notech_inv i_32937(.A(nbus_167[5]), .Z(n_28931));
	notech_inv i_32938(.A(nbus_167[6]), .Z(n_28932));
	notech_inv i_32939(.A(nbus_167[7]), .Z(n_28933));
	notech_inv i_32940(.A(nbus_167[8]), .Z(n_28934));
	notech_inv i_32941(.A(nbus_167[9]), .Z(n_28935));
	notech_inv i_32942(.A(nbus_167[10]), .Z(n_28936));
	notech_inv i_32943(.A(nbus_167[11]), .Z(n_28937));
	notech_inv i_32944(.A(nbus_167[12]), .Z(n_28938));
	notech_inv i_32945(.A(nbus_167[13]), .Z(n_28939));
	notech_inv i_32946(.A(nbus_167[14]), .Z(n_28940));
	notech_inv i_32947(.A(nbus_167[15]), .Z(n_28941));
	notech_inv i_32948(.A(nbus_167[16]), .Z(n_28942));
	notech_inv i_32949(.A(tsc[0]), .Z(n_28943));
	notech_inv i_32950(.A(tsc[1]), .Z(n_28944));
	notech_inv i_32951(.A(tsc[2]), .Z(n_28945));
	notech_inv i_32952(.A(tsc[3]), .Z(n_28946));
	notech_inv i_32953(.A(tsc[4]), .Z(n_28947));
	notech_inv i_32954(.A(tsc[5]), .Z(n_28948));
	notech_inv i_32955(.A(tsc[6]), .Z(n_28949));
	notech_inv i_32956(.A(tsc[8]), .Z(n_28950));
	notech_inv i_32957(.A(tsc[9]), .Z(n_28951));
	notech_inv i_32958(.A(tsc[12]), .Z(n_28952));
	notech_inv i_32959(.A(tsc[16]), .Z(n_28953));
	notech_inv i_32960(.A(tsc[17]), .Z(n_28954));
	notech_inv i_32961(.A(tsc[18]), .Z(n_28955));
	notech_inv i_32962(.A(tsc[19]), .Z(n_28956));
	notech_inv i_32963(.A(tsc[21]), .Z(n_28957));
	notech_inv i_32964(.A(tsc[26]), .Z(n_28958));
	notech_inv i_32965(.A(tsc[28]), .Z(n_28959));
	notech_inv i_32966(.A(tsc[29]), .Z(n_28960));
	notech_inv i_32967(.A(tsc[32]), .Z(n_28961));
	notech_inv i_32968(.A(tsc[33]), .Z(n_28962));
	notech_inv i_32969(.A(tsc[34]), .Z(n_28964));
	notech_inv i_32970(.A(tsc[35]), .Z(n_28965));
	notech_inv i_32971(.A(tsc[37]), .Z(n_28966));
	notech_inv i_32972(.A(tsc[39]), .Z(n_28967));
	notech_inv i_32973(.A(tsc[40]), .Z(n_28968));
	notech_inv i_32974(.A(tsc[48]), .Z(n_28970));
	notech_inv i_32975(.A(tsc[49]), .Z(n_28971));
	notech_inv i_32976(.A(tsc[50]), .Z(n_28972));
	notech_inv i_32977(.A(tsc[51]), .Z(n_28974));
	notech_inv i_32978(.A(tsc[52]), .Z(n_28976));
	notech_inv i_32979(.A(tsc[53]), .Z(n_28977));
	notech_inv i_32980(.A(tsc[55]), .Z(n_28978));
	notech_inv i_32981(.A(tsc[57]), .Z(n_28979));
	notech_inv i_32982(.A(tsc[58]), .Z(n_28980));
	notech_inv i_32983(.A(tsc[59]), .Z(n_28982));
	notech_inv i_32984(.A(tsc[60]), .Z(n_28983));
	notech_inv i_32985(.A(tsc[61]), .Z(n_28984));
	notech_inv i_32986(.A(nbus_161[0]), .Z(n_28985));
	notech_inv i_32987(.A(nbus_161[1]), .Z(n_28986));
	notech_inv i_32988(.A(nbus_161[2]), .Z(n_28989));
	notech_inv i_32989(.A(nbus_161[3]), .Z(n_28990));
	notech_inv i_32990(.A(nbus_161[4]), .Z(n_28991));
	notech_inv i_32991(.A(nbus_161[5]), .Z(n_28992));
	notech_inv i_32992(.A(nbus_161[6]), .Z(n_28993));
	notech_inv i_32993(.A(nbus_161[7]), .Z(n_28994));
	notech_inv i_32994(.A(nbus_161[8]), .Z(n_28995));
	notech_inv i_32995(.A(nbus_161[9]), .Z(n_28996));
	notech_inv i_32996(.A(nbus_161[10]), .Z(n_28997));
	notech_inv i_32997(.A(nbus_161[11]), .Z(n_28998));
	notech_inv i_32998(.A(nbus_161[12]), .Z(n_28999));
	notech_inv i_32999(.A(nbus_161[13]), .Z(n_29000));
	notech_inv i_33000(.A(nbus_161[14]), .Z(n_29001));
	notech_inv i_33001(.A(nbus_161[15]), .Z(n_29002));
	notech_inv i_33002(.A(mul64[0]), .Z(n_29003));
	notech_inv i_33003(.A(mul64[1]), .Z(n_29004));
	notech_inv i_33004(.A(mul64[2]), .Z(n_29005));
	notech_inv i_33005(.A(mul64[3]), .Z(n_29006));
	notech_inv i_33006(.A(mul64[4]), .Z(n_29007));
	notech_inv i_33007(.A(mul64[6]), .Z(n_29008));
	notech_inv i_33008(.A(mul64[7]), .Z(n_29009));
	notech_inv i_33009(.A(imm[34]), .Z(n_29010));
	notech_inv i_33010(.A(imm[3]), .Z(n_29011));
	notech_inv i_33011(.A(imm[21]), .Z(n_29012));
	notech_inv i_33012(.A(imm[44]), .Z(n_29013));
	notech_inv i_33013(.A(imm[12]), .Z(n_29014));
	notech_inv i_33014(.A(imm[25]), .Z(n_29015));
	notech_inv i_33015(.A(imm[4]), .Z(n_29016));
	notech_inv i_33017(.A(imm[5]), .Z(n_29017));
	notech_inv i_33018(.A(imm[17]), .Z(n_29018));
	notech_inv i_33020(.A(imm[19]), .Z(n_29019));
	notech_inv i_33021(.A(imm[20]), .Z(n_29020));
	notech_inv i_33022(.A(imm[6]), .Z(n_29021));
	notech_inv i_33023(.A(imm[7]), .Z(n_29022));
	notech_inv i_33024(.A(imm[8]), .Z(n_29023));
	notech_inv i_33025(.A(imm[9]), .Z(n_29024));
	notech_inv i_33026(.A(imm[11]), .Z(n_29025));
	notech_inv i_33027(.A(imm[13]), .Z(n_29026));
	notech_inv i_33028(.A(imm[14]), .Z(n_29027));
	notech_inv i_33029(.A(imm[15]), .Z(n_29028));
	notech_inv i_33030(.A(imm[22]), .Z(n_29029));
	notech_inv i_33031(.A(imm[31]), .Z(n_29030));
	notech_inv i_33032(.A(imm[30]), .Z(n_29031));
	notech_inv i_33033(.A(imm[26]), .Z(n_29032));
	notech_inv i_33034(.A(imm[10]), .Z(n_29033));
	notech_inv i_33035(.A(imm[27]), .Z(n_29034));
	notech_inv i_33036(.A(imm[32]), .Z(n_29035));
	notech_inv i_33037(.A(imm[33]), .Z(n_29036));
	notech_inv i_33038(.A(imm[35]), .Z(n_29037));
	notech_inv i_33042(.A(imm[36]), .Z(n_29038));
	notech_inv i_33046(.A(imm[40]), .Z(n_29039));
	notech_inv i_33047(.A(imm[41]), .Z(n_29040));
	notech_inv i_33048(.A(imm[42]), .Z(n_29041));
	notech_inv i_33050(.A(imm[43]), .Z(n_29042));
	notech_inv i_33051(.A(imm[45]), .Z(n_29043));
	notech_inv i_33053(.A(imm[46]), .Z(n_29044));
	notech_inv i_33054(.A(imm[47]), .Z(n_29045));
	notech_inv i_33055(.A(imm[18]), .Z(n_29046));
	notech_inv i_33057(.A(imm[16]), .Z(n_29047));
	notech_inv i_33059(.A(imm[23]), .Z(n_29048));
	notech_inv i_33060(.A(imm[24]), .Z(n_29049));
	notech_inv i_33062(.A(imm[28]), .Z(n_29050));
	notech_inv i_33063(.A(imm[29]), .Z(n_29051));
	notech_inv i_33064(.A(add_src[0]), .Z(n_29052));
	notech_inv i_33065(.A(add_src[1]), .Z(n_29053));
	notech_inv i_33067(.A(add_src[2]), .Z(n_29054));
	notech_inv i_33069(.A(add_src[5]), .Z(n_29055));
	notech_inv i_33070(.A(add_src[6]), .Z(n_29056));
	notech_inv i_33071(.A(add_src[7]), .Z(n_29060));
	notech_inv i_33072(.A(add_src[8]), .Z(n_29061));
	notech_inv i_33073(.A(add_src[9]), .Z(n_29062));
	notech_inv i_33074(.A(add_src[11]), .Z(n_29063));
	notech_inv i_33075(.A(add_src[12]), .Z(n_29064));
	notech_inv i_33076(.A(add_src[13]), .Z(n_29065));
	notech_inv i_33077(.A(add_src[14]), .Z(n_29066));
	notech_inv i_33078(.A(add_src[15]), .Z(n_29067));
	notech_inv i_33079(.A(add_src[16]), .Z(n_29069));
	notech_inv i_33080(.A(add_src[17]), .Z(n_29070));
	notech_inv i_33081(.A(add_src[18]), .Z(n_29072));
	notech_inv i_33082(.A(add_src[19]), .Z(n_29073));
	notech_inv i_33083(.A(add_src[20]), .Z(n_29074));
	notech_inv i_33084(.A(add_src[21]), .Z(n_29075));
	notech_inv i_33085(.A(add_src[22]), .Z(n_29076));
	notech_inv i_33086(.A(add_src[23]), .Z(n_29077));
	notech_inv i_33087(.A(add_src[24]), .Z(n_29078));
	notech_inv i_33088(.A(add_src[25]), .Z(n_29079));
	notech_inv i_33089(.A(add_src[26]), .Z(n_29080));
	notech_inv i_33090(.A(add_src[27]), .Z(n_29081));
	notech_inv i_33091(.A(add_src[28]), .Z(n_29082));
	notech_inv i_33092(.A(add_src[29]), .Z(n_29083));
	notech_inv i_33093(.A(add_src[30]), .Z(n_29084));
	notech_inv i_33094(.A(add_src[31]), .Z(n_29085));
	notech_inv i_33095(.A(nbus_166[0]), .Z(n_29086));
	notech_inv i_33096(.A(nbus_166[1]), .Z(n_29087));
	notech_inv i_33097(.A(nbus_166[2]), .Z(n_29088));
	notech_inv i_33098(.A(nbus_166[3]), .Z(n_29089));
	notech_inv i_33099(.A(nbus_166[4]), .Z(n_29090));
	notech_inv i_33100(.A(nbus_166[5]), .Z(n_29091));
	notech_inv i_33101(.A(nbus_166[6]), .Z(n_29092));
	notech_inv i_33102(.A(nbus_166[7]), .Z(n_29093));
	notech_inv i_33103(.A(nbus_166[8]), .Z(n_29094));
	notech_inv i_33104(.A(nbus_166[9]), .Z(n_29095));
	notech_inv i_33105(.A(nbus_166[10]), .Z(n_29096));
	notech_inv i_33106(.A(nbus_166[11]), .Z(n_29097));
	notech_inv i_33107(.A(nbus_166[12]), .Z(n_29098));
	notech_inv i_33108(.A(nbus_166[13]), .Z(n_29099));
	notech_inv i_33109(.A(nbus_166[14]), .Z(n_29100));
	notech_inv i_33110(.A(nbus_166[15]), .Z(n_29101));
	notech_inv i_33111(.A(nbus_166[16]), .Z(n_29102));
	notech_inv i_33112(.A(nbus_166[17]), .Z(n_29103));
	notech_inv i_33113(.A(nbus_166[18]), .Z(n_29104));
	notech_inv i_33114(.A(nbus_166[19]), .Z(n_29105));
	notech_inv i_33115(.A(nbus_166[20]), .Z(n_29106));
	notech_inv i_33116(.A(nbus_166[21]), .Z(n_29107));
	notech_inv i_33117(.A(nbus_166[22]), .Z(n_29108));
	notech_inv i_33118(.A(nbus_166[23]), .Z(n_29109));
	notech_inv i_33119(.A(nbus_166[24]), .Z(n_29110));
	notech_inv i_33120(.A(nbus_166[25]), .Z(n_29111));
	notech_inv i_33121(.A(nbus_166[26]), .Z(n_29112));
	notech_inv i_33122(.A(nbus_166[28]), .Z(n_29113));
	notech_inv i_33123(.A(nbus_166[29]), .Z(n_29114));
	notech_inv i_33124(.A(nbus_166[30]), .Z(n_29115));
	notech_inv i_33125(.A(nbus_166[32]), .Z(n_29116));
	notech_inv i_33126(.A(instrc[0]), .Z(n_29117));
	notech_inv i_33127(.A(instrc[8]), .Z(n_29118));
	notech_inv i_33128(.A(instrc[9]), .Z(n_29119));
	notech_inv i_33129(.A(instrc[10]), .Z(n_29120));
	notech_inv i_33130(.A(instrc[11]), .Z(n_29121));
	notech_inv i_33131(.A(instrc[12]), .Z(n_29122));
	notech_inv i_33132(.A(instrc[13]), .Z(n_29123));
	notech_inv i_33133(.A(instrc[14]), .Z(n_29124));
	notech_inv i_33134(.A(instrc[15]), .Z(n_29125));
	notech_inv i_33135(.A(instrc[16]), .Z(n_29127));
	notech_inv i_33136(.A(instrc[17]), .Z(n_29128));
	notech_inv i_33137(.A(instrc[18]), .Z(n_29129));
	notech_inv i_33138(.A(instrc[19]), .Z(n_29130));
	notech_inv i_33139(.A(instrc[20]), .Z(n_29131));
	notech_inv i_33140(.A(instrc[21]), .Z(n_29132));
	notech_inv i_33141(.A(instrc[22]), .Z(n_29133));
	notech_inv i_33142(.A(instrc[23]), .Z(n_29134));
	notech_inv i_33143(.A(instrc[24]), .Z(n_29135));
	notech_inv i_33144(.A(instrc[25]), .Z(n_29136));
	notech_inv i_33145(.A(instrc[26]), .Z(n_29137));
	notech_inv i_33146(.A(instrc[27]), .Z(n_29138));
	notech_inv i_33147(.A(instrc[28]), .Z(n_29139));
	notech_inv i_33148(.A(instrc[29]), .Z(n_29140));
	notech_inv i_33149(.A(instrc[30]), .Z(n_29141));
	notech_inv i_33150(.A(instrc[31]), .Z(n_29142));
	notech_inv i_33151(.A(instrc[32]), .Z(n_29143));
	notech_inv i_33152(.A(instrc[33]), .Z(n_29144));
	notech_inv i_33153(.A(instrc[34]), .Z(n_29145));
	notech_inv i_33154(.A(instrc[35]), .Z(n_29146));
	notech_inv i_33155(.A(instrc[36]), .Z(n_29147));
	notech_inv i_33156(.A(instrc[37]), .Z(n_29148));
	notech_inv i_33157(.A(instrc[38]), .Z(n_29149));
	notech_inv i_33158(.A(instrc[39]), .Z(n_29150));
	notech_inv i_33159(.A(instrc[40]), .Z(n_29151));
	notech_inv i_33160(.A(instrc[41]), .Z(n_29152));
	notech_inv i_33161(.A(instrc[42]), .Z(n_29153));
	notech_inv i_33162(.A(instrc[43]), .Z(n_29154));
	notech_inv i_33163(.A(instrc[44]), .Z(n_29155));
	notech_inv i_33164(.A(instrc[45]), .Z(n_29156));
	notech_inv i_33165(.A(instrc[46]), .Z(n_29157));
	notech_inv i_33166(.A(instrc[47]), .Z(n_29158));
	notech_inv i_33167(.A(instrc[48]), .Z(n_29159));
	notech_inv i_33168(.A(instrc[49]), .Z(n_29160));
	notech_inv i_33169(.A(instrc[50]), .Z(n_29161));
	notech_inv i_33170(.A(instrc[51]), .Z(n_29162));
	notech_inv i_33171(.A(instrc[52]), .Z(n_29163));
	notech_inv i_33172(.A(instrc[53]), .Z(n_29164));
	notech_inv i_33173(.A(instrc[54]), .Z(n_29165));
	notech_inv i_33174(.A(instrc[55]), .Z(n_29166));
	notech_inv i_33175(.A(instrc[72]), .Z(n_29167));
	notech_inv i_33177(.A(instrc[73]), .Z(n_29168));
	notech_inv i_33178(.A(instrc[74]), .Z(n_29169));
	notech_inv i_33180(.A(instrc[75]), .Z(n_29170));
	notech_inv i_33181(.A(instrc[76]), .Z(n_29171));
	notech_inv i_33182(.A(instrc[77]), .Z(n_29172));
	notech_inv i_33183(.A(instrc[78]), .Z(n_29173));
	notech_inv i_33184(.A(instrc[79]), .Z(n_29174));
	notech_inv i_33185(.A(instrc[108]), .Z(n_29175));
	notech_inv i_33186(.A(instrc[109]), .Z(n_29176));
	notech_inv i_33190(.A(n_59397), .Z(n_29177));
	notech_inv i_33191(.A(n_59373), .Z(n_29178));
	notech_inv i_33192(.A(n_60915), .Z(n_29179));
	notech_inv i_33193(.A(instrc[123]), .Z(n_29180));
	notech_inv i_33194(.A(nbus_160[3]), .Z(n_29181));
	notech_inv i_33195(.A(nbus_160[4]), .Z(n_29182));
	notech_inv i_33196(.A(nbus_160[5]), .Z(n_29183));
	notech_inv i_33197(.A(nbus_160[6]), .Z(n_29184));
	notech_inv i_33198(.A(nbus_160[7]), .Z(n_29185));
	notech_inv i_33199(.A(nbus_160[8]), .Z(n_29186));
	notech_inv i_33200(.A(nbus_160[9]), .Z(n_29187));
	notech_inv i_33201(.A(nbus_160[10]), .Z(n_29188));
	notech_inv i_33202(.A(nbus_160[11]), .Z(n_29189));
	notech_inv i_33203(.A(nbus_160[12]), .Z(n_29190));
	notech_inv i_33204(.A(nbus_160[13]), .Z(n_29191));
	notech_inv i_33205(.A(nbus_160[14]), .Z(n_29192));
	notech_inv i_33206(.A(nbus_160[15]), .Z(n_29194));
	notech_inv i_33207(.A(nbus_160[16]), .Z(n_29195));
	notech_inv i_33208(.A(nbus_160[17]), .Z(n_29197));
	notech_inv i_33209(.A(nbus_160[18]), .Z(n_29198));
	notech_inv i_33210(.A(nbus_160[19]), .Z(n_29199));
	notech_inv i_33211(.A(nbus_160[20]), .Z(n_29200));
	notech_inv i_33212(.A(nbus_160[21]), .Z(n_29202));
	notech_inv i_33213(.A(nbus_160[22]), .Z(n_29203));
	notech_inv i_33214(.A(nbus_160[23]), .Z(n_29205));
	notech_inv i_33215(.A(nbus_160[24]), .Z(n_29206));
	notech_inv i_33216(.A(nbus_160[25]), .Z(n_29208));
	notech_inv i_33217(.A(nbus_160[26]), .Z(n_29210));
	notech_inv i_33218(.A(nbus_160[27]), .Z(n_29211));
	notech_inv i_33219(.A(nbus_160[28]), .Z(n_29213));
	notech_inv i_33220(.A(nbus_160[29]), .Z(n_29214));
	notech_inv i_33221(.A(nbus_160[30]), .Z(n_29216));
	notech_inv i_33222(.A(nbus_160[31]), .Z(n_29217));
	notech_inv i_33223(.A(resb_shiftbox[8]), .Z(n_29218));
	notech_inv i_33224(.A(resb_shiftbox[9]), .Z(n_29222));
	notech_inv i_33225(.A(resb_shiftbox[10]), .Z(n_29226));
	notech_inv i_33226(.A(resb_shiftbox[11]), .Z(n_29227));
	notech_inv i_33227(.A(resb_shiftbox[12]), .Z(n_29228));
	notech_inv i_33228(.A(resb_shiftbox[13]), .Z(n_29229));
	notech_inv i_33229(.A(resb_shiftbox[14]), .Z(n_29231));
	notech_inv i_33230(.A(resb_shiftbox[15]), .Z(n_29232));
	notech_inv i_33231(.A(resb_shiftbox[16]), .Z(n_29233));
	notech_inv i_33232(.A(resb_shiftbox[17]), .Z(n_29234));
	notech_inv i_33233(.A(resb_shiftbox[18]), .Z(n_29235));
	notech_inv i_33234(.A(resb_shiftbox[19]), .Z(n_29236));
	notech_inv i_33235(.A(resb_shiftbox[20]), .Z(n_29237));
	notech_inv i_33236(.A(resb_shiftbox[21]), .Z(n_29238));
	notech_inv i_33237(.A(resb_shiftbox[22]), .Z(n_29239));
	notech_inv i_33238(.A(resb_shiftbox[23]), .Z(n_29241));
	notech_inv i_33239(.A(resb_shiftbox[24]), .Z(n_29242));
	notech_inv i_33240(.A(resb_shiftbox[25]), .Z(n_29243));
	notech_inv i_33241(.A(resb_shiftbox[26]), .Z(n_29244));
	notech_inv i_33242(.A(resb_shiftbox[27]), .Z(n_29245));
	notech_inv i_33243(.A(resb_shiftbox[28]), .Z(n_29246));
	notech_inv i_33244(.A(resb_shiftbox[29]), .Z(n_29247));
	notech_inv i_33245(.A(resb_shiftbox[30]), .Z(n_29248));
	notech_inv i_33246(.A(resb_shiftbox[31]), .Z(n_29249));
	notech_inv i_33247(.A(resb_shift4box[0]), .Z(n_29250));
	notech_inv i_33248(.A(resb_shift4box[1]), .Z(n_29251));
	notech_inv i_33249(.A(resb_shift4box[2]), .Z(n_29252));
	notech_inv i_33250(.A(resb_shift4box[3]), .Z(n_29253));
	notech_inv i_33251(.A(resb_shift4box[4]), .Z(n_29254));
	notech_inv i_33252(.A(resb_shift4box[8]), .Z(n_29255));
	notech_inv i_33253(.A(resb_shift4box[9]), .Z(n_29258));
	notech_inv i_33254(.A(resb_shift4box[10]), .Z(n_29261));
	notech_inv i_33255(.A(resb_shift4box[11]), .Z(n_29263));
	notech_inv i_33256(.A(resb_shift4box[12]), .Z(n_29264));
	notech_inv i_33257(.A(resb_shift4box[13]), .Z(n_29265));
	notech_inv i_33258(.A(resb_shift4box[14]), .Z(n_29266));
	notech_inv i_33259(.A(resb_shift4box[15]), .Z(n_29267));
	notech_inv i_33260(.A(resb_shift4box[16]), .Z(n_29268));
	notech_inv i_33262(.A(resb_shift4box[17]), .Z(n_29269));
	notech_inv i_33263(.A(resb_shift4box[18]), .Z(n_29270));
	notech_inv i_33264(.A(resb_shift4box[19]), .Z(n_29271));
	notech_inv i_33265(.A(resb_shift4box[20]), .Z(n_29272));
	notech_inv i_33267(.A(resb_shift4box[21]), .Z(n_29273));
	notech_inv i_33268(.A(resb_shift4box[22]), .Z(n_29274));
	notech_inv i_33269(.A(resb_shift4box[23]), .Z(n_29275));
	notech_inv i_33270(.A(resb_shift4box[24]), .Z(n_29276));
	notech_inv i_33271(.A(resb_shift4box[25]), .Z(n_29277));
	notech_inv i_33272(.A(resb_shift4box[26]), .Z(n_29278));
	notech_inv i_33273(.A(resb_shift4box[27]), .Z(n_29279));
	notech_inv i_33274(.A(resb_shift4box[28]), .Z(n_29280));
	notech_inv i_33275(.A(resb_shift4box[29]), .Z(n_29281));
	notech_inv i_33276(.A(resb_shift4box[30]), .Z(n_29283));
	notech_inv i_33277(.A(resb_shift4box[31]), .Z(n_29284));
	notech_inv i_33278(.A(Daddrs_8[0]), .Z(n_29285));
	notech_inv i_33279(.A(Daddrs_8[2]), .Z(n_29286));
	notech_inv i_33280(.A(Daddrs_8[3]), .Z(n_29287));
	notech_inv i_33281(.A(Daddrs_8[4]), .Z(n_29288));
	notech_inv i_33282(.A(Daddrs_8[5]), .Z(n_29289));
	notech_inv i_33283(.A(Daddrs_8[6]), .Z(n_29290));
	notech_inv i_33284(.A(Daddrs_8[7]), .Z(n_29291));
	notech_inv i_33285(.A(Daddrs_8[8]), .Z(n_29292));
	notech_inv i_33286(.A(Daddrs_8[9]), .Z(n_29293));
	notech_inv i_33287(.A(Daddrs_8[10]), .Z(n_29294));
	notech_inv i_33288(.A(Daddrs_8[11]), .Z(n_29295));
	notech_inv i_33289(.A(Daddrs_8[12]), .Z(n_29296));
	notech_inv i_33290(.A(Daddrs_8[13]), .Z(n_29297));
	notech_inv i_33291(.A(Daddrs_8[14]), .Z(n_29298));
	notech_inv i_33292(.A(Daddrs_8[15]), .Z(n_29299));
	notech_inv i_33293(.A(Daddrs_8[16]), .Z(n_29300));
	notech_inv i_33294(.A(Daddrs_8[17]), .Z(n_29301));
	notech_inv i_33295(.A(Daddrs_8[18]), .Z(n_29302));
	notech_inv i_33296(.A(Daddrs_8[19]), .Z(n_29303));
	notech_inv i_33297(.A(Daddrs_8[20]), .Z(n_29304));
	notech_inv i_33298(.A(Daddrs_8[21]), .Z(n_29305));
	notech_inv i_33299(.A(Daddrs_8[22]), .Z(n_29306));
	notech_inv i_33300(.A(Daddrs_8[23]), .Z(n_29307));
	notech_inv i_33301(.A(Daddrs_8[24]), .Z(n_29308));
	notech_inv i_33302(.A(Daddrs_8[25]), .Z(n_29309));
	notech_inv i_33303(.A(Daddrs_8[26]), .Z(n_29310));
	notech_inv i_33304(.A(Daddrs_8[27]), .Z(n_29311));
	notech_inv i_33305(.A(Daddrs_8[28]), .Z(n_29312));
	notech_inv i_33306(.A(Daddrs_8[29]), .Z(n_29313));
	notech_inv i_33307(.A(Daddrs_8[30]), .Z(n_29314));
	notech_inv i_33308(.A(Daddrs_8[31]), .Z(n_29315));
	notech_inv i_33309(.A(Daddrs_3[0]), .Z(n_29316));
	notech_inv i_33310(.A(Daddrs_3[1]), .Z(n_29317));
	notech_inv i_33311(.A(Daddrs_3[2]), .Z(n_29318));
	notech_inv i_33312(.A(Daddrs_3[3]), .Z(n_29319));
	notech_inv i_33313(.A(Daddrs_3[4]), .Z(n_29320));
	notech_inv i_33314(.A(Daddrs_3[5]), .Z(n_29321));
	notech_inv i_33315(.A(Daddrs_3[6]), .Z(n_29322));
	notech_inv i_33316(.A(Daddrs_3[7]), .Z(n_29323));
	notech_inv i_33317(.A(Daddrs_3[8]), .Z(n_29324));
	notech_inv i_33318(.A(Daddrs_3[9]), .Z(n_29325));
	notech_inv i_33319(.A(Daddrs_3[10]), .Z(n_29326));
	notech_inv i_33320(.A(Daddrs_3[12]), .Z(n_29327));
	notech_inv i_33321(.A(Daddrs_3[13]), .Z(n_29328));
	notech_inv i_33322(.A(Daddrs_3[14]), .Z(n_29329));
	notech_inv i_33323(.A(Daddrs_3[15]), .Z(n_29330));
	notech_inv i_33324(.A(Daddrs_3[16]), .Z(n_29331));
	notech_inv i_33325(.A(Daddrs_3[17]), .Z(n_29332));
	notech_inv i_33326(.A(Daddrs_3[18]), .Z(n_29333));
	notech_inv i_33327(.A(Daddrs_3[19]), .Z(n_29334));
	notech_inv i_33328(.A(Daddrs_3[20]), .Z(n_29335));
	notech_inv i_33329(.A(Daddrs_3[21]), .Z(n_29336));
	notech_inv i_33330(.A(Daddrs_3[22]), .Z(n_29337));
	notech_inv i_33331(.A(Daddrs_3[23]), .Z(n_29338));
	notech_inv i_33332(.A(Daddrs_3[24]), .Z(n_29339));
	notech_inv i_33333(.A(Daddrs_3[25]), .Z(n_29340));
	notech_inv i_33334(.A(Daddrs_3[26]), .Z(n_29341));
	notech_inv i_33335(.A(Daddrs_3[27]), .Z(n_29342));
	notech_inv i_33337(.A(Daddrs_3[28]), .Z(n_29343));
	notech_inv i_33338(.A(Daddrs_3[29]), .Z(n_29344));
	notech_inv i_33339(.A(Daddrs_3[30]), .Z(n_29345));
	notech_inv i_33340(.A(Daddrs_3[31]), .Z(n_29346));
	notech_inv i_33341(.A(Daddrs_1[0]), .Z(n_29347));
	notech_inv i_33342(.A(Daddrs_1[2]), .Z(n_29348));
	notech_inv i_33343(.A(Daddrs_1[3]), .Z(n_29349));
	notech_inv i_33344(.A(Daddrs_1[4]), .Z(n_29350));
	notech_inv i_33345(.A(Daddrs_1[5]), .Z(n_29351));
	notech_inv i_33346(.A(Daddrs_1[6]), .Z(n_29352));
	notech_inv i_33347(.A(Daddrs_1[7]), .Z(n_29353));
	notech_inv i_33348(.A(Daddrs_1[8]), .Z(n_29354));
	notech_inv i_33349(.A(Daddrs_1[9]), .Z(n_29355));
	notech_inv i_33350(.A(Daddrs_1[10]), .Z(n_29356));
	notech_inv i_33351(.A(Daddrs_1[11]), .Z(n_29357));
	notech_inv i_33352(.A(Daddrs_1[12]), .Z(n_29358));
	notech_inv i_33353(.A(Daddrs_1[13]), .Z(n_29359));
	notech_inv i_33354(.A(Daddrs_1[14]), .Z(n_29360));
	notech_inv i_33355(.A(Daddrs_1[15]), .Z(n_29361));
	notech_inv i_33356(.A(Daddrs_1[16]), .Z(n_29362));
	notech_inv i_33357(.A(Daddrs_1[17]), .Z(n_29363));
	notech_inv i_33358(.A(Daddrs_1[18]), .Z(n_29364));
	notech_inv i_33359(.A(Daddrs_1[19]), .Z(n_29365));
	notech_inv i_33360(.A(Daddrs_1[20]), .Z(n_29366));
	notech_inv i_33361(.A(Daddrs_1[21]), .Z(n_29367));
	notech_inv i_33362(.A(Daddrs_1[22]), .Z(n_29368));
	notech_inv i_33363(.A(Daddrs_1[23]), .Z(n_29369));
	notech_inv i_33364(.A(Daddrs_1[24]), .Z(n_29370));
	notech_inv i_33365(.A(Daddrs_1[25]), .Z(n_29371));
	notech_inv i_33366(.A(Daddrs_1[26]), .Z(n_29372));
	notech_inv i_33367(.A(Daddrs_1[27]), .Z(n_29373));
	notech_inv i_33368(.A(Daddrs_1[28]), .Z(n_29374));
	notech_inv i_33369(.A(Daddrs_1[29]), .Z(n_29375));
	notech_inv i_33370(.A(Daddrs_1[30]), .Z(n_29376));
	notech_inv i_33371(.A(Daddrs_1[31]), .Z(n_29377));
	notech_inv i_33372(.A(opc_14[0]), .Z(n_29378));
	notech_inv i_33373(.A(opc_14[1]), .Z(n_29379));
	notech_inv i_33374(.A(opc_14[2]), .Z(n_29380));
	notech_inv i_33375(.A(opc_14[3]), .Z(n_29381));
	notech_inv i_33376(.A(opc_14[4]), .Z(n_29382));
	notech_inv i_33377(.A(opc_14[5]), .Z(n_29383));
	notech_inv i_33378(.A(opc_14[6]), .Z(n_29384));
	notech_inv i_33380(.A(opc_14[7]), .Z(n_29385));
	notech_inv i_33381(.A(opc_14[8]), .Z(n_29386));
	notech_inv i_33382(.A(opc_14[9]), .Z(n_29387));
	notech_inv i_33383(.A(opc_14[10]), .Z(n_29388));
	notech_inv i_33384(.A(opc_14[11]), .Z(n_29389));
	notech_inv i_33385(.A(opc_14[12]), .Z(n_29390));
	notech_inv i_33386(.A(opc_14[13]), .Z(n_29391));
	notech_inv i_33387(.A(opc_14[14]), .Z(n_29392));
	notech_inv i_33388(.A(opc_14[15]), .Z(n_29393));
	notech_inv i_33389(.A(opc_14[16]), .Z(n_29394));
	notech_inv i_33390(.A(opc_14[17]), .Z(n_29395));
	notech_inv i_33391(.A(opc_14[18]), .Z(n_29396));
	notech_inv i_33392(.A(opc_14[19]), .Z(n_29397));
	notech_inv i_33393(.A(opc_14[20]), .Z(n_29398));
	notech_inv i_33394(.A(opc_14[21]), .Z(n_29399));
	notech_inv i_33395(.A(opc_14[22]), .Z(n_29400));
	notech_inv i_33396(.A(opc_14[23]), .Z(n_29401));
	notech_inv i_33398(.A(opc_14[24]), .Z(n_29402));
	notech_inv i_33399(.A(from_acu[0]), .Z(n_29403));
	notech_inv i_33400(.A(from_acu[1]), .Z(n_29404));
	notech_inv i_33401(.A(from_acu[2]), .Z(n_29405));
	notech_inv i_33402(.A(from_acu[3]), .Z(n_29406));
	notech_inv i_33403(.A(from_acu[4]), .Z(n_29407));
	notech_inv i_33404(.A(from_acu[5]), .Z(n_29408));
	notech_inv i_33405(.A(from_acu[6]), .Z(n_29409));
	notech_inv i_33406(.A(to_acu100236[0]), .Z(to_acu[0]));
	notech_inv i_33407(.A(to_acu100236[1]), .Z(to_acu[1]));
	notech_inv i_33408(.A(to_acu100236[2]), .Z(to_acu[2]));
	notech_inv i_33409(.A(to_acu100236[3]), .Z(to_acu[3]));
	notech_inv i_33410(.A(to_acu100236[4]), .Z(to_acu[4]));
	notech_inv i_33411(.A(to_acu100236[5]), .Z(to_acu[5]));
	notech_inv i_33412(.A(to_acu100236[6]), .Z(to_acu[6]));
	notech_inv i_33413(.A(to_acu100236[7]), .Z(to_acu[7]));
	notech_inv i_33414(.A(to_acu100236[8]), .Z(to_acu[8]));
	notech_inv i_33415(.A(to_acu100236[9]), .Z(to_acu[9]));
	notech_inv i_33416(.A(to_acu100236[10]), .Z(to_acu[10]));
	notech_inv i_33417(.A(to_acu100236[11]), .Z(to_acu[11]));
	notech_inv i_33418(.A(to_acu100236[12]), .Z(to_acu[12]));
	notech_inv i_33419(.A(to_acu100236[13]), .Z(to_acu[13]));
	notech_inv i_33420(.A(to_acu100236[14]), .Z(to_acu[14]));
	notech_inv i_33421(.A(to_acu100236[15]), .Z(to_acu[15]));
	notech_inv i_33422(.A(to_acu100236[16]), .Z(to_acu[16]));
	notech_inv i_33423(.A(to_acu100236[17]), .Z(to_acu[17]));
	notech_inv i_33424(.A(to_acu100236[18]), .Z(to_acu[18]));
	notech_inv i_33425(.A(to_acu100236[19]), .Z(to_acu[19]));
	notech_inv i_33426(.A(to_acu100236[20]), .Z(to_acu[20]));
	notech_inv i_33427(.A(to_acu100236[21]), .Z(to_acu[21]));
	notech_inv i_33428(.A(to_acu100236[22]), .Z(to_acu[22]));
	notech_inv i_33429(.A(to_acu100236[23]), .Z(to_acu[23]));
	notech_inv i_33430(.A(to_acu100236[24]), .Z(to_acu[24]));
	notech_inv i_33431(.A(to_acu100236[25]), .Z(to_acu[25]));
	notech_inv i_33432(.A(to_acu100236[26]), .Z(to_acu[26]));
	notech_inv i_33433(.A(to_acu100236[27]), .Z(to_acu[27]));
	notech_inv i_33434(.A(to_acu100236[28]), .Z(to_acu[28]));
	notech_inv i_33435(.A(to_acu100236[29]), .Z(to_acu[29]));
	notech_inv i_33436(.A(to_acu100236[30]), .Z(to_acu[30]));
	notech_inv i_33437(.A(to_acu100236[31]), .Z(to_acu[31]));
	notech_inv i_33438(.A(to_acu100236[32]), .Z(to_acu[32]));
	notech_inv i_33439(.A(to_acu100236[33]), .Z(to_acu[33]));
	notech_inv i_33440(.A(to_acu100236[34]), .Z(to_acu[34]));
	notech_inv i_33441(.A(to_acu100236[35]), .Z(to_acu[35]));
	notech_inv i_33442(.A(to_acu100236[36]), .Z(to_acu[36]));
	notech_inv i_33443(.A(to_acu100236[37]), .Z(to_acu[37]));
	notech_inv i_33444(.A(to_acu100236[38]), .Z(to_acu[38]));
	notech_inv i_33445(.A(to_acu100236[39]), .Z(to_acu[39]));
	notech_inv i_33446(.A(to_acu100236[40]), .Z(to_acu[40]));
	notech_inv i_33447(.A(to_acu100236[41]), .Z(to_acu[41]));
	notech_inv i_33448(.A(to_acu100236[42]), .Z(to_acu[42]));
	notech_inv i_33449(.A(to_acu100236[43]), .Z(to_acu[43]));
	notech_inv i_33450(.A(to_acu100236[44]), .Z(to_acu[44]));
	notech_inv i_33451(.A(to_acu100236[45]), .Z(to_acu[45]));
	notech_inv i_33452(.A(to_acu100236[46]), .Z(to_acu[46]));
	notech_inv i_33453(.A(to_acu100236[47]), .Z(to_acu[47]));
	notech_inv i_33454(.A(to_acu100236[48]), .Z(to_acu[48]));
	notech_inv i_33455(.A(to_acu100236[49]), .Z(to_acu[49]));
	notech_inv i_33456(.A(to_acu100236[50]), .Z(to_acu[50]));
	notech_inv i_33457(.A(to_acu100236[51]), .Z(to_acu[51]));
	notech_inv i_33458(.A(to_acu100236[52]), .Z(to_acu[52]));
	notech_inv i_33459(.A(to_acu100236[53]), .Z(to_acu[53]));
	notech_inv i_33460(.A(to_acu100236[54]), .Z(to_acu[54]));
	notech_inv i_33461(.A(to_acu100236[55]), .Z(to_acu[55]));
	notech_inv i_33462(.A(to_acu100236[56]), .Z(to_acu[56]));
	notech_inv i_33463(.A(to_acu100236[57]), .Z(to_acu[57]));
	notech_inv i_33464(.A(to_acu100236[58]), .Z(to_acu[58]));
	notech_inv i_33465(.A(to_acu100236[59]), .Z(to_acu[59]));
	notech_inv i_33466(.A(to_acu100236[60]), .Z(to_acu[60]));
	notech_inv i_33467(.A(to_acu100236[61]), .Z(to_acu[61]));
	notech_inv i_33468(.A(to_acu100236[62]), .Z(to_acu[62]));
	notech_inv i_33469(.A(to_acu100236[63]), .Z(to_acu[63]));
	notech_inv i_33470(.A(divq[0]), .Z(n_29474));
	notech_inv i_33471(.A(divq[1]), .Z(n_29475));
	notech_inv i_33472(.A(divq[2]), .Z(n_29476));
	notech_inv i_33473(.A(divq[3]), .Z(n_29477));
	notech_inv i_33474(.A(divq[4]), .Z(n_29478));
	notech_inv i_33475(.A(divq[5]), .Z(n_29479));
	notech_inv i_33476(.A(divq[6]), .Z(n_29480));
	notech_inv i_33477(.A(divq[7]), .Z(n_29481));
	notech_inv i_33478(.A(divq[8]), .Z(n_29482));
	notech_inv i_33479(.A(divq[9]), .Z(n_29483));
	notech_inv i_33480(.A(divq[10]), .Z(n_29484));
	notech_inv i_33481(.A(divq[11]), .Z(n_29485));
	notech_inv i_33482(.A(divq[12]), .Z(n_29486));
	notech_inv i_33483(.A(divq[13]), .Z(n_29487));
	notech_inv i_33484(.A(divq[14]), .Z(n_29488));
	notech_inv i_33485(.A(divq[15]), .Z(n_29489));
	notech_inv i_33486(.A(divq[16]), .Z(n_29490));
	notech_inv i_33487(.A(divq[17]), .Z(n_29491));
	notech_inv i_33488(.A(divq[18]), .Z(n_29492));
	notech_inv i_33489(.A(divq[19]), .Z(n_29493));
	notech_inv i_33490(.A(divq[20]), .Z(n_29494));
	notech_inv i_33491(.A(divq[21]), .Z(n_29495));
	notech_inv i_33492(.A(divq[22]), .Z(n_29496));
	notech_inv i_33493(.A(divq[23]), .Z(n_29497));
	notech_inv i_33494(.A(divq[24]), .Z(n_29498));
	notech_inv i_33495(.A(divq[25]), .Z(n_29499));
	notech_inv i_33496(.A(divq[26]), .Z(n_29500));
	notech_inv i_33497(.A(divq[27]), .Z(n_29501));
	notech_inv i_33498(.A(divq[28]), .Z(n_29502));
	notech_inv i_33499(.A(divq[29]), .Z(n_29503));
	notech_inv i_33500(.A(divq[30]), .Z(n_29504));
	notech_inv i_33501(.A(divq[31]), .Z(n_29505));
	notech_inv i_33502(.A(divq[32]), .Z(n_29506));
	notech_inv i_33503(.A(divq[33]), .Z(n_29507));
	notech_inv i_33504(.A(divq[34]), .Z(n_29508));
	notech_inv i_33505(.A(divq[35]), .Z(n_29509));
	notech_inv i_33506(.A(divq[36]), .Z(n_29510));
	notech_inv i_33507(.A(divq[37]), .Z(n_29511));
	notech_inv i_33508(.A(divq[38]), .Z(n_29512));
	notech_inv i_33509(.A(divq[39]), .Z(n_29513));
	notech_inv i_33510(.A(divq[40]), .Z(n_29514));
	notech_inv i_33511(.A(divq[41]), .Z(n_29515));
	notech_inv i_33512(.A(divq[42]), .Z(n_29516));
	notech_inv i_33513(.A(divq[43]), .Z(n_29517));
	notech_inv i_33514(.A(divq[44]), .Z(n_29518));
	notech_inv i_33515(.A(divq[45]), .Z(n_29519));
	notech_inv i_33516(.A(divq[46]), .Z(n_29520));
	notech_inv i_33517(.A(divq[47]), .Z(n_29521));
	notech_inv i_33518(.A(divq[48]), .Z(n_29522));
	notech_inv i_33519(.A(divq[49]), .Z(n_29523));
	notech_inv i_33520(.A(divq[50]), .Z(n_29524));
	notech_inv i_33521(.A(divq[51]), .Z(n_29525));
	notech_inv i_33522(.A(divq[52]), .Z(n_29526));
	notech_inv i_33523(.A(divq[53]), .Z(n_29527));
	notech_inv i_33524(.A(divq[54]), .Z(n_29528));
	notech_inv i_33525(.A(divq[55]), .Z(n_29529));
	notech_inv i_33526(.A(divq[56]), .Z(n_29530));
	notech_inv i_33527(.A(divq[57]), .Z(n_29531));
	notech_inv i_33528(.A(divq[58]), .Z(n_29532));
	notech_inv i_33529(.A(divq[59]), .Z(n_29533));
	notech_inv i_33530(.A(divq[60]), .Z(n_29534));
	notech_inv i_33531(.A(divq[61]), .Z(n_29535));
	notech_inv i_33532(.A(divq[62]), .Z(n_29536));
	notech_inv i_33533(.A(divq[63]), .Z(n_29537));
	notech_inv i_33534(.A(add_len_pc[0]), .Z(n_29538));
	notech_inv i_33535(.A(add_len_pc[1]), .Z(n_29539));
	notech_inv i_33536(.A(add_len_pc[2]), .Z(n_29540));
	notech_inv i_33537(.A(add_len_pc[3]), .Z(n_29541));
	notech_inv i_33538(.A(add_len_pc[4]), .Z(n_29542));
	notech_inv i_33539(.A(add_len_pc[5]), .Z(n_29543));
	notech_inv i_33540(.A(add_len_pc[7]), .Z(n_29544));
	notech_inv i_33541(.A(add_len_pc[8]), .Z(n_29545));
	notech_inv i_33542(.A(add_len_pc[9]), .Z(n_29546));
	notech_inv i_33543(.A(add_len_pc[10]), .Z(n_29547));
	notech_inv i_33544(.A(add_len_pc[11]), .Z(n_29548));
	notech_inv i_33545(.A(add_len_pc[12]), .Z(n_29549));
	notech_inv i_33546(.A(add_len_pc[13]), .Z(n_29550));
	notech_inv i_33547(.A(add_len_pc[14]), .Z(n_29551));
	notech_inv i_33548(.A(add_len_pc[15]), .Z(n_29552));
	notech_inv i_33549(.A(add_len_pc[21]), .Z(n_29553));
	notech_inv i_33550(.A(add_len_pc[30]), .Z(n_29554));
	notech_inv i_33551(.A(divr[0]), .Z(nbus_11328[0]));
	notech_inv i_33552(.A(divr[1]), .Z(nbus_11328[1]));
	notech_inv i_33553(.A(divr[2]), .Z(nbus_11328[2]));
	notech_inv i_33554(.A(divr[3]), .Z(nbus_11328[3]));
	notech_inv i_33555(.A(divr[4]), .Z(nbus_11328[4]));
	notech_inv i_33556(.A(divr[5]), .Z(nbus_11328[5]));
	notech_inv i_33557(.A(divr[6]), .Z(nbus_11328[6]));
	notech_inv i_33558(.A(divr[7]), .Z(nbus_11328[7]));
	notech_inv i_33559(.A(divr[8]), .Z(nbus_11328[8]));
	notech_inv i_33560(.A(divr[9]), .Z(nbus_11328[9]));
	notech_inv i_33561(.A(divr[10]), .Z(nbus_11328[10]));
	notech_inv i_33562(.A(divr[11]), .Z(nbus_11328[11]));
	notech_inv i_33563(.A(divr[12]), .Z(nbus_11328[12]));
	notech_inv i_33564(.A(divr[13]), .Z(nbus_11328[13]));
	notech_inv i_33565(.A(divr[14]), .Z(nbus_11328[14]));
	notech_inv i_33566(.A(divr[15]), .Z(nbus_11328[15]));
	notech_inv i_33567(.A(divr[16]), .Z(nbus_11328[16]));
	notech_inv i_33568(.A(divr[17]), .Z(nbus_11328[17]));
	notech_inv i_33569(.A(divr[18]), .Z(nbus_11328[18]));
	notech_inv i_33570(.A(divr[19]), .Z(nbus_11328[19]));
	notech_inv i_33571(.A(divr[20]), .Z(nbus_11328[20]));
	notech_inv i_33572(.A(divr[21]), .Z(nbus_11328[21]));
	notech_inv i_33573(.A(divr[22]), .Z(nbus_11328[22]));
	notech_inv i_33574(.A(divr[23]), .Z(nbus_11328[23]));
	notech_inv i_33575(.A(divr[24]), .Z(nbus_11328[24]));
	notech_inv i_33576(.A(divr[25]), .Z(nbus_11328[25]));
	notech_inv i_33577(.A(divr[26]), .Z(nbus_11328[26]));
	notech_inv i_33578(.A(divr[27]), .Z(nbus_11328[27]));
	notech_inv i_33579(.A(divr[28]), .Z(nbus_11328[28]));
	notech_inv i_33580(.A(divr[29]), .Z(nbus_11328[29]));
	notech_inv i_33581(.A(divr[30]), .Z(nbus_11328[30]));
	notech_inv i_33583(.A(divr[31]), .Z(nbus_11328[31]));
	notech_inv i_33584(.A(n_6364), .Z(n_29587));
	notech_inv i_33585(.A(n_7341), .Z(n_29588));
	notech_inv i_33586(.A(n_7303), .Z(n_29589));
	notech_inv i_33587(.A(n_7304), .Z(n_29590));
	notech_inv i_33588(.A(\regs_13_14[30] ), .Z(n_29591));
	notech_inv i_33589(.A(\opa_12[13] ), .Z(n_29592));
	notech_inv i_33590(.A(n_11432), .Z(n_29593));
	notech_inv i_33591(.A(n_6401), .Z(n_29594));
	notech_inv i_33592(.A(n_6402), .Z(n_29595));
	notech_inv i_33593(.A(\opa_12[11] ), .Z(n_29596));
	notech_inv i_33594(.A(n_7336), .Z(n_29597));
	notech_inv i_33595(.A(n_7335), .Z(n_29598));
	notech_inv i_33596(.A(n_7334), .Z(n_29600));
	notech_inv i_33597(.A(n_56172), .Z(n_29601));
	notech_inv i_33598(.A(n_7333), .Z(n_29602));
	notech_inv i_33599(.A(n_7375), .Z(n_29604));
	notech_inv i_33600(.A(\regs_1_0[28] ), .Z(n_29605));
	notech_inv i_33602(.A(\nbus_14523[26] ), .Z(n_29606));
	notech_inv i_33603(.A(\eflags[26] ), .Z(n_29607));
	notech_inv i_33604(.A(\nbus_14523[27] ), .Z(n_29608));
	notech_inv i_33605(.A(\eflags[27] ), .Z(n_29609));
	notech_inv i_33606(.A(\nbus_14523[28] ), .Z(n_29610));
	notech_inv i_33607(.A(\eflags[28] ), .Z(n_29611));
	notech_inv i_33608(.A(\nbus_14523[29] ), .Z(n_29612));
	notech_inv i_33609(.A(\eflags[29] ), .Z(n_29613));
	notech_inv i_33610(.A(\opa_12[7] ), .Z(n_29614));
	notech_inv i_33611(.A(\eflags[7] ), .Z(n_29615));
	notech_inv i_33612(.A(\nbus_14523[7] ), .Z(n_29616));
	notech_inv i_33614(.A(\nbus_14523[31] ), .Z(n_29617));
	notech_inv i_33615(.A(\eflags[31] ), .Z(n_29618));
	notech_inv i_33616(.A(\regs_13_14[31] ), .Z(n_29619));
	notech_inv i_33618(.A(\eflags[11] ), .Z(n_29620));
	notech_inv i_33619(.A(\nbus_14523[11] ), .Z(n_29621));
	notech_inv i_33620(.A(\eflags[13] ), .Z(n_29622));
	notech_inv i_33621(.A(\nbus_14523[13] ), .Z(n_29623));
	notech_inv i_33622(.A(\nbus_14523[30] ), .Z(n_29624));
	notech_inv i_33623(.A(\eflags[30] ), .Z(n_29625));
	notech_inv i_33624(.A(\opa_1[5] ), .Z(n_29626));
	notech_inv i_33625(.A(n_10906), .Z(n_29627));
	notech_inv i_33626(.A(instrc[97]), .Z(n_29628));
	notech_inv i_33627(.A(instrc[89]), .Z(n_29631));
	notech_inv i_33628(.A(instrc[124]), .Z(n_29632));
	notech_inv i_33629(.A(instrc[100]), .Z(n_29633));
	notech_inv i_33630(.A(instrc[92]), .Z(n_29634));
	notech_inv i_33631(.A(instrc[101]), .Z(n_29635));
	notech_inv i_33632(.A(instrc[93]), .Z(n_29636));
	notech_inv i_33633(.A(instrc[103]), .Z(n_29637));
	notech_inv i_33634(.A(instrc[95]), .Z(n_29638));
	notech_inv i_33635(.A(instrc[99]), .Z(n_29639));
	notech_inv i_33636(.A(instrc[91]), .Z(n_29640));
	notech_inv i_33637(.A(instrc[96]), .Z(n_29641));
	notech_inv i_33638(.A(instrc[88]), .Z(n_29642));
	notech_inv i_33639(.A(instrc[81]), .Z(n_29643));
	notech_inv i_33640(.A(instrc[82]), .Z(n_29644));
	notech_inv i_33641(.A(instrc[80]), .Z(n_29645));
	notech_inv i_33642(.A(instrc[83]), .Z(n_29646));
	notech_inv i_33643(.A(instrc[84]), .Z(n_29647));
	notech_inv i_33644(.A(instrc[86]), .Z(n_29648));
	notech_inv i_33645(.A(instrc[87]), .Z(n_29649));
	notech_inv i_33646(.A(instrc[85]), .Z(n_29650));
	notech_inv i_33647(.A(\opa_12[5] ), .Z(n_29651));
	notech_inv i_33648(.A(n_57064), .Z(n_29652));
	notech_inv i_33649(.A(n_57042), .Z(n_29653));
	notech_inv i_33650(.A(n_61136), .Z(n_29654));
	notech_inv i_33651(.A(read_ack), .Z(n_29655));
	notech_inv i_33652(.A(n_5221), .Z(n_29656));
	notech_inv i_33653(.A(n_5219), .Z(n_29657));
	notech_inv i_33654(.A(n_57082), .Z(n_29658));
	notech_inv i_33655(.A(\regs_13_14[29] ), .Z(n_29659));
	notech_inv i_33656(.A(\regs_13_14[26] ), .Z(n_29660));
	notech_inv i_33657(.A(\regs_13_14[27] ), .Z(n_29661));
	notech_inv i_33658(.A(\regs_13_14[28] ), .Z(n_29662));
	notech_inv i_33659(.A(instrc[127]), .Z(n_29663));
	notech_inv i_33660(.A(instrc[126]), .Z(n_29664));
	notech_inv i_33661(.A(instrc[102]), .Z(n_29665));
	notech_inv i_33662(.A(instrc[94]), .Z(n_29666));
	notech_inv i_33663(.A(instrc[98]), .Z(n_29667));
	notech_inv i_33664(.A(instrc[90]), .Z(n_29668));
	notech_inv i_33665(.A(\regs_1_0[21] ), .Z(n_29669));
	notech_inv i_33666(.A(\regs_1[14] ), .Z(n_29670));
	notech_inv i_33667(.A(n_8128), .Z(n_29671));
	notech_inv i_33668(.A(\regs_1[13] ), .Z(n_29672));
	notech_inv i_33669(.A(n_8127), .Z(n_29673));
	notech_inv i_33670(.A(\regs_1[12] ), .Z(n_29674));
	notech_inv i_33671(.A(n_8126), .Z(n_29675));
	notech_inv i_33672(.A(\regs_1[1] ), .Z(n_29676));
	notech_inv i_33673(.A(n_8115), .Z(n_29677));
	notech_inv i_33674(.A(\opa_12[1] ), .Z(n_29678));
	notech_inv i_33675(.A(\opa_12[12] ), .Z(n_29679));
	notech_inv i_33676(.A(\opa_12[14] ), .Z(n_29680));
	notech_inv i_33677(.A(\regs_13_14[21] ), .Z(n_29681));
	notech_inv i_33678(.A(n_8124), .Z(n_29682));
	notech_inv i_33679(.A(\regs_1[10] ), .Z(n_29683));
	notech_inv i_33680(.A(\opa_12[10] ), .Z(n_29684));
	notech_inv i_33681(.A(\regs_1_0[30] ), .Z(n_29685));
	notech_inv i_33682(.A(n_6407), .Z(n_29687));
	notech_inv i_33683(.A(n_6408), .Z(n_29689));
	notech_inv i_33684(.A(n_6405), .Z(n_29690));
	notech_inv i_33685(.A(n_6406), .Z(n_29691));
	notech_inv i_33686(.A(nCF_shiftbox), .Z(n_29692));
	notech_inv i_33687(.A(nCF_arithbox), .Z(n_29693));
	notech_inv i_33688(.A(n_7340), .Z(n_29695));
	notech_inv i_33689(.A(n_7339), .Z(n_29696));
	notech_inv i_33690(.A(n_7338), .Z(n_29697));
	notech_inv i_33691(.A(n_7337), .Z(n_29698));
	notech_inv i_33692(.A(n_7378), .Z(n_29699));
	notech_inv i_33693(.A(n_7377), .Z(n_29700));
	notech_inv i_33694(.A(n_11313), .Z(n_29701));
	notech_inv i_33695(.A(n_9887), .Z(n_29702));
	notech_inv i_33696(.A(n_11314), .Z(n_29704));
	notech_inv i_33697(.A(\regs_1_0[22] ), .Z(n_29705));
	notech_inv i_33698(.A(n_8116), .Z(n_29706));
	notech_inv i_33699(.A(\regs_1[2] ), .Z(n_29707));
	notech_inv i_33700(.A(\regs_13_14[22] ), .Z(n_29708));
	notech_inv i_33701(.A(\regs_1_0[18] ), .Z(n_29709));
	notech_inv i_33702(.A(\regs_13_14[16] ), .Z(n_29710));
	notech_inv i_33703(.A(\regs_13_14[18] ), .Z(n_29711));
	notech_inv i_33704(.A(\eflags[18] ), .Z(n_29712));
	notech_inv i_33705(.A(\nbus_14523[18] ), .Z(n_29713));
	notech_inv i_33706(.A(n_8120), .Z(n_29714));
	notech_inv i_33707(.A(\regs_1[6] ), .Z(n_29715));
	notech_inv i_33708(.A(n_8119), .Z(n_29716));
	notech_inv i_33709(.A(n_8117), .Z(n_29717));
	notech_inv i_33710(.A(\eflags[6] ), .Z(n_29718));
	notech_inv i_33711(.A(\nbus_14523[6] ), .Z(n_29719));
	notech_inv i_33712(.A(\nbus_14523[10] ), .Z(n_29720));
	notech_inv i_33713(.A(n_10908), .Z(n_29721));
	notech_inv i_33714(.A(\opa_1[7] ), .Z(n_29722));
	notech_inv i_33715(.A(\opa_12[6] ), .Z(n_29723));
	notech_inv i_33716(.A(\opa_1[6] ), .Z(n_29724));
	notech_inv i_33718(.A(\opa_12[4] ), .Z(n_29725));
	notech_inv i_33719(.A(n_10905), .Z(n_29726));
	notech_inv i_33721(.A(\opa_1[4] ), .Z(n_29727));
	notech_inv i_33722(.A(\opa_12[3] ), .Z(n_29728));
	notech_inv i_33724(.A(n_10904), .Z(n_29729));
	notech_inv i_33725(.A(\opa_1[3] ), .Z(n_29730));
	notech_inv i_33726(.A(n_10903), .Z(n_29731));
	notech_inv i_33727(.A(\opa_1[2] ), .Z(n_29732));
	notech_inv i_33728(.A(\opa_12[2] ), .Z(n_29733));
	notech_inv i_33729(.A(instrc[107]), .Z(n_29734));
	notech_inv i_33730(.A(instrc[104]), .Z(n_29735));
	notech_inv i_33731(.A(n_57369), .Z(n_29736));
	notech_inv i_33732(.A(instrc[105]), .Z(n_29737));
	notech_inv i_33733(.A(n_9229), .Z(n_29738));
	notech_inv i_33734(.A(n_9230), .Z(n_29739));
	notech_inv i_33735(.A(n_9231), .Z(n_29740));
	notech_inv i_33736(.A(n_328963506), .Z(n_29741));
	notech_inv i_33737(.A(\opa_12[0] ), .Z(n_29742));
	notech_inv i_33738(.A(\opa_12[9] ), .Z(n_29743));
	notech_inv i_33739(.A(readio_ack), .Z(n_29744));
	notech_inv i_33740(.A(n_8118), .Z(n_29745));
	notech_inv i_33741(.A(\regs_1[4] ), .Z(n_29746));
	notech_inv i_33742(.A(n_8121), .Z(n_29747));
	notech_inv i_33743(.A(\regs_1[7] ), .Z(n_29748));
	notech_inv i_33744(.A(n_8123), .Z(n_29749));
	notech_inv i_33745(.A(\regs_1[9] ), .Z(n_29750));
	notech_inv i_33746(.A(n_8125), .Z(n_29751));
	notech_inv i_33747(.A(\regs_1[11] ), .Z(n_29752));
	notech_inv i_33748(.A(\regs_1[15] ), .Z(n_29753));
	notech_inv i_33749(.A(\opa_12[15] ), .Z(n_29754));
	notech_inv i_33750(.A(n_8114), .Z(n_29755));
	notech_inv i_33751(.A(n_11431), .Z(n_29756));
	notech_inv i_33752(.A(n_11430), .Z(n_29757));
	notech_inv i_33753(.A(n_11429), .Z(n_29758));
	notech_inv i_33754(.A(n_6403), .Z(n_29759));
	notech_inv i_33755(.A(n_6404), .Z(n_29760));
	notech_inv i_33756(.A(n_7376), .Z(n_29761));
	notech_inv i_33757(.A(n_11309), .Z(n_29762));
	notech_inv i_33758(.A(n_9885), .Z(n_29763));
	notech_inv i_33759(.A(n_11310), .Z(n_29764));
	notech_inv i_33760(.A(\regs_13_14[23] ), .Z(n_29765));
	notech_inv i_33761(.A(\regs_13_14[24] ), .Z(n_29769));
	notech_inv i_33762(.A(\regs_13_14[25] ), .Z(n_29770));
	notech_inv i_33763(.A(start_up), .Z(n_29771));
	notech_inv i_33764(.A(\regs_13_14[17] ), .Z(n_29772));
	notech_inv i_33765(.A(\regs_13_14[19] ), .Z(n_29773));
	notech_inv i_33766(.A(\regs_13_14[20] ), .Z(n_29775));
	notech_inv i_33767(.A(n_11419), .Z(n_29776));
	notech_inv i_33768(.A(n_11420), .Z(n_29779));
	notech_inv i_33769(.A(n_11422), .Z(n_29780));
	notech_inv i_33770(.A(n_11423), .Z(n_29784));
	notech_inv i_33771(.A(n_11424), .Z(n_29785));
	notech_inv i_33772(.A(n_8122), .Z(n_29786));
	notech_inv i_33773(.A(\opa_12[8] ), .Z(n_29787));
	notech_inv i_33774(.A(\nbus_14523[9] ), .Z(n_29788));
	notech_inv i_33775(.A(ie), .Z(n_29789));
	notech_inv i_33776(.A(\nbus_14523[4] ), .Z(n_29790));
	notech_inv i_33777(.A(\eflags[4] ), .Z(n_29791));
	notech_inv i_33778(.A(\eflags[0] ), .Z(n_29792));
	notech_inv i_33779(.A(n_61515), .Z(n_29793));
	notech_inv i_33780(.A(n_7356), .Z(n_29794));
	notech_inv i_33781(.A(n_7360), .Z(n_29795));
	notech_inv i_33782(.A(n_7361), .Z(n_29796));
	notech_inv i_33783(.A(n_7363), .Z(n_29797));
	notech_inv i_33784(.A(n_7370), .Z(n_29798));
	notech_inv i_33785(.A(n_7379), .Z(n_29799));
	notech_inv i_33786(.A(n_7295), .Z(n_29800));
	notech_inv i_33787(.A(n_7296), .Z(n_29801));
	notech_inv i_33788(.A(n_7309), .Z(n_29802));
	notech_inv i_33789(.A(n_7310), .Z(n_29803));
	notech_inv i_33790(.A(n_7323), .Z(n_29804));
	notech_inv i_33791(.A(n_6352), .Z(n_29805));
	notech_inv i_33792(.A(n_6351), .Z(n_29806));
	notech_inv i_33793(.A(n_6358), .Z(n_29807));
	notech_inv i_33794(.A(n_6357), .Z(n_29808));
	notech_inv i_33795(.A(n_6368), .Z(n_29809));
	notech_inv i_33796(.A(n_6372), .Z(n_29810));
	notech_inv i_33797(.A(n_6371), .Z(n_29811));
	notech_inv i_33798(.A(n_6375), .Z(n_29812));
	notech_inv i_33799(.A(n_6376), .Z(n_29813));
	notech_inv i_33800(.A(n_6377), .Z(n_29814));
	notech_inv i_33801(.A(n_6378), .Z(n_29815));
	notech_inv i_33802(.A(n_6392), .Z(n_29816));
	notech_inv i_33803(.A(n_6391), .Z(n_29817));
	notech_inv i_33804(.A(n_6410), .Z(n_29818));
	notech_inv i_33805(.A(n_6409), .Z(n_29819));
	notech_inv i_33806(.A(n_7359), .Z(n_29820));
	notech_inv i_33807(.A(n_6349), .Z(n_29821));
	notech_inv i_33808(.A(n_6350), .Z(n_29822));
	notech_inv i_33809(.A(n_6370), .Z(n_29823));
	notech_inv i_33810(.A(n_6369), .Z(n_29824));
	notech_inv i_33811(.A(n_6374), .Z(n_29825));
	notech_inv i_33812(.A(n_6373), .Z(n_29826));
	notech_inv i_33813(.A(n_7374), .Z(n_29827));
	notech_inv i_33814(.A(n_6354), .Z(n_29828));
	notech_inv i_33815(.A(n_6353), .Z(n_29830));
	notech_inv i_33816(.A(n_6394), .Z(n_29831));
	notech_inv i_33817(.A(n_6396), .Z(n_29832));
	notech_inv i_33818(.A(n_6398), .Z(n_29833));
	notech_inv i_33819(.A(n_6400), .Z(n_29834));
	notech_inv i_33820(.A(\nbus_14523[22] ), .Z(n_29835));
	notech_inv i_33821(.A(\eflags[22] ), .Z(n_29837));
	notech_inv i_33822(.A(\nbus_14523[23] ), .Z(n_29838));
	notech_inv i_33823(.A(\eflags[23] ), .Z(n_29839));
	notech_inv i_33824(.A(\nbus_14523[24] ), .Z(n_29840));
	notech_inv i_33825(.A(\eflags[24] ), .Z(n_29841));
	notech_inv i_33826(.A(n_7365), .Z(n_29842));
	notech_inv i_33827(.A(n_7366), .Z(n_29843));
	notech_inv i_33828(.A(n_7367), .Z(n_29844));
	notech_inv i_33829(.A(n_7368), .Z(n_29845));
	notech_inv i_33830(.A(n_7369), .Z(n_29846));
	notech_inv i_33831(.A(n_6382), .Z(n_29847));
	notech_inv i_33832(.A(n_6384), .Z(n_29848));
	notech_inv i_33833(.A(n_6386), .Z(n_29849));
	notech_inv i_33834(.A(n_6388), .Z(n_29850));
	notech_inv i_33835(.A(n_6390), .Z(n_29851));
	notech_inv i_33836(.A(\nbus_14523[16] ), .Z(n_29852));
	notech_inv i_33837(.A(\eflags[16] ), .Z(n_29853));
	notech_inv i_33838(.A(\nbus_14523[21] ), .Z(n_29854));
	notech_inv i_33839(.A(\eflags[21] ), .Z(n_29855));
	notech_inv i_33840(.A(n_7354), .Z(n_29856));
	notech_inv i_33841(.A(n_6356), .Z(n_29857));
	notech_inv i_33842(.A(n_6360), .Z(n_29858));
	notech_inv i_33843(.A(\nbus_14523[5] ), .Z(n_29859));
	notech_inv i_33844(.A(\eflags[5] ), .Z(n_29860));
	notech_inv i_33845(.A(n_7357), .Z(n_29861));
	notech_inv i_33846(.A(n_6366), .Z(n_29862));
	notech_inv i_33847(.A(\nbus_14523[8] ), .Z(n_29863));
	notech_inv i_33848(.A(\eflags[8] ), .Z(n_29864));
	notech_inv i_33849(.A(\nbus_14523[15] ), .Z(n_29865));
	notech_inv i_33850(.A(\eflags[15] ), .Z(n_29866));
	notech_inv i_33851(.A(\nbus_14523[14] ), .Z(n_29867));
	notech_inv i_33852(.A(\eflags[14] ), .Z(n_29868));
	notech_inv i_33853(.A(\eflags[1] ), .Z(n_29869));
	notech_inv i_33854(.A(n_7362), .Z(n_29870));
	notech_inv i_33855(.A(n_7283), .Z(n_29871));
	notech_inv i_33856(.A(n_7289), .Z(n_29872));
	notech_inv i_33857(.A(n_7306), .Z(n_29873));
	notech_inv i_33858(.A(n_7305), .Z(n_29874));
	notech_inv i_33859(.A(n_7307), .Z(n_29875));
	notech_inv i_33860(.A(n_7308), .Z(n_29876));
	notech_inv i_33861(.A(n_7282), .Z(n_29877));
	notech_inv i_33862(.A(n_7281), .Z(n_29878));
	notech_inv i_33863(.A(n_7301), .Z(n_29879));
	notech_inv i_33864(.A(n_7302), .Z(n_29880));
	notech_inv i_33865(.A(\regs_1_0[25] ), .Z(n_29881));
	notech_inv i_33866(.A(n_7285), .Z(n_29882));
	notech_inv i_33867(.A(n_7286), .Z(n_29883));
	notech_inv i_33868(.A(n_7331), .Z(n_29884));
	notech_inv i_33869(.A(n_11428), .Z(n_29885));
	notech_inv i_33870(.A(\nbus_14523[25] ), .Z(n_29886));
	notech_inv i_33871(.A(\eflags[25] ), .Z(n_29887));
	notech_inv i_33872(.A(n_7313), .Z(n_29888));
	notech_inv i_33873(.A(n_7314), .Z(n_29889));
	notech_inv i_33874(.A(n_7287), .Z(n_29890));
	notech_inv i_33875(.A(n_7291), .Z(n_29891));
	notech_inv i_33876(.A(\nbus_14523[3] ), .Z(n_29892));
	notech_inv i_33877(.A(\eflags[3] ), .Z(n_29893));
	notech_inv i_33878(.A(n_7297), .Z(n_29894));
	notech_inv i_33879(.A(\nbus_14523[12] ), .Z(n_29896));
	notech_inv i_33880(.A(\eflags[12] ), .Z(n_29898));
	notech_inv i_33881(.A(n_9239), .Z(n_29899));
	notech_inv i_33882(.A(n_9240), .Z(n_29900));
	notech_inv i_33883(.A(n_9234), .Z(n_29901));
	notech_inv i_33884(.A(n_9235), .Z(n_29903));
	notech_inv i_33885(.A(n_346373943), .Z(n_29904));
	notech_inv i_33886(.A(n_7350), .Z(n_29906));
	notech_inv i_33887(.A(n_7353), .Z(n_29908));
	notech_inv i_33888(.A(\regs_1_0[23] ), .Z(n_29910));
	notech_inv i_33889(.A(\regs_1_0[24] ), .Z(n_29911));
	notech_inv i_33890(.A(n_7351), .Z(n_29913));
	notech_inv i_33891(.A(n_7371), .Z(n_29914));
	notech_inv i_33892(.A(n_7372), .Z(n_29916));
	notech_inv i_33893(.A(n_7373), .Z(n_29918));
	notech_inv i_33894(.A(n_7325), .Z(n_29926));
	notech_inv i_33895(.A(n_7327), .Z(n_29927));
	notech_inv i_33896(.A(n_7329), .Z(n_29928));
	notech_inv i_33897(.A(n_11405), .Z(n_29929));
	notech_inv i_33898(.A(\nbus_14523[2] ), .Z(n_29930));
	notech_inv i_33899(.A(\eflags[2] ), .Z(n_29931));
	notech_inv i_33900(.A(\regs_1_0[20] ), .Z(n_29932));
	notech_inv i_33901(.A(n_7315), .Z(n_29933));
	notech_inv i_33902(.A(n_7317), .Z(n_29935));
	notech_inv i_33903(.A(n_7319), .Z(n_29936));
	notech_inv i_33905(.A(n_7321), .Z(n_29937));
	notech_inv i_33906(.A(\nbus_14523[17] ), .Z(n_29938));
	notech_inv i_33907(.A(\eflags[17] ), .Z(n_29939));
	notech_inv i_33908(.A(n_11421), .Z(n_29940));
	notech_inv i_33910(.A(\nbus_14523[19] ), .Z(n_29941));
	notech_inv i_33911(.A(\eflags[19] ), .Z(n_29942));
	notech_inv i_33912(.A(\nbus_14523[20] ), .Z(n_29943));
	notech_inv i_33913(.A(\eflags[20] ), .Z(n_29944));
	notech_inv i_33914(.A(n_7352), .Z(n_29945));
	notech_inv i_33915(.A(n_11406), .Z(n_29946));
	notech_inv i_33916(.A(n_11408), .Z(n_29947));
	notech_inv i_33917(.A(n_11409), .Z(n_29948));
	notech_inv i_33918(.A(n_11410), .Z(n_29949));
	notech_inv i_33919(.A(n_11425), .Z(n_29950));
	notech_inv i_33920(.A(n_11426), .Z(n_29951));
	notech_inv i_33921(.A(n_11427), .Z(n_29952));
	notech_inv i_33922(.A(\opa_1[0] ), .Z(n_29953));
	notech_inv i_33923(.A(\opa_1[1] ), .Z(n_29955));
	notech_inv i_33925(.A(mul64[8]), .Z(n_29956));
	notech_inv i_33926(.A(\opa_1[8] ), .Z(n_29958));
	notech_inv i_33927(.A(n_10909), .Z(n_29959));
	notech_inv i_33928(.A(mul64[9]), .Z(n_29960));
	notech_inv i_33929(.A(\opa_1[9] ), .Z(n_29961));
	notech_inv i_33930(.A(n_10910), .Z(n_29962));
	notech_inv i_33931(.A(mul64[10]), .Z(n_29963));
	notech_inv i_33933(.A(\opa_1[10] ), .Z(n_29964));
	notech_inv i_33934(.A(n_10911), .Z(n_29965));
	notech_inv i_33935(.A(mul64[11]), .Z(n_29966));
	notech_inv i_33936(.A(\opa_1[11] ), .Z(n_29968));
	notech_inv i_33939(.A(n_10912), .Z(n_29969));
	notech_inv i_33940(.A(mul64[12]), .Z(n_29970));
	notech_inv i_33941(.A(\opa_1[12] ), .Z(n_29971));
	notech_inv i_33942(.A(n_10913), .Z(n_29972));
	notech_inv i_33943(.A(mul64[13]), .Z(n_29973));
	notech_inv i_33944(.A(\opa_1[13] ), .Z(n_29974));
	notech_inv i_33945(.A(n_10914), .Z(n_29975));
	notech_inv i_33946(.A(mul64[14]), .Z(n_29976));
	notech_inv i_33947(.A(\opa_1[14] ), .Z(n_29977));
	notech_inv i_33948(.A(n_10915), .Z(n_29978));
	notech_inv i_33949(.A(mul64[15]), .Z(n_29979));
	notech_inv i_33950(.A(\opa_1[15] ), .Z(n_29980));
	notech_inv i_33951(.A(n_10916), .Z(n_29981));
	notech_inv i_33952(.A(n_10917), .Z(n_29982));
	notech_inv i_33953(.A(mul64[16]), .Z(n_29983));
	notech_inv i_33954(.A(n_10918), .Z(n_29985));
	notech_inv i_33955(.A(mul64[17]), .Z(n_29986));
	notech_inv i_33956(.A(n_10919), .Z(n_29987));
	notech_inv i_33957(.A(mul64[18]), .Z(n_29988));
	notech_inv i_33958(.A(n_10920), .Z(n_29991));
	notech_inv i_33959(.A(mul64[19]), .Z(n_29994));
	notech_inv i_33960(.A(n_10921), .Z(n_29995));
	notech_inv i_33961(.A(mul64[20]), .Z(n_29996));
	notech_inv i_33962(.A(n_10922), .Z(n_29997));
	notech_inv i_33963(.A(mul64[21]), .Z(n_29998));
	notech_inv i_33964(.A(n_10923), .Z(n_29999));
	notech_inv i_33965(.A(mul64[22]), .Z(n_30000));
	notech_inv i_33966(.A(n_10924), .Z(n_30001));
	notech_inv i_33967(.A(mul64[23]), .Z(n_30002));
	notech_inv i_33968(.A(n_10925), .Z(n_30003));
	notech_inv i_33969(.A(mul64[24]), .Z(n_30004));
	notech_inv i_33970(.A(n_10926), .Z(n_30005));
	notech_inv i_33971(.A(mul64[25]), .Z(n_30006));
	notech_inv i_33972(.A(n_10927), .Z(n_30007));
	notech_inv i_33973(.A(mul64[26]), .Z(n_30008));
	notech_inv i_33974(.A(n_10928), .Z(n_30009));
	notech_inv i_33975(.A(mul64[27]), .Z(n_30010));
	notech_inv i_33976(.A(n_10929), .Z(n_30011));
	notech_inv i_33977(.A(mul64[28]), .Z(n_30012));
	notech_inv i_33978(.A(n_10930), .Z(n_30013));
	notech_inv i_33979(.A(mul64[29]), .Z(n_30014));
	notech_inv i_33980(.A(n_10931), .Z(n_30015));
	notech_inv i_33981(.A(mul64[30]), .Z(n_30016));
	notech_inv i_33982(.A(mul64[31]), .Z(n_30017));
	notech_inv i_33983(.A(nbus_11317_2100235), .Z(\nbus_11317[2] ));
	notech_inv i_33984(.A(n_9224), .Z(n_30019));
	notech_inv i_33985(.A(n_9225), .Z(n_30020));
	notech_inv i_33986(.A(n_9226), .Z(n_30021));
	notech_inv i_33987(.A(n_9219), .Z(n_30022));
	notech_inv i_33988(.A(n_9220), .Z(n_30023));
	notech_inv i_33989(.A(n_9221), .Z(n_30024));
	notech_inv i_33990(.A(n_349680997100234), .Z(n_349680997));
	notech_inv i_33991(.A(n_9214), .Z(n_30026));
	notech_inv i_33992(.A(n_9215), .Z(n_30027));
	notech_inv i_33993(.A(n_9216), .Z(n_30029));
	notech_inv i_33994(.A(n_11434), .Z(n_30031));
	notech_inv i_33995(.A(n_11403), .Z(n_30032));
	notech_inv i_33996(.A(n_9324), .Z(n_30033));
	notech_inv i_33997(.A(n_9325), .Z(n_30034));
	notech_inv i_33998(.A(n_9326), .Z(n_30035));
	notech_inv i_33999(.A(n_9289), .Z(n_30036));
	notech_inv i_34000(.A(n_9290), .Z(n_30037));
	notech_inv i_34001(.A(n_9291), .Z(n_30039));
	notech_inv i_34002(.A(n_9284), .Z(n_30040));
	notech_inv i_34003(.A(n_9285), .Z(n_30041));
	notech_inv i_34004(.A(n_9286), .Z(n_30042));
	notech_inv i_34005(.A(n_9279), .Z(n_30043));
	notech_inv i_34006(.A(n_9280), .Z(n_30044));
	notech_inv i_34007(.A(n_9281), .Z(n_30045));
	notech_inv i_34008(.A(n_9274), .Z(n_30046));
	notech_inv i_34009(.A(n_9275), .Z(n_30047));
	notech_inv i_34010(.A(n_9276), .Z(n_30048));
	notech_inv i_34011(.A(n_9269), .Z(n_30050));
	notech_inv i_34012(.A(n_9270), .Z(n_30051));
	notech_inv i_34013(.A(n_9271), .Z(n_30052));
	notech_inv i_34014(.A(n_9259), .Z(n_30053));
	notech_inv i_34015(.A(n_9260), .Z(n_30054));
	notech_inv i_34016(.A(n_9261), .Z(n_30055));
	notech_inv i_34017(.A(n_9254), .Z(n_30056));
	notech_inv i_34018(.A(n_9255), .Z(n_30057));
	notech_inv i_34019(.A(n_9256), .Z(n_30058));
	notech_inv i_34020(.A(n_9249), .Z(n_30059));
	notech_inv i_34021(.A(n_9250), .Z(n_30060));
	notech_inv i_34022(.A(n_9251), .Z(n_30061));
	notech_inv i_34023(.A(n_9244), .Z(n_30062));
	notech_inv i_34024(.A(n_9245), .Z(n_30063));
	notech_inv i_34025(.A(n_9246), .Z(n_30064));
	notech_inv i_34026(.A(n_9340), .Z(n_30065));
	notech_inv i_34027(.A(n_9339), .Z(n_30066));
	notech_inv i_34028(.A(n_9341), .Z(n_30067));
	notech_inv i_34029(.A(\nbus_11317[25] ), .Z(n_30068));
	notech_inv i_34030(.A(n_9345), .Z(n_30070));
	notech_inv i_34031(.A(n_9344), .Z(n_30071));
	notech_inv i_34032(.A(n_9346), .Z(n_30072));
	notech_inv i_34033(.A(\nbus_11317[26] ), .Z(n_30073));
	notech_inv i_34034(.A(n_9365), .Z(n_30074));
	notech_inv i_34035(.A(n_9364), .Z(n_30075));
	notech_inv i_34036(.A(n_9366), .Z(n_30076));
	notech_inv i_34037(.A(\nbus_11317[30] ), .Z(n_30077));
	notech_inv i_34038(.A(n_9372), .Z(n_30078));
	notech_inv i_34039(.A(n_9371), .Z(n_30079));
	notech_inv i_34040(.A(n_8149), .Z(n_30080));
	notech_inv i_34041(.A(n_11279), .Z(n_30081));
	notech_inv i_34042(.A(n_9870), .Z(n_30082));
	notech_inv i_34043(.A(n_11281), .Z(n_30083));
	notech_inv i_34044(.A(n_9871), .Z(n_30084));
	notech_inv i_34045(.A(n_11283), .Z(n_30085));
	notech_inv i_34046(.A(n_9872), .Z(n_30086));
	notech_inv i_34047(.A(n_11285), .Z(n_30087));
	notech_inv i_34048(.A(n_9873), .Z(n_30089));
	notech_inv i_34049(.A(n_11287), .Z(n_30090));
	notech_inv i_34050(.A(n_9874), .Z(n_30091));
	notech_inv i_34051(.A(n_11289), .Z(n_30092));
	notech_inv i_34052(.A(n_9875), .Z(n_30093));
	notech_inv i_34053(.A(n_11291), .Z(n_30094));
	notech_inv i_34054(.A(n_9876), .Z(n_30095));
	notech_inv i_34055(.A(n_11293), .Z(n_30096));
	notech_inv i_34057(.A(n_9877), .Z(n_30097));
	notech_inv i_34058(.A(n_11311), .Z(n_30098));
	notech_inv i_34059(.A(n_9886), .Z(n_30099));
	notech_inv i_34060(.A(n_9351), .Z(n_30101));
	notech_inv i_34061(.A(n_9349), .Z(n_30102));
	notech_inv i_34062(.A(n_9350), .Z(n_30103));
	notech_inv i_34063(.A(n_9266), .Z(n_30104));
	notech_inv i_34064(.A(n_11317), .Z(n_30105));
	notech_inv i_34065(.A(n_9889), .Z(n_30106));
	notech_inv i_34066(.A(n_11318), .Z(n_30107));
	notech_inv i_34070(.A(n_11315), .Z(n_30108));
	notech_inv i_34071(.A(n_9888), .Z(n_30110));
	notech_inv i_34072(.A(n_11316), .Z(n_30111));
	notech_inv i_34073(.A(n_11307), .Z(n_30112));
	notech_inv i_34074(.A(n_9884), .Z(n_30113));
	notech_inv i_34075(.A(n_11308), .Z(n_30114));
	notech_inv i_34076(.A(n_11305), .Z(n_30115));
	notech_inv i_34077(.A(n_9883), .Z(n_30116));
	notech_inv i_34078(.A(n_11306), .Z(n_30117));
	notech_inv i_34079(.A(n_11303), .Z(n_30118));
	notech_inv i_34080(.A(n_9882), .Z(n_30119));
	notech_inv i_34081(.A(n_11304), .Z(n_30120));
	notech_inv i_34082(.A(n_11301), .Z(n_30121));
	notech_inv i_34083(.A(n_9881), .Z(n_30122));
	notech_inv i_34084(.A(n_11302), .Z(n_30125));
	notech_inv i_34085(.A(n_11299), .Z(n_30127));
	notech_inv i_34086(.A(n_9880), .Z(n_30128));
	notech_inv i_34087(.A(n_11300), .Z(n_30129));
	notech_inv i_34088(.A(n_11297), .Z(n_30130));
	notech_inv i_34089(.A(n_9879), .Z(n_30131));
	notech_inv i_34090(.A(n_11298), .Z(n_30132));
	notech_inv i_34091(.A(n_11295), .Z(n_30133));
	notech_inv i_34092(.A(n_9878), .Z(n_30136));
	notech_inv i_34093(.A(n_11296), .Z(n_30137));
	notech_inv i_34094(.A(n_11275), .Z(n_30139));
	notech_inv i_34095(.A(n_9868), .Z(n_30140));
	notech_inv i_34096(.A(n_11276), .Z(n_30144));
	notech_inv i_3409795650(.A(n_11273), .Z(n_30145));
	notech_inv i_34098(.A(n_9867), .Z(n_30146));
	notech_inv i_34099(.A(n_11274), .Z(n_30147));
	notech_inv i_34100(.A(n_11271), .Z(n_30148));
	notech_inv i_34101(.A(n_9866), .Z(n_30149));
	notech_inv i_3410295649(.A(n_11272), .Z(n_30150));
	notech_inv i_34103(.A(n_11269), .Z(n_30151));
	notech_inv i_34104(.A(n_9865), .Z(n_30152));
	notech_inv i_34105(.A(n_11270), .Z(n_30153));
	notech_inv i_34106(.A(n_11267), .Z(n_30154));
	notech_inv i_3410795648(.A(n_9864), .Z(n_30155));
	notech_inv i_34108(.A(n_11268), .Z(n_30156));
	notech_inv i_34109(.A(n_11265), .Z(n_30157));
	notech_inv i_34110(.A(n_9863), .Z(n_30158));
	notech_inv i_34111(.A(n_11266), .Z(n_30159));
	notech_inv i_3411295647(.A(n_11263), .Z(n_30160));
	notech_inv i_34113(.A(n_9862), .Z(n_30161));
	notech_inv i_34114(.A(n_11264), .Z(n_30162));
	notech_inv i_34115(.A(n_11261), .Z(n_30163));
	notech_inv i_34116(.A(n_9861), .Z(n_30164));
	notech_inv i_3411795646(.A(n_11262), .Z(n_30165));
	notech_inv i_34118(.A(n_11259), .Z(n_30166));
	notech_inv i_34119(.A(n_9860), .Z(n_30167));
	notech_inv i_34120(.A(n_11260), .Z(n_30168));
	notech_inv i_34121(.A(\opc_5[8] ), .Z(n_30169));
	notech_inv i_3412295645(.A(n_8299), .Z(n_30170));
	notech_inv i_34123(.A(mul64[40]), .Z(n_30171));
	notech_inv i_34124(.A(mul64[63]), .Z(n_30172));
	notech_inv i_34125(.A(mul64[62]), .Z(n_30173));
	notech_inv i_34126(.A(mul64[61]), .Z(n_30174));
	notech_inv i_34127(.A(mul64[60]), .Z(n_30175));
	notech_inv i_34128(.A(mul64[59]), .Z(n_30176));
	notech_inv i_34129(.A(mul64[58]), .Z(n_30177));
	notech_inv i_34130(.A(mul64[57]), .Z(n_30178));
	notech_inv i_34131(.A(mul64[56]), .Z(n_30179));
	notech_inv i_34132(.A(mul64[55]), .Z(n_30180));
	notech_inv i_34133(.A(mul64[54]), .Z(n_30181));
	notech_inv i_34134(.A(mul64[53]), .Z(n_30182));
	notech_inv i_34135(.A(mul64[52]), .Z(n_30183));
	notech_inv i_34136(.A(mul64[51]), .Z(n_30184));
	notech_inv i_34138(.A(mul64[50]), .Z(n_30185));
	notech_inv i_34139(.A(mul64[49]), .Z(n_30186));
	notech_inv i_34140(.A(mul64[48]), .Z(n_30187));
	notech_inv i_34141(.A(mul64[47]), .Z(n_30188));
	notech_inv i_34142(.A(mul64[46]), .Z(n_30189));
	notech_inv i_34143(.A(mul64[45]), .Z(n_30190));
	notech_inv i_34144(.A(mul64[44]), .Z(n_30191));
	notech_inv i_34147(.A(mul64[43]), .Z(n_30192));
	notech_inv i_34148(.A(mul64[42]), .Z(n_30193));
	notech_inv i_34150(.A(mul64[41]), .Z(n_30194));
	notech_inv i_34151(.A(mul64[36]), .Z(n_30195));
	notech_inv i_34152(.A(mul64[35]), .Z(n_30196));
	notech_inv i_34153(.A(mul64[34]), .Z(n_30197));
	notech_inv i_34155(.A(mul64[33]), .Z(n_30198));
	notech_inv i_34156(.A(mul64[32]), .Z(n_30199));
	notech_inv i_34157(.A(mul64[39]), .Z(n_30200));
	notech_inv i_34158(.A(n_5185), .Z(n_30201));
	notech_inv i_34159(.A(n_5180), .Z(n_30202));
	notech_inv i_34160(.A(n_9359), .Z(n_30203));
	notech_inv i_34161(.A(n_9360), .Z(n_30204));
	notech_inv i_34162(.A(n_9361), .Z(n_30205));
	notech_inv i_34163(.A(n_9354), .Z(n_30206));
	notech_inv i_34164(.A(n_9355), .Z(n_30207));
	notech_inv i_34165(.A(n_9356), .Z(n_30208));
	notech_inv i_34166(.A(n_9334), .Z(n_30209));
	notech_inv i_34167(.A(n_9335), .Z(n_30210));
	notech_inv i_34168(.A(n_9336), .Z(n_30211));
	notech_inv i_34169(.A(n_9329), .Z(n_30212));
	notech_inv i_34170(.A(n_9330), .Z(n_30213));
	notech_inv i_34171(.A(n_9331), .Z(n_30214));
	notech_inv i_34172(.A(n_9319), .Z(n_30215));
	notech_inv i_34173(.A(n_9320), .Z(n_30216));
	notech_inv i_34174(.A(n_9321), .Z(n_30217));
	notech_inv i_34175(.A(n_9314), .Z(n_30218));
	notech_inv i_34176(.A(n_9315), .Z(n_30219));
	notech_inv i_34177(.A(n_9316), .Z(n_30220));
	notech_inv i_34178(.A(n_9309), .Z(n_30221));
	notech_inv i_34179(.A(n_9310), .Z(n_30222));
	notech_inv i_34180(.A(n_9311), .Z(n_30223));
	notech_inv i_34181(.A(n_9304), .Z(n_30224));
	notech_inv i_34182(.A(n_9305), .Z(n_30225));
	notech_inv i_34183(.A(n_9306), .Z(n_30226));
	notech_inv i_34184(.A(n_9299), .Z(n_30227));
	notech_inv i_34185(.A(n_9300), .Z(n_30228));
	notech_inv i_34186(.A(n_9301), .Z(n_30229));
	notech_inv i_34187(.A(n_9294), .Z(n_30230));
	notech_inv i_34188(.A(n_9295), .Z(n_30231));
	notech_inv i_34189(.A(n_9296), .Z(n_30232));
	notech_inv i_34190(.A(n_130392201), .Z(n_30233));
	notech_inv i_34191(.A(n_8130), .Z(n_30234));
	notech_inv i_34192(.A(n_8131), .Z(n_30235));
	notech_inv i_34193(.A(n_8132), .Z(n_30236));
	notech_inv i_34194(.A(n_8133), .Z(n_30237));
	notech_inv i_34195(.A(n_8134), .Z(n_30238));
	notech_inv i_34196(.A(n_8135), .Z(n_30239));
	notech_inv i_34197(.A(n_8136), .Z(n_30240));
	notech_inv i_34198(.A(n_8137), .Z(n_30241));
	notech_inv i_34199(.A(n_8138), .Z(n_30242));
	notech_inv i_34200(.A(n_8139), .Z(n_30243));
	notech_inv i_34201(.A(n_8140), .Z(n_30245));
	notech_inv i_34202(.A(n_8141), .Z(n_30247));
	notech_inv i_34203(.A(n_8142), .Z(n_30248));
	notech_inv i_34204(.A(n_8143), .Z(n_30249));
	notech_inv i_34205(.A(n_8144), .Z(n_30250));
	notech_inv i_34206(.A(n_8145), .Z(n_30252));
	notech_inv i_34207(.A(n_8146), .Z(n_30253));
	notech_inv i_34208(.A(n_8147), .Z(n_30255));
	notech_inv i_34209(.A(n_8148), .Z(n_30257));
	notech_inv i_34210(.A(n_8150), .Z(n_30259));
	notech_inv i_34211(.A(n_8151), .Z(n_30260));
	notech_inv i_34212(.A(n_8152), .Z(n_30262));
	notech_inv i_34213(.A(n_8153), .Z(n_30263));
	notech_inv i_34214(.A(n_8154), .Z(n_30265));
	notech_inv i_34215(.A(n_8155), .Z(n_30267));
	notech_inv i_34216(.A(n_8156), .Z(n_30271));
	notech_inv i_34217(.A(n_8157), .Z(n_30275));
	notech_inv i_34218(.A(n_8158), .Z(n_30276));
	notech_inv i_34219(.A(n_8159), .Z(n_30277));
	notech_inv i_34220(.A(n_8160), .Z(n_30279));
	notech_inv i_34221(.A(n_8161), .Z(n_30280));
	notech_inv i_34222(.A(n_8162), .Z(n_30281));
	notech_inv i_34223(.A(n_8163), .Z(n_30282));
	notech_inv i_34224(.A(n_8164), .Z(n_30283));
	notech_inv i_34225(.A(n_8165), .Z(n_30284));
	notech_inv i_34226(.A(n_8166), .Z(n_30285));
	notech_inv i_34227(.A(n_8167), .Z(n_30286));
	notech_inv i_34228(.A(n_8168), .Z(n_30287));
	notech_inv i_34229(.A(n_8169), .Z(n_30288));
	notech_inv i_34230(.A(n_8170), .Z(n_30289));
	notech_inv i_34231(.A(n_8171), .Z(n_30291));
	notech_inv i_34232(.A(n_8172), .Z(n_30292));
	notech_inv i_34233(.A(n_8173), .Z(n_30293));
	notech_inv i_34234(.A(n_8174), .Z(n_30295));
	notech_inv i_34235(.A(n_8175), .Z(n_30296));
	notech_inv i_34236(.A(n_8176), .Z(n_30297));
	notech_inv i_34237(.A(n_8177), .Z(n_30298));
	notech_inv i_34238(.A(n_8178), .Z(n_30302));
	notech_inv i_34239(.A(n_8179), .Z(n_30304));
	notech_inv i_34240(.A(n_8180), .Z(n_30307));
	notech_inv i_34241(.A(n_8181), .Z(n_30308));
	notech_inv i_34242(.A(n_8182), .Z(n_30309));
	notech_inv i_34244(.A(n_8183), .Z(n_30313));
	notech_inv i_34245(.A(n_8184), .Z(n_30314));
	notech_inv i_34247(.A(n_8185), .Z(n_30316));
	notech_inv i_34248(.A(n_8186), .Z(n_30317));
	notech_inv i_34249(.A(n_8187), .Z(n_30318));
	notech_inv i_34250(.A(n_8188), .Z(n_30319));
	notech_inv i_34251(.A(n_8189), .Z(n_30320));
	notech_inv i_34252(.A(n_8190), .Z(n_30321));
	notech_inv i_34253(.A(n_8191), .Z(n_30323));
	notech_inv i_34254(.A(n_8192), .Z(n_30324));
	notech_inv i_34255(.A(n_8193), .Z(n_30326));
	notech_inv i_34256(.A(n_8194), .Z(n_30327));
	notech_inv i_34257(.A(n_8195), .Z(n_30330));
	notech_inv i_34259(.A(n_8196), .Z(n_30331));
	notech_inv i_34260(.A(n_8197), .Z(n_30333));
	notech_inv i_34261(.A(n_8198), .Z(n_30334));
	notech_inv i_34262(.A(n_8199), .Z(n_30335));
	notech_inv i_34263(.A(n_8200), .Z(n_30336));
	notech_inv i_34266(.A(n_8201), .Z(n_30337));
	notech_inv i_34267(.A(n_8202), .Z(n_30338));
	notech_inv i_34268(.A(n_8203), .Z(n_30339));
	notech_inv i_34269(.A(n_8204), .Z(n_30340));
	notech_inv i_34270(.A(n_8205), .Z(n_30341));
	notech_inv i_34271(.A(n_8206), .Z(n_30343));
	notech_inv i_34272(.A(n_8207), .Z(n_30345));
	notech_inv i_34273(.A(n_8208), .Z(n_30346));
	notech_inv i_34274(.A(n_8209), .Z(n_30347));
	notech_inv i_34275(.A(n_8210), .Z(n_30348));
	notech_inv i_34276(.A(n_8211), .Z(n_30349));
	notech_inv i_34277(.A(n_8212), .Z(n_30351));
	notech_inv i_34278(.A(n_8213), .Z(n_30353));
	notech_inv i_34279(.A(n_8214), .Z(n_30354));
	notech_inv i_34280(.A(n_8215), .Z(n_30355));
	notech_inv i_34281(.A(n_8216), .Z(n_30356));
	notech_inv i_34282(.A(n_8217), .Z(n_30358));
	notech_inv i_34283(.A(n_8218), .Z(n_30360));
	notech_inv i_34284(.A(n_8219), .Z(n_30362));
	notech_inv i_34286(.A(n_8220), .Z(n_30363));
	notech_inv i_34288(.A(n_8221), .Z(n_30364));
	notech_inv i_34289(.A(n_8222), .Z(n_30367));
	notech_inv i_34290(.A(n_8223), .Z(n_30368));
	notech_inv i_34291(.A(n_8224), .Z(n_30369));
	notech_inv i_34292(.A(n_8225), .Z(n_30371));
	notech_inv i_34293(.A(n_8226), .Z(n_30372));
	notech_inv i_34294(.A(n_9858), .Z(n_30373));
	notech_inv i_34295(.A(n_9859), .Z(n_30375));
	notech_inv i_34296(.A(n_11258), .Z(n_30376));
	notech_inv i_34297(.A(n_8291), .Z(n_30377));
	notech_inv i_34298(.A(n_8324), .Z(n_30378));
	notech_inv i_34299(.A(n_8292), .Z(n_30379));
	notech_inv i_34300(.A(n_8325), .Z(n_30380));
	notech_inv i_34301(.A(\opc_1[1] ), .Z(n_30381));
	notech_inv i_34302(.A(n_8293), .Z(n_30382));
	notech_inv i_34303(.A(\opc_1[2] ), .Z(n_30383));
	notech_inv i_34304(.A(n_8326), .Z(n_30384));
	notech_inv i_34305(.A(n_8294), .Z(n_30385));
	notech_inv i_34306(.A(n_8327), .Z(n_30386));
	notech_inv i_34307(.A(n_8295), .Z(n_30388));
	notech_inv i_34308(.A(n_8328), .Z(n_30390));
	notech_inv i_34309(.A(\opc_1[4] ), .Z(n_30391));
	notech_inv i_34310(.A(\opc_5[9] ), .Z(n_30392));
	notech_inv i_34311(.A(n_8300), .Z(n_30393));
	notech_inv i_34312(.A(\opc_5[10] ), .Z(n_30394));
	notech_inv i_34313(.A(n_8301), .Z(n_30395));
	notech_inv i_34314(.A(\opc_5[11] ), .Z(n_30396));
	notech_inv i_34315(.A(n_8302), .Z(n_30397));
	notech_inv i_34316(.A(\opc_5[12] ), .Z(n_30398));
	notech_inv i_34317(.A(n_8303), .Z(n_30399));
	notech_inv i_34318(.A(\opc_5[13] ), .Z(n_30400));
	notech_inv i_34319(.A(n_8304), .Z(n_30401));
	notech_inv i_34320(.A(\opc_5[14] ), .Z(n_30402));
	notech_inv i_34321(.A(n_8305), .Z(n_30403));
	notech_inv i_34322(.A(n_8306), .Z(n_30404));
	notech_inv i_34323(.A(\opc_5[15] ), .Z(n_30405));
	notech_inv i_34324(.A(n_8307), .Z(n_30406));
	notech_inv i_34325(.A(\opc_5[16] ), .Z(n_30407));
	notech_inv i_34326(.A(n_8308), .Z(n_30408));
	notech_inv i_34327(.A(\opc_5[17] ), .Z(n_30409));
	notech_inv i_34328(.A(n_8309), .Z(n_30410));
	notech_inv i_34329(.A(\opc_5[18] ), .Z(n_30411));
	notech_inv i_34330(.A(n_8310), .Z(n_30412));
	notech_inv i_34331(.A(\opc_5[19] ), .Z(n_30413));
	notech_inv i_34332(.A(n_8311), .Z(n_30414));
	notech_inv i_34333(.A(\opc_5[20] ), .Z(n_30416));
	notech_inv i_34334(.A(n_8312), .Z(n_30417));
	notech_inv i_34335(.A(\opc_5[21] ), .Z(n_30418));
	notech_inv i_34336(.A(n_8313), .Z(n_30419));
	notech_inv i_34337(.A(\opc_5[22] ), .Z(n_30420));
	notech_inv i_34338(.A(n_8314), .Z(n_30421));
	notech_inv i_34339(.A(\opc_5[23] ), .Z(n_30422));
	notech_inv i_34340(.A(n_8315), .Z(n_30423));
	notech_inv i_34341(.A(\opc_5[24] ), .Z(n_30424));
	notech_inv i_34342(.A(n_8316), .Z(n_30425));
	notech_inv i_34343(.A(\opc_5[25] ), .Z(n_30426));
	notech_inv i_34344(.A(n_8317), .Z(n_30427));
	notech_inv i_34345(.A(\opc_5[26] ), .Z(n_30428));
	notech_inv i_34346(.A(n_8318), .Z(n_30429));
	notech_inv i_34347(.A(\opc_5[27] ), .Z(n_30430));
	notech_inv i_34348(.A(n_8319), .Z(n_30431));
	notech_inv i_34349(.A(\opc_5[28] ), .Z(n_30432));
	notech_inv i_34350(.A(n_8320), .Z(n_30433));
	notech_inv i_34351(.A(\opc_5[29] ), .Z(n_30434));
	notech_inv i_34352(.A(n_8321), .Z(n_30435));
	notech_inv i_34353(.A(\opc_5[30] ), .Z(n_30436));
	notech_inv i_34354(.A(n_8322), .Z(n_30437));
	notech_inv i_34355(.A(\opc_5[31] ), .Z(n_30438));
	notech_inv i_34356(.A(\opc_1[5] ), .Z(n_30439));
	notech_inv i_34357(.A(\opc_5[5] ), .Z(n_30440));
	notech_inv i_34358(.A(n_8296), .Z(n_30441));
	notech_inv i_34359(.A(\opc_1[6] ), .Z(n_30443));
	notech_inv i_34360(.A(\opc_5[6] ), .Z(n_30444));
	notech_inv i_34361(.A(n_8297), .Z(n_30445));
	notech_inv i_34362(.A(n_9869), .Z(n_30446));
	notech_inv i_34363(.A(n_5227), .Z(n_30448));
	notech_inv i_34364(.A(n_8298), .Z(n_30449));
	notech_inv i_34365(.A(\opc_5[7] ), .Z(n_30450));
	notech_inv i_34366(.A(\opc_1[7] ), .Z(n_30452));
	notech_inv i_34367(.A(n_11188), .Z(n_30453));
	notech_inv i_34368(.A(n_11187), .Z(n_30454));
	notech_inv i_34369(.A(n_11186), .Z(n_30456));
	notech_inv i_34370(.A(n_11184), .Z(n_30457));
	notech_inv i_34371(.A(n_11183), .Z(n_30458));
	notech_inv i_34372(.A(n_11182), .Z(n_30460));
	notech_inv i_34373(.A(n_11181), .Z(n_30462));
	notech_inv i_34374(.A(n_11180), .Z(n_30463));
	notech_inv i_34375(.A(n_11179), .Z(n_30465));
	notech_inv i_34376(.A(n_11178), .Z(n_30467));
	notech_inv i_34377(.A(n_11177), .Z(n_30468));
	notech_inv i_34378(.A(n_11176), .Z(n_30469));
	notech_inv i_34379(.A(n_11175), .Z(n_30471));
	notech_inv i_34380(.A(n_11174), .Z(n_30473));
	notech_inv i_34381(.A(n_11173), .Z(n_30474));
	notech_inv i_34382(.A(n_11172), .Z(n_30476));
	notech_inv i_34383(.A(n_11171), .Z(n_30477));
	notech_inv i_34384(.A(n_11170), .Z(n_30478));
	notech_inv i_34385(.A(n_11169), .Z(n_30479));
	notech_inv i_34386(.A(n_11168), .Z(n_30480));
	notech_inv i_34387(.A(n_11167), .Z(n_30482));
	notech_inv i_34388(.A(n_11166), .Z(n_30483));
	notech_inv i_34389(.A(n_11165), .Z(n_30484));
	notech_inv i_34390(.A(n_11164), .Z(n_30485));
	notech_inv i_34391(.A(n_11163), .Z(n_30486));
	notech_inv i_34392(.A(n_11162), .Z(n_30487));
	notech_inv i_34393(.A(n_11161), .Z(n_30488));
	notech_inv i_34394(.A(n_11160), .Z(n_30489));
	notech_inv i_34395(.A(n_11159), .Z(n_30490));
	notech_inv i_34396(.A(n_11158), .Z(n_30491));
	notech_inv i_34397(.A(n_11157), .Z(n_30492));
	notech_inv i_34398(.A(n_11156), .Z(n_30493));
	notech_inv i_34399(.A(n_11155), .Z(n_30494));
	notech_inv i_34400(.A(n_11154), .Z(n_30495));
	notech_inv i_34401(.A(n_11153), .Z(n_30496));
	notech_inv i_34402(.A(n_11152), .Z(n_30498));
	notech_inv i_34403(.A(n_11151), .Z(n_30499));
	notech_inv i_34404(.A(n_11150), .Z(n_30500));
	notech_inv i_34405(.A(n_11149), .Z(n_30501));
	notech_inv i_34406(.A(n_11148), .Z(n_30502));
	notech_inv i_34407(.A(n_11147), .Z(n_30503));
	notech_inv i_34408(.A(n_11146), .Z(n_30504));
	notech_inv i_34409(.A(n_11145), .Z(n_30505));
	notech_inv i_34410(.A(n_11144), .Z(n_30506));
	notech_inv i_34411(.A(n_11143), .Z(n_30507));
	notech_inv i_34412(.A(n_11142), .Z(n_30508));
	notech_inv i_34413(.A(n_11141), .Z(n_30509));
	notech_inv i_34414(.A(n_11140), .Z(n_30510));
	notech_inv i_34415(.A(n_11139), .Z(n_30511));
	notech_inv i_34416(.A(n_11138), .Z(n_30512));
	notech_inv i_34417(.A(n_11137), .Z(n_30513));
	notech_inv i_34418(.A(n_11136), .Z(n_30514));
	notech_inv i_34419(.A(n_11135), .Z(n_30515));
	notech_inv i_34420(.A(n_11134), .Z(n_30516));
	notech_inv i_34421(.A(n_11133), .Z(n_30517));
	notech_inv i_34422(.A(n_11132), .Z(n_30518));
	notech_inv i_34423(.A(n_11131), .Z(n_30519));
	notech_inv i_34424(.A(n_11130), .Z(n_30520));
	notech_inv i_34425(.A(n_11129), .Z(n_30521));
	notech_inv i_34426(.A(n_11128), .Z(n_30522));
	notech_inv i_34427(.A(n_11127), .Z(n_30523));
	notech_inv i_34428(.A(n_11126), .Z(n_30524));
	notech_inv i_34429(.A(n_11125), .Z(n_30525));
	notech_inv i_34430(.A(n_11114), .Z(n_30526));
	notech_inv i_34431(.A(n_11113), .Z(n_30527));
	notech_inv i_34432(.A(n_11091), .Z(n_30529));
	notech_inv i_34433(.A(n_11090), .Z(n_30530));
	notech_inv i_34434(.A(n_11089), .Z(n_30531));
	notech_inv i_34435(.A(n_11088), .Z(n_30532));
	notech_inv i_34436(.A(n_11087), .Z(n_30533));
	notech_inv i_34437(.A(n_11086), .Z(n_30534));
	notech_inv i_34438(.A(n_11085), .Z(n_30535));
	notech_inv i_34439(.A(n_11084), .Z(n_30536));
	notech_inv i_34440(.A(n_11083), .Z(n_30537));
	notech_inv i_34441(.A(n_11082), .Z(n_30538));
	notech_inv i_34442(.A(n_11081), .Z(n_30539));
	notech_inv i_34443(.A(n_11080), .Z(n_30540));
	notech_inv i_34444(.A(n_11079), .Z(n_30541));
	notech_inv i_34445(.A(n_11078), .Z(n_30542));
	notech_inv i_34446(.A(n_11077), .Z(n_30543));
	notech_inv i_34447(.A(n_11076), .Z(n_30544));
	notech_inv i_34448(.A(n_11075), .Z(n_30545));
	notech_inv i_34449(.A(n_11074), .Z(n_30546));
	notech_inv i_34450(.A(n_11073), .Z(n_30547));
	notech_inv i_34451(.A(n_11072), .Z(n_30548));
	notech_inv i_34452(.A(n_11069), .Z(n_30549));
	notech_inv i_34453(.A(n_11062), .Z(n_30550));
	notech_inv i_34454(.A(n_11061), .Z(n_30551));
	notech_inv i_34455(.A(n_11220), .Z(n_30552));
	notech_inv i_34456(.A(n_11219), .Z(n_30553));
	notech_inv i_34457(.A(n_11218), .Z(n_30554));
	notech_inv i_34458(.A(n_11217), .Z(n_30555));
	notech_inv i_34459(.A(n_11216), .Z(n_30556));
	notech_inv i_34460(.A(n_11215), .Z(n_30557));
	notech_inv i_34461(.A(n_11214), .Z(n_30558));
	notech_inv i_34462(.A(n_11213), .Z(n_30559));
	notech_inv i_34463(.A(n_11212), .Z(n_30560));
	notech_inv i_34464(.A(n_11211), .Z(n_30561));
	notech_inv i_34465(.A(n_11210), .Z(n_30562));
	notech_inv i_34466(.A(n_11209), .Z(n_30563));
	notech_inv i_34467(.A(n_11208), .Z(n_30564));
	notech_inv i_34469(.A(n_11207), .Z(n_30566));
	notech_inv i_34470(.A(n_11206), .Z(n_30567));
	notech_inv i_34471(.A(n_11205), .Z(n_30571));
	notech_inv i_34472(.A(n_11204), .Z(n_30572));
	notech_inv i_34473(.A(n_11203), .Z(n_30573));
	notech_inv i_34475(.A(n_11202), .Z(n_30574));
	notech_inv i_34476(.A(n_11201), .Z(n_30575));
	notech_inv i_34477(.A(n_11200), .Z(n_30576));
	notech_inv i_34478(.A(n_11199), .Z(n_30577));
	notech_inv i_34479(.A(n_11198), .Z(n_30578));
	notech_inv i_34480(.A(n_11197), .Z(n_30579));
	notech_inv i_34481(.A(n_11196), .Z(n_30580));
	notech_inv i_34482(.A(n_11195), .Z(n_30581));
	notech_inv i_34483(.A(n_11194), .Z(n_30585));
	notech_inv i_34485(.A(n_11193), .Z(n_30586));
	notech_inv i_34486(.A(n_11192), .Z(n_30587));
	notech_inv i_34489(.A(n_11191), .Z(n_30589));
	notech_inv i_34490(.A(n_11190), .Z(n_30590));
	notech_inv i_34491(.A(n_11189), .Z(n_30591));
	notech_inv i_34492(.A(n_11124), .Z(n_30592));
	notech_inv i_34493(.A(n_11123), .Z(n_30593));
	notech_inv i_34494(.A(n_11122), .Z(n_30595));
	notech_inv i_34495(.A(n_11121), .Z(n_30596));
	notech_inv i_34496(.A(n_11120), .Z(n_30597));
	notech_inv i_34497(.A(n_11119), .Z(n_30599));
	notech_inv i_34498(.A(n_11118), .Z(n_30600));
	notech_inv i_34499(.A(n_11117), .Z(n_30601));
	notech_inv i_34500(.A(n_11116), .Z(n_30602));
	notech_inv i_34501(.A(n_11115), .Z(n_30603));
	notech_inv i_34502(.A(n_11112), .Z(n_30604));
	notech_inv i_34503(.A(n_11111), .Z(n_30605));
	notech_inv i_34504(.A(n_11110), .Z(n_30608));
	notech_inv i_34505(.A(n_11109), .Z(n_30609));
	notech_inv i_34506(.A(n_11108), .Z(n_30610));
	notech_inv i_34507(.A(n_11107), .Z(n_30611));
	notech_inv i_34508(.A(n_11106), .Z(n_30612));
	notech_inv i_34509(.A(n_11105), .Z(n_30613));
	notech_inv i_34510(.A(n_11104), .Z(n_30614));
	notech_inv i_34511(.A(n_11103), .Z(n_30615));
	notech_inv i_34512(.A(n_11102), .Z(n_30616));
	notech_inv i_34513(.A(n_11101), .Z(n_30617));
	notech_inv i_34514(.A(n_11100), .Z(n_30618));
	notech_inv i_34515(.A(n_11099), .Z(n_30619));
	notech_inv i_34516(.A(n_11098), .Z(n_30620));
	notech_inv i_34517(.A(n_11097), .Z(n_30621));
	notech_inv i_34518(.A(n_11096), .Z(n_30622));
	notech_inv i_34519(.A(n_11095), .Z(n_30623));
	notech_inv i_34520(.A(n_11094), .Z(n_30624));
	notech_inv i_34521(.A(n_11093), .Z(n_30625));
	notech_inv i_34522(.A(n_11092), .Z(n_30626));
	notech_inv i_34523(.A(n_11071), .Z(n_30627));
	notech_inv i_34524(.A(n_11070), .Z(n_30628));
	notech_inv i_34525(.A(n_11068), .Z(n_30629));
	notech_inv i_34526(.A(n_11067), .Z(n_30630));
	notech_inv i_34527(.A(n_11066), .Z(n_30631));
	notech_inv i_34528(.A(n_11065), .Z(n_30632));
	notech_inv i_34529(.A(n_11063), .Z(n_30633));
	notech_inv i_34530(.A(n_11185), .Z(n_30634));
	notech_inv i_34531(.A(n_60769), .Z(n_30635));
	AWMUX_16_32_7 i_34097(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14523[31] , \nbus_14523[30] , \nbus_14523[29] , \nbus_14523[28] 
		, \nbus_14523[27] , \nbus_14523[26] , \nbus_14523[25] , \nbus_14523[24] 
		, \nbus_14523[23] , \nbus_14523[22] , \nbus_14523[21] , \nbus_14523[20] 
		, \nbus_14523[19] , \nbus_14523[18] , \nbus_14523[17] , \nbus_14523[16] 
		, \nbus_14523[15] , \nbus_14523[14] , \nbus_14523[13] , \nbus_14523[12] 
		, \nbus_14523[11] , \nbus_14523[10] , \nbus_14523[9] , \nbus_14523[8] 
		, \nbus_14523[7] , \nbus_14523[6] , \nbus_14523[5] , \nbus_14523[4] 
		, \nbus_14523[3] , \nbus_14523[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_56001, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, n_56172, ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[107], n_57361, instrc[105], instrc[104]}), .O0({n_11092
		, n_11091, n_11090, n_11089, n_11088, n_11087, n_11086, n_11085,
		 n_11084, n_11083, n_11082, n_11081, n_11080, n_11079, n_11078, n_11077
		, n_11076, n_11075, n_11074, n_11073, n_11072, n_11071, n_11070,
		 n_11069, n_11068, n_11067, n_11066, n_11065, n_11064, n_11063, n_11062
		, n_11061}));
	AWMUX_16_32_6 i_34102(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14523[31] , \nbus_14523[30] , \nbus_14523[29] , \nbus_14523[28] 
		, \nbus_14523[27] , \nbus_14523[26] , \nbus_14523[25] , \nbus_14523[24] 
		, \nbus_14523[23] , \nbus_14523[22] , \nbus_14523[21] , \nbus_14523[20] 
		, \nbus_14523[19] , \nbus_14523[18] , \nbus_14523[17] , \nbus_14523[16] 
		, \nbus_14523[15] , \nbus_14523[14] , \nbus_14523[13] , \nbus_14523[12] 
		, \nbus_14523[11] , \nbus_14523[10] , \nbus_14523[9] , \nbus_14523[8] 
		, \nbus_14523[7] , \nbus_14523[6] , \nbus_14523[5] , \nbus_14523[4] 
		, \nbus_14523[3] , \nbus_14523[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_56001, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, n_56172, ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[103], instrc[102], instrc[101], instrc[100]}), .O0
		({n_11124, n_11123, n_11122, n_11121, n_11120, n_11119, n_11118,
		 n_11117, n_11116, n_11115, n_11114, n_11113, n_11112, n_11111, n_11110
		, n_11109, n_11108, n_11107, n_11106, n_11105, n_11104, n_11103,
		 n_11102, n_11101, n_11100, n_11099, n_11098, n_11097, n_11096, n_11095
		, n_11094, n_11093}));
	AWMUX_16_32_5 i_34107(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14523[31] , \nbus_14523[30] , \nbus_14523[29] , \nbus_14523[28] 
		, \nbus_14523[27] , \nbus_14523[26] , \nbus_14523[25] , \nbus_14523[24] 
		, \nbus_14523[23] , \nbus_14523[22] , \nbus_14523[21] , \nbus_14523[20] 
		, \nbus_14523[19] , \nbus_14523[18] , \nbus_14523[17] , \nbus_14523[16] 
		, \nbus_14523[15] , \nbus_14523[14] , \nbus_14523[13] , \nbus_14523[12] 
		, \nbus_14523[11] , \nbus_14523[10] , \nbus_14523[9] , \nbus_14523[8] 
		, \nbus_14523[7] , \nbus_14523[6] , \nbus_14523[5] , \nbus_14523[4] 
		, \nbus_14523[3] , \nbus_14523[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_56001, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, n_56172, ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[99], instrc[98], instrc[97], instrc[96]}), .O0({n_11156
		, n_11155, n_11154, n_11153, n_11152, n_11151, n_11150, n_11149,
		 n_11148, n_11147, n_11146, n_11145, n_11144, n_11143, n_11142, n_11141
		, n_11140, n_11139, n_11138, n_11137, n_11136, n_11135, n_11134,
		 n_11133, n_11132, n_11131, n_11130, n_11129, n_11128, n_11127, n_11126
		, n_11125}));
	AWMUX_16_32_4 i_34112(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14523[31] , \nbus_14523[30] , \nbus_14523[29] , \nbus_14523[28] 
		, \nbus_14523[27] , \nbus_14523[26] , \nbus_14523[25] , \nbus_14523[24] 
		, \nbus_14523[23] , \nbus_14523[22] , \nbus_14523[21] , \nbus_14523[20] 
		, \nbus_14523[19] , \nbus_14523[18] , \nbus_14523[17] , \nbus_14523[16] 
		, \nbus_14523[15] , \nbus_14523[14] , \nbus_14523[13] , \nbus_14523[12] 
		, \nbus_14523[11] , \nbus_14523[10] , \nbus_14523[9] , \nbus_14523[8] 
		, \nbus_14523[7] , \nbus_14523[6] , \nbus_14523[5] , \nbus_14523[4] 
		, \nbus_14523[3] , \nbus_14523[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_56001, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, n_56172, ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[95], instrc[94], instrc[93], instrc[92]}), .O0({n_11188
		, n_11187, n_11186, n_11185, n_11184, n_11183, n_11182, n_11181,
		 n_11180, n_11179, n_11178, n_11177, n_11176, n_11175, n_11174, n_11173
		, n_11172, n_11171, n_11170, n_11169, n_11168, n_11167, n_11166,
		 n_11165, n_11164, n_11163, n_11162, n_11161, n_11160, n_11159, n_11158
		, n_11157}));
	AWMUX_16_32_3 i_34117(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14523[31] , \nbus_14523[30] , \nbus_14523[29] , \nbus_14523[28] 
		, \nbus_14523[27] , \nbus_14523[26] , \nbus_14523[25] , \nbus_14523[24] 
		, \nbus_14523[23] , \nbus_14523[22] , \nbus_14523[21] , \nbus_14523[20] 
		, \nbus_14523[19] , \nbus_14523[18] , \nbus_14523[17] , \nbus_14523[16] 
		, \nbus_14523[15] , \nbus_14523[14] , \nbus_14523[13] , \nbus_14523[12] 
		, \nbus_14523[11] , \nbus_14523[10] , \nbus_14523[9] , \nbus_14523[8] 
		, \nbus_14523[7] , \nbus_14523[6] , \nbus_14523[5] , \nbus_14523[4] 
		, \nbus_14523[3] , \nbus_14523[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_56001, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, n_56172, ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[91], instrc[90], instrc[89], instrc[88]}), .O0({n_11220
		, n_11219, n_11218, n_11217, n_11216, n_11215, n_11214, n_11213,
		 n_11212, n_11211, n_11210, n_11209, n_11208, n_11207, n_11206, n_11205
		, n_11204, n_11203, n_11202, n_11201, n_11200, n_11199, n_11198,
		 n_11197, n_11196, n_11195, n_11194, n_11193, n_11192, n_11191, n_11190
		, n_11189}));
	AWMUX_16_32_2 i_34122(.I0(write_data_25), .I1(write_data_26), .I2(write_data_27
		), .I3(write_data_28), .I4(write_data_29), .I5(write_data_30), .I6
		(write_data_31), .I7(write_data_32), .S(all_cnt), .O0(write_data_33
		));
	AWMUX_16_32_1 i_56887(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14523[31] , \nbus_14523[30] , \nbus_14523[29] , \nbus_14523[28] 
		, \nbus_14523[27] , \nbus_14523[26] , \nbus_14523[25] , \nbus_14523[24] 
		, \nbus_14523[23] , \nbus_14523[22] , \nbus_14523[21] , \nbus_14523[20] 
		, \nbus_14523[19] , \nbus_14523[18] , \nbus_14523[17] , \nbus_14523[16] 
		, \nbus_14523[15] , \nbus_14523[14] , \nbus_14523[13] , \nbus_14523[12] 
		, \nbus_14523[11] , \nbus_14523[10] , \nbus_14523[9] , \nbus_14523[8] 
		, \nbus_14523[7] , \nbus_14523[6] , \nbus_14523[5] , \nbus_14523[4] 
		, \nbus_14523[3] , \nbus_14523[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_56001, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, n_56172, ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[127], instrc[126], instrc[125], instrc[124]}), .O0
		({\regs_13_14[31] , \regs_13_14[30] , \regs_13_14[29] , \regs_13_14[28] 
		, \regs_13_14[27] , \regs_13_14[26] , \regs_13_14[25] , \regs_13_14[24] 
		, \regs_13_14[23] , \regs_13_14[22] , \regs_13_14[21] , \regs_13_14[20] 
		, \regs_13_14[19] , \regs_13_14[18] , \regs_13_14[17] , \regs_13_14[16] 
		, \opa_12[15] , \opa_12[14] , \opa_12[13] , \opa_12[12] , \opa_12[11] 
		, \opa_12[10] , \opa_12[9] , \opa_12[8] , \opa_12[7] , \opa_12[6] 
		, \opa_12[5] , \opa_12[4] , \opa_12[3] , \opa_12[2] , \opa_12[1] 
		, \opa_12[0] }));
	AWMUX_16_32_0 i_57241(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14523[31] , \nbus_14523[30] , \nbus_14523[29] , \nbus_14523[28] 
		, \nbus_14523[27] , \nbus_14523[26] , \nbus_14523[25] , \nbus_14523[24] 
		, \nbus_14523[23] , \nbus_14523[22] , \nbus_14523[21] , \nbus_14523[20] 
		, \nbus_14523[19] , \nbus_14523[18] , \nbus_14523[17] , \nbus_14523[16] 
		, \nbus_14523[15] , \nbus_14523[14] , \nbus_14523[13] , \nbus_14523[12] 
		, \nbus_14523[11] , \nbus_14523[10] , \nbus_14523[9] , \nbus_14523[8] 
		, \nbus_14523[7] , \nbus_14523[6] , \nbus_14523[5] , \nbus_14523[4] 
		, \nbus_14523[3] , \nbus_14523[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_56001, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, n_56172, ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({n_57042, n_57020, n_57078, n_57064}), .O0(opc_10));
	AWDP_INC_232 i_2388(.O0({n_5096, n_5094, n_5092, n_5090, n_5088, n_5086,
		 n_5084, n_5082, n_5080, n_5078, n_5076, n_5074, n_5072, n_5070,
		 n_5068, n_5066, n_5064, n_5062, n_5060, n_5058, n_5056, n_5054,
		 n_5052, n_5050, n_5048, n_5046, n_5044, n_5042, n_5040, n_5038,
		 n_5036, n_5034, n_5032, n_5030, n_5028, n_5026, n_5024, n_5022,
		 n_5020, n_5018, n_5016, n_5014, n_5012, n_5010, n_5008, n_5006,
		 n_5004, n_5002, n_5000, n_4998, n_4996, n_4994, n_4992, n_4990,
		 n_4988, n_4986, n_4984, n_4982, n_4980, n_4978, n_4976, n_4974,
		 n_4972, n_4970}), .tsc(tsc));
	AWDP_SUB_81 i_2342(.O0(regs_4_2), .regs_4(regs_4), .calc_sz({calc_sz[2],
		 n_58101, calc_sz[0]}));
	AWDP_ADD_114 i_2341(.O0({n_7380, n_7379, n_7378, n_7377, n_7376, n_7375,
		 n_7374, n_7373, n_7372, n_7371, n_7370, n_7369, n_7368, n_7367,
		 n_7366, n_7365, n_7364, n_7363, n_7362, n_7361, n_7360, n_7359,
		 n_7358, n_7357, n_7356, n_7355, n_7354, n_7353, n_7352, n_7351,
		 n_7350, n_7349}), .regs_4(regs_4), .calc_sz({calc_sz[2], n_58101
		, calc_sz[0]}));
	AWDP_ADD_67 i_2338(.O0({n_6411, n_6409, n_6407, n_6405, n_6403, n_6401, n_6399
		, n_6397, n_6395, n_6393, n_6391, n_6389, n_6387, n_6385, n_6383
		, n_6381, n_6379, n_6377, n_6375, n_6373, n_6371, n_6369, n_6367
		, n_6365, n_6363, n_6361, n_6359, n_6357, n_6355, n_6353, n_6351
		, n_6349}), .regs_7(regs_7), .opd({opd[31], opd[30], opd[29], opd
		[28], opd[27], opd[26], opd[25], opd[24], opd[23], opd[22], opd[
		21], opd[20], opd[19], opd[18], opd[17], opd[16], opd[15], opd[
		14], opd[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7],
		 opd[6], opd[5], n_59214, n_59222, n_59258, n_59240, n_59186})
		);
	AWDP_SUB_197 i_2337(.O0({n_6412, n_6410, n_6408, n_6406, n_6404, n_6402,
		 n_6400, n_6398, n_6396, n_6394, n_6392, n_6390, n_6388, n_6386,
		 n_6384, n_6382, n_6380, n_6378, n_6376, n_6374, n_6372, n_6370,
		 n_6368, n_6366, n_6364, n_6362, n_6360, n_6358, n_6356, n_6354,
		 n_6352, n_6350}), .regs_7(regs_7), .opd({opd[31], opd[30], opd[
		29], opd[28], opd[27], opd[26], opd[25], opd[24], opd[23], opd[
		22], opd[21], opd[20], opd[19], opd[18], opd[17], opd[16], opd[
		15], opd[14], opd[13], opd[12], opd[11], opd[10], opd[9], opd[8]
		, opd[7], opd[6], opd[5], n_59214, n_59222, n_59258, n_59240, n_59186
		}));
	shiftbox shiftbox(.shiftop({\opcode[3] , \opcode[2] , \opcode[1] , \opcode[0] 
		}), .calc_sz({calc_sz[3], calc_sz[2], n_58101, calc_sz[0]}), .ci
		(\eflags[0] ), .co(nCF_shiftbox), .co4(nCF_shift4box), .opa({opa
		[31], opa[30], opa[29], opa[28], opa[27], opa[26], opa[25], opa[
		24], opa[23], opa[22], opa[21], opa[20], opa[19], opa[18], opa[
		17], opa[16], n_60102, opa[14], opa[13], opa[12], opa[11], opa[
		10], opa[9], opa[8], n_60091, n_60082, opa[5], opa[4], opa[3], opa
		[2], opa[1], opa[0]}), .opb(opb), .resa(resa_shiftbox), .resb(resb_shiftbox
		), .resa4(resa_shift4box), .resb4(resb_shift4box));
	AWMUX_16_1 i_2321(.I0(\eflags[11] ), .I2(\eflags[0] ), .I4(\eflags[6] ),
		 .I6(\cond[6] ), .I8(\eflags[7] ), .I10(\eflags[2] ), .I12(\cond[12] 
		), .I14(\cond[14] ), .S({n_62892, n_62776, n_62864, n_62868}), .O0
		(cond_1));
	AWDP_ADD_5 i_2319(.add_len_pc32(add_len_pc32), .regs_14(regs_14), .lenpc
		(lenpc));
	AWDP_ADD_179 i_2318(.add_len_pc16({n_5175, n_5174, n_5173, n_5172, n_5171
		, n_5170, n_5169, n_5168, n_5167, n_5166, n_5165, n_5164, n_5163
		, n_5162, n_5161, n_5160}), .regs_14({regs_14[15], regs_14[14], regs_14
		[13], regs_14[12], regs_14[11], regs_14[10], regs_14[9], regs_14
		[8], regs_14[7], regs_14[6], regs_14[5], regs_14[4], regs_14[3],
		 regs_14[2], regs_14[1], regs_14[0]}), .lenpc({lenpc[15], lenpc[
		14], lenpc[13], lenpc[12], lenpc[11], lenpc[10], lenpc[9], lenpc
		[8], lenpc[7], lenpc[6], lenpc[5], lenpc[4], lenpc[3], lenpc[2],
		 lenpc[1], lenpc[0]}));
	AWDP_ADD_44 i_2313(.O0({n_11434, n_11433, n_11432, n_11431, n_11430, n_11429
		, n_11428, n_11427, n_11426, n_11425, n_11424, n_11423, n_11422,
		 n_11421, n_11420, n_11419, n_11418, n_11417, n_11416, n_11415, n_11414
		, n_11413, n_11412, n_11411, n_11410, n_11409, n_11408, n_11407,
		 n_11406, n_11405, n_11404, n_11403}), .I0({\nbus_11317[31] , \nbus_11317[30] 
		, \nbus_11317[29] , \nbus_11317[28] , n_328384274, \nbus_11317[26] 
		, \nbus_11317[25] , \nbus_11317[24] , \nbus_11317[23] , n_327984270
		, \nbus_11317[21] , \nbus_11317[20] , \nbus_11317[19] , \nbus_11317[18] 
		, \nbus_11317[17] , \nbus_11317[16] , n_327884269, n_327784268, n_327684267
		, n_327584266, n_327484265, \nbus_11317[10] , n_327384264, n_327284263
		, n_327184262, n_327084261, \nbus_11317[5] , n_346373943, n_328963506
		, \nbus_11317[2] , n_349680997, n_349580996}), .add_len_pc(add_len_pc
		));
	AWDP_EQ_111 i_2289(.O0({n_5179}), .mul64({mul64[63], mul64[62], mul64[61
		], mul64[60], mul64[59], mul64[58], mul64[57], mul64[56], mul64[
		55], mul64[54], mul64[53], mul64[52], mul64[51], mul64[50], mul64
		[49], mul64[48], mul64[47], mul64[46], mul64[45], mul64[44], mul64
		[43], mul64[42], mul64[41], mul64[40], mul64[39], mul64[38], mul64
		[37], mul64[36], mul64[35], mul64[34], mul64[33], mul64[32], mul64
		[31], mul64[30], mul64[29], mul64[28], mul64[27], mul64[26], mul64
		[25], mul64[24], mul64[23], mul64[22], mul64[21], mul64[20], mul64
		[19], mul64[18], mul64[17], mul64[16], mul64[15], mul64[14], mul64
		[13], mul64[12], mul64[11], mul64[10], mul64[9], mul64[8]}));
	AWDP_EQ_128 i_2288(.O0({n_5180}), .mul64({mul64[63], mul64[62], mul64[61
		], mul64[60], mul64[59], mul64[58], mul64[57], mul64[56], mul64[
		55], mul64[54], mul64[53], mul64[52], mul64[51], mul64[50], mul64
		[49], mul64[48], mul64[47], mul64[46], mul64[45], mul64[44], mul64
		[43], mul64[42], mul64[41], mul64[40], mul64[39], mul64[38], mul64
		[37], mul64[36], mul64[35], mul64[34], mul64[33], mul64[32], mul64
		[31], mul64[30], mul64[29], mul64[28], mul64[27], mul64[26], mul64
		[25], mul64[24], mul64[23], mul64[22], mul64[21], mul64[20], mul64
		[19], mul64[18], mul64[17], mul64[16]}));
	AWDP_EQ_231 i_2285(.O0({n_5183}), .mul64({mul64[63], mul64[62], mul64[61
		], mul64[60], mul64[59], mul64[58], mul64[57], mul64[56], mul64[
		55], mul64[54], mul64[53], mul64[52], mul64[51], mul64[50], mul64
		[49], mul64[48], mul64[47], mul64[46], mul64[45], mul64[44], mul64
		[43], mul64[42], mul64[41], mul64[40], mul64[39], mul64[38], mul64
		[37], mul64[36], mul64[35], mul64[34], mul64[33], mul64[32], mul64
		[31], mul64[30], mul64[29], mul64[28], mul64[27], mul64[26], mul64
		[25], mul64[24], mul64[23], mul64[22], mul64[21], mul64[20], mul64
		[19], mul64[18], mul64[17], mul64[16], mul64[15], mul64[14], mul64
		[13], mul64[12], mul64[11], mul64[10], mul64[9], mul64[8]}));
	AWDP_EQ_124 i_2283(.O0({n_5185}), .mul64({mul64[63], mul64[62], mul64[61
		], mul64[60], mul64[59], mul64[58], mul64[57], mul64[56], mul64[
		55], mul64[54], mul64[53], mul64[52], mul64[51], mul64[50], mul64
		[49], mul64[48], mul64[47], mul64[46], mul64[45], mul64[44], mul64
		[43], mul64[42], mul64[41], mul64[40], mul64[39], mul64[38], mul64
		[37], mul64[36], mul64[35], mul64[34], mul64[33], mul64[32], mul64
		[31], mul64[30], mul64[29], mul64[28], mul64[27], mul64[26], mul64
		[25], mul64[24], mul64[23], mul64[22], mul64[21], mul64[20], mul64
		[19], mul64[18], mul64[17], mul64[16]}));
	AWDP_EQ_222 i_2281(.O0({n_5187}), .mul64({mul64[63], mul64[62], mul64[61
		], mul64[60], mul64[59], mul64[58], mul64[57], mul64[56], mul64[
		55], mul64[54], mul64[53], mul64[52], mul64[51], mul64[50], mul64
		[49], mul64[48], mul64[47], mul64[46], mul64[45], mul64[44], mul64
		[43], mul64[42], mul64[41], mul64[40], mul64[39], mul64[38], mul64
		[37], mul64[36], mul64[35], mul64[34], mul64[33], mul64[32]}));
	AWDP_ADD_168 i_2275(.O0(nbus_157), .opa({opa[31], opa[30], opa[29], opa[
		28], opa[27], opa[26], opa[25], opa[24], opa[23], opa[22], opa[
		21], opa[20], opa[19], opa[18], opa[17], opa[16], n_60102, opa[
		14], opa[13], opa[12], opa[11], opa[10], opa[9], opa[8], n_60091
		, n_60082, opa[5], opa[4], opa[3], opa[2], opa[1], n_60072}), .opd
		({opd[31], opd[30], opd[29], opd[28], opd[27], opd[26], opd[25],
		 opd[24], opd[23], opd[22], opd[21], opd[20], opd[19], opd[18], opd
		[17], opd[16], opd[15], opd[14], opd[13], opd[12], opd[11], opd[
		10], opd[9], opd[8], opd[7], opd[6], opd[5], n_59214, n_59222, n_59258
		, n_59240, n_59186}));
	AWDP_ADD_21 i_2273(.O0(nbus_158), .opa({n_60102, opa[14], opa[13], opa[
		12], opa[11], opa[10], opa[9], opa[8], n_60091, n_60082, opa[5],
		 opa[4], opa[3], opa[2], opa[1], n_60072}), .opd({opd[15], opd[
		14], opd[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7],
		 opd[6], opd[5], opd[4], opd[3], opd[2], opd[1], opd[0]}));
	AWDP_ADD_121 i_2272(.O0(nbus_159), .opa({n_60091, n_60082, opa[5], opa[4
		], opa[3], opa[2], opa[1], n_60072}), .opd({opd[7], opd[6], opd[
		5], opd[4], opd[3], opd[2], opd[1], opd[0]}));
	AWDP_ADD_0 i_2271(.O0(nbus_160), .opb(opb), .I0({UNCONNECTED_000, 
		UNCONNECTED_001, UNCONNECTED_002, UNCONNECTED_003, 
		UNCONNECTED_004, UNCONNECTED_005, UNCONNECTED_006, 
		UNCONNECTED_007, UNCONNECTED_008, UNCONNECTED_009, 
		UNCONNECTED_010, UNCONNECTED_011, UNCONNECTED_012, n_57361, 
		UNCONNECTED_013, UNCONNECTED_014, UNCONNECTED_015, 
		UNCONNECTED_016, UNCONNECTED_017, UNCONNECTED_018, 
		UNCONNECTED_019, UNCONNECTED_020, UNCONNECTED_021, 
		UNCONNECTED_022, UNCONNECTED_023, UNCONNECTED_024, 
		UNCONNECTED_025, UNCONNECTED_026, UNCONNECTED_027, 
		UNCONNECTED_028, instrc[105], instrc[104]}));
	AWDP_ADD_109 i_2270(.O0(nbus_161), .opb({opb[15], opb[14], opb[13], opb[
		12], opb[11], opb[10], opb[9], opb[8], opb[7], opb[6], opb[5], opb
		[4], opb[3], opb[2], opb[1], opb[0]}), .I0({n_57361, 
		UNCONNECTED_029, UNCONNECTED_030, UNCONNECTED_031, 
		UNCONNECTED_032, UNCONNECTED_033, UNCONNECTED_034, 
		UNCONNECTED_035, UNCONNECTED_036, UNCONNECTED_037, 
		UNCONNECTED_038, UNCONNECTED_039, UNCONNECTED_040, 
		UNCONNECTED_041, instrc[105], instrc[104]}));
	AWDP_ADD_116 i_2269(.O0(nbus_162), .opa({opa[31], opa[30], opa[29], opa[
		28], opa[27], opa[26], opa[25], opa[24], opa[23], opa[22], opa[
		21], opa[20], opa[19], opa[18], opa[17], opa[16], n_60102, opa[
		14], opa[13], opa[12], opa[11], opa[10], opa[9], opa[8], n_60091
		, n_60082, opa[5], opa[4], opa[3], opa[2], opa[1], n_60072}), .I0
		({UNCONNECTED_042, UNCONNECTED_043, UNCONNECTED_044, 
		UNCONNECTED_045, UNCONNECTED_046, UNCONNECTED_047, 
		UNCONNECTED_048, UNCONNECTED_049, UNCONNECTED_050, 
		UNCONNECTED_051, UNCONNECTED_052, UNCONNECTED_053, n_57363, 
		UNCONNECTED_054, UNCONNECTED_055, UNCONNECTED_056, 
		UNCONNECTED_057, UNCONNECTED_058, UNCONNECTED_059, 
		UNCONNECTED_060, UNCONNECTED_061, UNCONNECTED_062, 
		UNCONNECTED_063, UNCONNECTED_064, UNCONNECTED_065, 
		UNCONNECTED_066, UNCONNECTED_067, UNCONNECTED_068, 
		UNCONNECTED_069, UNCONNECTED_070, instrc[105], instrc[104]}));
	AWDP_ADD_234 i_2268(.O0(nbus_163), .opa({n_60102, opa[14], opa[13], opa[
		12], opa[11], opa[10], opa[9], opa[8], n_60091, n_60082, opa[5],
		 opa[4], opa[3], opa[2], opa[1], n_60072}), .I0({UNCONNECTED_071
		, UNCONNECTED_072, n_57368, UNCONNECTED_073, UNCONNECTED_074, 
		UNCONNECTED_075, UNCONNECTED_076, UNCONNECTED_077, 
		UNCONNECTED_078, UNCONNECTED_079, UNCONNECTED_080, 
		UNCONNECTED_081, UNCONNECTED_082, UNCONNECTED_083, instrc[105], instrc
		[104]}));
	AWDP_SUB_206 i_2267(.O0(nbus_164), .opa({opa[31], opa[30], opa[29], opa[
		28], opa[27], opa[26], opa[25], opa[24], opa[23], opa[22], opa[
		21], opa[20], opa[19], opa[18], opa[17], opa[16], n_60102, opa[
		14], opa[13], opa[12], opa[11], opa[10], opa[9], opa[8], n_60091
		, n_60082, opa[5], opa[4], opa[3], opa[2], opa[1], n_60072}), .I0
		({UNCONNECTED_084, UNCONNECTED_085, UNCONNECTED_086, 
		UNCONNECTED_087, UNCONNECTED_088, UNCONNECTED_089, 
		UNCONNECTED_090, UNCONNECTED_091, UNCONNECTED_092, 
		UNCONNECTED_093, UNCONNECTED_094, UNCONNECTED_095, n_57361, 
		UNCONNECTED_096, UNCONNECTED_097, UNCONNECTED_098, 
		UNCONNECTED_099, UNCONNECTED_100, UNCONNECTED_101, 
		UNCONNECTED_102, UNCONNECTED_103, UNCONNECTED_104, 
		UNCONNECTED_105, UNCONNECTED_106, UNCONNECTED_107, 
		UNCONNECTED_108, UNCONNECTED_109, UNCONNECTED_110, 
		UNCONNECTED_111, UNCONNECTED_112, instrc[105], instrc[104]}));
	AWDP_SUB_129 i_2266(.O0(nbus_165), .opa({n_60102, opa[14], opa[13], opa[
		12], opa[11], opa[10], opa[9], opa[8], n_60091, n_60082, opa[5],
		 opa[4], opa[3], opa[2], opa[1], n_60072}), .I0({UNCONNECTED_113
		, UNCONNECTED_114, n_57363, UNCONNECTED_115, UNCONNECTED_116, 
		UNCONNECTED_117, UNCONNECTED_118, UNCONNECTED_119, 
		UNCONNECTED_120, UNCONNECTED_121, UNCONNECTED_122, 
		UNCONNECTED_123, UNCONNECTED_124, UNCONNECTED_125, instrc[105], instrc
		[104]}));
	AWDP_ADD_100 i_2265(.O0(nbus_166), .opd({opd[31], opd[30], opd[29], opd[
		28], opd[27], opd[26], opd[25], opd[24], opd[23], opd[22], opd[
		21], opd[20], opd[19], opd[18], opd[17], opd[16], opd[15], opd[
		14], opd[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7],
		 opd[6], opd[5], n_59214, n_59222, n_59258, n_59240, opd[0]}), .I0
		({UNCONNECTED_126, UNCONNECTED_127, UNCONNECTED_128, 
		UNCONNECTED_129, UNCONNECTED_130, UNCONNECTED_131, 
		UNCONNECTED_132, UNCONNECTED_133, UNCONNECTED_134, 
		UNCONNECTED_135, UNCONNECTED_136, UNCONNECTED_137, 
		UNCONNECTED_138, UNCONNECTED_139, UNCONNECTED_140, 
		UNCONNECTED_141, UNCONNECTED_142, UNCONNECTED_143, 
		UNCONNECTED_144, UNCONNECTED_145, UNCONNECTED_146, 
		UNCONNECTED_147, UNCONNECTED_148, UNCONNECTED_149, 
		UNCONNECTED_150, UNCONNECTED_151, UNCONNECTED_152, n_57363, 
		UNCONNECTED_153, UNCONNECTED_154, instrc[105], instrc[104]}));
	AWDP_ADD_149 i_2264(.O0(nbus_167), .opd({opd[15], opd[14], opd[13], opd[
		12], opd[11], opd[10], opd[9], opd[8], opd[7], opd[6], opd[5], n_59214
		, opd[3], opd[2], opd[1], n_59186}), .I0({UNCONNECTED_155, 
		UNCONNECTED_156, UNCONNECTED_157, UNCONNECTED_158, 
		UNCONNECTED_159, UNCONNECTED_160, UNCONNECTED_161, 
		UNCONNECTED_162, UNCONNECTED_163, UNCONNECTED_164, 
		UNCONNECTED_165, n_57362, UNCONNECTED_166, UNCONNECTED_167, instrc
		[105], instrc[104]}));
	AWDP_LSH_38 i_2263(.O0(nbus_11310), .opb({opb[4], opb[3], opb[2], opb[1]
		, opb[0]}));
	AWDP_ADD_69 i_2148(.O0({n_7343, n_7341, n_7339, n_7337, n_7335, n_7333, n_7331
		, n_7329, n_7327, n_7325, n_7323, n_7321, n_7319, n_7317, n_7315
		, n_7313, n_7311, n_7309, n_7307, n_7305, n_7303, n_7301, n_7299
		, n_7297, n_7295, n_7293, n_7291, n_7289, n_7287, n_7285, n_7283
		, n_7281}), .regs_6(regs_6), .opd({opd[31], opd[30], opd[29], opd
		[28], opd[27], opd[26], opd[25], opd[24], opd[23], opd[22], opd[
		21], opd[20], opd[19], opd[18], opd[17], opd[16], opd[15], opd[
		14], opd[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7],
		 opd[6], opd[5], n_59214, n_59222, n_59258, n_59240, n_59186})
		);
	AWDP_SUB_200 i_2147(.O0({n_7344, n_7342, n_7340, n_7338, n_7336, n_7334,
		 n_7332, n_7330, n_7328, n_7326, n_7324, n_7322, n_7320, n_7318,
		 n_7316, n_7314, n_7312, n_7310, n_7308, n_7306, n_7304, n_7302,
		 n_7300, n_7298, n_7296, n_7294, n_7292, n_7290, n_7288, n_7286,
		 n_7284, n_7282}), .regs_6(regs_6), .opd({opd[31], opd[30], opd[
		29], opd[28], opd[27], opd[26], opd[25], opd[24], opd[23], opd[
		22], opd[21], opd[20], opd[19], opd[18], opd[17], opd[16], opd[
		15], opd[14], opd[13], opd[12], opd[11], opd[10], opd[9], opd[8]
		, opd[7], opd[6], opd[5], n_59214, n_59222, n_59258, n_59240, n_59186
		}));
	AWDP_DEC_7 i_2117(.O0({\regs_1_0[31] , \regs_1_0[30] , \regs_1_0[29] , \regs_1_0[28] 
		, \regs_1_0[27] , \regs_1_0[26] , \regs_1_0[25] , \regs_1_0[24] 
		, \regs_1_0[23] , \regs_1_0[22] , \regs_1_0[21] , \regs_1_0[20] 
		, \regs_1_0[19] , \regs_1_0[18] , \regs_1_0[17] , \regs_1_0[16] 
		, n_8129, n_8128, n_8127, n_8126, n_8125, n_8124, n_8123, n_8122
		, n_8121, n_8120, n_8119, n_8118, n_8117, n_8116, n_8115, n_8114
		}), .ecx(ecx));
	AWDP_DEC_2 i_2116(.O0({\regs_1[15] , \regs_1[14] , \regs_1[13] , \regs_1[12] 
		, \regs_1[11] , \regs_1[10] , \regs_1[9] , \regs_1[8] , \regs_1[7] 
		, \regs_1[6] , \regs_1[5] , \regs_1[4] , \regs_1[3] , \regs_1[2] 
		, \regs_1[1] , \regs_1[0] }), .cx({ecx[15], ecx[14], ecx[13], ecx
		[12], ecx[11], ecx[10], ecx[9], ecx[8], ecx[7], ecx[6], ecx[5], ecx
		[4], ecx[3], ecx[2], ecx[1], ecx[0]}));
	AWDP_INC_212 i_2112(.O0({n_8193, n_8192, n_8191, n_8190, n_8189, n_8188,
		 n_8187, n_8186, n_8185, n_8184, n_8183, n_8182, n_8181, n_8180,
		 n_8179, n_8178, n_8177, n_8176, n_8175, n_8174, n_8173, n_8172,
		 n_8171, n_8170, n_8169, n_8168, n_8167, n_8166, n_8165, n_8164,
		 n_8163, n_8162, n_8161, n_8160, n_8159, n_8158, n_8157, n_8156,
		 n_8155, n_8154, n_8153, n_8152, n_8151, n_8150, n_8149, n_8148,
		 n_8147, n_8146, n_8145, n_8144, n_8143, n_8142, n_8141, n_8140,
		 n_8139, n_8138, n_8137, n_8136, n_8135, n_8134, n_8133, n_8132,
		 n_8131, n_8130}), .I0({nbus_11295[31], nbus_11295[30], nbus_11295
		[29], nbus_11295[28], n_57881, nbus_11295[26], nbus_11295[25], nbus_11295
		[24], nbus_11295[23], nbus_11295[22], nbus_11295[21], nbus_11295
		[20], nbus_11295[19], nbus_11295[18], nbus_11295[17], nbus_11295
		[16], nbus_11295[15], nbus_11295[14], nbus_11295[13], nbus_11295
		[12], nbus_11295[11], nbus_11295[10], nbus_11295[9], nbus_11295[
		8], nbus_11295[7], nbus_11295[6], nbus_11295[5], nbus_11295[4], n_57909
		, nbus_11295[2], nbus_11295[1], n_59717, n_59726, n_57828, n_57815
		, n_57802, n_57792, n_57783, n_57771, n_57761, n_57751, n_57742,
		 n_57733, n_57720, n_57707, n_57698, n_57689, n_57680, n_57671, n_57662
		, n_57653, n_57644, n_57635, n_57625, n_57613, n_57604, n_57957,
		 n_57592, n_57583, n_57574, n_57563, n_57552, n_57542, n_59742})
		);
	AWDP_INC_11111286 i_2109(.O0({UNCONNECTED_168, UNCONNECTED_169, 
		UNCONNECTED_170, UNCONNECTED_171, UNCONNECTED_172, 
		UNCONNECTED_173, UNCONNECTED_174, UNCONNECTED_175, 
		UNCONNECTED_176, UNCONNECTED_177, UNCONNECTED_178, 
		UNCONNECTED_179, UNCONNECTED_180, UNCONNECTED_181, 
		UNCONNECTED_182, UNCONNECTED_183, UNCONNECTED_184, 
		UNCONNECTED_185, UNCONNECTED_186, UNCONNECTED_187, 
		UNCONNECTED_188, UNCONNECTED_189, UNCONNECTED_190, 
		UNCONNECTED_191, UNCONNECTED_192, UNCONNECTED_193, 
		UNCONNECTED_194, UNCONNECTED_195, UNCONNECTED_196, 
		UNCONNECTED_197, UNCONNECTED_198, n_8226, n_8225, n_8224, n_8223
		, n_8222, n_8221, n_8220, n_8219, n_8218, n_8217, n_8216, n_8215
		, n_8214, n_8213, n_8212, n_8211, n_8210, n_8209, n_8208, n_8207
		, n_8206, n_8205, n_8204, n_8203, n_8202, n_8201, n_8200, n_8199
		, n_8198, n_8197, n_8196, n_8195, n_8194}), .I0({UNCONNECTED_199
		, UNCONNECTED_200, UNCONNECTED_201, UNCONNECTED_202, 
		UNCONNECTED_203, UNCONNECTED_204, UNCONNECTED_205, 
		UNCONNECTED_206, UNCONNECTED_207, UNCONNECTED_208, 
		UNCONNECTED_209, UNCONNECTED_210, UNCONNECTED_211, 
		UNCONNECTED_212, UNCONNECTED_213, UNCONNECTED_214, 
		UNCONNECTED_215, UNCONNECTED_216, UNCONNECTED_217, 
		UNCONNECTED_218, UNCONNECTED_219, UNCONNECTED_220, 
		UNCONNECTED_221, UNCONNECTED_222, UNCONNECTED_223, 
		UNCONNECTED_224, UNCONNECTED_225, UNCONNECTED_226, 
		UNCONNECTED_227, UNCONNECTED_228, UNCONNECTED_229, 
		UNCONNECTED_230, n_57837, n_55929, n_55956, n_55974, n_55938, n_55947
		, n_55965, n_56475, n_56347, n_56338, n_56329, n_56320, n_56311,
		 n_56302, n_56293, n_56284, n_56275, n_56248, n_56230, n_56221, n_56181
		, n_56154, n_56136, n_56118, n_56109, n_56082, n_56073, n_56064,
		 n_55983, n_55992, n_56010, n_56028}));
	AWDP_LE_215 i_2108(.O0({n_5219}), .divq(divq), .I0({UNCONNECTED_231, divr
		[63], divr[62], divr[61], divr[60], divr[59], divr[58], divr[57]
		, divr[56], divr[55], divr[54], divr[53], divr[52], divr[51], divr
		[50], divr[49], divr[48], divr[47], divr[46], divr[45], divr[44]
		, divr[43], divr[42], divr[41], divr[40], divr[39], divr[38], divr
		[37], divr[36], divr[35], divr[34], divr[33], divr[32], divr[31]
		, divr[30], divr[29], divr[28], divr[27], divr[26], divr[25], divr
		[24], divr[23], divr[22], divr[21], divr[20], divr[19], divr[18]
		, divr[17], divr[16], divr[15], divr[14], divr[13], divr[12], divr
		[11], divr[10], divr[9], divr[8], divr[7], divr[6], divr[5], divr
		[4], divr[3], divr[2], divr[1]}));
	AWDP_SUB_237 i_2105(.O0(divr_1), .divr(divr), .divq(divq));
	AWDP_GE_13 i_2103(.O0({n_5221}), .divr(divr), .divq(divq));
	AWDP_LSH_9 i_2102(.O0(nbus_11360), .opd({opd[5], n_59214, n_59222, n_59258
		, n_59240, n_59186}));
	AWDP_ADD_8 i_2101(.O0(opc_14), .opc({opc[31], opc[30], opc[29], opc[28],
		 opc[27], opc[26], opc[25], opc[24], opc[23], opc[22], opc[21], opc
		[20], opc[19], opc[18], opc[17], opc[16], opc[15], opc[14], opc[
		13], opc[12], opc[11], opc[10], opc[9], opc[8], opc[7], opc[6], opc
		[5], opc[4], opc[3], opc[2], opc[1], n_59735}), .I0(nbus_11360)
		);
	AWDP_INC_183 i_2095(.O0({n_8322, n_8321, n_8320, n_8319, n_8318, n_8317,
		 n_8316, n_8315, n_8314, n_8313, n_8312, n_8311, n_8310, n_8309,
		 n_8308, n_8307, n_8306, n_8305, n_8304, n_8303, n_8302, n_8301,
		 n_8300, n_8299, n_8298, n_8297, n_8296, n_8295, n_8294, n_8293,
		 n_8292, n_8291}), .I0(nbus_11328));
	AWDP_DEC_155 i_2092(.O0({\opc_1[7] , \opc_1[6] , \opc_1[5] , \opc_1[4] ,
		 \opc_1[3] , \opc_1[2] , \opc_1[1] , \opc_1[0] }), .opc({opc[7],
		 opc[6], opc[5], opc[4], opc[3], opc[2], opc[1], n_59735}));
	AWDP_DEC_83 i_2089(.O0({\opc_5[31] , \opc_5[30] , \opc_5[29] , \opc_5[28] 
		, \opc_5[27] , \opc_5[26] , \opc_5[25] , \opc_5[24] , \opc_5[23] 
		, \opc_5[22] , \opc_5[21] , \opc_5[20] , \opc_5[19] , \opc_5[18] 
		, \opc_5[17] , \opc_5[16] , \opc_5[15] , \opc_5[14] , \opc_5[13] 
		, \opc_5[12] , \opc_5[11] , \opc_5[10] , \opc_5[9] , \opc_5[8] ,
		 \opc_5[7] , \opc_5[6] , \opc_5[5] , n_8328, n_8327, n_8326, n_8325
		, n_8324}), .opc({opc[31], opc[30], opc[29], opc[28], opc[27], opc
		[26], opc[25], opc[24], opc[23], opc[22], opc[21], opc[20], opc[
		19], opc[18], opc[17], opc[16], opc[15], opc[14], opc[13], opc[
		12], opc[11], opc[10], opc[9], opc[8], opc[7], opc[6], opc[5], opc
		[4], opc[3], opc[2], opc[1], n_59735}));
	AWDP_EQ_158 i_2084(.O0({n_5227}), .I0({opb[31], opb[30], opb[29], opb[28
		], opb[27], opb[26], opb[25], opb[24], opb[23], opb[22], opb[21]
		, opb[20], opb[19], opb[18], opb[17], opb[16], opb[15], opb[14],
		 opb[13], opb[12], opb[11], opb[10], opb[9], opb[8], opb[7], opb
		[6], opb[5], opb[4], opb[3], opb[2], opb[1], opb[0], opc[31], opc
		[30], opc[29], opc[28], opc[27], opc[26], opc[25], opc[24], opc[
		23], opc[22], opc[21], opc[20], opc[19], opc[18], opc[17], opc[
		16], opc[15], opc[14], opc[13], opc[12], opc[11], opc[10], opc[9
		], opc[8], opc[7], opc[6], opc[5], opc[4], opc[3], opc[2], opc[1
		], n_59735}), .I1({regs_2[31], regs_2[30], regs_2[29], regs_2[28
		], regs_2[27], regs_2[26], regs_2[25], regs_2[24], regs_2[23], regs_2
		[22], regs_2[21], regs_2[20], regs_2[19], regs_2[18], regs_2[17]
		, regs_2[16], regs_2[15], regs_2[14], regs_2[13], regs_2[12], regs_2
		[11], regs_2[10], regs_2[9], regs_2[8], regs_2[7], regs_2[6], regs_2
		[5], regs_2[4], regs_2[3], regs_2[2], regs_2[1], regs_2[0], regs_0
		[31], regs_0[30], regs_0[29], regs_0[28], regs_0[27], regs_0[26]
		, regs_0[25], regs_0[24], regs_0[23], regs_0[22], regs_0[21], regs_0
		[20], regs_0[19], regs_0[18], regs_0[17], regs_0[16], regs_0[15]
		, regs_0[14], regs_0[13], regs_0[12], regs_0[11], regs_0[10], regs_0
		[9], regs_0[8], regs_0[7], regs_0[6], regs_0[5], regs_0[4], regs_0
		[3], regs_0[2], regs_0[1], regs_0[0]}));
	AWDP_INC_28 i_2076(.O0(opa_0), .I0({n_59726, n_57828, n_57815, n_57802, n_57792
		, n_57783, n_57771, n_57761, n_57751, n_57742, n_57733, n_57720,
		 n_57707, n_57698, n_57689, n_57680, n_57671, n_57662, n_57653, n_57644
		, n_57635, n_57625, n_57613, n_57604, n_57957, n_57592, n_57583,
		 n_57574, n_57563, n_57552, n_57542, n_59742}));
	AWDP_INC_167 i_2074(.O0({\opa_1[15] , \opa_1[14] , \opa_1[13] , \opa_1[12] 
		, \opa_1[11] , \opa_1[10] , \opa_1[9] , \opa_1[8] , \opa_1[7] , \opa_1[6] 
		, \opa_1[5] , \opa_1[4] , \opa_1[3] , \opa_1[2] , \opa_1[1] , \opa_1[0] 
		}), .I0({n_57671, n_57662, n_57653, n_57644, n_57635, n_57625, n_57613
		, n_57604, n_57957, n_57592, n_57583, n_57574, n_57563, n_57552,
		 n_57542, n_59742}));
	AWDP_INC_91 i_2063(.O0({n_10932, n_10931, n_10930, n_10929, n_10928, n_10927
		, n_10926, n_10925, n_10924, n_10923, n_10922, n_10921, n_10920,
		 n_10919, n_10918, n_10917, n_10916, n_10915, n_10914, n_10913, n_10912
		, n_10911, n_10910, n_10909, n_10908, n_10907, n_10906, n_10905,
		 n_10904, n_10903, n_10902, n_10901}), .I0({nbus_11295[31], nbus_11295
		[30], nbus_11295[29], nbus_11295[28], n_57881, nbus_11295[26], nbus_11295
		[25], nbus_11295[24], nbus_11295[23], nbus_11295[22], nbus_11295
		[21], nbus_11295[20], nbus_11295[19], nbus_11295[18], nbus_11295
		[17], nbus_11295[16], nbus_11295[15], nbus_11295[14], nbus_11295
		[13], nbus_11295[12], nbus_11295[11], nbus_11295[10], nbus_11295
		[9], nbus_11295[8], nbus_11295[7], nbus_11295[6], nbus_11295[5],
		 nbus_11295[4], n_57909, nbus_11295[2], nbus_11295[1], n_59717})
		);
	arithbox arithbox(.arithop({\opcode[3] , \opcode[2] , \opcode[1] , \opcode[0] 
		}), .calc_sz({calc_sz[3], calc_sz[2], n_58101, calc_sz[0]}), .ci
		(\eflags[0] ), .co(nCF_arithbox), .af(nAF_arithbox), .ai(\eflags[4] 
		), .sa(opas_arithbox), .sb(opbs_arithbox), .opa({opa[31], opa[30
		], opa[29], opa[28], opa[27], opa[26], opa[25], opa[24], opa[23]
		, opa[22], opa[21], opa[20], opa[19], opa[18], opa[17], opa[16],
		 n_60102, opa[14], opa[13], opa[12], opa[11], opa[10], opa[9], opa
		[8], n_60091, n_60082, opa[5], opa[4], opa[3], opa[2], opa[1], n_60072
		}), .opb(opb), .resa(resa_arithbox), .cmp(tcmp_arithbox));
	synthetic_op synthetic_op(.clk(clk), .sel({\opcode[2] , \opcode[1] , \opcode[0] 
		}), .opa32({opa[31], opa[30], opa[29], opa[28], opa[27], opa[26]
		, opa[25], opa[24], opa[23], opa[22], opa[21], opa[20], opa[19],
		 opa[18], opa[17], opa[16], n_60102, opa[14], opa[13], opa[12], opa
		[11], opa[10], opa[9], opa[8], n_60091, n_60082, opa[5], opa[4],
		 opa[3], opa[2], opa[1], n_60072}), .opb32(opb), .res64(mul64)
		);
	AWDP_ADD_40 i_2028(.O0({n_9369, n_9364, n_9359, n_9354, n_9349, n_9344, n_9339
		, n_9334, n_9329, n_9324, n_9319, n_9314, n_9309, n_9304, n_9299
		, n_9294, n_9289, n_9284, n_9279, n_9274, n_9269, n_9264, n_9259
		, n_9254, n_9249, n_9244, n_9239, n_9234, n_9229, n_9224, n_9219
		, n_9214}), .opb(opb), .I0({UNCONNECTED_232, UNCONNECTED_233, 
		UNCONNECTED_234, UNCONNECTED_235, UNCONNECTED_236, 
		UNCONNECTED_237, UNCONNECTED_238, UNCONNECTED_239, 
		UNCONNECTED_240, UNCONNECTED_241, UNCONNECTED_242, 
		UNCONNECTED_243, UNCONNECTED_244, UNCONNECTED_245, 
		UNCONNECTED_246, UNCONNECTED_247, UNCONNECTED_248, 
		UNCONNECTED_249, UNCONNECTED_250, UNCONNECTED_251, 
		UNCONNECTED_252, UNCONNECTED_253, UNCONNECTED_254, 
		UNCONNECTED_255, n_60091, n_60082, opa[5], opa[4], opa[3], opa[2
		], opa[1], n_60072}));
	AWDP_ADD_26 i_2026(.O0({n_9371, n_9365, n_9360, n_9355, n_9350, n_9345, n_9340
		, n_9335, n_9330, n_9325, n_9320, n_9315, n_9310, n_9305, n_9300
		, n_9295, n_9290, n_9285, n_9280, n_9275, n_9270, n_9265, n_9260
		, n_9255, n_9250, n_9245, n_9240, n_9235, n_9230, n_9225, n_9220
		, n_9215}), .opd(opd), .I0({UNCONNECTED_256, UNCONNECTED_257, 
		UNCONNECTED_258, opc[31], opc[30], opc[29], opc[28], opc[27], opc
		[26], opc[25], opc[24], opc[23], opc[22], opc[21], opc[20], opc[
		19], opc[18], opc[17], opc[16], opc[15], opc[14], opc[13], opc[
		12], opc[11], opc[10], opc[9], opc[8], opc[7], opc[6], opc[5], 
		UNCONNECTED_259, UNCONNECTED_260}));
	AWDP_ADD_123 i_2025(.O0({n_9372, n_9366, n_9361, n_9356, n_9351, n_9346,
		 n_9341, n_9336, n_9331, n_9326, n_9321, n_9316, n_9311, n_9306,
		 n_9301, n_9296, n_9291, n_9286, n_9281, n_9276, n_9271, n_9266,
		 n_9261, n_9256, n_9251, n_9246, n_9241, n_9236, n_9231, n_9226,
		 n_9221, n_9216}), .opd({opd[31], opd[30], opd[29], opd[28], opd
		[27], opd[26], opd[25], opd[24], opd[23], opd[22], opd[21], opd[
		20], opd[19], opd[18], opd[17], opd[16], opd[15], opd[14], opd[
		13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7], opd[6], opd
		[5], n_59214, n_59222, opd[2], n_59240, opd[0]}));
	AWDP_ADD_166 i_1992(.O0({n_5489, n_5487, n_5485, n_5483, n_5481, n_5479,
		 n_5477, n_5475, n_5473, n_5471, n_5469, n_5467, n_5465, n_5463,
		 n_5461, n_5459, n_5457, n_5455, n_5453, n_5451, n_5449, n_5447,
		 n_5445, n_5443, n_5441, n_5439, n_5437, n_5435, n_5433, n_5431,
		 n_5429, n_5427}), .ldtr(ldtr), .I0({gs[31], gs[30], gs[29], gs[
		28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs[
		20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs[
		12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], UNCONNECTED_261, UNCONNECTED_262, UNCONNECTED_263}));
	AWDP_ADD_169 i_1990(.O0({n_5490, n_5488, n_5486, n_5484, n_5482, n_5480,
		 n_5478, n_5476, n_5474, n_5472, n_5470, n_5468, n_5466, n_5464,
		 n_5462, n_5460, n_5458, n_5456, n_5454, n_5452, n_5450, n_5448,
		 n_5446, n_5444, n_5442, n_5440, n_5438, n_5436, n_5434, n_5432,
		 n_5430, n_5428}), .gdtr(gdtr), .I0({gs[31], gs[30], gs[29], gs[
		28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs[
		20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs[
		12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], UNCONNECTED_264, UNCONNECTED_265, UNCONNECTED_266}));
	AWDP_ADD_92 i_1987(.O0({n_11317, n_11315, n_11313, n_11311, n_11309, n_11307
		, n_11305, n_11303, n_11301, n_11299, n_11297, n_11295, n_11293,
		 n_11291, n_11289, n_11287, n_11285, n_11283, n_11281, n_11279, n_11277
		, n_11275, n_11273, n_11271, n_11269, n_11267, n_11265, n_11263,
		 n_11261, n_11259, n_11257, n_11255}), .idtr(idtr), .I0({instrc[
		95], instrc[94], instrc[93], instrc[92], instrc[91], instrc[90],
		 instrc[89], instrc[88], instrc[87], instrc[86], instrc[85], instrc
		[84], instrc[83], instrc[82], instrc[81], instrc[80], 
		UNCONNECTED_267, UNCONNECTED_268, UNCONNECTED_269}));
	AWDP_ADD_61 i_1985(.O0({n_11318, n_11316, n_11314, n_11312, n_11310, n_11308
		, n_11306, n_11304, n_11302, n_11300, n_11298, n_11296, n_11294,
		 n_11292, n_11290, n_11288, n_11286, n_11284, n_11282, n_11280, n_11278
		, n_11276, n_11274, n_11272, n_11270, n_11268, n_11266, n_11264,
		 n_11262, n_11260, n_11258, n_11256}), .gdtr(gdtr), .I0({\tr[15] 
		, \tr[14] , \tr[13] , \tr[12] , \tr[11] , \tr[10] , \tr[9] , \tr[8] 
		, \tr[7] , \tr[6] , \tr[5] , \tr[4] , \tr[3] , UNCONNECTED_270, 
		UNCONNECTED_271, UNCONNECTED_272}));
	AWDP_SUB_177 i_1984(.O0(Daddrs_8), .opd({opd[31], opd[30], opd[29], opd[
		28], opd[27], opd[26], opd[25], opd[24], opd[23], opd[22], opd[
		21], opd[20], opd[19], opd[18], opd[17], opd[16], opd[15], opd[
		14], opd[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7],
		 opd[6], opd[5], n_59214, n_59222, n_59258, n_59240, opd[0]}));
	AWDP_ADD_47 i_1983(.O0(Daddrs_1), .Daddrs(Daddr));
	AWDP_ADD_62 i_1982(.O0(Daddrs_3), .Daddrs(Daddr));
	AWDP_ADD_24 i_1980(.O0({n_9889, n_9888, n_9887, n_9886, n_9885, n_9884, n_9883
		, n_9882, n_9881, n_9880, n_9879, n_9878, n_9877, n_9876, n_9875
		, n_9874, n_9873, n_9872, n_9871, n_9870, n_9869, n_9868, n_9867
		, n_9866, n_9865, n_9864, n_9863, n_9862, n_9861, n_9860, n_9859
		, n_9858}), .opd(opd), .desc(desc));
	AWDP_ADD_102 i_1945(.O0({n_6084, n_6083, n_6082, n_6081, n_6080, n_6079,
		 n_6078, n_6077, n_6076, n_6075, n_6074, n_6073, n_6072, n_6071,
		 n_6070, n_6069, n_6068, n_6067, n_6066, n_6065, n_6064, n_6063,
		 n_6062, n_6061, n_6060, n_6059, n_6058, n_6057, n_6056, n_6055,
		 n_6054, n_6053}), .I0({UNCONNECTED_273, UNCONNECTED_274, 
		UNCONNECTED_275, UNCONNECTED_276, UNCONNECTED_277, 
		UNCONNECTED_278, UNCONNECTED_279, UNCONNECTED_280, 
		UNCONNECTED_281, UNCONNECTED_282, UNCONNECTED_283, 
		UNCONNECTED_284, UNCONNECTED_285, UNCONNECTED_286, 
		UNCONNECTED_287, UNCONNECTED_288, regs_14[15], regs_14[14], regs_14
		[13], regs_14[12], regs_14[11], regs_14[10], regs_14[9], regs_14
		[8], regs_14[7], regs_14[6], regs_14[5], regs_14[4], regs_14[3],
		 regs_14[2], regs_14[1], regs_14[0]}), .I1({\nbus_14523[27] , \nbus_14523[26] 
		, \nbus_14523[25] , \nbus_14523[24] , \nbus_14523[23] , \nbus_14523[22] 
		, \nbus_14523[21] , \nbus_14523[20] , \nbus_14523[19] , \nbus_14523[18] 
		, \nbus_14523[17] , \nbus_14523[16] , \nbus_14523[15] , \nbus_14523[14] 
		, \nbus_14523[13] , \nbus_14523[12] , \nbus_14523[11] , \nbus_14523[10] 
		, \nbus_14523[9] , \nbus_14523[8] , \nbus_14523[7] , \nbus_14523[6] 
		, \nbus_14523[5] , \nbus_14523[4] , \nbus_14523[3] , \nbus_14523[2] 
		, cs[1], cs[0], UNCONNECTED_289, UNCONNECTED_290, 
		UNCONNECTED_291, UNCONNECTED_292}));
endmodule
module cpu(clk, rstn, iack, int_cpu, ivect, cr0, cr2, icr2, cr3, cs, pg_fault, ipg_fault
		, useq_ptr, valid_len, queue, pg_en, pc_out, pc_req, read_req, write_req
		, read_ack, write_ack, flush_Itlb, flush_Dtlb, readio_req, writeio_req
		, readio_ack, writeio_ack, write_data, writeio_data, read_data, readio_data
		, write_sz, read_sz, io_add, Daddr, pt_fault, wr_fault);

	input clk;
	input rstn;
	output iack;
	input int_cpu;
	input [7:0] ivect;
	output [31:0] cr0;
	input [31:0] cr2;
	input [31:0] icr2;
	output [31:0] cr3;
	output [31:0] cs;
	input pg_fault;
	input ipg_fault;
	output [3:0] useq_ptr;
	input [5:0] valid_len;
	input [127:0] queue;
	output pg_en;
	output [31:0] pc_out;
	output pc_req;
	output read_req;
	output write_req;
	input read_ack;
	input write_ack;
	output flush_Itlb;
	output flush_Dtlb;
	output readio_req;
	output writeio_req;
	input readio_ack;
	input writeio_ack;
	output [31:0] write_data;
	output [31:0] writeio_data;
	input [31:0] read_data;
	input [31:0] readio_data;
	output [1:0] write_sz;
	output [1:0] read_sz;
	output [31:0] io_add;
	output [31:0] Daddr;
	input pt_fault;
	input wr_fault;

	wire [2:0] reps;
	wire [2:0] opz;
	wire [127:0] dec2vliw;
	wire [31:0] lenpc;
	wire [31:0] add_src;
	wire [7:0] from_acu;
	wire [63:0] to_acu;
	wire [210:0] deco2acu;



	vliw i_vliw(.clk(clk), .rstn(rstn), .instrc(dec2vliw), .ie(ie), .readio_data
		(readio_data), .io_add({UNCONNECTED_000, UNCONNECTED_001, 
		UNCONNECTED_002, UNCONNECTED_003, UNCONNECTED_004, 
		UNCONNECTED_005, UNCONNECTED_006, UNCONNECTED_007, 
		UNCONNECTED_008, UNCONNECTED_009, UNCONNECTED_010, 
		UNCONNECTED_011, UNCONNECTED_012, UNCONNECTED_013, 
		UNCONNECTED_014, UNCONNECTED_015, io_add[15], io_add[14], io_add
		[13], io_add[12], io_add[11], io_add[10], io_add[9], io_add[8], io_add
		[7], io_add[6], io_add[5], io_add[4], io_add[3], io_add[2], io_add
		[1], io_add[0]}), .writeio_data(writeio_data), .writeio_req(writeio_req
		), .readio_req(readio_req), .writeio_ack(writeio_ack), .readio_ack
		(readio_ack), .read_reqs(read_req), .read_ack(read_ack), .read_data
		(read_data), .over_seg({\over_seg[5] , UNCONNECTED_016, 
		UNCONNECTED_017, UNCONNECTED_018, UNCONNECTED_019, 
		UNCONNECTED_020}), .cr3({cr3[31], cr3[30], cr3[29], cr3[28], cr3
		[27], cr3[26], cr3[25], cr3[24], cr3[23], cr3[22], cr3[21], cr3[
		20], cr3[19], cr3[18], cr3[17], cr3[16], cr3[15], cr3[14], cr3[
		13], cr3[12], UNCONNECTED_021, UNCONNECTED_022, UNCONNECTED_023,
		 UNCONNECTED_024, UNCONNECTED_025, UNCONNECTED_026, 
		UNCONNECTED_027, UNCONNECTED_028, UNCONNECTED_029, 
		UNCONNECTED_030, UNCONNECTED_031, UNCONNECTED_032}), .cr2(cr2), 
		.icr2(icr2), .cr0({UNCONNECTED_033, UNCONNECTED_034, 
		UNCONNECTED_035, UNCONNECTED_036, UNCONNECTED_037, 
		UNCONNECTED_038, UNCONNECTED_039, UNCONNECTED_040, 
		UNCONNECTED_041, UNCONNECTED_042, UNCONNECTED_043, 
		UNCONNECTED_044, UNCONNECTED_045, UNCONNECTED_046, 
		UNCONNECTED_047, cr0[16], UNCONNECTED_048, UNCONNECTED_049, 
		UNCONNECTED_050, UNCONNECTED_051, UNCONNECTED_052, 
		UNCONNECTED_053, UNCONNECTED_054, UNCONNECTED_055, 
		UNCONNECTED_056, UNCONNECTED_057, UNCONNECTED_058, 
		UNCONNECTED_059, UNCONNECTED_060, \cr0[2] , UNCONNECTED_061, \cr0[0] 
		}), .write_reqs(write_req), .write_ack(write_ack), .write_data(write_data
		), .Daddr(Daddr), .write_sz(write_sz), .cs({UNCONNECTED_062, 
		UNCONNECTED_063, UNCONNECTED_064, UNCONNECTED_065, 
		UNCONNECTED_066, UNCONNECTED_067, UNCONNECTED_068, 
		UNCONNECTED_069, UNCONNECTED_070, UNCONNECTED_071, 
		UNCONNECTED_072, UNCONNECTED_073, UNCONNECTED_074, 
		UNCONNECTED_075, UNCONNECTED_076, UNCONNECTED_077, 
		UNCONNECTED_078, UNCONNECTED_079, UNCONNECTED_080, 
		UNCONNECTED_081, UNCONNECTED_082, UNCONNECTED_083, 
		UNCONNECTED_084, UNCONNECTED_085, UNCONNECTED_086, 
		UNCONNECTED_087, UNCONNECTED_088, UNCONNECTED_089, 
		UNCONNECTED_090, UNCONNECTED_091, cs[1], cs[0]}), .add_src(add_src
		), .from_acu(from_acu), .to_acu(to_acu), .pg_en(pg_en), .imm({
		UNCONNECTED_092, UNCONNECTED_093, UNCONNECTED_094, 
		UNCONNECTED_095, UNCONNECTED_096, UNCONNECTED_097, 
		UNCONNECTED_098, UNCONNECTED_099, UNCONNECTED_100, 
		UNCONNECTED_101, UNCONNECTED_102, UNCONNECTED_103, 
		UNCONNECTED_104, UNCONNECTED_105, UNCONNECTED_106, 
		UNCONNECTED_107, \imm[47] , \imm[46] , \imm[45] , \imm[44] , \imm[43] 
		, \imm[42] , \imm[41] , \imm[40] , \imm[39] , \imm[38] , \imm[37] 
		, \imm[36] , \imm[35] , \imm[34] , \imm[33] , \imm[32] , \imm[31] 
		, \imm[30] , \imm[29] , \imm[28] , \imm[27] , \imm[26] , \imm[25] 
		, \imm[24] , \imm[23] , \imm[22] , \imm[21] , \imm[20] , \imm[19] 
		, \imm[18] , \imm[17] , \imm[16] , \imm[15] , \imm[14] , \imm[13] 
		, \imm[12] , \imm[11] , \imm[10] , \imm[9] , \imm[8] , \imm[7] ,
		 \imm[6] , \imm[5] , \imm[4] , \imm[3] , \imm[2] , \imm[1] , \imm[0] 
		}), .lenpc(lenpc), .pc_out(pc_out), .pc_req(pc_req), .opz(opz), 
		.reps(reps), .flush_tlb(flush_Itlb), .flush_Dtlb(flush_Dtlb), .terminate
		(term), .start_up(st), .pg_fault(pg_fault), .ipg_fault(ipg_fault
		), .wr_fault(wr_fault), .pt_fault(pt_fault));
	acu i_acu(.clk(clk), .rstn(rstn), .from_regf(to_acu), .add_src(add_src),
		 .to_regf(from_acu), .from_dec(deco2acu), .db67(\cr0[0] ));
	deco i_deco(.clk(clk), .rstn(rstn), .useq_ptr(useq_ptr), .in128(queue), 
		.adz(\cr0[0] ), .pc_req(pc_req), .ivect(ivect), .int_main(int_cpu
		), .iack(iack), .ie(ie), .pg_fault(pg_fault), .ipg_fault(ipg_fault
		), .cpl({cs[1], cs[0]}), .cr0({UNCONNECTED_108, UNCONNECTED_109,
		 UNCONNECTED_110, UNCONNECTED_111, UNCONNECTED_112, 
		UNCONNECTED_113, UNCONNECTED_114, UNCONNECTED_115, 
		UNCONNECTED_116, UNCONNECTED_117, UNCONNECTED_118, 
		UNCONNECTED_119, UNCONNECTED_120, UNCONNECTED_121, 
		UNCONNECTED_122, UNCONNECTED_123, UNCONNECTED_124, 
		UNCONNECTED_125, UNCONNECTED_126, UNCONNECTED_127, 
		UNCONNECTED_128, UNCONNECTED_129, UNCONNECTED_130, 
		UNCONNECTED_131, UNCONNECTED_132, UNCONNECTED_133, 
		UNCONNECTED_134, UNCONNECTED_135, UNCONNECTED_136, \cr0[2] , 
		UNCONNECTED_137, UNCONNECTED_138}), .valid_len(valid_len), .to_vliw
		(dec2vliw), .lenpc_out(lenpc), .immediate({UNCONNECTED_139, 
		UNCONNECTED_140, UNCONNECTED_141, UNCONNECTED_142, 
		UNCONNECTED_143, UNCONNECTED_144, UNCONNECTED_145, 
		UNCONNECTED_146, UNCONNECTED_147, UNCONNECTED_148, 
		UNCONNECTED_149, UNCONNECTED_150, UNCONNECTED_151, 
		UNCONNECTED_152, UNCONNECTED_153, UNCONNECTED_154, \imm[47] , \imm[46] 
		, \imm[45] , \imm[44] , \imm[43] , \imm[42] , \imm[41] , \imm[40] 
		, \imm[39] , \imm[38] , \imm[37] , \imm[36] , \imm[35] , \imm[34] 
		, \imm[33] , \imm[32] , \imm[31] , \imm[30] , \imm[29] , \imm[28] 
		, \imm[27] , \imm[26] , \imm[25] , \imm[24] , \imm[23] , \imm[22] 
		, \imm[21] , \imm[20] , \imm[19] , \imm[18] , \imm[17] , \imm[16] 
		, \imm[15] , \imm[14] , \imm[13] , \imm[12] , \imm[11] , \imm[10] 
		, \imm[9] , \imm[8] , \imm[7] , \imm[6] , \imm[5] , \imm[4] , \imm[3] 
		, \imm[2] , \imm[1] , \imm[0] }), .to_acu(deco2acu), .operand_size
		(opz), .reps(reps), .over_seg({\over_seg[5] , UNCONNECTED_155, 
		UNCONNECTED_156, UNCONNECTED_157, UNCONNECTED_158, 
		UNCONNECTED_159}), .term(term), .start(st));
endmodule
module AWDP_ADD_10(O0, addr);

	output [31:0] O0;
	input [31:0] addr;

	wire \addr[4] ;
	wire \addr[5] ;
	wire \addr[6] ;
	wire \addr[7] ;
	wire \addr[8] ;
	wire \addr[9] ;
	wire \addr[10] ;
	wire \addr[11] ;
	wire \addr[12] ;
	wire \addr[13] ;
	wire \addr[14] ;
	wire \addr[15] ;
	wire \addr[16] ;
	wire \addr[17] ;
	wire \addr[18] ;
	wire \addr[19] ;
	wire \addr[20] ;
	wire \addr[21] ;
	wire \addr[22] ;
	wire \addr[23] ;
	wire \addr[24] ;
	wire \addr[25] ;
	wire \addr[26] ;
	wire \addr[27] ;
	wire \addr[28] ;
	wire \addr[29] ;
	wire \addr[30] ;
	wire \addr[31] ;


	assign O0[0] = addr[0];
	assign O0[1] = addr[1];
	assign O0[2] = addr[2];
	assign O0[3] = addr[3];
	assign \addr[4]  = addr[4];
	assign \addr[5]  = addr[5];
	assign \addr[6]  = addr[6];
	assign \addr[7]  = addr[7];
	assign \addr[8]  = addr[8];
	assign \addr[9]  = addr[9];
	assign \addr[10]  = addr[10];
	assign \addr[11]  = addr[11];
	assign \addr[12]  = addr[12];
	assign \addr[13]  = addr[13];
	assign \addr[14]  = addr[14];
	assign \addr[15]  = addr[15];
	assign \addr[16]  = addr[16];
	assign \addr[17]  = addr[17];
	assign \addr[18]  = addr[18];
	assign \addr[19]  = addr[19];
	assign \addr[20]  = addr[20];
	assign \addr[21]  = addr[21];
	assign \addr[22]  = addr[22];
	assign \addr[23]  = addr[23];
	assign \addr[24]  = addr[24];
	assign \addr[25]  = addr[25];
	assign \addr[26]  = addr[26];
	assign \addr[27]  = addr[27];
	assign \addr[28]  = addr[28];
	assign \addr[29]  = addr[29];
	assign \addr[30]  = addr[30];
	assign \addr[31]  = addr[31];

	notech_ha2 i_27(.A(\addr[31] ), .B(n_300), .Z(O0[31]));
	notech_ha2 i_26(.A(\addr[30] ), .B(n_298), .Z(O0[30]), .CO(n_300));
	notech_ha2 i_25(.A(\addr[29] ), .B(n_296), .Z(O0[29]), .CO(n_298));
	notech_ha2 i_24(.A(\addr[28] ), .B(n_294), .Z(O0[28]), .CO(n_296));
	notech_ha2 i_23(.A(\addr[27] ), .B(n_292), .Z(O0[27]), .CO(n_294));
	notech_ha2 i_22(.A(\addr[26] ), .B(n_290), .Z(O0[26]), .CO(n_292));
	notech_ha2 i_21(.A(\addr[25] ), .B(n_288), .Z(O0[25]), .CO(n_290));
	notech_ha2 i_20(.A(\addr[24] ), .B(n_286), .Z(O0[24]), .CO(n_288));
	notech_ha2 i_19(.A(\addr[23] ), .B(n_284), .Z(O0[23]), .CO(n_286));
	notech_ha2 i_18(.A(\addr[22] ), .B(n_282), .Z(O0[22]), .CO(n_284));
	notech_ha2 i_17(.A(\addr[21] ), .B(n_280), .Z(O0[21]), .CO(n_282));
	notech_ha2 i_16(.A(\addr[20] ), .B(n_278), .Z(O0[20]), .CO(n_280));
	notech_ha2 i_15(.A(\addr[19] ), .B(n_276), .Z(O0[19]), .CO(n_278));
	notech_ha2 i_14(.A(\addr[18] ), .B(n_274), .Z(O0[18]), .CO(n_276));
	notech_ha2 i_13(.A(\addr[17] ), .B(n_272), .Z(O0[17]), .CO(n_274));
	notech_ha2 i_12(.A(\addr[16] ), .B(n_270), .Z(O0[16]), .CO(n_272));
	notech_ha2 i_11(.A(\addr[15] ), .B(n_268), .Z(O0[15]), .CO(n_270));
	notech_ha2 i_10(.A(\addr[14] ), .B(n_266), .Z(O0[14]), .CO(n_268));
	notech_ha2 i_9(.A(\addr[13] ), .B(n_264), .Z(O0[13]), .CO(n_266));
	notech_ha2 i_8(.A(\addr[12] ), .B(n_262), .Z(O0[12]), .CO(n_264));
	notech_ha2 i_7(.A(\addr[11] ), .B(n_260), .Z(O0[11]), .CO(n_262));
	notech_ha2 i_6(.A(\addr[10] ), .B(n_258), .Z(O0[10]), .CO(n_260));
	notech_ha2 i_5(.A(\addr[9] ), .B(n_256), .Z(O0[9]), .CO(n_258));
	notech_ha2 i_4(.A(\addr[8] ), .B(n_254), .Z(O0[8]), .CO(n_256));
	notech_ha2 i_3(.A(\addr[7] ), .B(n_252), .Z(O0[7]), .CO(n_254));
	notech_ha2 i_2(.A(\addr[6] ), .B(n_250), .Z(O0[6]), .CO(n_252));
	notech_ha2 i_1(.A(\addr[5] ), .B(\addr[4] ), .Z(O0[5]), .CO(n_250));
	notech_inv i_0(.A(\addr[4] ), .Z(O0[4]));
endmodule
module AWDP_ADD_33(O0, addrshft, useq_ptr);
    output [6:0] O0;
    input [5:0] addrshft;
    input [3:0] useq_ptr;
    // Line 87
    wire [6:0] N875;
    // Line 58
    wire [6:0] O0;

    // Line 87
    assign N875 = useq_ptr + addrshft;
    // Line 58
    assign O0 = N875;
endmodule

module AWDP_EQ_2715865(O0, addr, addrf);
    output [0:0] O0;
    input [31:0] addr;
    input [31:0] addrf;
    // Line 58
    wire [0:0] O0;
    // Line 91
    wire [0:0] N881;

    // Line 58
    assign O0 = N881;
    // Line 91
    assign N881 = addr == addrf;
endmodule

module AWDP_EQ_3416052(O0, tagA, addr);
    output [0:0] O0;
    input [17:0] tagA;
    input [31:14] addr;
    // Line 134
    wire [0:0] N889;
    // Line 134
    wire [0:0] O0;

    // Line 134
    assign N889 = tagA == addr;
    // Line 134
    assign O0 = N889;
endmodule

module AWDP_INC_1315491(O0, purge_cnt);

	output [10:0] O0;
	input [10:0] purge_cnt;




	notech_ha2 i_10(.A(purge_cnt[10]), .B(n_106), .Z(O0[10]));
	notech_ha2 i_9(.A(purge_cnt[9]), .B(n_104), .Z(O0[9]), .CO(n_106));
	notech_ha2 i_8(.A(purge_cnt[8]), .B(n_102), .Z(O0[8]), .CO(n_104));
	notech_ha2 i_7(.A(purge_cnt[7]), .B(n_100), .Z(O0[7]), .CO(n_102));
	notech_ha2 i_6(.A(purge_cnt[6]), .B(n_98), .Z(O0[6]), .CO(n_100));
	notech_ha2 i_5(.A(purge_cnt[5]), .B(n_96), .Z(O0[5]), .CO(n_98));
	notech_ha2 i_4(.A(purge_cnt[4]), .B(n_94), .Z(O0[4]), .CO(n_96));
	notech_ha2 i_3(.A(purge_cnt[3]), .B(n_92), .Z(O0[3]), .CO(n_94));
	notech_ha2 i_2(.A(purge_cnt[2]), .B(n_90), .Z(O0[2]), .CO(n_92));
	notech_ha2 i_1(.A(purge_cnt[1]), .B(purge_cnt[0]), .Z(O0[1]), .CO(n_90)
		);
	notech_inv i_0(.A(purge_cnt[0]), .Z(O0[0]));
endmodule
module useq(iaddr, idata, code_req, code_ack, clk, rstn, useq_ptr, squeue, pc_in
		, pc_req, cs, pg_en, pg_fault, pc_pg_fault, valid_len, busy_ram
		);

	output [31:0] iaddr;
	input [127:0] idata;
	output code_req;
	input code_ack;
	input clk;
	input rstn;
	input [3:0] useq_ptr;
	output [127:0] squeue;
	input [31:0] pc_in;
	input pc_req;
	input [31:0] cs;
	input pg_en;
	input pg_fault;
	output pc_pg_fault;
	output [5:0] valid_len;
	input busy_ram;

	wire [1:0] wptr;
	wire [1:0] fault_wptr;
	wire [255:0] queue;
	wire [17:0] tagA;
	wire [3:0] tagV;
	wire [31:0] addr_0;
	wire [149:0] cacheD;
	wire [9:0] cacheA;
	wire [6:0] nbus_81;
	wire [10:0] purge_cnt;
	wire [5:0] addrshft;
	wire [31:0] addrf;

	supply0 AMBIT_GND;
	supply1 AMBIT_VDD;


	notech_inv i_16134(.A(n_62887), .Z(n_62888));
	notech_inv i_16133(.A(n_62882), .Z(n_62887));
	notech_inv i_16132(.A(n_62885), .Z(n_62886));
	notech_inv i_16131(.A(n_62878), .Z(n_62885));
	notech_inv i_16130(.A(n_62883), .Z(n_62884));
	notech_inv i_16129(.A(n_62876), .Z(n_62883));
	notech_inv i_16128(.A(n_62881), .Z(n_62882));
	notech_inv i_16127(.A(n_62884), .Z(n_62881));
	notech_inv i_16126(.A(n_62879), .Z(n_62880));
	notech_inv i_16125(.A(cacheD[148]), .Z(n_62879));
	notech_inv i_16124(.A(n_62877), .Z(n_62878));
	notech_inv i_16123(.A(n_62880), .Z(n_62877));
	notech_inv i_16122(.A(n_62875), .Z(n_62876));
	notech_inv i_16121(.A(n_62886), .Z(n_62875));
	notech_inv i_15992(.A(n_62745), .Z(n_62746));
	notech_inv i_15991(.A(n_62696), .Z(n_62745));
	notech_inv i_15950(.A(n_62703), .Z(n_62704));
	notech_inv i_15949(.A(n_62628), .Z(n_62703));
	notech_inv i_15948(.A(n_62701), .Z(n_62702));
	notech_inv i_15947(.A(n_62622), .Z(n_62701));
	notech_inv i_15946(.A(n_62699), .Z(n_62700));
	notech_inv i_15945(.A(n_62618), .Z(n_62699));
	notech_inv i_15944(.A(n_62697), .Z(n_62698));
	notech_inv i_15943(.A(n_62616), .Z(n_62697));
	notech_inv i_15942(.A(n_62695), .Z(n_62696));
	notech_inv i_15941(.A(n_62698), .Z(n_62695));
	notech_inv i_15878(.A(n_62631), .Z(n_62632));
	notech_inv i_15877(.A(n_62556), .Z(n_62631));
	notech_inv i_15876(.A(n_62629), .Z(n_62630));
	notech_inv i_15875(.A(n_62554), .Z(n_62629));
	notech_inv i_15874(.A(n_62627), .Z(n_62628));
	notech_inv i_15873(.A(n_62630), .Z(n_62627));
	notech_inv i_15872(.A(n_62625), .Z(n_62626));
	notech_inv i_15871(.A(n_62550), .Z(n_62625));
	notech_inv i_15870(.A(n_62623), .Z(n_62624));
	notech_inv i_15869(.A(n_62548), .Z(n_62623));
	notech_inv i_15868(.A(n_62621), .Z(n_62622));
	notech_inv i_15867(.A(n_62624), .Z(n_62621));
	notech_inv i_15866(.A(n_62619), .Z(n_62620));
	notech_inv i_15865(.A(n_62546), .Z(n_62619));
	notech_inv i_15864(.A(n_62617), .Z(n_62618));
	notech_inv i_15863(.A(n_62620), .Z(n_62617));
	notech_inv i_15862(.A(n_62615), .Z(n_62616));
	notech_inv i_15861(.A(n_62700), .Z(n_62615));
	notech_inv i_15804(.A(n_62557), .Z(n_62558));
	notech_inv i_15803(.A(clk), .Z(n_62557));
	notech_inv i_15802(.A(n_62555), .Z(n_62556));
	notech_inv i_15801(.A(n_62558), .Z(n_62555));
	notech_inv i_15800(.A(n_62553), .Z(n_62554));
	notech_inv i_15799(.A(n_62632), .Z(n_62553));
	notech_inv i_15798(.A(n_62551), .Z(n_62552));
	notech_inv i_15797(.A(n_62458), .Z(n_62551));
	notech_inv i_15796(.A(n_62549), .Z(n_62550));
	notech_inv i_15795(.A(n_62552), .Z(n_62549));
	notech_inv i_15794(.A(n_62547), .Z(n_62548));
	notech_inv i_15793(.A(n_62626), .Z(n_62547));
	notech_inv i_15792(.A(n_62545), .Z(n_62546));
	notech_inv i_15791(.A(n_62702), .Z(n_62545));
	notech_inv i_15703(.A(n_62457), .Z(n_62458));
	notech_inv i_15702(.A(n_62704), .Z(n_62457));
	notech_inv i_14328(.A(n_61356), .Z(n_61379));
	notech_inv i_14327(.A(n_61356), .Z(n_61378));
	notech_inv i_14326(.A(n_61356), .Z(n_61377));
	notech_inv i_14325(.A(n_61356), .Z(n_61376));
	notech_inv i_14324(.A(n_61356), .Z(n_61375));
	notech_inv i_14322(.A(n_61356), .Z(n_61373));
	notech_inv i_14321(.A(n_61356), .Z(n_61372));
	notech_inv i_14320(.A(n_61356), .Z(n_61371));
	notech_inv i_14319(.A(n_61356), .Z(n_61370));
	notech_inv i_14318(.A(n_61356), .Z(n_61369));
	notech_inv i_14316(.A(n_61356), .Z(n_61367));
	notech_inv i_14315(.A(n_61356), .Z(n_61366));
	notech_inv i_14314(.A(n_61356), .Z(n_61365));
	notech_inv i_14313(.A(n_61356), .Z(n_61364));
	notech_inv i_14312(.A(n_61356), .Z(n_61363));
	notech_inv i_14310(.A(n_61356), .Z(n_61361));
	notech_inv i_14309(.A(n_61356), .Z(n_61360));
	notech_inv i_14308(.A(n_61356), .Z(n_61359));
	notech_inv i_14307(.A(n_61356), .Z(n_61358));
	notech_inv i_14306(.A(n_61356), .Z(n_61357));
	notech_inv i_14305(.A(rstn), .Z(n_61356));
	notech_inv i_14304(.A(n_61350), .Z(n_61355));
	notech_inv i_14303(.A(n_61350), .Z(n_61354));
	notech_inv i_14302(.A(n_61350), .Z(n_61353));
	notech_inv i_14301(.A(n_61350), .Z(n_61352));
	notech_inv i_14300(.A(n_61350), .Z(n_61351));
	notech_inv i_14299(.A(rstn), .Z(n_61350));
	notech_inv i_13756(.A(n_141554120), .Z(n_60802));
	notech_inv i_13754(.A(n_141554120), .Z(n_60800));
	notech_inv i_13753(.A(n_141554120), .Z(n_60799));
	notech_inv i_13749(.A(n_141554120), .Z(n_60795));
	notech_inv i_13747(.A(n_141554120), .Z(n_60793));
	notech_inv i_13744(.A(n_141554120), .Z(n_60790));
	notech_inv i_13742(.A(n_141554120), .Z(n_60788));
	notech_inv i_13741(.A(n_141554120), .Z(n_60787));
	notech_inv i_13733(.A(n_60777), .Z(n_60778));
	notech_inv i_13732(.A(purge), .Z(n_60777));
	notech_inv i_13711(.A(n_60749), .Z(n_60754));
	notech_inv i_13707(.A(n_60749), .Z(n_60750));
	notech_inv i_13706(.A(pc_req), .Z(n_60749));
	notech_inv i_13693(.A(n_60641), .Z(n_60642));
	notech_inv i_13692(.A(n_141154116), .Z(n_60641));
	notech_inv i_13688(.A(n_60641), .Z(n_60637));
	notech_inv i_13684(.A(n_60641), .Z(n_60633));
	notech_inv i_13679(.A(n_60641), .Z(n_60628));
	notech_inv i_13675(.A(n_60641), .Z(n_60624));
	notech_inv i_13665(.A(n_60613), .Z(n_60614));
	notech_inv i_13664(.A(n_60594), .Z(n_60613));
	notech_inv i_13660(.A(n_60613), .Z(n_60609));
	notech_inv i_13656(.A(n_60613), .Z(n_60605));
	notech_inv i_13651(.A(n_60613), .Z(n_60600));
	notech_inv i_13647(.A(n_60613), .Z(n_60596));
	notech_inv i_13645(.A(n_60641), .Z(n_60594));
	notech_inv i_13637(.A(n_60585), .Z(n_60586));
	notech_inv i_13636(.A(n_60566), .Z(n_60585));
	notech_inv i_13632(.A(n_60585), .Z(n_60581));
	notech_inv i_13628(.A(n_60585), .Z(n_60577));
	notech_inv i_13623(.A(n_60585), .Z(n_60572));
	notech_inv i_13619(.A(n_60585), .Z(n_60568));
	notech_inv i_13617(.A(n_60641), .Z(n_60566));
	notech_inv i_13607(.A(n_60554), .Z(n_60555));
	notech_inv i_13606(.A(\nbus_93[0] ), .Z(n_60554));
	notech_inv i_13484(.A(n_140854113), .Z(n_60422));
	notech_inv i_13482(.A(n_140854113), .Z(n_60420));
	notech_inv i_13481(.A(n_140854113), .Z(n_60419));
	notech_inv i_13477(.A(n_140854113), .Z(n_60415));
	notech_inv i_13475(.A(n_140854113), .Z(n_60413));
	notech_inv i_13472(.A(n_140854113), .Z(n_60410));
	notech_inv i_13470(.A(n_140854113), .Z(n_60408));
	notech_inv i_13469(.A(n_140854113), .Z(n_60407));
	notech_inv i_12038(.A(n_58974), .Z(n_58987));
	notech_inv i_12036(.A(n_58974), .Z(n_58985));
	notech_inv i_12033(.A(n_58974), .Z(n_58982));
	notech_inv i_12031(.A(n_58974), .Z(n_58980));
	notech_inv i_12027(.A(n_58974), .Z(n_58976));
	notech_inv i_12026(.A(n_58974), .Z(n_58975));
	notech_inv i_12025(.A(n_2910), .Z(n_58974));
	notech_inv i_12023(.A(n_58955), .Z(n_58971));
	notech_inv i_12021(.A(n_58955), .Z(n_58969));
	notech_inv i_12020(.A(n_58955), .Z(n_58968));
	notech_inv i_12016(.A(n_58955), .Z(n_58964));
	notech_inv i_12014(.A(n_58955), .Z(n_58962));
	notech_inv i_12011(.A(n_58955), .Z(n_58959));
	notech_inv i_12009(.A(n_58955), .Z(n_58957));
	notech_inv i_12008(.A(n_58955), .Z(n_58956));
	notech_inv i_12007(.A(n_1277), .Z(n_58955));
	notech_inv i_12000(.A(n_58942), .Z(n_58947));
	notech_inv i_11996(.A(n_58942), .Z(n_58943));
	notech_inv i_11995(.A(n_2923), .Z(n_58942));
	notech_inv i_11992(.A(n_58923), .Z(n_58938));
	notech_inv i_11990(.A(n_58923), .Z(n_58936));
	notech_inv i_11985(.A(n_58923), .Z(n_58931));
	notech_inv i_11984(.A(n_58923), .Z(n_58930));
	notech_inv i_11978(.A(n_58923), .Z(n_58924));
	notech_inv i_11977(.A(n_1317), .Z(n_58923));
	notech_inv i_11975(.A(n_58902), .Z(n_58920));
	notech_inv i_11973(.A(n_58902), .Z(n_58918));
	notech_inv i_11970(.A(n_58902), .Z(n_58915));
	notech_inv i_11968(.A(n_58902), .Z(n_58913));
	notech_inv i_11965(.A(n_58902), .Z(n_58910));
	notech_inv i_11963(.A(n_58902), .Z(n_58908));
	notech_inv i_11960(.A(n_58902), .Z(n_58905));
	notech_inv i_11958(.A(n_58902), .Z(n_58903));
	notech_inv i_11957(.A(n_1285), .Z(n_58902));
	notech_inv i_11955(.A(n_58883), .Z(n_58899));
	notech_inv i_11953(.A(n_58883), .Z(n_58897));
	notech_inv i_11952(.A(n_58883), .Z(n_58896));
	notech_inv i_11948(.A(n_58883), .Z(n_58892));
	notech_inv i_11946(.A(n_58883), .Z(n_58890));
	notech_inv i_11943(.A(n_58883), .Z(n_58887));
	notech_inv i_11941(.A(n_58883), .Z(n_58885));
	notech_inv i_11940(.A(n_58883), .Z(n_58884));
	notech_inv i_11939(.A(n_1290), .Z(n_58883));
	notech_inv i_11937(.A(n_58864), .Z(n_58880));
	notech_inv i_11935(.A(n_58864), .Z(n_58878));
	notech_inv i_11934(.A(n_58864), .Z(n_58877));
	notech_inv i_11930(.A(n_58864), .Z(n_58873));
	notech_inv i_11928(.A(n_58864), .Z(n_58871));
	notech_inv i_11925(.A(n_58864), .Z(n_58868));
	notech_inv i_11923(.A(n_58864), .Z(n_58866));
	notech_inv i_11922(.A(n_58864), .Z(n_58865));
	notech_inv i_11921(.A(n_1280), .Z(n_58864));
	notech_inv i_11919(.A(n_58845), .Z(n_58861));
	notech_inv i_11917(.A(n_58845), .Z(n_58859));
	notech_inv i_11916(.A(n_58845), .Z(n_58858));
	notech_inv i_11912(.A(n_58845), .Z(n_58854));
	notech_inv i_11910(.A(n_58845), .Z(n_58852));
	notech_inv i_11907(.A(n_58845), .Z(n_58849));
	notech_inv i_11905(.A(n_58845), .Z(n_58847));
	notech_inv i_11904(.A(n_58845), .Z(n_58846));
	notech_inv i_11903(.A(n_1275), .Z(n_58845));
	notech_inv i_11896(.A(n_58832), .Z(n_58837));
	notech_inv i_11892(.A(n_58832), .Z(n_58833));
	notech_inv i_11891(.A(n_2046), .Z(n_58832));
	notech_inv i_11889(.A(n_58816), .Z(n_58829));
	notech_inv i_11887(.A(n_58816), .Z(n_58827));
	notech_inv i_11883(.A(n_58816), .Z(n_58823));
	notech_inv i_11882(.A(n_58816), .Z(n_58822));
	notech_inv i_11876(.A(n_1313), .Z(n_58816));
	notech_inv i_11869(.A(n_58803), .Z(n_58808));
	notech_inv i_11865(.A(n_58803), .Z(n_58804));
	notech_inv i_11864(.A(n_42899), .Z(n_58803));
	notech_inv i_11862(.A(n_58782), .Z(n_58800));
	notech_inv i_11860(.A(n_58782), .Z(n_58798));
	notech_inv i_11857(.A(n_58782), .Z(n_58795));
	notech_inv i_11855(.A(n_58782), .Z(n_58793));
	notech_inv i_11852(.A(n_58782), .Z(n_58790));
	notech_inv i_11850(.A(n_58782), .Z(n_58788));
	notech_inv i_11847(.A(n_58782), .Z(n_58785));
	notech_inv i_11845(.A(n_58782), .Z(n_58783));
	notech_inv i_11844(.A(n_1292), .Z(n_58782));
	notech_inv i_11842(.A(n_58761), .Z(n_58779));
	notech_inv i_11840(.A(n_58761), .Z(n_58777));
	notech_inv i_11837(.A(n_58761), .Z(n_58774));
	notech_inv i_11835(.A(n_58761), .Z(n_58772));
	notech_inv i_11832(.A(n_58761), .Z(n_58769));
	notech_inv i_11830(.A(n_58761), .Z(n_58767));
	notech_inv i_11827(.A(n_58761), .Z(n_58764));
	notech_inv i_11825(.A(n_58761), .Z(n_58762));
	notech_inv i_11824(.A(n_1302), .Z(n_58761));
	notech_inv i_11822(.A(n_58740), .Z(n_58758));
	notech_inv i_11820(.A(n_58740), .Z(n_58756));
	notech_inv i_11817(.A(n_58740), .Z(n_58753));
	notech_inv i_11815(.A(n_58740), .Z(n_58751));
	notech_inv i_11812(.A(n_58740), .Z(n_58748));
	notech_inv i_11810(.A(n_58740), .Z(n_58746));
	notech_inv i_11807(.A(n_58740), .Z(n_58743));
	notech_inv i_11805(.A(n_58740), .Z(n_58741));
	notech_inv i_11804(.A(n_1310), .Z(n_58740));
	notech_inv i_11802(.A(n_58719), .Z(n_58737));
	notech_inv i_11800(.A(n_58719), .Z(n_58735));
	notech_inv i_11797(.A(n_58719), .Z(n_58732));
	notech_inv i_11795(.A(n_58719), .Z(n_58730));
	notech_inv i_11792(.A(n_58719), .Z(n_58727));
	notech_inv i_11790(.A(n_58719), .Z(n_58725));
	notech_inv i_11787(.A(n_58719), .Z(n_58722));
	notech_inv i_11785(.A(n_58719), .Z(n_58720));
	notech_inv i_11784(.A(n_1297), .Z(n_58719));
	notech_inv i_11782(.A(n_58703), .Z(n_58716));
	notech_inv i_11780(.A(n_58703), .Z(n_58714));
	notech_inv i_11777(.A(n_58703), .Z(n_58711));
	notech_inv i_11775(.A(n_58703), .Z(n_58709));
	notech_inv i_11771(.A(n_58703), .Z(n_58705));
	notech_inv i_11769(.A(n_2886), .Z(n_58703));
	notech_inv i_11762(.A(n_58690), .Z(n_58695));
	notech_inv i_11758(.A(n_58690), .Z(n_58691));
	notech_inv i_11757(.A(n_2048), .Z(n_58690));
	notech_inv i_11750(.A(n_58677), .Z(n_58682));
	notech_inv i_11746(.A(n_58677), .Z(n_58678));
	notech_inv i_11745(.A(n_2047), .Z(n_58677));
	notech_inv i_11741(.A(n_58666), .Z(n_58672));
	notech_inv i_11736(.A(n_58666), .Z(n_58667));
	notech_inv i_11735(.A(n_2889), .Z(n_58666));
	notech_inv i_11733(.A(n_58645), .Z(n_58663));
	notech_inv i_11731(.A(n_58645), .Z(n_58661));
	notech_inv i_11728(.A(n_58645), .Z(n_58658));
	notech_inv i_11726(.A(n_58645), .Z(n_58656));
	notech_inv i_11723(.A(n_58645), .Z(n_58653));
	notech_inv i_11721(.A(n_58645), .Z(n_58651));
	notech_inv i_11718(.A(n_58645), .Z(n_58648));
	notech_inv i_11716(.A(n_58645), .Z(n_58646));
	notech_inv i_11715(.A(n_1287), .Z(n_58645));
	notech_inv i_11713(.A(n_58624), .Z(n_58642));
	notech_inv i_11711(.A(n_58624), .Z(n_58640));
	notech_inv i_11708(.A(n_58624), .Z(n_58637));
	notech_inv i_11706(.A(n_58624), .Z(n_58635));
	notech_inv i_11703(.A(n_58624), .Z(n_58632));
	notech_inv i_11701(.A(n_58624), .Z(n_58630));
	notech_inv i_11698(.A(n_58624), .Z(n_58627));
	notech_inv i_11696(.A(n_58624), .Z(n_58625));
	notech_inv i_11695(.A(n_1308), .Z(n_58624));
	notech_inv i_11693(.A(n_58605), .Z(n_58621));
	notech_inv i_11691(.A(n_58605), .Z(n_58619));
	notech_inv i_11690(.A(n_58605), .Z(n_58618));
	notech_inv i_11686(.A(n_58605), .Z(n_58614));
	notech_inv i_11684(.A(n_58605), .Z(n_58612));
	notech_inv i_11681(.A(n_58605), .Z(n_58609));
	notech_inv i_11679(.A(n_58605), .Z(n_58607));
	notech_inv i_11678(.A(n_58605), .Z(n_58606));
	notech_inv i_11677(.A(n_1304), .Z(n_58605));
	notech_inv i_11536(.A(n_58434), .Z(n_58447));
	notech_inv i_11534(.A(n_58434), .Z(n_58445));
	notech_inv i_11530(.A(n_58434), .Z(n_58441));
	notech_inv i_11524(.A(n_58434), .Z(n_58435));
	notech_inv i_11523(.A(n_1299), .Z(n_58434));
	notech_inv i_8527(.A(n_55169), .Z(n_55187));
	notech_inv i_8525(.A(n_55169), .Z(n_55185));
	notech_inv i_8522(.A(n_55169), .Z(n_55182));
	notech_inv i_8520(.A(n_55169), .Z(n_55180));
	notech_inv i_8517(.A(n_55169), .Z(n_55177));
	notech_inv i_8515(.A(n_55169), .Z(n_55175));
	notech_inv i_8512(.A(n_55169), .Z(n_55172));
	notech_inv i_8510(.A(n_55169), .Z(n_55170));
	notech_inv i_8509(.A(n_3780), .Z(n_55169));
	notech_inv i_8507(.A(n_55148), .Z(n_55166));
	notech_inv i_8505(.A(n_55148), .Z(n_55164));
	notech_inv i_8502(.A(n_55148), .Z(n_55161));
	notech_inv i_8500(.A(n_55148), .Z(n_55159));
	notech_inv i_8497(.A(n_55148), .Z(n_55156));
	notech_inv i_8495(.A(n_55148), .Z(n_55154));
	notech_inv i_8492(.A(n_55148), .Z(n_55151));
	notech_inv i_8490(.A(n_55148), .Z(n_55149));
	notech_inv i_8489(.A(n_3779), .Z(n_55148));
	notech_inv i_8487(.A(n_55127), .Z(n_55145));
	notech_inv i_8485(.A(n_55127), .Z(n_55143));
	notech_inv i_8482(.A(n_55127), .Z(n_55140));
	notech_inv i_8480(.A(n_55127), .Z(n_55138));
	notech_inv i_8477(.A(n_55127), .Z(n_55135));
	notech_inv i_8475(.A(n_55127), .Z(n_55133));
	notech_inv i_8472(.A(n_55127), .Z(n_55130));
	notech_inv i_8470(.A(n_55127), .Z(n_55128));
	notech_inv i_8469(.A(n_8165), .Z(n_55127));
	notech_and3 i_164577879(.A(n_2670), .B(n_2669), .C(n_1699), .Z(n_2672)
		);
	notech_ao4 i_164277882(.A(n_58968), .B(n_43060), .C(n_58774), .D(n_43091
		), .Z(n_2673));
	notech_ao4 i_164377881(.A(n_42963), .B(n_42899), .C(n_58795), .D(n_43123
		), .Z(n_2674));
	notech_ao4 i_166677858(.A(n_58896), .B(n_42988), .C(n_58915), .D(n_42980
		), .Z(n_2677));
	notech_ao4 i_166877856(.A(n_58753), .B(n_42996), .C(n_58732), .D(n_43012
		), .Z(n_2679));
	notech_ao4 i_167577849(.A(n_2048), .B(n_43046), .C(n_2047), .D(n_43109),
		 .Z(n_2681));
	notech_and4 i_167877846(.A(n_2677), .B(n_2679), .C(n_2681), .D(n_1702), 
		.Z(n_2682));
	notech_ao4 i_166977855(.A(n_58858), .B(n_43036), .C(n_58637), .D(n_43004
		), .Z(n_2683));
	notech_ao4 i_167077854(.A(n_58658), .B(n_43020), .C(n_58877), .D(n_43028
		), .Z(n_2684));
	notech_and3 i_167677848(.A(n_2684), .B(n_2683), .C(n_1715), .Z(n_2686)
		);
	notech_ao4 i_167377851(.A(n_58968), .B(n_43062), .C(n_58774), .D(n_43093
		), .Z(n_2687));
	notech_ao4 i_167477850(.A(n_42964), .B(n_42899), .C(n_58795), .D(n_43125
		), .Z(n_2688));
	notech_ao4 i_170977827(.A(n_58896), .B(n_42989), .C(n_58915), .D(n_42981
		), .Z(n_2691));
	notech_ao4 i_171177825(.A(n_58753), .B(n_42997), .C(n_58732), .D(n_43013
		), .Z(n_2693));
	notech_ao4 i_171877818(.A(n_2048), .B(n_43048), .C(n_2047), .D(n_43111),
		 .Z(n_2695));
	notech_and4 i_172177815(.A(n_2691), .B(n_2693), .C(n_2695), .D(n_1718), 
		.Z(n_2696));
	notech_ao4 i_171277824(.A(n_58858), .B(n_43037), .C(n_58637), .D(n_43005
		), .Z(n_2697));
	notech_ao4 i_171377823(.A(n_58658), .B(n_43021), .C(n_58877), .D(n_43029
		), .Z(n_2698));
	notech_and3 i_171977817(.A(n_2698), .B(n_2697), .C(n_1731), .Z(n_2700)
		);
	notech_ao4 i_171677820(.A(n_58968), .B(n_43064), .C(n_58774), .D(n_43095
		), .Z(n_2701));
	notech_ao4 i_171777819(.A(n_42965), .B(n_58808), .C(n_58795), .D(n_43127
		), .Z(n_2702));
	notech_ao4 i_175677796(.A(n_58896), .B(n_42990), .C(n_58915), .D(n_42982
		), .Z(n_2705));
	notech_ao4 i_175977794(.A(n_58753), .B(n_42998), .C(n_58732), .D(n_43014
		), .Z(n_2707));
	notech_ao4 i_176677787(.A(n_58695), .B(n_43050), .C(n_58682), .D(n_43113
		), .Z(n_2709));
	notech_and4 i_176977784(.A(n_2705), .B(n_2707), .C(n_2709), .D(n_1734), 
		.Z(n_2710));
	notech_ao4 i_176077793(.A(n_58858), .B(n_43038), .C(n_58637), .D(n_43006
		), .Z(n_2711));
	notech_ao4 i_176177792(.A(n_58658), .B(n_43022), .C(n_58877), .D(n_43030
		), .Z(n_271296494));
	notech_and3 i_176777786(.A(n_271296494), .B(n_2711), .C(n_1747), .Z(n_2714
		));
	notech_ao4 i_176477789(.A(n_58968), .B(n_43066), .C(n_58774), .D(n_43097
		), .Z(n_2716));
	notech_ao4 i_176577788(.A(n_42966), .B(n_42899), .C(n_58795), .D(n_43129
		), .Z(n_2717));
	notech_ao4 i_178877765(.A(n_58896), .B(n_42991), .C(n_58915), .D(n_42983
		), .Z(n_2720));
	notech_ao4 i_179077763(.A(n_58753), .B(n_42999), .C(n_58732), .D(n_43015
		), .Z(n_2722));
	notech_ao4 i_179777756(.A(n_2048), .B(n_43052), .C(n_2047), .D(n_43115),
		 .Z(n_2724));
	notech_and4 i_180677753(.A(n_2720), .B(n_2722), .C(n_2724), .D(n_1750), 
		.Z(n_2725));
	notech_ao4 i_179177762(.A(n_58858), .B(n_43039), .C(n_58637), .D(n_43007
		), .Z(n_2726));
	notech_ao4 i_179277761(.A(n_58658), .B(n_43023), .C(n_58877), .D(n_43031
		), .Z(n_2727));
	notech_and3 i_180477755(.A(n_2727), .B(n_2726), .C(n_1763), .Z(n_2729)
		);
	notech_ao4 i_179577758(.A(n_58968), .B(n_43068), .C(n_58774), .D(n_43099
		), .Z(n_273096495));
	notech_ao4 i_179677757(.A(n_42967), .B(n_42899), .C(n_58795), .D(n_43131
		), .Z(n_2731));
	notech_ao4 i_182677734(.A(n_58896), .B(n_43004), .C(n_58915), .D(n_42996
		), .Z(n_2734));
	notech_ao4 i_182877732(.A(n_58753), .B(n_43012), .C(n_58732), .D(n_43028
		), .Z(n_273696496));
	notech_ao4 i_183577725(.A(n_2048), .B(n_43078), .C(n_2047), .D(n_43141),
		 .Z(n_2738));
	notech_and4 i_183877722(.A(n_2734), .B(n_273696496), .C(n_2738), .D(n_1766
		), .Z(n_2739));
	notech_ao4 i_182977731(.A(n_58858), .B(n_43062), .C(n_58637), .D(n_43020
		), .Z(n_2740));
	notech_ao4 i_183077730(.A(n_58658), .B(n_43036), .C(n_58877), .D(n_43046
		), .Z(n_2741));
	notech_and3 i_183677724(.A(n_2741), .B(n_2740), .C(n_1779), .Z(n_274396497
		));
	notech_ao4 i_183377727(.A(n_58968), .B(n_43093), .C(n_58774), .D(n_43125
		), .Z(n_2744));
	notech_ao4 i_183477726(.A(n_42980), .B(n_42899), .C(n_58795), .D(n_43156
		), .Z(n_2745));
	notech_ao4 i_194977611(.A(n_60624), .B(n_43480), .C(n_60799), .D(n_43295
		), .Z(n_2748));
	notech_ao4 i_195377607(.A(n_60624), .B(n_43479), .C(n_60799), .D(n_43293
		), .Z(n_2749));
	notech_ao4 i_195777603(.A(n_60624), .B(n_43478), .C(n_60799), .D(n_43291
		), .Z(n_2750));
	notech_ao4 i_196177599(.A(n_60624), .B(n_43477), .C(n_60799), .D(n_43289
		), .Z(n_2751));
	notech_ao4 i_196577595(.A(n_60624), .B(n_43476), .C(n_60799), .D(n_43287
		), .Z(n_2752));
	notech_ao4 i_196977591(.A(n_60624), .B(n_43475), .C(n_60799), .D(n_43285
		), .Z(n_2753));
	notech_ao4 i_197377587(.A(n_60624), .B(n_43474), .C(n_60799), .D(n_43283
		), .Z(n_2754));
	notech_ao4 i_197777583(.A(n_60624), .B(n_43473), .C(n_60799), .D(n_43281
		), .Z(n_2755));
	notech_ao4 i_198177579(.A(n_60594), .B(n_43472), .C(n_60799), .D(n_43279
		), .Z(n_2756));
	notech_ao4 i_198577575(.A(n_60594), .B(n_43471), .C(n_60799), .D(n_43277
		), .Z(n_2757));
	notech_ao4 i_198977571(.A(n_60594), .B(n_43470), .C(n_60800), .D(n_43275
		), .Z(n_2758));
	notech_ao4 i_199377567(.A(n_60594), .B(n_43469), .C(n_60800), .D(n_43273
		), .Z(n_2759));
	notech_ao4 i_199777563(.A(n_60594), .B(n_43468), .C(n_60799), .D(n_43271
		), .Z(n_2760));
	notech_ao4 i_200177559(.A(n_60624), .B(n_43467), .C(n_60799), .D(n_43269
		), .Z(n_2761));
	notech_ao4 i_200577555(.A(n_60594), .B(n_43466), .C(n_60799), .D(n_43267
		), .Z(n_2762));
	notech_ao4 i_200977551(.A(n_60594), .B(n_43465), .C(n_60799), .D(n_43265
		), .Z(n_2763));
	notech_ao4 i_201377547(.A(n_60628), .B(n_43464), .C(n_60799), .D(n_43263
		), .Z(n_2764));
	notech_ao4 i_201777543(.A(n_60628), .B(n_43463), .C(n_60795), .D(n_43261
		), .Z(n_2765));
	notech_ao4 i_202177539(.A(n_60628), .B(n_43462), .C(n_60795), .D(n_43259
		), .Z(n_2766));
	notech_ao4 i_202577535(.A(n_60628), .B(n_43461), .C(n_60795), .D(n_43257
		), .Z(n_2767));
	notech_ao4 i_202977531(.A(n_60628), .B(n_43460), .C(n_60795), .D(n_43255
		), .Z(n_2768));
	notech_ao4 i_203377527(.A(n_60628), .B(n_43459), .C(n_60795), .D(n_43253
		), .Z(n_2769));
	notech_ao4 i_203777523(.A(n_60628), .B(n_43458), .C(n_60795), .D(n_43251
		), .Z(n_2770));
	notech_ao4 i_204177519(.A(n_60628), .B(n_43457), .C(n_60795), .D(n_43249
		), .Z(n_2771));
	notech_ao4 i_204577515(.A(n_60624), .B(n_43456), .C(n_60795), .D(n_43247
		), .Z(n_2772));
	notech_ao4 i_204977511(.A(n_60624), .B(n_43455), .C(n_60799), .D(n_43245
		), .Z(n_2773));
	notech_ao4 i_205377507(.A(n_60624), .B(n_43454), .C(n_60795), .D(n_43243
		), .Z(n_2774));
	notech_ao4 i_205877502(.A(n_60799), .B(n_43241), .C(n_60624), .D(n_43453
		), .Z(n_2775));
	notech_ao4 i_206277498(.A(n_60628), .B(n_43452), .C(n_60799), .D(n_43239
		), .Z(n_2776));
	notech_ao4 i_206677494(.A(n_60628), .B(n_43451), .C(n_60795), .D(n_43237
		), .Z(n_2777));
	notech_ao4 i_207177489(.A(n_60795), .B(n_43235), .C(n_60624), .D(n_43450
		), .Z(n_2778));
	notech_ao4 i_207577485(.A(n_60624), .B(n_43449), .C(n_60795), .D(n_43233
		), .Z(n_2779));
	notech_ao4 i_207977481(.A(n_60614), .B(n_43448), .C(n_60795), .D(n_43231
		), .Z(n_2781));
	notech_ao4 i_208377477(.A(n_60614), .B(n_43447), .C(n_60800), .D(n_43229
		), .Z(n_2782));
	notech_ao4 i_208777473(.A(n_60609), .B(n_43446), .C(n_60802), .D(n_43227
		), .Z(n_2783));
	notech_ao4 i_209277468(.A(n_60802), .B(n_43225), .C(n_60614), .D(n_43445
		), .Z(n_2784));
	notech_ao4 i_209777463(.A(n_60802), .B(n_43223), .C(n_60614), .D(n_43444
		), .Z(n_2785));
	notech_ao4 i_210177459(.A(n_60614), .B(n_43443), .C(n_60802), .D(n_43221
		), .Z(n_2787));
	notech_ao4 i_210677454(.A(n_60802), .B(n_43219), .C(n_60614), .D(n_43442
		), .Z(n_2788));
	notech_ao4 i_211177449(.A(n_60802), .B(n_43217), .C(n_60614), .D(n_43441
		), .Z(n_2789));
	notech_ao4 i_211677444(.A(n_60802), .B(n_43215), .C(n_60609), .D(n_43440
		), .Z(n_2790));
	notech_ao4 i_212177439(.A(n_60802), .B(n_43213), .C(n_60609), .D(n_43439
		), .Z(n_2791));
	notech_ao4 i_212677434(.A(n_60802), .B(n_43211), .C(n_60609), .D(n_43438
		), .Z(n_2793));
	notech_ao4 i_213177429(.A(n_60802), .B(n_43209), .C(n_60609), .D(n_43437
		), .Z(n_2794));
	notech_ao4 i_213677424(.A(n_60802), .B(n_43207), .C(n_60609), .D(n_43436
		), .Z(n_2796));
	notech_ao4 i_214177419(.A(n_60802), .B(n_43205), .C(n_60609), .D(n_43435
		), .Z(n_2797));
	notech_ao4 i_214677414(.A(n_60802), .B(n_43203), .C(n_60609), .D(n_43434
		), .Z(n_2799));
	notech_ao4 i_215477406(.A(n_60609), .B(n_43432), .C(n_60802), .D(n_43200
		), .Z(n_2800));
	notech_ao4 i_215877402(.A(n_60594), .B(n_43431), .C(n_60802), .D(n_43198
		), .Z(n_2801));
	notech_ao4 i_216277398(.A(n_60594), .B(n_43430), .C(n_60802), .D(n_43196
		), .Z(n_2802));
	notech_ao4 i_216677394(.A(n_60594), .B(n_43429), .C(n_60802), .D(n_43194
		), .Z(n_2803));
	notech_ao4 i_217077390(.A(n_60594), .B(n_43428), .C(n_60800), .D(n_43192
		), .Z(n_2805));
	notech_ao4 i_217477386(.A(n_60594), .B(n_43427), .C(n_60800), .D(n_43190
		), .Z(n_2806));
	notech_ao4 i_217877382(.A(n_60594), .B(n_43426), .C(n_60800), .D(n_43188
		), .Z(n_2807));
	notech_ao4 i_218277378(.A(n_60594), .B(n_43425), .C(n_60800), .D(n_43186
		), .Z(n_2808));
	notech_ao4 i_218677374(.A(n_60594), .B(n_43424), .C(n_60800), .D(n_43184
		), .Z(n_2809));
	notech_ao4 i_219077370(.A(n_60614), .B(n_43423), .C(n_60800), .D(n_43182
		), .Z(n_2811));
	notech_ao4 i_219477366(.A(n_60614), .B(n_43422), .C(n_60800), .D(n_43180
		), .Z(n_2812));
	notech_ao4 i_219877362(.A(n_60614), .B(n_43421), .C(n_60800), .D(n_43178
		), .Z(n_2813));
	notech_ao4 i_220277358(.A(n_60614), .B(n_43420), .C(n_60800), .D(n_43176
		), .Z(n_2814));
	notech_ao4 i_220677354(.A(n_60614), .B(n_43419), .C(n_60800), .D(n_43174
		), .Z(n_2815));
	notech_ao4 i_221077350(.A(n_60614), .B(n_43418), .C(n_60802), .D(n_43172
		), .Z(n_2817));
	notech_ao4 i_221477346(.A(n_60614), .B(n_43417), .C(n_60800), .D(n_43170
		), .Z(n_2818));
	notech_ao4 i_221877342(.A(n_60614), .B(n_43416), .C(n_60800), .D(n_43168
		), .Z(n_2819));
	notech_ao4 i_222277338(.A(n_60628), .B(n_43415), .C(n_60800), .D(n_43166
		), .Z(n_2820));
	notech_ao4 i_222677334(.A(n_60642), .B(n_43414), .C(n_60800), .D(n_43164
		), .Z(n_2821));
	notech_ao4 i_223477326(.A(n_60642), .B(n_43412), .C(n_60800), .D(n_43160
		), .Z(n_2823));
	notech_ao4 i_223877322(.A(n_60642), .B(n_43411), .C(n_60795), .D(n_43158
		), .Z(n_2824));
	notech_ao4 i_224677314(.A(n_60642), .B(n_43409), .C(n_60788), .D(n_43154
		), .Z(n_2825));
	notech_ao4 i_227077290(.A(n_60642), .B(n_43403), .C(n_60788), .D(n_43143
		), .Z(n_2826));
	notech_ao4 i_227477286(.A(n_60642), .B(n_43402), .C(n_60788), .D(n_43141
		), .Z(n_2827));
	notech_ao4 i_227877282(.A(n_60642), .B(n_43401), .C(n_60788), .D(n_43139
		), .Z(n_2829));
	notech_ao4 i_228277278(.A(n_60642), .B(n_43400), .C(n_60788), .D(n_43137
		), .Z(n_2830));
	notech_ao4 i_228677274(.A(n_60642), .B(n_43399), .C(n_60788), .D(n_43135
		), .Z(n_2831));
	notech_ao4 i_229077270(.A(n_60642), .B(n_43398), .C(n_60788), .D(n_43133
		), .Z(n_2832));
	notech_ao4 i_229477266(.A(n_60637), .B(n_43397), .C(n_60788), .D(n_43131
		), .Z(n_2833));
	notech_ao4 i_229877262(.A(n_60637), .B(n_43396), .C(n_60790), .D(n_43129
		), .Z(n_2835));
	notech_ao4 i_230277258(.A(n_60642), .B(n_43395), .C(n_60790), .D(n_43127
		), .Z(n_2836));
	notech_ao4 i_230677254(.A(n_60642), .B(n_43394), .C(n_60790), .D(n_43125
		), .Z(n_2837));
	notech_ao4 i_231077250(.A(n_60642), .B(n_43393), .C(n_60790), .D(n_43123
		), .Z(n_2838));
	notech_ao4 i_231477246(.A(n_60642), .B(n_43392), .C(n_60788), .D(n_43121
		), .Z(n_2839));
	notech_ao4 i_231877242(.A(n_141154116), .B(n_43391), .C(n_60788), .D(n_43119
		), .Z(n_2841));
	notech_ao4 i_232277238(.A(n_141154116), .B(n_43390), .C(n_60790), .D(n_43117
		), .Z(n_2842));
	notech_ao4 i_232677234(.A(n_141154116), .B(n_43389), .C(n_60790), .D(n_43115
		), .Z(n_2843));
	notech_ao4 i_233077230(.A(n_141154116), .B(n_43388), .C(n_60788), .D(n_43113
		), .Z(n_2844));
	notech_ao4 i_233477226(.A(n_141154116), .B(n_43387), .C(n_60787), .D(n_43111
		), .Z(n_2845));
	notech_ao4 i_233877222(.A(n_141154116), .B(n_43386), .C(n_60787), .D(n_43109
		), .Z(n_2847));
	notech_ao4 i_234277218(.A(n_141154116), .B(n_43385), .C(n_60787), .D(n_43107
		), .Z(n_2848));
	notech_ao4 i_234677214(.A(n_141154116), .B(n_43384), .C(n_60787), .D(n_43105
		), .Z(n_2849));
	notech_ao4 i_235077210(.A(n_141154116), .B(n_43383), .C(n_60787), .D(n_43103
		), .Z(n_2850));
	notech_ao4 i_235477206(.A(n_141154116), .B(n_43382), .C(n_60787), .D(n_43101
		), .Z(n_2851));
	notech_ao4 i_235877202(.A(n_60642), .B(n_43381), .C(n_60787), .D(n_43099
		), .Z(n_2853));
	notech_ao4 i_236277198(.A(n_141154116), .B(n_43380), .C(n_60787), .D(n_43097
		), .Z(n_2854));
	notech_ao4 i_236677194(.A(n_141154116), .B(n_43379), .C(n_60788), .D(n_43095
		), .Z(n_2855));
	notech_ao4 i_237077190(.A(n_141154116), .B(n_43378), .C(n_60788), .D(n_43093
		), .Z(n_2856));
	notech_ao4 i_237477186(.A(n_141154116), .B(n_43377), .C(n_60788), .D(n_43091
		), .Z(n_2857));
	notech_ao4 i_237877182(.A(n_141154116), .B(n_43376), .C(n_60788), .D(n_43089
		), .Z(n_2859));
	notech_ao4 i_238277178(.A(n_60633), .B(n_43375), .C(n_60788), .D(n_43087
		), .Z(n_2860));
	notech_ao4 i_239177169(.A(n_60787), .B(n_43084), .C(n_60633), .D(n_43373
		), .Z(n_2861));
	notech_ao4 i_239577165(.A(n_60633), .B(n_43372), .C(n_60788), .D(n_43082
		), .Z(n_2862));
	notech_ao4 i_239977161(.A(n_60633), .B(n_43371), .C(n_60788), .D(n_43080
		), .Z(n_2863));
	notech_ao4 i_240377157(.A(n_60633), .B(n_43370), .C(n_60790), .D(n_43078
		), .Z(n_2865));
	notech_ao4 i_240777153(.A(n_60633), .B(n_43369), .C(n_60793), .D(n_43076
		), .Z(n_2866));
	notech_ao4 i_241177149(.A(n_60633), .B(n_43368), .C(n_60793), .D(n_43074
		), .Z(n_2867));
	notech_ao4 i_241577145(.A(n_60633), .B(n_43367), .C(n_60793), .D(n_43072
		), .Z(n_2868));
	notech_ao4 i_241977141(.A(n_60628), .B(n_43366), .C(n_60793), .D(n_43070
		), .Z(n_2869));
	notech_ao4 i_242377137(.A(n_60628), .B(n_43365), .C(n_60793), .D(n_43068
		), .Z(n_2871));
	notech_ao4 i_242777133(.A(n_60628), .B(n_43364), .C(n_60793), .D(n_43066
		), .Z(n_2872));
	notech_ao4 i_243177129(.A(n_60628), .B(n_43363), .C(n_60793), .D(n_43064
		), .Z(n_2873));
	notech_ao4 i_243577125(.A(n_60633), .B(n_43362), .C(n_60793), .D(n_43062
		), .Z(n_2874));
	notech_ao4 i_243977121(.A(n_60633), .B(n_43361), .C(n_60795), .D(n_43060
		), .Z(n_2875));
	notech_ao4 i_244377117(.A(n_60633), .B(n_43360), .C(n_60795), .D(n_43058
		), .Z(n_2877));
	notech_ao4 i_244777113(.A(n_60633), .B(n_43359), .C(n_60795), .D(n_43056
		), .Z(n_2878));
	notech_ao4 i_245177109(.A(n_60637), .B(n_43358), .C(n_60795), .D(n_43054
		), .Z(n_2879));
	notech_ao4 i_245577105(.A(n_60637), .B(n_43357), .C(n_43052), .D(n_60793
		), .Z(n_2880));
	notech_ao4 i_245977101(.A(n_60637), .B(n_43356), .C(n_60793), .D(n_43050
		), .Z(n_2881));
	notech_ao4 i_246377097(.A(n_60637), .B(n_43355), .C(n_60793), .D(n_43048
		), .Z(n_2883));
	notech_ao4 i_246777093(.A(n_60637), .B(n_43354), .C(n_60793), .D(n_43046
		), .Z(n_2884));
	notech_ao4 i_247177089(.A(n_60637), .B(n_43353), .C(n_60793), .D(n_43044
		), .Z(n_2885));
	notech_and2 i_70(.A(addrshft[1]), .B(n_43296), .Z(n_2886));
	notech_and2 i_68(.A(n_43297), .B(n_43296), .Z(n_2887));
	notech_and2 i_71(.A(addrshft[0]), .B(n_43297), .Z(n_2889));
	notech_ao4 i_163977885(.A(n_58658), .B(n_43019), .C(n_58877), .D(n_43027
		), .Z(n_2670));
	notech_nao3 i_10(.A(addrshft[1]), .B(addrshft[0]), .C(n_58985), .Z(n_1277
		));
	notech_nao3 i_11(.A(n_43296), .B(n_43297), .C(n_58985), .Z(n_1280));
	notech_nao3 i_12(.A(addrshft[0]), .B(n_43297), .C(n_58982), .Z(n_1275)
		);
	notech_nao3 i_13(.A(addrshft[1]), .B(n_43296), .C(n_2923), .Z(n_1285));
	notech_nao3 i_14(.A(addrshft[1]), .B(addrshft[0]), .C(n_58947), .Z(n_1290
		));
	notech_nand2 i_2443(.A(queue[127]), .B(n_58827), .Z(n_2890));
	notech_nao3 i_2428(.A(n_58714), .B(queue[207]), .C(n_58982), .Z(n_2907)
		);
	notech_nand3 i_12825106(.A(n_2941), .B(n_2933), .C(n_2890), .Z(squeue[
		127]));
	notech_and2 i_61(.A(n_43300), .B(n_43301), .Z(n_2908));
	notech_or4 i_77(.A(addrshft[2]), .B(addrshft[4]), .C(addrshft[5]), .D(n_43299
		), .Z(n_2910));
	notech_nao3 i_1330845(.A(addrshft[1]), .B(n_43296), .C(n_58982), .Z(n_1329
		));
	notech_and4 i_80(.A(addrshft[3]), .B(addrshft[2]), .C(n_43301), .D(n_43300
		), .Z(n_2915));
	notech_or4 i_78(.A(addrshft[4]), .B(addrshft[5]), .C(addrshft[3]), .D(n_43298
		), .Z(n_2919));
	notech_and3 i_56(.A(n_2919), .B(n_58877), .C(n_58858), .Z(n_2921));
	notech_or4 i_84(.A(addrshft[4]), .B(addrshft[5]), .C(addrshft[3]), .D(addrshft
		[2]), .Z(n_2923));
	notech_nao3 i_1330800(.A(addrshft[0]), .B(n_43297), .C(n_2923), .Z(n_1317
		));
	notech_nao3 i_1330815(.A(n_43297), .B(n_43296), .C(n_2919), .Z(n_1310)
		);
	notech_nao3 i_43(.A(addrshft[0]), .B(n_43297), .C(n_2919), .Z(n_1308));
	notech_nand2 i_44(.A(n_2887), .B(n_2915), .Z(n_1304));
	notech_nao3 i_45(.A(addrshft[0]), .B(n_2915), .C(addrshft[1]), .Z(n_1302
		));
	notech_nao3 i_46(.A(addrshft[1]), .B(n_2915), .C(addrshft[0]), .Z(n_1299
		));
	notech_nao3 i_48(.A(addrshft[1]), .B(n_43296), .C(n_2919), .Z(n_1297));
	notech_nand3 i_49(.A(addrshft[1]), .B(addrshft[0]), .C(n_2915), .Z(n_1292
		));
	notech_nao3 i_51(.A(addrshft[1]), .B(addrshft[0]), .C(n_2919), .Z(n_1287
		));
	notech_ao4 i_2444(.A(n_58637), .B(n_43121), .C(n_58753), .D(n_43105), .Z
		(n_2927));
	notech_ao4 i_2445(.A(n_58774), .B(n_43247), .C(n_58618), .D(n_43231), .Z
		(n_2929));
	notech_ao4 i_2446(.A(n_58732), .B(n_43137), .C(n_58445), .D(n_43263), .Z
		(n_2931));
	notech_and4 i_2455(.A(n_2931), .B(n_2929), .C(n_2927), .D(n_2907), .Z(n_2933
		));
	notech_ao4 i_2447(.A(n_58896), .B(n_43089), .C(n_58795), .D(n_43279), .Z
		(n_2934));
	notech_ao4 i_2448(.A(n_58915), .B(n_43074), .C(n_58658), .D(n_43152), .Z
		(n_2935));
	notech_ao4 i_2449(.A(n_58877), .B(n_43168), .C(n_58936), .D(n_43058), .Z
		(n_2938));
	notech_ao4 i_2450(.A(n_58858), .B(n_43184), .C(n_58968), .D(n_43215), .Z
		(n_2939));
	notech_and4 i_2456(.A(n_2939), .B(n_2938), .C(n_2935), .D(n_2934), .Z(n_2941
		));
	notech_and2 i_170180074(.A(n_942), .B(n_937), .Z(n_4532));
	notech_ao4 i_163877886(.A(n_58858), .B(n_43035), .C(n_58637), .D(n_43003
		), .Z(n_2669));
	notech_nao3 i_159380071(.A(n_941), .B(n_2950), .C(n_42908), .Z(\nbus_93[0] 
		));
	notech_ao4 i_227155(.A(n_2945), .B(addrshft[1]), .C(n_948), .D(n_935), .Z
		(valid_len_1100256));
	notech_ao4 i_327156(.A(n_2945), .B(addrshft[2]), .C(n_948), .D(n_930), .Z
		(valid_len_2100255));
	notech_ao4 i_627159(.A(n_28356622), .B(n_43301), .C(n_924), .D(n_948), .Z
		(valid_len_5100254));
	notech_or4 i_3879313(.A(nbus_81[4]), .B(nbus_81[5]), .C(nbus_81[6]), .D(n_141254117
		), .Z(n_141154116));
	notech_ao4 i_627171(.A(n_950), .B(n_2944), .C(n_920), .D(n_43482), .Z(n_4675
		));
	notech_and3 i_579804(.A(n_43297), .B(n_43296), .C(n_43298), .Z(n_28656625
		));
	notech_or4 i_1179803(.A(addrshft[1]), .B(addrshft[0]), .C(addrshft[2]), 
		.D(addrshft[3]), .Z(n_28556624));
	notech_and4 i_164777877(.A(n_2663), .B(n_2665), .C(n_2667), .D(n_1686), 
		.Z(n_2668));
	notech_ao4 i_3479801(.A(wptr[0]), .B(n_42914), .C(n_948), .D(n_28556624)
		, .Z(n_28356622));
	notech_nand2 i_5486(.A(n_141554120), .B(n_43489), .Z(n_2944));
	notech_ao4 i_164477880(.A(n_2048), .B(n_43044), .C(n_2047), .D(n_43107),
		 .Z(n_2667));
	notech_nand2 i_330772(.A(wptr[1]), .B(n_42913), .Z(n_2945));
	notech_or4 i_2279292(.A(purge), .B(n_42907), .C(n_42897), .D(n_60754), .Z
		(n_2946));
	notech_nao3 i_7649(.A(pg_fault), .B(n_42910), .C(pc_pg_fault), .Z(n_2947
		));
	notech_ao4 i_163777887(.A(n_58753), .B(n_42995), .C(n_58732), .D(n_43011
		), .Z(n_2665));
	notech_nao3 i_4279314(.A(n_60790), .B(n_42914), .C(code_req), .Z(n_140854113
		));
	notech_and2 i_5487(.A(n_43489), .B(n_60790), .Z(n_2949));
	notech_or2 i_7479319(.A(n_951), .B(n_2946), .Z(n_2950));
	notech_nand2 i_7379350(.A(n_42914), .B(n_42913), .Z(n_2951));
	notech_ao4 i_163577889(.A(n_58915), .B(n_42979), .C(n_58896), .D(n_42987
		), .Z(n_2663));
	notech_nand2 i_5468(.A(n_62888), .B(n_2947), .Z(n_2993));
	notech_nao3 i_7653(.A(n_43481), .B(n_43482), .C(nbus_81[6]), .Z(n_141554120
		));
	notech_or2 i_7650(.A(n_8133), .B(n_42910), .Z(n_2995));
	notech_nand2 i_211487(.A(code_ack), .B(code_req), .Z(n_2997));
	notech_ao4 i_161177912(.A(n_42962), .B(n_58808), .C(n_58795), .D(n_43121
		), .Z(n_2660));
	notech_ao4 i_161077913(.A(n_58968), .B(n_43058), .C(n_58774), .D(n_43089
		), .Z(n_2659));
	notech_ao3 i_161377910(.A(n_2656), .B(n_2655), .C(n_1683), .Z(n_2658));
	notech_ao4 i_160777916(.A(n_58658), .B(n_43018), .C(n_58878), .D(n_43026
		), .Z(n_2656));
	notech_ao4 i_160677917(.A(n_58859), .B(n_43034), .C(n_58637), .D(n_43002
		), .Z(n_2655));
	notech_and4 i_161577908(.A(n_2649), .B(n_2651), .C(n_2653), .D(n_1670), 
		.Z(n_2654));
	notech_ao4 i_161277911(.A(n_58695), .B(n_43042), .C(n_58682), .D(n_43105
		), .Z(n_2653));
	notech_ao4 i_160577918(.A(n_58753), .B(n_42994), .C(n_58732), .D(n_43010
		), .Z(n_2651));
	notech_ao4 i_160377920(.A(n_58896), .B(n_42986), .C(n_58915), .D(n_42978
		), .Z(n_2649));
	notech_ao4 i_156877943(.A(n_42961), .B(n_58808), .C(n_58795), .D(n_43119
		), .Z(n_2646));
	notech_ao4 i_156777944(.A(n_58969), .B(n_43056), .C(n_58774), .D(n_43087
		), .Z(n_2645));
	notech_ao3 i_157077941(.A(n_2642), .B(n_2641), .C(n_1667), .Z(n_2644));
	notech_ao4 i_156477947(.A(n_58658), .B(n_43017), .C(n_58878), .D(n_43025
		), .Z(n_2642));
	notech_ao4 i_156377948(.A(n_58859), .B(n_43033), .C(n_58637), .D(n_43001
		), .Z(n_2641));
	notech_and4 i_157277939(.A(n_2635), .B(n_2637), .C(n_2639), .D(n_1654), 
		.Z(n_2640));
	notech_ao4 i_156977942(.A(n_58695), .B(n_43041), .C(n_58682), .D(n_43103
		), .Z(n_2639));
	notech_ao4 i_156277949(.A(n_58753), .B(n_42993), .C(n_58732), .D(n_43009
		), .Z(n_2637));
	notech_ao4 i_156077951(.A(n_58897), .B(n_42985), .C(n_58915), .D(n_42977
		), .Z(n_2635));
	notech_ao4 i_153777974(.A(n_42960), .B(n_58808), .C(n_58795), .D(n_43117
		), .Z(n_2632));
	notech_ao4 i_153677975(.A(n_58969), .B(n_43054), .C(n_58774), .D(n_43085
		), .Z(n_2631));
	notech_and3 i_153977972(.A(n_2628), .B(n_2627), .C(n_1651), .Z(n_2630)
		);
	notech_ao4 i_153377978(.A(n_58658), .B(n_43016), .C(n_58878), .D(n_43024
		), .Z(n_2628));
	notech_ao4 i_153277979(.A(n_58859), .B(n_43032), .C(n_58637), .D(n_43000
		), .Z(n_2627));
	notech_and4 i_154177970(.A(n_2621), .B(n_2623), .C(n_2625), .D(n_1638), 
		.Z(n_2626));
	notech_ao4 i_153877973(.A(n_58695), .B(n_43040), .C(n_58682), .D(n_43101
		), .Z(n_2625));
	notech_ao4 i_153177980(.A(n_58753), .B(n_42992), .C(n_58732), .D(n_43008
		), .Z(n_2623));
	notech_ao4 i_152977982(.A(n_58897), .B(n_42984), .C(n_58915), .D(n_42976
		), .Z(n_2621));
	notech_ao4 i_150678005(.A(n_42959), .B(n_58808), .C(n_58795), .D(n_43115
		), .Z(n_2618));
	notech_ao4 i_150578006(.A(n_58969), .B(n_43052), .C(n_58774), .D(n_43084
		), .Z(n_2617));
	notech_and3 i_150878003(.A(n_2614), .B(n_2613), .C(n_1635), .Z(n_2616)
		);
	notech_ao4 i_150278009(.A(n_58658), .B(n_43015), .C(n_58878), .D(n_43023
		), .Z(n_2614));
	notech_ao4 i_150178010(.A(n_58859), .B(n_43031), .C(n_58637), .D(n_42999
		), .Z(n_2613));
	notech_and4 i_151078001(.A(n_2607), .B(n_2609), .C(n_2611), .D(n_1622), 
		.Z(n_2612));
	notech_ao4 i_150778004(.A(n_58695), .B(n_43039), .C(n_58682), .D(n_43099
		), .Z(n_2611));
	notech_ao4 i_150078011(.A(n_58753), .B(n_42991), .C(n_58732), .D(n_43007
		), .Z(n_2609));
	notech_ao4 i_149778013(.A(n_58897), .B(n_42983), .C(n_58915), .D(n_42975
		), .Z(n_2607));
	notech_ao4 i_147178036(.A(n_42958), .B(n_58808), .C(n_58795), .D(n_43113
		), .Z(n_2604));
	notech_ao4 i_147078037(.A(n_58969), .B(n_43050), .C(n_58774), .D(n_43082
		), .Z(n_2603));
	notech_and3 i_147478034(.A(n_2600), .B(n_2599), .C(n_1619), .Z(n_2602)
		);
	notech_ao4 i_146778040(.A(n_58658), .B(n_43014), .C(n_58877), .D(n_43022
		), .Z(n_2600));
	notech_ao4 i_146578041(.A(n_58858), .B(n_43030), .C(n_58637), .D(n_42998
		), .Z(n_2599));
	notech_and4 i_147778032(.A(n_2593), .B(n_2595), .C(n_2597), .D(n_1606), 
		.Z(n_2598));
	notech_ao4 i_147378035(.A(n_58695), .B(n_43038), .C(n_58682), .D(n_43097
		), .Z(n_2597));
	notech_ao4 i_146478042(.A(n_58753), .B(n_42990), .C(n_58732), .D(n_43006
		), .Z(n_2595));
	notech_ao4 i_146178044(.A(n_58897), .B(n_42982), .C(n_58915), .D(n_42974
		), .Z(n_2593));
	notech_ao4 i_143178067(.A(n_42957), .B(n_58808), .C(n_58795), .D(n_43111
		), .Z(n_2590));
	notech_ao4 i_143078068(.A(n_58968), .B(n_43048), .C(n_58774), .D(n_43080
		), .Z(n_2589));
	notech_and3 i_143378065(.A(n_2586), .B(n_2585), .C(n_1603), .Z(n_2588)
		);
	notech_ao4 i_142778071(.A(n_58658), .B(n_43013), .C(n_58877), .D(n_43021
		), .Z(n_2586));
	notech_ao4 i_142678072(.A(n_58858), .B(n_43029), .C(n_58637), .D(n_42997
		), .Z(n_2585));
	notech_and4 i_143578063(.A(n_2579), .B(n_2581), .C(n_2583), .D(n_1590), 
		.Z(n_2584));
	notech_ao4 i_143278066(.A(n_58695), .B(n_43037), .C(n_58682), .D(n_43095
		), .Z(n_2583));
	notech_ao4 i_142578073(.A(n_58753), .B(n_42989), .C(n_58732), .D(n_43005
		), .Z(n_2581));
	notech_ao4 i_142378075(.A(n_58896), .B(n_42981), .C(n_58915), .D(n_42973
		), .Z(n_2579));
	notech_ao4 i_140078098(.A(n_42956), .B(n_42899), .C(n_58795), .D(n_43109
		), .Z(n_2576));
	notech_ao4 i_139978099(.A(n_58968), .B(n_43046), .C(n_58774), .D(n_43078
		), .Z(n_2575));
	notech_and3 i_140278096(.A(n_2572), .B(n_2571), .C(n_1587), .Z(n_2574)
		);
	notech_ao4 i_139678102(.A(n_58658), .B(n_43012), .C(n_58877), .D(n_43020
		), .Z(n_2572));
	notech_ao4 i_139578103(.A(n_58858), .B(n_43028), .C(n_58637), .D(n_42996
		), .Z(n_2571));
	notech_and4 i_140478094(.A(n_2565), .B(n_2567), .C(n_2569), .D(n_1574), 
		.Z(n_2570));
	notech_ao4 i_140178097(.A(n_2048), .B(n_43036), .C(n_2047), .D(n_43093),
		 .Z(n_2569));
	notech_ao4 i_139478104(.A(n_58753), .B(n_42988), .C(n_58732), .D(n_43004
		), .Z(n_2567));
	notech_ao4 i_139278106(.A(n_58896), .B(n_42980), .C(n_58915), .D(n_42972
		), .Z(n_2565));
	notech_ao4 i_136978129(.A(n_42955), .B(n_42899), .C(n_58795), .D(n_43107
		), .Z(n_2562));
	notech_ao4 i_136878130(.A(n_58968), .B(n_43044), .C(n_58774), .D(n_43076
		), .Z(n_2561));
	notech_and3 i_137178127(.A(n_2558), .B(n_2557), .C(n_1571), .Z(n_2560)
		);
	notech_ao4 i_136578133(.A(n_58658), .B(n_43011), .C(n_58877), .D(n_43019
		), .Z(n_2558));
	notech_ao4 i_136478134(.A(n_58858), .B(n_43027), .C(n_58637), .D(n_42995
		), .Z(n_2557));
	notech_and4 i_137378125(.A(n_2551), .B(n_2553), .C(n_2555), .D(n_1558), 
		.Z(n_2556));
	notech_ao4 i_137078128(.A(n_2048), .B(n_43035), .C(n_2047), .D(n_43091),
		 .Z(n_2555));
	notech_ao4 i_136378135(.A(n_58753), .B(n_42987), .C(n_58732), .D(n_43003
		), .Z(n_2553));
	notech_ao4 i_136178137(.A(n_58915), .B(n_42971), .C(n_58896), .D(n_42979
		), .Z(n_2551));
	notech_ao4 i_133878160(.A(n_42954), .B(n_42899), .C(n_58795), .D(n_43105
		), .Z(n_2548));
	notech_ao4 i_133778161(.A(n_58968), .B(n_43042), .C(n_58774), .D(n_43074
		), .Z(n_2547));
	notech_ao3 i_134078158(.A(n_2544), .B(n_2543), .C(n_1555), .Z(n_2546));
	notech_ao4 i_133478164(.A(n_58658), .B(n_43010), .C(n_58873), .D(n_43018
		), .Z(n_2544));
	notech_ao4 i_133378165(.A(n_58854), .B(n_43026), .C(n_58637), .D(n_42994
		), .Z(n_2543));
	notech_and4 i_134278156(.A(n_2537), .B(n_2539), .C(n_2541), .D(n_1542), 
		.Z(n_2542));
	notech_ao4 i_133978159(.A(n_2048), .B(n_43034), .C(n_2047), .D(n_43089),
		 .Z(n_2541));
	notech_ao4 i_133278166(.A(n_58753), .B(n_42986), .C(n_58732), .D(n_43002
		), .Z(n_2539));
	notech_ao4 i_133078168(.A(n_58896), .B(n_42978), .C(n_58915), .D(n_42970
		), .Z(n_2537));
	notech_ao4 i_130778191(.A(n_42953), .B(n_42899), .C(n_58793), .D(n_43103
		), .Z(n_2534));
	notech_ao4 i_130678192(.A(n_58964), .B(n_43041), .C(n_58772), .D(n_43072
		), .Z(n_2533));
	notech_ao3 i_130978189(.A(n_2530), .B(n_2529), .C(n_1539), .Z(n_2532));
	notech_ao4 i_130378195(.A(n_58656), .B(n_43009), .C(n_58873), .D(n_43017
		), .Z(n_2530));
	notech_ao4 i_130278196(.A(n_58854), .B(n_43025), .C(n_58635), .D(n_42993
		), .Z(n_2529));
	notech_and4 i_131178187(.A(n_2523), .B(n_2525), .C(n_2527), .D(n_1526), 
		.Z(n_2528));
	notech_ao4 i_130878190(.A(n_2048), .B(n_43033), .C(n_2047), .D(n_43087),
		 .Z(n_2527));
	notech_ao4 i_130178197(.A(n_58751), .B(n_42985), .C(n_58730), .D(n_43001
		), .Z(n_2525));
	notech_ao4 i_129978199(.A(n_58892), .B(n_42977), .C(n_58913), .D(n_42969
		), .Z(n_2523));
	notech_ao4 i_127678222(.A(n_42951), .B(n_42899), .C(n_58793), .D(n_43099
		), .Z(n_2520));
	notech_ao4 i_127578223(.A(n_58964), .B(n_43039), .C(n_58772), .D(n_43068
		), .Z(n_2519));
	notech_and3 i_127878220(.A(n_2516), .B(n_2515), .C(n_1523), .Z(n_2518)
		);
	notech_ao4 i_127278226(.A(n_58656), .B(n_43007), .C(n_58873), .D(n_43015
		), .Z(n_2516));
	notech_ao4 i_127178227(.A(n_58854), .B(n_43023), .C(n_58635), .D(n_42991
		), .Z(n_2515));
	notech_and4 i_128078218(.A(n_2509), .B(n_2511), .C(n_2513), .D(n_1510), 
		.Z(n_2514));
	notech_ao4 i_127778221(.A(n_2048), .B(n_43031), .C(n_2047), .D(n_43084),
		 .Z(n_2513));
	notech_ao4 i_127078228(.A(n_58751), .B(n_42983), .C(n_58730), .D(n_42999
		), .Z(n_2511));
	notech_ao4 i_126878230(.A(n_58892), .B(n_42975), .C(n_58913), .D(n_42967
		), .Z(n_2509));
	notech_ao4 i_124478253(.A(n_42950), .B(n_42899), .C(n_58793), .D(n_43097
		), .Z(n_2506));
	notech_ao4 i_124378254(.A(n_58964), .B(n_43038), .C(n_58772), .D(n_43066
		), .Z(n_2505));
	notech_and3 i_124678251(.A(n_2502), .B(n_2501), .C(n_1507), .Z(n_2504)
		);
	notech_ao4 i_124078257(.A(n_58656), .B(n_43006), .C(n_58873), .D(n_43014
		), .Z(n_2502));
	notech_ao4 i_123978258(.A(n_58854), .B(n_43022), .C(n_58635), .D(n_42990
		), .Z(n_2501));
	notech_and4 i_124878249(.A(n_2495), .B(n_2497), .C(n_2499), .D(n_1494), 
		.Z(n_2500));
	notech_ao4 i_124578252(.A(n_2048), .B(n_43030), .C(n_2047), .D(n_43082),
		 .Z(n_2499));
	notech_ao4 i_123878259(.A(n_58751), .B(n_42982), .C(n_58730), .D(n_42998
		), .Z(n_2497));
	notech_ao4 i_123678261(.A(n_58892), .B(n_42974), .C(n_58913), .D(n_42966
		), .Z(n_2495));
	notech_ao4 i_121378284(.A(n_42949), .B(n_42899), .C(n_58793), .D(n_43095
		), .Z(n_2492));
	notech_ao4 i_121278285(.A(n_58964), .B(n_43037), .C(n_58772), .D(n_43064
		), .Z(n_2491));
	notech_and3 i_121578282(.A(n_2488), .B(n_2487), .C(n_1491), .Z(n_2490)
		);
	notech_ao4 i_120978288(.A(n_58656), .B(n_43005), .C(n_58873), .D(n_43013
		), .Z(n_2488));
	notech_ao4 i_120878289(.A(n_58854), .B(n_43021), .C(n_58635), .D(n_42989
		), .Z(n_2487));
	notech_and4 i_121778280(.A(n_2481), .B(n_2483), .C(n_2485), .D(n_1478), 
		.Z(n_2486));
	notech_ao4 i_121478283(.A(n_2048), .B(n_43029), .C(n_2047), .D(n_43080),
		 .Z(n_2485));
	notech_ao4 i_120778290(.A(n_58751), .B(n_42981), .C(n_58730), .D(n_42997
		), .Z(n_2483));
	notech_ao4 i_120578292(.A(n_58892), .B(n_42973), .C(n_58913), .D(n_42965
		), .Z(n_2481));
	notech_ao4 i_117478315(.A(n_42948), .B(n_42899), .C(n_58793), .D(n_43093
		), .Z(n_2478));
	notech_ao4 i_117378316(.A(n_58964), .B(n_43036), .C(n_58772), .D(n_43062
		), .Z(n_2477));
	notech_and3 i_117778313(.A(n_2474), .B(n_2473), .C(n_1475), .Z(n_2476)
		);
	notech_ao4 i_116878319(.A(n_58656), .B(n_43004), .C(n_58873), .D(n_43012
		), .Z(n_2474));
	notech_ao4 i_116778320(.A(n_58854), .B(n_43020), .C(n_58635), .D(n_42988
		), .Z(n_2473));
	notech_and4 i_118078311(.A(n_2467), .B(n_2469), .C(n_2471), .D(n_1462), 
		.Z(n_2472));
	notech_ao4 i_117678314(.A(n_2048), .B(n_43028), .C(n_2047), .D(n_43078),
		 .Z(n_2471));
	notech_ao4 i_116578321(.A(n_58751), .B(n_42980), .C(n_58730), .D(n_42996
		), .Z(n_2469));
	notech_ao4 i_116278323(.A(n_58892), .B(n_42972), .C(n_58913), .D(n_42964
		), .Z(n_2467));
	notech_ao4 i_112878346(.A(n_42947), .B(n_42899), .C(n_58793), .D(n_43091
		), .Z(n_2464));
	notech_ao4 i_112678347(.A(n_58964), .B(n_43035), .C(n_58772), .D(n_43060
		), .Z(n_2463));
	notech_and3 i_113178344(.A(n_2460), .B(n_2459), .C(n_1459), .Z(n_2462)
		);
	notech_ao4 i_112278350(.A(n_58656), .B(n_43003), .C(n_58873), .D(n_43011
		), .Z(n_2460));
	notech_ao4 i_112078351(.A(n_58854), .B(n_43019), .C(n_58635), .D(n_42987
		), .Z(n_2459));
	notech_and4 i_113478342(.A(n_2453), .B(n_2455), .C(n_2457), .D(n_1446), 
		.Z(n_2458));
	notech_ao4 i_112978345(.A(n_2048), .B(n_43027), .C(n_2047), .D(n_43076),
		 .Z(n_2457));
	notech_ao4 i_111978352(.A(n_58751), .B(n_42979), .C(n_58730), .D(n_42995
		), .Z(n_2455));
	notech_ao4 i_111678354(.A(n_58913), .B(n_42963), .C(n_58892), .D(n_42971
		), .Z(n_2453));
	notech_ao4 i_108178377(.A(n_42946), .B(n_42899), .C(n_58793), .D(n_43089
		), .Z(n_2450));
	notech_ao4 i_108078378(.A(n_58964), .B(n_43034), .C(n_58772), .D(n_43058
		), .Z(n_2449));
	notech_ao3 i_108478375(.A(n_2446), .B(n_2445), .C(n_1443), .Z(n_2448));
	notech_ao4 i_107578381(.A(n_58656), .B(n_43002), .C(n_58873), .D(n_43010
		), .Z(n_2446));
	notech_ao4 i_107478382(.A(n_58854), .B(n_43018), .C(n_58635), .D(n_42986
		), .Z(n_2445));
	notech_and4 i_108778373(.A(n_2439), .B(n_2441), .C(n_2443), .D(n_1430), 
		.Z(n_2444));
	notech_ao4 i_108378376(.A(n_2048), .B(n_43026), .C(n_2047), .D(n_43074),
		 .Z(n_2443));
	notech_ao4 i_107278383(.A(n_58751), .B(n_42978), .C(n_58730), .D(n_42994
		), .Z(n_2441));
	notech_ao4 i_106978385(.A(n_58892), .B(n_42970), .C(n_58913), .D(n_42962
		), .Z(n_2439));
	notech_ao4 i_103578408(.A(n_42945), .B(n_42899), .C(n_58793), .D(n_43087
		), .Z(n_2436));
	notech_ao4 i_103378409(.A(n_58964), .B(n_43033), .C(n_58772), .D(n_43056
		), .Z(n_2435));
	notech_ao3 i_103878406(.A(n_2432), .B(n_2431), .C(n_1427), .Z(n_2434));
	notech_ao4 i_102978412(.A(n_58656), .B(n_43001), .C(n_58877), .D(n_43009
		), .Z(n_2432));
	notech_ao4 i_102778413(.A(n_58858), .B(n_43017), .C(n_58635), .D(n_42985
		), .Z(n_2431));
	notech_and4 i_104178404(.A(n_2425), .B(n_2427), .C(n_2429), .D(n_1414), 
		.Z(n_2430));
	notech_ao4 i_103678407(.A(n_2048), .B(n_43025), .C(n_2047), .D(n_43072),
		 .Z(n_2429));
	notech_ao4 i_102678414(.A(n_58751), .B(n_42977), .C(n_58730), .D(n_42993
		), .Z(n_2427));
	notech_ao4 i_102378416(.A(n_58892), .B(n_42969), .C(n_58913), .D(n_42961
		), .Z(n_2425));
	notech_ao4 i_98878439(.A(n_42943), .B(n_42899), .C(n_58793), .D(n_43084)
		, .Z(n_2422));
	notech_ao4 i_98778440(.A(n_58968), .B(n_43031), .C(n_58772), .D(n_43052)
		, .Z(n_2421));
	notech_and3 i_99178437(.A(n_2418), .B(n_2417), .C(n_1411), .Z(n_2420));
	notech_ao4 i_98278443(.A(n_58656), .B(n_42999), .C(n_58877), .D(n_43007)
		, .Z(n_2418));
	notech_ao4 i_98178444(.A(n_58858), .B(n_43015), .C(n_58635), .D(n_42983)
		, .Z(n_2417));
	notech_and4 i_99478435(.A(n_2411), .B(n_2413), .C(n_2415), .D(n_1398), .Z
		(n_2416));
	notech_ao4 i_99078438(.A(n_2048), .B(n_43023), .C(n_2047), .D(n_43068), 
		.Z(n_2415));
	notech_ao4 i_97978445(.A(n_58751), .B(n_42975), .C(n_58730), .D(n_42991)
		, .Z(n_2413));
	notech_ao4 i_97678447(.A(n_58896), .B(n_42967), .C(n_58913), .D(n_42959)
		, .Z(n_2411));
	notech_ao4 i_94278470(.A(n_42942), .B(n_42899), .C(n_58793), .D(n_43082)
		, .Z(n_240896491));
	notech_ao4 i_94078471(.A(n_58968), .B(n_43030), .C(n_58772), .D(n_43050)
		, .Z(n_240796490));
	notech_and3 i_94578468(.A(n_2404100081), .B(n_2403100082), .C(n_1395), .Z
		(n_2406100079));
	notech_ao4 i_93678474(.A(n_58656), .B(n_42998), .C(n_58877), .D(n_43006)
		, .Z(n_2404100081));
	notech_ao4 i_93478475(.A(n_58858), .B(n_43014), .C(n_58635), .D(n_42982)
		, .Z(n_2403100082));
	notech_and4 i_94878466(.A(n_2397100088), .B(n_2399100086), .C(n_2401100084
		), .D(n_1382), .Z(n_2402100083));
	notech_ao4 i_94378469(.A(n_2048), .B(n_43022), .C(n_2047), .D(n_43066), 
		.Z(n_2401100084));
	notech_ao4 i_93378476(.A(n_58751), .B(n_42974), .C(n_58730), .D(n_42990)
		, .Z(n_2399100086));
	notech_ao4 i_93078478(.A(n_58896), .B(n_42966), .C(n_58913), .D(n_42958)
		, .Z(n_2397100088));
	notech_ao4 i_89578501(.A(n_42941), .B(n_58804), .C(n_58793), .D(n_43080)
		, .Z(n_2393100091));
	notech_ao4 i_89478502(.A(n_58968), .B(n_43029), .C(n_58772), .D(n_43048)
		, .Z(n_2392100092));
	notech_and3 i_89878499(.A(n_2389100095), .B(n_2388100096), .C(n_1379), .Z
		(n_2391100093));
	notech_ao4 i_88978505(.A(n_58656), .B(n_42997), .C(n_58877), .D(n_43005)
		, .Z(n_2389100095));
	notech_ao4 i_88878506(.A(n_58858), .B(n_43013), .C(n_58635), .D(n_42981)
		, .Z(n_2388100096));
	notech_and4 i_90178497(.A(n_2382100100), .B(n_2384100098), .C(n_2386), .D
		(n_1366), .Z(n_2387));
	notech_ao4 i_89778500(.A(n_58691), .B(n_43021), .C(n_58678), .D(n_43064)
		, .Z(n_2386));
	notech_ao4 i_88678507(.A(n_58751), .B(n_42973), .C(n_58730), .D(n_42989)
		, .Z(n_2384100098));
	notech_ao4 i_88378509(.A(n_58896), .B(n_42965), .C(n_58913), .D(n_42957)
		, .Z(n_2382100100));
	notech_ao4 i_84978532(.A(n_42940), .B(n_58804), .C(n_58793), .D(n_43078)
		, .Z(n_2379100102));
	notech_ao4 i_84778533(.A(n_58968), .B(n_43028), .C(n_58772), .D(n_43046)
		, .Z(n_2378100103));
	notech_and3 i_85278530(.A(n_2375100105), .B(n_2374100106), .C(n_1363), .Z
		(n_2377100104));
	notech_ao4 i_84378536(.A(n_58656), .B(n_42996), .C(n_58873), .D(n_43004)
		, .Z(n_2375100105));
	notech_ao4 i_84178537(.A(n_58854), .B(n_43012), .C(n_58635), .D(n_42980)
		, .Z(n_2374100106));
	notech_and4 i_85578528(.A(n_2368100112), .B(n_2370100110), .C(n_2372100108
		), .D(n_1350), .Z(n_2373100107));
	notech_ao4 i_85078531(.A(n_58691), .B(n_43020), .C(n_58678), .D(n_43062)
		, .Z(n_2372100108));
	notech_ao4 i_84078538(.A(n_58751), .B(n_42972), .C(n_58730), .D(n_42988)
		, .Z(n_2370100110));
	notech_ao4 i_83778540(.A(n_58896), .B(n_42964), .C(n_58913), .D(n_42956)
		, .Z(n_2368100112));
	notech_ao4 i_77778563(.A(n_42939), .B(n_58804), .C(n_58793), .D(n_43076)
		, .Z(n_2365100115));
	notech_ao4 i_77678564(.A(n_58964), .B(n_43027), .C(n_58772), .D(n_43044)
		, .Z(n_2364100116));
	notech_and3 i_78378561(.A(n_2361100119), .B(n_236096489), .C(n_1347), .Z
		(n_2363100117));
	notech_ao4 i_77378567(.A(n_58656), .B(n_42995), .C(n_58873), .D(n_43003)
		, .Z(n_2361100119));
	notech_ao4 i_76478568(.A(n_58854), .B(n_43011), .C(n_58635), .D(n_42979)
		, .Z(n_236096489));
	notech_and4 i_78578559(.A(n_235496486), .B(n_235696487), .C(n_235896488)
		, .D(n_1334), .Z(n_2359100120));
	notech_ao4 i_77878562(.A(n_58691), .B(n_43019), .C(n_58678), .D(n_43060)
		, .Z(n_235896488));
	notech_ao4 i_76378569(.A(n_58751), .B(n_42971), .C(n_58730), .D(n_42987)
		, .Z(n_235696487));
	notech_ao4 i_75778571(.A(n_58913), .B(n_42955), .C(n_58892), .D(n_42963)
		, .Z(n_235496486));
	notech_ao4 i_73078594(.A(n_42938), .B(n_58804), .C(n_58793), .D(n_43074)
		, .Z(n_2351100124));
	notech_ao4 i_72978595(.A(n_58964), .B(n_43026), .C(n_58772), .D(n_43042)
		, .Z(n_235096484));
	notech_ao3 i_73278592(.A(n_2347100126), .B(n_234696482), .C(n_1331), .Z(n_2349100125
		));
	notech_ao4 i_72678598(.A(n_58656), .B(n_42994), .C(n_58877), .D(n_43002)
		, .Z(n_2347100126));
	notech_ao4 i_72578599(.A(n_58858), .B(n_43010), .C(n_42978), .D(n_58635)
		, .Z(n_234696482));
	notech_and4 i_73478590(.A(n_234096479), .B(n_234296480), .C(n_234496481)
		, .D(n_1316), .Z(n_2345100127));
	notech_ao4 i_73178593(.A(n_58691), .B(n_43018), .C(n_58678), .D(n_43058)
		, .Z(n_234496481));
	notech_ao4 i_72478600(.A(n_58751), .B(n_42970), .C(n_58730), .D(n_42986)
		, .Z(n_234296480));
	notech_ao4 i_72278602(.A(n_58892), .B(n_42962), .C(n_58913), .D(n_42954)
		, .Z(n_234096479));
	notech_ao4 i_69978625(.A(n_42937), .B(n_58804), .C(n_58793), .D(n_43072)
		, .Z(n_2337));
	notech_ao4 i_69878626(.A(n_58964), .B(n_43025), .C(n_58772), .D(n_43041)
		, .Z(n_2336));
	notech_ao3 i_70178623(.A(n_2333), .B(n_2332), .C(n_1312), .Z(n_2335));
	notech_ao4 i_69578629(.A(n_58656), .B(n_42993), .C(n_58877), .D(n_43001)
		, .Z(n_2333));
	notech_ao4 i_69478630(.A(n_58858), .B(n_43009), .C(n_58635), .D(n_42977)
		, .Z(n_2332));
	notech_and4 i_70378621(.A(n_2326), .B(n_2328), .C(n_2330), .D(n_1293), .Z
		(n_2331));
	notech_ao4 i_70078624(.A(n_58691), .B(n_43017), .C(n_58678), .D(n_43056)
		, .Z(n_2330));
	notech_ao4 i_69378631(.A(n_58751), .B(n_42969), .C(n_58730), .D(n_42985)
		, .Z(n_2328));
	notech_ao4 i_69178633(.A(n_58896), .B(n_42961), .C(n_58913), .D(n_42953)
		, .Z(n_2326));
	notech_ao4 i_66878656(.A(n_42936), .B(n_58804), .C(n_58793), .D(n_43070)
		, .Z(n_2323));
	notech_ao4 i_66778657(.A(n_58964), .B(n_43024), .C(n_58772), .D(n_43040)
		, .Z(n_2322));
	notech_and3 i_67078654(.A(n_2319), .B(n_2318), .C(n_1288), .Z(n_2321));
	notech_ao4 i_66478660(.A(n_58656), .B(n_42992), .C(n_58880), .D(n_43000)
		, .Z(n_2319));
	notech_ao4 i_66378661(.A(n_58861), .B(n_43008), .C(n_58635), .D(n_42976)
		, .Z(n_2318));
	notech_and4 i_67278652(.A(n_2312), .B(n_2314), .C(n_2316), .D(n_1270), .Z
		(n_2317));
	notech_ao4 i_66978655(.A(n_58691), .B(n_43016), .C(n_58678), .D(n_43054)
		, .Z(n_2316));
	notech_ao4 i_66278662(.A(n_58751), .B(n_42968), .C(n_58730), .D(n_42984)
		, .Z(n_2314));
	notech_ao4 i_66078664(.A(n_58896), .B(n_42960), .C(n_58913), .D(n_42952)
		, .Z(n_2312));
	notech_ao4 i_63678687(.A(n_58804), .B(n_42935), .C(n_58800), .D(n_43068)
		, .Z(n_2309));
	notech_ao4 i_63578688(.A(n_58971), .B(n_43023), .C(n_58779), .D(n_43039)
		, .Z(n_2308));
	notech_and3 i_63878685(.A(n_2305), .B(n_2304), .C(n_1267), .Z(n_2307));
	notech_ao4 i_63278691(.A(n_58663), .B(n_42991), .C(n_58880), .D(n_42999)
		, .Z(n_2305));
	notech_ao4 i_63178692(.A(n_58861), .B(n_43007), .C(n_58642), .D(n_42975)
		, .Z(n_2304));
	notech_and4 i_64078683(.A(n_2298), .B(n_2300), .C(n_2302), .D(n_1254), .Z
		(n_2303));
	notech_ao4 i_63778686(.A(n_58691), .B(n_43015), .C(n_58678), .D(n_43052)
		, .Z(n_2302));
	notech_ao4 i_63078693(.A(n_58758), .B(n_42967), .C(n_58737), .D(n_42983)
		, .Z(n_2300));
	notech_ao4 i_62878695(.A(n_58899), .B(n_42959), .C(n_58920), .D(n_42951)
		, .Z(n_2298));
	notech_ao4 i_60578718(.A(n_58804), .B(n_42934), .C(n_58800), .D(n_43066)
		, .Z(n_2295));
	notech_ao4 i_60478719(.A(n_58971), .B(n_43022), .C(n_58779), .D(n_43038)
		, .Z(n_2294));
	notech_and3 i_60778716(.A(n_2291), .B(n_2290), .C(n_1251), .Z(n_2293));
	notech_ao4 i_60178722(.A(n_58663), .B(n_42990), .C(n_58880), .D(n_42998)
		, .Z(n_2291));
	notech_ao4 i_60078723(.A(n_58861), .B(n_43006), .C(n_58642), .D(n_42974)
		, .Z(n_2290));
	notech_and4 i_60978714(.A(n_2284), .B(n_2286), .C(n_2288), .D(n_1238), .Z
		(n_2289));
	notech_ao4 i_60678717(.A(n_58691), .B(n_43014), .C(n_58678), .D(n_43050)
		, .Z(n_2288));
	notech_ao4 i_59978724(.A(n_58758), .B(n_42966), .C(n_58737), .D(n_42982)
		, .Z(n_2286));
	notech_ao4 i_59778726(.A(n_58899), .B(n_42958), .C(n_58920), .D(n_42950)
		, .Z(n_2284));
	notech_ao4 i_57478749(.A(n_58804), .B(n_42933), .C(n_58800), .D(n_43064)
		, .Z(n_2281));
	notech_ao4 i_57378750(.A(n_58971), .B(n_43021), .C(n_58779), .D(n_43037)
		, .Z(n_2280));
	notech_and3 i_57678747(.A(n_2277), .B(n_2276), .C(n_1235), .Z(n_2279));
	notech_ao4 i_57078753(.A(n_58663), .B(n_42989), .C(n_58880), .D(n_42997)
		, .Z(n_2277));
	notech_ao4 i_56978754(.A(n_58861), .B(n_43005), .C(n_58642), .D(n_42973)
		, .Z(n_2276));
	notech_and4 i_57878745(.A(n_2270), .B(n_2272), .C(n_2274), .D(n_1222), .Z
		(n_2275));
	notech_ao4 i_57578748(.A(n_58691), .B(n_43013), .C(n_58678), .D(n_43048)
		, .Z(n_2274));
	notech_ao4 i_56878755(.A(n_58758), .B(n_42965), .C(n_58737), .D(n_42981)
		, .Z(n_2272));
	notech_ao4 i_56678757(.A(n_58899), .B(n_42957), .C(n_58920), .D(n_42949)
		, .Z(n_2270));
	notech_ao4 i_54378780(.A(n_58804), .B(n_42932), .C(n_58800), .D(n_43062)
		, .Z(n_2267));
	notech_ao4 i_54278781(.A(n_58971), .B(n_43020), .C(n_58779), .D(n_43036)
		, .Z(n_2266));
	notech_and3 i_54578778(.A(n_2263), .B(n_2262), .C(n_1219), .Z(n_2265));
	notech_ao4 i_53978784(.A(n_58663), .B(n_42988), .C(n_58880), .D(n_42996)
		, .Z(n_2263));
	notech_ao4 i_53878785(.A(n_58861), .B(n_43004), .C(n_58642), .D(n_42972)
		, .Z(n_2262));
	notech_and4 i_54778776(.A(n_2256), .B(n_2258), .C(n_2260), .D(n_1206), .Z
		(n_2261));
	notech_ao4 i_54478779(.A(n_58691), .B(n_43012), .C(n_58678), .D(n_43046)
		, .Z(n_2260));
	notech_ao4 i_53778786(.A(n_58758), .B(n_42964), .C(n_58737), .D(n_42980)
		, .Z(n_2258));
	notech_ao4 i_53578788(.A(n_58899), .B(n_42956), .C(n_58920), .D(n_42948)
		, .Z(n_2256));
	notech_ao4 i_51278811(.A(n_42931), .B(n_58804), .C(n_58800), .D(n_43060)
		, .Z(n_2253));
	notech_ao4 i_51178812(.A(n_58971), .B(n_43019), .C(n_58779), .D(n_43035)
		, .Z(n_2252));
	notech_and3 i_51478809(.A(n_2249), .B(n_2248), .C(n_1203), .Z(n_2251));
	notech_ao4 i_50878815(.A(n_58663), .B(n_42987), .C(n_58880), .D(n_42995)
		, .Z(n_2249));
	notech_ao4 i_50778816(.A(n_58861), .B(n_43003), .C(n_58642), .D(n_42971)
		, .Z(n_2248));
	notech_and4 i_51678807(.A(n_2242), .B(n_2244), .C(n_2246), .D(n_1190), .Z
		(n_2247));
	notech_ao4 i_51378810(.A(n_58691), .B(n_43011), .C(n_58678), .D(n_43044)
		, .Z(n_2246));
	notech_ao4 i_50678817(.A(n_58758), .B(n_42963), .C(n_58737), .D(n_42979)
		, .Z(n_2244));
	notech_ao4 i_50478819(.A(n_58899), .B(n_42955), .C(n_58936), .D(n_42939)
		, .Z(n_2242));
	notech_ao4 i_48178842(.A(n_58804), .B(n_42930), .C(n_58800), .D(n_43058)
		, .Z(n_2239));
	notech_ao4 i_48078843(.A(n_58971), .B(n_43018), .C(n_58779), .D(n_43034)
		, .Z(n_2238));
	notech_ao3 i_48378840(.A(n_2235), .B(n_2234), .C(n_1187), .Z(n_2237));
	notech_ao4 i_47778846(.A(n_58663), .B(n_42986), .C(n_58880), .D(n_42994)
		, .Z(n_2235));
	notech_ao4 i_47678847(.A(n_58861), .B(n_43002), .C(n_58642), .D(n_42970)
		, .Z(n_2234));
	notech_and4 i_48578838(.A(n_2228), .B(n_2230), .C(n_2232), .D(n_1174), .Z
		(n_2233));
	notech_ao4 i_48278841(.A(n_58691), .B(n_43010), .C(n_58678), .D(n_43042)
		, .Z(n_2232));
	notech_ao4 i_47578848(.A(n_58758), .B(n_42962), .C(n_58737), .D(n_42978)
		, .Z(n_2230));
	notech_ao4 i_47378850(.A(n_58899), .B(n_42954), .C(n_58920), .D(n_42946)
		, .Z(n_2228));
	notech_ao4 i_45078873(.A(n_58804), .B(n_42929), .C(n_58800), .D(n_43054)
		, .Z(n_2225));
	notech_ao4 i_44978874(.A(n_58971), .B(n_43016), .C(n_58779), .D(n_43032)
		, .Z(n_2224));
	notech_and3 i_45278871(.A(n_2221), .B(n_2220), .C(n_1171), .Z(n_2223));
	notech_ao4 i_44678877(.A(n_58663), .B(n_42984), .C(n_58880), .D(n_42992)
		, .Z(n_2221));
	notech_ao4 i_44578878(.A(n_58861), .B(n_43000), .C(n_58642), .D(n_42968)
		, .Z(n_2220));
	notech_and4 i_45478869(.A(n_2214), .B(n_2216), .C(n_2218), .D(n_1157), .Z
		(n_2219));
	notech_ao4 i_45178872(.A(n_58691), .B(n_43008), .C(n_58678), .D(n_43040)
		, .Z(n_2218));
	notech_ao4 i_44478879(.A(n_58758), .B(n_42960), .C(n_58737), .D(n_42976)
		, .Z(n_2216));
	notech_ao4 i_44278881(.A(n_58899), .B(n_42952), .C(n_58920), .D(n_42944)
		, .Z(n_2214));
	notech_ao4 i_41978904(.A(n_58808), .B(n_42928), .C(n_58800), .D(n_43052)
		, .Z(n_2211));
	notech_ao4 i_41878905(.A(n_58971), .B(n_43015), .C(n_58779), .D(n_43031)
		, .Z(n_2210));
	notech_and3 i_42178902(.A(n_2207), .B(n_2206), .C(n_1152), .Z(n_2209));
	notech_ao4 i_41578908(.A(n_58663), .B(n_42983), .C(n_58880), .D(n_42991)
		, .Z(n_2207));
	notech_ao4 i_41478909(.A(n_58861), .B(n_42999), .C(n_58642), .D(n_42967)
		, .Z(n_2206));
	notech_and4 i_42378900(.A(n_2200), .B(n_2202), .C(n_2204), .D(n_1137), .Z
		(n_2205));
	notech_ao4 i_42078903(.A(n_58695), .B(n_43007), .C(n_58682), .D(n_43039)
		, .Z(n_2204));
	notech_ao4 i_41378910(.A(n_58758), .B(n_42959), .C(n_58737), .D(n_42975)
		, .Z(n_2202));
	notech_ao4 i_41178912(.A(n_58899), .B(n_42951), .C(n_58920), .D(n_42943)
		, .Z(n_2200));
	notech_ao4 i_38878935(.A(n_58808), .B(n_42927), .C(n_58800), .D(n_43050)
		, .Z(n_2197));
	notech_ao4 i_38778936(.A(n_58971), .B(n_43014), .C(n_58779), .D(n_43030)
		, .Z(n_2196));
	notech_and3 i_39078933(.A(n_2193), .B(n_2192), .C(n_1132), .Z(n_2195));
	notech_ao4 i_38478939(.A(n_58663), .B(n_42982), .C(n_58880), .D(n_42990)
		, .Z(n_2193));
	notech_ao4 i_38378940(.A(n_58861), .B(n_42998), .C(n_58642), .D(n_42966)
		, .Z(n_2192));
	notech_and4 i_39278931(.A(n_2186), .B(n_2188), .C(n_2190), .D(n_1119), .Z
		(n_2191));
	notech_ao4 i_38978934(.A(n_58695), .B(n_43006), .C(n_58682), .D(n_43038)
		, .Z(n_2190));
	notech_ao4 i_38278941(.A(n_58758), .B(n_42958), .C(n_58737), .D(n_42974)
		, .Z(n_2188));
	notech_ao4 i_38078943(.A(n_58899), .B(n_42950), .C(n_58920), .D(n_42942)
		, .Z(n_2186));
	notech_ao4 i_35778966(.A(n_58808), .B(n_42926), .C(n_58800), .D(n_43048)
		, .Z(n_2183));
	notech_ao4 i_35678967(.A(n_58971), .B(n_43013), .C(n_58779), .D(n_43029)
		, .Z(n_2182));
	notech_and3 i_35978964(.A(n_2179), .B(n_2178), .C(n_1116), .Z(n_2181));
	notech_ao4 i_35378970(.A(n_58663), .B(n_42981), .C(n_58880), .D(n_42989)
		, .Z(n_2179));
	notech_ao4 i_35278971(.A(n_58861), .B(n_42997), .C(n_58642), .D(n_42965)
		, .Z(n_2178));
	notech_and4 i_36178962(.A(n_2172), .B(n_2174), .C(n_2176), .D(n_1103), .Z
		(n_2177));
	notech_ao4 i_35878965(.A(n_58695), .B(n_43005), .C(n_58682), .D(n_43037)
		, .Z(n_2176));
	notech_ao4 i_35178972(.A(n_58758), .B(n_42957), .C(n_58737), .D(n_42973)
		, .Z(n_2174));
	notech_ao4 i_34978974(.A(n_58899), .B(n_42949), .C(n_58920), .D(n_42941)
		, .Z(n_2172));
	notech_ao4 i_32678997(.A(n_58808), .B(n_42925), .C(n_58800), .D(n_43046)
		, .Z(n_2169));
	notech_ao4 i_32578998(.A(n_58971), .B(n_43012), .C(n_58779), .D(n_43028)
		, .Z(n_2168));
	notech_and3 i_32878995(.A(n_2165), .B(n_2164), .C(n_1100), .Z(n_2167));
	notech_ao4 i_32279001(.A(n_58663), .B(n_42980), .C(n_58880), .D(n_42988)
		, .Z(n_2165));
	notech_ao4 i_32179002(.A(n_58861), .B(n_42996), .C(n_58642), .D(n_42964)
		, .Z(n_2164));
	notech_and4 i_33078993(.A(n_2158), .B(n_2160), .C(n_2162), .D(n_1087), .Z
		(n_2163));
	notech_ao4 i_32778996(.A(n_58695), .B(n_43004), .C(n_58682), .D(n_43036)
		, .Z(n_2162));
	notech_ao4 i_32079003(.A(n_58758), .B(n_42956), .C(n_58737), .D(n_42972)
		, .Z(n_2160));
	notech_ao4 i_31879005(.A(n_58899), .B(n_42948), .C(n_58920), .D(n_42940)
		, .Z(n_2158));
	notech_ao4 i_29579028(.A(n_42924), .B(n_58808), .C(n_58800), .D(n_43042)
		, .Z(n_2155));
	notech_ao4 i_29479029(.A(n_58971), .B(n_43010), .C(n_43026), .D(n_58779)
		, .Z(n_2154));
	notech_ao3 i_29779026(.A(n_2151), .B(n_2150), .C(n_1084), .Z(n_2153));
	notech_ao4 i_29179032(.A(n_42978), .B(n_58663), .C(n_58880), .D(n_42986)
		, .Z(n_2151));
	notech_ao4 i_29079033(.A(n_58861), .B(n_42994), .C(n_58642), .D(n_42962)
		, .Z(n_2150));
	notech_and4 i_29979024(.A(n_2144), .B(n_2146), .C(n_2148), .D(n_1071), .Z
		(n_2149));
	notech_ao4 i_29679027(.A(n_43002), .B(n_58695), .C(n_43034), .D(n_58682)
		, .Z(n_2148));
	notech_ao4 i_28979034(.A(n_58758), .B(n_42954), .C(n_58737), .D(n_42970)
		, .Z(n_2146));
	notech_ao4 i_28779036(.A(n_58899), .B(n_42946), .C(n_58920), .D(n_42938)
		, .Z(n_2144));
	notech_ao4 i_26479059(.A(n_58808), .B(n_42923), .C(n_58800), .D(n_43041)
		, .Z(n_2141));
	notech_ao4 i_26379060(.A(n_58971), .B(n_43009), .C(n_58779), .D(n_43025)
		, .Z(n_2140));
	notech_ao3 i_26679057(.A(n_2137), .B(n_2136), .C(n_1068), .Z(n_2139));
	notech_ao4 i_26079063(.A(n_58663), .B(n_42977), .C(n_58880), .D(n_42985)
		, .Z(n_2137));
	notech_ao4 i_25979064(.A(n_58861), .B(n_42993), .C(n_58642), .D(n_42961)
		, .Z(n_2136));
	notech_and4 i_26879055(.A(n_2130), .B(n_2132), .C(n_2134), .D(n_1055), .Z
		(n_2135));
	notech_ao4 i_26579058(.A(n_58695), .B(n_43001), .C(n_58682), .D(n_43033)
		, .Z(n_2134));
	notech_ao4 i_25879065(.A(n_58758), .B(n_42953), .C(n_58737), .D(n_42969)
		, .Z(n_2132));
	notech_ao4 i_25679067(.A(n_58899), .B(n_42945), .C(n_58920), .D(n_42937)
		, .Z(n_2130));
	notech_ao4 i_23379090(.A(n_58808), .B(n_42922), .C(n_58800), .D(n_43040)
		, .Z(n_2127));
	notech_ao4 i_23279091(.A(n_58971), .B(n_43008), .C(n_58779), .D(n_43024)
		, .Z(n_2126));
	notech_and3 i_23579088(.A(n_2123), .B(n_2122), .C(n_1052), .Z(n_2125));
	notech_ao4 i_22979094(.A(n_58663), .B(n_42976), .C(n_58880), .D(n_42984)
		, .Z(n_2123));
	notech_ao4 i_22879095(.A(n_58861), .B(n_42992), .C(n_58642), .D(n_42960)
		, .Z(n_2122));
	notech_and4 i_23779086(.A(n_2116), .B(n_2118), .C(n_2120), .D(n_1039), .Z
		(n_2121));
	notech_ao4 i_23479089(.A(n_58695), .B(n_43000), .C(n_58682), .D(n_43032)
		, .Z(n_2120));
	notech_ao4 i_22779096(.A(n_58758), .B(n_42952), .C(n_58737), .D(n_42968)
		, .Z(n_2118));
	notech_ao4 i_22579098(.A(n_58899), .B(n_42944), .C(n_58920), .D(n_42936)
		, .Z(n_2116));
	notech_ao4 i_20279121(.A(n_58804), .B(n_42921), .C(n_58800), .D(n_43039)
		, .Z(n_2113));
	notech_ao4 i_20179122(.A(n_58971), .B(n_43007), .C(n_58779), .D(n_43023)
		, .Z(n_2112));
	notech_and3 i_20479119(.A(n_2109), .B(n_2108), .C(n_1036), .Z(n_2111));
	notech_ao4 i_19879125(.A(n_58663), .B(n_42975), .C(n_58880), .D(n_42983)
		, .Z(n_2109));
	notech_ao4 i_19779126(.A(n_58861), .B(n_42991), .C(n_58642), .D(n_42959)
		, .Z(n_2108));
	notech_and4 i_20679117(.A(n_2102), .B(n_2104), .C(n_2106), .D(n_1023), .Z
		(n_2107));
	notech_ao4 i_20379120(.A(n_58691), .B(n_42999), .C(n_58678), .D(n_43031)
		, .Z(n_2106));
	notech_ao4 i_19679127(.A(n_58758), .B(n_42951), .C(n_58737), .D(n_42967)
		, .Z(n_2104));
	notech_ao4 i_19479129(.A(n_58899), .B(n_42943), .C(n_58920), .D(n_42935)
		, .Z(n_2102));
	notech_ao4 i_17179152(.A(n_58804), .B(n_42920), .C(n_58800), .D(n_43038)
		, .Z(n_2099));
	notech_ao4 i_17079153(.A(n_58971), .B(n_43006), .C(n_58779), .D(n_43022)
		, .Z(n_2098));
	notech_and3 i_17379150(.A(n_2095), .B(n_2094), .C(n_1020), .Z(n_2097));
	notech_ao4 i_16779156(.A(n_58663), .B(n_42974), .C(n_58878), .D(n_42982)
		, .Z(n_2095));
	notech_ao4 i_16679157(.A(n_58859), .B(n_42990), .C(n_58642), .D(n_42958)
		, .Z(n_2094));
	notech_and4 i_17579148(.A(n_2088), .B(n_2090), .C(n_2092), .D(n_1007), .Z
		(n_2093));
	notech_ao4 i_17279151(.A(n_58691), .B(n_42998), .C(n_58678), .D(n_43030)
		, .Z(n_2092));
	notech_ao4 i_16579158(.A(n_58758), .B(n_42950), .C(n_58737), .D(n_42966)
		, .Z(n_2090));
	notech_ao4 i_16379160(.A(n_58899), .B(n_42942), .C(n_58920), .D(n_42934)
		, .Z(n_2088));
	notech_ao4 i_14079183(.A(n_58808), .B(n_42919), .C(n_58798), .D(n_43037)
		, .Z(n_2085));
	notech_ao4 i_13979184(.A(n_58969), .B(n_43005), .C(n_58777), .D(n_43021)
		, .Z(n_2084));
	notech_and3 i_14279181(.A(n_2081), .B(n_2080), .C(n_1004), .Z(n_2083));
	notech_ao4 i_13679187(.A(n_58661), .B(n_42973), .C(n_58878), .D(n_42981)
		, .Z(n_2081));
	notech_ao4 i_13579188(.A(n_58859), .B(n_42989), .C(n_58640), .D(n_42957)
		, .Z(n_2080));
	notech_and4 i_14479179(.A(n_2074), .B(n_2076), .C(n_2078), .D(n_991), .Z
		(n_2079));
	notech_ao4 i_14179182(.A(n_58695), .B(n_42997), .C(n_58682), .D(n_43029)
		, .Z(n_2078));
	notech_ao4 i_13479189(.A(n_58756), .B(n_42949), .C(n_58735), .D(n_42965)
		, .Z(n_2076));
	notech_ao4 i_13279191(.A(n_58897), .B(n_42941), .C(n_58920), .D(n_42933)
		, .Z(n_2074));
	notech_ao4 i_10979214(.A(n_58808), .B(n_42918), .C(n_58798), .D(n_43036)
		, .Z(n_2071));
	notech_ao4 i_10879215(.A(n_58969), .B(n_43004), .C(n_58777), .D(n_43020)
		, .Z(n_2070));
	notech_and3 i_11179212(.A(n_2067), .B(n_2066), .C(n_988), .Z(n_2069));
	notech_ao4 i_10579218(.A(n_58661), .B(n_42972), .C(n_58878), .D(n_42980)
		, .Z(n_2067));
	notech_ao4 i_10479219(.A(n_58859), .B(n_42988), .C(n_58640), .D(n_42956)
		, .Z(n_2066));
	notech_and4 i_11379210(.A(n_2060), .B(n_2062), .C(n_2064), .D(n_975), .Z
		(n_2065));
	notech_ao4 i_11079213(.A(n_58695), .B(n_42996), .C(n_58682), .D(n_43028)
		, .Z(n_2064));
	notech_ao4 i_10379220(.A(n_58756), .B(n_42948), .C(n_58735), .D(n_42964)
		, .Z(n_2062));
	notech_ao4 i_10179222(.A(n_58897), .B(n_42940), .C(n_58918), .D(n_42932)
		, .Z(n_2060));
	notech_ao4 i_7779245(.A(n_58808), .B(n_42917), .C(n_58798), .D(n_43035),
		 .Z(n_2057));
	notech_and4 i_1079303(.A(n_58969), .B(n_2046), .C(n_1329), .D(n_42895), 
		.Z(n_1313));
	notech_ao4 i_7679246(.A(n_58969), .B(n_43003), .C(n_58777), .D(n_43019),
		 .Z(n_2056));
	notech_and3 i_7979243(.A(n_2053), .B(n_2052), .C(n_972), .Z(n_2055));
	notech_ao4 i_7079249(.A(n_58661), .B(n_42971), .C(n_58878), .D(n_42979),
		 .Z(n_2053));
	notech_ao4 i_6879250(.A(n_58859), .B(n_42987), .C(n_58640), .D(n_42955),
		 .Z(n_2052));
	notech_and4 i_8179241(.A(n_2042), .B(n_2044), .C(n_2049), .D(n_959), .Z(n_2050
		));
	notech_ao4 i_7879244(.A(n_58695), .B(n_42995), .C(n_58682), .D(n_43027),
		 .Z(n_2049));
	notech_nao3 i_1379301(.A(n_58714), .B(n_2046), .C(n_58985), .Z(n_2048)
		);
	notech_nand3 i_1279302(.A(n_58714), .B(n_58837), .C(n_2915), .Z(n_2047)
		);
	notech_and4 i_2079294(.A(n_58936), .B(n_58918), .C(n_58897), .D(n_2921),
		 .Z(n_2046));
	notech_ao4 i_6779251(.A(n_58756), .B(n_42947), .C(n_58735), .D(n_42963),
		 .Z(n_2044));
	notech_ao4 i_6479253(.A(n_58897), .B(n_42939), .C(n_58918), .D(n_42931),
		 .Z(n_2042));
	notech_or2 i_1779297(.A(pg_fault), .B(n_2037), .Z(n_2038));
	notech_nand2 i_1579299(.A(n_2396), .B(n_42903), .Z(n_2037));
	notech_nand2 i_3279282(.A(tagV[2]), .B(n_4676), .Z(n_2035));
	notech_nor2 i_1679298(.A(code_req), .B(wptr[1]), .Z(n_141254117));
	notech_nand3 i_1879296(.A(n_62888), .B(n_2947), .C(n_2995), .Z(n_2033)
		);
	notech_nand2 i_128389(.A(n_2885), .B(n_2030), .Z(n_2780));
	notech_nand2 i_246977091(.A(\queue_0[0] ), .B(n_60419), .Z(n_2030));
	notech_nand2 i_228390(.A(n_2884), .B(n_2028), .Z(n_2786));
	notech_nand2 i_246577095(.A(\queue_0[1] ), .B(n_60419), .Z(n_2028));
	notech_nand2 i_328391(.A(n_2883), .B(n_2026), .Z(n_2792));
	notech_nand2 i_246177099(.A(\queue_0[2] ), .B(n_60419), .Z(n_2026));
	notech_nand2 i_428392(.A(n_2881), .B(n_2024), .Z(n_2798));
	notech_nand2 i_245777103(.A(\queue_0[3] ), .B(n_60419), .Z(n_2024));
	notech_nand2 i_528393(.A(n_2880), .B(n_2022), .Z(n_2804));
	notech_nand2 i_245377107(.A(\queue_0[4] ), .B(n_60419), .Z(n_2022));
	notech_nand2 i_628394(.A(n_2879), .B(n_2020), .Z(n_2810));
	notech_nand2 i_244977111(.A(\queue_0[5] ), .B(n_60419), .Z(n_2020));
	notech_nand2 i_728395(.A(n_2878), .B(n_2018), .Z(n_2816));
	notech_nand2 i_244577115(.A(\queue_0[6] ), .B(n_60419), .Z(n_2018));
	notech_nand2 i_828396(.A(n_2877), .B(n_2016), .Z(n_2822));
	notech_nand2 i_244177119(.A(\queue_0[7] ), .B(n_60419), .Z(n_2016));
	notech_nand2 i_928397(.A(n_2875), .B(n_2014), .Z(n_2828));
	notech_nand2 i_243777123(.A(\queue_0[8] ), .B(n_60420), .Z(n_2014));
	notech_nand2 i_1028398(.A(n_2874), .B(n_2012), .Z(n_2834));
	notech_nand2 i_243377127(.A(\queue_0[9] ), .B(n_60419), .Z(n_2012));
	notech_nand2 i_1128399(.A(n_2873), .B(n_2010), .Z(n_2840));
	notech_nand2 i_242977131(.A(\queue_0[10] ), .B(n_60420), .Z(n_2010));
	notech_nand2 i_1228400(.A(n_2872), .B(n_2008), .Z(n_2846));
	notech_nand2 i_242577135(.A(\queue_0[11] ), .B(n_60420), .Z(n_2008));
	notech_nand2 i_1328401(.A(n_2871), .B(n_2006), .Z(n_2852));
	notech_nand2 i_242177139(.A(\queue_0[12] ), .B(n_60419), .Z(n_2006));
	notech_nand2 i_1428402(.A(n_2869), .B(n_2004), .Z(n_2858));
	notech_nand2 i_241777143(.A(\queue_0[13] ), .B(n_60419), .Z(n_2004));
	notech_nand2 i_1528403(.A(n_2868), .B(n_2002), .Z(n_2864));
	notech_nand2 i_241377147(.A(\queue_0[14] ), .B(n_60419), .Z(n_2002));
	notech_nand2 i_1628404(.A(n_2867), .B(n_2000), .Z(n_2870));
	notech_nand2 i_240977151(.A(\queue_0[15] ), .B(n_60419), .Z(n_2000));
	notech_nand2 i_1728405(.A(n_2866), .B(n_1998), .Z(n_2876));
	notech_nand2 i_240577155(.A(\queue_0[16] ), .B(n_60415), .Z(n_1998));
	notech_nand2 i_1828406(.A(n_2865), .B(n_1996), .Z(n_2882));
	notech_nand2 i_240177159(.A(\queue_0[17] ), .B(n_60415), .Z(n_1996));
	notech_nand2 i_1928407(.A(n_2863), .B(n_1994), .Z(n_2888));
	notech_nand2 i_239777163(.A(\queue_0[18] ), .B(n_60415), .Z(n_1994));
	notech_nand2 i_2028408(.A(n_2862), .B(n_1992), .Z(n_2894));
	notech_nand2 i_239377167(.A(\queue_0[19] ), .B(n_60415), .Z(n_1992));
	notech_nand2 i_2128409(.A(n_2861), .B(n_1989), .Z(n_2900));
	notech_nand2 i_238877172(.A(\queue_0[20] ), .B(n_60415), .Z(n_1989));
	notech_nand2 i_2328411(.A(n_2860), .B(n_1987), .Z(n_2912));
	notech_nand2 i_238077180(.A(\queue_0[22] ), .B(n_60415), .Z(n_1987));
	notech_nand2 i_2428412(.A(n_2859), .B(n_1985), .Z(n_2918));
	notech_nand2 i_237677184(.A(\queue_0[23] ), .B(n_60415), .Z(n_1985));
	notech_nand2 i_2528413(.A(n_2857), .B(n_1983), .Z(n_2924));
	notech_nand2 i_237277188(.A(\queue_0[24] ), .B(n_60415), .Z(n_1983));
	notech_nand2 i_2628414(.A(n_2856), .B(n_1981), .Z(n_2930));
	notech_nand2 i_236877192(.A(\queue_0[25] ), .B(n_60419), .Z(n_1981));
	notech_nand2 i_2728415(.A(n_2855), .B(n_1979), .Z(n_2936));
	notech_nand2 i_236477196(.A(\queue_0[26] ), .B(n_60419), .Z(n_1979));
	notech_nand2 i_2828416(.A(n_2854), .B(n_1977), .Z(n_2942));
	notech_nand2 i_236077200(.A(\queue_0[27] ), .B(n_60419), .Z(n_1977));
	notech_nand2 i_2928417(.A(n_2853), .B(n_1975), .Z(n_2948));
	notech_nand2 i_235677204(.A(\queue_0[28] ), .B(n_60419), .Z(n_1975));
	notech_nand2 i_3028418(.A(n_2851), .B(n_1973), .Z(n_2954));
	notech_nand2 i_235277208(.A(\queue_0[29] ), .B(n_60415), .Z(n_1973));
	notech_nand2 i_3128419(.A(n_2850), .B(n_1971), .Z(n_2960));
	notech_nand2 i_234877212(.A(\queue_0[30] ), .B(n_60415), .Z(n_1971));
	notech_nand2 i_3228420(.A(n_2849), .B(n_1969), .Z(n_2966));
	notech_nand2 i_234477216(.A(\queue_0[31] ), .B(n_60419), .Z(n_1969));
	notech_nand2 i_3328421(.A(n_2848), .B(n_1967), .Z(n_2972));
	notech_nand2 i_234077220(.A(\queue_0[32] ), .B(n_60415), .Z(n_1967));
	notech_nand2 i_3428422(.A(n_2847), .B(n_1965), .Z(n_2978));
	notech_nand2 i_233677224(.A(\queue_0[33] ), .B(n_60420), .Z(n_1965));
	notech_nand2 i_3528423(.A(n_2845), .B(n_1963), .Z(n_2984));
	notech_nand2 i_233277228(.A(\queue_0[34] ), .B(n_60422), .Z(n_1963));
	notech_nand2 i_3628424(.A(n_2844), .B(n_1961), .Z(n_2990));
	notech_nand2 i_232877232(.A(\queue_0[35] ), .B(n_60422), .Z(n_1961));
	notech_nand2 i_3728425(.A(n_2843), .B(n_1959), .Z(n_2996));
	notech_nand2 i_232477236(.A(\queue_0[36] ), .B(n_60422), .Z(n_1959));
	notech_nand2 i_3828426(.A(n_2842), .B(n_1957), .Z(n_3002));
	notech_nand2 i_232077240(.A(\queue_0[37] ), .B(n_60422), .Z(n_1957));
	notech_nand2 i_3928427(.A(n_2841), .B(n_1955), .Z(n_3008));
	notech_nand2 i_231677244(.A(\queue_0[38] ), .B(n_60422), .Z(n_1955));
	notech_nand2 i_4028428(.A(n_2839), .B(n_1953), .Z(n_3014));
	notech_nand2 i_231277248(.A(\queue_0[39] ), .B(n_60422), .Z(n_1953));
	notech_nand2 i_4128429(.A(n_2838), .B(n_1951), .Z(n_3020));
	notech_nand2 i_230877252(.A(\queue_0[40] ), .B(n_60422), .Z(n_1951));
	notech_nand2 i_4228430(.A(n_2837), .B(n_1949), .Z(n_3026));
	notech_nand2 i_230477256(.A(\queue_0[41] ), .B(n_60422), .Z(n_1949));
	notech_nand2 i_4328431(.A(n_2836), .B(n_1947), .Z(n_3032));
	notech_nand2 i_230077260(.A(\queue_0[42] ), .B(n_60422), .Z(n_1947));
	notech_nand2 i_4428432(.A(n_2835), .B(n_1945), .Z(n_3038));
	notech_nand2 i_229677264(.A(\queue_0[43] ), .B(n_60422), .Z(n_1945));
	notech_nand2 i_4528433(.A(n_2833), .B(n_1943), .Z(n_3044));
	notech_nand2 i_229277268(.A(\queue_0[44] ), .B(n_60422), .Z(n_1943));
	notech_nand2 i_4628434(.A(n_2832), .B(n_1941), .Z(n_3050));
	notech_nand2 i_228877272(.A(\queue_0[45] ), .B(n_60422), .Z(n_1941));
	notech_nand2 i_4728435(.A(n_2831), .B(n_1939), .Z(n_3056));
	notech_nand2 i_228477276(.A(\queue_0[46] ), .B(n_60422), .Z(n_1939));
	notech_nand2 i_4828436(.A(n_2830), .B(n_1937), .Z(n_3062));
	notech_nand2 i_228077280(.A(\queue_0[47] ), .B(n_60422), .Z(n_1937));
	notech_nand2 i_4928437(.A(n_2829), .B(n_1935), .Z(n_3068));
	notech_nand2 i_227677284(.A(\queue_0[48] ), .B(n_60422), .Z(n_1935));
	notech_nand2 i_5028438(.A(n_2827), .B(n_1933), .Z(n_3074));
	notech_nand2 i_227277288(.A(\queue_0[49] ), .B(n_60422), .Z(n_1933));
	notech_nand2 i_5128439(.A(n_2826), .B(n_1931), .Z(n_3080));
	notech_nand2 i_226877292(.A(\queue_0[50] ), .B(n_60420), .Z(n_1931));
	notech_nand2 i_5728445(.A(n_2825), .B(n_1929), .Z(n_3116));
	notech_nand2 i_224477316(.A(\queue_0[56] ), .B(n_60420), .Z(n_1929));
	notech_nand2 i_5928447(.A(n_2824), .B(n_1927), .Z(n_3128));
	notech_nand2 i_223677324(.A(\queue_0[58] ), .B(n_60420), .Z(n_1927));
	notech_nand2 i_6028448(.A(n_2823), .B(n_1925), .Z(n_3134));
	notech_nand2 i_223277328(.A(\queue_0[59] ), .B(n_60420), .Z(n_1925));
	notech_nand2 i_6228450(.A(n_2821), .B(n_1923), .Z(n_3146));
	notech_nand2 i_222477336(.A(\queue_0[61] ), .B(n_60420), .Z(n_1923));
	notech_nand2 i_6328451(.A(n_2820), .B(n_1921), .Z(n_3152));
	notech_nand2 i_222077340(.A(\queue_0[62] ), .B(n_60420), .Z(n_1921));
	notech_nand2 i_6428452(.A(n_2819), .B(n_1919), .Z(n_3158));
	notech_nand2 i_221677344(.A(\queue_0[63] ), .B(n_60420), .Z(n_1919));
	notech_nand2 i_6528453(.A(n_2818), .B(n_1917), .Z(n_3164));
	notech_nand2 i_221277348(.A(\queue_0[64] ), .B(n_60420), .Z(n_1917));
	notech_nand2 i_6628454(.A(n_2817), .B(n_1915), .Z(n_3170));
	notech_nand2 i_220877352(.A(\queue_0[65] ), .B(n_60420), .Z(n_1915));
	notech_nand2 i_6728455(.A(n_2815), .B(n_1913), .Z(n_3176));
	notech_nand2 i_220477356(.A(\queue_0[66] ), .B(n_60420), .Z(n_1913));
	notech_nand2 i_6828456(.A(n_2814), .B(n_1911), .Z(n_3182));
	notech_nand2 i_220077360(.A(\queue_0[67] ), .B(n_60422), .Z(n_1911));
	notech_nand2 i_6928457(.A(n_2813), .B(n_1909), .Z(n_3188));
	notech_nand2 i_219677364(.A(\queue_0[68] ), .B(n_60422), .Z(n_1909));
	notech_nand2 i_7028458(.A(n_2812), .B(n_1907), .Z(n_3194));
	notech_nand2 i_219277368(.A(\queue_0[69] ), .B(n_60420), .Z(n_1907));
	notech_nand2 i_7128459(.A(n_2811), .B(n_1905), .Z(n_3200));
	notech_nand2 i_218877372(.A(\queue_0[70] ), .B(n_60420), .Z(n_1905));
	notech_nand2 i_7228460(.A(n_2809), .B(n_1903), .Z(n_3206));
	notech_nand2 i_218477376(.A(\queue_0[71] ), .B(n_60420), .Z(n_1903));
	notech_nand2 i_7328461(.A(n_2808), .B(n_1901), .Z(n_3212));
	notech_nand2 i_218077380(.A(\queue_0[72] ), .B(n_60420), .Z(n_1901));
	notech_nand2 i_7428462(.A(n_2807), .B(n_1899), .Z(n_3218));
	notech_nand2 i_217677384(.A(\queue_0[73] ), .B(n_60408), .Z(n_1899));
	notech_nand2 i_7528463(.A(n_2806), .B(n_1897), .Z(n_3224));
	notech_nand2 i_217277388(.A(\queue_0[74] ), .B(n_60408), .Z(n_1897));
	notech_nand2 i_7628464(.A(n_2805), .B(n_1895), .Z(n_3230));
	notech_nand2 i_216877392(.A(\queue_0[75] ), .B(n_60408), .Z(n_1895));
	notech_nand2 i_7728465(.A(n_2803), .B(n_1893), .Z(n_3236));
	notech_nand2 i_216477396(.A(\queue_0[76] ), .B(n_60408), .Z(n_1893));
	notech_nand2 i_7828466(.A(n_2802), .B(n_1891), .Z(n_3242));
	notech_nand2 i_216077400(.A(\queue_0[77] ), .B(n_60408), .Z(n_1891));
	notech_nand2 i_7928467(.A(n_2801), .B(n_1889), .Z(n_3248));
	notech_nand2 i_215677404(.A(\queue_0[78] ), .B(n_60408), .Z(n_1889));
	notech_nand2 i_8028468(.A(n_2800), .B(n_1887), .Z(n_3254));
	notech_nand2 i_215277408(.A(\queue_0[79] ), .B(n_60408), .Z(n_1887));
	notech_nand2 i_8228470(.A(n_2799), .B(n_1884), .Z(n_3266));
	notech_nand2 i_214377417(.A(\queue_0[81] ), .B(n_60408), .Z(n_1884));
	notech_nand2 i_8328471(.A(n_2797), .B(n_1881), .Z(n_3272));
	notech_nand2 i_213877422(.A(\queue_0[82] ), .B(n_60410), .Z(n_1881));
	notech_nand2 i_8428472(.A(n_2796), .B(n_1878), .Z(n_3278));
	notech_nand2 i_213377427(.A(\queue_0[83] ), .B(n_60410), .Z(n_1878));
	notech_nand2 i_8528473(.A(n_2794), .B(n_1875), .Z(n_3284));
	notech_nand2 i_212877432(.A(\queue_0[84] ), .B(n_60410), .Z(n_1875));
	notech_nand2 i_8628474(.A(n_2793), .B(n_1872), .Z(n_3290));
	notech_nand2 i_212377437(.A(\queue_0[85] ), .B(n_60410), .Z(n_1872));
	notech_nand2 i_8728475(.A(n_2791), .B(n_1869), .Z(n_3296));
	notech_nand2 i_211877442(.A(\queue_0[86] ), .B(n_60410), .Z(n_1869));
	notech_nand2 i_8828476(.A(n_2790), .B(n_1866), .Z(n_3302));
	notech_nand2 i_211377447(.A(\queue_0[87] ), .B(n_60410), .Z(n_1866));
	notech_nand2 i_8928477(.A(n_2789), .B(n_1863), .Z(n_3308));
	notech_nand2 i_210877452(.A(\queue_0[88] ), .B(n_60410), .Z(n_1863));
	notech_nand2 i_9028478(.A(n_2788), .B(n_1860), .Z(n_3314));
	notech_nand2 i_210377457(.A(\queue_0[89] ), .B(n_60410), .Z(n_1860));
	notech_nand2 i_9128479(.A(n_2787), .B(n_1858), .Z(n_3320));
	notech_nand2 i_209977461(.A(\queue_0[90] ), .B(n_60407), .Z(n_1858));
	notech_nand2 i_9228480(.A(n_2785), .B(n_1855), .Z(n_3326));
	notech_nand2 i_209477466(.A(\queue_0[91] ), .B(n_60407), .Z(n_1855));
	notech_nand2 i_9328481(.A(n_2784), .B(n_1852), .Z(n_3332));
	notech_nand2 i_208977471(.A(\queue_0[92] ), .B(n_60407), .Z(n_1852));
	notech_nand2 i_9428482(.A(n_2783), .B(n_1850), .Z(n_3338));
	notech_nand2 i_208577475(.A(\queue_0[93] ), .B(n_60407), .Z(n_1850));
	notech_nand2 i_9528483(.A(n_2782), .B(n_1848), .Z(n_3344));
	notech_nand2 i_208177479(.A(\queue_0[94] ), .B(n_60407), .Z(n_1848));
	notech_nand2 i_9628484(.A(n_2781), .B(n_1846), .Z(n_3350));
	notech_nand2 i_207777483(.A(\queue_0[95] ), .B(n_60407), .Z(n_1846));
	notech_nand2 i_9728485(.A(n_2779), .B(n_1844), .Z(n_3356));
	notech_nand2 i_207377487(.A(\queue_0[96] ), .B(n_60407), .Z(n_1844));
	notech_nand2 i_9828486(.A(n_2778), .B(n_1841), .Z(n_3362));
	notech_nand2 i_206877492(.A(\queue_0[97] ), .B(n_60407), .Z(n_1841));
	notech_nand2 i_9928487(.A(n_2777), .B(n_1839), .Z(n_3368));
	notech_nand2 i_206477496(.A(\queue_0[98] ), .B(n_60408), .Z(n_1839));
	notech_nand2 i_10028488(.A(n_2776), .B(n_1837), .Z(n_3374));
	notech_nand2 i_206077500(.A(\queue_0[99] ), .B(n_60408), .Z(n_1837));
	notech_nand2 i_10128489(.A(n_2775), .B(n_1834), .Z(n_3380));
	notech_nand2 i_205577505(.A(\queue_0[100] ), .B(n_60408), .Z(n_1834));
	notech_nand2 i_10228490(.A(n_2774), .B(n_1832), .Z(n_3386));
	notech_nand2 i_205177509(.A(\queue_0[101] ), .B(n_60408), .Z(n_1832));
	notech_nand2 i_10328491(.A(n_2773), .B(n_1830), .Z(n_3392));
	notech_nand2 i_204777513(.A(\queue_0[102] ), .B(n_60408), .Z(n_1830));
	notech_nand2 i_10428492(.A(n_2772), .B(n_1828), .Z(n_3398));
	notech_nand2 i_204377517(.A(\queue_0[103] ), .B(n_60408), .Z(n_1828));
	notech_nand2 i_10528493(.A(n_2771), .B(n_1826), .Z(n_3404));
	notech_nand2 i_203977521(.A(\queue_0[104] ), .B(n_60408), .Z(n_1826));
	notech_nand2 i_10628494(.A(n_2770), .B(n_1824), .Z(n_3410));
	notech_nand2 i_203577525(.A(\queue_0[105] ), .B(n_60408), .Z(n_1824));
	notech_nand2 i_10728495(.A(n_2769), .B(n_1822), .Z(n_3416));
	notech_nand2 i_203177529(.A(\queue_0[106] ), .B(n_60410), .Z(n_1822));
	notech_nand2 i_10828496(.A(n_2768), .B(n_1820), .Z(n_3422));
	notech_nand2 i_202777533(.A(\queue_0[107] ), .B(n_60413), .Z(n_1820));
	notech_nand2 i_10928497(.A(n_2767), .B(n_1818), .Z(n_3428));
	notech_nand2 i_202377537(.A(\queue_0[108] ), .B(n_60413), .Z(n_1818));
	notech_nand2 i_11028498(.A(n_2766), .B(n_1816), .Z(n_3434));
	notech_nand2 i_201977541(.A(\queue_0[109] ), .B(n_60413), .Z(n_1816));
	notech_nand2 i_11128499(.A(n_2765), .B(n_1814), .Z(n_3440));
	notech_nand2 i_201577545(.A(\queue_0[110] ), .B(n_60413), .Z(n_1814));
	notech_nand2 i_11228500(.A(n_2764), .B(n_1812), .Z(n_3446));
	notech_nand2 i_201177549(.A(\queue_0[111] ), .B(n_60413), .Z(n_1812));
	notech_nand2 i_11328501(.A(n_2763), .B(n_1810), .Z(n_3452));
	notech_nand2 i_200777553(.A(\queue_0[112] ), .B(n_60413), .Z(n_1810));
	notech_nand2 i_11428502(.A(n_2762), .B(n_1808), .Z(n_3458));
	notech_nand2 i_200377557(.A(\queue_0[113] ), .B(n_60413), .Z(n_1808));
	notech_nand2 i_11528503(.A(n_2761), .B(n_1806), .Z(n_3464));
	notech_nand2 i_199977561(.A(\queue_0[114] ), .B(n_60413), .Z(n_1806));
	notech_nand2 i_11628504(.A(n_2760), .B(n_1804), .Z(n_3470));
	notech_nand2 i_199577565(.A(\queue_0[115] ), .B(n_60415), .Z(n_1804));
	notech_nand2 i_11728505(.A(n_2759), .B(n_1802), .Z(n_3476));
	notech_nand2 i_199177569(.A(\queue_0[116] ), .B(n_60415), .Z(n_1802));
	notech_nand2 i_11828506(.A(n_2758), .B(n_1800), .Z(n_3482));
	notech_nand2 i_198777573(.A(\queue_0[117] ), .B(n_60415), .Z(n_1800));
	notech_nand2 i_11928507(.A(n_2757), .B(n_1798), .Z(n_3488));
	notech_nand2 i_198377577(.A(\queue_0[118] ), .B(n_60415), .Z(n_1798));
	notech_nand2 i_12028508(.A(n_2756), .B(n_1796), .Z(n_3494));
	notech_nand2 i_197977581(.A(\queue_0[119] ), .B(n_60415), .Z(n_1796));
	notech_nand2 i_12128509(.A(n_2755), .B(n_1794), .Z(n_3500));
	notech_nand2 i_197577585(.A(\queue_0[120] ), .B(n_60413), .Z(n_1794));
	notech_nand2 i_12228510(.A(n_2754), .B(n_1792), .Z(n_3506));
	notech_nand2 i_197177589(.A(\queue_0[121] ), .B(n_60415), .Z(n_1792));
	notech_nand2 i_12328511(.A(n_2753), .B(n_1790), .Z(n_3512));
	notech_nand2 i_196777593(.A(\queue_0[122] ), .B(n_60415), .Z(n_1790));
	notech_nand2 i_12428512(.A(n_2752), .B(n_1788), .Z(n_3518));
	notech_nand2 i_196377597(.A(\queue_0[123] ), .B(n_60410), .Z(n_1788));
	notech_nand2 i_12528513(.A(n_2751), .B(n_1786), .Z(n_3524));
	notech_nand2 i_195977601(.A(\queue_0[124] ), .B(n_60410), .Z(n_1786));
	notech_nand2 i_12628514(.A(n_2750), .B(n_1784), .Z(n_3530));
	notech_nand2 i_195577605(.A(\queue_0[125] ), .B(n_60413), .Z(n_1784));
	notech_nand2 i_12728515(.A(n_2749), .B(n_1782), .Z(n_3536));
	notech_nand2 i_195177609(.A(\queue_0[126] ), .B(n_60410), .Z(n_1782));
	notech_nand2 i_12828516(.A(n_2748), .B(n_1780), .Z(n_3542));
	notech_nand2 i_194777613(.A(\queue_0[127] ), .B(n_60410), .Z(n_1780));
	notech_and4 i_6625044(.A(n_2745), .B(n_2744), .C(n_2739), .D(n_274396497
		), .Z(squeue_65100257));
	notech_nao3 i_182577735(.A(n_2046), .B(queue[161]), .C(n_58618), .Z(n_1779
		));
	notech_nao3 i_181177748(.A(n_58672), .B(queue[73]), .C(n_2923), .Z(n_1766
		));
	notech_and4 i_5325031(.A(n_2731), .B(n_273096495), .C(n_2725), .D(n_2729
		), .Z(squeue_52100258));
	notech_nao3 i_178777766(.A(n_2046), .B(queue[148]), .C(n_58618), .Z(n_1763
		));
	notech_nao3 i_177477779(.A(n_58672), .B(queue[60]), .C(n_2923), .Z(n_1750
		));
	notech_and4 i_5225030(.A(n_2717), .B(n_2716), .C(n_2710), .D(n_2714), .Z
		(squeue_51100259));
	notech_nao3 i_175477797(.A(n_2046), .B(queue[147]), .C(n_58618), .Z(n_1747
		));
	notech_nao3 i_172677810(.A(n_58672), .B(queue[59]), .C(n_58947), .Z(n_1734
		));
	notech_and4 i_5125029(.A(n_2702), .B(n_2701), .C(n_2696), .D(n_2700), .Z
		(squeue_50100260));
	notech_nao3 i_170877828(.A(n_58837), .B(queue[146]), .C(n_58618), .Z(n_1731
		));
	notech_nao3 i_168377841(.A(n_58672), .B(queue[58]), .C(n_58947), .Z(n_1718
		));
	notech_and4 i_5025028(.A(n_2688), .B(n_2687), .C(n_2682), .D(n_2686), .Z
		(squeue_49100261));
	notech_nao3 i_166577859(.A(n_58837), .B(queue[145]), .C(n_58618), .Z(n_1715
		));
	notech_nao3 i_165277872(.A(n_58672), .B(queue[57]), .C(n_58947), .Z(n_1702
		));
	notech_and4 i_4925027(.A(n_2674), .B(n_2673), .C(n_2668), .D(n_2672), .Z
		(squeue_48100262));
	notech_nao3 i_163477890(.A(n_58837), .B(queue[144]), .C(n_58618), .Z(n_1699
		));
	notech_nao3 i_162077903(.A(n_58672), .B(queue[56]), .C(n_58947), .Z(n_1686
		));
	notech_and4 i_4825026(.A(n_2660), .B(n_2659), .C(n_2654), .D(n_2658), .Z
		(squeue_47100263));
	notech_and4 i_160277921(.A(n_2887), .B(n_2915), .C(n_58837), .D(queue[
		143]), .Z(n_1683));
	notech_or2 i_157777934(.A(n_58936), .B(n_42970), .Z(n_1670));
	notech_and4 i_4725025(.A(n_2646), .B(n_2645), .C(n_2640), .D(n_2644), .Z
		(squeue_46100264));
	notech_and4 i_155977952(.A(n_2887), .B(n_2915), .C(n_58837), .D(queue[
		142]), .Z(n_1667));
	notech_or2 i_154677965(.A(n_58936), .B(n_42969), .Z(n_1654));
	notech_and4 i_4625024(.A(n_2632), .B(n_2631), .C(n_2626), .D(n_2630), .Z
		(squeue_45100265));
	notech_nao3 i_152877983(.A(n_58837), .B(queue[141]), .C(n_58619), .Z(n_1651
		));
	notech_nao3 i_151577996(.A(n_58672), .B(queue[53]), .C(n_58947), .Z(n_1638
		));
	notech_and4 i_4525023(.A(n_2618), .B(n_2617), .C(n_2612), .D(n_2616), .Z
		(squeue_44100266));
	notech_nao3 i_149678014(.A(n_58837), .B(queue[140]), .C(n_58619), .Z(n_1635
		));
	notech_nao3 i_148278027(.A(n_58672), .B(queue[52]), .C(n_58947), .Z(n_1622
		));
	notech_and4 i_4425022(.A(n_2604), .B(n_2603), .C(n_2598), .D(n_2602), .Z
		(squeue_43100267));
	notech_nao3 i_145978045(.A(n_2046), .B(queue[139]), .C(n_58619), .Z(n_1619
		));
	notech_nao3 i_144078058(.A(n_58672), .B(queue[51]), .C(n_2923), .Z(n_1606
		));
	notech_and4 i_4325021(.A(n_2590), .B(n_2589), .C(n_2584), .D(n_2588), .Z
		(squeue_42100268));
	notech_nao3 i_142278076(.A(n_2046), .B(queue[138]), .C(n_58618), .Z(n_1603
		));
	notech_nao3 i_140978089(.A(n_58672), .B(queue[50]), .C(n_2923), .Z(n_1590
		));
	notech_and4 i_4225020(.A(n_2576), .B(n_2575), .C(n_2570), .D(n_2574), .Z
		(squeue_41100269));
	notech_nao3 i_139178107(.A(n_2046), .B(queue[137]), .C(n_58618), .Z(n_1587
		));
	notech_nao3 i_137878120(.A(n_58672), .B(queue[49]), .C(n_2923), .Z(n_1574
		));
	notech_and4 i_4125019(.A(n_2562), .B(n_2561), .C(n_2556), .D(n_2560), .Z
		(squeue_40100270));
	notech_nao3 i_136078138(.A(n_2046), .B(queue[136]), .C(n_58618), .Z(n_1571
		));
	notech_nao3 i_134778151(.A(n_58672), .B(queue[48]), .C(n_2923), .Z(n_1558
		));
	notech_and4 i_4025018(.A(n_2548), .B(n_2547), .C(n_2542), .D(n_2546), .Z
		(squeue_39100271));
	notech_and4 i_132978169(.A(n_2887), .B(n_2915), .C(n_2046), .D(queue[135
		]), .Z(n_1555));
	notech_or2 i_131678182(.A(n_58936), .B(n_42962), .Z(n_1542));
	notech_and4 i_3925017(.A(n_2534), .B(n_2533), .C(n_2528), .D(n_2532), .Z
		(squeue_38100272));
	notech_and4 i_129878200(.A(n_2887), .B(n_2915), .C(n_2046), .D(queue[134
		]), .Z(n_1539));
	notech_or2 i_128578213(.A(n_58936), .B(n_42961), .Z(n_1526));
	notech_and4 i_3725015(.A(n_2520), .B(n_2519), .C(n_2514), .D(n_2518), .Z
		(squeue_36100273));
	notech_nao3 i_126778231(.A(n_2046), .B(queue[132]), .C(n_58618), .Z(n_1523
		));
	notech_nao3 i_125378244(.A(n_58672), .B(queue[44]), .C(n_2923), .Z(n_1510
		));
	notech_and4 i_3625014(.A(n_2506), .B(n_2505), .C(n_2500), .D(n_2504), .Z
		(squeue_35100274));
	notech_nao3 i_123578262(.A(n_2046), .B(queue[131]), .C(n_58618), .Z(n_1507
		));
	notech_nao3 i_122278275(.A(n_58672), .B(queue[43]), .C(n_2923), .Z(n_1494
		));
	notech_and4 i_3525013(.A(n_2492), .B(n_2491), .C(n_2486), .D(n_2490), .Z
		(squeue_34100275));
	notech_nao3 i_120478293(.A(n_2046), .B(queue[130]), .C(n_58614), .Z(n_1491
		));
	notech_nand3 i_26979568(.A(n_2037), .B(n_8137), .C(n_8133), .Z(n_133997809
		));
	notech_or4 i_3779798(.A(useq_ptr[3]), .B(useq_ptr[2]), .C(useq_ptr[1]), 
		.D(useq_ptr[0]), .Z(n_134097810));
	notech_nand3 i_27479563(.A(n_62888), .B(n_2947), .C(n_42897), .Z(n_134197811
		));
	notech_nao3 i_27079567(.A(n_60790), .B(n_134097810), .C(n_2946), .Z(n_134297812
		));
	notech_mux2 i_222655(.S(n_136597835), .A(n_2949), .B(n_42898), .Z(n_134997819
		));
	notech_nand2 i_214877412(.A(n_60410), .B(\queue_0[80] ), .Z(n_135097820)
		);
	notech_nand2 i_8128469(.A(n_136697836), .B(n_135097820), .Z(n_135297822)
		);
	notech_nand2 i_225677304(.A(n_60410), .B(\queue_0[53] ), .Z(n_135397823)
		);
	notech_nand2 i_5428442(.A(n_136797837), .B(n_135397823), .Z(n_135597825)
		);
	notech_nand2 i_226477296(.A(n_60410), .B(\queue_0[51] ), .Z(n_135697826)
		);
	notech_nand2 i_5228440(.A(n_136897838), .B(n_135697826), .Z(n_135897828)
		);
	notech_nand2 i_238477176(.A(n_60413), .B(\queue_0[21] ), .Z(n_135997829)
		);
	notech_nand2 i_2228410(.A(n_136997839), .B(n_135997829), .Z(n_136197831)
		);
	notech_xor2 i_2379291(.A(n_42914), .B(wptr[0]), .Z(n_136597835));
	notech_ao4 i_215077410(.A(n_60637), .B(n_43433), .C(n_60790), .D(n_43201
		), .Z(n_136697836));
	notech_ao4 i_225877302(.A(n_60790), .B(n_43148), .C(n_60637), .D(n_43406
		), .Z(n_136797837));
	notech_ao4 i_226677294(.A(n_60633), .B(n_43404), .C(n_60790), .D(n_43144
		), .Z(n_136897838));
	notech_ao4 i_238677174(.A(n_60637), .B(n_43374), .C(n_60790), .D(n_43085
		), .Z(n_136997839));
	notech_nand2 i_3094209(.A(queue[8]), .B(n_58827), .Z(n_137097840));
	notech_nao3 i_1594224(.A(n_58711), .B(queue[88]), .C(n_58985), .Z(n_138597855
		));
	notech_nand3 i_924987(.A(n_269299158), .B(n_268599151), .C(n_137097840),
		 .Z(squeue[8]));
	notech_nand2 i_8794225(.A(queue[14]), .B(n_58822), .Z(n_138797857));
	notech_nao3 i_6494240(.A(n_58711), .B(queue[94]), .C(n_58985), .Z(n_140297872
		));
	notech_nand3 i_1524993(.A(n_270699172), .B(n_269999165), .C(n_138797857)
		, .Z(squeue[14]));
	notech_nand2 i_11894241(.A(n_58827), .B(queue[29]), .Z(n_140497874));
	notech_nao3 i_10394256(.A(n_58714), .B(queue[109]), .C(n_58985), .Z(n_141997889
		));
	notech_nand3 i_3025008(.A(n_272199186), .B(n_271499179), .C(n_140497874)
		, .Z(squeue[29]));
	notech_nand2 i_14994257(.A(n_58827), .B(queue[37]), .Z(n_142197891));
	notech_nao3 i_13494272(.A(n_58714), .B(queue[117]), .C(n_58985), .Z(n_143697906
		));
	notech_nand3 i_3825016(.A(n_273599200), .B(n_272899193), .C(n_142197891)
		, .Z(squeue[37]));
	notech_nand2 i_18094273(.A(n_58827), .B(queue[53]), .Z(n_143897908));
	notech_nao3 i_16594288(.A(n_58714), .B(queue[133]), .C(n_58982), .Z(n_145397923
		));
	notech_nand3 i_5425032(.A(n_275099214), .B(n_274299207), .C(n_143897908)
		, .Z(squeue[53]));
	notech_nand2 i_21194289(.A(n_58827), .B(queue[54]), .Z(n_145597925));
	notech_nao3 i_19694304(.A(n_58714), .B(queue[134]), .C(n_58982), .Z(n_147097940
		));
	notech_nand3 i_5525033(.A(n_276499228), .B(n_275799221), .C(n_145597925)
		, .Z(squeue[54]));
	notech_nand2 i_24294305(.A(n_58827), .B(queue[55]), .Z(n_147297942));
	notech_nao3 i_22794320(.A(n_58714), .B(queue[135]), .C(n_58982), .Z(n_148797957
		));
	notech_nand3 i_5625034(.A(n_277899242), .B(n_277199235), .C(n_147297942)
		, .Z(squeue[55]));
	notech_nand2 i_27394321(.A(n_58827), .B(queue[56]), .Z(n_148997959));
	notech_nao3 i_25894336(.A(n_58711), .B(queue[136]), .C(n_58982), .Z(n_150497974
		));
	notech_nand3 i_5725035(.A(n_279299256), .B(n_278599249), .C(n_148997959)
		, .Z(squeue[56]));
	notech_nand2 i_30494337(.A(n_58822), .B(queue[57]), .Z(n_150697976));
	notech_nao3 i_28994352(.A(n_58711), .B(queue[137]), .C(n_58982), .Z(n_152197991
		));
	notech_nand3 i_5825036(.A(n_280699270), .B(n_279999263), .C(n_150697976)
		, .Z(squeue[57]));
	notech_nand2 i_33594353(.A(n_58822), .B(queue[58]), .Z(n_152397993));
	notech_nao3 i_32094368(.A(n_58711), .B(queue[138]), .C(n_58982), .Z(n_153898008
		));
	notech_nand3 i_5925037(.A(n_282099284), .B(n_281399277), .C(n_152397993)
		, .Z(squeue[58]));
	notech_nand2 i_36694369(.A(n_58822), .B(queue[59]), .Z(n_154098010));
	notech_nao3 i_35194384(.A(n_58711), .B(queue[139]), .C(n_58982), .Z(n_155598025
		));
	notech_nand3 i_6025038(.A(n_283499298), .B(n_282799291), .C(n_154098010)
		, .Z(squeue[59]));
	notech_nand2 i_39794385(.A(n_58822), .B(queue[60]), .Z(n_155798027));
	notech_nao3 i_38294400(.A(n_58711), .B(queue[140]), .C(n_58982), .Z(n_157298042
		));
	notech_nand3 i_6125039(.A(n_284899312), .B(n_284199305), .C(n_155798027)
		, .Z(squeue[60]));
	notech_nand2 i_42894401(.A(n_58822), .B(queue[61]), .Z(n_157498044));
	notech_nao3 i_41394416(.A(n_58711), .B(queue[141]), .C(n_58982), .Z(n_158998059
		));
	notech_nand3 i_6225040(.A(n_286299326), .B(n_285599319), .C(n_157498044)
		, .Z(squeue[61]));
	notech_nand2 i_45994417(.A(n_58822), .B(queue[62]), .Z(n_159198061));
	notech_nao3 i_44494432(.A(n_58711), .B(queue[142]), .C(n_58982), .Z(n_160698076
		));
	notech_nand3 i_6325041(.A(n_287699340), .B(n_286999333), .C(n_159198061)
		, .Z(squeue[62]));
	notech_nand2 i_49094433(.A(n_58822), .B(queue[63]), .Z(n_160898078));
	notech_nao3 i_47594448(.A(n_58711), .B(queue[143]), .C(n_58985), .Z(n_162398093
		));
	notech_nand3 i_6425042(.A(n_289099354), .B(n_288399347), .C(n_160898078)
		, .Z(squeue[63]));
	notech_nand2 i_52194449(.A(n_58822), .B(queue[64]), .Z(n_162598095));
	notech_nao3 i_50694464(.A(n_58711), .B(queue[144]), .C(n_58987), .Z(n_164098110
		));
	notech_nand3 i_6525043(.A(n_290499368), .B(n_289799361), .C(n_162598095)
		, .Z(squeue[64]));
	notech_nand2 i_55294465(.A(n_58822), .B(queue[66]), .Z(n_164298112));
	notech_nao3 i_53794480(.A(n_58711), .B(queue[146]), .C(n_58987), .Z(n_165798127
		));
	notech_nand3 i_6725045(.A(n_291999382), .B(n_291299375), .C(n_164298112)
		, .Z(squeue[66]));
	notech_nand2 i_58394481(.A(n_58822), .B(queue[67]), .Z(n_165998129));
	notech_nao3 i_56894496(.A(n_58716), .B(queue[147]), .C(n_58987), .Z(n_167498144
		));
	notech_nand3 i_6825046(.A(n_293399396), .B(n_292699389), .C(n_165998129)
		, .Z(squeue[67]));
	notech_nand2 i_61494497(.A(n_58827), .B(queue[68]), .Z(n_167698146));
	notech_nao3 i_59994511(.A(n_58716), .B(queue[148]), .C(n_58987), .Z(n_169198161
		));
	notech_nand3 i_6925047(.A(n_294799410), .B(n_294099403), .C(n_167698146)
		, .Z(squeue[68]));
	notech_nand2 i_64594512(.A(n_58829), .B(queue[69]), .Z(n_169398163));
	notech_nao3 i_63094525(.A(n_58716), .B(queue[149]), .C(n_58987), .Z(n_170898178
		));
	notech_nand3 i_7025048(.A(n_296199424), .B(n_295499417), .C(n_169398163)
		, .Z(squeue[69]));
	notech_nand2 i_67694526(.A(n_58829), .B(queue[70]), .Z(n_171098180));
	notech_nao3 i_66194541(.A(n_58716), .B(queue[150]), .C(n_58987), .Z(n_172598195
		));
	notech_nand3 i_7125049(.A(n_297699438), .B(n_296999431), .C(n_171098180)
		, .Z(squeue[70]));
	notech_nand2 i_70794542(.A(n_58829), .B(queue[71]), .Z(n_172798197));
	notech_nao3 i_69294557(.A(n_58716), .B(queue[151]), .C(n_58987), .Z(n_174298212
		));
	notech_nand3 i_7225050(.A(n_299599452), .B(n_298499445), .C(n_172798197)
		, .Z(squeue[71]));
	notech_nand2 i_73894558(.A(n_58829), .B(queue[72]), .Z(n_174498214));
	notech_nao3 i_72394573(.A(n_58716), .B(queue[152]), .C(n_58987), .Z(n_175998229
		));
	notech_nand3 i_7325051(.A(n_3012), .B(n_300299455), .C(n_174498214), .Z(squeue
		[72]));
	notech_nand2 i_76994574(.A(n_58829), .B(queue[73]), .Z(n_176198231));
	notech_nao3 i_75494589(.A(n_58716), .B(queue[153]), .C(n_58987), .Z(n_177698246
		));
	notech_nand3 i_7425052(.A(n_302699460), .B(n_3019), .C(n_176198231), .Z(squeue
		[73]));
	notech_nand2 i_80094590(.A(n_58829), .B(queue[74]), .Z(n_177898248));
	notech_nao3 i_78594605(.A(n_58716), .B(queue[154]), .C(n_58987), .Z(n_179398263
		));
	notech_nand3 i_7525053(.A(n_3040), .B(n_3033), .C(n_177898248), .Z(squeue
		[74]));
	notech_nand2 i_83194606(.A(n_58829), .B(queue[75]), .Z(n_179598265));
	notech_nao3 i_81694621(.A(n_58716), .B(queue[155]), .C(n_58985), .Z(n_181098280
		));
	notech_nand3 i_7625054(.A(n_305699465), .B(n_3049), .C(n_179598265), .Z(squeue
		[75]));
	notech_nand2 i_86294622(.A(n_58829), .B(queue[76]), .Z(n_181298282));
	notech_nao3 i_84794637(.A(n_58716), .B(queue[156]), .C(n_58985), .Z(n_182798297
		));
	notech_nand3 i_7725055(.A(n_3070), .B(n_3063), .C(n_181298282), .Z(squeue
		[76]));
	notech_nand2 i_89394638(.A(n_58829), .B(queue[77]), .Z(n_182998299));
	notech_nao3 i_87894653(.A(n_58714), .B(queue[157]), .C(n_58985), .Z(n_184498314
		));
	notech_nand3 i_7825056(.A(n_3084), .B(n_3077), .C(n_182998299), .Z(squeue
		[77]));
	notech_nand2 i_92494654(.A(n_58829), .B(queue[78]), .Z(n_184698316));
	notech_nao3 i_90994669(.A(n_58714), .B(queue[158]), .C(n_58985), .Z(n_186198331
		));
	notech_nand3 i_7925057(.A(n_3100), .B(n_309299470), .C(n_184698316), .Z(squeue
		[78]));
	notech_nand2 i_95594670(.A(n_58827), .B(queue[79]), .Z(n_186398333));
	notech_nao3 i_94094685(.A(n_58714), .B(queue[159]), .C(n_58985), .Z(n_187898348
		));
	notech_nand3 i_8025058(.A(n_3114), .B(n_3107), .C(n_186398333), .Z(squeue
		[79]));
	notech_nand2 i_986(.A(n_58827), .B(queue[80]), .Z(n_188098350));
	notech_nao3 i_97194699(.A(n_58714), .B(queue[160]), .C(n_58987), .Z(n_189598365
		));
	notech_nand3 i_8125059(.A(n_312899475), .B(n_3121), .C(n_188098350), .Z(squeue
		[80]));
	notech_nand2 i_1017(.A(n_58827), .B(queue[81]), .Z(n_189798367));
	notech_nao3 i_1002(.A(n_58714), .B(queue[161]), .C(n_58987), .Z(n_191298382
		));
	notech_nand3 i_8225060(.A(n_3142), .B(n_3135), .C(n_189798367), .Z(squeue
		[81]));
	notech_nand2 i_1048(.A(n_58827), .B(queue[82]), .Z(n_191498384));
	notech_nao3 i_1033(.A(n_58716), .B(queue[162]), .C(n_58987), .Z(n_192998399
		));
	notech_nand3 i_8325061(.A(n_3156), .B(n_3149), .C(n_191498384), .Z(squeue
		[82]));
	notech_nand2 i_1079(.A(n_58827), .B(queue[83]), .Z(n_193198401));
	notech_nao3 i_1064(.A(n_58716), .B(queue[163]), .C(n_58985), .Z(n_194698416
		));
	notech_nand3 i_8425062(.A(n_317099482), .B(n_3163), .C(n_193198401), .Z(squeue
		[83]));
	notech_nand2 i_1110(.A(n_58829), .B(queue[84]), .Z(n_194898418));
	notech_nao3 i_1095(.A(n_58716), .B(queue[164]), .C(n_58987), .Z(n_196398433
		));
	notech_nand3 i_8525063(.A(n_3184), .B(n_3177), .C(n_194898418), .Z(squeue
		[84]));
	notech_nand2 i_1141(.A(n_58829), .B(queue[85]), .Z(n_196598435));
	notech_nao3 i_1126(.A(n_58714), .B(queue[165]), .C(n_58982), .Z(n_198098450
		));
	notech_nand3 i_8625064(.A(n_3198), .B(n_3191), .C(n_196598435), .Z(squeue
		[85]));
	notech_nand2 i_1172(.A(n_58829), .B(queue[86]), .Z(n_198298452));
	notech_nao3 i_1157(.A(n_58716), .B(queue[166]), .C(n_58975), .Z(n_199798467
		));
	notech_nand3 i_8725065(.A(n_321299489), .B(n_3205), .C(n_198298452), .Z(squeue
		[86]));
	notech_nand2 i_1203(.A(n_58829), .B(queue[87]), .Z(n_199998469));
	notech_nao3 i_1188(.A(n_58711), .B(queue[167]), .C(n_58975), .Z(n_201498484
		));
	notech_nand3 i_8825066(.A(n_3226), .B(n_3219), .C(n_199998469), .Z(squeue
		[87]));
	notech_nand2 i_1234(.A(n_58822), .B(queue[88]), .Z(n_201698486));
	notech_nao3 i_1219(.A(n_58705), .B(queue[168]), .C(n_58976), .Z(n_203198501
		));
	notech_nand3 i_8925067(.A(n_3240), .B(n_3233), .C(n_201698486), .Z(squeue
		[88]));
	notech_nand2 i_1265(.A(n_58829), .B(queue[89]), .Z(n_203398503));
	notech_nao3 i_1250(.A(n_58705), .B(queue[169]), .C(n_58976), .Z(n_204898518
		));
	notech_nand3 i_9025068(.A(n_325499496), .B(n_3247), .C(n_203398503), .Z(squeue
		[89]));
	notech_nand2 i_1296(.A(n_58829), .B(queue[90]), .Z(n_205098520));
	notech_nao3 i_1281(.A(n_58705), .B(queue[170]), .C(n_58976), .Z(n_206598535
		));
	notech_nand3 i_9125069(.A(n_3269), .B(n_3262), .C(n_205098520), .Z(squeue
		[90]));
	notech_nand2 i_1327(.A(n_58823), .B(queue[91]), .Z(n_206798537));
	notech_nao3 i_1312(.A(n_58705), .B(queue[171]), .C(n_58975), .Z(n_208298552
		));
	notech_nand3 i_9225070(.A(n_3283), .B(n_3276), .C(n_206798537), .Z(squeue
		[91]));
	notech_nand2 i_1358(.A(n_58823), .B(queue[92]), .Z(n_208498554));
	notech_nao3 i_1343(.A(n_58705), .B(queue[172]), .C(n_58975), .Z(n_209998569
		));
	notech_nand3 i_9325071(.A(n_3297), .B(n_329099501), .C(n_208498554), .Z(squeue
		[92]));
	notech_nand2 i_1389(.A(n_58829), .B(queue[93]), .Z(n_210198571));
	notech_nao3 i_1374(.A(n_58705), .B(queue[173]), .C(n_58975), .Z(n_211698586
		));
	notech_nand3 i_9425072(.A(n_3311), .B(n_3304), .C(n_210198571), .Z(squeue
		[93]));
	notech_nand2 i_1420(.A(n_58829), .B(queue[94]), .Z(n_211898588));
	notech_nao3 i_1405(.A(n_58705), .B(queue[174]), .C(n_58975), .Z(n_213398603
		));
	notech_nand3 i_9525073(.A(n_3325), .B(n_3318), .C(n_211898588), .Z(squeue
		[94]));
	notech_nand2 i_1451(.A(n_58827), .B(queue[95]), .Z(n_213598605));
	notech_nao3 i_1436(.A(n_58705), .B(queue[175]), .C(n_58975), .Z(n_215098620
		));
	notech_nand3 i_9625074(.A(n_3339), .B(n_333299508), .C(n_213598605), .Z(squeue
		[95]));
	notech_nand2 i_1482(.A(n_58829), .B(queue[96]), .Z(n_215298622));
	notech_nao3 i_1467(.A(n_58705), .B(queue[176]), .C(n_58975), .Z(n_216798637
		));
	notech_nand3 i_9725075(.A(n_3353), .B(n_3346), .C(n_215298622), .Z(squeue
		[96]));
	notech_nand2 i_1513(.A(n_58829), .B(queue[97]), .Z(n_216998639));
	notech_nao3 i_1498(.A(n_58705), .B(queue[177]), .C(n_58975), .Z(n_218498654
		));
	notech_nand3 i_9825076(.A(n_3367), .B(n_3360), .C(n_216998639), .Z(squeue
		[97]));
	notech_nand2 i_1544(.A(n_58823), .B(queue[98]), .Z(n_218698656));
	notech_nao3 i_1529(.A(n_58714), .B(queue[178]), .C(n_58975), .Z(n_220198671
		));
	notech_nand3 i_9925077(.A(n_3381), .B(n_337499515), .C(n_218698656), .Z(squeue
		[98]));
	notech_nand2 i_1575(.A(n_58823), .B(queue[99]), .Z(n_220398673));
	notech_nao3 i_1560(.A(n_58714), .B(queue[179]), .C(n_58975), .Z(n_221898688
		));
	notech_nand3 i_10025078(.A(n_3395), .B(n_3388), .C(n_220398673), .Z(squeue
		[99]));
	notech_nand2 i_1606(.A(n_58823), .B(queue[100]), .Z(n_222098690));
	notech_nao3 i_1591(.A(n_58714), .B(queue[180]), .C(n_58975), .Z(n_223598705
		));
	notech_nand3 i_10125079(.A(n_3409), .B(n_3402), .C(n_222098690), .Z(squeue
		[100]));
	notech_nand2 i_1637(.A(n_58823), .B(queue[101]), .Z(n_223798707));
	notech_nao3 i_1622(.A(n_58714), .B(queue[181]), .C(n_58976), .Z(n_225298722
		));
	notech_nand3 i_10225080(.A(n_3423), .B(n_341699522), .C(n_223798707), .Z
		(squeue[101]));
	notech_nand2 i_1668(.A(n_58823), .B(queue[102]), .Z(n_225498724));
	notech_nao3 i_1653(.A(n_58714), .B(queue[182]), .C(n_58976), .Z(n_226998739
		));
	notech_nand3 i_10325081(.A(n_3437), .B(n_3430), .C(n_225498724), .Z(squeue
		[102]));
	notech_nand2 i_1699(.A(n_58823), .B(queue[103]), .Z(n_227198741));
	notech_nao3 i_1684(.A(n_58705), .B(queue[183]), .C(n_58976), .Z(n_228698756
		));
	notech_nand3 i_10425082(.A(n_3451), .B(n_3444), .C(n_227198741), .Z(squeue
		[103]));
	notech_nand2 i_1730(.A(n_58823), .B(queue[104]), .Z(n_228898758));
	notech_nao3 i_1715(.A(n_58705), .B(queue[184]), .C(n_58975), .Z(n_230398773
		));
	notech_nand3 i_10525083(.A(n_3465), .B(n_345899529), .C(n_228898758), .Z
		(squeue[104]));
	notech_nand2 i_1761(.A(n_58823), .B(queue[105]), .Z(n_230598775));
	notech_nao3 i_1746(.A(n_58705), .B(queue[185]), .C(n_58976), .Z(n_232098790
		));
	notech_nand3 i_10625084(.A(n_3479), .B(n_3472), .C(n_230598775), .Z(squeue
		[105]));
	notech_nand2 i_1792(.A(n_58823), .B(queue[106]), .Z(n_232298792));
	notech_nao3 i_1777(.A(n_58714), .B(queue[186]), .C(n_58975), .Z(n_233798807
		));
	notech_nand3 i_10725085(.A(n_3493), .B(n_3486), .C(n_232298792), .Z(squeue
		[106]));
	notech_nand2 i_1823(.A(n_58823), .B(queue[107]), .Z(n_233998809));
	notech_nao3 i_1808(.A(n_58705), .B(queue[187]), .C(n_58980), .Z(n_235498824
		));
	notech_nand3 i_10825086(.A(n_3507), .B(n_350099536), .C(n_233998809), .Z
		(squeue[107]));
	notech_nand2 i_1854(.A(n_58827), .B(queue[108]), .Z(n_235698826));
	notech_nao3 i_1839(.A(n_58709), .B(queue[188]), .C(n_58980), .Z(n_237198841
		));
	notech_nand3 i_10925087(.A(n_3521), .B(n_3514), .C(n_235698826), .Z(squeue
		[108]));
	notech_nand2 i_1885(.A(n_58823), .B(queue[109]), .Z(n_237398843));
	notech_nao3 i_1870(.A(n_58709), .B(queue[189]), .C(n_58980), .Z(n_238898858
		));
	notech_nand3 i_11025088(.A(n_3535), .B(n_3528), .C(n_237398843), .Z(squeue
		[109]));
	notech_nand2 i_1916(.A(n_58823), .B(queue[110]), .Z(n_239098860));
	notech_nao3 i_1901(.A(n_58709), .B(queue[190]), .C(n_58980), .Z(n_240598875
		));
	notech_nand3 i_11125089(.A(n_3549), .B(n_354299543), .C(n_239098860), .Z
		(squeue[110]));
	notech_nand2 i_1947(.A(n_58823), .B(queue[111]), .Z(n_2407));
	notech_nao3 i_1932(.A(n_58709), .B(queue[191]), .C(n_58980), .Z(n_242398889
		));
	notech_nand3 i_11225090(.A(n_3563), .B(n_3556), .C(n_2407), .Z(squeue[
		111]));
	notech_nand2 i_1978(.A(n_58823), .B(queue[112]), .Z(n_242598891));
	notech_nao3 i_1963(.A(n_58709), .B(queue[192]), .C(n_58980), .Z(n_244098906
		));
	notech_nand3 i_11325091(.A(n_3577), .B(n_3570), .C(n_242598891), .Z(squeue
		[112]));
	notech_nand2 i_2009(.A(n_58823), .B(queue[113]), .Z(n_244298908));
	notech_nao3 i_1994(.A(n_58709), .B(queue[193]), .C(n_58980), .Z(n_245798923
		));
	notech_nand3 i_11425092(.A(n_3591), .B(n_358499550), .C(n_244298908), .Z
		(squeue[113]));
	notech_nand2 i_2040(.A(n_58822), .B(queue[114]), .Z(n_245998925));
	notech_nao3 i_2025(.A(n_58711), .B(queue[194]), .C(n_58980), .Z(n_247498940
		));
	notech_nand3 i_11525093(.A(n_3605), .B(n_3598), .C(n_245998925), .Z(squeue
		[114]));
	notech_nand2 i_2071(.A(n_58822), .B(queue[115]), .Z(n_247698942));
	notech_nao3 i_2056(.A(n_58709), .B(queue[195]), .C(n_58980), .Z(n_249198957
		));
	notech_nand3 i_11625094(.A(n_3619), .B(n_3612), .C(n_247698942), .Z(squeue
		[115]));
	notech_nand2 i_2102(.A(n_58823), .B(queue[116]), .Z(n_249398959));
	notech_nao3 i_2087(.A(n_58709), .B(queue[196]), .C(n_58980), .Z(n_250898974
		));
	notech_nand3 i_11725095(.A(n_3633), .B(n_362699557), .C(n_249398959), .Z
		(squeue[116]));
	notech_nand2 i_2133(.A(n_58823), .B(queue[117]), .Z(n_251098976));
	notech_nao3 i_2118(.A(n_58709), .B(queue[197]), .C(n_58975), .Z(n_252598991
		));
	notech_nand3 i_11825096(.A(n_3647), .B(n_3640), .C(n_251098976), .Z(squeue
		[117]));
	notech_nand2 i_2164(.A(n_58822), .B(queue[118]), .Z(n_252798993));
	notech_nao3 i_2149(.A(n_58705), .B(queue[198]), .C(n_58975), .Z(n_254299008
		));
	notech_nand3 i_11925097(.A(n_3661), .B(n_3654), .C(n_252798993), .Z(squeue
		[118]));
	notech_nand2 i_2195(.A(n_58827), .B(queue[119]), .Z(n_254499010));
	notech_nao3 i_2180(.A(n_58705), .B(queue[199]), .C(n_58975), .Z(n_255999025
		));
	notech_nand3 i_12025098(.A(n_3676), .B(n_366899564), .C(n_254499010), .Z
		(squeue[119]));
	notech_nand2 i_2226(.A(n_58827), .B(queue[120]), .Z(n_256199027));
	notech_nao3 i_2211(.A(n_58705), .B(queue[200]), .C(n_58975), .Z(n_257699042
		));
	notech_nand3 i_12125099(.A(n_3690), .B(n_3683), .C(n_256199027), .Z(squeue
		[120]));
	notech_nand2 i_2257(.A(n_58827), .B(queue[121]), .Z(n_257899044));
	notech_nao3 i_2242(.A(n_58705), .B(queue[201]), .C(n_58975), .Z(n_259399059
		));
	notech_nand3 i_12225100(.A(n_370499569), .B(n_3697), .C(n_257899044), .Z
		(squeue[121]));
	notech_nand2 i_2288(.A(n_58827), .B(queue[122]), .Z(n_259599061));
	notech_nao3 i_2273(.A(n_58705), .B(queue[202]), .C(n_58980), .Z(n_261099076
		));
	notech_nand3 i_12325101(.A(n_3718), .B(n_3711), .C(n_259599061), .Z(squeue
		[122]));
	notech_nand2 i_2319(.A(n_58822), .B(queue[123]), .Z(n_261299078));
	notech_nao3 i_2304(.A(n_58709), .B(queue[203]), .C(n_58980), .Z(n_262799093
		));
	notech_nand3 i_12425102(.A(n_3732), .B(n_3725), .C(n_261299078), .Z(squeue
		[123]));
	notech_nand2 i_2350(.A(n_58822), .B(queue[124]), .Z(n_262999095));
	notech_nao3 i_2335(.A(n_58709), .B(queue[204]), .C(n_58980), .Z(n_264499110
		));
	notech_nand3 i_12525103(.A(n_374699576), .B(n_3739), .C(n_262999095), .Z
		(squeue[124]));
	notech_nand2 i_2381(.A(n_58822), .B(queue[125]), .Z(n_264699112));
	notech_nao3 i_2366(.A(n_58709), .B(queue[205]), .C(n_58975), .Z(n_266199127
		));
	notech_nand3 i_12625104(.A(n_3760), .B(n_3753), .C(n_264699112), .Z(squeue
		[125]));
	notech_nand2 i_2412(.A(n_58822), .B(queue[126]), .Z(n_266399129));
	notech_nao3 i_2397(.A(n_58709), .B(queue[206]), .C(n_58980), .Z(n_267899144
		));
	notech_nand3 i_12725105(.A(n_3774), .B(n_3767), .C(n_266399129), .Z(squeue
		[126]));
	notech_ao4 i_3194700(.A(n_58640), .B(n_42963), .C(n_58756), .D(n_42955),
		 .Z(n_268099146));
	notech_ao4 i_3294702(.A(n_58777), .B(n_43027), .C(n_58614), .D(n_43019),
		 .Z(n_268299148));
	notech_ao4 i_3494703(.A(n_58735), .B(n_42971), .C(n_58445), .D(n_43035),
		 .Z(n_268399149));
	notech_and4 i_5994705(.A(n_268399149), .B(n_268299148), .C(n_268099146),
		 .D(n_138597855), .Z(n_268599151));
	notech_ao4 i_3594706(.A(n_58897), .B(n_42947), .C(n_58798), .D(n_43044),
		 .Z(n_268699152));
	notech_ao4 i_3694707(.A(n_58918), .B(n_42939), .C(n_58661), .D(n_42979),
		 .Z(n_268799153));
	notech_ao4 i_3794709(.A(n_58878), .B(n_42987), .C(n_58936), .D(n_42931),
		 .Z(n_268999155));
	notech_ao4 i_3894710(.A(n_58859), .B(n_42995), .C(n_58969), .D(n_43011),
		 .Z(n_269099156));
	notech_and4 i_6094712(.A(n_269099156), .B(n_268999155), .C(n_268799153),
		 .D(n_268699152), .Z(n_269299158));
	notech_ao4 i_8894714(.A(n_58640), .B(n_42969), .C(n_58756), .D(n_42961),
		 .Z(n_269499160));
	notech_ao4 i_8994716(.A(n_58777), .B(n_43033), .C(n_58614), .D(n_43025),
		 .Z(n_269699162));
	notech_ao4 i_9094717(.A(n_58735), .B(n_42977), .C(n_43041), .D(n_58441),
		 .Z(n_269799163));
	notech_and4 i_9994719(.A(n_269799163), .B(n_269699162), .C(n_269499160),
		 .D(n_140297872), .Z(n_269999165));
	notech_ao4 i_9194720(.A(n_58897), .B(n_42953), .C(n_58798), .D(n_43056),
		 .Z(n_270099166));
	notech_ao4 i_9294721(.A(n_58918), .B(n_42945), .C(n_58661), .D(n_42985),
		 .Z(n_270199167));
	notech_ao4 i_9394723(.A(n_58878), .B(n_42993), .C(n_58936), .D(n_42937),
		 .Z(n_270399169));
	notech_ao4 i_9494724(.A(n_58859), .B(n_43001), .C(n_58969), .D(n_43017),
		 .Z(n_270499170));
	notech_and4 i_10094726(.A(n_270499170), .B(n_270399169), .C(n_270199167)
		, .D(n_270099166), .Z(n_270699172));
	notech_ao4 i_11994728(.A(n_58640), .B(n_42984), .C(n_58756), .D(n_42976)
		, .Z(n_270899174));
	notech_ao4 i_12094730(.A(n_58777), .B(n_43054), .C(n_58614), .D(n_43040)
		, .Z(n_271099176));
	notech_ao4 i_12194731(.A(n_58735), .B(n_42992), .C(n_58445), .D(n_43070)
		, .Z(n_271199177));
	notech_and4 i_13094733(.A(n_271199177), .B(n_271099176), .C(n_270899174)
		, .D(n_141997889), .Z(n_271499179));
	notech_ao4 i_12294734(.A(n_58897), .B(n_42968), .C(n_58798), .D(n_43085)
		, .Z(n_271599180));
	notech_ao4 i_12394735(.A(n_58918), .B(n_42960), .C(n_58661), .D(n_43000)
		, .Z(n_271699181));
	notech_ao4 i_12494737(.A(n_58878), .B(n_43008), .C(n_58936), .D(n_42952)
		, .Z(n_271899183));
	notech_ao4 i_12594738(.A(n_58859), .B(n_43016), .C(n_58969), .D(n_43032)
		, .Z(n_271999184));
	notech_and4 i_13194740(.A(n_271999184), .B(n_271899183), .C(n_271699181)
		, .D(n_271599180), .Z(n_272199186));
	notech_ao4 i_15094742(.A(n_58640), .B(n_42992), .C(n_58756), .D(n_42984)
		, .Z(n_272399188));
	notech_ao4 i_15194744(.A(n_58777), .B(n_43070), .C(n_58614), .D(n_43054)
		, .Z(n_272599190));
	notech_ao4 i_15294745(.A(n_58735), .B(n_43000), .C(n_58445), .D(n_43085)
		, .Z(n_272699191));
	notech_and4 i_16194747(.A(n_272699191), .B(n_272599190), .C(n_272399188)
		, .D(n_143697906), .Z(n_272899193));
	notech_ao4 i_15394748(.A(n_58897), .B(n_42976), .C(n_58798), .D(n_43101)
		, .Z(n_272999194));
	notech_ao4 i_15494749(.A(n_58918), .B(n_42968), .C(n_58661), .D(n_43008)
		, .Z(n_273099195));
	notech_ao4 i_15594751(.A(n_58878), .B(n_43016), .C(n_58936), .D(n_42960)
		, .Z(n_273299197));
	notech_ao4 i_15694752(.A(n_58859), .B(n_43024), .C(n_58969), .D(n_43040)
		, .Z(n_273399198));
	notech_and4 i_16294754(.A(n_273399198), .B(n_273299197), .C(n_273099195)
		, .D(n_272999194), .Z(n_273599200));
	notech_ao4 i_18194756(.A(n_58640), .B(n_43008), .C(n_58756), .D(n_43000)
		, .Z(n_273799202));
	notech_ao4 i_18294758(.A(n_58777), .B(n_43101), .C(n_58614), .D(n_43085)
		, .Z(n_273999204));
	notech_ao4 i_18394759(.A(n_58735), .B(n_43016), .C(n_58445), .D(n_43117)
		, .Z(n_274099205));
	notech_and4 i_19294761(.A(n_274099205), .B(n_273999204), .C(n_273799202)
		, .D(n_145397923), .Z(n_274299207));
	notech_ao4 i_18494762(.A(n_58897), .B(n_42992), .C(n_58798), .D(n_43133)
		, .Z(n_274399208));
	notech_ao4 i_18594763(.A(n_58918), .B(n_42984), .C(n_58661), .D(n_43024)
		, .Z(n_274499209));
	notech_ao4 i_18694765(.A(n_58878), .B(n_43032), .C(n_58931), .D(n_42976)
		, .Z(n_274799211));
	notech_ao4 i_18794766(.A(n_58859), .B(n_43040), .C(n_58969), .D(n_43070)
		, .Z(n_274899212));
	notech_and4 i_19394768(.A(n_274899212), .B(n_274799211), .C(n_274499209)
		, .D(n_274399208), .Z(n_275099214));
	notech_ao4 i_21294770(.A(n_58640), .B(n_43009), .C(n_58756), .D(n_43001)
		, .Z(n_275299216));
	notech_ao4 i_21394772(.A(n_58777), .B(n_43103), .C(n_58614), .D(n_43087)
		, .Z(n_275499218));
	notech_ao4 i_21494773(.A(n_58735), .B(n_43017), .C(n_58445), .D(n_43119)
		, .Z(n_275599219));
	notech_and4 i_22394775(.A(n_275599219), .B(n_275499218), .C(n_275299216)
		, .D(n_147097940), .Z(n_275799221));
	notech_ao4 i_21594776(.A(n_58897), .B(n_42993), .C(n_58798), .D(n_43135)
		, .Z(n_275899222));
	notech_ao4 i_21694777(.A(n_58918), .B(n_42985), .C(n_58661), .D(n_43025)
		, .Z(n_275999223));
	notech_ao4 i_21794779(.A(n_58878), .B(n_43033), .C(n_58931), .D(n_42977)
		, .Z(n_276199225));
	notech_ao4 i_21894780(.A(n_58859), .B(n_43041), .C(n_58969), .D(n_43072)
		, .Z(n_276299226));
	notech_and4 i_22494782(.A(n_276299226), .B(n_276199225), .C(n_275999223)
		, .D(n_275899222), .Z(n_276499228));
	notech_ao4 i_24394784(.A(n_58640), .B(n_43010), .C(n_58756), .D(n_43002)
		, .Z(n_276699230));
	notech_ao4 i_24494786(.A(n_58777), .B(n_43105), .C(n_58618), .D(n_43089)
		, .Z(n_276899232));
	notech_ao4 i_24594787(.A(n_58735), .B(n_43018), .C(n_58445), .D(n_43121)
		, .Z(n_276999233));
	notech_and4 i_25494789(.A(n_276999233), .B(n_276899232), .C(n_276699230)
		, .D(n_148797957), .Z(n_277199235));
	notech_ao4 i_24694790(.A(n_58899), .B(n_42994), .C(n_58798), .D(n_43137)
		, .Z(n_277299236));
	notech_ao4 i_24794791(.A(n_58918), .B(n_42986), .C(n_58661), .D(n_43026)
		, .Z(n_277399237));
	notech_ao4 i_24894793(.A(n_58880), .B(n_43034), .C(n_58931), .D(n_42978)
		, .Z(n_277599239));
	notech_ao4 i_24994794(.A(n_58861), .B(n_43042), .C(n_58971), .D(n_43074)
		, .Z(n_277699240));
	notech_and4 i_25594796(.A(n_277699240), .B(n_277599239), .C(n_277399237)
		, .D(n_277299236), .Z(n_277899242));
	notech_ao4 i_27494798(.A(n_58640), .B(n_43011), .C(n_58756), .D(n_43003)
		, .Z(n_278099244));
	notech_ao4 i_27594800(.A(n_58777), .B(n_43107), .C(n_58618), .D(n_43091)
		, .Z(n_278299246));
	notech_ao4 i_27694801(.A(n_58735), .B(n_43019), .C(n_58445), .D(n_43123)
		, .Z(n_278399247));
	notech_and4 i_28594803(.A(n_278399247), .B(n_278299246), .C(n_278099244)
		, .D(n_150497974), .Z(n_278599249));
	notech_ao4 i_27794804(.A(n_58899), .B(n_42995), .C(n_58798), .D(n_43139)
		, .Z(n_278699250));
	notech_ao4 i_27894805(.A(n_58918), .B(n_42987), .C(n_58661), .D(n_43027)
		, .Z(n_278799251));
	notech_ao4 i_27994807(.A(n_58880), .B(n_43035), .C(n_58931), .D(n_42979)
		, .Z(n_278999253));
	notech_ao4 i_28094808(.A(n_58861), .B(n_43044), .C(n_58971), .D(n_43076)
		, .Z(n_279099254));
	notech_and4 i_28694810(.A(n_279099254), .B(n_278999253), .C(n_278799251)
		, .D(n_278699250), .Z(n_279299256));
	notech_ao4 i_30594812(.A(n_58640), .B(n_43012), .C(n_58756), .D(n_43004)
		, .Z(n_279499258));
	notech_ao4 i_30694814(.A(n_58777), .B(n_43109), .C(n_58618), .D(n_43093)
		, .Z(n_279699260));
	notech_ao4 i_30794815(.A(n_58735), .B(n_43020), .C(n_58441), .D(n_43125)
		, .Z(n_279799261));
	notech_and4 i_31694817(.A(n_279799261), .B(n_279699260), .C(n_279499258)
		, .D(n_152197991), .Z(n_279999263));
	notech_ao4 i_30894818(.A(n_58897), .B(n_42996), .C(n_58798), .D(n_43141)
		, .Z(n_280099264));
	notech_ao4 i_30994819(.A(n_58918), .B(n_42988), .C(n_58661), .D(n_43028)
		, .Z(n_280199265));
	notech_ao4 i_31094821(.A(n_58878), .B(n_43036), .C(n_58931), .D(n_42980)
		, .Z(n_280399267));
	notech_ao4 i_31194822(.A(n_58859), .B(n_43046), .C(n_58969), .D(n_43078)
		, .Z(n_280499268));
	notech_and4 i_31794824(.A(n_280499268), .B(n_280399267), .C(n_280199265)
		, .D(n_280099264), .Z(n_280699270));
	notech_ao4 i_33694826(.A(n_58640), .B(n_43013), .C(n_58756), .D(n_43005)
		, .Z(n_280899272));
	notech_ao4 i_33794828(.A(n_58777), .B(n_43111), .C(n_58618), .D(n_43095)
		, .Z(n_281099274));
	notech_ao4 i_33894829(.A(n_58735), .B(n_43021), .C(n_58441), .D(n_43127)
		, .Z(n_281199275));
	notech_and4 i_34794831(.A(n_281199275), .B(n_281099274), .C(n_280899272)
		, .D(n_153898008), .Z(n_281399277));
	notech_ao4 i_33994832(.A(n_58897), .B(n_42997), .C(n_58798), .D(n_43143)
		, .Z(n_281499278));
	notech_ao4 i_34094833(.A(n_58918), .B(n_42989), .C(n_58661), .D(n_43029)
		, .Z(n_281599279));
	notech_ao4 i_34194835(.A(n_58878), .B(n_43037), .C(n_58931), .D(n_42981)
		, .Z(n_281799281));
	notech_ao4 i_34294836(.A(n_58859), .B(n_43048), .C(n_58969), .D(n_43080)
		, .Z(n_281899282));
	notech_and4 i_34894838(.A(n_281899282), .B(n_281799281), .C(n_281599279)
		, .D(n_281499278), .Z(n_282099284));
	notech_ao4 i_36794840(.A(n_58640), .B(n_43014), .C(n_58756), .D(n_43006)
		, .Z(n_282299286));
	notech_ao4 i_36894842(.A(n_58777), .B(n_43113), .C(n_58614), .D(n_43097)
		, .Z(n_282499288));
	notech_ao4 i_36994843(.A(n_58735), .B(n_43022), .C(n_58441), .D(n_43129)
		, .Z(n_282599289));
	notech_and4 i_37894845(.A(n_282599289), .B(n_282499288), .C(n_282299286)
		, .D(n_155598025), .Z(n_282799291));
	notech_ao4 i_37094846(.A(n_58897), .B(n_42998), .C(n_58798), .D(n_43144)
		, .Z(n_282899292));
	notech_ao4 i_37194847(.A(n_58918), .B(n_42990), .C(n_58661), .D(n_43030)
		, .Z(n_282999293));
	notech_ao4 i_37294849(.A(n_58878), .B(n_43038), .C(n_58936), .D(n_42982)
		, .Z(n_283199295));
	notech_ao4 i_37394850(.A(n_58859), .B(n_43050), .C(n_58969), .D(n_43082)
		, .Z(n_283299296));
	notech_and4 i_37994852(.A(n_283299296), .B(n_283199295), .C(n_282999293)
		, .D(n_282899292), .Z(n_283499298));
	notech_ao4 i_39894854(.A(n_58640), .B(n_43015), .C(n_58756), .D(n_43007)
		, .Z(n_283699300));
	notech_ao4 i_39994856(.A(n_58777), .B(n_43115), .C(n_58614), .D(n_43099)
		, .Z(n_283899302));
	notech_ao4 i_40094857(.A(n_58735), .B(n_43023), .C(n_58441), .D(n_43131)
		, .Z(n_283999303));
	notech_and4 i_40994859(.A(n_283999303), .B(n_283899302), .C(n_283699300)
		, .D(n_157298042), .Z(n_284199305));
	notech_ao4 i_40194860(.A(n_58897), .B(n_42999), .C(n_58798), .D(n_43146)
		, .Z(n_284299306));
	notech_ao4 i_40294861(.A(n_58918), .B(n_42991), .C(n_58661), .D(n_43031)
		, .Z(n_284399307));
	notech_ao4 i_40394863(.A(n_58878), .B(n_43039), .C(n_58936), .D(n_42983)
		, .Z(n_284599309));
	notech_ao4 i_40494864(.A(n_58859), .B(n_43052), .C(n_58969), .D(n_43084)
		, .Z(n_284699310));
	notech_and4 i_41094866(.A(n_284699310), .B(n_284599309), .C(n_284399307)
		, .D(n_284299306), .Z(n_284899312));
	notech_ao4 i_42994868(.A(n_58640), .B(n_43016), .C(n_58756), .D(n_43008)
		, .Z(n_285099314));
	notech_ao4 i_43094870(.A(n_58777), .B(n_43117), .C(n_58614), .D(n_43101)
		, .Z(n_285299316));
	notech_ao4 i_43194871(.A(n_58735), .B(n_43024), .C(n_58441), .D(n_43133)
		, .Z(n_285399317));
	notech_and4 i_44094873(.A(n_285399317), .B(n_285299316), .C(n_285099314)
		, .D(n_158998059), .Z(n_285599319));
	notech_ao4 i_43294874(.A(n_58892), .B(n_43000), .C(n_58798), .D(n_43148)
		, .Z(n_285699320));
	notech_ao4 i_43394875(.A(n_58918), .B(n_42992), .C(n_58661), .D(n_43032)
		, .Z(n_285799321));
	notech_ao4 i_43494877(.A(n_58873), .B(n_43040), .C(n_58936), .D(n_42984)
		, .Z(n_285999323));
	notech_ao4 i_43594878(.A(n_58854), .B(n_43054), .C(n_58964), .D(n_43085)
		, .Z(n_286099324));
	notech_and4 i_44194880(.A(n_286099324), .B(n_285999323), .C(n_285799321)
		, .D(n_285699320), .Z(n_286299326));
	notech_ao4 i_46094882(.A(n_58627), .B(n_43017), .C(n_58743), .D(n_43009)
		, .Z(n_286499328));
	notech_ao4 i_46194884(.A(n_58764), .B(n_43119), .C(n_58621), .D(n_43103)
		, .Z(n_286699330));
	notech_ao4 i_46294885(.A(n_58722), .B(n_43025), .C(n_58441), .D(n_43135)
		, .Z(n_286799331));
	notech_and4 i_47194887(.A(n_286799331), .B(n_286699330), .C(n_286499328)
		, .D(n_160698076), .Z(n_286999333));
	notech_ao4 i_46394888(.A(n_58885), .B(n_43001), .C(n_58785), .D(n_43150)
		, .Z(n_287099334));
	notech_ao4 i_46494889(.A(n_58905), .B(n_42993), .C(n_58648), .D(n_43033)
		, .Z(n_287199335));
	notech_ao4 i_46594891(.A(n_58866), .B(n_43041), .C(n_58931), .D(n_42985)
		, .Z(n_287399337));
	notech_ao4 i_46694892(.A(n_58847), .B(n_43056), .C(n_58957), .D(n_43087)
		, .Z(n_287499338));
	notech_and4 i_47294894(.A(n_287499338), .B(n_287399337), .C(n_287199335)
		, .D(n_287099334), .Z(n_287699340));
	notech_ao4 i_49194896(.A(n_58627), .B(n_43018), .C(n_58743), .D(n_43010)
		, .Z(n_287899342));
	notech_ao4 i_49294898(.A(n_58764), .B(n_43121), .C(n_58621), .D(n_43105)
		, .Z(n_288099344));
	notech_ao4 i_49394899(.A(n_58722), .B(n_43026), .C(n_58441), .D(n_43137)
		, .Z(n_288199345));
	notech_and4 i_50294901(.A(n_288199345), .B(n_288099344), .C(n_287899342)
		, .D(n_162398093), .Z(n_288399347));
	notech_ao4 i_49494902(.A(n_58885), .B(n_43002), .C(n_58785), .D(n_43152)
		, .Z(n_288499348));
	notech_ao4 i_49594903(.A(n_58905), .B(n_42994), .C(n_58648), .D(n_43034)
		, .Z(n_288599349));
	notech_ao4 i_49694905(.A(n_58866), .B(n_43042), .C(n_58931), .D(n_42986)
		, .Z(n_288799351));
	notech_ao4 i_49794906(.A(n_58847), .B(n_43058), .C(n_58957), .D(n_43089)
		, .Z(n_288899352));
	notech_and4 i_50394908(.A(n_288899352), .B(n_288799351), .C(n_288599349)
		, .D(n_288499348), .Z(n_289099354));
	notech_ao4 i_52294910(.A(n_58627), .B(n_43019), .C(n_58743), .D(n_43011)
		, .Z(n_289299356));
	notech_ao4 i_52394912(.A(n_58764), .B(n_43123), .C(n_58621), .D(n_43107)
		, .Z(n_289499358));
	notech_ao4 i_52494913(.A(n_58722), .B(n_43027), .C(n_58441), .D(n_43139)
		, .Z(n_289599359));
	notech_and4 i_53394915(.A(n_289599359), .B(n_289499358), .C(n_289299356)
		, .D(n_164098110), .Z(n_289799361));
	notech_ao4 i_52594916(.A(n_58885), .B(n_43003), .C(n_58785), .D(n_43154)
		, .Z(n_289899362));
	notech_ao4 i_52694917(.A(n_58905), .B(n_42995), .C(n_58648), .D(n_43035)
		, .Z(n_289999363));
	notech_ao4 i_52794919(.A(n_58866), .B(n_43044), .C(n_58938), .D(n_42987)
		, .Z(n_290199365));
	notech_ao4 i_52894920(.A(n_58847), .B(n_43060), .C(n_58957), .D(n_43091)
		, .Z(n_290299366));
	notech_and4 i_53494922(.A(n_290299366), .B(n_290199365), .C(n_289999363)
		, .D(n_289899362), .Z(n_290499368));
	notech_ao4 i_55394924(.A(n_58627), .B(n_43021), .C(n_58743), .D(n_43013)
		, .Z(n_290799370));
	notech_ao4 i_55494926(.A(n_58764), .B(n_43127), .C(n_58621), .D(n_43111)
		, .Z(n_290999372));
	notech_ao4 i_55594927(.A(n_58722), .B(n_43029), .C(n_58441), .D(n_43143)
		, .Z(n_291099373));
	notech_and4 i_56494929(.A(n_291099373), .B(n_290999372), .C(n_290799370)
		, .D(n_165798127), .Z(n_291299375));
	notech_ao4 i_55694930(.A(n_58885), .B(n_43005), .C(n_58785), .D(n_43158)
		, .Z(n_291399376));
	notech_ao4 i_55794931(.A(n_58905), .B(n_42997), .C(n_58648), .D(n_43037)
		, .Z(n_291499377));
	notech_ao4 i_55894933(.A(n_58866), .B(n_43048), .C(n_58938), .D(n_42989)
		, .Z(n_291699379));
	notech_ao4 i_55994934(.A(n_58847), .B(n_43064), .C(n_58957), .D(n_43095)
		, .Z(n_291799380));
	notech_and4 i_56594936(.A(n_291799380), .B(n_291699379), .C(n_291499377)
		, .D(n_291399376), .Z(n_291999382));
	notech_ao4 i_58494938(.A(n_58627), .B(n_43022), .C(n_58743), .D(n_43014)
		, .Z(n_292199384));
	notech_ao4 i_58594940(.A(n_58764), .B(n_43129), .C(n_58621), .D(n_43113)
		, .Z(n_292399386));
	notech_ao4 i_58694941(.A(n_58722), .B(n_43030), .C(n_58441), .D(n_43144)
		, .Z(n_292499387));
	notech_and4 i_59594943(.A(n_292499387), .B(n_292399386), .C(n_292199384)
		, .D(n_167498144), .Z(n_292699389));
	notech_ao4 i_58794944(.A(n_58885), .B(n_43006), .C(n_58785), .D(n_43160)
		, .Z(n_292799390));
	notech_ao4 i_58894945(.A(n_58905), .B(n_42998), .C(n_58648), .D(n_43038)
		, .Z(n_292899391));
	notech_ao4 i_58994947(.A(n_58866), .B(n_43050), .C(n_58938), .D(n_42990)
		, .Z(n_293099393));
	notech_ao4 i_59094948(.A(n_58847), .B(n_43066), .C(n_58957), .D(n_43097)
		, .Z(n_293199394));
	notech_and4 i_59694950(.A(n_293199394), .B(n_293099393), .C(n_292899391)
		, .D(n_292799390), .Z(n_293399396));
	notech_ao4 i_61594952(.A(n_58627), .B(n_43023), .C(n_58743), .D(n_43015)
		, .Z(n_293599398));
	notech_ao4 i_61694954(.A(n_58764), .B(n_43131), .C(n_58621), .D(n_43115)
		, .Z(n_293799400));
	notech_ao4 i_61794955(.A(n_58722), .B(n_43031), .C(n_58445), .D(n_43146)
		, .Z(n_293899401));
	notech_and4 i_62680080(.A(n_293899401), .B(n_293799400), .C(n_293599398)
		, .D(n_169198161), .Z(n_294099403));
	notech_ao4 i_61894957(.A(n_58885), .B(n_43007), .C(n_58785), .D(n_43162)
		, .Z(n_294199404));
	notech_ao4 i_61994958(.A(n_58905), .B(n_42999), .C(n_58648), .D(n_43039)
		, .Z(n_294299405));
	notech_ao4 i_62094960(.A(n_58866), .B(n_43052), .C(n_58938), .D(n_42991)
		, .Z(n_294499407));
	notech_ao4 i_62194961(.A(n_58847), .B(n_43068), .C(n_58957), .D(n_43099)
		, .Z(n_294599408));
	notech_and4 i_62794963(.A(n_294599408), .B(n_294499407), .C(n_294299405)
		, .D(n_294199404), .Z(n_294799410));
	notech_ao4 i_64694965(.A(n_58627), .B(n_43024), .C(n_58743), .D(n_43016)
		, .Z(n_294999412));
	notech_ao4 i_64794967(.A(n_58764), .B(n_43133), .C(n_58621), .D(n_43117)
		, .Z(n_295199414));
	notech_ao4 i_64894968(.A(n_58722), .B(n_43032), .C(n_58447), .D(n_43148)
		, .Z(n_295299415));
	notech_and4 i_65794970(.A(n_295299415), .B(n_295199414), .C(n_294999412)
		, .D(n_170898178), .Z(n_295499417));
	notech_ao4 i_64994971(.A(n_58885), .B(n_43008), .C(n_58785), .D(n_43164)
		, .Z(n_295599418));
	notech_ao4 i_65094972(.A(n_58905), .B(n_43000), .C(n_58648), .D(n_43040)
		, .Z(n_295699419));
	notech_ao4 i_65194974(.A(n_58866), .B(n_43054), .C(n_58938), .D(n_42992)
		, .Z(n_295899421));
	notech_ao4 i_65294975(.A(n_58847), .B(n_43070), .C(n_58957), .D(n_43101)
		, .Z(n_295999422));
	notech_and4 i_65894976(.A(n_295999422), .B(n_295899421), .C(n_295699419)
		, .D(n_295599418), .Z(n_296199424));
	notech_ao4 i_67794978(.A(n_58627), .B(n_43025), .C(n_58743), .D(n_43017)
		, .Z(n_296399426));
	notech_ao4 i_67894980(.A(n_58764), .B(n_43135), .C(n_58621), .D(n_43119)
		, .Z(n_296699428));
	notech_ao4 i_67994981(.A(n_58722), .B(n_43033), .C(n_58447), .D(n_43150)
		, .Z(n_296799429));
	notech_and4 i_68894983(.A(n_296799429), .B(n_296699428), .C(n_296399426)
		, .D(n_172598195), .Z(n_296999431));
	notech_ao4 i_68094984(.A(n_58885), .B(n_43009), .C(n_58785), .D(n_43166)
		, .Z(n_297099432));
	notech_ao4 i_68194985(.A(n_58905), .B(n_43001), .C(n_58648), .D(n_43041)
		, .Z(n_297199433));
	notech_ao4 i_68294987(.A(n_58866), .B(n_43056), .C(n_58938), .D(n_42993)
		, .Z(n_297399435));
	notech_ao4 i_68394988(.A(n_58847), .B(n_43072), .C(n_58957), .D(n_43103)
		, .Z(n_297499436));
	notech_and4 i_68994990(.A(n_297499436), .B(n_297399435), .C(n_297199433)
		, .D(n_297099432), .Z(n_297699438));
	notech_ao4 i_70894992(.A(n_58627), .B(n_43026), .C(n_58743), .D(n_43018)
		, .Z(n_297899440));
	notech_ao4 i_70994994(.A(n_58764), .B(n_43137), .C(n_58621), .D(n_43121)
		, .Z(n_298099442));
	notech_ao4 i_71094995(.A(n_58722), .B(n_43034), .C(n_58447), .D(n_43152)
		, .Z(n_298199443));
	notech_and4 i_71994997(.A(n_298199443), .B(n_298099442), .C(n_297899440)
		, .D(n_174298212), .Z(n_298499445));
	notech_ao4 i_71194998(.A(n_58887), .B(n_43010), .C(n_58785), .D(n_43168)
		, .Z(n_298699446));
	notech_ao4 i_71294999(.A(n_58905), .B(n_43002), .C(n_58648), .D(n_43042)
		, .Z(n_298899447));
	notech_ao4 i_71395001(.A(n_58868), .B(n_43058), .C(n_58938), .D(n_42994)
		, .Z(n_299099449));
	notech_ao4 i_71495002(.A(n_58849), .B(n_43074), .C(n_58959), .D(n_43105)
		, .Z(n_299299450));
	notech_and4 i_72095004(.A(n_299299450), .B(n_299099449), .C(n_298899447)
		, .D(n_298699446), .Z(n_299599452));
	notech_ao4 i_73995006(.A(n_58627), .B(n_43027), .C(n_58743), .D(n_43019)
		, .Z(n_299799454));
	notech_ao4 i_74095008(.A(n_58764), .B(n_43139), .C(n_58621), .D(n_43123)
		, .Z(n_2999));
	notech_ao4 i_74195009(.A(n_58722), .B(n_43035), .C(n_58447), .D(n_43154)
		, .Z(n_3000));
	notech_and4 i_75095011(.A(n_3000), .B(n_2999), .C(n_299799454), .D(n_175998229
		), .Z(n_300299455));
	notech_ao4 i_74295012(.A(n_58887), .B(n_43011), .C(n_58785), .D(n_43170)
		, .Z(n_3004));
	notech_ao4 i_74395013(.A(n_58905), .B(n_43003), .C(n_58648), .D(n_43044)
		, .Z(n_3005));
	notech_ao4 i_74495015(.A(n_58868), .B(n_43060), .C(n_58938), .D(n_42995)
		, .Z(n_3009));
	notech_ao4 i_74595016(.A(n_58849), .B(n_43076), .C(n_58959), .D(n_43107)
		, .Z(n_3010));
	notech_and4 i_75195018(.A(n_3010), .B(n_3009), .C(n_3005), .D(n_3004), .Z
		(n_3012));
	notech_ao4 i_77095020(.A(n_58627), .B(n_43028), .C(n_58743), .D(n_43020)
		, .Z(n_301499456));
	notech_ao4 i_77195022(.A(n_58764), .B(n_43141), .C(n_58621), .D(n_43125)
		, .Z(n_301699457));
	notech_ao4 i_77295023(.A(n_58722), .B(n_43036), .C(n_58447), .D(n_43156)
		, .Z(n_3017));
	notech_and4 i_78195025(.A(n_3017), .B(n_301699457), .C(n_301499456), .D(n_177698246
		), .Z(n_3019));
	notech_ao4 i_77395026(.A(n_58887), .B(n_43012), .C(n_58785), .D(n_43172)
		, .Z(n_302099459));
	notech_ao4 i_77495027(.A(n_58905), .B(n_43004), .C(n_58648), .D(n_43046)
		, .Z(n_3021));
	notech_ao4 i_77595029(.A(n_58868), .B(n_43062), .C(n_58938), .D(n_42996)
		, .Z(n_3023));
	notech_ao4 i_77695030(.A(n_58849), .B(n_43078), .C(n_58959), .D(n_43109)
		, .Z(n_3024));
	notech_and4 i_78295032(.A(n_3024), .B(n_3023), .C(n_3021), .D(n_302099459
		), .Z(n_302699460));
	notech_ao4 i_80195034(.A(n_58627), .B(n_43029), .C(n_58743), .D(n_43021)
		, .Z(n_3028));
	notech_ao4 i_80295036(.A(n_58764), .B(n_43143), .C(n_58621), .D(n_43127)
		, .Z(n_3030));
	notech_ao4 i_80395037(.A(n_58722), .B(n_43037), .C(n_58447), .D(n_43158)
		, .Z(n_3031));
	notech_and4 i_81295039(.A(n_3031), .B(n_3030), .C(n_3028), .D(n_179398263
		), .Z(n_3033));
	notech_ao4 i_80495040(.A(n_58887), .B(n_43013), .C(n_58785), .D(n_43174)
		, .Z(n_3034));
	notech_ao4 i_80595041(.A(n_58905), .B(n_43005), .C(n_58648), .D(n_43048)
		, .Z(n_3035));
	notech_ao4 i_80695043(.A(n_58868), .B(n_43064), .C(n_58938), .D(n_42997)
		, .Z(n_3037));
	notech_ao4 i_80795044(.A(n_58849), .B(n_43080), .C(n_58959), .D(n_43111)
		, .Z(n_303899462));
	notech_and4 i_81395046(.A(n_303899462), .B(n_3037), .C(n_3035), .D(n_3034
		), .Z(n_3040));
	notech_ao4 i_83295048(.A(n_58627), .B(n_43030), .C(n_58743), .D(n_43022)
		, .Z(n_3042));
	notech_ao4 i_83395050(.A(n_58764), .B(n_43144), .C(n_58621), .D(n_43129)
		, .Z(n_304499463));
	notech_ao4 i_83495051(.A(n_58722), .B(n_43038), .C(n_58447), .D(n_43160)
		, .Z(n_3045));
	notech_and4 i_84395053(.A(n_3045), .B(n_304499463), .C(n_3042), .D(n_181098280
		), .Z(n_3049));
	notech_ao4 i_83595054(.A(n_58887), .B(n_43014), .C(n_58785), .D(n_43176)
		, .Z(n_305099464));
	notech_ao4 i_83695055(.A(n_58905), .B(n_43006), .C(n_58648), .D(n_43050)
		, .Z(n_3051));
	notech_ao4 i_83795057(.A(n_58868), .B(n_43066), .C(n_58938), .D(n_42998)
		, .Z(n_3053));
	notech_ao4 i_83895058(.A(n_58849), .B(n_43082), .C(n_58959), .D(n_43113)
		, .Z(n_3054));
	notech_and4 i_84495060(.A(n_3054), .B(n_3053), .C(n_3051), .D(n_305099464
		), .Z(n_305699465));
	notech_ao4 i_86395062(.A(n_58627), .B(n_43031), .C(n_58743), .D(n_43023)
		, .Z(n_3058));
	notech_ao4 i_86495064(.A(n_58764), .B(n_43146), .C(n_58621), .D(n_43131)
		, .Z(n_3060));
	notech_ao4 i_86595065(.A(n_58722), .B(n_43039), .C(n_58447), .D(n_43162)
		, .Z(n_3061));
	notech_and4 i_87495067(.A(n_3061), .B(n_3060), .C(n_3058), .D(n_182798297
		), .Z(n_3063));
	notech_ao4 i_86695068(.A(n_58887), .B(n_43015), .C(n_58785), .D(n_43178)
		, .Z(n_3064));
	notech_ao4 i_86795069(.A(n_58905), .B(n_43007), .C(n_58648), .D(n_43052)
		, .Z(n_3065));
	notech_ao4 i_86895071(.A(n_58868), .B(n_43068), .C(n_58936), .D(n_42999)
		, .Z(n_3067));
	notech_ao4 i_86995072(.A(n_58849), .B(n_43084), .C(n_58957), .D(n_43115)
		, .Z(n_306899467));
	notech_and4 i_87595074(.A(n_306899467), .B(n_3067), .C(n_3065), .D(n_3064
		), .Z(n_3070));
	notech_ao4 i_89495076(.A(n_58627), .B(n_43032), .C(n_58743), .D(n_43024)
		, .Z(n_3072));
	notech_ao4 i_89595078(.A(n_58764), .B(n_43148), .C(n_58621), .D(n_43133)
		, .Z(n_307499468));
	notech_ao4 i_89695079(.A(n_58722), .B(n_43040), .C(n_58447), .D(n_43164)
		, .Z(n_3075));
	notech_and4 i_90595081(.A(n_3075), .B(n_307499468), .C(n_3072), .D(n_184498314
		), .Z(n_3077));
	notech_ao4 i_89795082(.A(n_58887), .B(n_43016), .C(n_58785), .D(n_43180)
		, .Z(n_3078));
	notech_ao4 i_89895083(.A(n_58905), .B(n_43008), .C(n_58648), .D(n_43054)
		, .Z(n_3079));
	notech_ao4 i_89995085(.A(n_58868), .B(n_43070), .C(n_58938), .D(n_43000)
		, .Z(n_3081));
	notech_ao4 i_90095086(.A(n_58849), .B(n_43085), .C(n_58959), .D(n_43117)
		, .Z(n_3082));
	notech_and4 i_90695088(.A(n_3082), .B(n_3081), .C(n_3079), .D(n_3078), .Z
		(n_3084));
	notech_ao4 i_92595090(.A(n_58627), .B(n_43033), .C(n_58743), .D(n_43025)
		, .Z(n_3087));
	notech_ao4 i_92695092(.A(n_58764), .B(n_43150), .C(n_58619), .D(n_43135)
		, .Z(n_3089));
	notech_ao4 i_92795093(.A(n_58722), .B(n_43041), .C(n_58447), .D(n_43166)
		, .Z(n_3090));
	notech_and4 i_93695095(.A(n_3090), .B(n_3089), .C(n_3087), .D(n_186198331
		), .Z(n_309299470));
	notech_ao4 i_92895096(.A(n_58887), .B(n_43017), .C(n_58785), .D(n_43182)
		, .Z(n_3093));
	notech_ao4 i_92995097(.A(n_58905), .B(n_43009), .C(n_58648), .D(n_43056)
		, .Z(n_3094));
	notech_ao4 i_93095099(.A(n_58868), .B(n_43072), .C(n_58936), .D(n_43001)
		, .Z(n_3096));
	notech_ao4 i_93195100(.A(n_58849), .B(n_43087), .C(n_58959), .D(n_43119)
		, .Z(n_3097));
	notech_and4 i_93795102(.A(n_3097), .B(n_3096), .C(n_3094), .D(n_3093), .Z
		(n_3100));
	notech_ao4 i_95695104(.A(n_58625), .B(n_43034), .C(n_58741), .D(n_43026)
		, .Z(n_3102));
	notech_ao4 i_95795106(.A(n_58762), .B(n_43152), .C(n_58619), .D(n_43137)
		, .Z(n_310499471));
	notech_ao4 i_95895107(.A(n_58720), .B(n_43042), .C(n_58445), .D(n_43168)
		, .Z(n_3105));
	notech_and4 i_96795109(.A(n_3105), .B(n_310499471), .C(n_3102), .D(n_187898348
		), .Z(n_3107));
	notech_ao4 i_95995110(.A(n_58884), .B(n_43018), .C(n_58783), .D(n_43184)
		, .Z(n_3108));
	notech_ao4 i_96095111(.A(n_58903), .B(n_43010), .C(n_58646), .D(n_43058)
		, .Z(n_3109));
	notech_ao4 i_96195113(.A(n_58865), .B(n_43074), .C(n_58936), .D(n_43002)
		, .Z(n_3111));
	notech_ao4 i_96295114(.A(n_58846), .B(n_43089), .C(n_58956), .D(n_43121)
		, .Z(n_3112));
	notech_and4 i_96895116(.A(n_3112), .B(n_3111), .C(n_3109), .D(n_3108), .Z
		(n_3114));
	notech_ao4 i_987(.A(n_58625), .B(n_43035), .C(n_58741), .D(n_43027), .Z(n_311699473
		));
	notech_ao4 i_988(.A(n_58762), .B(n_43154), .C(n_58619), .D(n_43139), .Z(n_3118
		));
	notech_ao4 i_989(.A(n_58720), .B(n_43044), .C(n_58445), .D(n_43170), .Z(n_3119
		));
	notech_and4 i_998(.A(n_3119), .B(n_3118), .C(n_311699473), .D(n_189598365
		), .Z(n_3121));
	notech_ao4 i_990(.A(n_58884), .B(n_43019), .C(n_58783), .D(n_43186), .Z(n_312299474
		));
	notech_ao4 i_991(.A(n_58903), .B(n_43011), .C(n_58646), .D(n_43060), .Z(n_3123
		));
	notech_ao4 i_992(.A(n_58865), .B(n_43076), .C(n_58936), .D(n_43003), .Z(n_3125
		));
	notech_ao4 i_993(.A(n_58846), .B(n_43091), .C(n_58956), .D(n_43123), .Z(n_3126
		));
	notech_and4 i_999(.A(n_3126), .B(n_3125), .C(n_3123), .D(n_312299474), .Z
		(n_312899475));
	notech_ao4 i_1018(.A(n_58625), .B(n_43036), .C(n_58741), .D(n_43028), .Z
		(n_3130));
	notech_ao4 i_1019(.A(n_58762), .B(n_43156), .C(n_58619), .D(n_43141), .Z
		(n_3132));
	notech_ao4 i_1020(.A(n_58720), .B(n_43046), .C(n_58445), .D(n_43172), .Z
		(n_3133));
	notech_and4 i_1029(.A(n_3133), .B(n_3132), .C(n_3130), .D(n_191298382), 
		.Z(n_3135));
	notech_ao4 i_1021(.A(n_58884), .B(n_43020), .C(n_58783), .D(n_43188), .Z
		(n_3136));
	notech_ao4 i_1022(.A(n_58903), .B(n_43012), .C(n_58646), .D(n_43062), .Z
		(n_3137));
	notech_ao4 i_1023(.A(n_58865), .B(n_43078), .C(n_58938), .D(n_43004), .Z
		(n_3139));
	notech_ao4 i_1024(.A(n_58846), .B(n_43093), .C(n_58956), .D(n_43125), .Z
		(n_314099477));
	notech_and4 i_1030(.A(n_314099477), .B(n_3139), .C(n_3137), .D(n_3136), 
		.Z(n_3142));
	notech_ao4 i_1049(.A(n_58625), .B(n_43037), .C(n_58741), .D(n_43029), .Z
		(n_3144));
	notech_ao4 i_1050(.A(n_58762), .B(n_43158), .C(n_58619), .D(n_43143), .Z
		(n_314699478));
	notech_ao4 i_1051(.A(n_58720), .B(n_43048), .C(n_58445), .D(n_43174), .Z
		(n_3147));
	notech_and4 i_1060(.A(n_3147), .B(n_314699478), .C(n_3144), .D(n_192998399
		), .Z(n_3149));
	notech_ao4 i_1052(.A(n_58884), .B(n_43021), .C(n_58783), .D(n_43190), .Z
		(n_3150));
	notech_ao4 i_1053(.A(n_58903), .B(n_43013), .C(n_58646), .D(n_43064), .Z
		(n_3151));
	notech_ao4 i_1054(.A(n_58865), .B(n_43080), .C(n_58938), .D(n_43005), .Z
		(n_3153));
	notech_ao4 i_1055(.A(n_58846), .B(n_43095), .C(n_58956), .D(n_43127), .Z
		(n_3154));
	notech_and4 i_1061(.A(n_3154), .B(n_3153), .C(n_3151), .D(n_3150), .Z(n_3156
		));
	notech_ao4 i_1080(.A(n_58625), .B(n_43038), .C(n_58741), .D(n_43030), .Z
		(n_315899480));
	notech_ao4 i_1081(.A(n_58762), .B(n_43160), .C(n_58619), .D(n_43144), .Z
		(n_3160));
	notech_ao4 i_1082(.A(n_58720), .B(n_43050), .C(n_58445), .D(n_43176), .Z
		(n_3161));
	notech_and4 i_1091(.A(n_3161), .B(n_3160), .C(n_315899480), .D(n_194698416
		), .Z(n_3163));
	notech_ao4 i_1083(.A(n_58884), .B(n_43022), .C(n_58783), .D(n_43192), .Z
		(n_316499481));
	notech_ao4 i_1084(.A(n_58903), .B(n_43014), .C(n_58646), .D(n_43066), .Z
		(n_3165));
	notech_ao4 i_1085(.A(n_58865), .B(n_43082), .C(n_58938), .D(n_43006), .Z
		(n_3167));
	notech_ao4 i_1086(.A(n_58846), .B(n_43097), .C(n_58956), .D(n_43129), .Z
		(n_3168));
	notech_and4 i_1092(.A(n_3168), .B(n_3167), .C(n_3165), .D(n_316499481), 
		.Z(n_317099482));
	notech_ao4 i_1111(.A(n_58625), .B(n_43039), .C(n_58741), .D(n_43031), .Z
		(n_3172));
	notech_ao4 i_1112(.A(n_58762), .B(n_43162), .C(n_58619), .D(n_43146), .Z
		(n_3174));
	notech_ao4 i_1113(.A(n_58720), .B(n_43052), .C(n_58447), .D(n_43178), .Z
		(n_3175));
	notech_and4 i_1122(.A(n_3175), .B(n_3174), .C(n_3172), .D(n_196398433), 
		.Z(n_3177));
	notech_ao4 i_1114(.A(n_58884), .B(n_43023), .C(n_58783), .D(n_43194), .Z
		(n_3178));
	notech_ao4 i_1115(.A(n_58903), .B(n_43015), .C(n_58646), .D(n_43068), .Z
		(n_3179));
	notech_ao4 i_1116(.A(n_58865), .B(n_43084), .C(n_58938), .D(n_43007), .Z
		(n_3181));
	notech_ao4 i_1117(.A(n_58846), .B(n_43099), .C(n_58956), .D(n_43131), .Z
		(n_318299484));
	notech_and4 i_1123(.A(n_318299484), .B(n_3181), .C(n_3179), .D(n_3178), 
		.Z(n_3184));
	notech_ao4 i_1142(.A(n_58625), .B(n_43040), .C(n_58741), .D(n_43032), .Z
		(n_3186));
	notech_ao4 i_1143(.A(n_58762), .B(n_43164), .C(n_58619), .D(n_43148), .Z
		(n_318899485));
	notech_ao4 i_1144(.A(n_58720), .B(n_43054), .C(n_58447), .D(n_43180), .Z
		(n_3189));
	notech_and4 i_1153(.A(n_3189), .B(n_318899485), .C(n_3186), .D(n_198098450
		), .Z(n_3191));
	notech_ao4 i_1145(.A(n_58884), .B(n_43024), .C(n_58783), .D(n_43196), .Z
		(n_3192));
	notech_ao4 i_1146(.A(n_58903), .B(n_43016), .C(n_58646), .D(n_43070), .Z
		(n_3193));
	notech_ao4 i_1147(.A(n_58865), .B(n_43085), .C(n_58938), .D(n_43008), .Z
		(n_3195));
	notech_ao4 i_1148(.A(n_58846), .B(n_43101), .C(n_58956), .D(n_43133), .Z
		(n_3196));
	notech_and4 i_1154(.A(n_3196), .B(n_3195), .C(n_3193), .D(n_3192), .Z(n_3198
		));
	notech_ao4 i_1173(.A(n_58625), .B(n_43041), .C(n_58741), .D(n_43033), .Z
		(n_320099487));
	notech_ao4 i_1174(.A(n_58762), .B(n_43166), .C(n_58619), .D(n_43150), .Z
		(n_3202));
	notech_ao4 i_1175(.A(n_58720), .B(n_43056), .C(n_58447), .D(n_43182), .Z
		(n_3203));
	notech_and4 i_1184(.A(n_3203), .B(n_3202), .C(n_320099487), .D(n_199798467
		), .Z(n_3205));
	notech_ao4 i_1176(.A(n_58884), .B(n_43025), .C(n_58783), .D(n_43198), .Z
		(n_320699488));
	notech_ao4 i_1177(.A(n_58903), .B(n_43017), .C(n_58646), .D(n_43072), .Z
		(n_3207));
	notech_ao4 i_1178(.A(n_58865), .B(n_43087), .C(n_58938), .D(n_43009), .Z
		(n_3209));
	notech_ao4 i_1179(.A(n_58846), .B(n_43103), .C(n_58956), .D(n_43135), .Z
		(n_3210));
	notech_and4 i_1185(.A(n_3210), .B(n_3209), .C(n_3207), .D(n_320699488), 
		.Z(n_321299489));
	notech_ao4 i_1204(.A(n_58625), .B(n_43042), .C(n_58741), .D(n_43034), .Z
		(n_3214));
	notech_ao4 i_1205(.A(n_58762), .B(n_43168), .C(n_58621), .D(n_43152), .Z
		(n_3216));
	notech_ao4 i_1206(.A(n_58720), .B(n_43058), .C(n_58447), .D(n_43184), .Z
		(n_3217));
	notech_and4 i_1215(.A(n_3217), .B(n_3216), .C(n_3214), .D(n_201498484), 
		.Z(n_3219));
	notech_ao4 i_1207(.A(n_58885), .B(n_43026), .C(n_58783), .D(n_43200), .Z
		(n_3220));
	notech_ao4 i_1208(.A(n_58903), .B(n_43018), .C(n_58646), .D(n_43074), .Z
		(n_3221));
	notech_ao4 i_1209(.A(n_58866), .B(n_43089), .C(n_58931), .D(n_43010), .Z
		(n_3223));
	notech_ao4 i_1210(.A(n_58847), .B(n_43105), .C(n_58957), .D(n_43137), .Z
		(n_322499491));
	notech_and4 i_1216(.A(n_322499491), .B(n_3223), .C(n_3221), .D(n_3220), 
		.Z(n_3226));
	notech_ao4 i_1235(.A(n_58625), .B(n_43044), .C(n_58741), .D(n_43035), .Z
		(n_3228));
	notech_ao4 i_1236(.A(n_58762), .B(n_43170), .C(n_58619), .D(n_43154), .Z
		(n_323099492));
	notech_ao4 i_1237(.A(n_58720), .B(n_43060), .C(n_58435), .D(n_43186), .Z
		(n_3231));
	notech_and4 i_1246(.A(n_3231), .B(n_323099492), .C(n_3228), .D(n_203198501
		), .Z(n_3233));
	notech_ao4 i_1238(.A(n_58885), .B(n_43027), .C(n_58783), .D(n_43201), .Z
		(n_3234));
	notech_ao4 i_1239(.A(n_58903), .B(n_43019), .C(n_58646), .D(n_43076), .Z
		(n_3235));
	notech_ao4 i_1240(.A(n_58866), .B(n_43091), .C(n_58924), .D(n_43011), .Z
		(n_3237));
	notech_ao4 i_1241(.A(n_58847), .B(n_43107), .C(n_58957), .D(n_43139), .Z
		(n_3238));
	notech_and4 i_1247(.A(n_3238), .B(n_3237), .C(n_3235), .D(n_3234), .Z(n_3240
		));
	notech_ao4 i_1266(.A(n_58625), .B(n_43046), .C(n_58741), .D(n_43036), .Z
		(n_324299494));
	notech_ao4 i_1267(.A(n_58762), .B(n_43172), .C(n_58619), .D(n_43156), .Z
		(n_3244));
	notech_ao4 i_1268(.A(n_58720), .B(n_43062), .C(n_58435), .D(n_43188), .Z
		(n_3245));
	notech_and4 i_1277(.A(n_3245), .B(n_3244), .C(n_324299494), .D(n_204898518
		), .Z(n_3247));
	notech_ao4 i_1269(.A(n_58885), .B(n_43028), .C(n_58783), .D(n_43203), .Z
		(n_324899495));
	notech_ao4 i_1270(.A(n_58903), .B(n_43020), .C(n_58646), .D(n_43078), .Z
		(n_3249));
	notech_ao4 i_1271(.A(n_58866), .B(n_43093), .C(n_58924), .D(n_43012), .Z
		(n_3251));
	notech_ao4 i_1272(.A(n_58847), .B(n_43109), .C(n_58957), .D(n_43141), .Z
		(n_3252));
	notech_and4 i_1278(.A(n_3252), .B(n_3251), .C(n_3249), .D(n_324899495), 
		.Z(n_325499496));
	notech_ao4 i_1297(.A(n_58625), .B(n_43048), .C(n_58741), .D(n_43037), .Z
		(n_3256));
	notech_ao4 i_1298(.A(n_58762), .B(n_43174), .C(n_58619), .D(n_43158), .Z
		(n_3258));
	notech_ao4 i_1299(.A(n_58720), .B(n_43064), .C(n_58435), .D(n_43190), .Z
		(n_3259));
	notech_and4 i_1308(.A(n_3259), .B(n_3258), .C(n_3256), .D(n_206598535), 
		.Z(n_3262));
	notech_ao4 i_1300(.A(n_58885), .B(n_43029), .C(n_58783), .D(n_43205), .Z
		(n_3263));
	notech_ao4 i_1301(.A(n_58903), .B(n_43021), .C(n_58646), .D(n_43080), .Z
		(n_3264));
	notech_ao4 i_1302(.A(n_58866), .B(n_43095), .C(n_58924), .D(n_43013), .Z
		(n_326699497));
	notech_ao4 i_1303(.A(n_58847), .B(n_43111), .C(n_58957), .D(n_43143), .Z
		(n_3267));
	notech_and4 i_1309(.A(n_3267), .B(n_326699497), .C(n_3264), .D(n_3263), 
		.Z(n_3269));
	notech_ao4 i_1328(.A(n_58625), .B(n_43050), .C(n_58741), .D(n_43038), .Z
		(n_3271));
	notech_ao4 i_1329(.A(n_58762), .B(n_43176), .C(n_58619), .D(n_43160), .Z
		(n_3273));
	notech_ao4 i_1330(.A(n_58720), .B(n_43066), .C(n_58435), .D(n_43192), .Z
		(n_3274));
	notech_and4 i_1339(.A(n_3274), .B(n_3273), .C(n_3271), .D(n_208298552), 
		.Z(n_3276));
	notech_ao4 i_1331(.A(n_58885), .B(n_43030), .C(n_58783), .D(n_43207), .Z
		(n_3277));
	notech_ao4 i_1332(.A(n_58903), .B(n_43022), .C(n_58646), .D(n_43082), .Z
		(n_327899499));
	notech_ao4 i_1333(.A(n_58866), .B(n_43097), .C(n_58924), .D(n_43014), .Z
		(n_3280));
	notech_ao4 i_1334(.A(n_58847), .B(n_43113), .C(n_58957), .D(n_43144), .Z
		(n_3281));
	notech_and4 i_1340(.A(n_3281), .B(n_3280), .C(n_327899499), .D(n_3277), 
		.Z(n_3283));
	notech_ao4 i_1359(.A(n_58625), .B(n_43052), .C(n_58741), .D(n_43039), .Z
		(n_3285));
	notech_ao4 i_1360(.A(n_58762), .B(n_43178), .C(n_58614), .D(n_43162), .Z
		(n_3287));
	notech_ao4 i_1361(.A(n_58720), .B(n_43068), .C(n_58435), .D(n_43194), .Z
		(n_3288));
	notech_and4 i_1370(.A(n_3288), .B(n_3287), .C(n_3285), .D(n_209998569), 
		.Z(n_329099501));
	notech_ao4 i_1362(.A(n_58885), .B(n_43031), .C(n_58783), .D(n_43209), .Z
		(n_3291));
	notech_ao4 i_1363(.A(n_58903), .B(n_43023), .C(n_58646), .D(n_43084), .Z
		(n_3292));
	notech_ao4 i_1364(.A(n_58866), .B(n_43099), .C(n_58924), .D(n_43015), .Z
		(n_3294));
	notech_ao4 i_1365(.A(n_58847), .B(n_43115), .C(n_58957), .D(n_43146), .Z
		(n_3295));
	notech_and4 i_1371(.A(n_3295), .B(n_3294), .C(n_3292), .D(n_3291), .Z(n_3297
		));
	notech_ao4 i_1390(.A(n_58625), .B(n_43054), .C(n_58741), .D(n_43040), .Z
		(n_3299));
	notech_ao4 i_1391(.A(n_58762), .B(n_43180), .C(n_58607), .D(n_43164), .Z
		(n_3301));
	notech_ao4 i_1392(.A(n_58720), .B(n_43070), .C(n_58435), .D(n_43196), .Z
		(n_330299503));
	notech_and4 i_1401(.A(n_330299503), .B(n_3301), .C(n_3299), .D(n_211698586
		), .Z(n_3304));
	notech_ao4 i_1393(.A(n_58885), .B(n_43032), .C(n_58783), .D(n_43211), .Z
		(n_3305));
	notech_ao4 i_1394(.A(n_58903), .B(n_43024), .C(n_58646), .D(n_43085), .Z
		(n_3306));
	notech_ao4 i_1395(.A(n_58866), .B(n_43101), .C(n_58924), .D(n_43016), .Z
		(n_330899504));
	notech_ao4 i_1396(.A(n_58847), .B(n_43117), .C(n_58957), .D(n_43148), .Z
		(n_3309));
	notech_and4 i_1402(.A(n_3309), .B(n_330899504), .C(n_3306), .D(n_3305), 
		.Z(n_3311));
	notech_ao4 i_1421(.A(n_58625), .B(n_43056), .C(n_58741), .D(n_43041), .Z
		(n_3313));
	notech_ao4 i_1422(.A(n_58762), .B(n_43182), .C(n_58607), .D(n_43166), .Z
		(n_3315));
	notech_ao4 i_1423(.A(n_58720), .B(n_43072), .C(n_58445), .D(n_43198), .Z
		(n_3316));
	notech_and4 i_1432(.A(n_3316), .B(n_3315), .C(n_3313), .D(n_213398603), 
		.Z(n_3318));
	notech_ao4 i_1424(.A(n_58885), .B(n_43033), .C(n_58783), .D(n_43213), .Z
		(n_3319));
	notech_ao4 i_1425(.A(n_58903), .B(n_43025), .C(n_58646), .D(n_43087), .Z
		(n_332099506));
	notech_ao4 i_1426(.A(n_58866), .B(n_43103), .C(n_58930), .D(n_43017), .Z
		(n_3322));
	notech_ao4 i_1427(.A(n_58847), .B(n_43119), .C(n_58957), .D(n_43150), .Z
		(n_3323));
	notech_and4 i_1433(.A(n_3323), .B(n_3322), .C(n_332099506), .D(n_3319), 
		.Z(n_3325));
	notech_ao4 i_1452(.A(n_58632), .B(n_43058), .C(n_58748), .D(n_43042), .Z
		(n_3327));
	notech_ao4 i_1453(.A(n_58769), .B(n_43184), .C(n_58609), .D(n_43168), .Z
		(n_3329));
	notech_ao4 i_1454(.A(n_58727), .B(n_43074), .C(n_58435), .D(n_43200), .Z
		(n_3330));
	notech_and4 i_1463(.A(n_3330), .B(n_3329), .C(n_3327), .D(n_215098620), 
		.Z(n_333299508));
	notech_ao4 i_1455(.A(n_58890), .B(n_43034), .C(n_58790), .D(n_43215), .Z
		(n_3333));
	notech_ao4 i_1456(.A(n_58910), .B(n_43026), .C(n_58653), .D(n_43089), .Z
		(n_3334));
	notech_ao4 i_1457(.A(n_58871), .B(n_43105), .C(n_58930), .D(n_43018), .Z
		(n_3336));
	notech_ao4 i_1458(.A(n_58852), .B(n_43121), .C(n_58962), .D(n_43152), .Z
		(n_3337));
	notech_and4 i_1464(.A(n_3337), .B(n_3336), .C(n_3334), .D(n_3333), .Z(n_3339
		));
	notech_ao4 i_1483(.A(n_58632), .B(n_43060), .C(n_58748), .D(n_43044), .Z
		(n_3341));
	notech_ao4 i_1484(.A(n_58769), .B(n_43186), .C(n_58607), .D(n_43170), .Z
		(n_3343));
	notech_ao4 i_1485(.A(n_58727), .B(n_43076), .C(n_58435), .D(n_43201), .Z
		(n_334499510));
	notech_and4 i_1494(.A(n_334499510), .B(n_3343), .C(n_3341), .D(n_216798637
		), .Z(n_3346));
	notech_ao4 i_1486(.A(n_58890), .B(n_43035), .C(n_58790), .D(n_43217), .Z
		(n_3347));
	notech_ao4 i_1487(.A(n_58910), .B(n_43027), .C(n_58653), .D(n_43091), .Z
		(n_3348));
	notech_ao4 i_1488(.A(n_58871), .B(n_43107), .C(n_58930), .D(n_43019), .Z
		(n_335099511));
	notech_ao4 i_1489(.A(n_58852), .B(n_43123), .C(n_58962), .D(n_43154), .Z
		(n_3351));
	notech_and4 i_1495(.A(n_3351), .B(n_335099511), .C(n_3348), .D(n_3347), 
		.Z(n_3353));
	notech_ao4 i_1514(.A(n_58632), .B(n_43062), .C(n_58748), .D(n_43046), .Z
		(n_3355));
	notech_ao4 i_1515(.A(n_58769), .B(n_43188), .C(n_58607), .D(n_43172), .Z
		(n_3357));
	notech_ao4 i_1516(.A(n_58727), .B(n_43078), .C(n_58435), .D(n_43203), .Z
		(n_3358));
	notech_and4 i_1525(.A(n_3358), .B(n_3357), .C(n_3355), .D(n_218498654), 
		.Z(n_3360));
	notech_ao4 i_1517(.A(n_58890), .B(n_43036), .C(n_58790), .D(n_43219), .Z
		(n_3361));
	notech_ao4 i_1518(.A(n_58910), .B(n_43028), .C(n_58653), .D(n_43093), .Z
		(n_336299513));
	notech_ao4 i_1519(.A(n_58871), .B(n_43109), .C(n_58930), .D(n_43020), .Z
		(n_3364));
	notech_ao4 i_1520(.A(n_58852), .B(n_43125), .C(n_58962), .D(n_43156), .Z
		(n_3365));
	notech_and4 i_1526(.A(n_3365), .B(n_3364), .C(n_336299513), .D(n_3361), 
		.Z(n_3367));
	notech_ao4 i_1545(.A(n_58632), .B(n_43064), .C(n_58748), .D(n_43048), .Z
		(n_3369));
	notech_ao4 i_1546(.A(n_58769), .B(n_43190), .C(n_58607), .D(n_43174), .Z
		(n_3371));
	notech_ao4 i_1547(.A(n_58727), .B(n_43080), .C(n_58435), .D(n_43205), .Z
		(n_3372));
	notech_and4 i_1556(.A(n_3372), .B(n_3371), .C(n_3369), .D(n_220198671), 
		.Z(n_337499515));
	notech_ao4 i_1548(.A(n_58890), .B(n_43037), .C(n_58790), .D(n_43221), .Z
		(n_3375));
	notech_ao4 i_1549(.A(n_58910), .B(n_43029), .C(n_58653), .D(n_43095), .Z
		(n_3376));
	notech_ao4 i_1550(.A(n_58871), .B(n_43111), .C(n_58930), .D(n_43021), .Z
		(n_3378));
	notech_ao4 i_1551(.A(n_58852), .B(n_43127), .C(n_58962), .D(n_43158), .Z
		(n_3379));
	notech_and4 i_1557(.A(n_3379), .B(n_3378), .C(n_3376), .D(n_3375), .Z(n_3381
		));
	notech_ao4 i_1576(.A(n_58632), .B(n_43066), .C(n_58748), .D(n_43050), .Z
		(n_3383));
	notech_ao4 i_1577(.A(n_58769), .B(n_43192), .C(n_58607), .D(n_43176), .Z
		(n_3385));
	notech_ao4 i_1578(.A(n_58727), .B(n_43082), .C(n_58435), .D(n_43207), .Z
		(n_338699517));
	notech_and4 i_1587(.A(n_338699517), .B(n_3385), .C(n_3383), .D(n_221898688
		), .Z(n_3388));
	notech_ao4 i_1579(.A(n_58890), .B(n_43038), .C(n_58790), .D(n_43223), .Z
		(n_3389));
	notech_ao4 i_1580(.A(n_58910), .B(n_43030), .C(n_58653), .D(n_43097), .Z
		(n_3390));
	notech_ao4 i_1581(.A(n_58871), .B(n_43113), .C(n_58924), .D(n_43022), .Z
		(n_339299518));
	notech_ao4 i_1582(.A(n_58852), .B(n_43129), .C(n_58962), .D(n_43160), .Z
		(n_3393));
	notech_and4 i_1588(.A(n_3393), .B(n_339299518), .C(n_3390), .D(n_3389), 
		.Z(n_3395));
	notech_ao4 i_1607(.A(n_58632), .B(n_43068), .C(n_58748), .D(n_43052), .Z
		(n_3397));
	notech_ao4 i_1608(.A(n_58769), .B(n_43194), .C(n_58609), .D(n_43178), .Z
		(n_3399));
	notech_ao4 i_1609(.A(n_58727), .B(n_43084), .C(n_58435), .D(n_43209), .Z
		(n_3400));
	notech_and4 i_1618(.A(n_3400), .B(n_3399), .C(n_3397), .D(n_223598705), 
		.Z(n_3402));
	notech_ao4 i_1610(.A(n_58890), .B(n_43039), .C(n_58790), .D(n_43225), .Z
		(n_3403));
	notech_ao4 i_1611(.A(n_58910), .B(n_43031), .C(n_58653), .D(n_43099), .Z
		(n_340499520));
	notech_ao4 i_1612(.A(n_58871), .B(n_43115), .C(n_58924), .D(n_43023), .Z
		(n_3406));
	notech_ao4 i_1613(.A(n_58852), .B(n_43131), .C(n_58962), .D(n_43162), .Z
		(n_3407));
	notech_and4 i_1619(.A(n_3407), .B(n_3406), .C(n_340499520), .D(n_3403), 
		.Z(n_3409));
	notech_ao4 i_1638(.A(n_58632), .B(n_43070), .C(n_58748), .D(n_43054), .Z
		(n_3411));
	notech_ao4 i_1639(.A(n_58769), .B(n_43196), .C(n_58609), .D(n_43180), .Z
		(n_3413));
	notech_ao4 i_1640(.A(n_58727), .B(n_43085), .C(n_58435), .D(n_43211), .Z
		(n_3414));
	notech_and4 i_1649(.A(n_3414), .B(n_3413), .C(n_3411), .D(n_225298722), 
		.Z(n_341699522));
	notech_ao4 i_1641(.A(n_58890), .B(n_43040), .C(n_58790), .D(n_43227), .Z
		(n_3417));
	notech_ao4 i_1642(.A(n_58910), .B(n_43032), .C(n_58653), .D(n_43101), .Z
		(n_3418));
	notech_ao4 i_1643(.A(n_58871), .B(n_43117), .C(n_58924), .D(n_43024), .Z
		(n_3420));
	notech_ao4 i_1644(.A(n_58852), .B(n_43133), .C(n_58962), .D(n_43164), .Z
		(n_3421));
	notech_and4 i_1650(.A(n_3421), .B(n_3420), .C(n_3418), .D(n_3417), .Z(n_3423
		));
	notech_ao4 i_1669(.A(n_58632), .B(n_43072), .C(n_58748), .D(n_43056), .Z
		(n_3425));
	notech_ao4 i_1670(.A(n_58769), .B(n_43198), .C(n_58609), .D(n_43182), .Z
		(n_3427));
	notech_ao4 i_1671(.A(n_58727), .B(n_43087), .C(n_58435), .D(n_43213), .Z
		(n_342899524));
	notech_and4 i_1680(.A(n_342899524), .B(n_3427), .C(n_3425), .D(n_226998739
		), .Z(n_3430));
	notech_ao4 i_1672(.A(n_58890), .B(n_43041), .C(n_58790), .D(n_43229), .Z
		(n_3431));
	notech_ao4 i_1673(.A(n_58910), .B(n_43033), .C(n_58653), .D(n_43103), .Z
		(n_3432));
	notech_ao4 i_1674(.A(n_58871), .B(n_43119), .C(n_58924), .D(n_43025), .Z
		(n_343499525));
	notech_ao4 i_1675(.A(n_58852), .B(n_43135), .C(n_58962), .D(n_43166), .Z
		(n_3435));
	notech_and4 i_1681(.A(n_3435), .B(n_343499525), .C(n_3432), .D(n_3431), 
		.Z(n_3437));
	notech_ao4 i_1700(.A(n_58632), .B(n_43074), .C(n_58748), .D(n_43058), .Z
		(n_3439));
	notech_ao4 i_1701(.A(n_58769), .B(n_43200), .C(n_58609), .D(n_43184), .Z
		(n_3441));
	notech_ao4 i_1702(.A(n_58727), .B(n_43089), .C(n_58435), .D(n_43215), .Z
		(n_3442));
	notech_and4 i_1711(.A(n_3442), .B(n_3441), .C(n_3439), .D(n_228698756), 
		.Z(n_3444));
	notech_ao4 i_1703(.A(n_58892), .B(n_43042), .C(n_58790), .D(n_43231), .Z
		(n_3445));
	notech_ao4 i_1704(.A(n_58910), .B(n_43034), .C(n_58653), .D(n_43105), .Z
		(n_344699527));
	notech_ao4 i_1705(.A(n_58873), .B(n_43121), .C(n_58924), .D(n_43026), .Z
		(n_3448));
	notech_ao4 i_1706(.A(n_58854), .B(n_43137), .C(n_58964), .D(n_43168), .Z
		(n_3449));
	notech_and4 i_1712(.A(n_3449), .B(n_3448), .C(n_344699527), .D(n_3445), 
		.Z(n_3451));
	notech_ao4 i_1731(.A(n_58632), .B(n_43076), .C(n_58748), .D(n_43060), .Z
		(n_3453));
	notech_ao4 i_1732(.A(n_58769), .B(n_43201), .C(n_58609), .D(n_43186), .Z
		(n_3455));
	notech_ao4 i_1733(.A(n_58727), .B(n_43091), .C(n_58435), .D(n_43217), .Z
		(n_3456));
	notech_and4 i_1742(.A(n_3456), .B(n_3455), .C(n_3453), .D(n_230398773), 
		.Z(n_345899529));
	notech_ao4 i_1734(.A(n_58892), .B(n_43044), .C(n_58790), .D(n_43233), .Z
		(n_3459));
	notech_ao4 i_1735(.A(n_58910), .B(n_43035), .C(n_58653), .D(n_43107), .Z
		(n_3460));
	notech_ao4 i_1736(.A(n_58873), .B(n_43123), .C(n_58924), .D(n_43027), .Z
		(n_3462));
	notech_ao4 i_1737(.A(n_58854), .B(n_43139), .C(n_58962), .D(n_43170), .Z
		(n_3463));
	notech_and4 i_1743(.A(n_3463), .B(n_3462), .C(n_3460), .D(n_3459), .Z(n_3465
		));
	notech_ao4 i_1762(.A(n_58632), .B(n_43078), .C(n_58748), .D(n_43062), .Z
		(n_3467));
	notech_ao4 i_1763(.A(n_58769), .B(n_43203), .C(n_58609), .D(n_43188), .Z
		(n_3469));
	notech_ao4 i_1764(.A(n_58727), .B(n_43093), .C(n_58435), .D(n_43219), .Z
		(n_347099531));
	notech_and4 i_1773(.A(n_347099531), .B(n_3469), .C(n_3467), .D(n_232098790
		), .Z(n_3472));
	notech_ao4 i_1765(.A(n_58892), .B(n_43046), .C(n_58790), .D(n_43235), .Z
		(n_3473));
	notech_ao4 i_1766(.A(n_58910), .B(n_43036), .C(n_58653), .D(n_43109), .Z
		(n_3474));
	notech_ao4 i_1767(.A(n_58873), .B(n_43125), .C(n_58924), .D(n_43028), .Z
		(n_347699532));
	notech_ao4 i_1768(.A(n_58854), .B(n_43141), .C(n_58964), .D(n_43172), .Z
		(n_3477));
	notech_and4 i_1774(.A(n_3477), .B(n_347699532), .C(n_3474), .D(n_3473), 
		.Z(n_3479));
	notech_ao4 i_1793(.A(n_58632), .B(n_43080), .C(n_58748), .D(n_43064), .Z
		(n_3481));
	notech_ao4 i_1794(.A(n_58769), .B(n_43205), .C(n_58609), .D(n_43190), .Z
		(n_3483));
	notech_ao4 i_1795(.A(n_58727), .B(n_43095), .C(n_58435), .D(n_43221), .Z
		(n_3484));
	notech_and4 i_1804(.A(n_3484), .B(n_3483), .C(n_3481), .D(n_233798807), 
		.Z(n_3486));
	notech_ao4 i_1796(.A(n_58892), .B(n_43048), .C(n_58790), .D(n_43237), .Z
		(n_3487));
	notech_ao4 i_1797(.A(n_58910), .B(n_43037), .C(n_58653), .D(n_43111), .Z
		(n_348899534));
	notech_ao4 i_1798(.A(n_58873), .B(n_43127), .C(n_58924), .D(n_43029), .Z
		(n_3490));
	notech_ao4 i_1799(.A(n_58854), .B(n_43143), .C(n_58964), .D(n_43174), .Z
		(n_3491));
	notech_and4 i_1805(.A(n_3491), .B(n_3490), .C(n_348899534), .D(n_3487), 
		.Z(n_3493));
	notech_ao4 i_1824(.A(n_58632), .B(n_43082), .C(n_58748), .D(n_43066), .Z
		(n_3495));
	notech_ao4 i_1825(.A(n_58769), .B(n_43207), .C(n_58607), .D(n_43192), .Z
		(n_3497));
	notech_ao4 i_1826(.A(n_58727), .B(n_43097), .C(n_58445), .D(n_43223), .Z
		(n_3498));
	notech_and4 i_1835(.A(n_3498), .B(n_3497), .C(n_3495), .D(n_235498824), 
		.Z(n_350099536));
	notech_ao4 i_1827(.A(n_58892), .B(n_43050), .C(n_58790), .D(n_43239), .Z
		(n_3501));
	notech_ao4 i_1828(.A(n_58910), .B(n_43038), .C(n_58653), .D(n_43113), .Z
		(n_3502));
	notech_ao4 i_1829(.A(n_58873), .B(n_43129), .C(n_58924), .D(n_43030), .Z
		(n_3504));
	notech_ao4 i_1830(.A(n_58854), .B(n_43144), .C(n_58962), .D(n_43176), .Z
		(n_3505));
	notech_and4 i_1836(.A(n_3505), .B(n_3504), .C(n_3502), .D(n_3501), .Z(n_3507
		));
	notech_ao4 i_1855(.A(n_58632), .B(n_43084), .C(n_58748), .D(n_43068), .Z
		(n_3509));
	notech_ao4 i_1856(.A(n_58769), .B(n_43209), .C(n_58606), .D(n_43194), .Z
		(n_3511));
	notech_ao4 i_1857(.A(n_58727), .B(n_43099), .C(n_58441), .D(n_43225), .Z
		(n_351299538));
	notech_and4 i_1866(.A(n_351299538), .B(n_3511), .C(n_3509), .D(n_237198841
		), .Z(n_3514));
	notech_ao4 i_1858(.A(n_58890), .B(n_43052), .C(n_58790), .D(n_43241), .Z
		(n_3515));
	notech_ao4 i_1859(.A(n_58910), .B(n_43039), .C(n_58653), .D(n_43115), .Z
		(n_3516));
	notech_ao4 i_1860(.A(n_58871), .B(n_43131), .C(n_58924), .D(n_43031), .Z
		(n_351899539));
	notech_ao4 i_1861(.A(n_58852), .B(n_43146), .C(n_58962), .D(n_43178), .Z
		(n_3519));
	notech_and4 i_1867(.A(n_3519), .B(n_351899539), .C(n_3516), .D(n_3515), 
		.Z(n_3521));
	notech_ao4 i_1886(.A(n_58632), .B(n_43085), .C(n_58748), .D(n_43070), .Z
		(n_3523));
	notech_ao4 i_1887(.A(n_58769), .B(n_43211), .C(n_58606), .D(n_43196), .Z
		(n_3525));
	notech_ao4 i_1888(.A(n_58727), .B(n_43101), .C(n_58441), .D(n_43227), .Z
		(n_3526));
	notech_and4 i_1897(.A(n_3526), .B(n_3525), .C(n_3523), .D(n_238898858), 
		.Z(n_3528));
	notech_ao4 i_1889(.A(n_58892), .B(n_43054), .C(n_58790), .D(n_43243), .Z
		(n_3529));
	notech_ao4 i_1890(.A(n_58910), .B(n_43040), .C(n_58653), .D(n_43117), .Z
		(n_353099541));
	notech_ao4 i_1891(.A(n_58873), .B(n_43133), .C(n_58924), .D(n_43032), .Z
		(n_3532));
	notech_ao4 i_1892(.A(n_58854), .B(n_43148), .C(n_58962), .D(n_43180), .Z
		(n_3533));
	notech_and4 i_1898(.A(n_3533), .B(n_3532), .C(n_353099541), .D(n_3529), 
		.Z(n_3535));
	notech_ao4 i_1917(.A(n_58632), .B(n_43087), .C(n_58748), .D(n_43072), .Z
		(n_3537));
	notech_ao4 i_1918(.A(n_58769), .B(n_43213), .C(n_58606), .D(n_43198), .Z
		(n_3539));
	notech_ao4 i_1919(.A(n_58727), .B(n_43103), .C(n_58441), .D(n_43229), .Z
		(n_3540));
	notech_and4 i_1928(.A(n_3540), .B(n_3539), .C(n_3537), .D(n_240598875), 
		.Z(n_354299543));
	notech_ao4 i_1920(.A(n_58892), .B(n_43056), .C(n_58790), .D(n_43245), .Z
		(n_3543));
	notech_ao4 i_1921(.A(n_58910), .B(n_43041), .C(n_58653), .D(n_43119), .Z
		(n_3544));
	notech_ao4 i_1922(.A(n_58873), .B(n_43135), .C(n_58931), .D(n_43033), .Z
		(n_3546));
	notech_ao4 i_1923(.A(n_58854), .B(n_43150), .C(n_58962), .D(n_43182), .Z
		(n_3547));
	notech_and4 i_1929(.A(n_3547), .B(n_3546), .C(n_3544), .D(n_3543), .Z(n_3549
		));
	notech_ao4 i_1948(.A(n_58630), .B(n_43089), .C(n_58746), .D(n_43074), .Z
		(n_3551));
	notech_ao4 i_1949(.A(n_58767), .B(n_43215), .C(n_58606), .D(n_43200), .Z
		(n_3553));
	notech_ao4 i_1950(.A(n_58725), .B(n_43105), .C(n_58441), .D(n_43231), .Z
		(n_355499545));
	notech_and4 i_1959(.A(n_355499545), .B(n_3553), .C(n_3551), .D(n_242398889
		), .Z(n_3556));
	notech_ao4 i_1951(.A(n_58887), .B(n_43058), .C(n_58788), .D(n_43247), .Z
		(n_3557));
	notech_ao4 i_1952(.A(n_58908), .B(n_43042), .C(n_58651), .D(n_43121), .Z
		(n_3558));
	notech_ao4 i_1953(.A(n_58868), .B(n_43137), .C(n_58931), .D(n_43034), .Z
		(n_356099546));
	notech_ao4 i_1954(.A(n_58849), .B(n_43152), .C(n_58959), .D(n_43184), .Z
		(n_3561));
	notech_and4 i_1960(.A(n_3561), .B(n_356099546), .C(n_3558), .D(n_3557), 
		.Z(n_3563));
	notech_ao4 i_1979(.A(n_58630), .B(n_43091), .C(n_58746), .D(n_43076), .Z
		(n_3565));
	notech_ao4 i_1980(.A(n_58767), .B(n_43217), .C(n_58606), .D(n_43201), .Z
		(n_3567));
	notech_ao4 i_1981(.A(n_58725), .B(n_43107), .C(n_58441), .D(n_43233), .Z
		(n_3568));
	notech_and4 i_1990(.A(n_3568), .B(n_3567), .C(n_3565), .D(n_244098906), 
		.Z(n_3570));
	notech_ao4 i_1982(.A(n_58887), .B(n_43060), .C(n_58788), .D(n_43249), .Z
		(n_3571));
	notech_ao4 i_1983(.A(n_58908), .B(n_43044), .C(n_58651), .D(n_43123), .Z
		(n_357299548));
	notech_ao4 i_1984(.A(n_58868), .B(n_43139), .C(n_58931), .D(n_43035), .Z
		(n_3574));
	notech_ao4 i_1985(.A(n_58849), .B(n_43154), .C(n_58959), .D(n_43186), .Z
		(n_3575));
	notech_and4 i_1991(.A(n_3575), .B(n_3574), .C(n_357299548), .D(n_3571), 
		.Z(n_3577));
	notech_ao4 i_2010(.A(n_58630), .B(n_43093), .C(n_58746), .D(n_43078), .Z
		(n_3579));
	notech_ao4 i_2011(.A(n_58767), .B(n_43219), .C(n_58606), .D(n_43203), .Z
		(n_3581));
	notech_ao4 i_2012(.A(n_58725), .B(n_43109), .C(n_58441), .D(n_43235), .Z
		(n_3582));
	notech_and4 i_2021(.A(n_3582), .B(n_3581), .C(n_3579), .D(n_245798923), 
		.Z(n_358499550));
	notech_ao4 i_2013(.A(n_58887), .B(n_43062), .C(n_58788), .D(n_43251), .Z
		(n_3585));
	notech_ao4 i_2014(.A(n_58908), .B(n_43046), .C(n_58651), .D(n_43125), .Z
		(n_3586));
	notech_ao4 i_2015(.A(n_58868), .B(n_43141), .C(n_58930), .D(n_43036), .Z
		(n_3588));
	notech_ao4 i_2016(.A(n_58849), .B(n_43156), .C(n_58959), .D(n_43188), .Z
		(n_3589));
	notech_and4 i_2022(.A(n_3589), .B(n_3588), .C(n_3586), .D(n_3585), .Z(n_3591
		));
	notech_ao4 i_2041(.A(n_58630), .B(n_43095), .C(n_58746), .D(n_43080), .Z
		(n_3593));
	notech_ao4 i_2042(.A(n_58767), .B(n_43221), .C(n_58606), .D(n_43205), .Z
		(n_3595));
	notech_ao4 i_2043(.A(n_58725), .B(n_43111), .C(n_58441), .D(n_43237), .Z
		(n_359699552));
	notech_and4 i_2052(.A(n_359699552), .B(n_3595), .C(n_3593), .D(n_247498940
		), .Z(n_3598));
	notech_ao4 i_2044(.A(n_58887), .B(n_43064), .C(n_58788), .D(n_43253), .Z
		(n_3599));
	notech_ao4 i_2045(.A(n_58908), .B(n_43048), .C(n_58651), .D(n_43127), .Z
		(n_3600));
	notech_ao4 i_2046(.A(n_58868), .B(n_43143), .C(n_58930), .D(n_43037), .Z
		(n_360299553));
	notech_ao4 i_2047(.A(n_58849), .B(n_43158), .C(n_58959), .D(n_43190), .Z
		(n_3603));
	notech_and4 i_2053(.A(n_3603), .B(n_360299553), .C(n_3600), .D(n_3599), 
		.Z(n_3605));
	notech_ao4 i_2072(.A(n_58630), .B(n_43097), .C(n_58746), .D(n_43082), .Z
		(n_3607));
	notech_ao4 i_2073(.A(n_58767), .B(n_43223), .C(n_58607), .D(n_43207), .Z
		(n_3609));
	notech_ao4 i_2074(.A(n_58725), .B(n_43113), .C(n_58441), .D(n_43239), .Z
		(n_3610));
	notech_and4 i_2083(.A(n_3610), .B(n_3609), .C(n_3607), .D(n_249198957), 
		.Z(n_3612));
	notech_ao4 i_2075(.A(n_58887), .B(n_43066), .C(n_58788), .D(n_43255), .Z
		(n_3613));
	notech_ao4 i_2076(.A(n_58908), .B(n_43050), .C(n_58651), .D(n_43129), .Z
		(n_361499555));
	notech_ao4 i_2077(.A(n_58868), .B(n_43144), .C(n_58931), .D(n_43038), .Z
		(n_3616));
	notech_ao4 i_2078(.A(n_58849), .B(n_43160), .C(n_58959), .D(n_43192), .Z
		(n_3617));
	notech_and4 i_2084(.A(n_3617), .B(n_3616), .C(n_361499555), .D(n_3613), 
		.Z(n_3619));
	notech_ao4 i_2103(.A(n_58630), .B(n_43099), .C(n_58746), .D(n_43084), .Z
		(n_3621));
	notech_ao4 i_2104(.A(n_58767), .B(n_43225), .C(n_58607), .D(n_43209), .Z
		(n_3623));
	notech_ao4 i_2105(.A(n_58725), .B(n_43115), .C(n_58441), .D(n_43241), .Z
		(n_3624));
	notech_and4 i_2114(.A(n_3624), .B(n_3623), .C(n_3621), .D(n_250898974), 
		.Z(n_362699557));
	notech_ao4 i_2106(.A(n_58887), .B(n_43068), .C(n_58788), .D(n_43257), .Z
		(n_3627));
	notech_ao4 i_2107(.A(n_58908), .B(n_43052), .C(n_58651), .D(n_43131), .Z
		(n_3628));
	notech_ao4 i_2108(.A(n_58868), .B(n_43146), .C(n_58931), .D(n_43039), .Z
		(n_3630));
	notech_ao4 i_2109(.A(n_58849), .B(n_43162), .C(n_58959), .D(n_43194), .Z
		(n_3631));
	notech_and4 i_2115(.A(n_3631), .B(n_3630), .C(n_3628), .D(n_3627), .Z(n_3633
		));
	notech_ao4 i_2134(.A(n_58630), .B(n_43101), .C(n_58746), .D(n_43085), .Z
		(n_3635));
	notech_ao4 i_2135(.A(n_58767), .B(n_43227), .C(n_58607), .D(n_43211), .Z
		(n_3637));
	notech_ao4 i_2136(.A(n_58725), .B(n_43117), .C(n_58447), .D(n_43243), .Z
		(n_363899559));
	notech_and4 i_2145(.A(n_363899559), .B(n_3637), .C(n_3635), .D(n_252598991
		), .Z(n_3640));
	notech_ao4 i_2137(.A(n_58887), .B(n_43070), .C(n_58788), .D(n_43259), .Z
		(n_3641));
	notech_ao4 i_2138(.A(n_58908), .B(n_43054), .C(n_58651), .D(n_43133), .Z
		(n_3642));
	notech_ao4 i_2139(.A(n_58868), .B(n_43148), .C(n_58931), .D(n_43040), .Z
		(n_364499560));
	notech_ao4 i_2140(.A(n_58849), .B(n_43164), .C(n_58959), .D(n_43196), .Z
		(n_3645));
	notech_and4 i_2146(.A(n_3645), .B(n_364499560), .C(n_3642), .D(n_3641), 
		.Z(n_3647));
	notech_ao4 i_2165(.A(n_58630), .B(n_43103), .C(n_58746), .D(n_43087), .Z
		(n_3649));
	notech_ao4 i_2166(.A(n_58767), .B(n_43229), .C(n_58607), .D(n_43213), .Z
		(n_3651));
	notech_ao4 i_2167(.A(n_58725), .B(n_43119), .C(n_58445), .D(n_43245), .Z
		(n_3652));
	notech_and4 i_2176(.A(n_3652), .B(n_3651), .C(n_3649), .D(n_254299008), 
		.Z(n_3654));
	notech_ao4 i_2168(.A(n_58887), .B(n_43072), .C(n_58788), .D(n_43261), .Z
		(n_3655));
	notech_ao4 i_2169(.A(n_58908), .B(n_43056), .C(n_58651), .D(n_43135), .Z
		(n_365699562));
	notech_ao4 i_2170(.A(n_58868), .B(n_43150), .C(n_58931), .D(n_43041), .Z
		(n_3658));
	notech_ao4 i_2171(.A(n_58849), .B(n_43166), .C(n_58959), .D(n_43198), .Z
		(n_3659));
	notech_and4 i_2177(.A(n_3659), .B(n_3658), .C(n_365699562), .D(n_3655), 
		.Z(n_3661));
	notech_ao4 i_2196(.A(n_58630), .B(n_43105), .C(n_58746), .D(n_43089), .Z
		(n_3663));
	notech_ao4 i_2197(.A(n_58767), .B(n_43231), .C(n_58607), .D(n_43215), .Z
		(n_3665));
	notech_ao4 i_2198(.A(n_58725), .B(n_43121), .C(n_58445), .D(n_43247), .Z
		(n_3666));
	notech_and4 i_2207(.A(n_3666), .B(n_3665), .C(n_3663), .D(n_255999025), 
		.Z(n_366899564));
	notech_ao4 i_2199(.A(n_58890), .B(n_43074), .C(n_58788), .D(n_43263), .Z
		(n_3669));
	notech_ao4 i_2200(.A(n_58908), .B(n_43058), .C(n_58651), .D(n_43137), .Z
		(n_3670));
	notech_ao4 i_2201(.A(n_58871), .B(n_43152), .C(n_58931), .D(n_43042), .Z
		(n_3672));
	notech_ao4 i_2202(.A(n_58852), .B(n_43168), .C(n_58962), .D(n_43200), .Z
		(n_3673));
	notech_and4 i_2208(.A(n_3673), .B(n_3672), .C(n_3670), .D(n_3669), .Z(n_3676
		));
	notech_ao4 i_2227(.A(n_58630), .B(n_43107), .C(n_58746), .D(n_43091), .Z
		(n_3678));
	notech_ao4 i_2228(.A(n_58767), .B(n_43233), .C(n_58607), .D(n_43217), .Z
		(n_368099565));
	notech_ao4 i_2229(.A(n_58725), .B(n_43123), .C(n_58445), .D(n_43249), .Z
		(n_3681));
	notech_and4 i_2238(.A(n_3681), .B(n_368099565), .C(n_3678), .D(n_257699042
		), .Z(n_3683));
	notech_ao4 i_2230(.A(n_58890), .B(n_43076), .C(n_58788), .D(n_43265), .Z
		(n_3684));
	notech_ao4 i_2231(.A(n_58908), .B(n_43060), .C(n_58651), .D(n_43139), .Z
		(n_3685));
	notech_ao4 i_2232(.A(n_58871), .B(n_43154), .C(n_58931), .D(n_43044), .Z
		(n_3687));
	notech_ao4 i_2233(.A(n_58852), .B(n_43170), .C(n_58962), .D(n_43201), .Z
		(n_3688));
	notech_and4 i_2239(.A(n_3688), .B(n_3687), .C(n_3685), .D(n_3684), .Z(n_3690
		));
	notech_ao4 i_2258(.A(n_58630), .B(n_43109), .C(n_58746), .D(n_43093), .Z
		(n_369299567));
	notech_ao4 i_2259(.A(n_58767), .B(n_43235), .C(n_58607), .D(n_43219), .Z
		(n_3694));
	notech_ao4 i_2260(.A(n_58725), .B(n_43125), .C(n_58445), .D(n_43251), .Z
		(n_3695));
	notech_and4 i_2269(.A(n_3695), .B(n_3694), .C(n_369299567), .D(n_259399059
		), .Z(n_3697));
	notech_ao4 i_2261(.A(n_58890), .B(n_43078), .C(n_58788), .D(n_43267), .Z
		(n_369899568));
	notech_ao4 i_2262(.A(n_58908), .B(n_43062), .C(n_58651), .D(n_43141), .Z
		(n_3699));
	notech_ao4 i_2263(.A(n_58871), .B(n_43156), .C(n_58930), .D(n_43046), .Z
		(n_3701));
	notech_ao4 i_2264(.A(n_58852), .B(n_43172), .C(n_58962), .D(n_43203), .Z
		(n_3702));
	notech_and4 i_2270(.A(n_3702), .B(n_3701), .C(n_3699), .D(n_369899568), 
		.Z(n_370499569));
	notech_ao4 i_2289(.A(n_58630), .B(n_43111), .C(n_58746), .D(n_43095), .Z
		(n_3706));
	notech_ao4 i_2290(.A(n_58767), .B(n_43237), .C(n_58612), .D(n_43221), .Z
		(n_3708));
	notech_ao4 i_2291(.A(n_58725), .B(n_43127), .C(n_58447), .D(n_43253), .Z
		(n_3709));
	notech_and4 i_2300(.A(n_3709), .B(n_3708), .C(n_3706), .D(n_261099076), 
		.Z(n_3711));
	notech_ao4 i_2292(.A(n_58890), .B(n_43080), .C(n_58788), .D(n_43269), .Z
		(n_3712));
	notech_ao4 i_2293(.A(n_58908), .B(n_43064), .C(n_58651), .D(n_43143), .Z
		(n_3713));
	notech_ao4 i_2294(.A(n_58871), .B(n_43158), .C(n_58930), .D(n_43048), .Z
		(n_3715));
	notech_ao4 i_2295(.A(n_58852), .B(n_43174), .C(n_58962), .D(n_43205), .Z
		(n_371699571));
	notech_and4 i_2301(.A(n_371699571), .B(n_3715), .C(n_3713), .D(n_3712), 
		.Z(n_3718));
	notech_ao4 i_2320(.A(n_58630), .B(n_43113), .C(n_58746), .D(n_43097), .Z
		(n_3720));
	notech_ao4 i_2321(.A(n_58767), .B(n_43239), .C(n_58612), .D(n_43223), .Z
		(n_372299572));
	notech_ao4 i_2322(.A(n_58725), .B(n_43129), .C(n_58447), .D(n_43255), .Z
		(n_3723));
	notech_and4 i_2331(.A(n_3723), .B(n_372299572), .C(n_3720), .D(n_262799093
		), .Z(n_3725));
	notech_ao4 i_2323(.A(n_58890), .B(n_43082), .C(n_58788), .D(n_43271), .Z
		(n_3726));
	notech_ao4 i_2324(.A(n_58908), .B(n_43066), .C(n_58651), .D(n_43144), .Z
		(n_3727));
	notech_ao4 i_2325(.A(n_58871), .B(n_43160), .C(n_58930), .D(n_43050), .Z
		(n_3729));
	notech_ao4 i_2326(.A(n_58852), .B(n_43176), .C(n_58959), .D(n_43207), .Z
		(n_3730));
	notech_and4 i_2332(.A(n_3730), .B(n_3729), .C(n_3727), .D(n_3726), .Z(n_3732
		));
	notech_ao4 i_2351(.A(n_58630), .B(n_43115), .C(n_58746), .D(n_43099), .Z
		(n_373499574));
	notech_ao4 i_2352(.A(n_58767), .B(n_43241), .C(n_58612), .D(n_43225), .Z
		(n_3736));
	notech_ao4 i_2353(.A(n_58725), .B(n_43131), .C(n_58447), .D(n_43257), .Z
		(n_3737));
	notech_and4 i_2362(.A(n_3737), .B(n_3736), .C(n_373499574), .D(n_264499110
		), .Z(n_3739));
	notech_ao4 i_2354(.A(n_58890), .B(n_43084), .C(n_58788), .D(n_43273), .Z
		(n_374099575));
	notech_ao4 i_2355(.A(n_58908), .B(n_43068), .C(n_58651), .D(n_43146), .Z
		(n_3741));
	notech_ao4 i_2356(.A(n_58871), .B(n_43162), .C(n_58930), .D(n_43052), .Z
		(n_3743));
	notech_ao4 i_2357(.A(n_58852), .B(n_43178), .C(n_58959), .D(n_43209), .Z
		(n_3744));
	notech_and4 i_2363(.A(n_3744), .B(n_3743), .C(n_3741), .D(n_374099575), 
		.Z(n_374699576));
	notech_ao4 i_2382(.A(n_58630), .B(n_43117), .C(n_58746), .D(n_43101), .Z
		(n_3748));
	notech_ao4 i_2383(.A(n_58767), .B(n_43243), .C(n_58612), .D(n_43227), .Z
		(n_3750));
	notech_ao4 i_2384(.A(n_58725), .B(n_43133), .C(n_58447), .D(n_43259), .Z
		(n_3751));
	notech_and4 i_2393(.A(n_3751), .B(n_3750), .C(n_3748), .D(n_266199127), 
		.Z(n_3753));
	notech_ao4 i_2385(.A(n_58890), .B(n_43085), .C(n_58788), .D(n_43275), .Z
		(n_3754));
	notech_ao4 i_2386(.A(n_58908), .B(n_43070), .C(n_58651), .D(n_43148), .Z
		(n_3755));
	notech_ao4 i_2387(.A(n_58871), .B(n_43164), .C(n_58930), .D(n_43054), .Z
		(n_3757));
	notech_ao4 i_2388(.A(n_58852), .B(n_43180), .C(n_58962), .D(n_43211), .Z
		(n_375899578));
	notech_and4 i_2394(.A(n_375899578), .B(n_3757), .C(n_3755), .D(n_3754), 
		.Z(n_3760));
	notech_ao4 i_2413(.A(n_58630), .B(n_43119), .C(n_58746), .D(n_43103), .Z
		(n_3762));
	notech_ao4 i_2414(.A(n_58767), .B(n_43245), .C(n_58612), .D(n_43229), .Z
		(n_376499579));
	notech_ao4 i_2415(.A(n_58725), .B(n_43135), .C(n_58447), .D(n_43261), .Z
		(n_3765));
	notech_and4 i_2424(.A(n_3765), .B(n_376499579), .C(n_3762), .D(n_267899144
		), .Z(n_3767));
	notech_ao4 i_2416(.A(n_58890), .B(n_43087), .C(n_58788), .D(n_43277), .Z
		(n_3768));
	notech_ao4 i_2417(.A(n_58908), .B(n_43072), .C(n_58651), .D(n_43150), .Z
		(n_3769));
	notech_ao4 i_2418(.A(n_58871), .B(n_43166), .C(n_58930), .D(n_43056), .Z
		(n_3771));
	notech_ao4 i_2419(.A(n_58852), .B(n_43182), .C(n_58959), .D(n_43213), .Z
		(n_3772));
	notech_and4 i_2425(.A(n_3772), .B(n_3771), .C(n_3769), .D(n_3768), .Z(n_3774
		));
	notech_and2 i_76280076(.A(n_942), .B(n_134197811), .Z(n_377699581));
	notech_ao3 i_180480073(.A(n_134297812), .B(n_8130), .C(n_8137), .Z(n_3777
		));
	notech_and2 i_77380072(.A(n_942), .B(n_133997809), .Z(n_3778));
	notech_ao4 i_81280070(.A(n_376156298), .B(n_2950), .C(n_60790), .D(n_2946
		), .Z(n_3779));
	notech_ao4 i_81180069(.A(n_2951), .B(n_2950), .C(n_60793), .D(n_2946), .Z
		(n_3780));
	notech_ao4 i_20928597(.A(n_60633), .B(n_43433), .C(n_55140), .D(n_43609)
		, .Z(n_3781));
	notech_ao4 i_18028568(.A(n_60633), .B(n_43404), .C(n_55140), .D(n_43610)
		, .Z(n_378299582));
	notech_ao4 i_15028538(.A(n_60637), .B(n_43374), .C(n_55140), .D(n_43611)
		, .Z(n_3783));
	notech_nand2 i_8379352(.A(n_42914), .B(wptr[0]), .Z(n_376156298));
	notech_nao3 i_118878306(.A(n_58672), .B(queue[42]), .C(n_2923), .Z(n_1478
		));
	notech_and4 i_3425012(.A(n_2478), .B(n_2477), .C(n_2472), .D(n_2476), .Z
		(squeue_33100276));
	notech_nao3 i_116178324(.A(n_2046), .B(queue[129]), .C(n_58612), .Z(n_1475
		));
	notech_nao3 i_114178337(.A(n_58672), .B(queue[41]), .C(n_2923), .Z(n_1462
		));
	notech_and4 i_3325011(.A(n_2464), .B(n_2463), .C(n_2458), .D(n_2462), .Z
		(squeue_32100277));
	notech_nao3 i_111478355(.A(n_2046), .B(queue[128]), .C(n_58612), .Z(n_1459
		));
	notech_nao3 i_109578368(.A(n_58672), .B(queue[40]), .C(n_2923), .Z(n_1446
		));
	notech_and4 i_3225010(.A(n_2450), .B(n_2449), .C(n_2444), .D(n_2448), .Z
		(squeue_31100278));
	notech_and4 i_106878386(.A(n_2887), .B(n_2915), .C(n_2046), .D(queue[127
		]), .Z(n_1443));
	notech_or2 i_104878399(.A(n_58930), .B(n_42954), .Z(n_1430));
	notech_and4 i_3125009(.A(n_2436), .B(n_2435), .C(n_2430), .D(n_2434), .Z
		(squeue_30100279));
	notech_and4 i_102178417(.A(n_2887), .B(n_2915), .C(n_2046), .D(queue[126
		]), .Z(n_1427));
	notech_or2 i_100278430(.A(n_58930), .B(n_42953), .Z(n_1414));
	notech_and4 i_2925007(.A(n_2422), .B(n_2421), .C(n_2416), .D(n_2420), .Z
		(squeue_28100280));
	notech_nao3 i_97578448(.A(n_58837), .B(queue[124]), .C(n_58614), .Z(n_1411
		));
	notech_nao3 i_95578461(.A(n_58672), .B(queue[36]), .C(n_2923), .Z(n_1398
		));
	notech_and4 i_2825006(.A(n_240896491), .B(n_240796490), .C(n_2402100083)
		, .D(n_2406100079), .Z(squeue_27100281));
	notech_nao3 i_92878479(.A(n_58833), .B(queue[123]), .C(n_58614), .Z(n_1395
		));
	notech_nand3 i_4379793(.A(code_ack), .B(code_req), .C(n_8629), .Z(n_6899651
		));
	notech_and3 i_22279615(.A(n_141554120), .B(n_43489), .C(n_43481), .Z(n_24299825
		));
	notech_xor2 i_4179795(.A(addrshft[3]), .B(n_28656625), .Z(n_24799830));
	notech_and2 i_5411(.A(addr_0[0]), .B(n_43489), .Z(n_27499857));
	notech_and2 i_5413(.A(addr_0[1]), .B(n_43489), .Z(n_27599858));
	notech_and2 i_5414(.A(addr_0[2]), .B(n_43489), .Z(n_27699859));
	notech_and2 i_5415(.A(addr_0[3]), .B(n_43489), .Z(n_27799860));
	notech_and2 i_5434(.A(n_2340), .B(n_43352), .Z(n_27899861));
	notech_and2 i_5435(.A(n_2342), .B(n_43352), .Z(n_27999862));
	notech_and2 i_5436(.A(n_2344), .B(n_43352), .Z(n_28099863));
	notech_and2 i_5437(.A(n_2346), .B(n_43352), .Z(n_28199864));
	notech_and2 i_5438(.A(n_2348), .B(n_43352), .Z(n_28299865));
	notech_and2 i_5439(.A(n_2350), .B(n_43352), .Z(n_28399866));
	notech_and2 i_5440(.A(n_2352), .B(n_43352), .Z(n_28499867));
	notech_and2 i_5441(.A(n_2354), .B(n_43352), .Z(n_28599868));
	notech_and2 i_5442(.A(n_2356), .B(n_43352), .Z(n_28699869));
	notech_and2 i_5443(.A(n_2358), .B(n_43352), .Z(n_28799870));
	notech_and2 i_5444(.A(n_2360), .B(n_43352), .Z(n_28899871));
	notech_and2 i_5446(.A(n_62888), .B(n_6899651), .Z(codeWEN));
	notech_and2 i_374479828(.A(idata[0]), .B(n_62884), .Z(cacheD[0]));
	notech_and2 i_374379829(.A(idata[1]), .B(n_62876), .Z(cacheD[1]));
	notech_and2 i_374279830(.A(idata[2]), .B(n_62882), .Z(cacheD[2]));
	notech_and2 i_374179831(.A(idata[3]), .B(n_62884), .Z(cacheD[3]));
	notech_and2 i_374079832(.A(idata[4]), .B(n_62884), .Z(cacheD[4]));
	notech_and2 i_373979833(.A(idata[5]), .B(n_62876), .Z(cacheD[5]));
	notech_and2 i_373879834(.A(idata[6]), .B(n_62876), .Z(cacheD[6]));
	notech_and2 i_373779835(.A(idata[7]), .B(n_62876), .Z(cacheD[7]));
	notech_and2 i_373679836(.A(idata[8]), .B(n_62876), .Z(cacheD[8]));
	notech_and2 i_373579837(.A(idata[9]), .B(n_62876), .Z(cacheD[9]));
	notech_and2 i_373479838(.A(idata[10]), .B(n_62876), .Z(cacheD[10]));
	notech_and2 i_373379839(.A(idata[11]), .B(n_62876), .Z(cacheD[11]));
	notech_and2 i_373279840(.A(idata[12]), .B(n_62876), .Z(cacheD[12]));
	notech_and2 i_373179841(.A(idata[13]), .B(n_62882), .Z(cacheD[13]));
	notech_and2 i_373079842(.A(idata[14]), .B(n_62884), .Z(cacheD[14]));
	notech_and2 i_372979843(.A(idata[15]), .B(n_62884), .Z(cacheD[15]));
	notech_and2 i_372879844(.A(idata[16]), .B(n_62882), .Z(cacheD[16]));
	notech_and2 i_372779845(.A(idata[17]), .B(n_62884), .Z(cacheD[17]));
	notech_and2 i_372679846(.A(idata[18]), .B(n_62882), .Z(cacheD[18]));
	notech_and2 i_372579847(.A(idata[19]), .B(n_62882), .Z(cacheD[19]));
	notech_and2 i_372479848(.A(idata[20]), .B(n_62884), .Z(cacheD[20]));
	notech_and2 i_372379849(.A(idata[21]), .B(n_62888), .Z(cacheD[21]));
	notech_and2 i_372279850(.A(idata[22]), .B(n_62884), .Z(cacheD[22]));
	notech_and2 i_372179851(.A(idata[23]), .B(n_62884), .Z(cacheD[23]));
	notech_and2 i_372079852(.A(idata[24]), .B(n_62884), .Z(cacheD[24]));
	notech_and2 i_371979853(.A(idata[25]), .B(n_62884), .Z(cacheD[25]));
	notech_and2 i_371879854(.A(idata[26]), .B(n_62884), .Z(cacheD[26]));
	notech_and2 i_371779855(.A(idata[27]), .B(n_62884), .Z(cacheD[27]));
	notech_and2 i_371679856(.A(idata[28]), .B(n_62884), .Z(cacheD[28]));
	notech_and2 i_371579857(.A(idata[29]), .B(n_62884), .Z(cacheD[29]));
	notech_and2 i_371479858(.A(idata[30]), .B(n_62884), .Z(cacheD[30]));
	notech_and2 i_371379859(.A(idata[31]), .B(n_62884), .Z(cacheD[31]));
	notech_and2 i_371279860(.A(idata[32]), .B(n_62884), .Z(cacheD[32]));
	notech_and2 i_371179861(.A(idata[33]), .B(n_62888), .Z(cacheD[33]));
	notech_and2 i_371079862(.A(idata[34]), .B(n_62882), .Z(cacheD[34]));
	notech_and2 i_370979863(.A(idata[35]), .B(n_62882), .Z(cacheD[35]));
	notech_and2 i_370879864(.A(idata[36]), .B(n_62882), .Z(cacheD[36]));
	notech_and2 i_370779865(.A(idata[37]), .B(n_62882), .Z(cacheD[37]));
	notech_and2 i_370679866(.A(idata[38]), .B(n_62882), .Z(cacheD[38]));
	notech_and2 i_370579867(.A(idata[39]), .B(n_62882), .Z(cacheD[39]));
	notech_and2 i_370479868(.A(idata[40]), .B(n_62882), .Z(cacheD[40]));
	notech_and2 i_370379869(.A(idata[41]), .B(n_62882), .Z(cacheD[41]));
	notech_and2 i_370279870(.A(idata[42]), .B(n_62882), .Z(cacheD[42]));
	notech_and2 i_370179871(.A(idata[43]), .B(n_62888), .Z(cacheD[43]));
	notech_and2 i_370079872(.A(idata[44]), .B(n_62888), .Z(cacheD[44]));
	notech_and2 i_369979873(.A(idata[45]), .B(n_62888), .Z(cacheD[45]));
	notech_and2 i_369879874(.A(idata[46]), .B(n_62888), .Z(cacheD[46]));
	notech_and2 i_369779875(.A(idata[47]), .B(n_62888), .Z(cacheD[47]));
	notech_and2 i_369679876(.A(idata[48]), .B(n_62888), .Z(cacheD[48]));
	notech_and2 i_369579877(.A(idata[49]), .B(n_62888), .Z(cacheD[49]));
	notech_and2 i_369479878(.A(idata[50]), .B(n_62888), .Z(cacheD[50]));
	notech_and2 i_369379879(.A(idata[51]), .B(n_62888), .Z(cacheD[51]));
	notech_and2 i_369279880(.A(n_62888), .B(idata[52]), .Z(cacheD[52]));
	notech_and2 i_369179881(.A(idata[53]), .B(n_62882), .Z(cacheD[53]));
	notech_and2 i_369079882(.A(n_62888), .B(idata[54]), .Z(cacheD[54]));
	notech_and2 i_368979883(.A(n_62888), .B(idata[55]), .Z(cacheD[55]));
	notech_and2 i_368879884(.A(idata[56]), .B(n_62882), .Z(cacheD[56]));
	notech_and2 i_368779885(.A(n_62888), .B(idata[57]), .Z(cacheD[57]));
	notech_and2 i_368679886(.A(idata[58]), .B(n_62882), .Z(cacheD[58]));
	notech_and2 i_368579887(.A(idata[59]), .B(n_62882), .Z(cacheD[59]));
	notech_and2 i_368479888(.A(n_62888), .B(idata[60]), .Z(cacheD[60]));
	notech_and2 i_368379889(.A(idata[61]), .B(n_62882), .Z(cacheD[61]));
	notech_and2 i_368279890(.A(idata[62]), .B(n_62876), .Z(cacheD[62]));
	notech_and2 i_368179891(.A(idata[63]), .B(n_62876), .Z(cacheD[63]));
	notech_and2 i_368079892(.A(idata[64]), .B(n_62876), .Z(cacheD[64]));
	notech_and2 i_367979893(.A(idata[65]), .B(n_62876), .Z(cacheD[65]));
	notech_and2 i_367879894(.A(idata[66]), .B(n_62876), .Z(cacheD[66]));
	notech_and2 i_367779895(.A(idata[67]), .B(n_62876), .Z(cacheD[67]));
	notech_and2 i_367679896(.A(idata[68]), .B(n_62876), .Z(cacheD[68]));
	notech_and2 i_367579897(.A(idata[69]), .B(n_62876), .Z(cacheD[69]));
	notech_and2 i_367479898(.A(idata[70]), .B(n_62876), .Z(cacheD[70]));
	notech_and2 i_367379899(.A(idata[71]), .B(n_62884), .Z(cacheD[71]));
	notech_and2 i_367279900(.A(idata[72]), .B(n_62878), .Z(cacheD[72]));
	notech_and2 i_367179901(.A(idata[73]), .B(n_62878), .Z(cacheD[73]));
	notech_and2 i_367079902(.A(idata[74]), .B(n_62878), .Z(cacheD[74]));
	notech_and2 i_366979903(.A(idata[75]), .B(n_62878), .Z(cacheD[75]));
	notech_and2 i_366879904(.A(idata[76]), .B(n_62878), .Z(cacheD[76]));
	notech_and2 i_366779905(.A(idata[77]), .B(n_62878), .Z(cacheD[77]));
	notech_and2 i_366679906(.A(idata[78]), .B(n_62878), .Z(cacheD[78]));
	notech_and2 i_366579907(.A(idata[79]), .B(n_62878), .Z(cacheD[79]));
	notech_and2 i_366479908(.A(idata[80]), .B(n_62878), .Z(cacheD[80]));
	notech_and2 i_366379909(.A(idata[81]), .B(n_62878), .Z(cacheD[81]));
	notech_and2 i_366279910(.A(idata[82]), .B(n_62878), .Z(cacheD[82]));
	notech_and2 i_366179911(.A(idata[83]), .B(n_62878), .Z(cacheD[83]));
	notech_and2 i_366079912(.A(idata[84]), .B(n_62878), .Z(cacheD[84]));
	notech_and2 i_365979913(.A(idata[85]), .B(n_62878), .Z(cacheD[85]));
	notech_and2 i_365879914(.A(idata[86]), .B(n_62878), .Z(cacheD[86]));
	notech_and2 i_365779915(.A(idata[87]), .B(n_62878), .Z(cacheD[87]));
	notech_and2 i_365679916(.A(idata[88]), .B(n_62878), .Z(cacheD[88]));
	notech_and2 i_365579917(.A(idata[89]), .B(n_62878), .Z(cacheD[89]));
	notech_and2 i_365479918(.A(idata[90]), .B(n_62886), .Z(cacheD[90]));
	notech_and2 i_365379919(.A(idata[91]), .B(n_62886), .Z(cacheD[91]));
	notech_and2 i_365279920(.A(idata[92]), .B(n_62886), .Z(cacheD[92]));
	notech_and2 i_365179921(.A(idata[93]), .B(n_62886), .Z(cacheD[93]));
	notech_and2 i_365079922(.A(idata[94]), .B(n_62886), .Z(cacheD[94]));
	notech_and2 i_364979923(.A(idata[95]), .B(n_62886), .Z(cacheD[95]));
	notech_and2 i_364879924(.A(idata[96]), .B(n_62886), .Z(cacheD[96]));
	notech_and2 i_364779925(.A(idata[97]), .B(n_62886), .Z(cacheD[97]));
	notech_and2 i_364679926(.A(idata[98]), .B(n_62886), .Z(cacheD[98]));
	notech_and2 i_364579927(.A(idata[99]), .B(n_62886), .Z(cacheD[99]));
	notech_and2 i_364479928(.A(idata[100]), .B(n_62886), .Z(cacheD[100]));
	notech_and2 i_364379929(.A(idata[101]), .B(n_62886), .Z(cacheD[101]));
	notech_and2 i_364279930(.A(idata[102]), .B(n_62886), .Z(cacheD[102]));
	notech_and2 i_364179931(.A(idata[103]), .B(n_62886), .Z(cacheD[103]));
	notech_and2 i_364079932(.A(idata[104]), .B(n_62886), .Z(cacheD[104]));
	notech_and2 i_363979933(.A(idata[105]), .B(n_62886), .Z(cacheD[105]));
	notech_and2 i_363879934(.A(idata[106]), .B(n_62886), .Z(cacheD[106]));
	notech_and2 i_363779935(.A(idata[107]), .B(n_62886), .Z(cacheD[107]));
	notech_and2 i_363679936(.A(idata[108]), .B(n_62878), .Z(cacheD[108]));
	notech_and2 i_363579937(.A(idata[109]), .B(n_62886), .Z(cacheD[109]));
	notech_and2 i_363479938(.A(idata[110]), .B(n_62880), .Z(cacheD[110]));
	notech_and2 i_363379939(.A(idata[111]), .B(n_62880), .Z(cacheD[111]));
	notech_and2 i_363279940(.A(idata[112]), .B(n_62880), .Z(cacheD[112]));
	notech_and2 i_363179941(.A(idata[113]), .B(n_62880), .Z(cacheD[113]));
	notech_and2 i_363079942(.A(idata[114]), .B(n_62880), .Z(cacheD[114]));
	notech_and2 i_362979943(.A(idata[115]), .B(n_62880), .Z(cacheD[115]));
	notech_and2 i_362879944(.A(idata[116]), .B(n_62880), .Z(cacheD[116]));
	notech_and2 i_362779945(.A(idata[117]), .B(n_62880), .Z(cacheD[117]));
	notech_and2 i_362679946(.A(idata[118]), .B(n_62880), .Z(cacheD[118]));
	notech_and2 i_362579947(.A(idata[119]), .B(n_62880), .Z(cacheD[119]));
	notech_and2 i_362479948(.A(idata[120]), .B(n_62880), .Z(cacheD[120]));
	notech_and2 i_362379949(.A(idata[121]), .B(n_62880), .Z(cacheD[121]));
	notech_and2 i_362279950(.A(idata[122]), .B(n_62880), .Z(cacheD[122]));
	notech_and2 i_362179951(.A(idata[123]), .B(n_62880), .Z(cacheD[123]));
	notech_and2 i_362079952(.A(idata[124]), .B(n_62880), .Z(cacheD[124]));
	notech_and2 i_361979953(.A(idata[125]), .B(n_62880), .Z(cacheD[125]));
	notech_and2 i_361879954(.A(idata[126]), .B(n_62880), .Z(cacheD[126]));
	notech_and2 i_361779955(.A(idata[127]), .B(n_62880), .Z(cacheD[127]));
	notech_and2 i_361679956(.A(iaddr[14]), .B(n_62880), .Z(cacheD[128]));
	notech_and2 i_361579957(.A(iaddr[15]), .B(cacheD[148]), .Z(cacheD[129])
		);
	notech_and2 i_361479958(.A(iaddr[16]), .B(cacheD[148]), .Z(cacheD[130])
		);
	notech_and2 i_361379959(.A(iaddr[17]), .B(cacheD[148]), .Z(cacheD[131])
		);
	notech_and2 i_361279960(.A(iaddr[18]), .B(cacheD[148]), .Z(cacheD[132])
		);
	notech_and2 i_361179961(.A(iaddr[19]), .B(cacheD[148]), .Z(cacheD[133])
		);
	notech_and2 i_361079962(.A(iaddr[20]), .B(cacheD[148]), .Z(cacheD[134])
		);
	notech_and2 i_360979963(.A(iaddr[21]), .B(cacheD[148]), .Z(cacheD[135])
		);
	notech_and2 i_360879964(.A(iaddr[22]), .B(cacheD[148]), .Z(cacheD[136])
		);
	notech_and2 i_360779965(.A(iaddr[23]), .B(cacheD[148]), .Z(cacheD[137])
		);
	notech_and2 i_360679966(.A(iaddr[24]), .B(cacheD[148]), .Z(cacheD[138])
		);
	notech_and2 i_360579967(.A(iaddr[25]), .B(cacheD[148]), .Z(cacheD[139])
		);
	notech_and2 i_360479968(.A(iaddr[26]), .B(cacheD[148]), .Z(cacheD[140])
		);
	notech_and2 i_360379969(.A(iaddr[27]), .B(cacheD[148]), .Z(cacheD[141])
		);
	notech_and2 i_360279970(.A(iaddr[28]), .B(cacheD[148]), .Z(cacheD[142])
		);
	notech_and2 i_360179971(.A(iaddr[29]), .B(cacheD[148]), .Z(cacheD[143])
		);
	notech_and2 i_360079972(.A(iaddr[30]), .B(cacheD[148]), .Z(cacheD[144])
		);
	notech_and2 i_359979973(.A(iaddr[31]), .B(cacheD[148]), .Z(cacheD[145])
		);
	notech_mux2 i_327168(.S(n_60754), .A(nbus_81[2]), .B(pc_in[2]), .Z(n_4657
		));
	notech_ao4 i_222659(.A(n_487100070), .B(n_488100071), .C(n_2947), .D(n_42914
		), .Z(n_2736));
	notech_mux2 i_1179315(.S(n_60754), .A(addr_0[10]), .B(pc_in[10]), .Z(n_4391
		));
	notech_ao4 i_22928617(.A(n_60637), .B(n_43453), .C(n_55140), .D(n_43517)
		, .Z(n_4148));
	notech_ao4 i_22628614(.A(n_60637), .B(n_43450), .C(n_55140), .D(n_43520)
		, .Z(n_4130));
	notech_ao4 i_22128609(.A(n_60637), .B(n_43445), .C(n_55140), .D(n_43525)
		, .Z(n_4100));
	notech_ao4 i_22028608(.A(n_60581), .B(n_43444), .C(n_55140), .D(n_43526)
		, .Z(n_4094));
	notech_ao4 i_21828606(.A(n_60581), .B(n_43442), .C(n_55140), .D(n_43528)
		, .Z(n_4082));
	notech_ao4 i_21728605(.A(n_60581), .B(n_43441), .C(n_55140), .D(n_43529)
		, .Z(n_4076));
	notech_ao4 i_21628604(.A(n_60581), .B(n_43440), .C(n_55140), .D(n_43530)
		, .Z(n_4070));
	notech_ao4 i_21528603(.A(n_60581), .B(n_43439), .C(n_55140), .D(n_43531)
		, .Z(n_4064));
	notech_ao4 i_21428602(.A(n_60581), .B(n_43438), .C(n_55140), .D(n_43532)
		, .Z(n_4058));
	notech_ao4 i_21328601(.A(n_60581), .B(n_43437), .C(n_55140), .D(n_43533)
		, .Z(n_4052));
	notech_ao4 i_21228600(.A(n_60581), .B(n_43436), .C(n_55140), .D(n_43534)
		, .Z(n_4046));
	notech_ao4 i_21128599(.A(n_60577), .B(n_43435), .C(n_55140), .D(n_43535)
		, .Z(n_4040));
	notech_ao4 i_21028598(.A(n_60577), .B(n_43434), .C(n_55140), .D(n_43536)
		, .Z(n_4034));
	notech_and2 i_3779351(.A(n_60793), .B(n_140854113), .Z(n_8165));
	notech_ao4 i_14928537(.A(n_60577), .B(n_43373), .C(n_55138), .D(n_43588)
		, .Z(n_3668));
	notech_nand2 i_222877332(.A(\queue_0[60] ), .B(n_60413), .Z(n_472100055)
		);
	notech_nand2 i_6128449(.A(n_489100072), .B(n_472100055), .Z(n_3140));
	notech_nand2 i_224077320(.A(\queue_0[57] ), .B(n_60413), .Z(n_474100057)
		);
	notech_nand2 i_5828446(.A(n_490100073), .B(n_474100057), .Z(n_3122));
	notech_nand2 i_224877312(.A(\queue_0[55] ), .B(n_60413), .Z(n_476100059)
		);
	notech_nand2 i_5628444(.A(n_491100074), .B(n_476100059), .Z(n_3110));
	notech_nand2 i_225277308(.A(\queue_0[54] ), .B(n_60413), .Z(n_478100061)
		);
	notech_nand2 i_5528443(.A(n_492100075), .B(n_478100061), .Z(n_3104));
	notech_nand2 i_226077300(.A(\queue_0[52] ), .B(n_60413), .Z(n_480100063)
		);
	notech_nand2 i_5328441(.A(n_493100076), .B(n_480100063), .Z(n_3092));
	notech_nand2 i_1979295(.A(n_43489), .B(n_2947), .Z(n_487100070));
	notech_nand2 i_189077670(.A(fault_wptr[1]), .B(fault_wptr[0]), .Z(n_488100071
		));
	notech_ao4 i_223077330(.A(n_60577), .B(n_43413), .C(n_60793), .D(n_43162
		), .Z(n_489100072));
	notech_ao4 i_224277318(.A(n_60581), .B(n_43410), .C(n_60793), .D(n_43156
		), .Z(n_490100073));
	notech_ao4 i_225077310(.A(n_60581), .B(n_43408), .C(n_60790), .D(n_43152
		), .Z(n_491100074));
	notech_ao4 i_225477306(.A(n_60577), .B(n_43407), .C(n_60790), .D(n_43150
		), .Z(n_492100075));
	notech_ao4 i_226277298(.A(n_60581), .B(n_43405), .C(n_60793), .D(n_43146
		), .Z(n_493100076));
	notech_ao4 i_78380075(.A(n_2033), .B(n_43489), .C(n_2993), .D(n_2995), .Z
		(n_2743));
	notech_mux2 i_180068(.S(purge), .A(iaddr[4]), .B(purge_cnt[0]), .Z(cacheA
		[0]));
	notech_mux2 i_211494(.S(purge), .A(iaddr[5]), .B(purge_cnt[1]), .Z(cacheA
		[1]));
	notech_mux2 i_380067(.S(purge), .A(iaddr[6]), .B(purge_cnt[2]), .Z(cacheA
		[2]));
	notech_mux2 i_480066(.S(purge), .A(iaddr[7]), .B(purge_cnt[3]), .Z(cacheA
		[3]));
	notech_mux2 i_511495(.S(purge), .A(iaddr[8]), .B(purge_cnt[4]), .Z(cacheA
		[4]));
	notech_mux2 i_680065(.S(purge), .A(iaddr[9]), .B(purge_cnt[5]), .Z(cacheA
		[5]));
	notech_mux2 i_780064(.S(purge), .A(iaddr[10]), .B(purge_cnt[6]), .Z(cacheA
		[6]));
	notech_mux2 i_880063(.S(purge), .A(iaddr[11]), .B(purge_cnt[7]), .Z(cacheA
		[7]));
	notech_mux2 i_980062(.S(purge), .A(iaddr[12]), .B(purge_cnt[8]), .Z(cacheA
		[8]));
	notech_mux2 i_1080061(.S(purge), .A(iaddr[13]), .B(purge_cnt[9]), .Z(cacheA
		[9]));
	notech_mux2 i_127154(.S(addrshft[0]), .A(n_2945), .B(n_948), .Z(valid_len_0100253
		));
	notech_ao4 i_427157(.A(addrshft[3]), .B(n_2945), .C(n_948), .D(n_24799830
		), .Z(valid_len_3100252));
	notech_nor2 i_527158(.A(n_28356622), .B(addrshft[4]), .Z(valid_len[4])
		);
	notech_mux2 i_427169(.S(n_60754), .A(nbus_81[3]), .B(pc_in[3]), .Z(n_4663
		));
	notech_mux2 i_227167(.S(n_60754), .A(nbus_81[1]), .B(pc_in[1]), .Z(n_4651
		));
	notech_mux2 i_127166(.S(n_60754), .A(nbus_81[0]), .B(pc_in[0]), .Z(n_4645
		));
	notech_ao4 i_122658(.A(fault_wptr[0]), .B(n_487100070), .C(n_2947), .D(n_42913
		), .Z(n_2730));
	notech_mux2 i_3279826(.S(n_60754), .A(addr_0[31]), .B(pc_in[31]), .Z(n_4517
		));
	notech_mux2 i_3179825(.S(n_60754), .A(addr_0[30]), .B(pc_in[30]), .Z(n_4511
		));
	notech_mux2 i_3079824(.S(n_60754), .A(addr_0[29]), .B(pc_in[29]), .Z(n_4505
		));
	notech_mux2 i_2979823(.S(n_60754), .A(addr_0[28]), .B(pc_in[28]), .Z(n_4499
		));
	notech_mux2 i_2879822(.S(n_60754), .A(addr_0[27]), .B(pc_in[27]), .Z(n_4493
		));
	notech_mux2 i_2779821(.S(n_60754), .A(addr_0[26]), .B(pc_in[26]), .Z(n_4487
		));
	notech_mux2 i_2679820(.S(n_60754), .A(addr_0[25]), .B(pc_in[25]), .Z(n_4481
		));
	notech_mux2 i_2579819(.S(n_60754), .A(addr_0[24]), .B(pc_in[24]), .Z(n_4475
		));
	notech_mux2 i_2479818(.S(n_60754), .A(addr_0[23]), .B(pc_in[23]), .Z(n_4469
		));
	notech_mux2 i_2379817(.S(n_60754), .A(addr_0[22]), .B(pc_in[22]), .Z(n_4463
		));
	notech_mux2 i_2279816(.S(n_60754), .A(addr_0[21]), .B(pc_in[21]), .Z(n_4457
		));
	notech_mux2 i_2179815(.S(n_60754), .A(addr_0[20]), .B(pc_in[20]), .Z(n_4451
		));
	notech_mux2 i_2079814(.S(n_60750), .A(addr_0[19]), .B(pc_in[19]), .Z(n_4445
		));
	notech_mux2 i_1979813(.S(n_60750), .A(addr_0[18]), .B(pc_in[18]), .Z(n_4439
		));
	notech_mux2 i_1879812(.S(n_60750), .A(addr_0[17]), .B(pc_in[17]), .Z(n_4433
		));
	notech_mux2 i_1779811(.S(n_60750), .A(addr_0[16]), .B(pc_in[16]), .Z(n_4427
		));
	notech_mux2 i_1679810(.S(n_60750), .A(addr_0[15]), .B(pc_in[15]), .Z(n_4421
		));
	notech_mux2 i_1579809(.S(n_60750), .A(addr_0[14]), .B(pc_in[14]), .Z(n_4415
		));
	notech_mux2 i_1479808(.S(n_60750), .A(addr_0[13]), .B(pc_in[13]), .Z(n_4409
		));
	notech_mux2 i_1379807(.S(n_60750), .A(addr_0[12]), .B(pc_in[12]), .Z(n_4403
		));
	notech_mux2 i_1279806(.S(n_60750), .A(addr_0[11]), .B(pc_in[11]), .Z(n_4397
		));
	notech_mux2 i_1011669(.S(n_60750), .A(addr_0[9]), .B(pc_in[9]), .Z(n_4385
		));
	notech_mux2 i_911668(.S(n_60750), .A(addr_0[8]), .B(pc_in[8]), .Z(n_4379
		));
	notech_mux2 i_811667(.S(n_60750), .A(addr_0[7]), .B(pc_in[7]), .Z(n_4373
		));
	notech_mux2 i_711666(.S(n_60750), .A(addr_0[6]), .B(pc_in[6]), .Z(n_4367
		));
	notech_mux2 i_611665(.S(n_60750), .A(addr_0[5]), .B(pc_in[5]), .Z(n_4361
		));
	notech_mux2 i_511664(.S(n_60750), .A(addr_0[4]), .B(pc_in[4]), .Z(n_4355
		));
	notech_ao4 i_25628644(.A(n_55138), .B(n_43490), .C(n_60586), .D(n_43480)
		, .Z(n_4310));
	notech_ao4 i_25528643(.A(n_55138), .B(n_43491), .C(n_60586), .D(n_43479)
		, .Z(n_4304));
	notech_ao4 i_25428642(.A(n_55138), .B(n_43492), .C(n_60586), .D(n_43478)
		, .Z(n_4298));
	notech_ao4 i_25328641(.A(n_55138), .B(n_43493), .C(n_60586), .D(n_43477)
		, .Z(n_4292));
	notech_ao4 i_25228640(.A(n_55138), .B(n_43494), .C(n_60586), .D(n_43476)
		, .Z(n_4286));
	notech_ao4 i_25128639(.A(n_55138), .B(n_43495), .C(n_60586), .D(n_43475)
		, .Z(n_4280));
	notech_ao4 i_25028638(.A(n_55138), .B(n_43496), .C(n_60586), .D(n_43474)
		, .Z(n_4274));
	notech_ao4 i_24928637(.A(n_55138), .B(n_43497), .C(n_60586), .D(n_43473)
		, .Z(n_4268));
	notech_ao4 i_24828636(.A(n_55138), .B(n_43498), .C(n_60586), .D(n_43472)
		, .Z(n_4262));
	notech_ao4 i_24728635(.A(n_55138), .B(n_43499), .C(n_60586), .D(n_43471)
		, .Z(n_4256));
	notech_ao4 i_24628634(.A(n_55138), .B(n_43500), .C(n_60581), .D(n_43470)
		, .Z(n_4250));
	notech_ao4 i_24528633(.A(n_55138), .B(n_43501), .C(n_60586), .D(n_43469)
		, .Z(n_4244));
	notech_ao4 i_24428632(.A(n_55138), .B(n_43502), .C(n_60586), .D(n_43468)
		, .Z(n_4238));
	notech_ao4 i_24328631(.A(n_55138), .B(n_43503), .C(n_60586), .D(n_43467)
		, .Z(n_4232));
	notech_ao4 i_24228630(.A(n_55138), .B(n_43504), .C(n_60586), .D(n_43466)
		, .Z(n_4226));
	notech_ao4 i_24128629(.A(n_55145), .B(n_43505), .C(n_60586), .D(n_43465)
		, .Z(n_4220));
	notech_ao4 i_24028628(.A(n_55145), .B(n_43506), .C(n_60568), .D(n_43464)
		, .Z(n_4214));
	notech_ao4 i_23928627(.A(n_55145), .B(n_43507), .C(n_60568), .D(n_43463)
		, .Z(n_4208));
	notech_ao4 i_23828626(.A(n_55145), .B(n_43508), .C(n_60568), .D(n_43462)
		, .Z(n_4202));
	notech_ao4 i_23728625(.A(n_55145), .B(n_43509), .C(n_60568), .D(n_43461)
		, .Z(n_4196));
	notech_ao4 i_23628624(.A(n_55145), .B(n_43510), .C(n_60572), .D(n_43460)
		, .Z(n_4190));
	notech_ao4 i_23528623(.A(n_55145), .B(n_43511), .C(n_60572), .D(n_43459)
		, .Z(n_4184));
	notech_ao4 i_23428622(.A(n_55145), .B(n_43512), .C(n_60568), .D(n_43458)
		, .Z(n_4178));
	notech_ao4 i_23328621(.A(n_55145), .B(n_43513), .C(n_60572), .D(n_43457)
		, .Z(n_4172));
	notech_ao4 i_23228620(.A(n_55145), .B(n_43514), .C(n_60568), .D(n_43456)
		, .Z(n_4166));
	notech_ao4 i_23128619(.A(n_55145), .B(n_43515), .C(n_60568), .D(n_43455)
		, .Z(n_4160));
	notech_ao4 i_23028618(.A(n_55145), .B(n_43516), .C(n_60568), .D(n_43454)
		, .Z(n_4154));
	notech_ao4 i_22828616(.A(n_60568), .B(n_43452), .C(n_55145), .D(n_43518)
		, .Z(n_4142));
	notech_ao4 i_22728615(.A(n_60568), .B(n_43451), .C(n_55145), .D(n_43519)
		, .Z(n_4136));
	notech_ao4 i_22528613(.A(n_60568), .B(n_43449), .C(n_55145), .D(n_43521)
		, .Z(n_4124));
	notech_ao4 i_22428612(.A(n_60568), .B(n_43448), .C(n_55145), .D(n_43522)
		, .Z(n_4118));
	notech_ao4 i_22328611(.A(n_60568), .B(n_43447), .C(n_55143), .D(n_43523)
		, .Z(n_4112));
	notech_ao4 i_22228610(.A(n_60577), .B(n_43446), .C(n_55143), .D(n_43524)
		, .Z(n_4106));
	notech_ao4 i_21928607(.A(n_60577), .B(n_43443), .C(n_55143), .D(n_43527)
		, .Z(n_4088));
	notech_ao4 i_20828596(.A(n_60572), .B(n_43432), .C(n_55143), .D(n_43537)
		, .Z(n_4022));
	notech_ao4 i_20728595(.A(n_60577), .B(n_43431), .C(n_55143), .D(n_43538)
		, .Z(n_4016));
	notech_ao4 i_20628594(.A(n_60577), .B(n_43430), .C(n_55143), .D(n_43539)
		, .Z(n_4010));
	notech_ao4 i_20528593(.A(n_60577), .B(n_43429), .C(n_55143), .D(n_43540)
		, .Z(n_4004));
	notech_ao4 i_20428592(.A(n_60577), .B(n_43428), .C(n_55143), .D(n_43541)
		, .Z(n_3998));
	notech_ao4 i_20328591(.A(n_60577), .B(n_43427), .C(n_55143), .D(n_43542)
		, .Z(n_3992));
	notech_ao4 i_20228590(.A(n_60572), .B(n_43426), .C(n_55143), .D(n_43543)
		, .Z(n_3986));
	notech_ao4 i_20128589(.A(n_60572), .B(n_43425), .C(n_55143), .D(n_43544)
		, .Z(n_3980));
	notech_ao4 i_20028588(.A(n_60572), .B(n_43424), .C(n_55143), .D(n_43545)
		, .Z(n_3974));
	notech_ao4 i_19928587(.A(n_60572), .B(n_43423), .C(n_55143), .D(n_43546)
		, .Z(n_3968));
	notech_ao4 i_19828586(.A(n_60572), .B(n_43422), .C(n_55143), .D(n_43547)
		, .Z(n_3962));
	notech_ao4 i_19728585(.A(n_60572), .B(n_43421), .C(n_55143), .D(n_43548)
		, .Z(n_3956));
	notech_ao4 i_19628584(.A(n_60572), .B(n_43420), .C(n_55143), .D(n_43549)
		, .Z(n_3950));
	notech_ao4 i_19528583(.A(n_60572), .B(n_43419), .C(n_55130), .D(n_43550)
		, .Z(n_3944));
	notech_ao4 i_19428582(.A(n_60566), .B(n_43418), .C(n_55130), .D(n_43551)
		, .Z(n_3938));
	notech_ao4 i_19328581(.A(n_60600), .B(n_43417), .C(n_55130), .D(n_43552)
		, .Z(n_3932));
	notech_ao4 i_19228580(.A(n_60605), .B(n_43416), .C(n_55130), .D(n_43553)
		, .Z(n_3926));
	notech_ao4 i_19128579(.A(n_60600), .B(n_43415), .C(n_55130), .D(n_43554)
		, .Z(n_3920));
	notech_ao4 i_19028578(.A(n_60600), .B(n_43414), .C(n_55130), .D(n_43555)
		, .Z(n_3914));
	notech_ao4 i_18928577(.A(n_60605), .B(n_43413), .C(n_55130), .D(n_43617)
		, .Z(n_3908));
	notech_ao4 i_18828576(.A(n_60605), .B(n_43412), .C(n_55130), .D(n_43556)
		, .Z(n_3902));
	notech_ao4 i_18728575(.A(n_60605), .B(n_43411), .C(n_55130), .D(n_43557)
		, .Z(n_3896));
	notech_ao4 i_18628574(.A(n_60605), .B(n_43410), .C(n_55130), .D(n_43616)
		, .Z(n_3890));
	notech_ao4 i_18528573(.A(n_60600), .B(n_43409), .C(n_55130), .D(n_43558)
		, .Z(n_3884));
	notech_ao4 i_18428572(.A(n_60600), .B(n_43408), .C(n_55130), .D(n_43615)
		, .Z(n_3878));
	notech_ao4 i_18328571(.A(n_60600), .B(n_43407), .C(n_55130), .D(n_43614)
		, .Z(n_3872));
	notech_ao4 i_18228570(.A(n_55130), .B(n_43612), .C(n_60600), .D(n_43406)
		, .Z(n_3866));
	notech_ao4 i_18128569(.A(n_60600), .B(n_43405), .C(n_55130), .D(n_43613)
		, .Z(n_3860));
	notech_ao4 i_17928567(.A(n_60600), .B(n_43403), .C(n_55130), .D(n_43559)
		, .Z(n_3848));
	notech_ao4 i_17828566(.A(n_60600), .B(n_43402), .C(n_55128), .D(n_43560)
		, .Z(n_3842));
	notech_ao4 i_17728565(.A(n_60600), .B(n_43401), .C(n_55128), .D(n_43561)
		, .Z(n_3836));
	notech_ao4 i_17628564(.A(n_60609), .B(n_43400), .C(n_55128), .D(n_43562)
		, .Z(n_3830));
	notech_ao4 i_17528563(.A(n_60609), .B(n_43399), .C(n_55128), .D(n_43563)
		, .Z(n_3824));
	notech_ao4 i_17428562(.A(n_60605), .B(n_43398), .C(n_55128), .D(n_43564)
		, .Z(n_3818));
	notech_ao4 i_17328561(.A(n_60605), .B(n_43397), .C(n_55128), .D(n_43565)
		, .Z(n_3812));
	notech_ao4 i_17228560(.A(n_60609), .B(n_43396), .C(n_55128), .D(n_43566)
		, .Z(n_3806));
	notech_ao4 i_17128559(.A(n_60609), .B(n_43395), .C(n_55128), .D(n_43567)
		, .Z(n_3800));
	notech_ao4 i_17028558(.A(n_60609), .B(n_43394), .C(n_55128), .D(n_43568)
		, .Z(n_3794));
	notech_ao4 i_16928557(.A(n_60609), .B(n_43393), .C(n_55128), .D(n_43569)
		, .Z(n_3788));
	notech_ao4 i_16828556(.A(n_60605), .B(n_43392), .C(n_55128), .D(n_43570)
		, .Z(n_3782));
	notech_ao4 i_16728555(.A(n_60605), .B(n_43391), .C(n_55128), .D(n_43571)
		, .Z(n_3776));
	notech_ao4 i_16628554(.A(n_60605), .B(n_43390), .C(n_55128), .D(n_43572)
		, .Z(n_3770));
	notech_ao4 i_16528553(.A(n_60605), .B(n_43389), .C(n_55128), .D(n_43573)
		, .Z(n_3764));
	notech_ao4 i_16428552(.A(n_60605), .B(n_43388), .C(n_55128), .D(n_43574)
		, .Z(n_3758));
	notech_ao4 i_16328551(.A(n_60605), .B(n_43387), .C(n_55128), .D(n_43575)
		, .Z(n_3752));
	notech_ao4 i_16228550(.A(n_60605), .B(n_43386), .C(n_55135), .D(n_43576)
		, .Z(n_3746));
	notech_ao4 i_16128549(.A(n_60605), .B(n_43385), .C(n_55135), .D(n_43577)
		, .Z(n_3740));
	notech_ao4 i_16028548(.A(n_60566), .B(n_43384), .C(n_55135), .D(n_43578)
		, .Z(n_3734));
	notech_ao4 i_15928547(.A(n_60566), .B(n_43383), .C(n_55135), .D(n_43579)
		, .Z(n_3728));
	notech_ao4 i_15828546(.A(n_60566), .B(n_43382), .C(n_55135), .D(n_43580)
		, .Z(n_3722));
	notech_ao4 i_15728545(.A(n_60566), .B(n_43381), .C(n_55135), .D(n_43581)
		, .Z(n_3716));
	notech_ao4 i_15628544(.A(n_60596), .B(n_43380), .C(n_55135), .D(n_43582)
		, .Z(n_3710));
	notech_ao4 i_15528543(.A(n_60596), .B(n_43379), .C(n_55135), .D(n_43583)
		, .Z(n_3704));
	notech_ao4 i_15428542(.A(n_60566), .B(n_43378), .C(n_55135), .D(n_43584)
		, .Z(n_3698));
	notech_ao4 i_15328541(.A(n_60596), .B(n_43377), .C(n_55135), .D(n_43585)
		, .Z(n_3692));
	notech_ao4 i_15228540(.A(n_60566), .B(n_43376), .C(n_55135), .D(n_43586)
		, .Z(n_3686));
	notech_ao4 i_15128539(.A(n_60566), .B(n_43375), .C(n_55135), .D(n_43587)
		, .Z(n_3680));
	notech_ao4 i_14828536(.A(n_60566), .B(n_43372), .C(n_55135), .D(n_43589)
		, .Z(n_3662));
	notech_ao4 i_14728535(.A(n_60566), .B(n_43371), .C(n_55135), .D(n_43590)
		, .Z(n_3656));
	notech_ao4 i_14628534(.A(n_60566), .B(n_43370), .C(n_55135), .D(n_43591)
		, .Z(n_3650));
	notech_ao4 i_14528533(.A(n_60566), .B(n_43369), .C(n_55135), .D(n_43592)
		, .Z(n_3644));
	notech_ao4 i_14428532(.A(n_60566), .B(n_43368), .C(n_55133), .D(n_43593)
		, .Z(n_3638));
	notech_ao4 i_14328531(.A(n_60566), .B(n_43367), .C(n_55133), .D(n_43594)
		, .Z(n_3632));
	notech_ao4 i_14228530(.A(n_60596), .B(n_43366), .C(n_55133), .D(n_43595)
		, .Z(n_3626));
	notech_ao4 i_14128529(.A(n_60596), .B(n_43365), .C(n_55133), .D(n_43596)
		, .Z(n_3620));
	notech_ao4 i_14028528(.A(n_60596), .B(n_43364), .C(n_55133), .D(n_43597)
		, .Z(n_3614));
	notech_ao4 i_13928527(.A(n_60596), .B(n_43363), .C(n_55133), .D(n_43598)
		, .Z(n_3608));
	notech_ao4 i_13828526(.A(n_60600), .B(n_43362), .C(n_55133), .D(n_43599)
		, .Z(n_3602));
	notech_ao4 i_13728525(.A(n_55133), .B(n_43600), .C(n_60600), .D(n_43361)
		, .Z(n_3596));
	notech_ao4 i_13628524(.A(n_60600), .B(n_43360), .C(n_55133), .D(n_43601)
		, .Z(n_3590));
	notech_ao4 i_13528523(.A(n_60600), .B(n_43359), .C(n_55133), .D(n_43602)
		, .Z(n_3584));
	notech_ao4 i_13428522(.A(n_60596), .B(n_43358), .C(n_55133), .D(n_43603)
		, .Z(n_3578));
	notech_ao4 i_13328521(.A(n_60596), .B(n_43357), .C(n_55133), .D(n_43604)
		, .Z(n_3572));
	notech_ao4 i_13228520(.A(n_60596), .B(n_43356), .C(n_55133), .D(n_43605)
		, .Z(n_3566));
	notech_ao4 i_13128519(.A(n_60596), .B(n_43355), .C(n_55133), .D(n_43606)
		, .Z(n_3560));
	notech_ao4 i_13028518(.A(n_60596), .B(n_43354), .C(n_55133), .D(n_43607)
		, .Z(n_3554));
	notech_ao4 i_12928517(.A(n_60596), .B(n_43353), .C(n_55133), .D(n_43608)
		, .Z(n_3548));
	notech_nao3 i_90978492(.A(n_58672), .B(queue[35]), .C(n_2923), .Z(n_1382
		));
	notech_and4 i_2725005(.A(n_2393100091), .B(n_2392100092), .C(n_2387), .D
		(n_2391100093), .Z(squeue_26100282));
	notech_nao3 i_88278510(.A(n_58833), .B(queue[122]), .C(n_58614), .Z(n_1379
		));
	notech_nao3 i_86278523(.A(n_58672), .B(queue[34]), .C(n_58943), .Z(n_1366
		));
	notech_and4 i_2625004(.A(n_2379100102), .B(n_2378100103), .C(n_2373100107
		), .D(n_2377100104), .Z(squeue_25100283));
	notech_nao3 i_83578541(.A(n_58833), .B(queue[121]), .C(n_58614), .Z(n_1363
		));
	notech_nao3 i_81678554(.A(n_58667), .B(queue[33]), .C(n_58943), .Z(n_1350
		));
	notech_and4 i_2525003(.A(n_2365100115), .B(n_2364100116), .C(n_2359100120
		), .D(n_2363100117), .Z(squeue_24100284));
	notech_nao3 i_75678572(.A(n_58833), .B(queue[120]), .C(n_58612), .Z(n_1347
		));
	notech_nao3 i_73978585(.A(n_58667), .B(queue[32]), .C(n_58943), .Z(n_1334
		));
	notech_and4 i_2425002(.A(n_2351100124), .B(n_235096484), .C(n_2345100127
		), .D(n_2349100125), .Z(squeue_23100285));
	notech_and4 i_72178603(.A(n_2887), .B(n_2915), .C(n_58833), .D(queue[119
		]), .Z(n_1331));
	notech_or2 i_70878616(.A(n_58930), .B(n_42946), .Z(n_1316));
	notech_and4 i_2325001(.A(n_2337), .B(n_2336), .C(n_2331), .D(n_2335), .Z
		(squeue_22100286));
	notech_and4 i_69078634(.A(n_2887), .B(n_2915), .C(n_58833), .D(queue[118
		]), .Z(n_1312));
	notech_nao3 i_67778647(.A(n_58667), .B(queue[30]), .C(n_58947), .Z(n_1293
		));
	notech_and4 i_2225000(.A(n_2323), .B(n_2322), .C(n_2317), .D(n_2321), .Z
		(squeue_21100287));
	notech_nao3 i_65878665(.A(n_58833), .B(queue[117]), .C(n_58612), .Z(n_1288
		));
	notech_nao3 i_64578678(.A(n_58667), .B(queue[29]), .C(n_58947), .Z(n_1270
		));
	notech_and4 i_2124999(.A(n_2309), .B(n_2308), .C(n_2303), .D(n_2307), .Z
		(squeue_20100288));
	notech_nao3 i_62778696(.A(n_58833), .B(queue[116]), .C(n_58614), .Z(n_1267
		));
	notech_nao3 i_61478709(.A(n_58667), .B(queue[28]), .C(n_58943), .Z(n_1254
		));
	notech_and4 i_2024998(.A(n_2295), .B(n_2294), .C(n_2289), .D(n_2293), .Z
		(squeue_19100289));
	notech_nao3 i_59678727(.A(n_58833), .B(queue[115]), .C(n_58612), .Z(n_1251
		));
	notech_nao3 i_58378740(.A(n_58667), .B(queue[27]), .C(n_58943), .Z(n_1238
		));
	notech_and4 i_1924997(.A(n_2281), .B(n_2280), .C(n_2275), .D(n_2279), .Z
		(squeue_18100290));
	notech_nao3 i_56578758(.A(n_58833), .B(queue[114]), .C(n_58609), .Z(n_1235
		));
	notech_nao3 i_55278771(.A(n_58667), .B(queue[26]), .C(n_58943), .Z(n_1222
		));
	notech_and4 i_1824996(.A(n_2267), .B(n_2266), .C(n_2261), .D(n_2265), .Z
		(squeue_17100291));
	notech_nao3 i_53478789(.A(n_58833), .B(queue[113]), .C(n_58609), .Z(n_1219
		));
	notech_nor2 i_5416(.A(n_60750), .B(wptr[0]), .Z(n_494100077));
	notech_reg purge_cnt_reg_0(.CP(n_62458), .D(n_40953), .CD(n_61370), .Q(purge_cnt
		[0]));
	notech_mux2 i_54565(.S(purge), .A(purge_cnt[0]), .B(n_27899861), .Z(n_40953
		));
	notech_reg purge_cnt_reg_1(.CP(n_62458), .D(n_40959), .CD(n_61370), .Q(purge_cnt
		[1]));
	notech_mux2 i_54573(.S(purge), .A(purge_cnt[1]), .B(n_27999862), .Z(n_40959
		));
	notech_reg purge_cnt_reg_2(.CP(n_62458), .D(n_40965), .CD(n_61370), .Q(purge_cnt
		[2]));
	notech_mux2 i_54581(.S(n_60778), .A(purge_cnt[2]), .B(n_28099863), .Z(n_40965
		));
	notech_reg purge_cnt_reg_3(.CP(n_62458), .D(n_40971), .CD(n_61370), .Q(purge_cnt
		[3]));
	notech_mux2 i_54589(.S(n_60778), .A(purge_cnt[3]), .B(n_28199864), .Z(n_40971
		));
	notech_reg purge_cnt_reg_4(.CP(n_62458), .D(n_40977), .CD(n_61370), .Q(purge_cnt
		[4]));
	notech_mux2 i_54597(.S(n_60778), .A(purge_cnt[4]), .B(n_28299865), .Z(n_40977
		));
	notech_reg purge_cnt_reg_5(.CP(n_62458), .D(n_40983), .CD(n_61371), .Q(purge_cnt
		[5]));
	notech_mux2 i_54605(.S(n_60778), .A(purge_cnt[5]), .B(n_28399866), .Z(n_40983
		));
	notech_reg purge_cnt_reg_6(.CP(n_62458), .D(n_40989), .CD(n_61371), .Q(purge_cnt
		[6]));
	notech_mux2 i_54613(.S(n_60778), .A(purge_cnt[6]), .B(n_28499867), .Z(n_40989
		));
	notech_reg purge_cnt_reg_7(.CP(n_62458), .D(n_40995), .CD(n_61371), .Q(purge_cnt
		[7]));
	notech_mux2 i_54621(.S(n_60778), .A(purge_cnt[7]), .B(n_28599868), .Z(n_40995
		));
	notech_reg purge_cnt_reg_8(.CP(n_62458), .D(n_41001), .CD(n_61370), .Q(purge_cnt
		[8]));
	notech_mux2 i_54629(.S(n_60778), .A(purge_cnt[8]), .B(n_28699869), .Z(n_41001
		));
	notech_reg purge_cnt_reg_9(.CP(n_62458), .D(n_41007), .CD(n_61371), .Q(purge_cnt
		[9]));
	notech_mux2 i_54637(.S(n_60778), .A(purge_cnt[9]), .B(n_28799870), .Z(n_41007
		));
	notech_reg purge_cnt_reg_10(.CP(n_62458), .D(n_41013), .CD(n_61370), .Q(purge_cnt
		[10]));
	notech_mux2 i_54645(.S(n_60778), .A(purge_cnt[10]), .B(n_28899871), .Z(n_41013
		));
	notech_reg_set purge_reg(.CP(n_62552), .D(n_41022), .SD(n_61370), .Q(purge
		));
	notech_nor2 i_54655(.A(purge_cnt[10]), .B(cacheD[148]), .Z(n_41022));
	notech_nao3 i_52178802(.A(n_58667), .B(queue[25]), .C(n_58943), .Z(n_1206
		));
	notech_reg fault_wptr_en_reg(.CP(n_62552), .D(n_41025), .CD(n_61370), .Q
		(fault_wptr_en));
	notech_mux2 i_54661(.S(n_377699581), .A(n_42907), .B(fault_wptr_en), .Z(n_41025
		));
	notech_reg pc_pg_fault_reg(.CP(n_62552), .D(n_41031), .CD(n_61369), .Q(pc_pg_fault
		));
	notech_mux2 i_54669(.S(n_42911), .A(pc_pg_fault), .B(n_42897), .Z(n_41031
		));
	notech_reg code_req_reg(.CP(n_62552), .D(n_41037), .CD(n_61369), .Q(code_req
		));
	notech_nand2 i_54677(.A(n_41039), .B(n_41040), .Z(n_41037));
	notech_or4 i_54678(.A(code_req), .B(n_487100070), .C(wptr[1]), .D(n_4532
		), .Z(n_41039));
	notech_nand3 i_54679(.A(n_942), .B(code_req), .C(n_937), .Z(n_41040));
	notech_and4 i_1724995(.A(n_2253), .B(n_2252), .C(n_2247), .D(n_2251), .Z
		(squeue_16100292));
	notech_reg addrshft_reg_0(.CP(n_62552), .D(n_41043), .CD(n_61369), .Q(addrshft
		[0]));
	notech_mux2 i_54685(.S(n_3777), .A(n_4645), .B(addrshft[0]), .Z(n_41043)
		);
	notech_nao3 i_50378820(.A(n_58833), .B(queue[112]), .C(n_58609), .Z(n_1203
		));
	notech_reg addrshft_reg_1(.CP(n_62552), .D(n_41049), .CD(n_61370), .Q(addrshft
		[1]));
	notech_mux2 i_54693(.S(n_3777), .A(n_4651), .B(addrshft[1]), .Z(n_41049)
		);
	notech_reg addrshft_reg_2(.CP(n_62552), .D(n_41055), .CD(n_61370), .Q(addrshft
		[2]));
	notech_mux2 i_54701(.S(n_3777), .A(n_4657), .B(addrshft[2]), .Z(n_41055)
		);
	notech_reg addrshft_reg_3(.CP(n_62552), .D(n_41061), .CD(n_61370), .Q(addrshft
		[3]));
	notech_mux2 i_54709(.S(n_3777), .A(n_4663), .B(addrshft[3]), .Z(n_41061)
		);
	notech_reg addrshft_reg_4(.CP(n_62552), .D(n_41067), .CD(n_61370), .Q(addrshft
		[4]));
	notech_mux2 i_54717(.S(n_3777), .A(n_24299825), .B(addrshft[4]), .Z(n_41067
		));
	notech_reg addrshft_reg_5(.CP(n_62552), .D(n_41073), .CD(n_61370), .Q(addrshft
		[5]));
	notech_mux2 i_54725(.S(n_3777), .A(n_42912), .B(addrshft[5]), .Z(n_41073
		));
	notech_reg wptr_reg_0(.CP(n_62552), .D(n_41079), .CD(n_61371), .Q(wptr[0
		]));
	notech_mux2 i_54733(.S(\nbus_94[0] ), .A(wptr[0]), .B(n_494100077), .Z(n_41079
		));
	notech_reg wptr_reg_1(.CP(n_62552), .D(n_41085), .CD(n_61372), .Q(wptr[1
		]));
	notech_mux2 i_54741(.S(\nbus_94[0] ), .A(wptr[1]), .B(n_134997819), .Z(n_41085
		));
	notech_reg fault_wptr_reg_0(.CP(n_62552), .D(n_41091), .CD(n_61372), .Q(fault_wptr
		[0]));
	notech_mux2 i_54749(.S(n_3778), .A(n_42915), .B(fault_wptr[0]), .Z(n_41091
		));
	notech_reg fault_wptr_reg_1(.CP(n_62552), .D(n_41097), .CD(n_61372), .Q(fault_wptr
		[1]));
	notech_mux2 i_54757(.S(n_3778), .A(n_42916), .B(fault_wptr[1]), .Z(n_41097
		));
	notech_reg addr_reg_0(.CP(n_62552), .D(n_41103), .CD(n_61372), .Q(iaddr[
		0]));
	notech_mux2 i_54765(.S(\nbus_93[0] ), .A(iaddr[0]), .B(n_27499857), .Z(n_41103
		));
	notech_reg addr_reg_1(.CP(n_62552), .D(n_41109), .CD(n_61372), .Q(iaddr[
		1]));
	notech_mux2 i_54773(.S(\nbus_93[0] ), .A(iaddr[1]), .B(n_27599858), .Z(n_41109
		));
	notech_reg addr_reg_2(.CP(n_62552), .D(n_41115), .CD(n_61372), .Q(iaddr[
		2]));
	notech_mux2 i_54781(.S(\nbus_93[0] ), .A(iaddr[2]), .B(n_27699859), .Z(n_41115
		));
	notech_reg addr_reg_3(.CP(n_62552), .D(n_41121), .CD(n_61372), .Q(iaddr[
		3]));
	notech_mux2 i_54789(.S(\nbus_93[0] ), .A(iaddr[3]), .B(n_27799860), .Z(n_41121
		));
	notech_nao3 i_49078833(.A(n_58709), .B(queue[32]), .C(n_58943), .Z(n_1190
		));
	notech_reg addr_reg_4(.CP(n_62552), .D(n_41127), .CD(n_61372), .Q(iaddr[
		4]));
	notech_mux2 i_54797(.S(\nbus_93[0] ), .A(iaddr[4]), .B(n_4355), .Z(n_41127
		));
	notech_reg addr_reg_5(.CP(n_62550), .D(n_41133), .CD(n_61372), .Q(iaddr[
		5]));
	notech_mux2 i_54805(.S(\nbus_93[0] ), .A(iaddr[5]), .B(n_4361), .Z(n_41133
		));
	notech_reg addr_reg_6(.CP(n_62550), .D(n_41139), .CD(n_61372), .Q(iaddr[
		6]));
	notech_mux2 i_54813(.S(\nbus_93[0] ), .A(iaddr[6]), .B(n_4367), .Z(n_41139
		));
	notech_and4 i_1624994(.A(n_2239), .B(n_2238), .C(n_2233), .D(n_2237), .Z
		(squeue_15100293));
	notech_reg addr_reg_7(.CP(n_62626), .D(n_41145), .CD(n_61372), .Q(iaddr[
		7]));
	notech_mux2 i_54821(.S(\nbus_93[0] ), .A(iaddr[7]), .B(n_4373), .Z(n_41145
		));
	notech_and4 i_47278851(.A(n_2887), .B(n_2915), .C(n_58833), .D(queue[111
		]), .Z(n_1187));
	notech_reg addr_reg_8(.CP(n_62626), .D(n_41151), .CD(n_61371), .Q(iaddr[
		8]));
	notech_mux2 i_54829(.S(\nbus_93[0] ), .A(iaddr[8]), .B(n_4379), .Z(n_41151
		));
	notech_reg addr_reg_9(.CP(n_62626), .D(n_41157), .CD(n_61371), .Q(iaddr[
		9]));
	notech_mux2 i_54837(.S(\nbus_93[0] ), .A(iaddr[9]), .B(n_4385), .Z(n_41157
		));
	notech_reg_set addr_reg_10(.CP(n_62626), .D(n_41163), .SD(n_61371), .Q(iaddr
		[10]));
	notech_mux2 i_54845(.S(\nbus_93[0] ), .A(iaddr[10]), .B(n_4391), .Z(n_41163
		));
	notech_reg_set addr_reg_11(.CP(n_62626), .D(n_41169), .SD(n_61371), .Q(iaddr
		[11]));
	notech_mux2 i_54853(.S(\nbus_93[0] ), .A(iaddr[11]), .B(n_4397), .Z(n_41169
		));
	notech_reg_set addr_reg_12(.CP(n_62626), .D(n_41175), .SD(n_61371), .Q(iaddr
		[12]));
	notech_mux2 i_54861(.S(\nbus_93[0] ), .A(iaddr[12]), .B(n_4403), .Z(n_41175
		));
	notech_reg_set addr_reg_13(.CP(n_62626), .D(n_41181), .SD(n_61371), .Q(iaddr
		[13]));
	notech_mux2 i_54869(.S(\nbus_93[0] ), .A(iaddr[13]), .B(n_4409), .Z(n_41181
		));
	notech_reg_set addr_reg_14(.CP(n_62626), .D(n_41187), .SD(n_61372), .Q(iaddr
		[14]));
	notech_mux2 i_54877(.S(\nbus_93[0] ), .A(iaddr[14]), .B(n_4415), .Z(n_41187
		));
	notech_reg_set addr_reg_15(.CP(n_62626), .D(n_41193), .SD(n_61371), .Q(iaddr
		[15]));
	notech_mux2 i_54885(.S(\nbus_93[0] ), .A(iaddr[15]), .B(n_4421), .Z(n_41193
		));
	notech_reg_set addr_reg_16(.CP(n_62626), .D(n_41199), .SD(n_61371), .Q(iaddr
		[16]));
	notech_mux2 i_54893(.S(n_60555), .A(iaddr[16]), .B(n_4427), .Z(n_41199)
		);
	notech_reg_set addr_reg_17(.CP(n_62626), .D(n_41205), .SD(n_61371), .Q(iaddr
		[17]));
	notech_mux2 i_54901(.S(n_60555), .A(iaddr[17]), .B(n_4433), .Z(n_41205)
		);
	notech_reg_set addr_reg_18(.CP(n_62626), .D(n_41211), .SD(n_61366), .Q(iaddr
		[18]));
	notech_mux2 i_54909(.S(n_60555), .A(iaddr[18]), .B(n_4439), .Z(n_41211)
		);
	notech_reg_set addr_reg_19(.CP(n_62626), .D(n_41217), .SD(n_61366), .Q(iaddr
		[19]));
	notech_mux2 i_54917(.S(n_60555), .A(iaddr[19]), .B(n_4445), .Z(n_41217)
		);
	notech_reg addr_reg_20(.CP(n_62626), .D(n_41223), .CD(n_61366), .Q(iaddr
		[20]));
	notech_mux2 i_54925(.S(n_60555), .A(iaddr[20]), .B(n_4451), .Z(n_41223)
		);
	notech_or2 i_45978864(.A(n_58930), .B(n_42938), .Z(n_1174));
	notech_reg addr_reg_21(.CP(n_62626), .D(n_41229), .CD(n_61366), .Q(iaddr
		[21]));
	notech_mux2 i_54933(.S(n_60555), .A(iaddr[21]), .B(n_4457), .Z(n_41229)
		);
	notech_reg addr_reg_22(.CP(n_62626), .D(n_41235), .CD(n_61366), .Q(iaddr
		[22]));
	notech_mux2 i_54941(.S(n_60555), .A(iaddr[22]), .B(n_4463), .Z(n_41235)
		);
	notech_reg addr_reg_23(.CP(n_62626), .D(n_41241), .CD(n_61367), .Q(iaddr
		[23]));
	notech_mux2 i_54949(.S(n_60555), .A(iaddr[23]), .B(n_4469), .Z(n_41241)
		);
	notech_and4 i_1424992(.A(n_2225), .B(n_2224), .C(n_2219), .D(n_2223), .Z
		(squeue_13100294));
	notech_reg addr_reg_24(.CP(n_62626), .D(n_41247), .CD(n_61367), .Q(iaddr
		[24]));
	notech_mux2 i_54957(.S(n_60555), .A(iaddr[24]), .B(n_4475), .Z(n_41247)
		);
	notech_nao3 i_44178882(.A(n_58837), .B(queue[109]), .C(n_58609), .Z(n_1171
		));
	notech_reg addr_reg_25(.CP(n_62550), .D(n_41253), .CD(n_61367), .Q(iaddr
		[25]));
	notech_mux2 i_54965(.S(n_60555), .A(iaddr[25]), .B(n_4481), .Z(n_41253)
		);
	notech_reg addr_reg_26(.CP(n_62550), .D(n_41259), .CD(n_61366), .Q(iaddr
		[26]));
	notech_mux2 i_54973(.S(n_60555), .A(iaddr[26]), .B(n_4487), .Z(n_41259)
		);
	notech_reg addr_reg_27(.CP(n_62550), .D(n_41265), .CD(n_61366), .Q(iaddr
		[27]));
	notech_mux2 i_54981(.S(n_60555), .A(iaddr[27]), .B(n_4493), .Z(n_41265)
		);
	notech_reg addr_reg_28(.CP(n_62550), .D(n_41271), .CD(n_61366), .Q(iaddr
		[28]));
	notech_mux2 i_54989(.S(n_60555), .A(iaddr[28]), .B(n_4499), .Z(n_41271)
		);
	notech_reg addr_reg_29(.CP(n_62550), .D(n_41277), .CD(n_61365), .Q(iaddr
		[29]));
	notech_mux2 i_54997(.S(n_60555), .A(iaddr[29]), .B(n_4505), .Z(n_41277)
		);
	notech_reg addr_reg_30(.CP(n_62550), .D(n_41283), .CD(n_61366), .Q(iaddr
		[30]));
	notech_mux2 i_55005(.S(n_60555), .A(iaddr[30]), .B(n_4511), .Z(n_41283)
		);
	notech_reg addr_reg_31(.CP(n_62550), .D(n_41289), .CD(n_61365), .Q(iaddr
		[31]));
	notech_mux2 i_55013(.S(n_60555), .A(iaddr[31]), .B(n_4517), .Z(n_41289)
		);
	notech_reg addrf_reg_0(.CP(n_62550), .D(iaddr[0]), .CD(n_61365), .Q(addrf
		[0]));
	notech_reg addrf_reg_1(.CP(n_62550), .D(iaddr[1]), .CD(n_61365), .Q(addrf
		[1]));
	notech_reg addrf_reg_2(.CP(n_62626), .D(iaddr[2]), .CD(n_61366), .Q(addrf
		[2]));
	notech_reg addrf_reg_3(.CP(n_62622), .D(iaddr[3]), .CD(n_61366), .Q(addrf
		[3]));
	notech_reg addrf_reg_4(.CP(n_62548), .D(iaddr[4]), .CD(n_61366), .Q(addrf
		[4]));
	notech_reg addrf_reg_5(.CP(n_62622), .D(iaddr[5]), .CD(n_61366), .Q(addrf
		[5]));
	notech_reg addrf_reg_6(.CP(n_62622), .D(iaddr[6]), .CD(n_61366), .Q(addrf
		[6]));
	notech_reg addrf_reg_7(.CP(n_62622), .D(iaddr[7]), .CD(n_61367), .Q(addrf
		[7]));
	notech_reg addrf_reg_8(.CP(n_62622), .D(iaddr[8]), .CD(n_61369), .Q(addrf
		[8]));
	notech_reg addrf_reg_9(.CP(n_62622), .D(iaddr[9]), .CD(n_61369), .Q(addrf
		[9]));
	notech_reg addrf_reg_10(.CP(n_62622), .D(iaddr[10]), .CD(n_61369), .Q(addrf
		[10]));
	notech_reg addrf_reg_11(.CP(n_62622), .D(iaddr[11]), .CD(n_61369), .Q(addrf
		[11]));
	notech_reg addrf_reg_12(.CP(n_62622), .D(iaddr[12]), .CD(n_61369), .Q(addrf
		[12]));
	notech_reg addrf_reg_13(.CP(n_62622), .D(iaddr[13]), .CD(n_61369), .Q(addrf
		[13]));
	notech_reg addrf_reg_14(.CP(n_62622), .D(iaddr[14]), .CD(n_61369), .Q(addrf
		[14]));
	notech_reg addrf_reg_15(.CP(n_62702), .D(iaddr[15]), .CD(n_61369), .Q(addrf
		[15]));
	notech_reg addrf_reg_16(.CP(n_62702), .D(iaddr[16]), .CD(n_61369), .Q(addrf
		[16]));
	notech_reg addrf_reg_17(.CP(n_62702), .D(iaddr[17]), .CD(n_61369), .Q(addrf
		[17]));
	notech_reg addrf_reg_18(.CP(n_62702), .D(iaddr[18]), .CD(n_61369), .Q(addrf
		[18]));
	notech_reg addrf_reg_19(.CP(n_62702), .D(iaddr[19]), .CD(n_61367), .Q(addrf
		[19]));
	notech_reg addrf_reg_20(.CP(n_62702), .D(iaddr[20]), .CD(n_61367), .Q(addrf
		[20]));
	notech_reg addrf_reg_21(.CP(n_62702), .D(iaddr[21]), .CD(n_61367), .Q(addrf
		[21]));
	notech_reg addrf_reg_22(.CP(n_62702), .D(iaddr[22]), .CD(n_61367), .Q(addrf
		[22]));
	notech_reg addrf_reg_23(.CP(n_62702), .D(iaddr[23]), .CD(n_61367), .Q(addrf
		[23]));
	notech_reg addrf_reg_24(.CP(n_62702), .D(iaddr[24]), .CD(n_61367), .Q(addrf
		[24]));
	notech_reg addrf_reg_25(.CP(n_62702), .D(iaddr[25]), .CD(n_61367), .Q(addrf
		[25]));
	notech_reg addrf_reg_26(.CP(n_62702), .D(iaddr[26]), .CD(n_61367), .Q(addrf
		[26]));
	notech_reg addrf_reg_27(.CP(n_62702), .D(iaddr[27]), .CD(n_61367), .Q(addrf
		[27]));
	notech_reg addrf_reg_28(.CP(n_62702), .D(iaddr[28]), .CD(n_61367), .Q(addrf
		[28]));
	notech_reg addrf_reg_29(.CP(n_62702), .D(iaddr[29]), .CD(n_61377), .Q(addrf
		[29]));
	notech_reg addrf_reg_30(.CP(n_62702), .D(iaddr[30]), .CD(n_61378), .Q(addrf
		[30]));
	notech_reg addrf_reg_31(.CP(n_62702), .D(iaddr[31]), .CD(n_61377), .Q(addrf
		[31]));
	notech_reg queue_reg_0(.CP(n_62702), .D(n_41359), .CD(n_61377), .Q(queue
		[0]));
	notech_mux2 i_55149(.S(n_55182), .A(n_2780), .B(queue[0]), .Z(n_41359)
		);
	notech_reg queue_reg_1(.CP(n_62622), .D(n_41365), .CD(n_61377), .Q(queue
		[1]));
	notech_mux2 i_55157(.S(n_55182), .A(n_2786), .B(queue[1]), .Z(n_41365)
		);
	notech_reg queue_reg_2(.CP(n_62548), .D(n_41371), .CD(n_61378), .Q(queue
		[2]));
	notech_mux2 i_55165(.S(n_55182), .A(n_2792), .B(queue[2]), .Z(n_41371)
		);
	notech_reg queue_reg_3(.CP(n_62624), .D(n_41377), .CD(n_61378), .Q(queue
		[3]));
	notech_mux2 i_55173(.S(n_55182), .A(n_2798), .B(queue[3]), .Z(n_41377)
		);
	notech_reg queue_reg_4(.CP(n_62624), .D(n_41383), .CD(n_61378), .Q(queue
		[4]));
	notech_mux2 i_55181(.S(n_55182), .A(n_2804), .B(queue[4]), .Z(n_41383)
		);
	notech_reg queue_reg_5(.CP(n_62624), .D(n_41389), .CD(n_61378), .Q(queue
		[5]));
	notech_mux2 i_55189(.S(n_55182), .A(n_2810), .B(queue[5]), .Z(n_41389)
		);
	notech_nao3 i_42878895(.A(n_58667), .B(queue[21]), .C(n_58943), .Z(n_1157
		));
	notech_reg queue_reg_6(.CP(n_62624), .D(n_41395), .CD(n_61378), .Q(queue
		[6]));
	notech_mux2 i_55197(.S(n_55182), .A(n_2816), .B(queue[6]), .Z(n_41395)
		);
	notech_reg queue_reg_7(.CP(n_62624), .D(n_41401), .CD(n_61377), .Q(queue
		[7]));
	notech_mux2 i_55205(.S(n_55182), .A(n_2822), .B(queue[7]), .Z(n_41401)
		);
	notech_reg queue_reg_8(.CP(n_62624), .D(n_41407), .CD(n_61377), .Q(queue
		[8]));
	notech_mux2 i_55213(.S(n_55182), .A(n_2828), .B(queue[8]), .Z(n_41407)
		);
	notech_and4 i_1324991(.A(n_2211), .B(n_2210), .C(n_2205), .D(n_2209), .Z
		(squeue_12100295));
	notech_reg queue_reg_9(.CP(n_62624), .D(n_41413), .CD(n_61377), .Q(queue
		[9]));
	notech_mux2 i_55221(.S(n_55182), .A(n_2834), .B(queue[9]), .Z(n_41413)
		);
	notech_nao3 i_41078913(.A(n_58837), .B(queue[108]), .C(n_58609), .Z(n_1152
		));
	notech_reg queue_reg_10(.CP(n_62624), .D(n_41419), .CD(n_61377), .Q(queue
		[10]));
	notech_mux2 i_55229(.S(n_55182), .A(n_2840), .B(queue[10]), .Z(n_41419)
		);
	notech_reg queue_reg_11(.CP(n_62624), .D(n_41425), .CD(n_61376), .Q(queue
		[11]));
	notech_mux2 i_55237(.S(n_55182), .A(n_2846), .B(queue[11]), .Z(n_41425)
		);
	notech_reg queue_reg_12(.CP(n_62624), .D(n_41431), .CD(n_61377), .Q(queue
		[12]));
	notech_mux2 i_55245(.S(n_55182), .A(n_2852), .B(queue[12]), .Z(n_41431)
		);
	notech_reg queue_reg_13(.CP(n_62624), .D(n_41437), .CD(n_61377), .Q(queue
		[13]));
	notech_mux2 i_55253(.S(n_55182), .A(n_2858), .B(queue[13]), .Z(n_41437)
		);
	notech_reg queue_reg_14(.CP(n_62624), .D(n_41443), .CD(n_61377), .Q(queue
		[14]));
	notech_mux2 i_55261(.S(n_55182), .A(n_2864), .B(queue[14]), .Z(n_41443)
		);
	notech_reg queue_reg_15(.CP(n_62624), .D(n_41449), .CD(n_61377), .Q(queue
		[15]));
	notech_mux2 i_55269(.S(n_55182), .A(n_2870), .B(queue[15]), .Z(n_41449)
		);
	notech_reg queue_reg_16(.CP(n_62624), .D(n_41455), .CD(n_61377), .Q(queue
		[16]));
	notech_mux2 i_55277(.S(n_55180), .A(n_2876), .B(queue[16]), .Z(n_41455)
		);
	notech_reg queue_reg_17(.CP(n_62624), .D(n_41461), .CD(n_61377), .Q(queue
		[17]));
	notech_mux2 i_55285(.S(n_55180), .A(n_2882), .B(queue[17]), .Z(n_41461)
		);
	notech_reg queue_reg_18(.CP(n_62624), .D(n_41467), .CD(n_61378), .Q(queue
		[18]));
	notech_mux2 i_55293(.S(n_55180), .A(n_2888), .B(queue[18]), .Z(n_41467)
		);
	notech_reg queue_reg_19(.CP(n_62624), .D(n_41473), .CD(n_61379), .Q(queue
		[19]));
	notech_mux2 i_55301(.S(n_55180), .A(n_2894), .B(queue[19]), .Z(n_41473)
		);
	notech_reg queue_reg_20(.CP(n_62624), .D(n_41479), .CD(n_61379), .Q(queue
		[20]));
	notech_mux2 i_55309(.S(n_55180), .A(n_2900), .B(queue[20]), .Z(n_41479)
		);
	notech_reg queue_reg_21(.CP(n_62624), .D(n_41485), .CD(n_61379), .Q(queue
		[21]));
	notech_mux2 i_55317(.S(n_55180), .A(n_136197831), .B(queue[21]), .Z(n_41485
		));
	notech_reg queue_reg_22(.CP(n_62548), .D(n_41491), .CD(n_61379), .Q(queue
		[22]));
	notech_mux2 i_55325(.S(n_55180), .A(n_2912), .B(queue[22]), .Z(n_41491)
		);
	notech_nao3 i_39778926(.A(n_58667), .B(queue[20]), .C(n_58947), .Z(n_1137
		));
	notech_reg queue_reg_23(.CP(n_62548), .D(n_41497), .CD(n_61379), .Q(queue
		[23]));
	notech_mux2 i_55333(.S(n_55180), .A(n_2918), .B(queue[23]), .Z(n_41497)
		);
	notech_reg queue_reg_24(.CP(n_62548), .D(n_41503), .CD(n_61379), .Q(queue
		[24]));
	notech_mux2 i_55341(.S(n_55180), .A(n_2924), .B(queue[24]), .Z(n_41503)
		);
	notech_reg queue_reg_25(.CP(n_62548), .D(n_41509), .CD(n_61379), .Q(queue
		[25]));
	notech_mux2 i_55349(.S(n_55180), .A(n_2930), .B(queue[25]), .Z(n_41509)
		);
	notech_and4 i_1224990(.A(n_2197), .B(n_2196), .C(n_2191), .D(n_2195), .Z
		(squeue_11100296));
	notech_reg queue_reg_26(.CP(n_62548), .D(n_41515), .CD(n_61379), .Q(queue
		[26]));
	notech_mux2 i_55357(.S(n_55180), .A(n_2936), .B(queue[26]), .Z(n_41515)
		);
	notech_nao3 i_37978944(.A(n_58837), .B(queue[107]), .C(n_58609), .Z(n_1132
		));
	notech_reg queue_reg_27(.CP(n_62548), .D(n_41521), .CD(n_61379), .Q(queue
		[27]));
	notech_mux2 i_55365(.S(n_55180), .A(n_2942), .B(queue[27]), .Z(n_41521)
		);
	notech_reg queue_reg_28(.CP(n_62548), .D(n_41527), .CD(n_61379), .Q(queue
		[28]));
	notech_mux2 i_55373(.S(n_55180), .A(n_2948), .B(queue[28]), .Z(n_41527)
		);
	notech_reg queue_reg_29(.CP(n_62548), .D(n_41533), .CD(n_61379), .Q(queue
		[29]));
	notech_mux2 i_55381(.S(n_55180), .A(n_2954), .B(queue[29]), .Z(n_41533)
		);
	notech_reg queue_reg_30(.CP(n_62548), .D(n_41539), .CD(n_61378), .Q(queue
		[30]));
	notech_mux2 i_55389(.S(n_55180), .A(n_2960), .B(queue[30]), .Z(n_41539)
		);
	notech_reg queue_reg_31(.CP(n_62702), .D(n_41545), .CD(n_61378), .Q(queue
		[31]));
	notech_mux2 i_55397(.S(n_55180), .A(n_2966), .B(queue[31]), .Z(n_41545)
		);
	notech_reg queue_reg_32(.CP(n_62616), .D(n_41551), .CD(n_61378), .Q(queue
		[32]));
	notech_mux2 i_55405(.S(n_55187), .A(n_2972), .B(queue[32]), .Z(n_41551)
		);
	notech_reg queue_reg_33(.CP(n_62616), .D(n_41557), .CD(n_61378), .Q(queue
		[33]));
	notech_mux2 i_55413(.S(n_55187), .A(n_2978), .B(queue[33]), .Z(n_41557)
		);
	notech_reg queue_reg_34(.CP(n_62616), .D(n_41563), .CD(n_61378), .Q(queue
		[34]));
	notech_mux2 i_55421(.S(n_55187), .A(n_2984), .B(queue[34]), .Z(n_41563)
		);
	notech_reg queue_reg_35(.CP(n_62616), .D(n_41569), .CD(n_61379), .Q(queue
		[35]));
	notech_mux2 i_55429(.S(n_55187), .A(n_2990), .B(queue[35]), .Z(n_41569)
		);
	notech_reg queue_reg_36(.CP(n_62616), .D(n_41575), .CD(n_61379), .Q(queue
		[36]));
	notech_mux2 i_55437(.S(n_55187), .A(n_2996), .B(queue[36]), .Z(n_41575)
		);
	notech_reg queue_reg_37(.CP(n_62616), .D(n_41581), .CD(n_61379), .Q(queue
		[37]));
	notech_mux2 i_55445(.S(n_55187), .A(n_3002), .B(queue[37]), .Z(n_41581)
		);
	notech_reg queue_reg_38(.CP(n_62616), .D(n_41587), .CD(n_61378), .Q(queue
		[38]));
	notech_mux2 i_55453(.S(n_55187), .A(n_3008), .B(queue[38]), .Z(n_41587)
		);
	notech_reg queue_reg_39(.CP(n_62616), .D(n_41593), .CD(n_61378), .Q(queue
		[39]));
	notech_mux2 i_55461(.S(n_55187), .A(n_3014), .B(queue[39]), .Z(n_41593)
		);
	notech_nao3 i_36678957(.A(n_58667), .B(queue[19]), .C(n_58947), .Z(n_1119
		));
	notech_reg queue_reg_40(.CP(n_62616), .D(n_41599), .CD(n_61373), .Q(queue
		[40]));
	notech_mux2 i_55469(.S(n_55187), .A(n_3020), .B(queue[40]), .Z(n_41599)
		);
	notech_reg queue_reg_41(.CP(n_62616), .D(n_41605), .CD(n_61373), .Q(queue
		[41]));
	notech_mux2 i_55477(.S(n_55187), .A(n_3026), .B(queue[41]), .Z(n_41605)
		);
	notech_reg queue_reg_42(.CP(n_62616), .D(n_41611), .CD(n_61373), .Q(queue
		[42]));
	notech_mux2 i_55485(.S(n_55187), .A(n_3032), .B(queue[42]), .Z(n_41611)
		);
	notech_and4 i_1124989(.A(n_2183), .B(n_2182), .C(n_2177), .D(n_2181), .Z
		(squeue_10100297));
	notech_reg queue_reg_43(.CP(n_62698), .D(n_41617), .CD(n_61373), .Q(queue
		[43]));
	notech_mux2 i_55493(.S(n_55187), .A(n_3038), .B(queue[43]), .Z(n_41617)
		);
	notech_nao3 i_34878975(.A(n_58837), .B(queue[106]), .C(n_58609), .Z(n_1116
		));
	notech_reg queue_reg_44(.CP(n_62698), .D(n_41623), .CD(n_61373), .Q(queue
		[44]));
	notech_mux2 i_55501(.S(n_55187), .A(n_3044), .B(queue[44]), .Z(n_41623)
		);
	notech_reg queue_reg_45(.CP(n_62698), .D(n_41629), .CD(n_61375), .Q(queue
		[45]));
	notech_mux2 i_55509(.S(n_55187), .A(n_3050), .B(queue[45]), .Z(n_41629)
		);
	notech_reg queue_reg_46(.CP(n_62698), .D(n_41635), .CD(n_61375), .Q(queue
		[46]));
	notech_mux2 i_55517(.S(n_55187), .A(n_3056), .B(queue[46]), .Z(n_41635)
		);
	notech_reg queue_reg_47(.CP(n_62698), .D(n_41641), .CD(n_61375), .Q(queue
		[47]));
	notech_mux2 i_55525(.S(n_55187), .A(n_3062), .B(queue[47]), .Z(n_41641)
		);
	notech_reg queue_reg_48(.CP(n_62698), .D(n_41647), .CD(n_61375), .Q(queue
		[48]));
	notech_mux2 i_55533(.S(n_55185), .A(n_3068), .B(queue[48]), .Z(n_41647)
		);
	notech_reg queue_reg_49(.CP(n_62698), .D(n_41653), .CD(n_61375), .Q(queue
		[49]));
	notech_mux2 i_55541(.S(n_55185), .A(n_3074), .B(queue[49]), .Z(n_41653)
		);
	notech_reg queue_reg_50(.CP(n_62698), .D(n_41659), .CD(n_61373), .Q(queue
		[50]));
	notech_mux2 i_55549(.S(n_55185), .A(n_3080), .B(queue[50]), .Z(n_41659)
		);
	notech_reg queue_reg_51(.CP(n_62698), .D(n_41665), .CD(n_61373), .Q(queue
		[51]));
	notech_mux2 i_55557(.S(n_55185), .A(n_135897828), .B(queue[51]), .Z(n_41665
		));
	notech_reg queue_reg_52(.CP(n_62698), .D(n_41671), .CD(n_61373), .Q(queue
		[52]));
	notech_mux2 i_55565(.S(n_55185), .A(n_3092), .B(queue[52]), .Z(n_41671)
		);
	notech_reg queue_reg_53(.CP(n_62698), .D(n_41677), .CD(n_61373), .Q(queue
		[53]));
	notech_mux2 i_55573(.S(n_55185), .A(n_135597825), .B(queue[53]), .Z(n_41677
		));
	notech_reg queue_reg_54(.CP(n_62698), .D(n_41683), .CD(n_61372), .Q(queue
		[54]));
	notech_mux2 i_55581(.S(n_55185), .A(n_3104), .B(queue[54]), .Z(n_41683)
		);
	notech_reg queue_reg_55(.CP(n_62698), .D(n_41689), .CD(n_61372), .Q(queue
		[55]));
	notech_mux2 i_55589(.S(n_55185), .A(n_3110), .B(queue[55]), .Z(n_41689)
		);
	notech_reg queue_reg_56(.CP(n_62698), .D(n_41695), .CD(n_61373), .Q(queue
		[56]));
	notech_mux2 i_55597(.S(n_55185), .A(n_3116), .B(queue[56]), .Z(n_41695)
		);
	notech_nao3 i_33578988(.A(n_58667), .B(queue[18]), .C(n_58947), .Z(n_1103
		));
	notech_reg queue_reg_57(.CP(n_62698), .D(n_41701), .CD(n_61373), .Q(queue
		[57]));
	notech_mux2 i_55605(.S(n_55185), .A(n_3122), .B(queue[57]), .Z(n_41701)
		);
	notech_reg queue_reg_58(.CP(n_62698), .D(n_41707), .CD(n_61373), .Q(queue
		[58]));
	notech_mux2 i_55613(.S(n_55185), .A(n_3128), .B(queue[58]), .Z(n_41707)
		);
	notech_reg queue_reg_59(.CP(n_62698), .D(n_41713), .CD(n_61373), .Q(queue
		[59]));
	notech_mux2 i_55621(.S(n_55185), .A(n_3134), .B(queue[59]), .Z(n_41713)
		);
	notech_and4 i_1024988(.A(n_2169), .B(n_2168), .C(n_2163), .D(n_2167), .Z
		(squeue_9100298));
	notech_reg queue_reg_60(.CP(n_62698), .D(n_41719), .CD(n_61373), .Q(queue
		[60]));
	notech_mux2 i_55629(.S(n_55185), .A(n_3140), .B(queue[60]), .Z(n_41719)
		);
	notech_nao3 i_31779006(.A(n_58837), .B(queue[105]), .C(n_58612), .Z(n_1100
		));
	notech_reg queue_reg_61(.CP(n_62698), .D(n_41725), .CD(n_61375), .Q(queue
		[61]));
	notech_mux2 i_55637(.S(n_55185), .A(n_3146), .B(queue[61]), .Z(n_41725)
		);
	notech_reg queue_reg_62(.CP(n_62746), .D(n_41731), .CD(n_61376), .Q(queue
		[62]));
	notech_mux2 i_55645(.S(n_55185), .A(n_3152), .B(queue[62]), .Z(n_41731)
		);
	notech_reg queue_reg_63(.CP(n_62746), .D(n_41737), .CD(n_61376), .Q(queue
		[63]));
	notech_mux2 i_55653(.S(n_55185), .A(n_3158), .B(queue[63]), .Z(n_41737)
		);
	notech_reg queue_reg_64(.CP(n_62746), .D(n_41743), .CD(n_61376), .Q(queue
		[64]));
	notech_mux2 i_55661(.S(n_55172), .A(n_3164), .B(queue[64]), .Z(n_41743)
		);
	notech_reg queue_reg_65(.CP(n_62746), .D(n_41749), .CD(n_61376), .Q(queue
		[65]));
	notech_mux2 i_55669(.S(n_55172), .A(n_3170), .B(queue[65]), .Z(n_41749)
		);
	notech_reg queue_reg_66(.CP(n_62746), .D(n_41755), .CD(n_61376), .Q(queue
		[66]));
	notech_mux2 i_55677(.S(n_55172), .A(n_3176), .B(queue[66]), .Z(n_41755)
		);
	notech_reg queue_reg_67(.CP(n_62746), .D(n_41761), .CD(n_61376), .Q(queue
		[67]));
	notech_mux2 i_55685(.S(n_55172), .A(n_3182), .B(queue[67]), .Z(n_41761)
		);
	notech_reg queue_reg_68(.CP(n_62746), .D(n_41767), .CD(n_61376), .Q(queue
		[68]));
	notech_mux2 i_55693(.S(n_55172), .A(n_3188), .B(queue[68]), .Z(n_41767)
		);
	notech_reg queue_reg_69(.CP(n_62746), .D(n_41773), .CD(n_61376), .Q(queue
		[69]));
	notech_mux2 i_55701(.S(n_55172), .A(n_3194), .B(queue[69]), .Z(n_41773)
		);
	notech_reg queue_reg_70(.CP(n_62746), .D(n_41779), .CD(n_61376), .Q(queue
		[70]));
	notech_mux2 i_55709(.S(n_55172), .A(n_3200), .B(queue[70]), .Z(n_41779)
		);
	notech_reg queue_reg_71(.CP(n_62746), .D(n_41785), .CD(n_61376), .Q(queue
		[71]));
	notech_mux2 i_55717(.S(n_55172), .A(n_3206), .B(queue[71]), .Z(n_41785)
		);
	notech_reg queue_reg_72(.CP(n_62746), .D(n_41791), .CD(n_61376), .Q(queue
		[72]));
	notech_mux2 i_55725(.S(n_55172), .A(n_3212), .B(queue[72]), .Z(n_41791)
		);
	notech_reg queue_reg_73(.CP(n_62746), .D(n_41797), .CD(n_61375), .Q(queue
		[73]));
	notech_mux2 i_55733(.S(n_55172), .A(n_3218), .B(queue[73]), .Z(n_41797)
		);
	notech_nao3 i_30479019(.A(n_58667), .B(queue[17]), .C(n_58947), .Z(n_1087
		));
	notech_reg queue_reg_74(.CP(n_62746), .D(n_41803), .CD(n_61375), .Q(queue
		[74]));
	notech_mux2 i_55741(.S(n_55172), .A(n_3224), .B(queue[74]), .Z(n_41803)
		);
	notech_reg queue_reg_75(.CP(n_62746), .D(n_41809), .CD(n_61375), .Q(queue
		[75]));
	notech_mux2 i_55749(.S(n_55172), .A(n_3230), .B(queue[75]), .Z(n_41809)
		);
	notech_reg queue_reg_76(.CP(n_62746), .D(n_41815), .CD(n_61375), .Q(queue
		[76]));
	notech_mux2 i_55757(.S(n_55172), .A(n_3236), .B(queue[76]), .Z(n_41815)
		);
	notech_and4 i_824986(.A(n_2155), .B(n_2154), .C(n_2149), .D(n_2153), .Z(squeue_7100299
		));
	notech_reg queue_reg_77(.CP(n_62746), .D(n_41821), .CD(n_61375), .Q(queue
		[77]));
	notech_mux2 i_55765(.S(n_55172), .A(n_3242), .B(queue[77]), .Z(n_41821)
		);
	notech_and4 i_28679037(.A(n_2887), .B(n_2915), .C(n_58837), .D(queue[103
		]), .Z(n_1084));
	notech_reg queue_reg_78(.CP(n_62746), .D(n_41827), .CD(n_61376), .Q(queue
		[78]));
	notech_mux2 i_55773(.S(n_55172), .A(n_3248), .B(queue[78]), .Z(n_41827)
		);
	notech_reg queue_reg_79(.CP(n_62746), .D(n_41833), .CD(n_61376), .Q(queue
		[79]));
	notech_mux2 i_55781(.S(n_55172), .A(n_3254), .B(queue[79]), .Z(n_41833)
		);
	notech_reg queue_reg_80(.CP(n_62746), .D(n_41839), .CD(n_61375), .Q(queue
		[80]));
	notech_mux2 i_55789(.S(n_55170), .A(n_135297822), .B(queue[80]), .Z(n_41839
		));
	notech_reg queue_reg_81(.CP(n_62746), .D(n_41845), .CD(n_61375), .Q(queue
		[81]));
	notech_mux2 i_55797(.S(n_55170), .A(n_3266), .B(queue[81]), .Z(n_41845)
		);
	notech_reg queue_reg_82(.CP(n_62696), .D(n_41851), .CD(n_61375), .Q(queue
		[82]));
	notech_mux2 i_55805(.S(n_55170), .A(n_3272), .B(queue[82]), .Z(n_41851)
		);
	notech_reg queue_reg_83(.CP(n_62696), .D(n_41857), .CD(n_61365), .Q(queue
		[83]));
	notech_mux2 i_55813(.S(n_55170), .A(n_3278), .B(queue[83]), .Z(n_41857)
		);
	notech_reg queue_reg_84(.CP(n_62696), .D(n_41863), .CD(n_61355), .Q(queue
		[84]));
	notech_mux2 i_55821(.S(n_55170), .A(n_3284), .B(queue[84]), .Z(n_41863)
		);
	notech_reg queue_reg_85(.CP(n_62696), .D(n_41869), .CD(n_61355), .Q(queue
		[85]));
	notech_mux2 i_55829(.S(n_55170), .A(n_3290), .B(queue[85]), .Z(n_41869)
		);
	notech_reg queue_reg_86(.CP(n_62696), .D(n_41875), .CD(n_61355), .Q(queue
		[86]));
	notech_mux2 i_55837(.S(n_55170), .A(n_3296), .B(queue[86]), .Z(n_41875)
		);
	notech_reg queue_reg_87(.CP(n_62696), .D(n_41881), .CD(n_61355), .Q(queue
		[87]));
	notech_mux2 i_55845(.S(n_55170), .A(n_3302), .B(queue[87]), .Z(n_41881)
		);
	notech_reg queue_reg_88(.CP(n_62696), .D(n_41887), .CD(n_61355), .Q(queue
		[88]));
	notech_mux2 i_55853(.S(n_55170), .A(n_3308), .B(queue[88]), .Z(n_41887)
		);
	notech_reg queue_reg_89(.CP(n_62696), .D(n_41893), .CD(n_61355), .Q(queue
		[89]));
	notech_mux2 i_55861(.S(n_55170), .A(n_3314), .B(queue[89]), .Z(n_41893)
		);
	notech_reg queue_reg_90(.CP(n_62696), .D(n_41899), .CD(n_61355), .Q(queue
		[90]));
	notech_mux2 i_55869(.S(n_55170), .A(n_3320), .B(queue[90]), .Z(n_41899)
		);
	notech_or2 i_27379050(.A(n_58930), .B(n_42930), .Z(n_1071));
	notech_reg queue_reg_91(.CP(n_62696), .D(n_41905), .CD(n_61355), .Q(queue
		[91]));
	notech_mux2 i_55877(.S(n_55170), .A(n_3326), .B(queue[91]), .Z(n_41905)
		);
	notech_reg queue_reg_92(.CP(n_62696), .D(n_41911), .CD(n_61355), .Q(queue
		[92]));
	notech_mux2 i_55885(.S(n_55170), .A(n_3332), .B(queue[92]), .Z(n_41911)
		);
	notech_reg queue_reg_93(.CP(n_62696), .D(n_41917), .CD(n_61355), .Q(queue
		[93]));
	notech_mux2 i_55893(.S(n_55170), .A(n_3338), .B(queue[93]), .Z(n_41917)
		);
	notech_and4 i_724985(.A(n_2141), .B(n_2140), .C(n_2135), .D(n_2139), .Z(squeue_6100300
		));
	notech_reg queue_reg_94(.CP(n_62700), .D(n_41923), .CD(n_61355), .Q(queue
		[94]));
	notech_mux2 i_55901(.S(n_55170), .A(n_3344), .B(queue[94]), .Z(n_41923)
		);
	notech_and4 i_25579068(.A(n_58837), .B(n_2887), .C(n_2915), .D(queue[102
		]), .Z(n_1068));
	notech_reg queue_reg_95(.CP(n_62618), .D(n_41929), .CD(n_61354), .Q(queue
		[95]));
	notech_mux2 i_55909(.S(n_55170), .A(n_3350), .B(queue[95]), .Z(n_41929)
		);
	notech_reg queue_reg_96(.CP(n_62618), .D(n_41935), .CD(n_61354), .Q(queue
		[96]));
	notech_mux2 i_55917(.S(n_55177), .A(n_3356), .B(queue[96]), .Z(n_41935)
		);
	notech_reg queue_reg_97(.CP(n_62618), .D(n_41941), .CD(n_61354), .Q(queue
		[97]));
	notech_mux2 i_55925(.S(n_55177), .A(n_3362), .B(queue[97]), .Z(n_41941)
		);
	notech_reg queue_reg_98(.CP(n_62618), .D(n_41947), .CD(n_61354), .Q(queue
		[98]));
	notech_mux2 i_55933(.S(n_55177), .A(n_3368), .B(queue[98]), .Z(n_41947)
		);
	notech_reg queue_reg_99(.CP(n_62618), .D(n_41953), .CD(n_61354), .Q(queue
		[99]));
	notech_mux2 i_55941(.S(n_55177), .A(n_3374), .B(queue[99]), .Z(n_41953)
		);
	notech_reg queue_reg_100(.CP(n_62618), .D(n_41959), .CD(n_61354), .Q(queue
		[100]));
	notech_mux2 i_55949(.S(n_55177), .A(n_3380), .B(queue[100]), .Z(n_41959)
		);
	notech_reg queue_reg_101(.CP(n_62618), .D(n_41965), .CD(n_61355), .Q(queue
		[101]));
	notech_mux2 i_55957(.S(n_55177), .A(n_3386), .B(queue[101]), .Z(n_41965)
		);
	notech_reg queue_reg_102(.CP(n_62618), .D(n_41971), .CD(n_61354), .Q(queue
		[102]));
	notech_mux2 i_55965(.S(n_55177), .A(n_3392), .B(queue[102]), .Z(n_41971)
		);
	notech_reg queue_reg_103(.CP(n_62618), .D(n_41977), .CD(n_61354), .Q(queue
		[103]));
	notech_mux2 i_55973(.S(n_55177), .A(n_3398), .B(queue[103]), .Z(n_41977)
		);
	notech_reg queue_reg_104(.CP(n_62700), .D(n_41983), .CD(n_61354), .Q(queue
		[104]));
	notech_mux2 i_55981(.S(n_55177), .A(n_3404), .B(queue[104]), .Z(n_41983)
		);
	notech_reg queue_reg_105(.CP(n_62700), .D(n_41989), .CD(n_61355), .Q(queue
		[105]));
	notech_mux2 i_55989(.S(n_55177), .A(n_3410), .B(queue[105]), .Z(n_41989)
		);
	notech_reg queue_reg_106(.CP(n_62700), .D(n_41995), .CD(n_61358), .Q(queue
		[106]));
	notech_mux2 i_55997(.S(n_55177), .A(n_3416), .B(queue[106]), .Z(n_41995)
		);
	notech_reg queue_reg_107(.CP(n_62700), .D(n_42001), .CD(n_61358), .Q(queue
		[107]));
	notech_mux2 i_56005(.S(n_55177), .A(n_3422), .B(queue[107]), .Z(n_42001)
		);
	notech_nao3 i_24279081(.A(queue[14]), .B(n_58667), .C(n_58947), .Z(n_1055
		));
	notech_reg queue_reg_108(.CP(n_62700), .D(n_42007), .CD(n_61357), .Q(queue
		[108]));
	notech_mux2 i_56013(.S(n_55177), .A(n_3428), .B(queue[108]), .Z(n_42007)
		);
	notech_reg queue_reg_109(.CP(n_62700), .D(n_42013), .CD(n_61357), .Q(queue
		[109]));
	notech_mux2 i_56021(.S(n_55177), .A(n_3434), .B(queue[109]), .Z(n_42013)
		);
	notech_reg queue_reg_110(.CP(n_62700), .D(n_42019), .CD(n_61357), .Q(queue
		[110]));
	notech_mux2 i_56029(.S(n_55177), .A(n_3440), .B(queue[110]), .Z(n_42019)
		);
	notech_and4 i_624984(.A(n_2127), .B(n_2126), .C(n_2121), .D(n_2125), .Z(squeue_5100301
		));
	notech_reg queue_reg_111(.CP(n_62700), .D(n_42025), .CD(n_61358), .Q(queue
		[111]));
	notech_mux2 i_56037(.S(n_55177), .A(n_3446), .B(queue[111]), .Z(n_42025)
		);
	notech_nao3 i_22479099(.A(n_58833), .B(queue[101]), .C(n_58612), .Z(n_1052
		));
	notech_reg queue_reg_112(.CP(n_62700), .D(n_42031), .CD(n_61358), .Q(queue
		[112]));
	notech_mux2 i_56045(.S(n_55175), .A(n_3452), .B(queue[112]), .Z(n_42031)
		);
	notech_reg queue_reg_113(.CP(n_62700), .D(n_42037), .CD(n_61358), .Q(queue
		[113]));
	notech_mux2 i_56053(.S(n_55175), .A(n_3458), .B(queue[113]), .Z(n_42037)
		);
	notech_reg queue_reg_114(.CP(n_62700), .D(n_42043), .CD(n_61358), .Q(queue
		[114]));
	notech_mux2 i_56061(.S(n_55175), .A(n_3464), .B(queue[114]), .Z(n_42043)
		);
	notech_reg queue_reg_115(.CP(n_62700), .D(n_42049), .CD(n_61358), .Q(queue
		[115]));
	notech_mux2 i_56069(.S(n_55175), .A(n_3470), .B(queue[115]), .Z(n_42049)
		);
	notech_reg queue_reg_116(.CP(n_62700), .D(n_42055), .CD(n_61357), .Q(queue
		[116]));
	notech_mux2 i_56077(.S(n_55175), .A(n_3476), .B(queue[116]), .Z(n_42055)
		);
	notech_reg queue_reg_117(.CP(n_62700), .D(n_42061), .CD(n_61357), .Q(queue
		[117]));
	notech_mux2 i_56085(.S(n_55175), .A(n_3482), .B(queue[117]), .Z(n_42061)
		);
	notech_reg queue_reg_118(.CP(n_62700), .D(n_42067), .CD(n_61357), .Q(queue
		[118]));
	notech_mux2 i_56093(.S(n_55175), .A(n_3488), .B(queue[118]), .Z(n_42067)
		);
	notech_reg queue_reg_119(.CP(n_62700), .D(n_42073), .CD(n_61357), .Q(queue
		[119]));
	notech_mux2 i_56101(.S(n_55175), .A(n_3494), .B(queue[119]), .Z(n_42073)
		);
	notech_reg queue_reg_120(.CP(n_62700), .D(n_42079), .CD(n_61357), .Q(queue
		[120]));
	notech_mux2 i_56109(.S(n_55175), .A(n_3500), .B(queue[120]), .Z(n_42079)
		);
	notech_reg queue_reg_121(.CP(n_62700), .D(n_42085), .CD(n_61357), .Q(queue
		[121]));
	notech_mux2 i_56117(.S(n_55175), .A(n_3506), .B(queue[121]), .Z(n_42085)
		);
	notech_reg queue_reg_122(.CP(n_62618), .D(n_42091), .CD(n_61357), .Q(queue
		[122]));
	notech_mux2 i_56125(.S(n_55175), .A(n_3512), .B(queue[122]), .Z(n_42091)
		);
	notech_reg queue_reg_123(.CP(n_62618), .D(n_42097), .CD(n_61357), .Q(queue
		[123]));
	notech_mux2 i_56133(.S(n_55175), .A(n_3518), .B(queue[123]), .Z(n_42097)
		);
	notech_reg queue_reg_124(.CP(n_62620), .D(n_42103), .CD(n_61357), .Q(queue
		[124]));
	notech_mux2 i_56141(.S(n_55175), .A(n_3524), .B(queue[124]), .Z(n_42103)
		);
	notech_nao3 i_21179112(.A(n_58667), .B(queue[13]), .C(n_58947), .Z(n_1039
		));
	notech_reg queue_reg_125(.CP(n_62620), .D(n_42109), .CD(n_61357), .Q(queue
		[125]));
	notech_mux2 i_56149(.S(n_55175), .A(n_3530), .B(queue[125]), .Z(n_42109)
		);
	notech_reg queue_reg_126(.CP(n_62620), .D(n_42115), .CD(n_61357), .Q(queue
		[126]));
	notech_mux2 i_56157(.S(n_55175), .A(n_3536), .B(queue[126]), .Z(n_42115)
		);
	notech_reg queue_reg_127(.CP(n_62620), .D(n_42121), .CD(n_61352), .Q(queue
		[127]));
	notech_mux2 i_56165(.S(n_55175), .A(n_3542), .B(queue[127]), .Z(n_42121)
		);
	notech_and4 i_524983(.A(n_2113), .B(n_2112), .C(n_2107), .D(n_2111), .Z(squeue_4100302
		));
	notech_reg queue_reg_128(.CP(n_62620), .D(n_42127), .CD(n_61352), .Q(queue
		[128]));
	notech_mux2 i_56173(.S(n_55161), .A(n_43043), .B(queue[128]), .Z(n_42127
		));
	notech_nao3 i_19379130(.A(n_58833), .B(queue[100]), .C(n_58612), .Z(n_1036
		));
	notech_reg queue_reg_129(.CP(n_62620), .D(n_42133), .CD(n_61352), .Q(queue
		[129]));
	notech_mux2 i_56181(.S(n_55161), .A(n_43045), .B(queue[129]), .Z(n_42133
		));
	notech_reg queue_reg_130(.CP(n_62620), .D(n_42139), .CD(n_61351), .Q(queue
		[130]));
	notech_mux2 i_56189(.S(n_55161), .A(n_43047), .B(queue[130]), .Z(n_42139
		));
	notech_reg queue_reg_131(.CP(n_62620), .D(n_42145), .CD(n_61351), .Q(queue
		[131]));
	notech_mux2 i_56197(.S(n_55161), .A(n_43049), .B(queue[131]), .Z(n_42145
		));
	notech_reg queue_reg_132(.CP(n_62620), .D(n_42151), .CD(n_61352), .Q(queue
		[132]));
	notech_mux2 i_56205(.S(n_55161), .A(n_43051), .B(queue[132]), .Z(n_42151
		));
	notech_reg queue_reg_133(.CP(n_62620), .D(n_42157), .CD(n_61352), .Q(queue
		[133]));
	notech_mux2 i_56213(.S(n_55161), .A(n_43053), .B(queue[133]), .Z(n_42157
		));
	notech_reg queue_reg_134(.CP(n_62620), .D(n_42163), .CD(n_61352), .Q(queue
		[134]));
	notech_mux2 i_56221(.S(n_55161), .A(n_43055), .B(queue[134]), .Z(n_42163
		));
	notech_reg queue_reg_135(.CP(n_62620), .D(n_42169), .CD(n_61352), .Q(queue
		[135]));
	notech_mux2 i_56229(.S(n_55161), .A(n_43057), .B(queue[135]), .Z(n_42169
		));
	notech_reg queue_reg_136(.CP(n_62620), .D(n_42175), .CD(n_61352), .Q(queue
		[136]));
	notech_mux2 i_56237(.S(n_55161), .A(n_43059), .B(queue[136]), .Z(n_42175
		));
	notech_reg queue_reg_137(.CP(n_62620), .D(n_42181), .CD(n_61351), .Q(queue
		[137]));
	notech_mux2 i_56245(.S(n_55161), .A(n_43061), .B(queue[137]), .Z(n_42181
		));
	notech_reg queue_reg_138(.CP(n_62620), .D(n_42187), .CD(n_61351), .Q(queue
		[138]));
	notech_mux2 i_56253(.S(n_55161), .A(n_43063), .B(queue[138]), .Z(n_42187
		));
	notech_reg queue_reg_139(.CP(n_62620), .D(n_42193), .CD(n_61351), .Q(queue
		[139]));
	notech_mux2 i_56261(.S(n_55161), .A(n_43065), .B(queue[139]), .Z(n_42193
		));
	notech_reg queue_reg_140(.CP(n_62620), .D(n_42199), .CD(n_61351), .Q(queue
		[140]));
	notech_mux2 i_56269(.S(n_55161), .A(n_43067), .B(queue[140]), .Z(n_42199
		));
	notech_reg queue_reg_141(.CP(n_62620), .D(n_42205), .CD(n_61351), .Q(queue
		[141]));
	notech_mux2 i_56277(.S(n_55161), .A(n_43069), .B(queue[141]), .Z(n_42205
		));
	notech_nao3 i_18079143(.A(n_58667), .B(queue[12]), .C(n_58947), .Z(n_1023
		));
	notech_reg queue_reg_142(.CP(n_62620), .D(n_42211), .CD(n_61351), .Q(queue
		[142]));
	notech_mux2 i_56285(.S(n_55161), .A(n_43071), .B(queue[142]), .Z(n_42211
		));
	notech_reg queue_reg_143(.CP(n_62546), .D(n_42217), .CD(n_61351), .Q(queue
		[143]));
	notech_mux2 i_56293(.S(n_55161), .A(n_43073), .B(queue[143]), .Z(n_42217
		));
	notech_reg queue_reg_144(.CP(n_62546), .D(n_42223), .CD(n_61351), .Q(queue
		[144]));
	notech_mux2 i_56301(.S(n_55159), .A(n_43075), .B(queue[144]), .Z(n_42223
		));
	notech_and4 i_424982(.A(n_2099), .B(n_2098), .C(n_2093), .D(n_2097), .Z(squeue_3100303
		));
	notech_reg queue_reg_145(.CP(n_62546), .D(n_42229), .CD(n_61351), .Q(queue
		[145]));
	notech_mux2 i_56309(.S(n_55159), .A(n_43077), .B(queue[145]), .Z(n_42229
		));
	notech_nao3 i_16279161(.A(n_58833), .B(queue[99]), .C(n_58612), .Z(n_1020
		));
	notech_reg queue_reg_146(.CP(n_62546), .D(n_42235), .CD(n_61351), .Q(queue
		[146]));
	notech_mux2 i_56317(.S(n_55159), .A(n_43079), .B(queue[146]), .Z(n_42235
		));
	notech_reg queue_reg_147(.CP(n_62546), .D(n_42241), .CD(n_61351), .Q(queue
		[147]));
	notech_mux2 i_56325(.S(n_55159), .A(n_43081), .B(queue[147]), .Z(n_42241
		));
	notech_reg queue_reg_148(.CP(n_62546), .D(n_42247), .CD(n_61352), .Q(queue
		[148]));
	notech_mux2 i_56333(.S(n_55159), .A(n_43083), .B(queue[148]), .Z(n_42247
		));
	notech_reg queue_reg_149(.CP(n_62546), .D(n_42253), .CD(n_61353), .Q(queue
		[149]));
	notech_mux2 i_56341(.S(n_55159), .A(n_42902), .B(queue[149]), .Z(n_42253
		));
	notech_reg queue_reg_150(.CP(n_62546), .D(n_42259), .CD(n_61353), .Q(queue
		[150]));
	notech_mux2 i_56349(.S(n_55159), .A(n_43086), .B(queue[150]), .Z(n_42259
		));
	notech_reg queue_reg_151(.CP(n_62546), .D(n_42265), .CD(n_61353), .Q(queue
		[151]));
	notech_mux2 i_56357(.S(n_55159), .A(n_43088), .B(queue[151]), .Z(n_42265
		));
	notech_reg queue_reg_152(.CP(n_62546), .D(n_42271), .CD(n_61353), .Q(queue
		[152]));
	notech_mux2 i_56365(.S(n_55159), .A(n_43090), .B(queue[152]), .Z(n_42271
		));
	notech_reg queue_reg_153(.CP(n_62546), .D(n_42277), .CD(n_61353), .Q(queue
		[153]));
	notech_mux2 i_56373(.S(n_55159), .A(n_43092), .B(queue[153]), .Z(n_42277
		));
	notech_reg queue_reg_154(.CP(n_62628), .D(n_42283), .CD(n_61354), .Q(queue
		[154]));
	notech_mux2 i_56381(.S(n_55159), .A(n_43094), .B(queue[154]), .Z(n_42283
		));
	notech_reg queue_reg_155(.CP(clk), .D(n_42289), .CD(n_61354), .Q(queue[
		155]));
	notech_mux2 i_56389(.S(n_55159), .A(n_43096), .B(queue[155]), .Z(n_42289
		));
	notech_reg queue_reg_156(.CP(clk), .D(n_42295), .CD(n_61354), .Q(queue[
		156]));
	notech_mux2 i_56397(.S(n_55159), .A(n_43098), .B(queue[156]), .Z(n_42295
		));
	notech_reg queue_reg_157(.CP(clk), .D(n_42301), .CD(n_61353), .Q(queue[
		157]));
	notech_mux2 i_56405(.S(n_55159), .A(n_43100), .B(queue[157]), .Z(n_42301
		));
	notech_reg queue_reg_158(.CP(clk), .D(n_42307), .CD(n_61354), .Q(queue[
		158]));
	notech_mux2 i_56413(.S(n_55159), .A(n_43102), .B(queue[158]), .Z(n_42307
		));
	notech_nao3 i_14979174(.A(n_58667), .B(queue[11]), .C(n_58947), .Z(n_1007
		));
	notech_reg queue_reg_159(.CP(n_62558), .D(n_42313), .CD(n_61353), .Q(queue
		[159]));
	notech_mux2 i_56421(.S(n_55159), .A(n_43104), .B(queue[159]), .Z(n_42313
		));
	notech_reg queue_reg_160(.CP(n_62558), .D(n_42319), .CD(n_61352), .Q(queue
		[160]));
	notech_mux2 i_56429(.S(n_55166), .A(n_43106), .B(queue[160]), .Z(n_42319
		));
	notech_reg queue_reg_161(.CP(n_62558), .D(n_42325), .CD(n_61353), .Q(queue
		[161]));
	notech_mux2 i_56437(.S(n_55166), .A(n_43108), .B(queue[161]), .Z(n_42325
		));
	notech_and4 i_324981(.A(n_2085), .B(n_2084), .C(n_2079), .D(n_2083), .Z(squeue_2100304
		));
	notech_reg queue_reg_162(.CP(n_62558), .D(n_42331), .CD(n_61352), .Q(queue
		[162]));
	notech_mux2 i_56445(.S(n_55166), .A(n_43110), .B(queue[162]), .Z(n_42331
		));
	notech_nao3 i_13179192(.A(n_58837), .B(queue[98]), .C(n_58609), .Z(n_1004
		));
	notech_reg queue_reg_163(.CP(n_62558), .D(n_42337), .CD(n_61352), .Q(queue
		[163]));
	notech_mux2 i_56453(.S(n_55166), .A(n_43112), .B(queue[163]), .Z(n_42337
		));
	notech_reg queue_reg_164(.CP(n_62558), .D(n_42343), .CD(n_61352), .Q(queue
		[164]));
	notech_mux2 i_56461(.S(n_55166), .A(n_43114), .B(queue[164]), .Z(n_42343
		));
	notech_reg queue_reg_165(.CP(n_62558), .D(n_42349), .CD(n_61353), .Q(queue
		[165]));
	notech_mux2 i_56469(.S(n_55166), .A(n_43116), .B(queue[165]), .Z(n_42349
		));
	notech_reg queue_reg_166(.CP(n_62558), .D(n_42355), .CD(n_61353), .Q(queue
		[166]));
	notech_mux2 i_56477(.S(n_55166), .A(n_43118), .B(queue[166]), .Z(n_42355
		));
	notech_reg queue_reg_167(.CP(n_62558), .D(n_42361), .CD(n_61353), .Q(queue
		[167]));
	notech_mux2 i_56485(.S(n_55166), .A(n_43120), .B(queue[167]), .Z(n_42361
		));
	notech_reg queue_reg_168(.CP(n_62558), .D(n_42367), .CD(n_61353), .Q(queue
		[168]));
	notech_mux2 i_56493(.S(n_55166), .A(n_43122), .B(queue[168]), .Z(n_42367
		));
	notech_reg queue_reg_169(.CP(n_62558), .D(n_42373), .CD(n_61353), .Q(queue
		[169]));
	notech_mux2 i_56501(.S(n_55166), .A(n_43124), .B(queue[169]), .Z(n_42373
		));
	notech_reg queue_reg_170(.CP(n_62558), .D(n_42379), .CD(n_61363), .Q(queue
		[170]));
	notech_mux2 i_56509(.S(n_55166), .A(n_43126), .B(queue[170]), .Z(n_42379
		));
	notech_reg queue_reg_171(.CP(n_62558), .D(n_42385), .CD(n_61363), .Q(queue
		[171]));
	notech_mux2 i_56517(.S(n_55166), .A(n_43128), .B(queue[171]), .Z(n_42385
		));
	notech_reg queue_reg_172(.CP(n_62558), .D(n_42391), .CD(n_61363), .Q(queue
		[172]));
	notech_mux2 i_56525(.S(n_55166), .A(n_43130), .B(queue[172]), .Z(n_42391
		));
	notech_reg queue_reg_173(.CP(n_62558), .D(n_42397), .CD(n_61363), .Q(queue
		[173]));
	notech_mux2 i_56533(.S(n_55166), .A(n_43132), .B(queue[173]), .Z(n_42397
		));
	notech_reg queue_reg_174(.CP(n_62558), .D(n_42403), .CD(n_61363), .Q(queue
		[174]));
	notech_mux2 i_56541(.S(n_55166), .A(n_43134), .B(queue[174]), .Z(n_42403
		));
	notech_reg queue_reg_175(.CP(n_62558), .D(n_42409), .CD(n_61363), .Q(queue
		[175]));
	notech_mux2 i_56549(.S(n_55166), .A(n_43136), .B(queue[175]), .Z(n_42409
		));
	notech_nao3 i_11879205(.A(n_58667), .B(queue[10]), .C(n_58947), .Z(n_991
		));
	notech_reg queue_reg_176(.CP(n_62558), .D(n_42415), .CD(n_61364), .Q(queue
		[176]));
	notech_mux2 i_56557(.S(n_55164), .A(n_43138), .B(queue[176]), .Z(n_42415
		));
	notech_reg queue_reg_177(.CP(n_62558), .D(n_42421), .CD(n_61363), .Q(queue
		[177]));
	notech_mux2 i_56565(.S(n_55164), .A(n_43140), .B(queue[177]), .Z(n_42421
		));
	notech_reg queue_reg_178(.CP(n_62632), .D(n_42427), .CD(n_61363), .Q(queue
		[178]));
	notech_mux2 i_56573(.S(n_55164), .A(n_43142), .B(queue[178]), .Z(n_42427
		));
	notech_and4 i_224980(.A(n_2071), .B(n_2070), .C(n_2065), .D(n_2069), .Z(squeue_1100305
		));
	notech_reg queue_reg_179(.CP(n_62556), .D(n_42433), .CD(n_61363), .Q(queue
		[179]));
	notech_mux2 i_56581(.S(n_55164), .A(n_42901), .B(queue[179]), .Z(n_42433
		));
	notech_nao3 i_10079223(.A(n_58837), .B(queue[97]), .C(n_58612), .Z(n_988
		));
	notech_reg queue_reg_180(.CP(n_62632), .D(n_42439), .CD(n_61363), .Q(queue
		[180]));
	notech_mux2 i_56589(.S(n_55164), .A(n_43145), .B(queue[180]), .Z(n_42439
		));
	notech_reg queue_reg_181(.CP(n_62632), .D(n_42445), .CD(n_61361), .Q(queue
		[181]));
	notech_mux2 i_56597(.S(n_55164), .A(n_43147), .B(queue[181]), .Z(n_42445
		));
	notech_reg queue_reg_182(.CP(n_62632), .D(n_42451), .CD(n_61361), .Q(queue
		[182]));
	notech_mux2 i_56605(.S(n_55164), .A(n_43149), .B(queue[182]), .Z(n_42451
		));
	notech_reg queue_reg_183(.CP(n_62632), .D(n_42457), .CD(n_61361), .Q(queue
		[183]));
	notech_mux2 i_56613(.S(n_55164), .A(n_43151), .B(queue[183]), .Z(n_42457
		));
	notech_reg queue_reg_184(.CP(n_62632), .D(n_42463), .CD(n_61361), .Q(queue
		[184]));
	notech_mux2 i_56621(.S(n_55164), .A(n_43153), .B(queue[184]), .Z(n_42463
		));
	notech_reg queue_reg_185(.CP(n_62632), .D(n_42469), .CD(n_61361), .Q(queue
		[185]));
	notech_mux2 i_56629(.S(n_55164), .A(n_43155), .B(queue[185]), .Z(n_42469
		));
	notech_reg queue_reg_186(.CP(n_62632), .D(n_42475), .CD(n_61363), .Q(queue
		[186]));
	notech_mux2 i_56637(.S(n_55164), .A(n_43157), .B(queue[186]), .Z(n_42475
		));
	notech_reg queue_reg_187(.CP(n_62632), .D(n_42481), .CD(n_61363), .Q(queue
		[187]));
	notech_mux2 i_56645(.S(n_55164), .A(n_43159), .B(queue[187]), .Z(n_42481
		));
	notech_reg queue_reg_188(.CP(n_62632), .D(n_42487), .CD(n_61363), .Q(queue
		[188]));
	notech_mux2 i_56653(.S(n_55164), .A(n_43161), .B(queue[188]), .Z(n_42487
		));
	notech_reg queue_reg_189(.CP(n_62632), .D(n_42493), .CD(n_61361), .Q(queue
		[189]));
	notech_mux2 i_56661(.S(n_55164), .A(n_43163), .B(queue[189]), .Z(n_42493
		));
	notech_reg queue_reg_190(.CP(n_62632), .D(n_42499), .CD(n_61363), .Q(queue
		[190]));
	notech_mux2 i_56669(.S(n_55164), .A(n_43165), .B(queue[190]), .Z(n_42499
		));
	notech_reg queue_reg_191(.CP(n_62632), .D(n_42505), .CD(n_61364), .Q(queue
		[191]));
	notech_mux2 i_56677(.S(n_55164), .A(n_43167), .B(queue[191]), .Z(n_42505
		));
	notech_reg queue_reg_192(.CP(n_62632), .D(n_42511), .CD(n_61365), .Q(queue
		[192]));
	notech_mux2 i_56685(.S(n_55151), .A(n_43169), .B(queue[192]), .Z(n_42511
		));
	notech_nao3 i_8779236(.A(n_58667), .B(queue[9]), .C(n_58947), .Z(n_975)
		);
	notech_reg queue_reg_193(.CP(n_62632), .D(n_42517), .CD(n_61365), .Q(queue
		[193]));
	notech_mux2 i_56693(.S(n_55151), .A(n_43171), .B(queue[193]), .Z(n_42517
		));
	notech_reg queue_reg_194(.CP(n_62632), .D(n_42523), .CD(n_61365), .Q(queue
		[194]));
	notech_mux2 i_56701(.S(n_55151), .A(n_43173), .B(queue[194]), .Z(n_42523
		));
	notech_reg queue_reg_195(.CP(n_62632), .D(n_42529), .CD(n_61364), .Q(queue
		[195]));
	notech_mux2 i_56709(.S(n_55151), .A(n_43175), .B(queue[195]), .Z(n_42529
		));
	notech_and4 i_124979(.A(n_2057), .B(n_2056), .C(n_2050), .D(n_2055), .Z(squeue_0100306
		));
	notech_reg queue_reg_196(.CP(n_62632), .D(n_42535), .CD(n_61365), .Q(queue
		[196]));
	notech_mux2 i_56717(.S(n_55151), .A(n_43177), .B(queue[196]), .Z(n_42535
		));
	notech_nao3 i_6379254(.A(n_58833), .B(queue[96]), .C(n_58612), .Z(n_972)
		);
	notech_reg queue_reg_197(.CP(n_62632), .D(n_42541), .CD(n_61365), .Q(queue
		[197]));
	notech_mux2 i_56725(.S(n_55151), .A(n_43179), .B(queue[197]), .Z(n_42541
		));
	notech_reg queue_reg_198(.CP(n_62556), .D(n_42547), .CD(n_61365), .Q(queue
		[198]));
	notech_mux2 i_56733(.S(n_55151), .A(n_43181), .B(queue[198]), .Z(n_42547
		));
	notech_reg queue_reg_199(.CP(n_62556), .D(n_42553), .CD(n_61365), .Q(queue
		[199]));
	notech_mux2 i_56741(.S(n_55151), .A(n_43183), .B(queue[199]), .Z(n_42553
		));
	notech_reg queue_reg_200(.CP(n_62556), .D(n_42559), .CD(n_61365), .Q(queue
		[200]));
	notech_mux2 i_56749(.S(n_55151), .A(n_43185), .B(queue[200]), .Z(n_42559
		));
	notech_reg queue_reg_201(.CP(n_62556), .D(n_42565), .CD(n_61365), .Q(queue
		[201]));
	notech_mux2 i_56757(.S(n_55151), .A(n_43187), .B(queue[201]), .Z(n_42565
		));
	notech_reg queue_reg_202(.CP(n_62556), .D(n_42571), .CD(n_61364), .Q(queue
		[202]));
	notech_mux2 i_56765(.S(n_55151), .A(n_43189), .B(queue[202]), .Z(n_42571
		));
	notech_reg queue_reg_203(.CP(n_62556), .D(n_42577), .CD(n_61364), .Q(queue
		[203]));
	notech_mux2 i_56773(.S(n_55151), .A(n_43191), .B(queue[203]), .Z(n_42577
		));
	notech_reg queue_reg_204(.CP(clk), .D(n_42583), .CD(n_61364), .Q(queue[
		204]));
	notech_mux2 i_56781(.S(n_55151), .A(n_43193), .B(queue[204]), .Z(n_42583
		));
	notech_reg queue_reg_205(.CP(n_62554), .D(n_42589), .CD(n_61364), .Q(queue
		[205]));
	notech_mux2 i_56789(.S(n_55151), .A(n_43195), .B(queue[205]), .Z(n_42589
		));
	notech_reg queue_reg_206(.CP(n_62628), .D(n_42595), .CD(n_61364), .Q(queue
		[206]));
	notech_mux2 i_56797(.S(n_55151), .A(n_43197), .B(queue[206]), .Z(n_42595
		));
	notech_reg queue_reg_207(.CP(n_62628), .D(n_42601), .CD(n_61364), .Q(queue
		[207]));
	notech_mux2 i_56805(.S(n_55151), .A(n_43199), .B(queue[207]), .Z(n_42601
		));
	notech_reg queue_reg_208(.CP(n_62628), .D(n_42607), .CD(n_61364), .Q(queue
		[208]));
	notech_mux2 i_56813(.S(n_55149), .A(n_42900), .B(queue[208]), .Z(n_42607
		));
	notech_reg queue_reg_209(.CP(n_62628), .D(n_42613), .CD(n_61364), .Q(queue
		[209]));
	notech_mux2 i_56821(.S(n_55149), .A(n_43202), .B(queue[209]), .Z(n_42613
		));
	notech_nao3 i_5079267(.A(n_58667), .B(queue[8]), .C(n_58947), .Z(n_959)
		);
	notech_reg queue_reg_210(.CP(n_62628), .D(n_42619), .CD(n_61364), .Q(queue
		[210]));
	notech_mux2 i_56829(.S(n_55149), .A(n_43204), .B(queue[210]), .Z(n_42619
		));
	notech_reg queue_reg_211(.CP(n_62704), .D(n_42625), .CD(n_61364), .Q(queue
		[211]));
	notech_mux2 i_56837(.S(n_55149), .A(n_43206), .B(queue[211]), .Z(n_42625
		));
	notech_reg queue_reg_212(.CP(n_62704), .D(n_42631), .CD(n_61364), .Q(queue
		[212]));
	notech_mux2 i_56845(.S(n_55149), .A(n_43208), .B(queue[212]), .Z(n_42631
		));
	notech_or4 i_175279354(.A(n_42908), .B(n_955), .C(n_956), .D(n_42896), .Z
		(\nbus_94[0] ));
	notech_reg queue_reg_213(.CP(n_62704), .D(n_42637), .CD(n_61359), .Q(queue
		[213]));
	notech_mux2 i_56853(.S(n_55149), .A(n_43210), .B(queue[213]), .Z(n_42637
		));
	notech_ao3 i_4379274(.A(pg_fault), .B(n_60413), .C(n_2946), .Z(n_956));
	notech_reg queue_reg_214(.CP(n_62704), .D(n_42643), .CD(n_61359), .Q(queue
		[214]));
	notech_mux2 i_56861(.S(n_55149), .A(n_43212), .B(queue[214]), .Z(n_42643
		));
	notech_and3 i_4179275(.A(n_2037), .B(n_2951), .C(n_8137), .Z(n_955));
	notech_reg queue_reg_215(.CP(n_62704), .D(n_42649), .CD(n_61359), .Q(queue
		[215]));
	notech_mux2 i_56869(.S(n_55149), .A(n_43214), .B(queue[215]), .Z(n_42649
		));
	notech_or4 i_7279318(.A(n_60778), .B(n_42907), .C(n_42897), .D(n_43489),
		 .Z(n_8130));
	notech_reg queue_reg_216(.CP(n_62704), .D(n_42655), .CD(n_61359), .Q(queue
		[216]));
	notech_mux2 i_56877(.S(n_55149), .A(n_43216), .B(queue[216]), .Z(n_42655
		));
	notech_nor2 i_6579316(.A(n_60790), .B(n_2946), .Z(n_8137));
	notech_reg queue_reg_217(.CP(n_62704), .D(n_42661), .CD(n_61359), .Q(queue
		[217]));
	notech_mux2 i_56885(.S(n_55149), .A(n_43218), .B(queue[217]), .Z(n_42661
		));
	notech_reg queue_reg_218(.CP(n_62704), .D(n_42667), .CD(n_61359), .Q(queue
		[218]));
	notech_mux2 i_56893(.S(n_55149), .A(n_43220), .B(queue[218]), .Z(n_42667
		));
	notech_reg queue_reg_219(.CP(n_62704), .D(n_42673), .CD(n_61359), .Q(queue
		[219]));
	notech_mux2 i_56901(.S(n_55149), .A(n_43222), .B(queue[219]), .Z(n_42673
		));
	notech_ao4 i_3579279(.A(n_140854113), .B(n_2038), .C(n_2997), .D(n_60596
		), .Z(n_951));
	notech_reg queue_reg_220(.CP(n_62704), .D(n_42679), .CD(n_61359), .Q(queue
		[220]));
	notech_mux2 i_56909(.S(n_55149), .A(n_43224), .B(queue[220]), .Z(n_42679
		));
	notech_or2 i_6979317(.A(fault_wptr[1]), .B(fault_wptr[0]), .Z(n_8133));
	notech_reg queue_reg_221(.CP(n_62704), .D(n_42685), .CD(n_61359), .Q(queue
		[221]));
	notech_mux2 i_56917(.S(n_55149), .A(n_43226), .B(queue[221]), .Z(n_42685
		));
	notech_nand2 i_5430(.A(n_43481), .B(n_43482), .Z(n_950));
	notech_reg queue_reg_222(.CP(n_62704), .D(n_42691), .CD(n_61359), .Q(queue
		[222]));
	notech_mux2 i_56925(.S(n_55149), .A(n_43228), .B(queue[222]), .Z(n_42691
		));
	notech_or4 i_7655(.A(tagV[1]), .B(tagV[0]), .C(tagV[3]), .D(n_2035), .Z(n_8629
		));
	notech_reg queue_reg_223(.CP(n_62704), .D(n_42697), .CD(n_61359), .Q(queue
		[223]));
	notech_mux2 i_56933(.S(n_55149), .A(n_43230), .B(queue[223]), .Z(n_42697
		));
	notech_nand2 i_43979398(.A(addrshft[4]), .B(n_43301), .Z(n_949));
	notech_reg queue_reg_224(.CP(n_62704), .D(n_42703), .CD(n_61358), .Q(queue
		[224]));
	notech_mux2 i_56941(.S(n_55156), .A(n_43232), .B(queue[224]), .Z(n_42703
		));
	notech_nand3 i_6279805(.A(wptr[0]), .B(n_42914), .C(n_2908), .Z(n_948)
		);
	notech_reg queue_reg_225(.CP(n_62704), .D(n_42709), .CD(n_61358), .Q(queue
		[225]));
	notech_mux2 i_56949(.S(n_55156), .A(n_43234), .B(queue[225]), .Z(n_42709
		));
	notech_reg queue_reg_226(.CP(n_62704), .D(n_42715), .CD(n_61358), .Q(queue
		[226]));
	notech_mux2 i_56957(.S(n_55156), .A(n_43236), .B(queue[226]), .Z(n_42715
		));
	notech_reg queue_reg_227(.CP(n_62704), .D(n_42721), .CD(n_61358), .Q(queue
		[227]));
	notech_mux2 i_56965(.S(n_55156), .A(n_43238), .B(queue[227]), .Z(n_42721
		));
	notech_nand2 i_44679391(.A(n_2396), .B(n_43488), .Z(n_945));
	notech_reg queue_reg_228(.CP(n_62704), .D(n_42727), .CD(n_61358), .Q(queue
		[228]));
	notech_mux2 i_56973(.S(n_55156), .A(n_43240), .B(queue[228]), .Z(n_42727
		));
	notech_nao3 i_44879389(.A(n_8629), .B(n_60413), .C(pg_fault), .Z(n_944)
		);
	notech_reg queue_reg_229(.CP(n_62628), .D(n_42733), .CD(n_61359), .Q(queue
		[229]));
	notech_mux2 i_56981(.S(n_55156), .A(n_43242), .B(queue[229]), .Z(n_42733
		));
	notech_reg queue_reg_230(.CP(n_62704), .D(n_42739), .CD(n_61359), .Q(queue
		[230]));
	notech_mux2 i_56989(.S(n_55156), .A(n_43244), .B(queue[230]), .Z(n_42739
		));
	notech_ao4 i_3379802(.A(n_2033), .B(n_43489), .C(n_60778), .D(n_2947), .Z
		(n_942));
	notech_reg queue_reg_231(.CP(n_62630), .D(n_42745), .CD(n_61359), .Q(queue
		[231]));
	notech_mux2 i_56997(.S(n_55156), .A(n_43246), .B(queue[231]), .Z(n_42745
		));
	notech_nao3 i_26879569(.A(n_2396), .B(n_8137), .C(n_8629), .Z(n_941));
	notech_reg queue_reg_232(.CP(n_62630), .D(n_42751), .CD(n_61358), .Q(queue
		[232]));
	notech_mux2 i_57005(.S(n_55156), .A(n_43248), .B(queue[232]), .Z(n_42751
		));
	notech_reg queue_reg_233(.CP(n_62630), .D(n_42757), .CD(n_61358), .Q(queue
		[233]));
	notech_mux2 i_57013(.S(n_55156), .A(n_43250), .B(queue[233]), .Z(n_42757
		));
	notech_reg queue_reg_234(.CP(n_62630), .D(n_42763), .CD(n_61360), .Q(queue
		[234]));
	notech_mux2 i_57021(.S(n_55156), .A(n_43252), .B(queue[234]), .Z(n_42763
		));
	notech_ao4 i_3679799(.A(n_60596), .B(n_2997), .C(n_945), .D(n_944), .Z(n_938
		));
	notech_reg queue_reg_235(.CP(n_62630), .D(n_42769), .CD(n_61361), .Q(queue
		[235]));
	notech_mux2 i_57029(.S(n_55156), .A(n_43254), .B(queue[235]), .Z(n_42769
		));
	notech_or2 i_27179566(.A(n_938), .B(n_2946), .Z(n_937));
	notech_reg queue_reg_236(.CP(n_62630), .D(n_42775), .CD(n_61361), .Q(queue
		[236]));
	notech_mux2 i_57037(.S(n_55156), .A(n_43256), .B(queue[236]), .Z(n_42775
		));
	notech_reg queue_reg_237(.CP(n_62630), .D(n_42781), .CD(n_61361), .Q(queue
		[237]));
	notech_mux2 i_57045(.S(n_55156), .A(n_43258), .B(queue[237]), .Z(n_42781
		));
	notech_xor2 i_3979797(.A(n_43296), .B(addrshft[1]), .Z(n_935));
	notech_reg queue_reg_238(.CP(n_62630), .D(n_42787), .CD(n_61360), .Q(queue
		[238]));
	notech_mux2 i_57053(.S(n_55156), .A(n_43260), .B(queue[238]), .Z(n_42787
		));
	notech_reg queue_reg_239(.CP(n_62630), .D(n_42793), .CD(n_61360), .Q(queue
		[239]));
	notech_mux2 i_57061(.S(n_55156), .A(n_43262), .B(queue[239]), .Z(n_42793
		));
	notech_reg queue_reg_240(.CP(n_62630), .D(n_42799), .CD(n_61361), .Q(queue
		[240]));
	notech_mux2 i_57069(.S(n_55154), .A(n_43264), .B(queue[240]), .Z(n_42799
		));
	notech_reg queue_reg_241(.CP(n_62630), .D(n_42805), .CD(n_61361), .Q(queue
		[241]));
	notech_mux2 i_57077(.S(n_55154), .A(n_43266), .B(queue[241]), .Z(n_42805
		));
	notech_reg queue_reg_242(.CP(n_62630), .D(n_42811), .CD(n_61361), .Q(queue
		[242]));
	notech_mux2 i_57085(.S(n_55154), .A(n_43268), .B(queue[242]), .Z(n_42811
		));
	notech_xor2 i_4079796(.A(addrshft[2]), .B(n_2887), .Z(n_930));
	notech_reg queue_reg_243(.CP(n_62630), .D(n_42817), .CD(n_61361), .Q(queue
		[243]));
	notech_mux2 i_57093(.S(n_55154), .A(n_43270), .B(queue[243]), .Z(n_42817
		));
	notech_reg queue_reg_244(.CP(n_62630), .D(n_42823), .CD(n_61361), .Q(queue
		[244]));
	notech_mux2 i_57101(.S(n_55154), .A(n_43272), .B(queue[244]), .Z(n_42823
		));
	notech_reg queue_reg_245(.CP(n_62630), .D(n_42829), .CD(n_61360), .Q(queue
		[245]));
	notech_mux2 i_57109(.S(n_55154), .A(n_43274), .B(queue[245]), .Z(n_42829
		));
	notech_reg queue_reg_246(.CP(n_62630), .D(n_42835), .CD(n_61360), .Q(queue
		[246]));
	notech_mux2 i_57117(.S(n_55154), .A(n_43276), .B(queue[246]), .Z(n_42835
		));
	notech_reg queue_reg_247(.CP(n_62630), .D(n_42841), .CD(n_61360), .Q(queue
		[247]));
	notech_mux2 i_57125(.S(n_55154), .A(n_43278), .B(queue[247]), .Z(n_42841
		));
	notech_reg queue_reg_248(.CP(n_62630), .D(n_42847), .CD(n_61360), .Q(queue
		[248]));
	notech_mux2 i_57133(.S(n_55154), .A(n_43280), .B(queue[248]), .Z(n_42847
		));
	notech_ao4 i_4279794(.A(addrshft[4]), .B(n_43301), .C(n_949), .D(n_42904
		), .Z(n_924));
	notech_reg queue_reg_249(.CP(n_62630), .D(n_42853), .CD(n_61360), .Q(queue
		[249]));
	notech_mux2 i_57141(.S(n_55154), .A(n_43282), .B(queue[249]), .Z(n_42853
		));
	notech_reg queue_reg_250(.CP(n_62554), .D(n_42859), .CD(n_61360), .Q(queue
		[250]));
	notech_mux2 i_57149(.S(n_55154), .A(n_43284), .B(queue[250]), .Z(n_42859
		));
	notech_reg queue_reg_251(.CP(n_62554), .D(n_42865), .CD(n_61360), .Q(queue
		[251]));
	notech_mux2 i_57157(.S(n_55154), .A(n_43286), .B(queue[251]), .Z(n_42865
		));
	notech_reg queue_reg_252(.CP(n_62554), .D(n_42871), .CD(n_61360), .Q(queue
		[252]));
	notech_mux2 i_57165(.S(n_55154), .A(n_43288), .B(queue[252]), .Z(n_42871
		));
	notech_ao4 i_4479792(.A(n_60750), .B(n_141554120), .C(n_2944), .D(n_43481
		), .Z(n_920));
	notech_reg queue_reg_253(.CP(n_62554), .D(n_42877), .CD(n_61360), .Q(queue
		[253]));
	notech_mux2 i_57173(.S(n_55154), .A(n_43290), .B(queue[253]), .Z(n_42877
		));
	notech_reg queue_reg_254(.CP(clk), .D(n_42883), .CD(n_61360), .Q(queue[
		254]));
	notech_mux2 i_57181(.S(n_55154), .A(n_43292), .B(queue[254]), .Z(n_42883
		));
	notech_reg queue_reg_255(.CP(n_62554), .D(n_42889), .CD(n_61360), .Q(queue
		[255]));
	notech_mux2 i_57189(.S(n_55154), .A(n_43294), .B(queue[255]), .Z(n_42889
		));
	notech_inv i_60228(.A(n_2915), .Z(n_42895));
	notech_inv i_60229(.A(n_2950), .Z(n_42896));
	notech_inv i_60230(.A(n_2995), .Z(n_42897));
	notech_inv i_60231(.A(n_2944), .Z(n_42898));
	notech_inv i_60232(.A(n_58822), .Z(n_42899));
	notech_inv i_60233(.A(n_3781), .Z(n_42900));
	notech_inv i_60234(.A(n_378299582), .Z(n_42901));
	notech_inv i_60235(.A(n_3783), .Z(n_42902));
	notech_inv i_60236(.A(n_8629), .Z(n_42903));
	notech_inv i_60237(.A(n_28556624), .Z(n_42904));
	notech_inv i_60240(.A(n_2947), .Z(n_42907));
	notech_inv i_60241(.A(n_8130), .Z(n_42908));
	notech_inv i_60242(.A(n_60778), .Z(cacheD[148]));
	notech_inv i_60243(.A(fault_wptr_en), .Z(n_42910));
	notech_inv i_60244(.A(n_2743), .Z(n_42911));
	notech_inv i_60245(.A(n_4675), .Z(n_42912));
	notech_inv i_60246(.A(wptr[0]), .Z(n_42913));
	notech_inv i_60247(.A(wptr[1]), .Z(n_42914));
	notech_inv i_60248(.A(n_2730), .Z(n_42915));
	notech_inv i_60249(.A(n_2736), .Z(n_42916));
	notech_inv i_60250(.A(queue[0]), .Z(n_42917));
	notech_inv i_60251(.A(queue[1]), .Z(n_42918));
	notech_inv i_60252(.A(queue[2]), .Z(n_42919));
	notech_inv i_60253(.A(queue[3]), .Z(n_42920));
	notech_inv i_60254(.A(queue[4]), .Z(n_42921));
	notech_inv i_60255(.A(queue[5]), .Z(n_42922));
	notech_inv i_60256(.A(queue[6]), .Z(n_42923));
	notech_inv i_60257(.A(queue[7]), .Z(n_42924));
	notech_inv i_60258(.A(queue[9]), .Z(n_42925));
	notech_inv i_60259(.A(queue[10]), .Z(n_42926));
	notech_inv i_60260(.A(queue[11]), .Z(n_42927));
	notech_inv i_60261(.A(queue[12]), .Z(n_42928));
	notech_inv i_60262(.A(queue[13]), .Z(n_42929));
	notech_inv i_60263(.A(queue[15]), .Z(n_42930));
	notech_inv i_60264(.A(queue[16]), .Z(n_42931));
	notech_inv i_60265(.A(queue[17]), .Z(n_42932));
	notech_inv i_60266(.A(queue[18]), .Z(n_42933));
	notech_inv i_60267(.A(queue[19]), .Z(n_42934));
	notech_inv i_60268(.A(queue[20]), .Z(n_42935));
	notech_inv i_60269(.A(queue[21]), .Z(n_42936));
	notech_inv i_60270(.A(queue[22]), .Z(n_42937));
	notech_inv i_60271(.A(queue[23]), .Z(n_42938));
	notech_inv i_60272(.A(queue[24]), .Z(n_42939));
	notech_inv i_60273(.A(queue[25]), .Z(n_42940));
	notech_inv i_60274(.A(queue[26]), .Z(n_42941));
	notech_inv i_60275(.A(queue[27]), .Z(n_42942));
	notech_inv i_60276(.A(queue[28]), .Z(n_42943));
	notech_inv i_60277(.A(queue[29]), .Z(n_42944));
	notech_inv i_60278(.A(queue[30]), .Z(n_42945));
	notech_inv i_60279(.A(queue[31]), .Z(n_42946));
	notech_inv i_60280(.A(queue[32]), .Z(n_42947));
	notech_inv i_60281(.A(queue[33]), .Z(n_42948));
	notech_inv i_60282(.A(queue[34]), .Z(n_42949));
	notech_inv i_60283(.A(queue[35]), .Z(n_42950));
	notech_inv i_60284(.A(queue[36]), .Z(n_42951));
	notech_inv i_60285(.A(queue[37]), .Z(n_42952));
	notech_inv i_60286(.A(queue[38]), .Z(n_42953));
	notech_inv i_60287(.A(queue[39]), .Z(n_42954));
	notech_inv i_60288(.A(queue[40]), .Z(n_42955));
	notech_inv i_60289(.A(queue[41]), .Z(n_42956));
	notech_inv i_60290(.A(queue[42]), .Z(n_42957));
	notech_inv i_60291(.A(queue[43]), .Z(n_42958));
	notech_inv i_60292(.A(queue[44]), .Z(n_42959));
	notech_inv i_60293(.A(queue[45]), .Z(n_42960));
	notech_inv i_60294(.A(queue[46]), .Z(n_42961));
	notech_inv i_60295(.A(queue[47]), .Z(n_42962));
	notech_inv i_60296(.A(queue[48]), .Z(n_42963));
	notech_inv i_60297(.A(queue[49]), .Z(n_42964));
	notech_inv i_60298(.A(queue[50]), .Z(n_42965));
	notech_inv i_60299(.A(queue[51]), .Z(n_42966));
	notech_inv i_60300(.A(queue[52]), .Z(n_42967));
	notech_inv i_60301(.A(queue[53]), .Z(n_42968));
	notech_inv i_60302(.A(queue[54]), .Z(n_42969));
	notech_inv i_60303(.A(queue[55]), .Z(n_42970));
	notech_inv i_60304(.A(queue[56]), .Z(n_42971));
	notech_inv i_60305(.A(queue[57]), .Z(n_42972));
	notech_inv i_60306(.A(queue[58]), .Z(n_42973));
	notech_inv i_60307(.A(queue[59]), .Z(n_42974));
	notech_inv i_60308(.A(queue[60]), .Z(n_42975));
	notech_inv i_60309(.A(queue[61]), .Z(n_42976));
	notech_inv i_60310(.A(queue[62]), .Z(n_42977));
	notech_inv i_60311(.A(queue[63]), .Z(n_42978));
	notech_inv i_60312(.A(queue[64]), .Z(n_42979));
	notech_inv i_60313(.A(queue[65]), .Z(n_42980));
	notech_inv i_60314(.A(queue[66]), .Z(n_42981));
	notech_inv i_60315(.A(queue[67]), .Z(n_42982));
	notech_inv i_60316(.A(queue[68]), .Z(n_42983));
	notech_inv i_60317(.A(queue[69]), .Z(n_42984));
	notech_inv i_60318(.A(queue[70]), .Z(n_42985));
	notech_inv i_60319(.A(queue[71]), .Z(n_42986));
	notech_inv i_60320(.A(queue[72]), .Z(n_42987));
	notech_inv i_60321(.A(queue[73]), .Z(n_42988));
	notech_inv i_60322(.A(queue[74]), .Z(n_42989));
	notech_inv i_60323(.A(queue[75]), .Z(n_42990));
	notech_inv i_60324(.A(queue[76]), .Z(n_42991));
	notech_inv i_60325(.A(queue[77]), .Z(n_42992));
	notech_inv i_60326(.A(queue[78]), .Z(n_42993));
	notech_inv i_60327(.A(queue[79]), .Z(n_42994));
	notech_inv i_60328(.A(queue[80]), .Z(n_42995));
	notech_inv i_60329(.A(queue[81]), .Z(n_42996));
	notech_inv i_60330(.A(queue[82]), .Z(n_42997));
	notech_inv i_60331(.A(queue[83]), .Z(n_42998));
	notech_inv i_60332(.A(queue[84]), .Z(n_42999));
	notech_inv i_60333(.A(queue[85]), .Z(n_43000));
	notech_inv i_60334(.A(queue[86]), .Z(n_43001));
	notech_inv i_60335(.A(queue[87]), .Z(n_43002));
	notech_inv i_60336(.A(queue[88]), .Z(n_43003));
	notech_inv i_60337(.A(queue[89]), .Z(n_43004));
	notech_inv i_60338(.A(queue[90]), .Z(n_43005));
	notech_inv i_60339(.A(queue[91]), .Z(n_43006));
	notech_inv i_60340(.A(queue[92]), .Z(n_43007));
	notech_inv i_60341(.A(queue[93]), .Z(n_43008));
	notech_inv i_60342(.A(queue[94]), .Z(n_43009));
	notech_inv i_60343(.A(queue[95]), .Z(n_43010));
	notech_inv i_60344(.A(queue[96]), .Z(n_43011));
	notech_inv i_60345(.A(queue[97]), .Z(n_43012));
	notech_inv i_60346(.A(queue[98]), .Z(n_43013));
	notech_inv i_60347(.A(queue[99]), .Z(n_43014));
	notech_inv i_60348(.A(queue[100]), .Z(n_43015));
	notech_inv i_60349(.A(queue[101]), .Z(n_43016));
	notech_inv i_60350(.A(queue[102]), .Z(n_43017));
	notech_inv i_60351(.A(queue[103]), .Z(n_43018));
	notech_inv i_60352(.A(queue[104]), .Z(n_43019));
	notech_inv i_60353(.A(queue[105]), .Z(n_43020));
	notech_inv i_60354(.A(queue[106]), .Z(n_43021));
	notech_inv i_60355(.A(queue[107]), .Z(n_43022));
	notech_inv i_60356(.A(queue[108]), .Z(n_43023));
	notech_inv i_60357(.A(queue[109]), .Z(n_43024));
	notech_inv i_60358(.A(queue[110]), .Z(n_43025));
	notech_inv i_60359(.A(queue[111]), .Z(n_43026));
	notech_inv i_60360(.A(queue[112]), .Z(n_43027));
	notech_inv i_60361(.A(queue[113]), .Z(n_43028));
	notech_inv i_60362(.A(queue[114]), .Z(n_43029));
	notech_inv i_60363(.A(queue[115]), .Z(n_43030));
	notech_inv i_60364(.A(queue[116]), .Z(n_43031));
	notech_inv i_60365(.A(queue[117]), .Z(n_43032));
	notech_inv i_60366(.A(queue[118]), .Z(n_43033));
	notech_inv i_60367(.A(queue[119]), .Z(n_43034));
	notech_inv i_60368(.A(queue[120]), .Z(n_43035));
	notech_inv i_60369(.A(queue[121]), .Z(n_43036));
	notech_inv i_60370(.A(queue[122]), .Z(n_43037));
	notech_inv i_60371(.A(queue[123]), .Z(n_43038));
	notech_inv i_60372(.A(queue[124]), .Z(n_43039));
	notech_inv i_60373(.A(queue[125]), .Z(n_43040));
	notech_inv i_60374(.A(queue[126]), .Z(n_43041));
	notech_inv i_60375(.A(queue[127]), .Z(n_43042));
	notech_inv i_60376(.A(n_3548), .Z(n_43043));
	notech_inv i_60377(.A(queue[128]), .Z(n_43044));
	notech_inv i_60378(.A(n_3554), .Z(n_43045));
	notech_inv i_60379(.A(queue[129]), .Z(n_43046));
	notech_inv i_60380(.A(n_3560), .Z(n_43047));
	notech_inv i_60381(.A(queue[130]), .Z(n_43048));
	notech_inv i_60382(.A(n_3566), .Z(n_43049));
	notech_inv i_60383(.A(queue[131]), .Z(n_43050));
	notech_inv i_60384(.A(n_3572), .Z(n_43051));
	notech_inv i_60385(.A(queue[132]), .Z(n_43052));
	notech_inv i_60386(.A(n_3578), .Z(n_43053));
	notech_inv i_60387(.A(queue[133]), .Z(n_43054));
	notech_inv i_60388(.A(n_3584), .Z(n_43055));
	notech_inv i_60389(.A(queue[134]), .Z(n_43056));
	notech_inv i_60390(.A(n_3590), .Z(n_43057));
	notech_inv i_60391(.A(queue[135]), .Z(n_43058));
	notech_inv i_60392(.A(n_3596), .Z(n_43059));
	notech_inv i_60393(.A(queue[136]), .Z(n_43060));
	notech_inv i_60394(.A(n_3602), .Z(n_43061));
	notech_inv i_60395(.A(queue[137]), .Z(n_43062));
	notech_inv i_60396(.A(n_3608), .Z(n_43063));
	notech_inv i_60397(.A(queue[138]), .Z(n_43064));
	notech_inv i_60398(.A(n_3614), .Z(n_43065));
	notech_inv i_60399(.A(queue[139]), .Z(n_43066));
	notech_inv i_60400(.A(n_3620), .Z(n_43067));
	notech_inv i_60401(.A(queue[140]), .Z(n_43068));
	notech_inv i_60402(.A(n_3626), .Z(n_43069));
	notech_inv i_60403(.A(queue[141]), .Z(n_43070));
	notech_inv i_60404(.A(n_3632), .Z(n_43071));
	notech_inv i_60405(.A(queue[142]), .Z(n_43072));
	notech_inv i_60406(.A(n_3638), .Z(n_43073));
	notech_inv i_60407(.A(queue[143]), .Z(n_43074));
	notech_inv i_60408(.A(n_3644), .Z(n_43075));
	notech_inv i_60409(.A(queue[144]), .Z(n_43076));
	notech_inv i_60410(.A(n_3650), .Z(n_43077));
	notech_inv i_60411(.A(queue[145]), .Z(n_43078));
	notech_inv i_60412(.A(n_3656), .Z(n_43079));
	notech_inv i_60413(.A(queue[146]), .Z(n_43080));
	notech_inv i_60414(.A(n_3662), .Z(n_43081));
	notech_inv i_60415(.A(queue[147]), .Z(n_43082));
	notech_inv i_60416(.A(n_3668), .Z(n_43083));
	notech_inv i_60417(.A(queue[148]), .Z(n_43084));
	notech_inv i_60418(.A(queue[149]), .Z(n_43085));
	notech_inv i_60419(.A(n_3680), .Z(n_43086));
	notech_inv i_60420(.A(queue[150]), .Z(n_43087));
	notech_inv i_60421(.A(n_3686), .Z(n_43088));
	notech_inv i_60422(.A(queue[151]), .Z(n_43089));
	notech_inv i_60423(.A(n_3692), .Z(n_43090));
	notech_inv i_60424(.A(queue[152]), .Z(n_43091));
	notech_inv i_60425(.A(n_3698), .Z(n_43092));
	notech_inv i_60426(.A(queue[153]), .Z(n_43093));
	notech_inv i_60427(.A(n_3704), .Z(n_43094));
	notech_inv i_60428(.A(queue[154]), .Z(n_43095));
	notech_inv i_60429(.A(n_3710), .Z(n_43096));
	notech_inv i_60430(.A(queue[155]), .Z(n_43097));
	notech_inv i_60431(.A(n_3716), .Z(n_43098));
	notech_inv i_60432(.A(queue[156]), .Z(n_43099));
	notech_inv i_60433(.A(n_3722), .Z(n_43100));
	notech_inv i_60434(.A(queue[157]), .Z(n_43101));
	notech_inv i_60435(.A(n_3728), .Z(n_43102));
	notech_inv i_60436(.A(queue[158]), .Z(n_43103));
	notech_inv i_60437(.A(n_3734), .Z(n_43104));
	notech_inv i_60438(.A(queue[159]), .Z(n_43105));
	notech_inv i_60439(.A(n_3740), .Z(n_43106));
	notech_inv i_60440(.A(queue[160]), .Z(n_43107));
	notech_inv i_60441(.A(n_3746), .Z(n_43108));
	notech_inv i_60442(.A(queue[161]), .Z(n_43109));
	notech_inv i_60443(.A(n_3752), .Z(n_43110));
	notech_inv i_60444(.A(queue[162]), .Z(n_43111));
	notech_inv i_60445(.A(n_3758), .Z(n_43112));
	notech_inv i_60446(.A(queue[163]), .Z(n_43113));
	notech_inv i_60447(.A(n_3764), .Z(n_43114));
	notech_inv i_60448(.A(queue[164]), .Z(n_43115));
	notech_inv i_60449(.A(n_3770), .Z(n_43116));
	notech_inv i_60450(.A(queue[165]), .Z(n_43117));
	notech_inv i_60451(.A(n_3776), .Z(n_43118));
	notech_inv i_60452(.A(queue[166]), .Z(n_43119));
	notech_inv i_60453(.A(n_3782), .Z(n_43120));
	notech_inv i_60454(.A(queue[167]), .Z(n_43121));
	notech_inv i_60455(.A(n_3788), .Z(n_43122));
	notech_inv i_60456(.A(queue[168]), .Z(n_43123));
	notech_inv i_60457(.A(n_3794), .Z(n_43124));
	notech_inv i_60458(.A(queue[169]), .Z(n_43125));
	notech_inv i_60459(.A(n_3800), .Z(n_43126));
	notech_inv i_60460(.A(queue[170]), .Z(n_43127));
	notech_inv i_60461(.A(n_3806), .Z(n_43128));
	notech_inv i_60462(.A(queue[171]), .Z(n_43129));
	notech_inv i_60463(.A(n_3812), .Z(n_43130));
	notech_inv i_60464(.A(queue[172]), .Z(n_43131));
	notech_inv i_60465(.A(n_3818), .Z(n_43132));
	notech_inv i_60466(.A(queue[173]), .Z(n_43133));
	notech_inv i_60467(.A(n_3824), .Z(n_43134));
	notech_inv i_60468(.A(queue[174]), .Z(n_43135));
	notech_inv i_60469(.A(n_3830), .Z(n_43136));
	notech_inv i_60470(.A(queue[175]), .Z(n_43137));
	notech_inv i_60471(.A(n_3836), .Z(n_43138));
	notech_inv i_60472(.A(queue[176]), .Z(n_43139));
	notech_inv i_60473(.A(n_3842), .Z(n_43140));
	notech_inv i_60474(.A(queue[177]), .Z(n_43141));
	notech_inv i_60475(.A(n_3848), .Z(n_43142));
	notech_inv i_60476(.A(queue[178]), .Z(n_43143));
	notech_inv i_60477(.A(queue[179]), .Z(n_43144));
	notech_inv i_60478(.A(n_3860), .Z(n_43145));
	notech_inv i_60479(.A(queue[180]), .Z(n_43146));
	notech_inv i_60480(.A(n_3866), .Z(n_43147));
	notech_inv i_60481(.A(queue[181]), .Z(n_43148));
	notech_inv i_60482(.A(n_3872), .Z(n_43149));
	notech_inv i_60483(.A(queue[182]), .Z(n_43150));
	notech_inv i_60484(.A(n_3878), .Z(n_43151));
	notech_inv i_60485(.A(queue[183]), .Z(n_43152));
	notech_inv i_60486(.A(n_3884), .Z(n_43153));
	notech_inv i_60487(.A(queue[184]), .Z(n_43154));
	notech_inv i_60488(.A(n_3890), .Z(n_43155));
	notech_inv i_60489(.A(queue[185]), .Z(n_43156));
	notech_inv i_60490(.A(n_3896), .Z(n_43157));
	notech_inv i_60491(.A(queue[186]), .Z(n_43158));
	notech_inv i_60492(.A(n_3902), .Z(n_43159));
	notech_inv i_60493(.A(queue[187]), .Z(n_43160));
	notech_inv i_60494(.A(n_3908), .Z(n_43161));
	notech_inv i_60495(.A(queue[188]), .Z(n_43162));
	notech_inv i_60496(.A(n_3914), .Z(n_43163));
	notech_inv i_60497(.A(queue[189]), .Z(n_43164));
	notech_inv i_60498(.A(n_3920), .Z(n_43165));
	notech_inv i_60499(.A(queue[190]), .Z(n_43166));
	notech_inv i_60500(.A(n_3926), .Z(n_43167));
	notech_inv i_60501(.A(queue[191]), .Z(n_43168));
	notech_inv i_60502(.A(n_3932), .Z(n_43169));
	notech_inv i_60503(.A(queue[192]), .Z(n_43170));
	notech_inv i_60504(.A(n_3938), .Z(n_43171));
	notech_inv i_60505(.A(queue[193]), .Z(n_43172));
	notech_inv i_60506(.A(n_3944), .Z(n_43173));
	notech_inv i_60507(.A(queue[194]), .Z(n_43174));
	notech_inv i_60508(.A(n_3950), .Z(n_43175));
	notech_inv i_60509(.A(queue[195]), .Z(n_43176));
	notech_inv i_60510(.A(n_3956), .Z(n_43177));
	notech_inv i_60511(.A(queue[196]), .Z(n_43178));
	notech_inv i_60512(.A(n_3962), .Z(n_43179));
	notech_inv i_60513(.A(queue[197]), .Z(n_43180));
	notech_inv i_60514(.A(n_3968), .Z(n_43181));
	notech_inv i_60515(.A(queue[198]), .Z(n_43182));
	notech_inv i_60516(.A(n_3974), .Z(n_43183));
	notech_inv i_60517(.A(queue[199]), .Z(n_43184));
	notech_inv i_60518(.A(n_3980), .Z(n_43185));
	notech_inv i_60519(.A(queue[200]), .Z(n_43186));
	notech_inv i_60520(.A(n_3986), .Z(n_43187));
	notech_inv i_60521(.A(queue[201]), .Z(n_43188));
	notech_inv i_60522(.A(n_3992), .Z(n_43189));
	notech_inv i_60523(.A(queue[202]), .Z(n_43190));
	notech_inv i_60524(.A(n_3998), .Z(n_43191));
	notech_inv i_60525(.A(queue[203]), .Z(n_43192));
	notech_inv i_60526(.A(n_4004), .Z(n_43193));
	notech_inv i_60527(.A(queue[204]), .Z(n_43194));
	notech_inv i_60528(.A(n_4010), .Z(n_43195));
	notech_inv i_60529(.A(queue[205]), .Z(n_43196));
	notech_inv i_60530(.A(n_4016), .Z(n_43197));
	notech_inv i_60531(.A(queue[206]), .Z(n_43198));
	notech_inv i_60532(.A(n_4022), .Z(n_43199));
	notech_inv i_60533(.A(queue[207]), .Z(n_43200));
	notech_inv i_60534(.A(queue[208]), .Z(n_43201));
	notech_inv i_60535(.A(n_4034), .Z(n_43202));
	notech_inv i_60536(.A(queue[209]), .Z(n_43203));
	notech_inv i_60537(.A(n_4040), .Z(n_43204));
	notech_inv i_60538(.A(queue[210]), .Z(n_43205));
	notech_inv i_60539(.A(n_4046), .Z(n_43206));
	notech_inv i_60540(.A(queue[211]), .Z(n_43207));
	notech_inv i_60541(.A(n_4052), .Z(n_43208));
	notech_inv i_60542(.A(queue[212]), .Z(n_43209));
	notech_inv i_60543(.A(n_4058), .Z(n_43210));
	notech_inv i_60544(.A(queue[213]), .Z(n_43211));
	notech_inv i_60545(.A(n_4064), .Z(n_43212));
	notech_inv i_60546(.A(queue[214]), .Z(n_43213));
	notech_inv i_60547(.A(n_4070), .Z(n_43214));
	notech_inv i_60548(.A(queue[215]), .Z(n_43215));
	notech_inv i_60549(.A(n_4076), .Z(n_43216));
	notech_inv i_60550(.A(queue[216]), .Z(n_43217));
	notech_inv i_60551(.A(n_4082), .Z(n_43218));
	notech_inv i_60552(.A(queue[217]), .Z(n_43219));
	notech_inv i_60553(.A(n_4088), .Z(n_43220));
	notech_inv i_60554(.A(queue[218]), .Z(n_43221));
	notech_inv i_60555(.A(n_4094), .Z(n_43222));
	notech_inv i_60556(.A(queue[219]), .Z(n_43223));
	notech_inv i_60557(.A(n_4100), .Z(n_43224));
	notech_inv i_60558(.A(queue[220]), .Z(n_43225));
	notech_inv i_60559(.A(n_4106), .Z(n_43226));
	notech_inv i_60560(.A(queue[221]), .Z(n_43227));
	notech_inv i_60561(.A(n_4112), .Z(n_43228));
	notech_inv i_60562(.A(queue[222]), .Z(n_43229));
	notech_inv i_60563(.A(n_4118), .Z(n_43230));
	notech_inv i_60564(.A(queue[223]), .Z(n_43231));
	notech_inv i_60565(.A(n_4124), .Z(n_43232));
	notech_inv i_60566(.A(queue[224]), .Z(n_43233));
	notech_inv i_60567(.A(n_4130), .Z(n_43234));
	notech_inv i_60568(.A(queue[225]), .Z(n_43235));
	notech_inv i_60569(.A(n_4136), .Z(n_43236));
	notech_inv i_60570(.A(queue[226]), .Z(n_43237));
	notech_inv i_60571(.A(n_4142), .Z(n_43238));
	notech_inv i_60572(.A(queue[227]), .Z(n_43239));
	notech_inv i_60573(.A(n_4148), .Z(n_43240));
	notech_inv i_60574(.A(queue[228]), .Z(n_43241));
	notech_inv i_60575(.A(n_4154), .Z(n_43242));
	notech_inv i_60576(.A(queue[229]), .Z(n_43243));
	notech_inv i_60577(.A(n_4160), .Z(n_43244));
	notech_inv i_60578(.A(queue[230]), .Z(n_43245));
	notech_inv i_60579(.A(n_4166), .Z(n_43246));
	notech_inv i_60580(.A(queue[231]), .Z(n_43247));
	notech_inv i_60581(.A(n_4172), .Z(n_43248));
	notech_inv i_60582(.A(queue[232]), .Z(n_43249));
	notech_inv i_60583(.A(n_4178), .Z(n_43250));
	notech_inv i_60584(.A(queue[233]), .Z(n_43251));
	notech_inv i_60585(.A(n_4184), .Z(n_43252));
	notech_inv i_60586(.A(queue[234]), .Z(n_43253));
	notech_inv i_60587(.A(n_4190), .Z(n_43254));
	notech_inv i_60588(.A(queue[235]), .Z(n_43255));
	notech_inv i_60589(.A(n_4196), .Z(n_43256));
	notech_inv i_60590(.A(queue[236]), .Z(n_43257));
	notech_inv i_60591(.A(n_4202), .Z(n_43258));
	notech_inv i_60592(.A(queue[237]), .Z(n_43259));
	notech_inv i_60593(.A(n_4208), .Z(n_43260));
	notech_inv i_60594(.A(queue[238]), .Z(n_43261));
	notech_inv i_60595(.A(n_4214), .Z(n_43262));
	notech_inv i_60596(.A(queue[239]), .Z(n_43263));
	notech_inv i_60597(.A(n_4220), .Z(n_43264));
	notech_inv i_60598(.A(queue[240]), .Z(n_43265));
	notech_inv i_60599(.A(n_4226), .Z(n_43266));
	notech_inv i_60600(.A(queue[241]), .Z(n_43267));
	notech_inv i_60601(.A(n_4232), .Z(n_43268));
	notech_inv i_60602(.A(queue[242]), .Z(n_43269));
	notech_inv i_60603(.A(n_4238), .Z(n_43270));
	notech_inv i_60604(.A(queue[243]), .Z(n_43271));
	notech_inv i_60605(.A(n_4244), .Z(n_43272));
	notech_inv i_60606(.A(queue[244]), .Z(n_43273));
	notech_inv i_60607(.A(n_4250), .Z(n_43274));
	notech_inv i_60608(.A(queue[245]), .Z(n_43275));
	notech_inv i_60609(.A(n_4256), .Z(n_43276));
	notech_inv i_60610(.A(queue[246]), .Z(n_43277));
	notech_inv i_60611(.A(n_4262), .Z(n_43278));
	notech_inv i_60612(.A(queue[247]), .Z(n_43279));
	notech_inv i_60613(.A(n_4268), .Z(n_43280));
	notech_inv i_60614(.A(queue[248]), .Z(n_43281));
	notech_inv i_60615(.A(n_4274), .Z(n_43282));
	notech_inv i_60616(.A(queue[249]), .Z(n_43283));
	notech_inv i_60617(.A(n_4280), .Z(n_43284));
	notech_inv i_60618(.A(queue[250]), .Z(n_43285));
	notech_inv i_60619(.A(n_4286), .Z(n_43286));
	notech_inv i_60620(.A(queue[251]), .Z(n_43287));
	notech_inv i_60621(.A(n_4292), .Z(n_43288));
	notech_inv i_60622(.A(queue[252]), .Z(n_43289));
	notech_inv i_60623(.A(n_4298), .Z(n_43290));
	notech_inv i_60624(.A(queue[253]), .Z(n_43291));
	notech_inv i_60625(.A(n_4304), .Z(n_43292));
	notech_inv i_60626(.A(queue[254]), .Z(n_43293));
	notech_inv i_60627(.A(n_4310), .Z(n_43294));
	notech_inv i_60628(.A(queue[255]), .Z(n_43295));
	notech_inv i_60629(.A(addrshft[0]), .Z(n_43296));
	notech_inv i_60630(.A(addrshft[1]), .Z(n_43297));
	notech_inv i_60631(.A(addrshft[2]), .Z(n_43298));
	notech_inv i_60632(.A(addrshft[3]), .Z(n_43299));
	notech_inv i_60633(.A(addrshft[4]), .Z(n_43300));
	notech_inv i_60634(.A(addrshft[5]), .Z(n_43301));
	notech_inv i_60635(.A(squeue_0100306), .Z(squeue[0]));
	notech_inv i_60636(.A(squeue_1100305), .Z(squeue[1]));
	notech_inv i_60637(.A(squeue_2100304), .Z(squeue[2]));
	notech_inv i_60638(.A(squeue_3100303), .Z(squeue[3]));
	notech_inv i_60639(.A(squeue_4100302), .Z(squeue[4]));
	notech_inv i_60640(.A(squeue_5100301), .Z(squeue[5]));
	notech_inv i_60641(.A(squeue_6100300), .Z(squeue[6]));
	notech_inv i_60642(.A(squeue_7100299), .Z(squeue[7]));
	notech_inv i_60643(.A(squeue_9100298), .Z(squeue[9]));
	notech_inv i_60644(.A(squeue_10100297), .Z(squeue[10]));
	notech_inv i_60645(.A(squeue_11100296), .Z(squeue[11]));
	notech_inv i_60646(.A(squeue_12100295), .Z(squeue[12]));
	notech_inv i_60647(.A(squeue_13100294), .Z(squeue[13]));
	notech_inv i_60648(.A(squeue_15100293), .Z(squeue[15]));
	notech_inv i_60649(.A(squeue_16100292), .Z(squeue[16]));
	notech_inv i_60650(.A(squeue_17100291), .Z(squeue[17]));
	notech_inv i_60651(.A(squeue_18100290), .Z(squeue[18]));
	notech_inv i_60652(.A(squeue_19100289), .Z(squeue[19]));
	notech_inv i_60653(.A(squeue_20100288), .Z(squeue[20]));
	notech_inv i_60654(.A(squeue_21100287), .Z(squeue[21]));
	notech_inv i_60655(.A(squeue_22100286), .Z(squeue[22]));
	notech_inv i_60656(.A(squeue_23100285), .Z(squeue[23]));
	notech_inv i_60657(.A(squeue_24100284), .Z(squeue[24]));
	notech_inv i_60658(.A(squeue_25100283), .Z(squeue[25]));
	notech_inv i_60659(.A(squeue_26100282), .Z(squeue[26]));
	notech_inv i_60660(.A(squeue_27100281), .Z(squeue[27]));
	notech_inv i_60661(.A(squeue_28100280), .Z(squeue[28]));
	notech_inv i_60662(.A(squeue_30100279), .Z(squeue[30]));
	notech_inv i_60663(.A(squeue_31100278), .Z(squeue[31]));
	notech_inv i_60664(.A(squeue_32100277), .Z(squeue[32]));
	notech_inv i_60665(.A(squeue_33100276), .Z(squeue[33]));
	notech_inv i_60666(.A(squeue_34100275), .Z(squeue[34]));
	notech_inv i_60667(.A(squeue_35100274), .Z(squeue[35]));
	notech_inv i_60668(.A(squeue_36100273), .Z(squeue[36]));
	notech_inv i_60669(.A(squeue_38100272), .Z(squeue[38]));
	notech_inv i_60670(.A(squeue_39100271), .Z(squeue[39]));
	notech_inv i_60671(.A(squeue_40100270), .Z(squeue[40]));
	notech_inv i_60672(.A(squeue_41100269), .Z(squeue[41]));
	notech_inv i_60673(.A(squeue_42100268), .Z(squeue[42]));
	notech_inv i_60674(.A(squeue_43100267), .Z(squeue[43]));
	notech_inv i_60675(.A(squeue_44100266), .Z(squeue[44]));
	notech_inv i_60676(.A(squeue_45100265), .Z(squeue[45]));
	notech_inv i_60677(.A(squeue_46100264), .Z(squeue[46]));
	notech_inv i_60678(.A(squeue_47100263), .Z(squeue[47]));
	notech_inv i_60679(.A(squeue_48100262), .Z(squeue[48]));
	notech_inv i_60680(.A(squeue_49100261), .Z(squeue[49]));
	notech_inv i_60681(.A(squeue_50100260), .Z(squeue[50]));
	notech_inv i_60682(.A(squeue_51100259), .Z(squeue[51]));
	notech_inv i_60683(.A(squeue_52100258), .Z(squeue[52]));
	notech_inv i_60684(.A(squeue_65100257), .Z(squeue[65]));
	notech_inv i_60685(.A(purge_cnt[10]), .Z(n_43352));
	notech_inv i_60686(.A(idata[0]), .Z(n_43353));
	notech_inv i_60687(.A(idata[1]), .Z(n_43354));
	notech_inv i_60688(.A(idata[2]), .Z(n_43355));
	notech_inv i_60689(.A(idata[3]), .Z(n_43356));
	notech_inv i_60690(.A(idata[4]), .Z(n_43357));
	notech_inv i_60691(.A(idata[5]), .Z(n_43358));
	notech_inv i_60692(.A(idata[6]), .Z(n_43359));
	notech_inv i_60693(.A(idata[7]), .Z(n_43360));
	notech_inv i_60694(.A(idata[8]), .Z(n_43361));
	notech_inv i_60695(.A(idata[9]), .Z(n_43362));
	notech_inv i_60696(.A(idata[10]), .Z(n_43363));
	notech_inv i_60697(.A(idata[11]), .Z(n_43364));
	notech_inv i_60698(.A(idata[12]), .Z(n_43365));
	notech_inv i_60699(.A(idata[13]), .Z(n_43366));
	notech_inv i_60700(.A(idata[14]), .Z(n_43367));
	notech_inv i_60701(.A(idata[15]), .Z(n_43368));
	notech_inv i_60702(.A(idata[16]), .Z(n_43369));
	notech_inv i_60703(.A(idata[17]), .Z(n_43370));
	notech_inv i_60704(.A(idata[18]), .Z(n_43371));
	notech_inv i_60705(.A(idata[19]), .Z(n_43372));
	notech_inv i_60706(.A(idata[20]), .Z(n_43373));
	notech_inv i_60707(.A(idata[21]), .Z(n_43374));
	notech_inv i_60708(.A(idata[22]), .Z(n_43375));
	notech_inv i_60709(.A(idata[23]), .Z(n_43376));
	notech_inv i_60710(.A(idata[24]), .Z(n_43377));
	notech_inv i_60711(.A(idata[25]), .Z(n_43378));
	notech_inv i_60712(.A(idata[26]), .Z(n_43379));
	notech_inv i_60713(.A(idata[27]), .Z(n_43380));
	notech_inv i_60714(.A(idata[28]), .Z(n_43381));
	notech_inv i_60715(.A(idata[29]), .Z(n_43382));
	notech_inv i_60716(.A(idata[30]), .Z(n_43383));
	notech_inv i_60717(.A(idata[31]), .Z(n_43384));
	notech_inv i_60718(.A(idata[32]), .Z(n_43385));
	notech_inv i_60719(.A(idata[33]), .Z(n_43386));
	notech_inv i_60720(.A(idata[34]), .Z(n_43387));
	notech_inv i_60721(.A(idata[35]), .Z(n_43388));
	notech_inv i_60722(.A(idata[36]), .Z(n_43389));
	notech_inv i_60723(.A(idata[37]), .Z(n_43390));
	notech_inv i_60724(.A(idata[38]), .Z(n_43391));
	notech_inv i_60725(.A(idata[39]), .Z(n_43392));
	notech_inv i_60726(.A(idata[40]), .Z(n_43393));
	notech_inv i_60727(.A(idata[41]), .Z(n_43394));
	notech_inv i_60728(.A(idata[42]), .Z(n_43395));
	notech_inv i_60729(.A(idata[43]), .Z(n_43396));
	notech_inv i_60730(.A(idata[44]), .Z(n_43397));
	notech_inv i_60731(.A(idata[45]), .Z(n_43398));
	notech_inv i_60732(.A(idata[46]), .Z(n_43399));
	notech_inv i_60733(.A(idata[47]), .Z(n_43400));
	notech_inv i_60734(.A(idata[48]), .Z(n_43401));
	notech_inv i_60735(.A(idata[49]), .Z(n_43402));
	notech_inv i_60736(.A(idata[50]), .Z(n_43403));
	notech_inv i_60737(.A(idata[51]), .Z(n_43404));
	notech_inv i_60738(.A(idata[52]), .Z(n_43405));
	notech_inv i_60739(.A(idata[53]), .Z(n_43406));
	notech_inv i_60740(.A(idata[54]), .Z(n_43407));
	notech_inv i_60741(.A(idata[55]), .Z(n_43408));
	notech_inv i_60742(.A(idata[56]), .Z(n_43409));
	notech_inv i_60743(.A(idata[57]), .Z(n_43410));
	notech_inv i_60744(.A(idata[58]), .Z(n_43411));
	notech_inv i_60745(.A(idata[59]), .Z(n_43412));
	notech_inv i_60746(.A(idata[60]), .Z(n_43413));
	notech_inv i_60747(.A(idata[61]), .Z(n_43414));
	notech_inv i_60748(.A(idata[62]), .Z(n_43415));
	notech_inv i_60749(.A(idata[63]), .Z(n_43416));
	notech_inv i_60750(.A(idata[64]), .Z(n_43417));
	notech_inv i_60751(.A(idata[65]), .Z(n_43418));
	notech_inv i_60752(.A(idata[66]), .Z(n_43419));
	notech_inv i_60753(.A(idata[67]), .Z(n_43420));
	notech_inv i_60754(.A(idata[68]), .Z(n_43421));
	notech_inv i_60755(.A(idata[69]), .Z(n_43422));
	notech_inv i_60756(.A(idata[70]), .Z(n_43423));
	notech_inv i_60757(.A(idata[71]), .Z(n_43424));
	notech_inv i_60758(.A(idata[72]), .Z(n_43425));
	notech_inv i_60759(.A(idata[73]), .Z(n_43426));
	notech_inv i_60760(.A(idata[74]), .Z(n_43427));
	notech_inv i_60761(.A(idata[75]), .Z(n_43428));
	notech_inv i_60762(.A(idata[76]), .Z(n_43429));
	notech_inv i_60763(.A(idata[77]), .Z(n_43430));
	notech_inv i_60764(.A(idata[78]), .Z(n_43431));
	notech_inv i_60765(.A(idata[79]), .Z(n_43432));
	notech_inv i_60766(.A(idata[80]), .Z(n_43433));
	notech_inv i_60767(.A(idata[81]), .Z(n_43434));
	notech_inv i_60768(.A(idata[82]), .Z(n_43435));
	notech_inv i_60769(.A(idata[83]), .Z(n_43436));
	notech_inv i_60770(.A(idata[84]), .Z(n_43437));
	notech_inv i_60771(.A(idata[85]), .Z(n_43438));
	notech_inv i_60772(.A(idata[86]), .Z(n_43439));
	notech_inv i_60773(.A(idata[87]), .Z(n_43440));
	notech_inv i_60774(.A(idata[88]), .Z(n_43441));
	notech_inv i_60775(.A(idata[89]), .Z(n_43442));
	notech_inv i_60776(.A(idata[90]), .Z(n_43443));
	notech_inv i_60777(.A(idata[91]), .Z(n_43444));
	notech_inv i_60778(.A(idata[92]), .Z(n_43445));
	notech_inv i_60779(.A(idata[93]), .Z(n_43446));
	notech_inv i_60780(.A(idata[94]), .Z(n_43447));
	notech_inv i_60781(.A(idata[95]), .Z(n_43448));
	notech_inv i_60782(.A(idata[96]), .Z(n_43449));
	notech_inv i_60783(.A(idata[97]), .Z(n_43450));
	notech_inv i_60784(.A(idata[98]), .Z(n_43451));
	notech_inv i_60785(.A(idata[99]), .Z(n_43452));
	notech_inv i_60786(.A(idata[100]), .Z(n_43453));
	notech_inv i_60787(.A(idata[101]), .Z(n_43454));
	notech_inv i_60788(.A(idata[102]), .Z(n_43455));
	notech_inv i_60789(.A(idata[103]), .Z(n_43456));
	notech_inv i_60790(.A(idata[104]), .Z(n_43457));
	notech_inv i_60791(.A(idata[105]), .Z(n_43458));
	notech_inv i_60792(.A(idata[106]), .Z(n_43459));
	notech_inv i_60793(.A(idata[107]), .Z(n_43460));
	notech_inv i_60794(.A(idata[108]), .Z(n_43461));
	notech_inv i_60795(.A(idata[109]), .Z(n_43462));
	notech_inv i_60796(.A(idata[110]), .Z(n_43463));
	notech_inv i_60797(.A(idata[111]), .Z(n_43464));
	notech_inv i_60798(.A(idata[112]), .Z(n_43465));
	notech_inv i_60799(.A(idata[113]), .Z(n_43466));
	notech_inv i_60800(.A(idata[114]), .Z(n_43467));
	notech_inv i_60801(.A(idata[115]), .Z(n_43468));
	notech_inv i_60802(.A(idata[116]), .Z(n_43469));
	notech_inv i_60803(.A(idata[117]), .Z(n_43470));
	notech_inv i_60804(.A(idata[118]), .Z(n_43471));
	notech_inv i_60805(.A(idata[119]), .Z(n_43472));
	notech_inv i_60806(.A(idata[120]), .Z(n_43473));
	notech_inv i_60807(.A(idata[121]), .Z(n_43474));
	notech_inv i_60808(.A(idata[122]), .Z(n_43475));
	notech_inv i_60809(.A(idata[123]), .Z(n_43476));
	notech_inv i_60810(.A(idata[124]), .Z(n_43477));
	notech_inv i_60811(.A(idata[125]), .Z(n_43478));
	notech_inv i_60812(.A(idata[126]), .Z(n_43479));
	notech_inv i_60813(.A(idata[127]), .Z(n_43480));
	notech_inv i_60814(.A(nbus_81[4]), .Z(n_43481));
	notech_inv i_60815(.A(nbus_81[5]), .Z(n_43482));
	notech_inv i_60816(.A(valid_len_0100253), .Z(valid_len[0]));
	notech_inv i_60817(.A(valid_len_1100256), .Z(valid_len[1]));
	notech_inv i_60818(.A(valid_len_2100255), .Z(valid_len[2]));
	notech_inv i_60819(.A(valid_len_3100252), .Z(valid_len[3]));
	notech_inv i_60820(.A(valid_len_5100254), .Z(valid_len[5]));
	notech_inv i_60821(.A(busy_ram), .Z(n_43488));
	notech_inv i_60822(.A(n_60750), .Z(n_43489));
	notech_inv i_60823(.A(\queue_0[127] ), .Z(n_43490));
	notech_inv i_60824(.A(\queue_0[126] ), .Z(n_43491));
	notech_inv i_60825(.A(\queue_0[125] ), .Z(n_43492));
	notech_inv i_60826(.A(\queue_0[124] ), .Z(n_43493));
	notech_inv i_60827(.A(\queue_0[123] ), .Z(n_43494));
	notech_inv i_60828(.A(\queue_0[122] ), .Z(n_43495));
	notech_inv i_60829(.A(\queue_0[121] ), .Z(n_43496));
	notech_inv i_60830(.A(\queue_0[120] ), .Z(n_43497));
	notech_inv i_60831(.A(\queue_0[119] ), .Z(n_43498));
	notech_inv i_60832(.A(\queue_0[118] ), .Z(n_43499));
	notech_inv i_60833(.A(\queue_0[117] ), .Z(n_43500));
	notech_inv i_60834(.A(\queue_0[116] ), .Z(n_43501));
	notech_inv i_60835(.A(\queue_0[115] ), .Z(n_43502));
	notech_inv i_60836(.A(\queue_0[114] ), .Z(n_43503));
	notech_inv i_60837(.A(\queue_0[113] ), .Z(n_43504));
	notech_inv i_60838(.A(\queue_0[112] ), .Z(n_43505));
	notech_inv i_60839(.A(\queue_0[111] ), .Z(n_43506));
	notech_inv i_60840(.A(\queue_0[110] ), .Z(n_43507));
	notech_inv i_60841(.A(\queue_0[109] ), .Z(n_43508));
	notech_inv i_60842(.A(\queue_0[108] ), .Z(n_43509));
	notech_inv i_60843(.A(\queue_0[107] ), .Z(n_43510));
	notech_inv i_60844(.A(\queue_0[106] ), .Z(n_43511));
	notech_inv i_60845(.A(\queue_0[105] ), .Z(n_43512));
	notech_inv i_60846(.A(\queue_0[104] ), .Z(n_43513));
	notech_inv i_60847(.A(\queue_0[103] ), .Z(n_43514));
	notech_inv i_60848(.A(\queue_0[102] ), .Z(n_43515));
	notech_inv i_60849(.A(\queue_0[101] ), .Z(n_43516));
	notech_inv i_60850(.A(\queue_0[100] ), .Z(n_43517));
	notech_inv i_60851(.A(\queue_0[99] ), .Z(n_43518));
	notech_inv i_60852(.A(\queue_0[98] ), .Z(n_43519));
	notech_inv i_60853(.A(\queue_0[97] ), .Z(n_43520));
	notech_inv i_60854(.A(\queue_0[96] ), .Z(n_43521));
	notech_inv i_60855(.A(\queue_0[95] ), .Z(n_43522));
	notech_inv i_60856(.A(\queue_0[94] ), .Z(n_43523));
	notech_inv i_60857(.A(\queue_0[93] ), .Z(n_43524));
	notech_inv i_60858(.A(\queue_0[92] ), .Z(n_43525));
	notech_inv i_60859(.A(\queue_0[91] ), .Z(n_43526));
	notech_inv i_60860(.A(\queue_0[90] ), .Z(n_43527));
	notech_inv i_60861(.A(\queue_0[89] ), .Z(n_43528));
	notech_inv i_60862(.A(\queue_0[88] ), .Z(n_43529));
	notech_inv i_60863(.A(\queue_0[87] ), .Z(n_43530));
	notech_inv i_60864(.A(\queue_0[86] ), .Z(n_43531));
	notech_inv i_60865(.A(\queue_0[85] ), .Z(n_43532));
	notech_inv i_60866(.A(\queue_0[84] ), .Z(n_43533));
	notech_inv i_60867(.A(\queue_0[83] ), .Z(n_43534));
	notech_inv i_60868(.A(\queue_0[82] ), .Z(n_43535));
	notech_inv i_60869(.A(\queue_0[81] ), .Z(n_43536));
	notech_inv i_60870(.A(\queue_0[79] ), .Z(n_43537));
	notech_inv i_60871(.A(\queue_0[78] ), .Z(n_43538));
	notech_inv i_60872(.A(\queue_0[77] ), .Z(n_43539));
	notech_inv i_60873(.A(\queue_0[76] ), .Z(n_43540));
	notech_inv i_60874(.A(\queue_0[75] ), .Z(n_43541));
	notech_inv i_60875(.A(\queue_0[74] ), .Z(n_43542));
	notech_inv i_60876(.A(\queue_0[73] ), .Z(n_43543));
	notech_inv i_60877(.A(\queue_0[72] ), .Z(n_43544));
	notech_inv i_60878(.A(\queue_0[71] ), .Z(n_43545));
	notech_inv i_60879(.A(\queue_0[70] ), .Z(n_43546));
	notech_inv i_60880(.A(\queue_0[69] ), .Z(n_43547));
	notech_inv i_60881(.A(\queue_0[68] ), .Z(n_43548));
	notech_inv i_60882(.A(\queue_0[67] ), .Z(n_43549));
	notech_inv i_60883(.A(\queue_0[66] ), .Z(n_43550));
	notech_inv i_60884(.A(\queue_0[65] ), .Z(n_43551));
	notech_inv i_60885(.A(\queue_0[64] ), .Z(n_43552));
	notech_inv i_60886(.A(\queue_0[63] ), .Z(n_43553));
	notech_inv i_60887(.A(\queue_0[62] ), .Z(n_43554));
	notech_inv i_60888(.A(\queue_0[61] ), .Z(n_43555));
	notech_inv i_60889(.A(\queue_0[59] ), .Z(n_43556));
	notech_inv i_60890(.A(\queue_0[58] ), .Z(n_43557));
	notech_inv i_60891(.A(\queue_0[56] ), .Z(n_43558));
	notech_inv i_60892(.A(\queue_0[50] ), .Z(n_43559));
	notech_inv i_60893(.A(\queue_0[49] ), .Z(n_43560));
	notech_inv i_60894(.A(\queue_0[48] ), .Z(n_43561));
	notech_inv i_60895(.A(\queue_0[47] ), .Z(n_43562));
	notech_inv i_60896(.A(\queue_0[46] ), .Z(n_43563));
	notech_inv i_60897(.A(\queue_0[45] ), .Z(n_43564));
	notech_inv i_60898(.A(\queue_0[44] ), .Z(n_43565));
	notech_inv i_60899(.A(\queue_0[43] ), .Z(n_43566));
	notech_inv i_60900(.A(\queue_0[42] ), .Z(n_43567));
	notech_inv i_60901(.A(\queue_0[41] ), .Z(n_43568));
	notech_inv i_60902(.A(\queue_0[40] ), .Z(n_43569));
	notech_inv i_60903(.A(\queue_0[39] ), .Z(n_43570));
	notech_inv i_60904(.A(\queue_0[38] ), .Z(n_43571));
	notech_inv i_60905(.A(\queue_0[37] ), .Z(n_43572));
	notech_inv i_60906(.A(\queue_0[36] ), .Z(n_43573));
	notech_inv i_60907(.A(\queue_0[35] ), .Z(n_43574));
	notech_inv i_60908(.A(\queue_0[34] ), .Z(n_43575));
	notech_inv i_60909(.A(\queue_0[33] ), .Z(n_43576));
	notech_inv i_60910(.A(\queue_0[32] ), .Z(n_43577));
	notech_inv i_60911(.A(\queue_0[31] ), .Z(n_43578));
	notech_inv i_60912(.A(\queue_0[30] ), .Z(n_43579));
	notech_inv i_60913(.A(\queue_0[29] ), .Z(n_43580));
	notech_inv i_60914(.A(\queue_0[28] ), .Z(n_43581));
	notech_inv i_60915(.A(\queue_0[27] ), .Z(n_43582));
	notech_inv i_60916(.A(\queue_0[26] ), .Z(n_43583));
	notech_inv i_60917(.A(\queue_0[25] ), .Z(n_43584));
	notech_inv i_60918(.A(\queue_0[24] ), .Z(n_43585));
	notech_inv i_60919(.A(\queue_0[23] ), .Z(n_43586));
	notech_inv i_60920(.A(\queue_0[22] ), .Z(n_43587));
	notech_inv i_60921(.A(\queue_0[20] ), .Z(n_43588));
	notech_inv i_60922(.A(\queue_0[19] ), .Z(n_43589));
	notech_inv i_60923(.A(\queue_0[18] ), .Z(n_43590));
	notech_inv i_60924(.A(\queue_0[17] ), .Z(n_43591));
	notech_inv i_60925(.A(\queue_0[16] ), .Z(n_43592));
	notech_inv i_60926(.A(\queue_0[15] ), .Z(n_43593));
	notech_inv i_60927(.A(\queue_0[14] ), .Z(n_43594));
	notech_inv i_60928(.A(\queue_0[13] ), .Z(n_43595));
	notech_inv i_60929(.A(\queue_0[12] ), .Z(n_43596));
	notech_inv i_60930(.A(\queue_0[11] ), .Z(n_43597));
	notech_inv i_60931(.A(\queue_0[10] ), .Z(n_43598));
	notech_inv i_60932(.A(\queue_0[9] ), .Z(n_43599));
	notech_inv i_60933(.A(\queue_0[8] ), .Z(n_43600));
	notech_inv i_60934(.A(\queue_0[7] ), .Z(n_43601));
	notech_inv i_60935(.A(\queue_0[6] ), .Z(n_43602));
	notech_inv i_60936(.A(\queue_0[5] ), .Z(n_43603));
	notech_inv i_60937(.A(\queue_0[4] ), .Z(n_43604));
	notech_inv i_60938(.A(\queue_0[3] ), .Z(n_43605));
	notech_inv i_60939(.A(\queue_0[2] ), .Z(n_43606));
	notech_inv i_60940(.A(\queue_0[1] ), .Z(n_43607));
	notech_inv i_60941(.A(\queue_0[0] ), .Z(n_43608));
	notech_inv i_60942(.A(\queue_0[80] ), .Z(n_43609));
	notech_inv i_60943(.A(\queue_0[51] ), .Z(n_43610));
	notech_inv i_60944(.A(\queue_0[21] ), .Z(n_43611));
	notech_inv i_60945(.A(\queue_0[53] ), .Z(n_43612));
	notech_inv i_60946(.A(\queue_0[52] ), .Z(n_43613));
	notech_inv i_60947(.A(\queue_0[54] ), .Z(n_43614));
	notech_inv i_60948(.A(\queue_0[55] ), .Z(n_43615));
	notech_inv i_60949(.A(\queue_0[57] ), .Z(n_43616));
	notech_inv i_60950(.A(\queue_0[60] ), .Z(n_43617));
	AWDP_INC_1315491 i_656(.O0({n_2360, n_2358, n_2356, n_2354, n_2352, n_2350
		, n_2348, n_2346, n_2344, n_2342, n_2340}), .purge_cnt(purge_cnt
		));
	AWDP_EQ_3416052 i_641(.O0({n_4676}), .tagA(tagA), .addr({iaddr[31], iaddr
		[30], iaddr[29], iaddr[28], iaddr[27], iaddr[26], iaddr[25], iaddr
		[24], iaddr[23], iaddr[22], iaddr[21], iaddr[20], iaddr[19], iaddr
		[18], iaddr[17], iaddr[16], iaddr[15], iaddr[14]}));
	AWDP_EQ_2715865 i_636(.O0({n_2396}), .addr(iaddr), .addrf(addrf));
	AWDP_ADD_33 i_626(.O0(nbus_81), .addrshft(addrshft), .useq_ptr(useq_ptr)
		);
	AWDP_ADD_10 i_612(.O0(addr_0), .addr(iaddr));
	datacache c1(.clk(clk), .A(cacheA), .D({AMBIT_GND, cacheD[148], 
		AMBIT_GND, AMBIT_GND, cacheD[145], cacheD[144], cacheD[143], cacheD
		[142], cacheD[141], cacheD[140], cacheD[139], cacheD[138], cacheD
		[137], cacheD[136], cacheD[135], cacheD[134], cacheD[133], cacheD
		[132], cacheD[131], cacheD[130], cacheD[129], cacheD[128], cacheD
		[127], cacheD[126], cacheD[125], cacheD[124], cacheD[123], cacheD
		[122], cacheD[121], cacheD[120], cacheD[119], cacheD[118], cacheD
		[117], cacheD[116], cacheD[115], cacheD[114], cacheD[113], cacheD
		[112], cacheD[111], cacheD[110], cacheD[109], cacheD[108], cacheD
		[107], cacheD[106], cacheD[105], cacheD[104], cacheD[103], cacheD
		[102], cacheD[101], cacheD[100], cacheD[99], cacheD[98], cacheD[
		97], cacheD[96], cacheD[95], cacheD[94], cacheD[93], cacheD[92],
		 cacheD[91], cacheD[90], cacheD[89], cacheD[88], cacheD[87], cacheD
		[86], cacheD[85], cacheD[84], cacheD[83], cacheD[82], cacheD[81]
		, cacheD[80], cacheD[79], cacheD[78], cacheD[77], cacheD[76], cacheD
		[75], cacheD[74], cacheD[73], cacheD[72], cacheD[71], cacheD[70]
		, cacheD[69], cacheD[68], cacheD[67], cacheD[66], cacheD[65], cacheD
		[64], cacheD[63], cacheD[62], cacheD[61], cacheD[60], cacheD[59]
		, cacheD[58], cacheD[57], cacheD[56], cacheD[55], cacheD[54], cacheD
		[53], cacheD[52], cacheD[51], cacheD[50], cacheD[49], cacheD[48]
		, cacheD[47], cacheD[46], cacheD[45], cacheD[44], cacheD[43], cacheD
		[42], cacheD[41], cacheD[40], cacheD[39], cacheD[38], cacheD[37]
		, cacheD[36], cacheD[35], cacheD[34], cacheD[33], cacheD[32], cacheD
		[31], cacheD[30], cacheD[29], cacheD[28], cacheD[27], cacheD[26]
		, cacheD[25], cacheD[24], cacheD[23], cacheD[22], cacheD[21], cacheD
		[20], cacheD[19], cacheD[18], cacheD[17], cacheD[16], cacheD[15]
		, cacheD[14], cacheD[13], cacheD[12], cacheD[11], cacheD[10], cacheD
		[9], cacheD[8], cacheD[7], cacheD[6], cacheD[5], cacheD[4], cacheD
		[3], cacheD[2], cacheD[1], cacheD[0]}), .Q({tagV[3], tagV[2], tagV
		[1], tagV[0], tagA[17], tagA[16], tagA[15], tagA[14], tagA[13], tagA
		[12], tagA[11], tagA[10], tagA[9], tagA[8], tagA[7], tagA[6], tagA
		[5], tagA[4], tagA[3], tagA[2], tagA[1], tagA[0], \queue_0[127] 
		, \queue_0[126] , \queue_0[125] , \queue_0[124] , \queue_0[123] 
		, \queue_0[122] , \queue_0[121] , \queue_0[120] , \queue_0[119] 
		, \queue_0[118] , \queue_0[117] , \queue_0[116] , \queue_0[115] 
		, \queue_0[114] , \queue_0[113] , \queue_0[112] , \queue_0[111] 
		, \queue_0[110] , \queue_0[109] , \queue_0[108] , \queue_0[107] 
		, \queue_0[106] , \queue_0[105] , \queue_0[104] , \queue_0[103] 
		, \queue_0[102] , \queue_0[101] , \queue_0[100] , \queue_0[99] ,
		 \queue_0[98] , \queue_0[97] , \queue_0[96] , \queue_0[95] , \queue_0[94] 
		, \queue_0[93] , \queue_0[92] , \queue_0[91] , \queue_0[90] , \queue_0[89] 
		, \queue_0[88] , \queue_0[87] , \queue_0[86] , \queue_0[85] , \queue_0[84] 
		, \queue_0[83] , \queue_0[82] , \queue_0[81] , \queue_0[80] , \queue_0[79] 
		, \queue_0[78] , \queue_0[77] , \queue_0[76] , \queue_0[75] , \queue_0[74] 
		, \queue_0[73] , \queue_0[72] , \queue_0[71] , \queue_0[70] , \queue_0[69] 
		, \queue_0[68] , \queue_0[67] , \queue_0[66] , \queue_0[65] , \queue_0[64] 
		, \queue_0[63] , \queue_0[62] , \queue_0[61] , \queue_0[60] , \queue_0[59] 
		, \queue_0[58] , \queue_0[57] , \queue_0[56] , \queue_0[55] , \queue_0[54] 
		, \queue_0[53] , \queue_0[52] , \queue_0[51] , \queue_0[50] , \queue_0[49] 
		, \queue_0[48] , \queue_0[47] , \queue_0[46] , \queue_0[45] , \queue_0[44] 
		, \queue_0[43] , \queue_0[42] , \queue_0[41] , \queue_0[40] , \queue_0[39] 
		, \queue_0[38] , \queue_0[37] , \queue_0[36] , \queue_0[35] , \queue_0[34] 
		, \queue_0[33] , \queue_0[32] , \queue_0[31] , \queue_0[30] , \queue_0[29] 
		, \queue_0[28] , \queue_0[27] , \queue_0[26] , \queue_0[25] , \queue_0[24] 
		, \queue_0[23] , \queue_0[22] , \queue_0[21] , \queue_0[20] , \queue_0[19] 
		, \queue_0[18] , \queue_0[17] , \queue_0[16] , \queue_0[15] , \queue_0[14] 
		, \queue_0[13] , \queue_0[12] , \queue_0[11] , \queue_0[10] , \queue_0[9] 
		, \queue_0[8] , \queue_0[7] , \queue_0[6] , \queue_0[5] , \queue_0[4] 
		, \queue_0[3] , \queue_0[2] , \queue_0[1] , \queue_0[0] }), .WEN
		(codeWEN), .M({AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, 
		AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD
		, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, 
		AMBIT_VDD}));
endmodule
module core(clk, rstn, ivect, int_main, iack, code_addr, code_data, code_req, code_ack
		, code_wreq, code_wack, code_wdata, readio_data, io_add, writeio_data
		, writeio_req, readio_req, writeio_ack, readio_ack, write_req, write_ack
		, write_data, write_sz, read_sz, write_msk, read_req, read_ack, read_data
		, Daddr, busy_ram, ipg_fault, outstanding);

	input clk;
	input rstn;
	input [7:0] ivect;
	input int_main;
	output iack;
	output [31:0] code_addr;
	input [127:0] code_data;
	output code_req;
	input code_ack;
	output code_wreq;
	input code_wack;
	output [31:0] code_wdata;
	input [31:0] readio_data;
	output [31:0] io_add;
	output [31:0] writeio_data;
	output writeio_req;
	output readio_req;
	input writeio_ack;
	input readio_ack;
	output write_req;
	input write_ack;
	output [31:0] write_data;
	output [1:0] write_sz;
	output [1:0] read_sz;
	output [3:0] write_msk;
	output read_req;
	input read_ack;
	input [31:0] read_data;
	output [31:0] Daddr;
	input busy_ram;
	output ipg_fault;
	output outstanding;

	wire [31:0] write_data_realign;
	wire [31:0] read_data_realign;
	wire [31:0] Daddr_realign;
	wire [5:0] valid_len;
	wire [1:0] int_write_sz;
	wire [31:0] iwrite_data;
	wire [31:0] int_code_addr;
	wire [31:0] icr2;
	wire [31:0] cr2;
	wire [31:0] pc_out;
	wire [31:0] int_Daddr;
	wire [3:0] useq_ptr;
	wire [127:0] queue;
	wire [1:0] nbus_14524;



	realign i_realign(.clk(clk), .rstn(rstn), .write_msk_out(write_msk), .addr_in
		(Daddr_realign), .addr_out({Daddr[31], Daddr[30], Daddr[29], Daddr
		[28], Daddr[27], Daddr[26], Daddr[25], Daddr[24], Daddr[23], Daddr
		[22], Daddr[21], Daddr[20], Daddr[19], Daddr[18], Daddr[17], Daddr
		[16], Daddr[15], Daddr[14], Daddr[13], Daddr[12], Daddr[11], Daddr
		[10], Daddr[9], Daddr[8], Daddr[7], Daddr[6], Daddr[5], Daddr[4]
		, Daddr[3], Daddr[2], UNCONNECTED_000, UNCONNECTED_001}), .write_sz_in
		(nbus_14524), .write_req_in(write_req_realign), .write_req_out(write_req
		), .write_ack_in(write_ack), .write_ack_out(write_ack_realign), 
		.read_req_in(read_req_realign), .read_req_out(read_req), .read_ack_in
		(read_ack), .read_ack_out(read_ack_realign), .read_data_in(read_data
		), .read_data_out(read_data_realign), .write_data_in(write_data_realign
		), .write_data_out(write_data));
	Itlb i_Itlb(.clk(clk), .rstn(rstn), .addr_phys({code_addr[31], code_addr
		[30], code_addr[29], code_addr[28], code_addr[27], code_addr[26]
		, code_addr[25], code_addr[24], code_addr[23], code_addr[22], code_addr
		[21], code_addr[20], code_addr[19], code_addr[18], code_addr[17]
		, code_addr[16], code_addr[15], code_addr[14], code_addr[13], code_addr
		[12], code_addr[11], code_addr[10], code_addr[9], code_addr[8], code_addr
		[7], code_addr[6], code_addr[5], code_addr[4], code_addr[3], code_addr
		[2], UNCONNECTED_002, UNCONNECTED_003}), .cr3({\cr3[31] , \cr3[30] 
		, \cr3[29] , \cr3[28] , \cr3[27] , \cr3[26] , \cr3[25] , \cr3[24] 
		, \cr3[23] , \cr3[22] , \cr3[21] , \cr3[20] , \cr3[19] , \cr3[18] 
		, \cr3[17] , \cr3[16] , \cr3[15] , \cr3[14] , \cr3[13] , \cr3[12] 
		, UNCONNECTED_004, UNCONNECTED_005, UNCONNECTED_006, 
		UNCONNECTED_007, UNCONNECTED_008, UNCONNECTED_009, 
		UNCONNECTED_010, UNCONNECTED_011, UNCONNECTED_012, 
		UNCONNECTED_013, UNCONNECTED_014, UNCONNECTED_015}), .data_miss(
		{code_data[31], code_data[30], code_data[29], code_data[28], code_data
		[27], code_data[26], code_data[25], code_data[24], code_data[23]
		, code_data[22], code_data[21], code_data[20], code_data[19], code_data
		[18], code_data[17], code_data[16], code_data[15], code_data[14]
		, code_data[13], code_data[12], UNCONNECTED_016, UNCONNECTED_017
		, UNCONNECTED_018, UNCONNECTED_019, code_data[7], code_data[6], code_data
		[5], code_data[4], code_data[3], code_data[2], code_data[1], code_data
		[0]}), .iDaddr(int_code_addr), .pg_en(pg_en), .owrite_data({
		UNCONNECTED_020, UNCONNECTED_021, UNCONNECTED_022, 
		UNCONNECTED_023, UNCONNECTED_024, UNCONNECTED_025, 
		UNCONNECTED_026, UNCONNECTED_027, UNCONNECTED_028, 
		UNCONNECTED_029, UNCONNECTED_030, UNCONNECTED_031, 
		UNCONNECTED_032, UNCONNECTED_033, UNCONNECTED_034, 
		UNCONNECTED_035, UNCONNECTED_036, UNCONNECTED_037, 
		UNCONNECTED_038, UNCONNECTED_039, UNCONNECTED_040, 
		UNCONNECTED_041, UNCONNECTED_042, UNCONNECTED_043, code_wdata[7]
		, code_wdata[6], code_wdata[5], code_wdata[4], code_wdata[3], code_wdata
		[2], code_wdata[1], code_wdata[0]}), .iread_req(int_code_req), .iread_ack
		(code_ack), .iwrite_ack(code_wack), .oread_req(code_req), .oread_ack
		(int_code_ack), .owrite_req(code_wreq), .pg_fault(n_3107), .cr2(icr2
		), .flush_tlb(flush_Itlb), .busy_ram(busy_ram));
	Dtlb i_Dtlb(.clk(clk), .rstn(rstn), .addr_phys(Daddr_realign), .cr3({\cr3[31] 
		, \cr3[30] , \cr3[29] , \cr3[28] , \cr3[27] , \cr3[26] , \cr3[25] 
		, \cr3[24] , \cr3[23] , \cr3[22] , \cr3[21] , \cr3[20] , \cr3[19] 
		, \cr3[18] , \cr3[17] , \cr3[16] , \cr3[15] , \cr3[14] , \cr3[13] 
		, \cr3[12] , UNCONNECTED_044, UNCONNECTED_045, UNCONNECTED_046, 
		UNCONNECTED_047, UNCONNECTED_048, UNCONNECTED_049, 
		UNCONNECTED_050, UNCONNECTED_051, UNCONNECTED_052, 
		UNCONNECTED_053, UNCONNECTED_054, UNCONNECTED_055}), .cr0({
		UNCONNECTED_056, UNCONNECTED_057, UNCONNECTED_058, 
		UNCONNECTED_059, UNCONNECTED_060, UNCONNECTED_061, 
		UNCONNECTED_062, UNCONNECTED_063, UNCONNECTED_064, 
		UNCONNECTED_065, UNCONNECTED_066, UNCONNECTED_067, 
		UNCONNECTED_068, UNCONNECTED_069, UNCONNECTED_070, \cr0[16] , 
		UNCONNECTED_071, UNCONNECTED_072, UNCONNECTED_073, 
		UNCONNECTED_074, UNCONNECTED_075, UNCONNECTED_076, 
		UNCONNECTED_077, UNCONNECTED_078, UNCONNECTED_079, 
		UNCONNECTED_080, UNCONNECTED_081, UNCONNECTED_082, 
		UNCONNECTED_083, UNCONNECTED_084, UNCONNECTED_085, 
		UNCONNECTED_086}), .data_miss(read_data_realign), .iDaddr(int_Daddr
		), .pg_en(pg_en), .iwrite_data(iwrite_data), .owrite_data(write_data_realign
		), .iread_req(int_read_req), .iread_ack(read_ack_realign), .iwrite_req
		(int_write_req), .iwrite_ack(write_ack_realign), .iwrite_sz(int_write_sz
		), .owrite_sz(nbus_14524), .oread_req(read_req_realign), .oread_ack
		(int_read_ack), .owrite_req(write_req_realign), .owrite_ack(int_write_ack
		), .pg_fault(pg_fault), .wr_fault(wr_fault), .cr2(cr2), .flush_tlb
		(flush_Dtlb), .cs({UNCONNECTED_087, UNCONNECTED_088, 
		UNCONNECTED_089, UNCONNECTED_090, UNCONNECTED_091, 
		UNCONNECTED_092, UNCONNECTED_093, UNCONNECTED_094, 
		UNCONNECTED_095, UNCONNECTED_096, UNCONNECTED_097, 
		UNCONNECTED_098, UNCONNECTED_099, UNCONNECTED_100, 
		UNCONNECTED_101, UNCONNECTED_102, UNCONNECTED_103, 
		UNCONNECTED_104, UNCONNECTED_105, UNCONNECTED_106, 
		UNCONNECTED_107, UNCONNECTED_108, UNCONNECTED_109, 
		UNCONNECTED_110, UNCONNECTED_111, UNCONNECTED_112, 
		UNCONNECTED_113, UNCONNECTED_114, UNCONNECTED_115, 
		UNCONNECTED_116, \cs[1] , \cs[0] }), .pt_fault(pt_fault), .busy_ram
		(busy_ram));
	cpu i_cpu(.clk(clk), .rstn(rstn), .iack(iack), .int_cpu(int_main), .ivect
		(ivect), .cr0({UNCONNECTED_117, UNCONNECTED_118, UNCONNECTED_119
		, UNCONNECTED_120, UNCONNECTED_121, UNCONNECTED_122, 
		UNCONNECTED_123, UNCONNECTED_124, UNCONNECTED_125, 
		UNCONNECTED_126, UNCONNECTED_127, UNCONNECTED_128, 
		UNCONNECTED_129, UNCONNECTED_130, UNCONNECTED_131, \cr0[16] , 
		UNCONNECTED_132, UNCONNECTED_133, UNCONNECTED_134, 
		UNCONNECTED_135, UNCONNECTED_136, UNCONNECTED_137, 
		UNCONNECTED_138, UNCONNECTED_139, UNCONNECTED_140, 
		UNCONNECTED_141, UNCONNECTED_142, UNCONNECTED_143, 
		UNCONNECTED_144, UNCONNECTED_145, UNCONNECTED_146, 
		UNCONNECTED_147}), .cr2(cr2), .icr2(icr2), .cr3({\cr3[31] , \cr3[30] 
		, \cr3[29] , \cr3[28] , \cr3[27] , \cr3[26] , \cr3[25] , \cr3[24] 
		, \cr3[23] , \cr3[22] , \cr3[21] , \cr3[20] , \cr3[19] , \cr3[18] 
		, \cr3[17] , \cr3[16] , \cr3[15] , \cr3[14] , \cr3[13] , \cr3[12] 
		, UNCONNECTED_148, UNCONNECTED_149, UNCONNECTED_150, 
		UNCONNECTED_151, UNCONNECTED_152, UNCONNECTED_153, 
		UNCONNECTED_154, UNCONNECTED_155, UNCONNECTED_156, 
		UNCONNECTED_157, UNCONNECTED_158, UNCONNECTED_159}), .cs({
		UNCONNECTED_160, UNCONNECTED_161, UNCONNECTED_162, 
		UNCONNECTED_163, UNCONNECTED_164, UNCONNECTED_165, 
		UNCONNECTED_166, UNCONNECTED_167, UNCONNECTED_168, 
		UNCONNECTED_169, UNCONNECTED_170, UNCONNECTED_171, 
		UNCONNECTED_172, UNCONNECTED_173, UNCONNECTED_174, 
		UNCONNECTED_175, UNCONNECTED_176, UNCONNECTED_177, 
		UNCONNECTED_178, UNCONNECTED_179, UNCONNECTED_180, 
		UNCONNECTED_181, UNCONNECTED_182, UNCONNECTED_183, 
		UNCONNECTED_184, UNCONNECTED_185, UNCONNECTED_186, 
		UNCONNECTED_187, UNCONNECTED_188, UNCONNECTED_189, \cs[1] , \cs[0] 
		}), .pg_fault(pg_fault), .ipg_fault(pc_pg_fault), .useq_ptr(useq_ptr
		), .valid_len(valid_len), .queue(queue), .pg_en(pg_en), .pc_out(pc_out
		), .pc_req(pc_req), .read_req(int_read_req), .write_req(int_write_req
		), .read_ack(int_read_ack), .write_ack(int_write_ack), .flush_Itlb
		(flush_Itlb), .flush_Dtlb(flush_Dtlb), .readio_req(readio_req), 
		.writeio_req(writeio_req), .readio_ack(readio_ack), .writeio_ack
		(writeio_ack), .write_data(iwrite_data), .writeio_data(writeio_data
		), .read_data(read_data_realign), .readio_data(readio_data), .write_sz
		(int_write_sz), .io_add({UNCONNECTED_190, UNCONNECTED_191, 
		UNCONNECTED_192, UNCONNECTED_193, UNCONNECTED_194, 
		UNCONNECTED_195, UNCONNECTED_196, UNCONNECTED_197, 
		UNCONNECTED_198, UNCONNECTED_199, UNCONNECTED_200, 
		UNCONNECTED_201, UNCONNECTED_202, UNCONNECTED_203, 
		UNCONNECTED_204, UNCONNECTED_205, io_add[15], io_add[14], io_add
		[13], io_add[12], io_add[11], io_add[10], io_add[9], io_add[8], io_add
		[7], io_add[6], io_add[5], io_add[4], io_add[3], io_add[2], io_add
		[1], io_add[0]}), .Daddr(int_Daddr), .pt_fault(pt_fault), .wr_fault
		(wr_fault));
	useq i_useq(.iaddr(int_code_addr), .idata(code_data), .code_req(int_code_req
		), .code_ack(int_code_ack), .clk(clk), .rstn(rstn), .useq_ptr(useq_ptr
		), .squeue(queue), .pc_in(pc_out), .pc_req(pc_req), .pg_fault(n_3107
		), .pc_pg_fault(pc_pg_fault), .valid_len(valid_len), .busy_ram(busy_ram
		));
endmodule
module v586(m00_AXI_RSTN, m00_AXI_CLK, m00_AXI_AWADDR, m00_AXI_AWVALID, m00_AXI_AWREADY
		, m00_AXI_AWBURST, m00_AXI_AWLEN, m00_AXI_AWSIZE, m00_AXI_ARADDR
		, m00_AXI_ARVALID, m00_AXI_ARREADY, m00_AXI_ARBURST, m00_AXI_ARLEN
		, m00_AXI_ARSIZE, m00_AXI_WDATA, m00_AXI_WVALID, m00_AXI_WREADY,
		 m00_AXI_WSTRB, m00_AXI_WLAST, m00_AXI_RDATA, m00_AXI_RVALID, m00_AXI_RREADY
		, m00_AXI_RLAST, m00_AXI_BVALID, m00_AXI_BREADY, m01_AXI_AWADDR,
		 m01_AXI_AWVALID, m01_AXI_AWREADY, m01_AXI_AWBURST, m01_AXI_AWLEN
		, m01_AXI_AWSIZE, m01_AXI_ARADDR, m01_AXI_ARVALID, m01_AXI_ARREADY
		, m01_AXI_ARBURST, m01_AXI_ARLEN, m01_AXI_ARSIZE, m01_AXI_WDATA,
		 m01_AXI_WVALID, m01_AXI_WREADY, m01_AXI_WSTRB, m01_AXI_WLAST, m01_AXI_RDATA
		, m01_AXI_RVALID, m01_AXI_RREADY, m01_AXI_RLAST, m01_AXI_BVALID,
		 m01_AXI_BREADY, int_pic, iack, ivect, debug);

	input m00_AXI_RSTN;
	input m00_AXI_CLK;
	output [31:0] m00_AXI_AWADDR;
	output m00_AXI_AWVALID;
	input m00_AXI_AWREADY;
	output [1:0] m00_AXI_AWBURST;
	output [7:0] m00_AXI_AWLEN;
	output [2:0] m00_AXI_AWSIZE;
	output [31:0] m00_AXI_ARADDR;
	output m00_AXI_ARVALID;
	input m00_AXI_ARREADY;
	output [1:0] m00_AXI_ARBURST;
	output [7:0] m00_AXI_ARLEN;
	output [2:0] m00_AXI_ARSIZE;
	output [31:0] m00_AXI_WDATA;
	output m00_AXI_WVALID;
	input m00_AXI_WREADY;
	output [3:0] m00_AXI_WSTRB;
	output m00_AXI_WLAST;
	input [31:0] m00_AXI_RDATA;
	input m00_AXI_RVALID;
	output m00_AXI_RREADY;
	input m00_AXI_RLAST;
	input m00_AXI_BVALID;
	output m00_AXI_BREADY;
	output [31:0] m01_AXI_AWADDR;
	output m01_AXI_AWVALID;
	input m01_AXI_AWREADY;
	output [1:0] m01_AXI_AWBURST;
	output [7:0] m01_AXI_AWLEN;
	output [2:0] m01_AXI_AWSIZE;
	output [31:0] m01_AXI_ARADDR;
	output m01_AXI_ARVALID;
	input m01_AXI_ARREADY;
	output [1:0] m01_AXI_ARBURST;
	output [7:0] m01_AXI_ARLEN;
	output [2:0] m01_AXI_ARSIZE;
	output [31:0] m01_AXI_WDATA;
	output m01_AXI_WVALID;
	input m01_AXI_WREADY;
	output [3:0] m01_AXI_WSTRB;
	output m01_AXI_WLAST;
	input [31:0] m01_AXI_RDATA;
	input m01_AXI_RVALID;
	output m01_AXI_RREADY;
	input m01_AXI_RLAST;
	input m01_AXI_BVALID;
	output m01_AXI_BREADY;
	input int_pic;
	output iack;
	input [7:0] ivect;
	output [4:0] debug;

	wire [3:0] write_msk;
	wire [31:0] writeio_data;
	wire [31:0] readio_data;
	wire [31:0] read_data;
	wire [31:0] write_data;
	wire [127:0] code_data;

	assign m00_AXI_BREADY = 1'b1;
	assign m01_AXI_AWBURST[1] = 1'b0;
	assign m01_AXI_AWBURST[0] = 1'b1;
	assign m01_AXI_AWLEN[7] = 1'b0;
	assign m01_AXI_AWLEN[6] = 1'b0;
	assign m01_AXI_AWLEN[5] = 1'b0;
	assign m01_AXI_AWLEN[4] = 1'b0;
	assign m01_AXI_AWLEN[3] = 1'b0;
	assign m01_AXI_AWLEN[2] = 1'b0;
	assign m01_AXI_AWLEN[1] = 1'b0;
	assign m01_AXI_AWLEN[0] = 1'b0;
	assign m01_AXI_AWSIZE[2] = 1'b0;
	assign m01_AXI_AWSIZE[1] = 1'b1;
	assign m01_AXI_AWSIZE[0] = 1'b0;
	assign m01_AXI_ARBURST[1] = 1'b0;
	assign m01_AXI_ARBURST[0] = 1'b1;
	assign m01_AXI_ARLEN[7] = 1'b0;
	assign m01_AXI_ARLEN[6] = 1'b0;
	assign m01_AXI_ARLEN[5] = 1'b0;
	assign m01_AXI_ARLEN[4] = 1'b0;
	assign m01_AXI_ARLEN[3] = 1'b0;
	assign m01_AXI_ARLEN[2] = 1'b0;
	assign m01_AXI_ARLEN[1] = 1'b0;
	assign m01_AXI_ARLEN[0] = 1'b0;
	assign m01_AXI_ARSIZE[2] = 1'b0;
	assign m01_AXI_ARSIZE[1] = 1'b1;
	assign m01_AXI_ARSIZE[0] = 1'b0;
	assign m01_AXI_WSTRB[3] = 1'b0;
	assign m01_AXI_WSTRB[2] = 1'b0;
	assign m01_AXI_WSTRB[1] = 1'b0;
	assign m01_AXI_WSTRB[0] = 1'b1;


	notech_inv i_15593(.A(n_62346), .Z(n_62348));
	notech_inv i_15592(.A(n_62346), .Z(n_62347));
	notech_inv i_15591(.A(m00_AXI_CLK), .Z(n_62346));
	biu32_axi ubiu(.rstn(m00_AXI_RSTN), .clk(n_62347), .write_req(write_req)
		, .write_ack(write_ack), .write_data(write_data), .write_msk(write_msk
		), .read_req(read_req), .read_ack(read_ack), .read_data(read_data
		), .Daddr({\Daddr[31] , \Daddr[30] , \Daddr[29] , \Daddr[28] , \Daddr[27] 
		, \Daddr[26] , \Daddr[25] , \Daddr[24] , \Daddr[23] , \Daddr[22] 
		, \Daddr[21] , \Daddr[20] , \Daddr[19] , \Daddr[18] , \Daddr[17] 
		, \Daddr[16] , \Daddr[15] , \Daddr[14] , \Daddr[13] , \Daddr[12] 
		, \Daddr[11] , \Daddr[10] , \Daddr[9] , \Daddr[8] , \Daddr[7] , \Daddr[6] 
		, \Daddr[5] , \Daddr[4] , \Daddr[3] , \Daddr[2] , 
		UNCONNECTED_000, UNCONNECTED_001}), .code_req(code_req), .code_ack
		(code_ack), .code_data(code_data), .code_addr({\code_addr[31] , \code_addr[30] 
		, \code_addr[29] , \code_addr[28] , \code_addr[27] , \code_addr[26] 
		, \code_addr[25] , \code_addr[24] , \code_addr[23] , \code_addr[22] 
		, \code_addr[21] , \code_addr[20] , \code_addr[19] , \code_addr[18] 
		, \code_addr[17] , \code_addr[16] , \code_addr[15] , \code_addr[14] 
		, \code_addr[13] , \code_addr[12] , \code_addr[11] , \code_addr[10] 
		, \code_addr[9] , \code_addr[8] , \code_addr[7] , \code_addr[6] 
		, \code_addr[5] , \code_addr[4] , \code_addr[3] , \code_addr[2] 
		, UNCONNECTED_002, UNCONNECTED_003}), .code_wreq(code_wreq), .code_wack
		(code_wack), .code_wdata({UNCONNECTED_004, UNCONNECTED_005, 
		UNCONNECTED_006, UNCONNECTED_007, UNCONNECTED_008, 
		UNCONNECTED_009, UNCONNECTED_010, UNCONNECTED_011, 
		UNCONNECTED_012, UNCONNECTED_013, UNCONNECTED_014, 
		UNCONNECTED_015, UNCONNECTED_016, UNCONNECTED_017, 
		UNCONNECTED_018, UNCONNECTED_019, UNCONNECTED_020, 
		UNCONNECTED_021, UNCONNECTED_022, UNCONNECTED_023, 
		UNCONNECTED_024, UNCONNECTED_025, UNCONNECTED_026, 
		UNCONNECTED_027, \code_wdata[7] , \code_wdata[6] , \code_wdata[5] 
		, \code_wdata[4] , \code_wdata[3] , \code_wdata[2] , \code_wdata[1] 
		, \code_wdata[0] }), .readio_req(readio_req), .writeio_req(writeio_req
		), .readio_ack(readio_ack), .writeio_ack(writeio_ack), .writeio_data
		(writeio_data), .readio_data(readio_data), .io_add({
		UNCONNECTED_028, UNCONNECTED_029, UNCONNECTED_030, 
		UNCONNECTED_031, UNCONNECTED_032, UNCONNECTED_033, 
		UNCONNECTED_034, UNCONNECTED_035, UNCONNECTED_036, 
		UNCONNECTED_037, UNCONNECTED_038, UNCONNECTED_039, 
		UNCONNECTED_040, UNCONNECTED_041, UNCONNECTED_042, 
		UNCONNECTED_043, \io_add[15] , \io_add[14] , \io_add[13] , \io_add[12] 
		, \io_add[11] , \io_add[10] , \io_add[9] , \io_add[8] , \io_add[7] 
		, \io_add[6] , \io_add[5] , \io_add[4] , \io_add[3] , \io_add[2] 
		, \io_add[1] , \io_add[0] }), .axi_AW(m00_AXI_AWADDR), .axi_AWVALID
		(m00_AXI_AWVALID), .axi_AWREADY(m00_AXI_AWREADY), .axi_AWBURST(m00_AXI_AWBURST
		), .axi_AWLEN(m00_AXI_AWLEN), .axi_AWSIZE(m00_AXI_AWSIZE), .axi_W
		(m00_AXI_WDATA), .axi_WVALID(m00_AXI_WVALID), .axi_WREADY(m00_AXI_WREADY
		), .axi_WSTRB(m00_AXI_WSTRB), .axi_WLAST(m00_AXI_WLAST), .axi_AR
		(m00_AXI_ARADDR), .axi_ARVALID(m00_AXI_ARVALID), .axi_ARREADY(m00_AXI_ARREADY
		), .axi_ARBURST(m00_AXI_ARBURST), .axi_ARLEN(m00_AXI_ARLEN), .axi_ARSIZE
		(m00_AXI_ARSIZE), .axi_R(m00_AXI_RDATA), .axi_RVALID(m00_AXI_RVALID
		), .axi_RREADY(m00_AXI_RREADY), .axi_RLAST(m00_AXI_RLAST), .axi_io_AW
		(m01_AXI_AWADDR), .axi_io_AWVALID(m01_AXI_AWVALID), .axi_io_AWREADY
		(m01_AXI_AWREADY), .axi_io_W(m01_AXI_WDATA), .axi_io_WVALID(m01_AXI_WVALID
		), .axi_io_WREADY(m01_AXI_WREADY), .axi_io_WLAST(m01_AXI_WLAST),
		 .axi_io_AR(m01_AXI_ARADDR), .axi_io_ARVALID(m01_AXI_ARVALID), .axi_io_ARREADY
		(m01_AXI_ARREADY), .axi_io_R(m01_AXI_RDATA), .axi_io_RVALID(m01_AXI_RVALID
		), .axi_io_RREADY(m01_AXI_RREADY), .busy(busy_ram));
	core ucore(.clk(n_62348), .rstn(m00_AXI_RSTN), .ivect(ivect), .int_main(int_pic
		), .iack(iack), .code_addr({\code_addr[31] , \code_addr[30] , \code_addr[29] 
		, \code_addr[28] , \code_addr[27] , \code_addr[26] , \code_addr[25] 
		, \code_addr[24] , \code_addr[23] , \code_addr[22] , \code_addr[21] 
		, \code_addr[20] , \code_addr[19] , \code_addr[18] , \code_addr[17] 
		, \code_addr[16] , \code_addr[15] , \code_addr[14] , \code_addr[13] 
		, \code_addr[12] , \code_addr[11] , \code_addr[10] , \code_addr[9] 
		, \code_addr[8] , \code_addr[7] , \code_addr[6] , \code_addr[5] 
		, \code_addr[4] , \code_addr[3] , \code_addr[2] , 
		UNCONNECTED_044, UNCONNECTED_045}), .code_data(code_data), .code_req
		(code_req), .code_ack(code_ack), .code_wreq(code_wreq), .code_wack
		(code_wack), .code_wdata({UNCONNECTED_046, UNCONNECTED_047, 
		UNCONNECTED_048, UNCONNECTED_049, UNCONNECTED_050, 
		UNCONNECTED_051, UNCONNECTED_052, UNCONNECTED_053, 
		UNCONNECTED_054, UNCONNECTED_055, UNCONNECTED_056, 
		UNCONNECTED_057, UNCONNECTED_058, UNCONNECTED_059, 
		UNCONNECTED_060, UNCONNECTED_061, UNCONNECTED_062, 
		UNCONNECTED_063, UNCONNECTED_064, UNCONNECTED_065, 
		UNCONNECTED_066, UNCONNECTED_067, UNCONNECTED_068, 
		UNCONNECTED_069, \code_wdata[7] , \code_wdata[6] , \code_wdata[5] 
		, \code_wdata[4] , \code_wdata[3] , \code_wdata[2] , \code_wdata[1] 
		, \code_wdata[0] }), .readio_data(readio_data), .io_add({
		UNCONNECTED_070, UNCONNECTED_071, UNCONNECTED_072, 
		UNCONNECTED_073, UNCONNECTED_074, UNCONNECTED_075, 
		UNCONNECTED_076, UNCONNECTED_077, UNCONNECTED_078, 
		UNCONNECTED_079, UNCONNECTED_080, UNCONNECTED_081, 
		UNCONNECTED_082, UNCONNECTED_083, UNCONNECTED_084, 
		UNCONNECTED_085, \io_add[15] , \io_add[14] , \io_add[13] , \io_add[12] 
		, \io_add[11] , \io_add[10] , \io_add[9] , \io_add[8] , \io_add[7] 
		, \io_add[6] , \io_add[5] , \io_add[4] , \io_add[3] , \io_add[2] 
		, \io_add[1] , \io_add[0] }), .writeio_data(writeio_data), .writeio_req
		(writeio_req), .readio_req(readio_req), .writeio_ack(writeio_ack
		), .readio_ack(readio_ack), .write_req(write_req), .write_ack(write_ack
		), .write_data(write_data), .write_msk(write_msk), .read_req(read_req
		), .read_ack(read_ack), .read_data(read_data), .Daddr({\Daddr[31] 
		, \Daddr[30] , \Daddr[29] , \Daddr[28] , \Daddr[27] , \Daddr[26] 
		, \Daddr[25] , \Daddr[24] , \Daddr[23] , \Daddr[22] , \Daddr[21] 
		, \Daddr[20] , \Daddr[19] , \Daddr[18] , \Daddr[17] , \Daddr[16] 
		, \Daddr[15] , \Daddr[14] , \Daddr[13] , \Daddr[12] , \Daddr[11] 
		, \Daddr[10] , \Daddr[9] , \Daddr[8] , \Daddr[7] , \Daddr[6] , \Daddr[5] 
		, \Daddr[4] , \Daddr[3] , \Daddr[2] , UNCONNECTED_086, 
		UNCONNECTED_087}), .busy_ram(busy_ram));
endmodule
