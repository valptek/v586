/* verilator lint_off IMPLICIT */
/* verilator lint_off UNDRIVEN */
/* verilator lint_off UNUSED */
/* verilator lint_off UNOPTFLAT */

module psram_axi(MEM_ADDR_OUT, MEM_CEN, MEM_OEN, MEM_WEN, MEM_BEN, MEM_ADV, MEM_CRE
		, MEM_DATA_I, MEM_DATA_O, MEM_DATA_T, s00_axi_aclk, s00_axi_aresetn
		, s00_axi_awid, s00_axi_awaddr, s00_axi_awlen, s00_axi_awsize, s00_axi_awburst
		, s00_axi_awlock, s00_axi_awcache, s00_axi_awprot, s00_axi_awqos
		, s00_axi_awregion, s00_axi_awuser, s00_axi_awvalid, s00_axi_awready
		, s00_axi_wdata, s00_axi_wstrb, s00_axi_wlast, s00_axi_wuser, s00_axi_wvalid
		, s00_axi_wready, s00_axi_bid, s00_axi_bresp, s00_axi_buser, s00_axi_bvalid
		, s00_axi_bready, s00_axi_arid, s00_axi_araddr, s00_axi_arlen, s00_axi_arsize
		, s00_axi_arburst, s00_axi_arlock, s00_axi_arcache, s00_axi_arprot
		, s00_axi_arqos, s00_axi_arregion, s00_axi_aruser, s00_axi_arvalid
		, s00_axi_arready, s00_axi_rid, s00_axi_rdata, s00_axi_rresp, s00_axi_rlast
		, s00_axi_ruser, s00_axi_rvalid, s00_axi_rready);

	output [22:0] MEM_ADDR_OUT;
	output MEM_CEN;
	output MEM_OEN;
	output MEM_WEN;
	output [1:0] MEM_BEN;
	output MEM_ADV;
	output MEM_CRE;
	input [15:0] MEM_DATA_I;
	output [15:0] MEM_DATA_O;
	output [15:0] MEM_DATA_T;
	input s00_axi_aclk;
	input s00_axi_aresetn;
	input [1:0] s00_axi_awid;
	input [23:0] s00_axi_awaddr;
	input [7:0] s00_axi_awlen;
	input [2:0] s00_axi_awsize;
	input [1:0] s00_axi_awburst;
	input s00_axi_awlock;
	input [3:0] s00_axi_awcache;
	input [2:0] s00_axi_awprot;
	input [3:0] s00_axi_awqos;
	input [3:0] s00_axi_awregion;
	input [1:0] s00_axi_awuser;
	input s00_axi_awvalid;
	output s00_axi_awready;
	input [31:0] s00_axi_wdata;
	input [3:0] s00_axi_wstrb;
	input s00_axi_wlast;
	input [1:0] s00_axi_wuser;
	input s00_axi_wvalid;
	output s00_axi_wready;
	output [1:0] s00_axi_bid;
	output [1:0] s00_axi_bresp;
	output [1:0] s00_axi_buser;
	output s00_axi_bvalid;
	input s00_axi_bready;
	input [1:0] s00_axi_arid;
	input [23:0] s00_axi_araddr;
	input [7:0] s00_axi_arlen;
	input [2:0] s00_axi_arsize;
	input [1:0] s00_axi_arburst;
	input s00_axi_arlock;
	input [3:0] s00_axi_arcache;
	input [2:0] s00_axi_arprot;
	input [3:0] s00_axi_arqos;
	input [3:0] s00_axi_arregion;
	input [1:0] s00_axi_aruser;
	input s00_axi_arvalid;
	output s00_axi_arready;
	output [1:0] s00_axi_rid;
	output [31:0] s00_axi_rdata;
	output [1:0] s00_axi_rresp;
	output s00_axi_rlast;
	output [1:0] s00_axi_ruser;
	output s00_axi_rvalid;
	input s00_axi_rready;

	wire [8:0] i_psram_sub_AsyncPSRAMinst_ce_cycle_counter;
	wire [6:0] i_psram_sub_AsyncPSRAMinst_waitcount;
	wire [18:0] i_psram_sub_AsyncPSRAMinst_last_page_read;
	wire [1:0] i_psram_sub_AsyncPSRAMinst_state;
	wire [6:0] i_psram_sub_AsyncPSRAMinst_cycle_time;
	wire [1:0] i_psram_sub_mem_byte_en;
	wire [22:0] i_psram_sub_mem_addr;
	wire [23:0] i_psram_sub_axi_awaddr;
	wire [23:0] i_psram_sub_axi_araddr;
	wire [15:0] i_psram_sub_mem_data_wr;
	wire [23:0] i_psram_sub_function_sub;
	wire [23:0] i_psram_sub_function_sub_0;
	wire [22:0] i_psram_sub_function_plus_2;
	wire [7:0] i_psram_sub_axi_awlen;
	wire [7:0] i_psram_sub_axi_awlen_cntr;
	wire [7:0] i_psram_sub_axi_arlen;
	wire [7:0] i_psram_sub_axi_arlen_cntr;
	wire [2:0] i_psram_sub_state;
	wire [2:0] i_psram_sub_state_5;
	wire \MEM_DATA_T[0] ;

	assign s00_axi_buser[1] = 1'b0;
	assign s00_axi_buser[0] = 1'b0;
	assign s00_axi_ruser[1] = 1'b0;
	assign s00_axi_ruser[0] = 1'b0;

	assign s00_axi_rid[0] = s00_axi_arid[0];
	assign s00_axi_rid[1] = s00_axi_arid[1];
	assign s00_axi_bid[0] = s00_axi_awid[0];
	assign s00_axi_bid[1] = s00_axi_awid[1];
	assign MEM_DATA_T[15] = \MEM_DATA_T[0] ;
	assign MEM_DATA_T[14] = \MEM_DATA_T[0] ;
	assign MEM_DATA_T[13] = \MEM_DATA_T[0] ;
	assign MEM_DATA_T[12] = \MEM_DATA_T[0] ;
	assign MEM_DATA_T[11] = \MEM_DATA_T[0] ;
	assign MEM_DATA_T[10] = \MEM_DATA_T[0] ;
	assign MEM_DATA_T[9] = \MEM_DATA_T[0] ;
	assign MEM_DATA_T[8] = \MEM_DATA_T[0] ;
	assign MEM_DATA_T[7] = \MEM_DATA_T[0] ;
	assign MEM_DATA_T[6] = \MEM_DATA_T[0] ;
	assign MEM_DATA_T[5] = \MEM_DATA_T[0] ;
	assign MEM_DATA_T[4] = \MEM_DATA_T[0] ;
	assign MEM_DATA_T[3] = \MEM_DATA_T[0] ;
	assign MEM_DATA_T[2] = \MEM_DATA_T[0] ;
	assign MEM_DATA_T[1] = \MEM_DATA_T[0] ;
	assign MEM_DATA_T[0] = \MEM_DATA_T[0] ;

	notech_inv i_02687(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[0]), .Z
		(i_psram_sub_AsyncPSRAMinst_n_107));
	notech_nand2 i_12686(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[0]),
		 .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[1]), .Z(n_55));
	notech_nand2 i_22685(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[1]),
		 .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[2]), .Z(n_56));
	notech_nand2 i_32684(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[2]),
		 .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[3]), .Z(n_57));
	notech_nand2 i_42683(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[3]),
		 .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[4]), .Z(n_58));
	notech_nand2 i_52682(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[4]),
		 .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[5]), .Z(n_59));
	notech_nand2 i_62681(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[5]),
		 .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[6]), .Z(n_60));
	notech_nand2 i_72680(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[6]),
		 .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[7]), .Z(n_61));
	notech_inv i_92679(.A(i_psram_sub_AsyncPSRAMinst_n_107), .Z(n_63));
	notech_inv i_102678(.A(n_55), .Z(n_100));
	notech_nor2 i_112677(.A(i_psram_sub_AsyncPSRAMinst_n_107), .B(n_56), .Z(n_65
		));
	notech_nor2 i_122676(.A(n_55), .B(n_57), .Z(n_66));
	notech_nor2 i_132675(.A(n_56), .B(n_58), .Z(n_67));
	notech_nor2 i_142674(.A(n_57), .B(n_59), .Z(n_68));
	notech_nor2 i_152673(.A(n_58), .B(n_60), .Z(n_69));
	notech_nor2 i_162672(.A(n_59), .B(n_61), .Z(n_70));
	notech_nand2 i_222671(.A(n_63), .B(n_67), .Z(n_76));
	notech_nand2 i_232670(.A(n_100), .B(n_68), .Z(n_77));
	notech_nand2 i_242669(.A(n_65), .B(n_69), .Z(n_78));
	notech_nand2 i_252668(.A(n_66), .B(n_70), .Z(n_79));
	notech_inv i_312667(.A(n_76), .Z(n_85));
	notech_inv i_322666(.A(n_77), .Z(n_86));
	notech_inv i_332665(.A(n_78), .Z(n_87));
	notech_inv i_342664(.A(n_79), .Z(n_108));
	notech_xor2 i_372663(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[1]),
		 .B(n_63), .Z(i_psram_sub_AsyncPSRAMinst_n_108));
	notech_xor2 i_382662(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[2]),
		 .B(n_100), .Z(i_psram_sub_AsyncPSRAMinst_n_109));
	notech_xor2 i_392661(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[3]),
		 .B(n_65), .Z(i_psram_sub_AsyncPSRAMinst_n_110));
	notech_xor2 i_402660(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[4]),
		 .B(n_66), .Z(i_psram_sub_AsyncPSRAMinst_n_111));
	notech_xor2 i_412659(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[5]),
		 .B(n_85), .Z(i_psram_sub_AsyncPSRAMinst_n_112));
	notech_xor2 i_422658(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[6]),
		 .B(n_86), .Z(i_psram_sub_AsyncPSRAMinst_n_113));
	notech_xor2 i_432657(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[7]),
		 .B(n_87), .Z(i_psram_sub_AsyncPSRAMinst_n_114));
	notech_xor2 i_442656(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[8]),
		 .B(n_108), .Z(i_psram_sub_AsyncPSRAMinst_n_115));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2606(.A(i_psram_sub_command), .Z
		(i_psram_sub_AsyncPSRAMinst_n_2970));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2605(.A(MEM_OEN), .Z(\MEM_DATA_T[0] 
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2604(.A(MEM_CEN), .Z(i_psram_sub_AsyncPSRAMinst_n_2968
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2603(.A(s00_axi_aresetn), .Z(i_psram_sub_AsyncPSRAMinst_n_2967
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2602(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[7]), .Z(i_psram_sub_AsyncPSRAMinst_n_2966));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2601(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[6]), .Z(i_psram_sub_AsyncPSRAMinst_n_2965));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2600(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[5]), .Z(i_psram_sub_AsyncPSRAMinst_n_2964));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2599(.A(MEM_ADDR_OUT[22]), .Z(i_psram_sub_AsyncPSRAMinst_n_2963
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2598(.A(MEM_ADDR_OUT[21]), .Z(i_psram_sub_AsyncPSRAMinst_n_2962
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2597(.A(MEM_ADDR_OUT[20]), .Z(i_psram_sub_AsyncPSRAMinst_n_2961
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2596(.A(MEM_ADDR_OUT[19]), .Z(i_psram_sub_AsyncPSRAMinst_n_2960
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2595(.A(MEM_ADDR_OUT[18]), .Z(i_psram_sub_AsyncPSRAMinst_n_2959
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2594(.A(MEM_ADDR_OUT[17]), .Z(i_psram_sub_AsyncPSRAMinst_n_2958
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2593(.A(MEM_ADDR_OUT[16]), .Z(i_psram_sub_AsyncPSRAMinst_n_2957
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2592(.A(MEM_ADDR_OUT[15]), .Z(i_psram_sub_AsyncPSRAMinst_n_2956
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2591(.A(MEM_ADDR_OUT[14]), .Z(i_psram_sub_AsyncPSRAMinst_n_2955
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2590(.A(MEM_ADDR_OUT[13]), .Z(i_psram_sub_AsyncPSRAMinst_n_2954
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2589(.A(MEM_ADDR_OUT[12]), .Z(i_psram_sub_AsyncPSRAMinst_n_2953
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2588(.A(MEM_ADDR_OUT[11]), .Z(i_psram_sub_AsyncPSRAMinst_n_2952
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2587(.A(MEM_ADDR_OUT[10]), .Z(i_psram_sub_AsyncPSRAMinst_n_2951
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2586(.A(MEM_ADDR_OUT[9]), .Z(i_psram_sub_AsyncPSRAMinst_n_2950
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2585(.A(MEM_ADDR_OUT[8]), .Z(i_psram_sub_AsyncPSRAMinst_n_2949
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2584(.A(MEM_ADDR_OUT[6]), .Z(i_psram_sub_AsyncPSRAMinst_n_2948
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2583(.A(MEM_ADDR_OUT[5]), .Z(i_psram_sub_AsyncPSRAMinst_n_2947
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2582(.A(MEM_ADDR_OUT[3]), .Z(i_psram_sub_AsyncPSRAMinst_n_2946
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2581(.A(MEM_ADDR_OUT[2]), .Z(i_psram_sub_AsyncPSRAMinst_n_2945
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2580(.A(MEM_ADDR_OUT[1]), .Z(i_psram_sub_AsyncPSRAMinst_n_2944
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2579(.A(MEM_ADDR_OUT[0]), .Z(i_psram_sub_AsyncPSRAMinst_n_2943
		));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2578(.A(i_psram_sub_mem_addr[22]
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2942));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2577(.A(i_psram_sub_mem_addr[21]
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2941));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2576(.A(i_psram_sub_mem_addr[20]
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2940));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2575(.A(i_psram_sub_mem_addr[19]
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2939));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2574(.A(i_psram_sub_mem_addr[18]
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2938));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2573(.A(i_psram_sub_mem_addr[17]
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2937));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2572(.A(i_psram_sub_mem_addr[16]
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2936));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2571(.A(i_psram_sub_mem_addr[15]
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2935));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2570(.A(i_psram_sub_mem_addr[14]
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2934));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2569(.A(i_psram_sub_mem_addr[13]
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2933));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2568(.A(i_psram_sub_mem_addr[12]
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2932));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2567(.A(i_psram_sub_mem_addr[11]
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2931));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2566(.A(i_psram_sub_mem_addr[10]
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2930));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2565(.A(i_psram_sub_mem_addr[9])
		, .Z(i_psram_sub_AsyncPSRAMinst_n_2929));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2564(.A(i_psram_sub_mem_addr[8])
		, .Z(i_psram_sub_AsyncPSRAMinst_n_2928));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2563(.A(i_psram_sub_mem_addr[6])
		, .Z(i_psram_sub_AsyncPSRAMinst_n_2927));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2562(.A(i_psram_sub_mem_addr[5])
		, .Z(i_psram_sub_AsyncPSRAMinst_n_2926));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2561(.A(i_psram_sub_mem_addr[3])
		, .Z(i_psram_sub_AsyncPSRAMinst_n_2925));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2560(.A(i_psram_sub_mem_addr[2])
		, .Z(i_psram_sub_AsyncPSRAMinst_n_2924));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2559(.A(i_psram_sub_mem_addr[1])
		, .Z(i_psram_sub_AsyncPSRAMinst_n_2923));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2558(.A(i_psram_sub_mem_addr[0])
		, .Z(i_psram_sub_AsyncPSRAMinst_n_2922));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2557(.A(i_psram_sub_AsyncPSRAMinst_cen_old
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2921));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2556(.A(i_psram_sub_AsyncPSRAMinst_state
		[1]), .Z(i_psram_sub_AsyncPSRAMinst_n_2920));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2555(.A(i_psram_sub_AsyncPSRAMinst_state
		[0]), .Z(i_psram_sub_AsyncPSRAMinst_n_2919));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2554(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[5]), .Z(i_psram_sub_AsyncPSRAMinst_n_2918));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2553(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[4]), .Z(i_psram_sub_AsyncPSRAMinst_n_2917));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2552(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[3]), .Z(i_psram_sub_AsyncPSRAMinst_n_2916));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2551(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[2]), .Z(i_psram_sub_AsyncPSRAMinst_n_2915));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2550(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[1]), .Z(i_psram_sub_AsyncPSRAMinst_n_2914));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2549(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[0]), .Z(i_psram_sub_AsyncPSRAMinst_n_2913));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2548(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[6]), .Z(i_psram_sub_AsyncPSRAMinst_n_2912));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2547(.A(i_psram_sub_AsyncPSRAMinst_n_549
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2911));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2546(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[5]), .Z(i_psram_sub_AsyncPSRAMinst_n_2910));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2545(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[4]), .Z(i_psram_sub_AsyncPSRAMinst_n_2909));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2544(.A(i_psram_sub_AsyncPSRAMinst_n_539
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2908));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2543(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[3]), .Z(i_psram_sub_AsyncPSRAMinst_n_2907));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2542(.A(i_psram_sub_AsyncPSRAMinst_n_534
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2906));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2541(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[2]), .Z(i_psram_sub_AsyncPSRAMinst_n_2905));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2540(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[1]), .Z(i_psram_sub_AsyncPSRAMinst_n_2904));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2539(.A(i_psram_sub_AsyncPSRAMinst_last_page_read
		[16]), .Z(i_psram_sub_AsyncPSRAMinst_n_2903));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2538(.A(i_psram_sub_AsyncPSRAMinst_last_page_read
		[15]), .Z(i_psram_sub_AsyncPSRAMinst_n_2902));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2537(.A(i_psram_sub_AsyncPSRAMinst_last_page_read
		[11]), .Z(i_psram_sub_AsyncPSRAMinst_n_2901));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2536(.A(i_psram_sub_AsyncPSRAMinst_last_page_read
		[10]), .Z(i_psram_sub_AsyncPSRAMinst_n_2900));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2535(.A(i_psram_sub_AsyncPSRAMinst_n_379
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2899));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2534(.A(i_psram_sub_AsyncPSRAMinst_last_page_read
		[6]), .Z(i_psram_sub_AsyncPSRAMinst_n_2898));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2533(.A(i_psram_sub_AsyncPSRAMinst_last_page_read
		[5]), .Z(i_psram_sub_AsyncPSRAMinst_n_2897));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2532(.A(i_psram_sub_AsyncPSRAMinst_last_page_read
		[1]), .Z(i_psram_sub_AsyncPSRAMinst_n_2896));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2531(.A(i_psram_sub_AsyncPSRAMinst_last_page_read
		[0]), .Z(i_psram_sub_AsyncPSRAMinst_n_2895));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2530(.A(i_psram_sub_AsyncPSRAMinst_n_791
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2894));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2529(.A(i_psram_sub_AsyncPSRAMinst_n_786
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2893));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2528(.A(i_psram_sub_AsyncPSRAMinst_n_781
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2892));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2527(.A(i_psram_sub_AsyncPSRAMinst_n_776
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2891));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2526(.A(i_psram_sub_AsyncPSRAMinst_n_771
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2890));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2525(.A(i_psram_sub_AsyncPSRAMinst_n_766
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2889));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2524(.A(i_psram_sub_AsyncPSRAMinst_n_761
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2888));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2523(.A(i_psram_sub_AsyncPSRAMinst_n_756
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2887));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2522(.A(i_psram_sub_AsyncPSRAMinst_n_751
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2886));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2521(.A(i_psram_sub_AsyncPSRAMinst_n_746
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2885));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2520(.A(i_psram_sub_AsyncPSRAMinst_n_741
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2884));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2519(.A(i_psram_sub_AsyncPSRAMinst_n_736
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2883));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2518(.A(i_psram_sub_AsyncPSRAMinst_n_731
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2882));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2517(.A(i_psram_sub_AsyncPSRAMinst_n_726
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2881));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2516(.A(i_psram_sub_AsyncPSRAMinst_n_721
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2880));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2515(.A(i_psram_sub_AsyncPSRAMinst_n_711
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2879));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2514(.A(i_psram_sub_AsyncPSRAMinst_n_706
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2878));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2513(.A(i_psram_sub_AsyncPSRAMinst_n_696
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2877));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2512(.A(i_psram_sub_AsyncPSRAMinst_n_691
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2876));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2511(.A(i_psram_sub_AsyncPSRAMinst_n_686
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2875));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2510(.A(i_psram_sub_AsyncPSRAMinst_n_681
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2874));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2509(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2873));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2508(.A(i_psram_sub_AsyncPSRAMinst_n_508
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2872));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2507(.A(i_psram_sub_AsyncPSRAMinst_n_505
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2871));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2506(.A(i_psram_sub_AsyncPSRAMinst_n_274
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2870));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2505(.A(i_psram_sub_AsyncPSRAMinst_n_642
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2869));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2504(.A(i_psram_sub_AsyncPSRAMinst_n_568
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2868));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2503(.A(i_psram_sub_AsyncPSRAMinst_n_247
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2867));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2502(.A(i_psram_sub_AsyncPSRAMinst_n_559
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2866));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2501(.A(i_psram_sub_AsyncPSRAMinst_n_446
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2865));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2500(.A(i_psram_sub_AsyncPSRAMinst_n_542
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2864));
	notech_inv i_psram_sub_AsyncPSRAMinst_i_2499(.A(i_psram_sub_AsyncPSRAMinst_n_637
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2863));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_2047(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_BEN[0]), .B(i_psram_sub_AsyncPSRAMinst_n_187), .Z(i_psram_sub_AsyncPSRAMinst_n_2857
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_LBN_reg(.CP(s00_axi_aclk),
		 .D(i_psram_sub_AsyncPSRAMinst_n_2857), .SD(1'b1), .Q(MEM_BEN[0]
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_15(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[15]), .SD(1'b1), .Q(MEM_DATA_O[15]
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_14(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[14]), .SD(1'b1), .Q(MEM_DATA_O[14]
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_13(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[13]), .SD(1'b1), .Q(MEM_DATA_O[13]
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_12(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[12]), .SD(1'b1), .Q(MEM_DATA_O[12]
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_11(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[11]), .SD(1'b1), .Q(MEM_DATA_O[11]
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_10(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[10]), .SD(1'b1), .Q(MEM_DATA_O[10]
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_9(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[9]), .SD(1'b1), .Q(MEM_DATA_O[9])
		);
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_8(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[8]), .SD(1'b1), .Q(MEM_DATA_O[8])
		);
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_7(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[7]), .SD(1'b1), .Q(MEM_DATA_O[7])
		);
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_6(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[6]), .SD(1'b1), .Q(MEM_DATA_O[6])
		);
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_5(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[5]), .SD(1'b1), .Q(MEM_DATA_O[5])
		);
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_4(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[4]), .SD(1'b1), .Q(MEM_DATA_O[4])
		);
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_3(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[3]), .SD(1'b1), .Q(MEM_DATA_O[3])
		);
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_2(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[2]), .SD(1'b1), .Q(MEM_DATA_O[2])
		);
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_1(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[1]), .SD(1'b1), .Q(MEM_DATA_O[1])
		);
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_DATA_O_reg_0(.CP(s00_axi_aclk
		), .D(i_psram_sub_mem_data_wr[0]), .SD(1'b1), .Q(MEM_DATA_O[0])
		);
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1975(.S(i_psram_sub_AsyncPSRAMinst_n_422
		), .A(i_psram_sub_mem_idle), .B(i_psram_sub_AsyncPSRAMinst_n_423
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2819));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_idle_reg(.CP(s00_axi_aclk)
		, .D(i_psram_sub_AsyncPSRAMinst_n_2819), .SD(1'b1), .Q(i_psram_sub_mem_idle
		));
	notech_nao3 i_psram_sub_AsyncPSRAMinst_i_102(.A(s00_axi_aresetn), .B(i_psram_sub_AsyncPSRAMinst_n_2867
		), .C(i_psram_sub_AsyncPSRAMinst_n_232), .Z(\i_psram_sub_AsyncPSRAMinst_state_3[1] 
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1967(.S(i_psram_sub_AsyncPSRAMinst_n_422
		), .A(MEM_CRE), .B(i_psram_sub_AsyncPSRAMinst_n_490), .Z(i_psram_sub_AsyncPSRAMinst_n_2813
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_CRE_reg(.CP(s00_axi_aclk),
		 .D(i_psram_sub_AsyncPSRAMinst_n_2813), .SD(1'b1), .Q(MEM_CRE)
		);
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1959(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_BEN[1]), .B(i_psram_sub_AsyncPSRAMinst_n_443), .Z(i_psram_sub_AsyncPSRAMinst_n_2807
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_UBN_reg(.CP(s00_axi_aclk),
		 .D(i_psram_sub_AsyncPSRAMinst_n_2807), .SD(1'b1), .Q(MEM_BEN[1]
		));
	notech_nao3 i_psram_sub_AsyncPSRAMinst_i_100(.A(s00_axi_aresetn), .B(i_psram_sub_AsyncPSRAMinst_n_235
		), .C(i_psram_sub_AsyncPSRAMinst_n_351), .Z(i_psram_sub_AsyncPSRAMinst_n_187
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1951(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[31] ), .B(i_psram_sub_AsyncPSRAMinst_n_376
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2801));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_15(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2801), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[31] 
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_99(.A(i_psram_sub_AsyncPSRAMinst_state
		[0]), .B(s00_axi_aresetn), .Z(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1943(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[30] ), .B(i_psram_sub_AsyncPSRAMinst_n_374
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2795));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_14(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2795), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[30] 
		));
	notech_nao3 i_psram_sub_AsyncPSRAMinst_i_98(.A(s00_axi_aresetn), .B(i_psram_sub_AsyncPSRAMinst_n_2919
		), .C(i_psram_sub_AsyncPSRAMinst_n_351), .Z(i_psram_sub_AsyncPSRAMinst_n_423
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1935(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[29] ), .B(i_psram_sub_AsyncPSRAMinst_n_373
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2789));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_13(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2789), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[29] 
		));
	notech_nand3 i_psram_sub_AsyncPSRAMinst_i_97(.A(i_psram_sub_AsyncPSRAMinst_state
		[0]), .B(i_psram_sub_AsyncPSRAMinst_n_238), .C(s00_axi_aresetn),
		 .Z(i_psram_sub_AsyncPSRAMinst_n_422));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1927(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[28] ), .B(i_psram_sub_AsyncPSRAMinst_n_372
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2783));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_12(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2783), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[28] 
		));
	notech_nao3 i_psram_sub_AsyncPSRAMinst_i_95(.A(s00_axi_aresetn), .B(i_psram_sub_AsyncPSRAMinst_n_236
		), .C(i_psram_sub_AsyncPSRAMinst_n_351), .Z(i_psram_sub_AsyncPSRAMinst_n_443
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1919(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[27] ), .B(i_psram_sub_AsyncPSRAMinst_n_371
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2777));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_11(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2777), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[27] 
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_93(.A(s00_axi_aresetn), .B(i_psram_sub_AsyncPSRAMinst_n_237
		), .Z(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] ));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1911(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[26] ), .B(i_psram_sub_AsyncPSRAMinst_n_369
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2771));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_10(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2771), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[26] 
		));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_73(.A(i_psram_sub_AsyncPSRAMinst_n_451
		), .B(i_psram_sub_AsyncPSRAMinst_state[0]), .Z(i_psram_sub_AsyncPSRAMinst_n_663
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1903(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[25] ), .B(i_psram_sub_AsyncPSRAMinst_n_368
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2765));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_9(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2765), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[25] 
		));
	notech_nao3 i_psram_sub_AsyncPSRAMinst_i_72(.A(i_psram_sub_command), .B(i_psram_sub_AsyncPSRAMinst_n_2919
		), .C(i_psram_sub_AsyncPSRAMinst_n_498), .Z(i_psram_sub_AsyncPSRAMinst_n_803
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1895(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[24] ), .B(i_psram_sub_AsyncPSRAMinst_n_367
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2759));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_8(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2759), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[24] 
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_69(.A(i_psram_sub_AsyncPSRAMinst_n_379
		), .B(i_psram_sub_AsyncPSRAMinst_n_239), .Z(i_psram_sub_AsyncPSRAMinst_n_194
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1887(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[23] ), .B(i_psram_sub_AsyncPSRAMinst_n_366
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2753));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_7(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2753), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[23] 
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_65(.A(i_psram_sub_AsyncPSRAMinst_n_379
		), .B(i_psram_sub_AsyncPSRAMinst_n_240), .Z(i_psram_sub_AsyncPSRAMinst_n_209
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1879(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[22] ), .B(i_psram_sub_AsyncPSRAMinst_n_364
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2747));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_6(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2747), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[22] 
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_64(.A(i_psram_sub_AsyncPSRAMinst_n_379
		), .B(i_psram_sub_AsyncPSRAMinst_n_241), .Z(i_psram_sub_AsyncPSRAMinst_n_214
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1871(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[21] ), .B(i_psram_sub_AsyncPSRAMinst_n_363
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2741));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_5(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2741), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[21] 
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_63(.A(i_psram_sub_AsyncPSRAMinst_n_379
		), .B(i_psram_sub_AsyncPSRAMinst_n_242), .Z(i_psram_sub_AsyncPSRAMinst_n_219
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1863(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[20] ), .B(i_psram_sub_AsyncPSRAMinst_n_362
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2735));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_4(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2735), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[20] 
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_62(.A(i_psram_sub_AsyncPSRAMinst_n_379
		), .B(i_psram_sub_AsyncPSRAMinst_n_243), .Z(i_psram_sub_AsyncPSRAMinst_n_224
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1855(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[19] ), .B(i_psram_sub_AsyncPSRAMinst_n_361
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2729));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_3(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2729), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[19] 
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_61(.A(i_psram_sub_AsyncPSRAMinst_n_379
		), .B(i_psram_sub_AsyncPSRAMinst_n_244), .Z(i_psram_sub_AsyncPSRAMinst_n_229
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1847(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[18] ), .B(i_psram_sub_AsyncPSRAMinst_n_359
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2723));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_2(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2723), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[18] 
		));
	notech_or4 i_psram_sub_AsyncPSRAMinst_i_59(.A(i_psram_sub_AsyncPSRAMinst_n_2967
		), .B(i_psram_sub_AsyncPSRAMinst_n_383), .C(i_psram_sub_AsyncPSRAMinst_n_382
		), .D(i_psram_sub_AsyncPSRAMinst_n_247), .Z(i_psram_sub_AsyncPSRAMinst_n_564
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1839(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[17] ), .B(i_psram_sub_AsyncPSRAMinst_n_358
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2717));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_1(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2717), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[17] 
		));
	notech_or4 i_psram_sub_AsyncPSRAMinst_i_58(.A(i_psram_sub_AsyncPSRAMinst_state
		[1]), .B(i_psram_sub_AsyncPSRAMinst_n_2919), .C(i_psram_sub_AsyncPSRAMinst_n_2967
		), .D(i_psram_sub_AsyncPSRAMinst_n_2869), .Z(i_psram_sub_AsyncPSRAMinst_n_563
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1831(.S(\i_psram_sub_AsyncPSRAMinst_nbus_19[0] 
		), .A(\i_psram_sub_axi_rdata_0[16] ), .B(i_psram_sub_AsyncPSRAMinst_n_357
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2711));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_data_rd_i_reg_0(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2711), .SD(1'b1), .Q(\i_psram_sub_axi_rdata_0[16] 
		));
	notech_nand3 i_psram_sub_AsyncPSRAMinst_i_57(.A(s00_axi_aresetn), .B(i_psram_sub_AsyncPSRAMinst_n_2920
		), .C(i_psram_sub_AsyncPSRAMinst_n_253), .Z(i_psram_sub_AsyncPSRAMinst_n_473
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1823(.S(i_psram_sub_AsyncPSRAMinst_n_422
		), .A(MEM_WEN), .B(i_psram_sub_AsyncPSRAMinst_n_663), .Z(i_psram_sub_AsyncPSRAMinst_n_2705
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_MEM_WEN_reg(.CP(s00_axi_aclk),
		 .D(i_psram_sub_AsyncPSRAMinst_n_2705), .SD(1'b1), .Q(MEM_WEN)
		);
	notech_or4 i_psram_sub_AsyncPSRAMinst_i_56(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_cem_time_expired), .C(i_psram_sub_AsyncPSRAMinst_n_2863
		), .D(i_psram_sub_AsyncPSRAMinst_n_2970), .Z(i_psram_sub_AsyncPSRAMinst_n_484
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1815(.S(i_psram_sub_AsyncPSRAMinst_n_422
		), .A(MEM_OEN), .B(i_psram_sub_AsyncPSRAMinst_n_803), .Z(i_psram_sub_AsyncPSRAMinst_n_2699
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_oen_i_reg(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2699), .SD(1'b1), .Q(MEM_OEN)
		);
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_55(.A(i_psram_sub_AsyncPSRAMinst_n_522
		), .B(i_psram_sub_AsyncPSRAMinst_n_255), .Z(i_psram_sub_AsyncPSRAMinst_n_519
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1807(.S(MEM_CEN), .A(i_psram_sub_AsyncPSRAMinst_n_2899
		), .B(i_psram_sub_AsyncPSRAMinst_cem_time_expired), .Z(i_psram_sub_AsyncPSRAMinst_n_2693
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_cem_time_expired_reg(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2693), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_cem_time_expired
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_54(.A(s00_axi_aresetn), .B(i_psram_sub_AsyncPSRAMinst_n_493
		), .Z(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] ));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1799(.S(MEM_CEN), .A(i_psram_sub_AsyncPSRAMinst_n_381
		), .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[8]), .Z(i_psram_sub_AsyncPSRAMinst_n_2687
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_ce_cycle_counter_reg_8(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2687), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[8]));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_53(.A(i_psram_sub_AsyncPSRAMinst_n_258
		), .B(i_psram_sub_AsyncPSRAMinst_n_256), .Z(i_psram_sub_AsyncPSRAMinst_n_524
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1791(.S(MEM_CEN), .A(i_psram_sub_AsyncPSRAMinst_n_229
		), .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[7]), .Z(i_psram_sub_AsyncPSRAMinst_n_2681
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_ce_cycle_counter_reg_7(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2681), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[7]));
	notech_nao3 i_psram_sub_AsyncPSRAMinst_i_52(.A(i_psram_sub_AsyncPSRAMinst_n_262
		), .B(i_psram_sub_AsyncPSRAMinst_n_438), .C(i_psram_sub_AsyncPSRAMinst_n_437
		), .Z(i_psram_sub_AsyncPSRAMinst_n_529));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1783(.S(MEM_CEN), .A(i_psram_sub_AsyncPSRAMinst_n_224
		), .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[6]), .Z(i_psram_sub_AsyncPSRAMinst_n_2675
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_ce_cycle_counter_reg_6(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2675), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[6]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_51(.A(i_psram_sub_AsyncPSRAMinst_n_269
		), .B(i_psram_sub_AsyncPSRAMinst_n_2907), .C(i_psram_sub_AsyncPSRAMinst_n_561
		), .D(i_psram_sub_AsyncPSRAMinst_n_555), .Z(i_psram_sub_AsyncPSRAMinst_n_534
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1775(.S(MEM_CEN), .A(i_psram_sub_AsyncPSRAMinst_n_219
		), .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[5]), .Z(i_psram_sub_AsyncPSRAMinst_n_2669
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_ce_cycle_counter_reg_5(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2669), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[5]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_50(.A(i_psram_sub_AsyncPSRAMinst_n_278
		), .B(i_psram_sub_AsyncPSRAMinst_n_2909), .C(i_psram_sub_AsyncPSRAMinst_n_551
		), .D(i_psram_sub_AsyncPSRAMinst_n_553), .Z(i_psram_sub_AsyncPSRAMinst_n_539
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1767(.S(MEM_CEN), .A(i_psram_sub_AsyncPSRAMinst_n_214
		), .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[4]), .Z(i_psram_sub_AsyncPSRAMinst_n_2663
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_ce_cycle_counter_reg_4(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2663), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[4]));
	notech_or4 i_psram_sub_AsyncPSRAMinst_i_49(.A(i_psram_sub_AsyncPSRAMinst_n_450
		), .B(i_psram_sub_AsyncPSRAMinst_n_449), .C(i_psram_sub_AsyncPSRAMinst_n_448
		), .D(i_psram_sub_AsyncPSRAMinst_n_452), .Z(i_psram_sub_AsyncPSRAMinst_n_544
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1759(.S(MEM_CEN), .A(i_psram_sub_AsyncPSRAMinst_n_209
		), .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[3]), .Z(i_psram_sub_AsyncPSRAMinst_n_2657
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_ce_cycle_counter_reg_3(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2657), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[3]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_48(.A(i_psram_sub_AsyncPSRAMinst_n_291
		), .B(i_psram_sub_AsyncPSRAMinst_n_2912), .C(i_psram_sub_AsyncPSRAMinst_n_516
		), .D(i_psram_sub_AsyncPSRAMinst_n_509), .Z(i_psram_sub_AsyncPSRAMinst_n_549
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1751(.S(MEM_CEN), .A(i_psram_sub_AsyncPSRAMinst_n_378
		), .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[2]), .Z(i_psram_sub_AsyncPSRAMinst_n_2651
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_ce_cycle_counter_reg_2(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2651), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[2]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_26(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2922), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2943), .Z(i_psram_sub_AsyncPSRAMinst_n_681
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1743(.S(MEM_CEN), .A(i_psram_sub_AsyncPSRAMinst_n_377
		), .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[1]), .Z(i_psram_sub_AsyncPSRAMinst_n_2645
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_ce_cycle_counter_reg_1(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2645), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[1]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_25(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2923), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2944), .Z(i_psram_sub_AsyncPSRAMinst_n_686
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1735(.S(MEM_CEN), .A(i_psram_sub_AsyncPSRAMinst_n_194
		), .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[0]), .Z(i_psram_sub_AsyncPSRAMinst_n_2639
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_ce_cycle_counter_reg_0(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2639), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[0]));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_cen_old_reg(.CP(s00_axi_aclk),
		 .D(MEM_CEN), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_cen_old)
		);
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_24(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2924), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2945), .Z(i_psram_sub_AsyncPSRAMinst_n_691
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1723(.S(i_psram_sub_AsyncPSRAMinst_n_563
		), .A(MEM_CEN), .B(i_psram_sub_AsyncPSRAMinst_n_564), .Z(i_psram_sub_AsyncPSRAMinst_n_2631
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_cen_i_reg(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2631), .SD(1'b1), .Q(MEM_CEN)
		);
	notech_reg_set i_psram_sub_AsyncPSRAMinst_state_reg_1(.CP(s00_axi_aclk),
		 .D(\i_psram_sub_AsyncPSRAMinst_state_3[1] ), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_state
		[1]));
	notech_nao3 i_psram_sub_AsyncPSRAMinst_i_1716(.A(i_psram_sub_AsyncPSRAMinst_n_664
		), .B(1'b1), .C(i_psram_sub_AsyncPSRAMinst_n_490), .Z(i_psram_sub_AsyncPSRAMinst_n_2628
		));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_state_reg_0(.CP(s00_axi_aclk),
		 .D(i_psram_sub_AsyncPSRAMinst_n_2628), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_state
		[0]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_23(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2925), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2946), .Z(i_psram_sub_AsyncPSRAMinst_n_696
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_1709(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[6]), .B(i_psram_sub_AsyncPSRAMinst_state[0]), .C(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2624));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_cycle_time_reg_6(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2624), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_cycle_time
		[6]));
	notech_nao3 i_psram_sub_AsyncPSRAMinst_i_22(.A(i_psram_sub_AsyncPSRAMinst_n_487
		), .B(i_psram_sub_AsyncPSRAMinst_n_486), .C(i_psram_sub_AsyncPSRAMinst_n_490
		), .Z(i_psram_sub_AsyncPSRAMinst_n_701));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_1701(.A(i_psram_sub_AsyncPSRAMinst_state
		[0]), .B(s00_axi_aresetn), .C(i_psram_sub_AsyncPSRAMinst_cycle_time
		[5]), .Z(i_psram_sub_AsyncPSRAMinst_n_2618));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_cycle_time_reg_5(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2618), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_cycle_time
		[5]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_21(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2926), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2947), .Z(i_psram_sub_AsyncPSRAMinst_n_706
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_1693(.A(i_psram_sub_AsyncPSRAMinst_state
		[0]), .B(s00_axi_aresetn), .C(i_psram_sub_AsyncPSRAMinst_cycle_time
		[4]), .Z(i_psram_sub_AsyncPSRAMinst_n_2612));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_cycle_time_reg_4(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2612), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_cycle_time
		[4]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_20(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2927), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2948), .Z(i_psram_sub_AsyncPSRAMinst_n_711
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_1685(.A(i_psram_sub_AsyncPSRAMinst_state
		[0]), .B(s00_axi_aresetn), .C(i_psram_sub_AsyncPSRAMinst_cycle_time
		[3]), .Z(i_psram_sub_AsyncPSRAMinst_n_2606));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_cycle_time_reg_3(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2606), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_cycle_time
		[3]));
	notech_nao3 i_psram_sub_AsyncPSRAMinst_i_19(.A(i_psram_sub_AsyncPSRAMinst_n_489
		), .B(i_psram_sub_AsyncPSRAMinst_n_488), .C(i_psram_sub_AsyncPSRAMinst_n_490
		), .Z(i_psram_sub_AsyncPSRAMinst_n_716));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1675(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_cycle_time[2]), .B(i_psram_sub_AsyncPSRAMinst_n_484
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2597));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_cycle_time_reg_2(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2597), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_cycle_time
		[2]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_18(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2928), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2949), .Z(i_psram_sub_AsyncPSRAMinst_n_721
		));
	notech_nand3 i_psram_sub_AsyncPSRAMinst_i_1667(.A(i_psram_sub_AsyncPSRAMinst_state
		[0]), .B(s00_axi_aresetn), .C(i_psram_sub_AsyncPSRAMinst_n_2914)
		, .Z(i_psram_sub_AsyncPSRAMinst_n_2591));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_cycle_time_reg_1(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2591), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_cycle_time
		[1]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_17(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2929), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2950), .Z(i_psram_sub_AsyncPSRAMinst_n_726
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1659(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_cycle_time[0]), .B(i_psram_sub_AsyncPSRAMinst_n_473
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2585));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_cycle_time_reg_0(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2585), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_cycle_time
		[0]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_16(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2930), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2951), .Z(i_psram_sub_AsyncPSRAMinst_n_731
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1651(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_waitcount[6]), .B(i_psram_sub_AsyncPSRAMinst_n_2911
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2579));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_waitcount_reg_6(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2579), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_waitcount
		[6]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_15(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2931), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2952), .Z(i_psram_sub_AsyncPSRAMinst_n_736
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1643(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_waitcount[5]), .B(i_psram_sub_AsyncPSRAMinst_n_544
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2573));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_waitcount_reg_5(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2573), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_waitcount
		[5]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_14(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2932), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2953), .Z(i_psram_sub_AsyncPSRAMinst_n_741
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1635(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_waitcount[4]), .B(i_psram_sub_AsyncPSRAMinst_n_2908
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2567));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_waitcount_reg_4(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2567), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_waitcount
		[4]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_13(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2933), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2954), .Z(i_psram_sub_AsyncPSRAMinst_n_746
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1627(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_waitcount[3]), .B(i_psram_sub_AsyncPSRAMinst_n_2906
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2561));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_waitcount_reg_3(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2561), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_waitcount
		[3]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_12(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2934), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2955), .Z(i_psram_sub_AsyncPSRAMinst_n_751
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1619(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_waitcount[2]), .B(i_psram_sub_AsyncPSRAMinst_n_529
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2555));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_waitcount_reg_2(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2555), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_waitcount
		[2]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_11(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2935), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2956), .Z(i_psram_sub_AsyncPSRAMinst_n_756
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1611(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_waitcount[1]), .B(i_psram_sub_AsyncPSRAMinst_n_524
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2549));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_waitcount_reg_1(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2549), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_waitcount
		[1]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_10(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2936), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2957), .Z(i_psram_sub_AsyncPSRAMinst_n_761
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1603(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_waitcount[0]), .B(i_psram_sub_AsyncPSRAMinst_n_519
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2543));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_waitcount_reg_0(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2543), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_waitcount
		[0]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_9(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2937), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2958), .Z(i_psram_sub_AsyncPSRAMinst_n_766
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1595(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[18]), .B(i_psram_sub_AsyncPSRAMinst_n_485
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2537));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_18(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2537), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[18]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_8(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2938), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2959), .Z(i_psram_sub_AsyncPSRAMinst_n_771
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1587(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[17]), .B(i_psram_sub_AsyncPSRAMinst_n_483
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2531));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_17(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2531), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[17]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_7(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2939), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2960), .Z(i_psram_sub_AsyncPSRAMinst_n_776
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1579(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[16]), .B(i_psram_sub_AsyncPSRAMinst_n_482
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2525));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_16(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2525), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[16]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_6(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2940), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2961), .Z(i_psram_sub_AsyncPSRAMinst_n_781
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1571(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[15]), .B(i_psram_sub_AsyncPSRAMinst_n_481
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2519));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_15(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2519), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[15]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_5(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2941), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2962), .Z(i_psram_sub_AsyncPSRAMinst_n_786
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1563(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[14]), .B(i_psram_sub_AsyncPSRAMinst_n_480
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2513));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_14(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2513), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[14]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_4(.A(i_psram_sub_AsyncPSRAMinst_n_498
		), .B(i_psram_sub_AsyncPSRAMinst_n_2942), .C(i_psram_sub_AsyncPSRAMinst_n_497
		), .D(i_psram_sub_AsyncPSRAMinst_n_2963), .Z(i_psram_sub_AsyncPSRAMinst_n_791
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1555(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[13]), .B(i_psram_sub_AsyncPSRAMinst_n_479
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2507));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_13(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2507), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[13]));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_3(.A(i_psram_sub_AsyncPSRAMinst_n_348
		), .B(i_psram_sub_AsyncPSRAMinst_n_349), .Z(i_psram_sub_AsyncPSRAMinst_n_674
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1547(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[12]), .B(i_psram_sub_AsyncPSRAMinst_n_478
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2501));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_12(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2501), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[12]));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_2(.A(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .B(i_psram_sub_AsyncPSRAMinst_n_351), .Z(i_psram_sub_AsyncPSRAMinst_n_673
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1539(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[11]), .B(i_psram_sub_AsyncPSRAMinst_n_477
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2495));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_11(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2495), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[11]));
	notech_nao3 i_psram_sub_AsyncPSRAMinst_i_1(.A(s00_axi_aresetn), .B(i_psram_sub_AsyncPSRAMinst_n_352
		), .C(i_psram_sub_AsyncPSRAMinst_n_351), .Z(i_psram_sub_AsyncPSRAMinst_n_451
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1531(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[10]), .B(i_psram_sub_AsyncPSRAMinst_n_476
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2489));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_10(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2489), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[10]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_400(.A(i_psram_sub_AsyncPSRAMinst_state
		[0]), .B(i_psram_sub_AsyncPSRAMinst_n_500), .C(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .D(i_psram_sub_AsyncPSRAMinst_n_233), .Z(i_psram_sub_AsyncPSRAMinst_n_664
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1523(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[9]), .B(i_psram_sub_AsyncPSRAMinst_n_475
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2483));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_9(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2483), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[9]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1515(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[8]), .B(i_psram_sub_AsyncPSRAMinst_n_474
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2477));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_8(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2477), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[8]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1507(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[7]), .B(i_psram_sub_AsyncPSRAMinst_n_472
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2471));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_7(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2471), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[7]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1499(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[6]), .B(i_psram_sub_AsyncPSRAMinst_n_471
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2465));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_6(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2465), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[6]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1491(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[5]), .B(i_psram_sub_AsyncPSRAMinst_n_470
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2459));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_5(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2459), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[5]));
	notech_or4 i_psram_sub_AsyncPSRAMinst_i_121(.A(i_psram_sub_AsyncPSRAMinst_n_657
		), .B(i_psram_sub_AsyncPSRAMinst_n_652), .C(i_psram_sub_AsyncPSRAMinst_n_2965
		), .D(i_psram_sub_AsyncPSRAMinst_n_2964), .Z(i_psram_sub_AsyncPSRAMinst_n_658
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1483(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[4]), .B(i_psram_sub_AsyncPSRAMinst_n_469
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2453));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_4(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2453), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[4]));
	notech_or4 i_psram_sub_AsyncPSRAMinst_i_426(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[2]), .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[1]), .C(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[8]), .D(i_psram_sub_AsyncPSRAMinst_n_2966), .Z(i_psram_sub_AsyncPSRAMinst_n_657
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1475(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[3]), .B(i_psram_sub_AsyncPSRAMinst_n_468
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2447));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_3(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2447), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[3]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1467(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[2]), .B(i_psram_sub_AsyncPSRAMinst_n_467
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2441));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_2(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2441), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[2]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1459(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[1]), .B(i_psram_sub_AsyncPSRAMinst_n_466
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2435));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_1(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2435), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[1]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1451(.S(\i_psram_sub_AsyncPSRAMinst_nbus_15[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_last_page_read[0]), .B(i_psram_sub_AsyncPSRAMinst_n_465
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2429));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_last_page_read_reg_0(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2429), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_last_page_read
		[0]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1443(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[22]), .B(i_psram_sub_AsyncPSRAMinst_n_2894), 
		.Z(i_psram_sub_AsyncPSRAMinst_n_2423));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_22(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2423), .SD(1'b1), .Q(MEM_ADDR_OUT
		[22]));
	notech_nand3 i_psram_sub_AsyncPSRAMinst_i_429(.A(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[3]), .B(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter[0]), .C(i_psram_sub_AsyncPSRAMinst_ce_cycle_counter
		[4]), .Z(i_psram_sub_AsyncPSRAMinst_n_652));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1435(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[21]), .B(i_psram_sub_AsyncPSRAMinst_n_2893), 
		.Z(i_psram_sub_AsyncPSRAMinst_n_2417));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_21(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2417), .SD(1'b1), .Q(MEM_ADDR_OUT
		[21]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1427(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[20]), .B(i_psram_sub_AsyncPSRAMinst_n_2892), 
		.Z(i_psram_sub_AsyncPSRAMinst_n_2411));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_20(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2411), .SD(1'b1), .Q(MEM_ADDR_OUT
		[20]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1419(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[19]), .B(i_psram_sub_AsyncPSRAMinst_n_2891), 
		.Z(i_psram_sub_AsyncPSRAMinst_n_2405));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_19(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2405), .SD(1'b1), .Q(MEM_ADDR_OUT
		[19]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1411(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[18]), .B(i_psram_sub_AsyncPSRAMinst_n_2890), 
		.Z(i_psram_sub_AsyncPSRAMinst_n_2399));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_18(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2399), .SD(1'b1), .Q(MEM_ADDR_OUT
		[18]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1403(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[17]), .B(i_psram_sub_AsyncPSRAMinst_n_2889), 
		.Z(i_psram_sub_AsyncPSRAMinst_n_2393));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_17(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2393), .SD(1'b1), .Q(MEM_ADDR_OUT
		[17]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1395(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[16]), .B(i_psram_sub_AsyncPSRAMinst_n_2888), 
		.Z(i_psram_sub_AsyncPSRAMinst_n_2387));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_16(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2387), .SD(1'b1), .Q(MEM_ADDR_OUT
		[16]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1387(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[15]), .B(i_psram_sub_AsyncPSRAMinst_n_2887), 
		.Z(i_psram_sub_AsyncPSRAMinst_n_2381));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_15(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2381), .SD(1'b1), .Q(MEM_ADDR_OUT
		[15]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1379(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[14]), .B(i_psram_sub_AsyncPSRAMinst_n_2886), 
		.Z(i_psram_sub_AsyncPSRAMinst_n_2375));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_14(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2375), .SD(1'b1), .Q(MEM_ADDR_OUT
		[14]));
	notech_or4 i_psram_sub_AsyncPSRAMinst_i_133(.A(i_psram_sub_AsyncPSRAMinst_n_386
		), .B(i_psram_sub_AsyncPSRAMinst_n_384), .C(i_psram_sub_AsyncPSRAMinst_n_436
		), .D(i_psram_sub_AsyncPSRAMinst_n_568), .Z(i_psram_sub_AsyncPSRAMinst_n_642
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1371(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[13]), .B(i_psram_sub_AsyncPSRAMinst_n_2885), 
		.Z(i_psram_sub_AsyncPSRAMinst_n_2369));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_13(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2369), .SD(1'b1), .Q(MEM_ADDR_OUT
		[13]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1363(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[12]), .B(i_psram_sub_AsyncPSRAMinst_n_2884), 
		.Z(i_psram_sub_AsyncPSRAMinst_n_2363));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_12(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2363), .SD(1'b1), .Q(MEM_ADDR_OUT
		[12]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1355(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[11]), .B(i_psram_sub_AsyncPSRAMinst_n_2883), 
		.Z(i_psram_sub_AsyncPSRAMinst_n_2357));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_11(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2357), .SD(1'b1), .Q(MEM_ADDR_OUT
		[11]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1347(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[10]), .B(i_psram_sub_AsyncPSRAMinst_n_2882), 
		.Z(i_psram_sub_AsyncPSRAMinst_n_2351));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_10(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2351), .SD(1'b1), .Q(MEM_ADDR_OUT
		[10]));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_104(.A(i_psram_sub_AsyncPSRAMinst_n_634
		), .B(i_psram_sub_AsyncPSRAMinst_n_624), .C(i_psram_sub_AsyncPSRAMinst_n_612
		), .D(i_psram_sub_AsyncPSRAMinst_n_601), .Z(i_psram_sub_AsyncPSRAMinst_n_637
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1339(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[9]), .B(i_psram_sub_AsyncPSRAMinst_n_2881), .Z
		(i_psram_sub_AsyncPSRAMinst_n_2345));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_9(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2345), .SD(1'b1), .Q(MEM_ADDR_OUT
		[9]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1331(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[8]), .B(i_psram_sub_AsyncPSRAMinst_n_2880), .Z
		(i_psram_sub_AsyncPSRAMinst_n_2339));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_8(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2339), .SD(1'b1), .Q(MEM_ADDR_OUT
		[8]));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_447(.A(i_psram_sub_AsyncPSRAMinst_page_valid
		), .B(i_psram_sub_AsyncPSRAMinst_n_631), .C(i_psram_sub_AsyncPSRAMinst_n_387
		), .D(i_psram_sub_AsyncPSRAMinst_n_629), .Z(i_psram_sub_AsyncPSRAMinst_n_634
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1323(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[7]), .B(i_psram_sub_AsyncPSRAMinst_n_716), .Z
		(i_psram_sub_AsyncPSRAMinst_n_2333));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_7(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2333), .SD(1'b1), .Q(MEM_ADDR_OUT
		[7]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1315(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[6]), .B(i_psram_sub_AsyncPSRAMinst_n_2879), .Z
		(i_psram_sub_AsyncPSRAMinst_n_2327));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_6(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2327), .SD(1'b1), .Q(MEM_ADDR_OUT
		[6]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1307(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[5]), .B(i_psram_sub_AsyncPSRAMinst_n_2878), .Z
		(i_psram_sub_AsyncPSRAMinst_n_2321));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_5(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2321), .SD(1'b1), .Q(MEM_ADDR_OUT
		[5]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_441(.A(i_psram_sub_mem_addr[4]),
		 .B(i_psram_sub_AsyncPSRAMinst_n_2895), .C(i_psram_sub_AsyncPSRAMinst_n_2926
		), .D(i_psram_sub_AsyncPSRAMinst_last_page_read[1]), .Z(i_psram_sub_AsyncPSRAMinst_n_631
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1299(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[4]), .B(i_psram_sub_AsyncPSRAMinst_n_701), .Z
		(i_psram_sub_AsyncPSRAMinst_n_2315));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_4(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2315), .SD(1'b1), .Q(MEM_ADDR_OUT
		[4]));
	notech_ao3 i_psram_sub_AsyncPSRAMinst_i_446(.A(i_psram_sub_AsyncPSRAMinst_n_628
		), .B(i_psram_sub_AsyncPSRAMinst_n_396), .C(i_psram_sub_AsyncPSRAMinst_n_626
		), .Z(i_psram_sub_AsyncPSRAMinst_n_629));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1291(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[3]), .B(i_psram_sub_AsyncPSRAMinst_n_2877), .Z
		(i_psram_sub_AsyncPSRAMinst_n_2309));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_3(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2309), .SD(1'b1), .Q(MEM_ADDR_OUT
		[3]));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_443(.A(i_psram_sub_mem_addr[5]),
		 .B(i_psram_sub_AsyncPSRAMinst_n_2896), .C(i_psram_sub_AsyncPSRAMinst_last_page_read
		[2]), .D(i_psram_sub_AsyncPSRAMinst_n_2927), .Z(i_psram_sub_AsyncPSRAMinst_n_628
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1283(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[2]), .B(i_psram_sub_AsyncPSRAMinst_n_2876), .Z
		(i_psram_sub_AsyncPSRAMinst_n_2303));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_2(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2303), .SD(1'b1), .Q(MEM_ADDR_OUT
		[2]));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1275(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[1]), .B(i_psram_sub_AsyncPSRAMinst_n_2875), .Z
		(i_psram_sub_AsyncPSRAMinst_n_2297));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_1(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2297), .SD(1'b1), .Q(MEM_ADDR_OUT
		[1]));
	notech_xor2 i_psram_sub_AsyncPSRAMinst_i_444(.A(i_psram_sub_mem_addr[7])
		, .B(i_psram_sub_AsyncPSRAMinst_last_page_read[3]), .Z(i_psram_sub_AsyncPSRAMinst_n_626
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1267(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(MEM_ADDR_OUT[0]), .B(i_psram_sub_AsyncPSRAMinst_n_2874), .Z
		(i_psram_sub_AsyncPSRAMinst_n_2291));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_mem_addr_out_i_reg_0(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2291), .SD(1'b1), .Q(MEM_ADDR_OUT
		[0]));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_456(.A(i_psram_sub_AsyncPSRAMinst_n_619
		), .B(i_psram_sub_AsyncPSRAMinst_n_402), .C(i_psram_sub_AsyncPSRAMinst_n_622
		), .D(i_psram_sub_AsyncPSRAMinst_n_618), .Z(i_psram_sub_AsyncPSRAMinst_n_624
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1259(.S(i_psram_sub_AsyncPSRAMinst_n_673
		), .A(i_psram_sub_AsyncPSRAMinst_page_valid), .B(i_psram_sub_AsyncPSRAMinst_n_674
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2285));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_page_valid_reg(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2285), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_page_valid
		));
	notech_mux2 i_psram_sub_AsyncPSRAMinst_i_1251(.S(\i_psram_sub_AsyncPSRAMinst_nbus_16[0] 
		), .A(i_psram_sub_AsyncPSRAMinst_current_cmd), .B(i_psram_sub_AsyncPSRAMinst_n_451
		), .Z(i_psram_sub_AsyncPSRAMinst_n_2279));
	notech_reg_set i_psram_sub_AsyncPSRAMinst_current_cmd_reg(.CP(s00_axi_aclk
		), .D(i_psram_sub_AsyncPSRAMinst_n_2279), .SD(1'b1), .Q(i_psram_sub_AsyncPSRAMinst_current_cmd
		));
	notech_xor2 i_psram_sub_AsyncPSRAMinst_i_448(.A(i_psram_sub_AsyncPSRAMinst_n_2928
		), .B(i_psram_sub_AsyncPSRAMinst_last_page_read[4]), .Z(i_psram_sub_AsyncPSRAMinst_n_622
		));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_449(.A(i_psram_sub_mem_addr[9]),
		 .B(i_psram_sub_AsyncPSRAMinst_n_2897), .C(i_psram_sub_AsyncPSRAMinst_n_2930
		), .D(i_psram_sub_AsyncPSRAMinst_last_page_read[6]), .Z(i_psram_sub_AsyncPSRAMinst_n_619
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_455(.A(i_psram_sub_AsyncPSRAMinst_n_617
		), .B(i_psram_sub_AsyncPSRAMinst_n_408), .C(i_psram_sub_AsyncPSRAMinst_n_614
		), .Z(i_psram_sub_AsyncPSRAMinst_n_618));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_452(.A(i_psram_sub_mem_addr[10])
		, .B(i_psram_sub_AsyncPSRAMinst_n_2898), .C(i_psram_sub_AsyncPSRAMinst_last_page_read
		[7]), .D(i_psram_sub_AsyncPSRAMinst_n_2931), .Z(i_psram_sub_AsyncPSRAMinst_n_617
		));
	notech_xor2 i_psram_sub_AsyncPSRAMinst_i_453(.A(i_psram_sub_AsyncPSRAMinst_n_2932
		), .B(i_psram_sub_AsyncPSRAMinst_last_page_read[8]), .Z(i_psram_sub_AsyncPSRAMinst_n_614
		));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_466(.A(i_psram_sub_AsyncPSRAMinst_n_607
		), .B(i_psram_sub_AsyncPSRAMinst_n_414), .C(i_psram_sub_AsyncPSRAMinst_n_609
		), .D(i_psram_sub_AsyncPSRAMinst_n_606), .Z(i_psram_sub_AsyncPSRAMinst_n_612
		));
	notech_xor2 i_psram_sub_AsyncPSRAMinst_i_458(.A(i_psram_sub_AsyncPSRAMinst_n_2933
		), .B(i_psram_sub_AsyncPSRAMinst_last_page_read[9]), .Z(i_psram_sub_AsyncPSRAMinst_n_609
		));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_459(.A(i_psram_sub_mem_addr[14])
		, .B(i_psram_sub_AsyncPSRAMinst_n_2900), .C(i_psram_sub_AsyncPSRAMinst_n_2935
		), .D(i_psram_sub_AsyncPSRAMinst_last_page_read[11]), .Z(i_psram_sub_AsyncPSRAMinst_n_607
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_465(.A(i_psram_sub_AsyncPSRAMinst_n_604
		), .B(i_psram_sub_AsyncPSRAMinst_n_419), .C(i_psram_sub_AsyncPSRAMinst_n_602
		), .Z(i_psram_sub_AsyncPSRAMinst_n_606));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_462(.A(i_psram_sub_mem_addr[15])
		, .B(i_psram_sub_AsyncPSRAMinst_n_2901), .C(i_psram_sub_AsyncPSRAMinst_last_page_read
		[12]), .D(i_psram_sub_AsyncPSRAMinst_n_2936), .Z(i_psram_sub_AsyncPSRAMinst_n_604
		));
	notech_xor2 i_psram_sub_AsyncPSRAMinst_i_463(.A(i_psram_sub_AsyncPSRAMinst_n_2937
		), .B(i_psram_sub_AsyncPSRAMinst_last_page_read[13]), .Z(i_psram_sub_AsyncPSRAMinst_n_602
		));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_475(.A(i_psram_sub_AsyncPSRAMinst_n_596
		), .B(i_psram_sub_AsyncPSRAMinst_n_426), .C(i_psram_sub_AsyncPSRAMinst_n_598
		), .D(i_psram_sub_AsyncPSRAMinst_n_594), .Z(i_psram_sub_AsyncPSRAMinst_n_601
		));
	notech_xor2 i_psram_sub_AsyncPSRAMinst_i_467(.A(i_psram_sub_AsyncPSRAMinst_n_2938
		), .B(i_psram_sub_AsyncPSRAMinst_last_page_read[14]), .Z(i_psram_sub_AsyncPSRAMinst_n_598
		));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_468(.A(i_psram_sub_mem_addr[19])
		, .B(i_psram_sub_AsyncPSRAMinst_n_2902), .C(i_psram_sub_AsyncPSRAMinst_n_2940
		), .D(i_psram_sub_AsyncPSRAMinst_last_page_read[16]), .Z(i_psram_sub_AsyncPSRAMinst_n_596
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_474(.A(i_psram_sub_AsyncPSRAMinst_n_593
		), .B(i_psram_sub_AsyncPSRAMinst_n_431), .C(i_psram_sub_AsyncPSRAMinst_n_591
		), .Z(i_psram_sub_AsyncPSRAMinst_n_594));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_471(.A(i_psram_sub_mem_addr[20])
		, .B(i_psram_sub_AsyncPSRAMinst_n_2903), .C(i_psram_sub_AsyncPSRAMinst_last_page_read
		[17]), .D(i_psram_sub_AsyncPSRAMinst_n_2941), .Z(i_psram_sub_AsyncPSRAMinst_n_593
		));
	notech_xor2 i_psram_sub_AsyncPSRAMinst_i_472(.A(i_psram_sub_AsyncPSRAMinst_n_2942
		), .B(i_psram_sub_AsyncPSRAMinst_last_page_read[18]), .Z(i_psram_sub_AsyncPSRAMinst_n_591
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_116(.A(i_psram_sub_AsyncPSRAMinst_n_2866
		), .B(i_psram_sub_AsyncPSRAMinst_n_586), .C(i_psram_sub_AsyncPSRAMinst_n_432
		), .Z(i_psram_sub_AsyncPSRAMinst_n_588));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_478(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[2]), .B(i_psram_sub_AsyncPSRAMinst_n_2915), .C(i_psram_sub_AsyncPSRAMinst_n_2916
		), .D(i_psram_sub_AsyncPSRAMinst_waitcount[3]), .Z(i_psram_sub_AsyncPSRAMinst_n_586
		));
	notech_nand3 i_psram_sub_AsyncPSRAMinst_i_110(.A(i_psram_sub_AsyncPSRAMinst_n_441
		), .B(i_psram_sub_AsyncPSRAMinst_n_433), .C(i_psram_sub_AsyncPSRAMinst_n_2866
		), .Z(i_psram_sub_AsyncPSRAMinst_n_568));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_497(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[3]), .B(i_psram_sub_AsyncPSRAMinst_n_2913), .Z(i_psram_sub_AsyncPSRAMinst_n_562
		));
	notech_nao3 i_psram_sub_AsyncPSRAMinst_i_499(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[0]), .B(s00_axi_aresetn), .C(i_psram_sub_AsyncPSRAMinst_n_442),
		 .Z(i_psram_sub_AsyncPSRAMinst_n_561));
	notech_or4 i_psram_sub_AsyncPSRAMinst_i_105(.A(i_psram_sub_AsyncPSRAMinst_n_2864
		), .B(i_psram_sub_AsyncPSRAMinst_n_444), .C(i_psram_sub_AsyncPSRAMinst_n_445
		), .D(i_psram_sub_AsyncPSRAMinst_n_2865), .Z(i_psram_sub_AsyncPSRAMinst_n_559
		));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_137(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[0]), .B(s00_axi_aresetn), .Z(i_psram_sub_AsyncPSRAMinst_n_556)
		);
	notech_nand3 i_psram_sub_AsyncPSRAMinst_i_500(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[2]), .B(i_psram_sub_AsyncPSRAMinst_waitcount[1]), .C(i_psram_sub_AsyncPSRAMinst_n_2907
		), .Z(i_psram_sub_AsyncPSRAMinst_n_555));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_505(.A(i_psram_sub_AsyncPSRAMinst_n_507
		), .B(i_psram_sub_AsyncPSRAMinst_n_447), .Z(i_psram_sub_AsyncPSRAMinst_n_553
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_506(.A(s00_axi_aresetn), .B(i_psram_sub_AsyncPSRAMinst_n_2909
		), .Z(i_psram_sub_AsyncPSRAMinst_n_551));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_513(.A(i_psram_sub_AsyncPSRAMinst_n_2864
		), .B(i_psram_sub_AsyncPSRAMinst_n_2916), .Z(i_psram_sub_AsyncPSRAMinst_n_543
		));
	notech_xor2 i_psram_sub_AsyncPSRAMinst_i_103(.A(i_psram_sub_AsyncPSRAMinst_n_2912
		), .B(i_psram_sub_AsyncPSRAMinst_cycle_time[6]), .Z(i_psram_sub_AsyncPSRAMinst_n_542
		));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_516(.A(i_psram_sub_AsyncPSRAMinst_n_2872
		), .B(i_psram_sub_AsyncPSRAMinst_cycle_time[6]), .C(i_psram_sub_AsyncPSRAMinst_waitcount
		[5]), .D(i_psram_sub_AsyncPSRAMinst_n_293), .Z(i_psram_sub_AsyncPSRAMinst_n_538
		));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_517(.A(i_psram_sub_AsyncPSRAMinst_n_294
		), .B(i_psram_sub_AsyncPSRAMinst_waitcount[4]), .C(i_psram_sub_AsyncPSRAMinst_n_507
		), .D(i_psram_sub_AsyncPSRAMinst_n_446), .Z(i_psram_sub_AsyncPSRAMinst_n_533
		));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_115(.A(i_psram_sub_AsyncPSRAMinst_n_463
		), .B(i_psram_sub_AsyncPSRAMinst_n_441), .C(i_psram_sub_AsyncPSRAMinst_n_462
		), .D(i_psram_sub_AsyncPSRAMinst_n_461), .Z(i_psram_sub_AsyncPSRAMinst_n_532
		));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_518(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[3]), .B(i_psram_sub_AsyncPSRAMinst_n_295), .C(i_psram_sub_AsyncPSRAMinst_n_2871
		), .D(i_psram_sub_AsyncPSRAMinst_n_441), .Z(i_psram_sub_AsyncPSRAMinst_n_530
		));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_130(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[2]), .B(i_psram_sub_AsyncPSRAMinst_n_299), .C(i_psram_sub_AsyncPSRAMinst_waitcount
		[1]), .D(i_psram_sub_AsyncPSRAMinst_n_297), .Z(i_psram_sub_AsyncPSRAMinst_n_526
		));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_134(.A(i_psram_sub_AsyncPSRAMinst_n_231
		), .B(i_psram_sub_AsyncPSRAMinst_n_518), .Z(i_psram_sub_AsyncPSRAMinst_n_522
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_107(.A(i_psram_sub_AsyncPSRAMinst_n_463
		), .B(i_psram_sub_AsyncPSRAMinst_n_441), .C(i_psram_sub_AsyncPSRAMinst_n_462
		), .Z(i_psram_sub_AsyncPSRAMinst_n_521));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_119(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[0]), .B(i_psram_sub_AsyncPSRAMinst_n_2967), .Z(i_psram_sub_AsyncPSRAMinst_n_518
		));
	notech_nao3 i_psram_sub_AsyncPSRAMinst_i_528(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[5]), .B(s00_axi_aresetn), .C(i_psram_sub_AsyncPSRAMinst_n_464),
		 .Z(i_psram_sub_AsyncPSRAMinst_n_516));
	notech_nor2 i_psram_sub_AsyncPSRAMinst_i_530(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[6]), .B(i_psram_sub_AsyncPSRAMinst_n_514), .Z(i_psram_sub_AsyncPSRAMinst_n_515
		));
	notech_nand3 i_psram_sub_AsyncPSRAMinst_i_117(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[1]), .B(i_psram_sub_AsyncPSRAMinst_cycle_time[0]), .C(i_psram_sub_AsyncPSRAMinst_cycle_time
		[2]), .Z(i_psram_sub_AsyncPSRAMinst_n_514));
	notech_nand3 i_psram_sub_AsyncPSRAMinst_i_529(.A(i_psram_sub_AsyncPSRAMinst_n_507
		), .B(i_psram_sub_AsyncPSRAMinst_waitcount[4]), .C(i_psram_sub_AsyncPSRAMinst_n_2912
		), .Z(i_psram_sub_AsyncPSRAMinst_n_509));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_114(.A(i_psram_sub_AsyncPSRAMinst_n_507
		), .B(i_psram_sub_AsyncPSRAMinst_waitcount[4]), .Z(i_psram_sub_AsyncPSRAMinst_n_508
		));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_106(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[0]), .B(i_psram_sub_AsyncPSRAMinst_waitcount[2]), .C(i_psram_sub_AsyncPSRAMinst_waitcount
		[1]), .D(i_psram_sub_AsyncPSRAMinst_waitcount[3]), .Z(i_psram_sub_AsyncPSRAMinst_n_507
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_113(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[2]), .B(i_psram_sub_AsyncPSRAMinst_waitcount[1]), .Z(i_psram_sub_AsyncPSRAMinst_n_505
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_136(.A(i_psram_sub_go), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_500));
	notech_nand3 i_psram_sub_AsyncPSRAMinst_i_131(.A(i_psram_sub_go), .B(s00_axi_aresetn
		), .C(i_psram_sub_AsyncPSRAMinst_n_2920), .Z(i_psram_sub_AsyncPSRAMinst_n_498
		));
	notech_nao3 i_psram_sub_AsyncPSRAMinst_i_132(.A(s00_axi_aresetn), .B(i_psram_sub_AsyncPSRAMinst_n_2920
		), .C(i_psram_sub_go), .Z(i_psram_sub_AsyncPSRAMinst_n_497));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_139(.A(i_psram_sub_AsyncPSRAMinst_state
		[0]), .B(i_psram_sub_AsyncPSRAMinst_n_2920), .Z(i_psram_sub_AsyncPSRAMinst_n_493
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_140(.A(i_psram_sub_AsyncPSRAMinst_cem_time_expired
		), .B(i_psram_sub_AsyncPSRAMinst_n_2968), .Z(i_psram_sub_AsyncPSRAMinst_n_491
		));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_96(.A(i_psram_sub_AsyncPSRAMinst_state
		[1]), .B(s00_axi_aresetn), .Z(i_psram_sub_AsyncPSRAMinst_n_490)
		);
	notech_nand3 i_psram_sub_AsyncPSRAMinst_i_341(.A(i_psram_sub_go), .B(i_psram_sub_mem_addr
		[7]), .C(s00_axi_aresetn), .Z(i_psram_sub_AsyncPSRAMinst_n_489)
		);
	notech_nao3 i_psram_sub_AsyncPSRAMinst_i_340(.A(MEM_ADDR_OUT[7]), .B(s00_axi_aresetn
		), .C(i_psram_sub_go), .Z(i_psram_sub_AsyncPSRAMinst_n_488));
	notech_nand3 i_psram_sub_AsyncPSRAMinst_i_335(.A(i_psram_sub_go), .B(i_psram_sub_mem_addr
		[4]), .C(s00_axi_aresetn), .Z(i_psram_sub_AsyncPSRAMinst_n_487)
		);
	notech_nao3 i_psram_sub_AsyncPSRAMinst_i_334(.A(MEM_ADDR_OUT[4]), .B(s00_axi_aresetn
		), .C(i_psram_sub_go), .Z(i_psram_sub_AsyncPSRAMinst_n_486));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_27(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[22]), .Z(i_psram_sub_AsyncPSRAMinst_n_485
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_28(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[21]), .Z(i_psram_sub_AsyncPSRAMinst_n_483
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_291590(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[20]), .Z(i_psram_sub_AsyncPSRAMinst_n_482
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_31(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[19]), .Z(i_psram_sub_AsyncPSRAMinst_n_481
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_32(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[18]), .Z(i_psram_sub_AsyncPSRAMinst_n_480
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_33(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[17]), .Z(i_psram_sub_AsyncPSRAMinst_n_479
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_34(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[16]), .Z(i_psram_sub_AsyncPSRAMinst_n_478
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_35(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[15]), .Z(i_psram_sub_AsyncPSRAMinst_n_477
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_36(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[14]), .Z(i_psram_sub_AsyncPSRAMinst_n_476
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_37(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[13]), .Z(i_psram_sub_AsyncPSRAMinst_n_475
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_38(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[12]), .Z(i_psram_sub_AsyncPSRAMinst_n_474
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_39(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[11]), .Z(i_psram_sub_AsyncPSRAMinst_n_472
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_40(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[10]), .Z(i_psram_sub_AsyncPSRAMinst_n_471
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_41(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[9]), .Z(i_psram_sub_AsyncPSRAMinst_n_470
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_42(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[8]), .Z(i_psram_sub_AsyncPSRAMinst_n_469
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_43(.A(MEM_ADDR_OUT[7]), .B(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .C(s00_axi_aresetn), .Z(i_psram_sub_AsyncPSRAMinst_n_468));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_44(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[6]), .Z(i_psram_sub_AsyncPSRAMinst_n_467
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_45(.A(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .B(s00_axi_aresetn), .C(MEM_ADDR_OUT[5]), .Z(i_psram_sub_AsyncPSRAMinst_n_466
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_46(.A(MEM_ADDR_OUT[4]), .B(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .C(s00_axi_aresetn), .Z(i_psram_sub_AsyncPSRAMinst_n_465));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_143(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[4]), .B(i_psram_sub_AsyncPSRAMinst_cycle_time[3]), .C(i_psram_sub_AsyncPSRAMinst_cycle_time
		[5]), .D(i_psram_sub_AsyncPSRAMinst_n_515), .Z(i_psram_sub_AsyncPSRAMinst_n_464
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_129(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[2]), .B(i_psram_sub_AsyncPSRAMinst_n_2915), .Z(i_psram_sub_AsyncPSRAMinst_n_463
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_126(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[1]), .B(i_psram_sub_AsyncPSRAMinst_n_2914), .Z(i_psram_sub_AsyncPSRAMinst_n_462
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_127(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[0]), .B(i_psram_sub_AsyncPSRAMinst_n_2913), .Z(i_psram_sub_AsyncPSRAMinst_n_461
		));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_310(.A(i_psram_sub_AsyncPSRAMinst_n_292
		), .B(i_psram_sub_AsyncPSRAMinst_n_2967), .Z(i_psram_sub_AsyncPSRAMinst_n_454
		));
	notech_or4 i_psram_sub_AsyncPSRAMinst_i_146(.A(i_psram_sub_AsyncPSRAMinst_n_514
		), .B(i_psram_sub_AsyncPSRAMinst_n_543), .C(i_psram_sub_AsyncPSRAMinst_cycle_time
		[5]), .D(i_psram_sub_AsyncPSRAMinst_n_2917), .Z(i_psram_sub_AsyncPSRAMinst_n_453
		));
	notech_ao3 i_psram_sub_AsyncPSRAMinst_i_303(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[5]), .B(s00_axi_aresetn), .C(i_psram_sub_AsyncPSRAMinst_n_285),
		 .Z(i_psram_sub_AsyncPSRAMinst_n_452));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_302(.A(i_psram_sub_AsyncPSRAMinst_n_453
		), .B(i_psram_sub_AsyncPSRAMinst_n_2872), .C(s00_axi_aresetn), .D
		(i_psram_sub_AsyncPSRAMinst_n_2910), .Z(i_psram_sub_AsyncPSRAMinst_n_450
		));
	notech_nor2 i_psram_sub_AsyncPSRAMinst_i_304(.A(i_psram_sub_AsyncPSRAMinst_n_522
		), .B(i_psram_sub_AsyncPSRAMinst_n_2910), .Z(i_psram_sub_AsyncPSRAMinst_n_449
		));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_125(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[5]), .B(s00_axi_aresetn), .C(i_psram_sub_AsyncPSRAMinst_n_508),
		 .D(i_psram_sub_AsyncPSRAMinst_n_2918), .Z(i_psram_sub_AsyncPSRAMinst_n_448
		));
	notech_or4 i_psram_sub_AsyncPSRAMinst_i_149(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[4]), .B(i_psram_sub_AsyncPSRAMinst_n_514), .C(i_psram_sub_AsyncPSRAMinst_n_543
		), .D(i_psram_sub_AsyncPSRAMinst_n_444), .Z(i_psram_sub_AsyncPSRAMinst_n_447
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_295(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[4]), .B(i_psram_sub_AsyncPSRAMinst_n_2917), .Z(i_psram_sub_AsyncPSRAMinst_n_446
		));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_294(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[4]), .B(i_psram_sub_AsyncPSRAMinst_n_2909), .Z(i_psram_sub_AsyncPSRAMinst_n_445
		));
	notech_xor2 i_psram_sub_AsyncPSRAMinst_i_109(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[5]), .B(i_psram_sub_AsyncPSRAMinst_waitcount[5]), .Z(i_psram_sub_AsyncPSRAMinst_n_444
		));
	notech_ao3 i_psram_sub_AsyncPSRAMinst_i_153(.A(i_psram_sub_AsyncPSRAMinst_n_2866
		), .B(i_psram_sub_AsyncPSRAMinst_n_2916), .C(i_psram_sub_AsyncPSRAMinst_n_514
		), .Z(i_psram_sub_AsyncPSRAMinst_n_442));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_280(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[3]), .B(i_psram_sub_AsyncPSRAMinst_n_2916), .Z(i_psram_sub_AsyncPSRAMinst_n_441
		));
	notech_or4 i_psram_sub_AsyncPSRAMinst_i_158(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[2]), .B(i_psram_sub_AsyncPSRAMinst_n_568), .C(i_psram_sub_AsyncPSRAMinst_n_2914
		), .D(i_psram_sub_AsyncPSRAMinst_n_2913), .Z(i_psram_sub_AsyncPSRAMinst_n_440
		));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_159(.A(i_psram_sub_AsyncPSRAMinst_n_461
		), .B(i_psram_sub_AsyncPSRAMinst_cycle_time[2]), .C(i_psram_sub_AsyncPSRAMinst_n_2868
		), .D(i_psram_sub_AsyncPSRAMinst_n_2914), .Z(i_psram_sub_AsyncPSRAMinst_n_439
		));
	notech_or4 i_psram_sub_AsyncPSRAMinst_i_275(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[1]), .B(i_psram_sub_AsyncPSRAMinst_n_439), .C(i_psram_sub_AsyncPSRAMinst_n_2967
		), .D(i_psram_sub_AsyncPSRAMinst_n_2905), .Z(i_psram_sub_AsyncPSRAMinst_n_438
		));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_274(.A(i_psram_sub_AsyncPSRAMinst_n_440
		), .B(i_psram_sub_AsyncPSRAMinst_n_556), .C(i_psram_sub_AsyncPSRAMinst_waitcount
		[1]), .D(i_psram_sub_AsyncPSRAMinst_n_2905), .Z(i_psram_sub_AsyncPSRAMinst_n_437
		));
	notech_xor2 i_psram_sub_AsyncPSRAMinst_i_111(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[2]), .B(i_psram_sub_AsyncPSRAMinst_waitcount[2]), .Z(i_psram_sub_AsyncPSRAMinst_n_436
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_267(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[3]), .B(i_psram_sub_AsyncPSRAMinst_n_2907), .Z(i_psram_sub_AsyncPSRAMinst_n_433
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_269(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[1]), .B(i_psram_sub_AsyncPSRAMinst_n_2904), .Z(i_psram_sub_AsyncPSRAMinst_n_432
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_225(.A(i_psram_sub_AsyncPSRAMinst_last_page_read
		[17]), .B(i_psram_sub_AsyncPSRAMinst_n_2941), .Z(i_psram_sub_AsyncPSRAMinst_n_431
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_230(.A(i_psram_sub_mem_addr[19
		]), .B(i_psram_sub_AsyncPSRAMinst_n_2902), .Z(i_psram_sub_AsyncPSRAMinst_n_426
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_235(.A(i_psram_sub_AsyncPSRAMinst_last_page_read
		[12]), .B(i_psram_sub_AsyncPSRAMinst_n_2936), .Z(i_psram_sub_AsyncPSRAMinst_n_419
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_240(.A(i_psram_sub_mem_addr[14
		]), .B(i_psram_sub_AsyncPSRAMinst_n_2900), .Z(i_psram_sub_AsyncPSRAMinst_n_414
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_248(.A(i_psram_sub_AsyncPSRAMinst_last_page_read
		[7]), .B(i_psram_sub_AsyncPSRAMinst_n_2931), .Z(i_psram_sub_AsyncPSRAMinst_n_408
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_255(.A(i_psram_sub_mem_addr[9]
		), .B(i_psram_sub_AsyncPSRAMinst_n_2897), .Z(i_psram_sub_AsyncPSRAMinst_n_402
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_260(.A(i_psram_sub_AsyncPSRAMinst_last_page_read
		[2]), .B(i_psram_sub_AsyncPSRAMinst_n_2927), .Z(i_psram_sub_AsyncPSRAMinst_n_396
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_265(.A(i_psram_sub_mem_addr[4]
		), .B(i_psram_sub_AsyncPSRAMinst_n_2895), .Z(i_psram_sub_AsyncPSRAMinst_n_387
		));
	notech_xor2 i_psram_sub_AsyncPSRAMinst_i_176(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[0]), .B(i_psram_sub_AsyncPSRAMinst_waitcount[0]), .Z(i_psram_sub_AsyncPSRAMinst_n_386
		));
	notech_xor2 i_psram_sub_AsyncPSRAMinst_i_175(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[1]), .B(i_psram_sub_AsyncPSRAMinst_waitcount[1]), .Z(i_psram_sub_AsyncPSRAMinst_n_384
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_195(.A(i_psram_sub_AsyncPSRAMinst_state
		[0]), .B(i_psram_sub_AsyncPSRAMinst_n_2920), .C(i_psram_sub_AsyncPSRAMinst_n_2873
		), .Z(i_psram_sub_AsyncPSRAMinst_n_383));
	notech_ao3 i_psram_sub_AsyncPSRAMinst_i_194(.A(i_psram_sub_AsyncPSRAMinst_n_2919
		), .B(i_psram_sub_AsyncPSRAMinst_n_245), .C(i_psram_sub_AsyncPSRAMinst_state
		[1]), .Z(i_psram_sub_AsyncPSRAMinst_n_382));
	notech_ao3 i_psram_sub_AsyncPSRAMinst_i_60(.A(i_psram_sub_AsyncPSRAMinst_n_115
		), .B(i_psram_sub_AsyncPSRAMinst_n_658), .C(i_psram_sub_AsyncPSRAMinst_cen_old
		), .Z(i_psram_sub_AsyncPSRAMinst_n_381));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_71(.A(i_psram_sub_AsyncPSRAMinst_cen_old
		), .B(i_psram_sub_AsyncPSRAMinst_n_658), .Z(i_psram_sub_AsyncPSRAMinst_n_379
		));
	notech_ao3 i_psram_sub_AsyncPSRAMinst_i_66(.A(i_psram_sub_AsyncPSRAMinst_n_109
		), .B(i_psram_sub_AsyncPSRAMinst_n_658), .C(i_psram_sub_AsyncPSRAMinst_cen_old
		), .Z(i_psram_sub_AsyncPSRAMinst_n_378));
	notech_ao3 i_psram_sub_AsyncPSRAMinst_i_67(.A(i_psram_sub_AsyncPSRAMinst_n_108
		), .B(i_psram_sub_AsyncPSRAMinst_n_658), .C(i_psram_sub_AsyncPSRAMinst_cen_old
		), .Z(i_psram_sub_AsyncPSRAMinst_n_377));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_177(.A(i_psram_sub_AsyncPSRAMinst_n_463
		), .B(i_psram_sub_AsyncPSRAMinst_n_441), .C(i_psram_sub_AsyncPSRAMinst_n_462
		), .D(i_psram_sub_AsyncPSRAMinst_n_2913), .Z(i_psram_sub_AsyncPSRAMinst_n_231
		));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_178(.A(i_psram_sub_go), .B(i_psram_sub_AsyncPSRAMinst_cem_time_expired
		), .C(i_psram_sub_AsyncPSRAMinst_n_2919), .D(i_psram_sub_AsyncPSRAMinst_n_2920
		), .Z(i_psram_sub_AsyncPSRAMinst_n_232));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_167(.A(i_psram_sub_AsyncPSRAMinst_n_532
		), .B(i_psram_sub_AsyncPSRAMinst_n_356), .C(i_psram_sub_AsyncPSRAMinst_n_588
		), .Z(i_psram_sub_AsyncPSRAMinst_n_233));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_184(.A(i_psram_sub_mem_byte_en
		[0]), .B(i_psram_sub_AsyncPSRAMinst_n_2920), .Z(i_psram_sub_AsyncPSRAMinst_n_235
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_185(.A(i_psram_sub_mem_byte_en
		[1]), .B(i_psram_sub_AsyncPSRAMinst_n_2920), .Z(i_psram_sub_AsyncPSRAMinst_n_236
		));
	notech_or4 i_psram_sub_AsyncPSRAMinst_i_186(.A(i_psram_sub_AsyncPSRAMinst_n_642
		), .B(i_psram_sub_AsyncPSRAMinst_state[1]), .C(i_psram_sub_AsyncPSRAMinst_n_2873
		), .D(i_psram_sub_AsyncPSRAMinst_n_2919), .Z(i_psram_sub_AsyncPSRAMinst_n_237
		));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_187(.A(i_psram_sub_AsyncPSRAMinst_state
		[1]), .B(i_psram_sub_AsyncPSRAMinst_n_642), .Z(i_psram_sub_AsyncPSRAMinst_n_238
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_188(.A(i_psram_sub_AsyncPSRAMinst_n_107
		), .B(i_psram_sub_AsyncPSRAMinst_n_2921), .Z(i_psram_sub_AsyncPSRAMinst_n_239
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_189(.A(i_psram_sub_AsyncPSRAMinst_n_110
		), .B(i_psram_sub_AsyncPSRAMinst_n_2921), .Z(i_psram_sub_AsyncPSRAMinst_n_240
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_190(.A(i_psram_sub_AsyncPSRAMinst_n_111
		), .B(i_psram_sub_AsyncPSRAMinst_n_2921), .Z(i_psram_sub_AsyncPSRAMinst_n_241
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_191(.A(i_psram_sub_AsyncPSRAMinst_n_112
		), .B(i_psram_sub_AsyncPSRAMinst_n_2921), .Z(i_psram_sub_AsyncPSRAMinst_n_242
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_192(.A(i_psram_sub_AsyncPSRAMinst_n_113
		), .B(i_psram_sub_AsyncPSRAMinst_n_2921), .Z(i_psram_sub_AsyncPSRAMinst_n_243
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_193(.A(i_psram_sub_AsyncPSRAMinst_n_114
		), .B(i_psram_sub_AsyncPSRAMinst_n_2921), .Z(i_psram_sub_AsyncPSRAMinst_n_244
		));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_163(.A(i_psram_sub_AsyncPSRAMinst_cem_time_expired
		), .B(i_psram_sub_AsyncPSRAMinst_n_246), .Z(i_psram_sub_AsyncPSRAMinst_n_245
		));
	notech_nor2 i_psram_sub_AsyncPSRAMinst_i_196(.A(i_psram_sub_go), .B(i_psram_sub_AsyncPSRAMinst_n_2968
		), .Z(i_psram_sub_AsyncPSRAMinst_n_246));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_197(.A(i_psram_sub_go), .B(i_psram_sub_AsyncPSRAMinst_n_2919
		), .C(i_psram_sub_AsyncPSRAMinst_n_2920), .D(i_psram_sub_AsyncPSRAMinst_n_248
		), .Z(i_psram_sub_AsyncPSRAMinst_n_247));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_171(.A(i_psram_sub_command), .B
		(i_psram_sub_AsyncPSRAMinst_n_637), .Z(i_psram_sub_AsyncPSRAMinst_n_248
		));
	notech_nand3 i_psram_sub_AsyncPSRAMinst_i_219(.A(i_psram_sub_go), .B(i_psram_sub_command
		), .C(i_psram_sub_AsyncPSRAMinst_n_254), .Z(i_psram_sub_AsyncPSRAMinst_n_253
		));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_162(.A(i_psram_sub_AsyncPSRAMinst_cem_time_expired
		), .B(i_psram_sub_AsyncPSRAMinst_n_2863), .Z(i_psram_sub_AsyncPSRAMinst_n_254
		));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_266(.A(i_psram_sub_AsyncPSRAMinst_n_588
		), .B(i_psram_sub_AsyncPSRAMinst_n_518), .Z(i_psram_sub_AsyncPSRAMinst_n_255
		));
	notech_ao3 i_psram_sub_AsyncPSRAMinst_i_270(.A(i_psram_sub_AsyncPSRAMinst_n_257
		), .B(i_psram_sub_AsyncPSRAMinst_waitcount[1]), .C(i_psram_sub_AsyncPSRAMinst_n_518
		), .Z(i_psram_sub_AsyncPSRAMinst_n_256));
	notech_or4 i_psram_sub_AsyncPSRAMinst_i_160(.A(i_psram_sub_AsyncPSRAMinst_n_436
		), .B(i_psram_sub_AsyncPSRAMinst_n_568), .C(i_psram_sub_AsyncPSRAMinst_n_2914
		), .D(i_psram_sub_AsyncPSRAMinst_cycle_time[0]), .Z(i_psram_sub_AsyncPSRAMinst_n_257
		));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_271(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[0]), .B(s00_axi_aresetn), .C(i_psram_sub_AsyncPSRAMinst_n_259),
		 .D(i_psram_sub_AsyncPSRAMinst_n_2904), .Z(i_psram_sub_AsyncPSRAMinst_n_258
		));
	notech_or4 i_psram_sub_AsyncPSRAMinst_i_161(.A(i_psram_sub_AsyncPSRAMinst_n_436
		), .B(i_psram_sub_AsyncPSRAMinst_n_568), .C(i_psram_sub_AsyncPSRAMinst_n_2913
		), .D(i_psram_sub_AsyncPSRAMinst_cycle_time[1]), .Z(i_psram_sub_AsyncPSRAMinst_n_259
		));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_276(.A(i_psram_sub_AsyncPSRAMinst_n_263
		), .B(i_psram_sub_AsyncPSRAMinst_n_518), .Z(i_psram_sub_AsyncPSRAMinst_n_262
		));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_156(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[1]), .B(i_psram_sub_AsyncPSRAMinst_n_505), .C(i_psram_sub_AsyncPSRAMinst_n_2905
		), .D(i_psram_sub_AsyncPSRAMinst_n_265), .Z(i_psram_sub_AsyncPSRAMinst_n_263
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_157(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[2]), .B(i_psram_sub_AsyncPSRAMinst_n_2913), .C(i_psram_sub_AsyncPSRAMinst_n_2868
		), .Z(i_psram_sub_AsyncPSRAMinst_n_265));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_151(.A(i_psram_sub_AsyncPSRAMinst_n_273
		), .B(i_psram_sub_AsyncPSRAMinst_n_518), .C(i_psram_sub_AsyncPSRAMinst_n_2967
		), .D(i_psram_sub_AsyncPSRAMinst_n_271), .Z(i_psram_sub_AsyncPSRAMinst_n_269
		));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_152(.A(i_psram_sub_AsyncPSRAMinst_n_526
		), .B(i_psram_sub_AsyncPSRAMinst_n_2870), .Z(i_psram_sub_AsyncPSRAMinst_n_271
		));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_155(.A(i_psram_sub_AsyncPSRAMinst_n_463
		), .B(i_psram_sub_AsyncPSRAMinst_n_462), .C(i_psram_sub_AsyncPSRAMinst_n_2866
		), .D(i_psram_sub_AsyncPSRAMinst_n_562), .Z(i_psram_sub_AsyncPSRAMinst_n_273
		));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_293(.A(i_psram_sub_AsyncPSRAMinst_n_2905
		), .B(i_psram_sub_AsyncPSRAMinst_n_2904), .C(i_psram_sub_AsyncPSRAMinst_n_2916
		), .D(i_psram_sub_AsyncPSRAMinst_n_559), .Z(i_psram_sub_AsyncPSRAMinst_n_274
		));
	notech_ao4 i_psram_sub_AsyncPSRAMinst_i_147(.A(i_psram_sub_AsyncPSRAMinst_n_518
		), .B(i_psram_sub_AsyncPSRAMinst_n_231), .C(i_psram_sub_AsyncPSRAMinst_n_280
		), .D(i_psram_sub_AsyncPSRAMinst_n_2967), .Z(i_psram_sub_AsyncPSRAMinst_n_278
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_148(.A(i_psram_sub_AsyncPSRAMinst_n_526
		), .B(i_psram_sub_AsyncPSRAMinst_n_530), .C(i_psram_sub_AsyncPSRAMinst_n_281
		), .Z(i_psram_sub_AsyncPSRAMinst_n_280));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_299(.A(i_psram_sub_AsyncPSRAMinst_n_507
		), .B(i_psram_sub_AsyncPSRAMinst_n_282), .Z(i_psram_sub_AsyncPSRAMinst_n_281
		));
	notech_ao3 i_psram_sub_AsyncPSRAMinst_i_150(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[4]), .B(i_psram_sub_AsyncPSRAMinst_n_542), .C(i_psram_sub_AsyncPSRAMinst_n_444
		), .Z(i_psram_sub_AsyncPSRAMinst_n_282));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_145(.A(i_psram_sub_AsyncPSRAMinst_n_526
		), .B(i_psram_sub_AsyncPSRAMinst_n_530), .C(i_psram_sub_AsyncPSRAMinst_n_533
		), .D(i_psram_sub_AsyncPSRAMinst_n_286), .Z(i_psram_sub_AsyncPSRAMinst_n_285
		));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_305(.A(i_psram_sub_AsyncPSRAMinst_n_508
		), .B(i_psram_sub_AsyncPSRAMinst_n_2864), .Z(i_psram_sub_AsyncPSRAMinst_n_286
		));
	notech_ao3 i_psram_sub_AsyncPSRAMinst_i_141(.A(i_psram_sub_AsyncPSRAMinst_n_522
		), .B(i_psram_sub_AsyncPSRAMinst_n_454), .C(i_psram_sub_AsyncPSRAMinst_n_448
		), .Z(i_psram_sub_AsyncPSRAMinst_n_291));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_142(.A(i_psram_sub_AsyncPSRAMinst_n_526
		), .B(i_psram_sub_AsyncPSRAMinst_n_530), .C(i_psram_sub_AsyncPSRAMinst_n_533
		), .D(i_psram_sub_AsyncPSRAMinst_n_538), .Z(i_psram_sub_AsyncPSRAMinst_n_292
		));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_144(.A(i_psram_sub_AsyncPSRAMinst_cycle_time
		[6]), .B(i_psram_sub_AsyncPSRAMinst_n_446), .C(i_psram_sub_AsyncPSRAMinst_n_532
		), .D(i_psram_sub_AsyncPSRAMinst_n_2918), .Z(i_psram_sub_AsyncPSRAMinst_n_293
		));
	notech_ao3 i_psram_sub_AsyncPSRAMinst_i_170(.A(i_psram_sub_AsyncPSRAMinst_n_461
		), .B(i_psram_sub_AsyncPSRAMinst_n_521), .C(i_psram_sub_AsyncPSRAMinst_cycle_time
		[4]), .Z(i_psram_sub_AsyncPSRAMinst_n_294));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_172(.A(i_psram_sub_AsyncPSRAMinst_n_463
		), .B(i_psram_sub_AsyncPSRAMinst_n_461), .C(i_psram_sub_AsyncPSRAMinst_n_462
		), .D(i_psram_sub_AsyncPSRAMinst_n_2916), .Z(i_psram_sub_AsyncPSRAMinst_n_295
		));
	notech_ao3 i_psram_sub_AsyncPSRAMinst_i_173(.A(i_psram_sub_AsyncPSRAMinst_n_461
		), .B(i_psram_sub_AsyncPSRAMinst_n_463), .C(i_psram_sub_AsyncPSRAMinst_cycle_time
		[1]), .Z(i_psram_sub_AsyncPSRAMinst_n_297));
	notech_ao3 i_psram_sub_AsyncPSRAMinst_i_174(.A(i_psram_sub_AsyncPSRAMinst_n_462
		), .B(i_psram_sub_AsyncPSRAMinst_n_461), .C(i_psram_sub_AsyncPSRAMinst_cycle_time
		[2]), .Z(i_psram_sub_AsyncPSRAMinst_n_299));
	notech_and4 i_psram_sub_AsyncPSRAMinst_i_393(.A(i_psram_sub_AsyncPSRAMinst_page_valid
		), .B(i_psram_sub_AsyncPSRAMinst_n_491), .C(s00_axi_aresetn), .D
		(i_psram_sub_AsyncPSRAMinst_n_2919), .Z(i_psram_sub_AsyncPSRAMinst_n_348
		));
	notech_and3 i_psram_sub_AsyncPSRAMinst_i_396(.A(i_psram_sub_AsyncPSRAMinst_state
		[0]), .B(s00_axi_aresetn), .C(i_psram_sub_AsyncPSRAMinst_current_cmd
		), .Z(i_psram_sub_AsyncPSRAMinst_n_349));
	notech_nor2 i_psram_sub_AsyncPSRAMinst_i_397(.A(i_psram_sub_go), .B(i_psram_sub_AsyncPSRAMinst_state
		[1]), .Z(i_psram_sub_AsyncPSRAMinst_n_351));
	notech_nand2 i_psram_sub_AsyncPSRAMinst_i_398(.A(i_psram_sub_command), .B
		(i_psram_sub_AsyncPSRAMinst_n_2920), .Z(i_psram_sub_AsyncPSRAMinst_n_352
		));
	notech_or2 i_psram_sub_AsyncPSRAMinst_i_183(.A(i_psram_sub_AsyncPSRAMinst_waitcount
		[0]), .B(i_psram_sub_AsyncPSRAMinst_n_2913), .Z(i_psram_sub_AsyncPSRAMinst_n_356
		));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_94(.A(MEM_DATA_I[0]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_357));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_92(.A(MEM_DATA_I[1]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_358));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_91(.A(MEM_DATA_I[2]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_359));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_90(.A(MEM_DATA_I[3]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_361));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_89(.A(MEM_DATA_I[4]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_362));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_88(.A(MEM_DATA_I[5]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_363));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_87(.A(MEM_DATA_I[6]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_364));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_86(.A(MEM_DATA_I[7]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_366));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_85(.A(MEM_DATA_I[8]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_367));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_84(.A(MEM_DATA_I[9]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_368));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_83(.A(MEM_DATA_I[10]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_369));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_82(.A(MEM_DATA_I[11]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_371));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_81(.A(MEM_DATA_I[12]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_372));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_79(.A(MEM_DATA_I[13]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_373));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_76(.A(MEM_DATA_I[14]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_374));
	notech_and2 i_psram_sub_AsyncPSRAMinst_i_75(.A(MEM_DATA_I[15]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_AsyncPSRAMinst_n_376));
	notech_inv i_02655(.A(i_psram_sub_mem_addr[0]), .Z(i_psram_sub_function_plus_2
		[0]));
	notech_nand2 i_12654(.A(i_psram_sub_mem_addr[0]), .B(i_psram_sub_mem_addr
		[1]), .Z(n_1391736));
	notech_nand2 i_22653(.A(i_psram_sub_mem_addr[1]), .B(i_psram_sub_mem_addr
		[2]), .Z(n_1401735));
	notech_nand2 i_32652(.A(i_psram_sub_mem_addr[2]), .B(i_psram_sub_mem_addr
		[3]), .Z(n_1411734));
	notech_nand2 i_42651(.A(i_psram_sub_mem_addr[3]), .B(i_psram_sub_mem_addr
		[4]), .Z(n_1421733));
	notech_nand2 i_52650(.A(i_psram_sub_mem_addr[4]), .B(i_psram_sub_mem_addr
		[5]), .Z(n_1431732));
	notech_nand2 i_62649(.A(i_psram_sub_mem_addr[5]), .B(i_psram_sub_mem_addr
		[6]), .Z(n_1441731));
	notech_nand2 i_72648(.A(i_psram_sub_mem_addr[6]), .B(i_psram_sub_mem_addr
		[7]), .Z(n_1451730));
	notech_nand2 i_82647(.A(i_psram_sub_mem_addr[7]), .B(i_psram_sub_mem_addr
		[8]), .Z(n_1461729));
	notech_nand2 i_92646(.A(i_psram_sub_mem_addr[8]), .B(i_psram_sub_mem_addr
		[9]), .Z(n_1471728));
	notech_nand2 i_102645(.A(i_psram_sub_mem_addr[9]), .B(i_psram_sub_mem_addr
		[10]), .Z(n_1481727));
	notech_nand2 i_112644(.A(i_psram_sub_mem_addr[10]), .B(i_psram_sub_mem_addr
		[11]), .Z(n_1491726));
	notech_nand2 i_122643(.A(i_psram_sub_mem_addr[11]), .B(i_psram_sub_mem_addr
		[12]), .Z(n_1501725));
	notech_nand2 i_132642(.A(i_psram_sub_mem_addr[12]), .B(i_psram_sub_mem_addr
		[13]), .Z(n_1511724));
	notech_nand2 i_142641(.A(i_psram_sub_mem_addr[13]), .B(i_psram_sub_mem_addr
		[14]), .Z(n_1521723));
	notech_nand2 i_152640(.A(i_psram_sub_mem_addr[14]), .B(i_psram_sub_mem_addr
		[15]), .Z(n_153));
	notech_nand2 i_162639(.A(i_psram_sub_mem_addr[15]), .B(i_psram_sub_mem_addr
		[16]), .Z(n_1541722));
	notech_nand2 i_172638(.A(i_psram_sub_mem_addr[16]), .B(i_psram_sub_mem_addr
		[17]), .Z(n_155));
	notech_nand2 i_182637(.A(i_psram_sub_mem_addr[17]), .B(i_psram_sub_mem_addr
		[18]), .Z(n_1561721));
	notech_nand2 i_192636(.A(i_psram_sub_mem_addr[18]), .B(i_psram_sub_mem_addr
		[19]), .Z(n_1571720));
	notech_nand2 i_202635(.A(i_psram_sub_mem_addr[19]), .B(i_psram_sub_mem_addr
		[20]), .Z(n_1581719));
	notech_nand2 i_21(.A(i_psram_sub_mem_addr[20]), .B(i_psram_sub_mem_addr[
		21]), .Z(n_1591718));
	notech_inv i_232634(.A(i_psram_sub_function_plus_2[0]), .Z(n_1611717));
	notech_inv i_242633(.A(n_1391736), .Z(n_2771716));
	notech_nor2 i_252632(.A(i_psram_sub_function_plus_2[0]), .B(n_1401735), 
		.Z(n_1631715));
	notech_nor2 i_262631(.A(n_1391736), .B(n_1411734), .Z(n_1641714));
	notech_nor2 i_272630(.A(n_1401735), .B(n_1421733), .Z(n_1651713));
	notech_nor2 i_282629(.A(n_1411734), .B(n_1431732), .Z(n_1661712));
	notech_nor2 i_292628(.A(n_1421733), .B(n_1441731), .Z(n_1671711));
	notech_nor2 i_302627(.A(n_1431732), .B(n_1451730), .Z(n_1681710));
	notech_nor2 i_312626(.A(n_1441731), .B(n_1461729), .Z(n_1691709));
	notech_nor2 i_322625(.A(n_1451730), .B(n_1471728), .Z(n_1701708));
	notech_nor2 i_332624(.A(n_1461729), .B(n_1481727), .Z(n_1711707));
	notech_nor2 i_342623(.A(n_1471728), .B(n_1491726), .Z(n_1721706));
	notech_nor2 i_352622(.A(n_1481727), .B(n_1501725), .Z(n_1731705));
	notech_nor2 i_362621(.A(n_1491726), .B(n_1511724), .Z(n_1741704));
	notech_nor2 i_372620(.A(n_1501725), .B(n_1521723), .Z(n_175));
	notech_nor2 i_382619(.A(n_1511724), .B(n_153), .Z(n_1761703));
	notech_nor2 i_392618(.A(n_1521723), .B(n_1541722), .Z(n_1771702));
	notech_nor2 i_402617(.A(n_153), .B(n_155), .Z(n_1781701));
	notech_nor2 i_412616(.A(n_1541722), .B(n_1561721), .Z(n_179));
	notech_nor2 i_422615(.A(n_155), .B(n_1571720), .Z(n_1801700));
	notech_nor2 i_43(.A(n_1561721), .B(n_1581719), .Z(n_1811699));
	notech_nor2 i_442614(.A(n_1571720), .B(n_1591718), .Z(n_1821698));
	notech_inv i_462613(.A(n_1611717), .Z(n_1841697));
	notech_inv i_472612(.A(n_2771716), .Z(n_1851696));
	notech_inv i_482611(.A(n_1631715), .Z(n_1861695));
	notech_inv i_492610(.A(n_1641714), .Z(n_2781694));
	notech_nand2 i_502609(.A(n_1611717), .B(n_1651713), .Z(n_1881693));
	notech_nand2 i_512608(.A(n_2771716), .B(n_1661712), .Z(n_1891692));
	notech_nand2 i_522607(.A(n_1631715), .B(n_1671711), .Z(n_1901691));
	notech_nand2 i_532606(.A(n_1641714), .B(n_1681710), .Z(n_1911690));
	notech_nand2 i_542605(.A(n_1651713), .B(n_1691709), .Z(n_1921689));
	notech_nand2 i_552604(.A(n_1661712), .B(n_1701708), .Z(n_1931688));
	notech_nand2 i_562603(.A(n_1671711), .B(n_1711707), .Z(n_1941687));
	notech_nand2 i_572602(.A(n_1681710), .B(n_1721706), .Z(n_1951686));
	notech_nand2 i_582601(.A(n_1691709), .B(n_1731705), .Z(n_1961685));
	notech_nand2 i_592600(.A(n_1701708), .B(n_1741704), .Z(n_197));
	notech_nand2 i_602599(.A(n_1711707), .B(n_175), .Z(n_1981684));
	notech_nand2 i_612598(.A(n_1721706), .B(n_1761703), .Z(n_1991683));
	notech_nand2 i_622597(.A(n_1731705), .B(n_1771702), .Z(n_2001682));
	notech_nand2 i_632596(.A(n_1741704), .B(n_1781701), .Z(n_2011681));
	notech_nand2 i_642595(.A(n_175), .B(n_179), .Z(n_2021680));
	notech_nand2 i_652594(.A(n_1761703), .B(n_1801700), .Z(n_203));
	notech_nand2 i_662593(.A(n_1771702), .B(n_1811699), .Z(n_204));
	notech_nand2 i_672592(.A(n_1781701), .B(n_1821698), .Z(n_205));
	notech_inv i_692591(.A(n_1841697), .Z(n_2071679));
	notech_inv i_702590(.A(n_1851696), .Z(n_2081678));
	notech_inv i_71(.A(n_1861695), .Z(n_2091677));
	notech_inv i_722589(.A(n_2781694), .Z(n_2101676));
	notech_inv i_73(.A(n_1881693), .Z(n_2111675));
	notech_inv i_742588(.A(n_1891692), .Z(n_2121674));
	notech_nor2 i_772587(.A(n_1841697), .B(n_1921689), .Z(n_2151673));
	notech_nor2 i_782586(.A(n_1851696), .B(n_1931688), .Z(n_2161672));
	notech_nor2 i_792585(.A(n_1861695), .B(n_1941687), .Z(n_2171671));
	notech_nor2 i_802584(.A(n_2781694), .B(n_1951686), .Z(n_2181670));
	notech_nor2 i_812583(.A(n_1881693), .B(n_1961685), .Z(n_2191669));
	notech_nor2 i_822582(.A(n_1891692), .B(n_197), .Z(n_2201668));
	notech_nor2 i_832581(.A(n_1901691), .B(n_1981684), .Z(n_2211667));
	notech_nor2 i_842580(.A(n_1911690), .B(n_1991683), .Z(n_2221666));
	notech_nor2 i_852579(.A(n_1921689), .B(n_2001682), .Z(n_2231665));
	notech_nor2 i_862578(.A(n_1931688), .B(n_2011681), .Z(n_2241664));
	notech_nor2 i_872577(.A(n_1941687), .B(n_2021680), .Z(n_2251663));
	notech_nor2 i_882576(.A(n_1951686), .B(n_203), .Z(n_226));
	notech_nor2 i_892575(.A(n_1961685), .B(n_204), .Z(n_227));
	notech_nor2 i_902574(.A(n_197), .B(n_205), .Z(n_2281662));
	notech_inv i_922573(.A(n_2071679), .Z(n_2301661));
	notech_inv i_93(.A(n_2081678), .Z(n_2311660));
	notech_inv i_94(.A(n_2091677), .Z(n_2321659));
	notech_inv i_95(.A(n_2101676), .Z(n_2331658));
	notech_inv i_962572(.A(n_2111675), .Z(n_2341657));
	notech_inv i_972571(.A(n_2121674), .Z(n_235));
	notech_inv i_1002570(.A(n_2151673), .Z(n_2381656));
	notech_inv i_1012569(.A(n_2161672), .Z(n_2391655));
	notech_inv i_1022568(.A(n_2171671), .Z(n_2401654));
	notech_inv i_1032567(.A(n_2181670), .Z(n_241));
	notech_inv i_1042566(.A(n_2191669), .Z(n_2421653));
	notech_inv i_1052565(.A(n_2201668), .Z(n_2431652));
	notech_inv i_1062564(.A(n_2211667), .Z(n_2441651));
	notech_inv i_1072563(.A(n_2221666), .Z(n_2821650));
	notech_nand2 i_1082562(.A(n_2071679), .B(n_2231665), .Z(n_2461649));
	notech_nand2 i_109(.A(n_2081678), .B(n_2241664), .Z(n_2471648));
	notech_nand2 i_110(.A(n_2091677), .B(n_2251663), .Z(n_2481647));
	notech_nand2 i_111(.A(n_2101676), .B(n_226), .Z(n_2491646));
	notech_nand2 i_112(.A(n_2111675), .B(n_227), .Z(n_250));
	notech_nand2 i_113(.A(n_2121674), .B(n_2281662), .Z(n_251));
	notech_inv i_1382561(.A(n_2301661), .Z(n_2861645));
	notech_inv i_1392560(.A(i_psram_sub_mem_addr[1]), .Z(n_2891644));
	notech_nand2 i_1402559(.A(n_2891644), .B(n_2301661), .Z(n_2901643));
	notech_nand2 i_1412558(.A(i_psram_sub_mem_addr[1]), .B(n_2861645), .Z(n_2871642
		));
	notech_nand2 i_1422557(.A(n_2871642), .B(n_2901643), .Z(n_2881641));
	notech_inv i_1432556(.A(n_2881641), .Z(i_psram_sub_function_plus_2[1])
		);
	notech_inv i_1442555(.A(n_2311660), .Z(n_2911640));
	notech_inv i_1452554(.A(i_psram_sub_mem_addr[2]), .Z(n_2941639));
	notech_nand2 i_1462553(.A(n_2941639), .B(n_2311660), .Z(n_2951638));
	notech_nand2 i_1472552(.A(i_psram_sub_mem_addr[2]), .B(n_2911640), .Z(n_2921637
		));
	notech_nand2 i_1482551(.A(n_2921637), .B(n_2951638), .Z(n_2931636));
	notech_inv i_1492550(.A(n_2931636), .Z(i_psram_sub_function_plus_2[2])
		);
	notech_inv i_1502549(.A(n_2321659), .Z(n_2961635));
	notech_inv i_1512548(.A(i_psram_sub_mem_addr[3]), .Z(n_2991634));
	notech_nand2 i_1522547(.A(n_2991634), .B(n_2321659), .Z(n_3001633));
	notech_nand2 i_1532546(.A(i_psram_sub_mem_addr[3]), .B(n_2961635), .Z(n_2971632
		));
	notech_nand2 i_1542545(.A(n_2971632), .B(n_3001633), .Z(n_2981631));
	notech_inv i_1552544(.A(n_2981631), .Z(i_psram_sub_function_plus_2[3])
		);
	notech_inv i_1562543(.A(n_2331658), .Z(n_3011630));
	notech_inv i_1572542(.A(i_psram_sub_mem_addr[4]), .Z(n_3041629));
	notech_nand2 i_1582541(.A(n_3041629), .B(n_2331658), .Z(n_3051628));
	notech_nand2 i_1592540(.A(i_psram_sub_mem_addr[4]), .B(n_3011630), .Z(n_3021627
		));
	notech_nand2 i_1602539(.A(n_3021627), .B(n_3051628), .Z(n_3031626));
	notech_inv i_1612538(.A(n_3031626), .Z(i_psram_sub_function_plus_2[4])
		);
	notech_inv i_1622537(.A(n_2341657), .Z(n_3061625));
	notech_inv i_1632536(.A(i_psram_sub_mem_addr[5]), .Z(n_3091624));
	notech_nand2 i_1642535(.A(n_3091624), .B(n_2341657), .Z(n_3101623));
	notech_nand2 i_1652534(.A(i_psram_sub_mem_addr[5]), .B(n_3061625), .Z(n_3071622
		));
	notech_nand2 i_1662533(.A(n_3071622), .B(n_3101623), .Z(n_3081621));
	notech_inv i_1672532(.A(n_3081621), .Z(i_psram_sub_function_plus_2[5])
		);
	notech_inv i_1682531(.A(n_235), .Z(n_3111620));
	notech_inv i_1692530(.A(i_psram_sub_mem_addr[6]), .Z(n_3141619));
	notech_nand2 i_1702529(.A(n_3141619), .B(n_235), .Z(n_3151618));
	notech_nand2 i_1712528(.A(i_psram_sub_mem_addr[6]), .B(n_3111620), .Z(n_3121617
		));
	notech_nand2 i_1722527(.A(n_3121617), .B(n_3151618), .Z(n_3131616));
	notech_inv i_1732526(.A(n_3131616), .Z(i_psram_sub_function_plus_2[6])
		);
	notech_inv i_1742525(.A(n_1901691), .Z(n_3161615));
	notech_inv i_1752524(.A(i_psram_sub_mem_addr[7]), .Z(n_3191614));
	notech_nand2 i_1762523(.A(n_3191614), .B(n_1901691), .Z(n_3201613));
	notech_nand2 i_1772522(.A(i_psram_sub_mem_addr[7]), .B(n_3161615), .Z(n_3171612
		));
	notech_nand2 i_1782521(.A(n_3171612), .B(n_3201613), .Z(n_3181611));
	notech_inv i_1792520(.A(n_3181611), .Z(i_psram_sub_function_plus_2[7])
		);
	notech_inv i_1802519(.A(n_1911690), .Z(n_3211610));
	notech_inv i_1812518(.A(i_psram_sub_mem_addr[8]), .Z(n_3241609));
	notech_nand2 i_1822517(.A(n_3241609), .B(n_1911690), .Z(n_3251608));
	notech_nand2 i_1832516(.A(i_psram_sub_mem_addr[8]), .B(n_3211610), .Z(n_3221607
		));
	notech_nand2 i_1842515(.A(n_3221607), .B(n_3251608), .Z(n_3231606));
	notech_inv i_1852514(.A(n_3231606), .Z(i_psram_sub_function_plus_2[8])
		);
	notech_inv i_1862513(.A(n_2381656), .Z(n_3261605));
	notech_inv i_1872512(.A(i_psram_sub_mem_addr[9]), .Z(n_3291604));
	notech_nand2 i_1882511(.A(n_3291604), .B(n_2381656), .Z(n_3301603));
	notech_nand2 i_1892510(.A(i_psram_sub_mem_addr[9]), .B(n_3261605), .Z(n_3271602
		));
	notech_nand2 i_1902509(.A(n_3271602), .B(n_3301603), .Z(n_3281601));
	notech_inv i_1912508(.A(n_3281601), .Z(i_psram_sub_function_plus_2[9])
		);
	notech_inv i_1922507(.A(n_2391655), .Z(n_3311600));
	notech_inv i_1932506(.A(i_psram_sub_mem_addr[10]), .Z(n_3341599));
	notech_nand2 i_1942505(.A(n_3341599), .B(n_2391655), .Z(n_3351598));
	notech_nand2 i_1952504(.A(i_psram_sub_mem_addr[10]), .B(n_3311600), .Z(n_3321597
		));
	notech_nand2 i_1962503(.A(n_3321597), .B(n_3351598), .Z(n_3331596));
	notech_inv i_1972502(.A(n_3331596), .Z(i_psram_sub_function_plus_2[10])
		);
	notech_inv i_1982501(.A(n_2401654), .Z(n_3361595));
	notech_inv i_1992500(.A(i_psram_sub_mem_addr[11]), .Z(n_3391594));
	notech_nand2 i_2002499(.A(n_3391594), .B(n_2401654), .Z(n_3401593));
	notech_nand2 i_2012498(.A(i_psram_sub_mem_addr[11]), .B(n_3361595), .Z(n_3371592
		));
	notech_nand2 i_2022497(.A(n_3371592), .B(n_3401593), .Z(n_3381591));
	notech_inv i_2032496(.A(n_3381591), .Z(i_psram_sub_function_plus_2[11])
		);
	notech_inv i_2042495(.A(n_241), .Z(n_3411590));
	notech_inv i_2052494(.A(i_psram_sub_mem_addr[12]), .Z(n_3441589));
	notech_nand2 i_2062493(.A(n_3441589), .B(n_241), .Z(n_3451588));
	notech_nand2 i_2072492(.A(i_psram_sub_mem_addr[12]), .B(n_3411590), .Z(n_3421587
		));
	notech_nand2 i_2082491(.A(n_3421587), .B(n_3451588), .Z(n_3431586));
	notech_inv i_2092490(.A(n_3431586), .Z(i_psram_sub_function_plus_2[12])
		);
	notech_inv i_2102489(.A(n_2421653), .Z(n_3461585));
	notech_inv i_2112488(.A(i_psram_sub_mem_addr[13]), .Z(n_3491584));
	notech_nand2 i_2122487(.A(n_3491584), .B(n_2421653), .Z(n_3501583));
	notech_nand2 i_2132486(.A(i_psram_sub_mem_addr[13]), .B(n_3461585), .Z(n_3471582
		));
	notech_nand2 i_2142485(.A(n_3471582), .B(n_3501583), .Z(n_3481581));
	notech_inv i_2152484(.A(n_3481581), .Z(i_psram_sub_function_plus_2[13])
		);
	notech_inv i_2162483(.A(n_2431652), .Z(n_3511580));
	notech_inv i_2172482(.A(i_psram_sub_mem_addr[14]), .Z(n_3541579));
	notech_nand2 i_2182481(.A(n_3541579), .B(n_2431652), .Z(n_3551578));
	notech_nand2 i_2192480(.A(i_psram_sub_mem_addr[14]), .B(n_3511580), .Z(n_3521577
		));
	notech_nand2 i_2202479(.A(n_3521577), .B(n_3551578), .Z(n_3531576));
	notech_inv i_2212478(.A(n_3531576), .Z(i_psram_sub_function_plus_2[14])
		);
	notech_inv i_2222477(.A(n_2441651), .Z(n_3561575));
	notech_inv i_2232476(.A(i_psram_sub_mem_addr[15]), .Z(n_3591574));
	notech_nand2 i_2242475(.A(n_3591574), .B(n_2441651), .Z(n_3601573));
	notech_nand2 i_2252474(.A(i_psram_sub_mem_addr[15]), .B(n_3561575), .Z(n_3571572
		));
	notech_nand2 i_2262473(.A(n_3571572), .B(n_3601573), .Z(n_3581571));
	notech_inv i_2272472(.A(n_3581571), .Z(i_psram_sub_function_plus_2[15])
		);
	notech_inv i_2282471(.A(n_2821650), .Z(n_3611570));
	notech_inv i_2292470(.A(i_psram_sub_mem_addr[16]), .Z(n_3641569));
	notech_nand2 i_2302469(.A(n_3641569), .B(n_2821650), .Z(n_3651568));
	notech_nand2 i_2312468(.A(i_psram_sub_mem_addr[16]), .B(n_3611570), .Z(n_3621567
		));
	notech_nand2 i_2322467(.A(n_3621567), .B(n_3651568), .Z(n_3631566));
	notech_inv i_2332466(.A(n_3631566), .Z(i_psram_sub_function_plus_2[16])
		);
	notech_inv i_2342465(.A(n_2461649), .Z(n_3661565));
	notech_inv i_2352464(.A(i_psram_sub_mem_addr[17]), .Z(n_3691564));
	notech_nand2 i_2362463(.A(n_3691564), .B(n_2461649), .Z(n_3701563));
	notech_nand2 i_2372462(.A(i_psram_sub_mem_addr[17]), .B(n_3661565), .Z(n_3671562
		));
	notech_nand2 i_2382461(.A(n_3671562), .B(n_3701563), .Z(n_3681561));
	notech_inv i_2392460(.A(n_3681561), .Z(i_psram_sub_function_plus_2[17])
		);
	notech_inv i_2402459(.A(n_2471648), .Z(n_3711560));
	notech_inv i_2412458(.A(i_psram_sub_mem_addr[18]), .Z(n_3741559));
	notech_nand2 i_2422457(.A(n_3741559), .B(n_2471648), .Z(n_3751558));
	notech_nand2 i_2432456(.A(i_psram_sub_mem_addr[18]), .B(n_3711560), .Z(n_3721557
		));
	notech_nand2 i_2442455(.A(n_3721557), .B(n_3751558), .Z(n_3731556));
	notech_inv i_2452454(.A(n_3731556), .Z(i_psram_sub_function_plus_2[18])
		);
	notech_inv i_2462453(.A(n_2481647), .Z(n_3761555));
	notech_inv i_2472452(.A(i_psram_sub_mem_addr[19]), .Z(n_3791554));
	notech_nand2 i_2482451(.A(n_3791554), .B(n_2481647), .Z(n_3801553));
	notech_nand2 i_2492450(.A(i_psram_sub_mem_addr[19]), .B(n_3761555), .Z(n_3771552
		));
	notech_nand2 i_2502449(.A(n_3771552), .B(n_3801553), .Z(n_3781551));
	notech_inv i_2512448(.A(n_3781551), .Z(i_psram_sub_function_plus_2[19])
		);
	notech_inv i_2522447(.A(n_2491646), .Z(n_381));
	notech_inv i_2532446(.A(i_psram_sub_mem_addr[20]), .Z(n_384));
	notech_nand2 i_2542445(.A(n_384), .B(n_2491646), .Z(n_385));
	notech_nand2 i_2552444(.A(i_psram_sub_mem_addr[20]), .B(n_381), .Z(n_382
		));
	notech_nand2 i_2562443(.A(n_382), .B(n_385), .Z(n_383));
	notech_inv i_2572442(.A(n_383), .Z(i_psram_sub_function_plus_2[20]));
	notech_inv i_258(.A(n_250), .Z(n_3861550));
	notech_inv i_259(.A(i_psram_sub_mem_addr[21]), .Z(n_3891549));
	notech_nand2 i_260(.A(n_3891549), .B(n_250), .Z(n_3901548));
	notech_nand2 i_261(.A(i_psram_sub_mem_addr[21]), .B(n_3861550), .Z(n_3871547
		));
	notech_nand2 i_262(.A(n_3871547), .B(n_3901548), .Z(n_3881546));
	notech_inv i_263(.A(n_3881546), .Z(i_psram_sub_function_plus_2[21]));
	notech_inv i_2642441(.A(n_251), .Z(n_3911545));
	notech_inv i_2652440(.A(i_psram_sub_mem_addr[22]), .Z(n_3941544));
	notech_nand2 i_2662439(.A(n_3941544), .B(n_251), .Z(n_3951543));
	notech_nand2 i_2672438(.A(i_psram_sub_mem_addr[22]), .B(n_3911545), .Z(n_3921542
		));
	notech_nand2 i_2682437(.A(n_3921542), .B(n_3951543), .Z(n_3931541));
	notech_inv i_269(.A(n_3931541), .Z(i_psram_sub_function_plus_2[22]));
	notech_inv i_122436(.A(n_2491525), .Z(n_3711414));
	notech_inv i_172435(.A(n_4181343), .Z(n_4691274));
	notech_inv i_492434(.A(n_2421532), .Z(n_3631422));
	notech_inv i_591707(.A(n_2421532), .Z(n_6251413));
	notech_inv i_592433(.A(i_psram_sub_axi_awaddr[1]), .Z(n_2651524));
	notech_inv i_602432(.A(i_psram_sub_axi_awaddr[10]), .Z(n_2741515));
	notech_inv i_611706(.A(n_6421389), .Z(n_6901309));
	notech_inv i_612431(.A(i_psram_sub_axi_awaddr[11]), .Z(n_2751514));
	notech_inv i_621705(.A(i_psram_sub_axi_awaddr[11]), .Z(n_6021456));
	notech_inv i_622430(.A(i_psram_sub_axi_awaddr[12]), .Z(n_2761513));
	notech_inv i_631704(.A(n_6011455), .Z(n_6491378));
	notech_inv i_632429(.A(i_psram_sub_axi_awaddr[13]), .Z(n_2771512));
	notech_inv i_641703(.A(i_psram_sub_axi_awaddr[13]), .Z(n_6061450));
	notech_inv i_642428(.A(i_psram_sub_axi_awaddr[14]), .Z(n_2781511));
	notech_inv i_651702(.A(n_6891308), .Z(n_7371232));
	notech_inv i_652427(.A(i_psram_sub_axi_awaddr[15]), .Z(n_2791510));
	notech_inv i_661701(.A(i_psram_sub_axi_awaddr[15]), .Z(n_6101444));
	notech_inv i_662426(.A(i_psram_sub_axi_awaddr[16]), .Z(n_2801509));
	notech_inv i_671700(.A(n_6091443), .Z(n_6571366));
	notech_inv i_672425(.A(i_psram_sub_axi_awaddr[17]), .Z(n_2811508));
	notech_inv i_681699(.A(i_psram_sub_axi_awaddr[17]), .Z(n_6141438));
	notech_inv i_682424(.A(i_psram_sub_axi_awaddr[18]), .Z(n_2821507));
	notech_inv i_691698(.A(n_6581365), .Z(n_7061285));
	notech_inv i_692423(.A(i_psram_sub_axi_awaddr[19]), .Z(n_2831506));
	notech_inv i_701697(.A(i_psram_sub_axi_awaddr[19]), .Z(n_6181432));
	notech_inv i_702422(.A(i_psram_sub_axi_awaddr[20]), .Z(n_2841505));
	notech_inv i_711696(.A(n_6171431), .Z(n_6651354));
	notech_inv i_711695(.A(i_psram_sub_axi_awaddr[21]), .Z(n_2851504));
	notech_inv i_741694(.A(i_psram_sub_axi_awaddr[21]), .Z(n_6221426));
	notech_inv i_741693(.A(i_psram_sub_axi_awaddr[22]), .Z(n_2861503));
	notech_inv i_741692(.A(n_4171344), .Z(n_4681275));
	notech_inv i_761691(.A(n_6401392), .Z(n_6881312));
	notech_inv i_761690(.A(i_psram_sub_axi_awaddr[10]), .Z(n_6001459));
	notech_inv i_761689(.A(n_5991458), .Z(n_6471381));
	notech_inv i_761688(.A(i_psram_sub_axi_awaddr[12]), .Z(n_6041453));
	notech_inv i_761687(.A(n_6871311), .Z(n_7351235));
	notech_inv i_761686(.A(i_psram_sub_axi_awaddr[14]), .Z(n_6081447));
	notech_inv i_761685(.A(n_6071446), .Z(n_6551369));
	notech_inv i_761684(.A(i_psram_sub_axi_awaddr[16]), .Z(n_6121441));
	notech_inv i_761683(.A(n_6561368), .Z(n_7041288));
	notech_inv i_761682(.A(i_psram_sub_axi_awaddr[18]), .Z(n_6161435));
	notech_inv i_761681(.A(n_6151434), .Z(n_6631357));
	notech_inv i_761680(.A(i_psram_sub_axi_awaddr[20]), .Z(n_6201429));
	notech_inv i_741679(.A(n_4671276), .Z(n_5221224));
	notech_inv i_761678(.A(n_5971461), .Z(n_6451384));
	notech_inv i_761677(.A(n_6851314), .Z(n_7331238));
	notech_inv i_761676(.A(n_6051449), .Z(n_6531372));
	notech_inv i_761675(.A(n_6541371), .Z(n_7021291));
	notech_inv i_761674(.A(n_6131437), .Z(n_6611360));
	notech_inv i_741673(.A(n_3701415), .Z(n_4191342));
	notech_inv i_741672(.A(n_4661277), .Z(n_5211225));
	notech_inv i_741671(.A(n_3641421), .Z(n_4111350));
	notech_inv i_761670(.A(n_5951463), .Z(n_6431387));
	notech_inv i_761669(.A(n_6831317), .Z(n_7311241));
	notech_inv i_761668(.A(n_6031452), .Z(n_6511375));
	notech_inv i_761667(.A(n_6521374), .Z(n_7001294));
	notech_inv i_761666(.A(n_6111440), .Z(n_6591363));
	notech_inv i_741665(.A(n_4651278), .Z(n_5201226));
	notech_inv i_761664(.A(n_6811320), .Z(n_7291244));
	notech_inv i_761663(.A(n_6501377), .Z(n_6981297));
	notech_inv i_761662(.A(n_4641279), .Z(n_7441213));
	notech_inv i_761661(.A(n_6791323), .Z(n_7271247));
	notech_inv i_761660(.A(n_6481380), .Z(n_6961300));
	notech_inv i_741659(.A(n_2491525), .Z(n_4711273));
	notech_inv i_761658(.A(n_6461383), .Z(n_6941303));
	notech_inv i_762421(.A(n_6441386), .Z(n_6921306));
	notech_inv i_741657(.A(n_2941500), .Z(n_7671193));
	notech_inv i_742420(.A(i_psram_sub_axi_awaddr[1]), .Z(n_7621194));
	notech_inv i_1250(.A(i_psram_sub_axi_awaddr[0]), .Z(n_7571195));
	notech_inv i_22419(.A(s00_axi_awlen[0]), .Z(n_2181540));
	notech_inv i_32418(.A(s00_axi_awlen[1]), .Z(n_2191539));
	notech_inv i_42417(.A(s00_axi_awlen[2]), .Z(n_2201538));
	notech_inv i_52416(.A(s00_axi_awlen[3]), .Z(n_2211537));
	notech_inv i_62415(.A(s00_axi_awlen[4]), .Z(n_2221536));
	notech_inv i_72414(.A(s00_axi_awlen[5]), .Z(n_2231535));
	notech_inv i_82413(.A(s00_axi_awlen[6]), .Z(n_2241534));
	notech_inv i_92412(.A(s00_axi_awlen[7]), .Z(n_2251533));
	notech_nor2 i_262411(.A(i_psram_sub_axi_awaddr[2]), .B(n_2181540), .Z(n_2421532
		));
	notech_nor2 i_272410(.A(i_psram_sub_axi_awaddr[3]), .B(n_2191539), .Z(n_2431531
		));
	notech_nor2 i_282409(.A(i_psram_sub_axi_awaddr[4]), .B(n_2201538), .Z(n_2441530
		));
	notech_nor2 i_292408(.A(i_psram_sub_axi_awaddr[5]), .B(n_2211537), .Z(n_2451529
		));
	notech_nor2 i_302407(.A(i_psram_sub_axi_awaddr[6]), .B(n_2221536), .Z(n_2461528
		));
	notech_nor2 i_312406(.A(i_psram_sub_axi_awaddr[7]), .B(n_2231535), .Z(n_2471527
		));
	notech_nor2 i_322405(.A(i_psram_sub_axi_awaddr[8]), .B(n_2241534), .Z(n_2481526
		));
	notech_nor2 i_332404(.A(i_psram_sub_axi_awaddr[9]), .B(n_2251533), .Z(n_2491525
		));
	notech_nand2 i_502403(.A(i_psram_sub_axi_awaddr[2]), .B(n_2181540), .Z(n_2661523
		));
	notech_nand2 i_512402(.A(i_psram_sub_axi_awaddr[3]), .B(n_2191539), .Z(n_2671522
		));
	notech_nand2 i_522401(.A(i_psram_sub_axi_awaddr[4]), .B(n_2201538), .Z(n_2681521
		));
	notech_nand2 i_532400(.A(i_psram_sub_axi_awaddr[5]), .B(n_2211537), .Z(n_2691520
		));
	notech_nand2 i_542399(.A(i_psram_sub_axi_awaddr[6]), .B(n_2221536), .Z(n_2701519
		));
	notech_nand2 i_552398(.A(i_psram_sub_axi_awaddr[7]), .B(n_2231535), .Z(n_2711518
		));
	notech_nand2 i_562397(.A(i_psram_sub_axi_awaddr[8]), .B(n_2241534), .Z(n_2721517
		));
	notech_nand2 i_572396(.A(i_psram_sub_axi_awaddr[9]), .B(n_2251533), .Z(n_2731516
		));
	notech_inv i_722395(.A(i_psram_sub_axi_awaddr[0]), .Z(n_2881502));
	notech_inv i_772394(.A(n_2421532), .Z(n_2931501));
	notech_nand2 i_782393(.A(n_2931501), .B(n_2661523), .Z(n_2941500));
	notech_inv i_792392(.A(n_2431531), .Z(n_2951499));
	notech_nand2 i_802391(.A(n_2951499), .B(n_2671522), .Z(n_2961498));
	notech_inv i_812390(.A(n_2441530), .Z(n_2971497));
	notech_nand2 i_822389(.A(n_2971497), .B(n_2681521), .Z(n_2981496));
	notech_inv i_832388(.A(n_2451529), .Z(n_2991495));
	notech_nand2 i_842387(.A(n_2991495), .B(n_2691520), .Z(n_3001494));
	notech_inv i_852386(.A(n_2461528), .Z(n_3011493));
	notech_nand2 i_862385(.A(n_3011493), .B(n_2701519), .Z(n_3021492));
	notech_inv i_872384(.A(n_2471527), .Z(n_3031491));
	notech_nand2 i_882383(.A(n_3031491), .B(n_2711518), .Z(n_3041490));
	notech_inv i_892382(.A(n_2481526), .Z(n_3051489));
	notech_nand2 i_902381(.A(n_3051489), .B(n_2721517), .Z(n_3061488));
	notech_inv i_912380(.A(n_2491525), .Z(n_3071487));
	notech_nand2 i_922379(.A(n_3071487), .B(n_2731516), .Z(n_3081486));
	notech_or2 i_3602378(.A(n_2421532), .B(n_2651524), .Z(n_5821485));
	notech_and2 i_3612377(.A(n_5821485), .B(n_2661523), .Z(n_5811484));
	notech_inv i_3622376(.A(n_5811484), .Z(n_3391483));
	notech_or2 i_3632375(.A(n_2431531), .B(n_2661523), .Z(n_5841482));
	notech_and2 i_3642374(.A(n_5841482), .B(n_2671522), .Z(n_5831481));
	notech_inv i_3652373(.A(n_5831481), .Z(n_3401480));
	notech_or2 i_3662372(.A(n_2441530), .B(n_2671522), .Z(n_5861479));
	notech_and2 i_3672371(.A(n_5861479), .B(n_2681521), .Z(n_5851478));
	notech_inv i_3682370(.A(n_5851478), .Z(n_3411477));
	notech_or2 i_3692369(.A(n_2451529), .B(n_2681521), .Z(n_5881476));
	notech_and2 i_3702368(.A(n_5881476), .B(n_2691520), .Z(n_5871475));
	notech_inv i_3712367(.A(n_5871475), .Z(n_3421474));
	notech_or2 i_3722366(.A(n_2461528), .B(n_2691520), .Z(n_5901473));
	notech_and2 i_3732365(.A(n_5901473), .B(n_2701519), .Z(n_5891472));
	notech_inv i_3742364(.A(n_5891472), .Z(n_3431471));
	notech_or2 i_3752363(.A(n_2471527), .B(n_2701519), .Z(n_5921470));
	notech_and2 i_3762362(.A(n_5921470), .B(n_2711518), .Z(n_5911469));
	notech_inv i_3772361(.A(n_5911469), .Z(n_3441468));
	notech_or2 i_3782360(.A(n_2481526), .B(n_2711518), .Z(n_5941467));
	notech_and2 i_3792359(.A(n_5941467), .B(n_2721517), .Z(n_5931466));
	notech_inv i_3802358(.A(n_5931466), .Z(n_3451465));
	notech_or2 i_3812357(.A(n_2491525), .B(n_2721517), .Z(n_5961464));
	notech_and2 i_3822356(.A(n_5961464), .B(n_2731516), .Z(n_5951463));
	notech_inv i_3832355(.A(n_5951463), .Z(n_3461462));
	notech_and2 i_3852354(.A(n_2731516), .B(n_2741515), .Z(n_5971461));
	notech_inv i_3862353(.A(n_5971461), .Z(n_3471460));
	notech_and2 i_3882352(.A(n_6001459), .B(n_2751514), .Z(n_5991458));
	notech_inv i_3892351(.A(n_5991458), .Z(n_3481457));
	notech_and2 i_3912350(.A(n_6021456), .B(n_2761513), .Z(n_6011455));
	notech_inv i_3922349(.A(n_6011455), .Z(n_3491454));
	notech_and2 i_3942348(.A(n_6041453), .B(n_2771512), .Z(n_6031452));
	notech_inv i_3952347(.A(n_6031452), .Z(n_3501451));
	notech_and2 i_3972346(.A(n_6061450), .B(n_2781511), .Z(n_6051449));
	notech_inv i_3982345(.A(n_6051449), .Z(n_3511448));
	notech_and2 i_4002344(.A(n_6081447), .B(n_2791510), .Z(n_6071446));
	notech_inv i_4012343(.A(n_6071446), .Z(n_3521445));
	notech_and2 i_4032342(.A(n_6101444), .B(n_2801509), .Z(n_6091443));
	notech_inv i_4042341(.A(n_6091443), .Z(n_3531442));
	notech_and2 i_4062340(.A(n_6121441), .B(n_2811508), .Z(n_6111440));
	notech_inv i_4072339(.A(n_6111440), .Z(n_3541439));
	notech_and2 i_4092338(.A(n_6141438), .B(n_2821507), .Z(n_6131437));
	notech_inv i_4102337(.A(n_6131437), .Z(n_3551436));
	notech_and2 i_4122336(.A(n_6161435), .B(n_2831506), .Z(n_6151434));
	notech_inv i_4132335(.A(n_6151434), .Z(n_3561433));
	notech_and2 i_4152334(.A(n_6181432), .B(n_2841505), .Z(n_6171431));
	notech_inv i_4162333(.A(n_6171431), .Z(n_3571430));
	notech_and2 i_4182332(.A(n_6201429), .B(n_2851504), .Z(n_6191428));
	notech_inv i_4192331(.A(n_6191428), .Z(n_3581427));
	notech_and2 i_4212330(.A(n_6221426), .B(n_2861503), .Z(n_6211425));
	notech_inv i_4222329(.A(n_6211425), .Z(n_3591424));
	notech_inv i_1442328(.A(n_2881502), .Z(n_3601423));
	notech_nor2 i_1482327(.A(n_2421532), .B(n_2431531), .Z(n_3641421));
	notech_nor2 i_1492326(.A(n_2431531), .B(n_2441530), .Z(n_3651420));
	notech_nor2 i_1502325(.A(n_2441530), .B(n_2451529), .Z(n_3661419));
	notech_nor2 i_1512324(.A(n_2451529), .B(n_2461528), .Z(n_3671418));
	notech_nor2 i_1522323(.A(n_2461528), .B(n_2471527), .Z(n_3681417));
	notech_nor2 i_1532322(.A(n_2471527), .B(n_2481526), .Z(n_3691416));
	notech_nor2 i_1542321(.A(n_2481526), .B(n_2491525), .Z(n_3701415));
	notech_or2 i_4272320(.A(n_6251413), .B(n_3391483), .Z(n_6261412));
	notech_inv i_4282319(.A(n_6261412), .Z(n_3861411));
	notech_or2 i_4302318(.A(n_3641421), .B(n_3401480), .Z(n_6281410));
	notech_inv i_4312317(.A(n_6281410), .Z(n_3871409));
	notech_and2 i_4322316(.A(n_3651420), .B(n_3391483), .Z(n_6291408));
	notech_or2 i_4332315(.A(n_6291408), .B(n_3411477), .Z(n_6301407));
	notech_inv i_4342314(.A(n_6301407), .Z(n_3881406));
	notech_and2 i_4352313(.A(n_3661419), .B(n_3401480), .Z(n_6311405));
	notech_or2 i_4362312(.A(n_6311405), .B(n_3421474), .Z(n_6321404));
	notech_inv i_4372311(.A(n_6321404), .Z(n_3891403));
	notech_and2 i_4382310(.A(n_3671418), .B(n_3411477), .Z(n_6331402));
	notech_or2 i_4392309(.A(n_6331402), .B(n_3431471), .Z(n_6341401));
	notech_inv i_4402308(.A(n_6341401), .Z(n_3901400));
	notech_and2 i_4412307(.A(n_3681417), .B(n_3421474), .Z(n_6351399));
	notech_or2 i_4422306(.A(n_6351399), .B(n_3441468), .Z(n_6361398));
	notech_inv i_4432305(.A(n_6361398), .Z(n_3911397));
	notech_and2 i_4442304(.A(n_3691416), .B(n_3431471), .Z(n_6371396));
	notech_or2 i_4452303(.A(n_6371396), .B(n_3451465), .Z(n_6381395));
	notech_inv i_4462302(.A(n_6381395), .Z(n_3921394));
	notech_and2 i_4472301(.A(n_3701415), .B(n_3441468), .Z(n_6391393));
	notech_or2 i_4482300(.A(n_6391393), .B(n_3461462), .Z(n_6401392));
	notech_inv i_4492299(.A(n_6401392), .Z(n_3931391));
	notech_and2 i_4502298(.A(n_3711414), .B(n_3451465), .Z(n_6411390));
	notech_or2 i_4512297(.A(n_6411390), .B(n_3471460), .Z(n_6421389));
	notech_inv i_4522296(.A(n_6421389), .Z(n_3941388));
	notech_or2 i_4542295(.A(n_6431387), .B(n_3481457), .Z(n_6441386));
	notech_inv i_4552294(.A(n_6441386), .Z(n_3951385));
	notech_or2 i_4572293(.A(n_6451384), .B(n_3491454), .Z(n_6461383));
	notech_inv i_4582292(.A(n_6461383), .Z(n_3961382));
	notech_or2 i_4602291(.A(n_6471381), .B(n_3501451), .Z(n_6481380));
	notech_inv i_4612290(.A(n_6481380), .Z(n_3971379));
	notech_or2 i_4632289(.A(n_6491378), .B(n_3511448), .Z(n_6501377));
	notech_inv i_4642288(.A(n_6501377), .Z(n_3981376));
	notech_or2 i_4662287(.A(n_6511375), .B(n_3521445), .Z(n_6521374));
	notech_inv i_4672286(.A(n_6521374), .Z(n_3991373));
	notech_or2 i_4692285(.A(n_6531372), .B(n_3531442), .Z(n_6541371));
	notech_inv i_4702284(.A(n_6541371), .Z(n_4001370));
	notech_or2 i_4722283(.A(n_6551369), .B(n_3541439), .Z(n_6561368));
	notech_inv i_4732282(.A(n_6561368), .Z(n_4011367));
	notech_or2 i_4752281(.A(n_6571366), .B(n_3551436), .Z(n_6581365));
	notech_inv i_4762280(.A(n_6581365), .Z(n_4021364));
	notech_or2 i_4782279(.A(n_6591363), .B(n_3561433), .Z(n_6601362));
	notech_inv i_4792278(.A(n_6601362), .Z(n_4031361));
	notech_or2 i_4812277(.A(n_6611360), .B(n_3571430), .Z(n_6621359));
	notech_inv i_4822276(.A(n_6621359), .Z(n_4041358));
	notech_or2 i_4842275(.A(n_6631357), .B(n_3581427), .Z(n_6641356));
	notech_inv i_4852274(.A(n_6641356), .Z(n_4051355));
	notech_or2 i_4872273(.A(n_6651354), .B(n_3591424), .Z(n_6661353));
	notech_inv i_4882272(.A(n_6661353), .Z(n_4061352));
	notech_inv i_1912271(.A(n_3601423), .Z(n_4071351));
	notech_nand2 i_1962270(.A(n_3631422), .B(n_3651420), .Z(n_4121349));
	notech_nand2 i_1972269(.A(n_3641421), .B(n_3661419), .Z(n_4131348));
	notech_nand2 i_1982268(.A(n_3651420), .B(n_3671418), .Z(n_4141347));
	notech_nand2 i_1992267(.A(n_3661419), .B(n_3681417), .Z(n_4151346));
	notech_nand2 i_2002266(.A(n_3671418), .B(n_3691416), .Z(n_4161345));
	notech_nand2 i_2012265(.A(n_3681417), .B(n_3701415), .Z(n_4171344));
	notech_nand2 i_2022264(.A(n_3691416), .B(n_3711414), .Z(n_4181343));
	notech_inv i_2172263(.A(n_3861411), .Z(n_4331341));
	notech_or2 i_4892262(.A(n_4111350), .B(n_4071351), .Z(n_6681340));
	notech_and2 i_4902261(.A(n_6681340), .B(n_3871409), .Z(n_6671339));
	notech_inv i_4912260(.A(n_6671339), .Z(n_4341338));
	notech_and2 i_4932259(.A(n_4121349), .B(n_3881406), .Z(n_6691337));
	notech_inv i_4942258(.A(n_6691337), .Z(n_4351336));
	notech_and2 i_4962257(.A(n_4131348), .B(n_3891403), .Z(n_6711335));
	notech_inv i_4972256(.A(n_6711335), .Z(n_4361334));
	notech_or2 i_4982255(.A(n_4141347), .B(n_3861411), .Z(n_6741333));
	notech_and2 i_4992254(.A(n_6741333), .B(n_3901400), .Z(n_6731332));
	notech_inv i_5002253(.A(n_6731332), .Z(n_4371331));
	notech_or2 i_5012252(.A(n_4151346), .B(n_3871409), .Z(n_6761330));
	notech_and2 i_5022251(.A(n_6761330), .B(n_3911397), .Z(n_6751329));
	notech_inv i_5032250(.A(n_6751329), .Z(n_4381328));
	notech_or2 i_5042249(.A(n_4161345), .B(n_3881406), .Z(n_6781327));
	notech_and2 i_5052248(.A(n_6781327), .B(n_3921394), .Z(n_6771326));
	notech_inv i_5062247(.A(n_6771326), .Z(n_4391325));
	notech_or2 i_5072246(.A(n_4171344), .B(n_3891403), .Z(n_6801324));
	notech_and2 i_5082245(.A(n_6801324), .B(n_3931391), .Z(n_6791323));
	notech_inv i_5092244(.A(n_6791323), .Z(n_4401322));
	notech_or2 i_5102243(.A(n_4181343), .B(n_3901400), .Z(n_6821321));
	notech_and2 i_5112242(.A(n_6821321), .B(n_3941388), .Z(n_6811320));
	notech_inv i_5122241(.A(n_6811320), .Z(n_4411319));
	notech_or2 i_5132240(.A(n_4191342), .B(n_3911397), .Z(n_6841318));
	notech_and2 i_5142239(.A(n_6841318), .B(n_3951385), .Z(n_6831317));
	notech_inv i_5152238(.A(n_6831317), .Z(n_4421316));
	notech_or2 i_5162237(.A(n_2491525), .B(n_3921394), .Z(n_6861315));
	notech_and2 i_5172236(.A(n_6861315), .B(n_3961382), .Z(n_6851314));
	notech_inv i_5182235(.A(n_6851314), .Z(n_4431313));
	notech_and2 i_5202234(.A(n_6881312), .B(n_3971379), .Z(n_6871311));
	notech_inv i_5212233(.A(n_6871311), .Z(n_4441310));
	notech_and2 i_5232232(.A(n_6901309), .B(n_3981376), .Z(n_6891308));
	notech_inv i_5242231(.A(n_6891308), .Z(n_4451307));
	notech_and2 i_5262230(.A(n_6921306), .B(n_3991373), .Z(n_6911305));
	notech_inv i_5272229(.A(n_6911305), .Z(n_4461304));
	notech_and2 i_5292228(.A(n_6941303), .B(n_4001370), .Z(n_6931302));
	notech_inv i_5302227(.A(n_6931302), .Z(n_4471301));
	notech_and2 i_5322226(.A(n_6961300), .B(n_4011367), .Z(n_6951299));
	notech_inv i_5332225(.A(n_6951299), .Z(n_4481298));
	notech_and2 i_5352224(.A(n_6981297), .B(n_4021364), .Z(n_6971296));
	notech_inv i_5362223(.A(n_6971296), .Z(n_4491295));
	notech_and2 i_5382222(.A(n_7001294), .B(n_4031361), .Z(n_6991293));
	notech_inv i_5392221(.A(n_6991293), .Z(n_4501292));
	notech_and2 i_5412220(.A(n_7021291), .B(n_4041358), .Z(n_7011290));
	notech_inv i_5422219(.A(n_7011290), .Z(n_4511289));
	notech_and2 i_5442218(.A(n_7041288), .B(n_4051355), .Z(n_7031287));
	notech_inv i_5452217(.A(n_7031287), .Z(n_4521286));
	notech_and2 i_5472216(.A(n_7061285), .B(n_4061352), .Z(n_7051284));
	notech_inv i_5482215(.A(n_7051284), .Z(n_4531283));
	notech_inv i_2382214(.A(n_4071351), .Z(n_4541282));
	notech_nor2 i_2462213(.A(n_4111350), .B(n_4151346), .Z(n_4621281));
	notech_nor2 i_2472212(.A(n_4121349), .B(n_4161345), .Z(n_4631280));
	notech_nor2 i_2482211(.A(n_4131348), .B(n_4171344), .Z(n_4641279));
	notech_nor2 i_2492210(.A(n_4141347), .B(n_4181343), .Z(n_4651278));
	notech_nor2 i_2502209(.A(n_4151346), .B(n_4191342), .Z(n_4661277));
	notech_nor2 i_2512208(.A(n_4161345), .B(n_2491525), .Z(n_4671276));
	notech_inv i_2642207(.A(n_4331341), .Z(n_4801272));
	notech_inv i_2652206(.A(n_4341338), .Z(n_4811271));
	notech_inv i_2662205(.A(n_4351336), .Z(n_4821270));
	notech_inv i_2672204(.A(n_4361334), .Z(n_4831269));
	notech_inv i_2682203(.A(n_4371331), .Z(n_4841268));
	notech_and2 i_5492202(.A(n_4621281), .B(n_4541282), .Z(n_7071267));
	notech_or2 i_5502201(.A(n_7071267), .B(n_4381328), .Z(n_7081266));
	notech_or2 i_5532200(.A(n_4631280), .B(n_4391325), .Z(n_7101265));
	notech_or2 i_5562199(.A(n_4641279), .B(n_4401322), .Z(n_7121264));
	notech_and2 i_5582198(.A(n_4651278), .B(n_4331341), .Z(n_7131263));
	notech_or2 i_5592197(.A(n_7131263), .B(n_4411319), .Z(n_7141262));
	notech_and2 i_5612196(.A(n_4661277), .B(n_4341338), .Z(n_7151261));
	notech_or2 i_5622195(.A(n_7151261), .B(n_4421316), .Z(n_7161260));
	notech_and2 i_5642194(.A(n_4671276), .B(n_4351336), .Z(n_7171259));
	notech_or2 i_5652193(.A(n_7171259), .B(n_4431313), .Z(n_7181258));
	notech_and2 i_5672192(.A(n_4681275), .B(n_4361334), .Z(n_7191257));
	notech_or2 i_5682191(.A(n_7191257), .B(n_4441310), .Z(n_7201256));
	notech_and2 i_5702190(.A(n_4691274), .B(n_4371331), .Z(n_7211255));
	notech_or2 i_5712189(.A(n_7211255), .B(n_4451307), .Z(n_7221254));
	notech_and2 i_5732188(.A(n_3701415), .B(n_4381328), .Z(n_7231253));
	notech_or2 i_5742187(.A(n_7231253), .B(n_4461304), .Z(n_7241252));
	notech_inv i_5752186(.A(n_7241252), .Z(n_4931251));
	notech_and2 i_5762185(.A(n_4711273), .B(n_4391325), .Z(n_7251250));
	notech_or2 i_5772184(.A(n_7251250), .B(n_4471301), .Z(n_7261249));
	notech_inv i_5782183(.A(n_7261249), .Z(n_4941248));
	notech_or2 i_5802182(.A(n_7271247), .B(n_4481298), .Z(n_7281246));
	notech_inv i_5812181(.A(n_7281246), .Z(n_4951245));
	notech_or2 i_5832180(.A(n_7291244), .B(n_4491295), .Z(n_7301243));
	notech_inv i_5842179(.A(n_7301243), .Z(n_4961242));
	notech_or2 i_5862178(.A(n_7311241), .B(n_4501292), .Z(n_7321240));
	notech_inv i_5872177(.A(n_7321240), .Z(n_4971239));
	notech_or2 i_5892176(.A(n_7331238), .B(n_4511289), .Z(n_7341237));
	notech_inv i_5902175(.A(n_7341237), .Z(n_4981236));
	notech_or2 i_5922174(.A(n_7351235), .B(n_4521286), .Z(n_7361234));
	notech_inv i_5932173(.A(n_7361234), .Z(n_4991233));
	notech_or2 i_5952172(.A(n_7371232), .B(n_4531283), .Z(n_7381231));
	notech_inv i_5962171(.A(n_7381231), .Z(n_5001230));
	notech_inv i_2852170(.A(n_4541282), .Z(n_5011229));
	notech_nand2 i_3012169(.A(n_4621281), .B(n_3701415), .Z(n_5171228));
	notech_nand2 i_3022168(.A(n_4631280), .B(n_4711273), .Z(n_5181227));
	notech_inv i_3112167(.A(n_4801272), .Z(n_5271223));
	notech_inv i_3122166(.A(n_4811271), .Z(n_5281222));
	notech_inv i_3132165(.A(n_4821270), .Z(n_5291221));
	notech_inv i_3142164(.A(n_4831269), .Z(n_5301220));
	notech_inv i_3152163(.A(n_4841268), .Z(n_5311219));
	notech_or2 i_5972162(.A(n_5171228), .B(n_5011229), .Z(n_7401218));
	notech_and2 i_5982161(.A(n_7401218), .B(n_4931251), .Z(n_7391217));
	notech_inv i_5992160(.A(n_7391217), .Z(n_5401216));
	notech_and2 i_6012159(.A(n_5181227), .B(n_4941248), .Z(n_7411215));
	notech_inv i_6022158(.A(n_7411215), .Z(n_5411214));
	notech_and2 i_6042157(.A(n_7441213), .B(n_4951245), .Z(n_7431212));
	notech_inv i_6052156(.A(n_7431212), .Z(n_5421211));
	notech_or2 i_6062155(.A(n_5201226), .B(n_4801272), .Z(n_7461210));
	notech_and2 i_6072154(.A(n_7461210), .B(n_4961242), .Z(n_7451209));
	notech_inv i_6082153(.A(n_7451209), .Z(n_5431208));
	notech_or2 i_6092152(.A(n_5211225), .B(n_4811271), .Z(n_7481207));
	notech_and2 i_6102151(.A(n_7481207), .B(n_4971239), .Z(n_7471206));
	notech_inv i_6112150(.A(n_7471206), .Z(n_5441205));
	notech_or2 i_6122149(.A(n_5221224), .B(n_4821270), .Z(n_7501204));
	notech_and2 i_6132148(.A(n_7501204), .B(n_4981236), .Z(n_7491203));
	notech_inv i_6142147(.A(n_7491203), .Z(n_5451202));
	notech_or2 i_6152146(.A(n_4171344), .B(n_4831269), .Z(n_7521201));
	notech_and2 i_6162145(.A(n_7521201), .B(n_4991233), .Z(n_7511200));
	notech_inv i_6172144(.A(n_7511200), .Z(n_5461199));
	notech_or2 i_6182143(.A(n_4181343), .B(n_4841268), .Z(n_7541198));
	notech_and2 i_6192142(.A(n_7541198), .B(n_5001230), .Z(n_7531197));
	notech_inv i_6202141(.A(n_7531197), .Z(n_5471196));
	notech_inv i_6262140(.A(n_7571195), .Z(i_psram_sub_function_sub_0[0]));
	notech_inv i_6322139(.A(n_7621194), .Z(i_psram_sub_function_sub_0[1]));
	notech_inv i_6382138(.A(n_7671193), .Z(i_psram_sub_function_sub_0[2]));
	notech_inv i_6392137(.A(n_5271223), .Z(n_7701192));
	notech_inv i_6402136(.A(n_2961498), .Z(n_7731191));
	notech_nand2 i_6412135(.A(n_7731191), .B(n_5271223), .Z(n_7741190));
	notech_nand2 i_6422134(.A(n_2961498), .B(n_7701192), .Z(n_7711189));
	notech_nand2 i_6432133(.A(n_7711189), .B(n_7741190), .Z(n_7721188));
	notech_inv i_6442132(.A(n_7721188), .Z(i_psram_sub_function_sub_0[3]));
	notech_inv i_6452131(.A(n_5281222), .Z(n_7751187));
	notech_inv i_6462130(.A(n_2981496), .Z(n_7781186));
	notech_nand2 i_6472129(.A(n_7781186), .B(n_5281222), .Z(n_7791185));
	notech_nand2 i_6482128(.A(n_2981496), .B(n_7751187), .Z(n_7761184));
	notech_nand2 i_6492127(.A(n_7761184), .B(n_7791185), .Z(n_7771183));
	notech_inv i_6502126(.A(n_7771183), .Z(i_psram_sub_function_sub_0[4]));
	notech_inv i_6512125(.A(n_5291221), .Z(n_7801182));
	notech_inv i_6522124(.A(n_3001494), .Z(n_7831181));
	notech_nand2 i_6532123(.A(n_7831181), .B(n_5291221), .Z(n_7841180));
	notech_nand2 i_6542122(.A(n_3001494), .B(n_7801182), .Z(n_7811179));
	notech_nand2 i_6552121(.A(n_7811179), .B(n_7841180), .Z(n_7821178));
	notech_inv i_6562120(.A(n_7821178), .Z(i_psram_sub_function_sub_0[5]));
	notech_inv i_6572119(.A(n_5301220), .Z(n_7851177));
	notech_inv i_6582118(.A(n_3021492), .Z(n_7881176));
	notech_nand2 i_6592117(.A(n_7881176), .B(n_5301220), .Z(n_7891175));
	notech_nand2 i_6602116(.A(n_3021492), .B(n_7851177), .Z(n_7861174));
	notech_nand2 i_6612115(.A(n_7861174), .B(n_7891175), .Z(n_7871173));
	notech_inv i_6622114(.A(n_7871173), .Z(i_psram_sub_function_sub_0[6]));
	notech_inv i_6632113(.A(n_5311219), .Z(n_7901172));
	notech_inv i_6642112(.A(n_3041490), .Z(n_7931171));
	notech_nand2 i_6652111(.A(n_7931171), .B(n_5311219), .Z(n_7941170));
	notech_nand2 i_6662110(.A(n_3041490), .B(n_7901172), .Z(n_7911169));
	notech_nand2 i_6672109(.A(n_7911169), .B(n_7941170), .Z(n_7921168));
	notech_inv i_6682108(.A(n_7921168), .Z(i_psram_sub_function_sub_0[7]));
	notech_inv i_6692107(.A(n_7081266), .Z(n_7951167));
	notech_inv i_6702106(.A(n_3061488), .Z(n_7981166));
	notech_nand2 i_6712105(.A(n_7981166), .B(n_7081266), .Z(n_7991165));
	notech_nand2 i_6722104(.A(n_3061488), .B(n_7951167), .Z(n_7961164));
	notech_nand2 i_6732103(.A(n_7961164), .B(n_7991165), .Z(n_7971163));
	notech_inv i_6742102(.A(n_7971163), .Z(i_psram_sub_function_sub_0[8]));
	notech_inv i_6752101(.A(n_7101265), .Z(n_8001162));
	notech_inv i_6762100(.A(n_3081486), .Z(n_8031161));
	notech_nand2 i_6772099(.A(n_8031161), .B(n_7101265), .Z(n_8041160));
	notech_nand2 i_6782098(.A(n_3081486), .B(n_8001162), .Z(n_8011159));
	notech_nand2 i_6792097(.A(n_8011159), .B(n_8041160), .Z(n_8021158));
	notech_inv i_6802096(.A(n_8021158), .Z(i_psram_sub_function_sub_0[9]));
	notech_inv i_6812095(.A(n_7121264), .Z(n_8051157));
	notech_inv i_6822094(.A(i_psram_sub_axi_awaddr[10]), .Z(n_8081156));
	notech_nand2 i_6832093(.A(n_8081156), .B(n_7121264), .Z(n_8091155));
	notech_nand2 i_6842092(.A(i_psram_sub_axi_awaddr[10]), .B(n_8051157), .Z
		(n_8061154));
	notech_nand2 i_6852091(.A(n_8061154), .B(n_8091155), .Z(n_8071153));
	notech_inv i_6862090(.A(n_8071153), .Z(i_psram_sub_function_sub_0[10])
		);
	notech_inv i_6872089(.A(n_7141262), .Z(n_8101152));
	notech_inv i_6882088(.A(i_psram_sub_axi_awaddr[11]), .Z(n_8131151));
	notech_nand2 i_6892087(.A(n_8131151), .B(n_7141262), .Z(n_8141150));
	notech_nand2 i_6902086(.A(i_psram_sub_axi_awaddr[11]), .B(n_8101152), .Z
		(n_8111149));
	notech_nand2 i_6912085(.A(n_8111149), .B(n_8141150), .Z(n_8121148));
	notech_inv i_6922084(.A(n_8121148), .Z(i_psram_sub_function_sub_0[11])
		);
	notech_inv i_6932083(.A(n_7161260), .Z(n_8151147));
	notech_inv i_6942082(.A(i_psram_sub_axi_awaddr[12]), .Z(n_8181146));
	notech_nand2 i_6952081(.A(n_8181146), .B(n_7161260), .Z(n_8191145));
	notech_nand2 i_6962080(.A(i_psram_sub_axi_awaddr[12]), .B(n_8151147), .Z
		(n_8161144));
	notech_nand2 i_6972079(.A(n_8161144), .B(n_8191145), .Z(n_8171143));
	notech_inv i_6982078(.A(n_8171143), .Z(i_psram_sub_function_sub_0[12])
		);
	notech_inv i_6992077(.A(n_7181258), .Z(n_8201142));
	notech_inv i_7002076(.A(i_psram_sub_axi_awaddr[13]), .Z(n_8231141));
	notech_nand2 i_7012075(.A(n_8231141), .B(n_7181258), .Z(n_8241140));
	notech_nand2 i_7022074(.A(i_psram_sub_axi_awaddr[13]), .B(n_8201142), .Z
		(n_8211139));
	notech_nand2 i_7032073(.A(n_8211139), .B(n_8241140), .Z(n_8221138));
	notech_inv i_7042072(.A(n_8221138), .Z(i_psram_sub_function_sub_0[13])
		);
	notech_inv i_7052071(.A(n_7201256), .Z(n_8251137));
	notech_inv i_7062070(.A(i_psram_sub_axi_awaddr[14]), .Z(n_8281136));
	notech_nand2 i_7072069(.A(n_8281136), .B(n_7201256), .Z(n_8291135));
	notech_nand2 i_7082068(.A(i_psram_sub_axi_awaddr[14]), .B(n_8251137), .Z
		(n_8261134));
	notech_nand2 i_7092067(.A(n_8261134), .B(n_8291135), .Z(n_8271133));
	notech_inv i_7102066(.A(n_8271133), .Z(i_psram_sub_function_sub_0[14])
		);
	notech_inv i_7112065(.A(n_7221254), .Z(n_8301132));
	notech_inv i_7122064(.A(i_psram_sub_axi_awaddr[15]), .Z(n_8331131));
	notech_nand2 i_7132063(.A(n_8331131), .B(n_7221254), .Z(n_8341130));
	notech_nand2 i_7142062(.A(i_psram_sub_axi_awaddr[15]), .B(n_8301132), .Z
		(n_8311129));
	notech_nand2 i_7152061(.A(n_8311129), .B(n_8341130), .Z(n_8321128));
	notech_inv i_7162060(.A(n_8321128), .Z(i_psram_sub_function_sub_0[15])
		);
	notech_inv i_7172059(.A(n_5401216), .Z(n_8351127));
	notech_inv i_7182058(.A(i_psram_sub_axi_awaddr[16]), .Z(n_8381126));
	notech_nand2 i_7192057(.A(n_8381126), .B(n_5401216), .Z(n_8391125));
	notech_nand2 i_7202056(.A(i_psram_sub_axi_awaddr[16]), .B(n_8351127), .Z
		(n_8361124));
	notech_nand2 i_7212055(.A(n_8361124), .B(n_8391125), .Z(n_8371123));
	notech_inv i_7222054(.A(n_8371123), .Z(i_psram_sub_function_sub_0[16])
		);
	notech_inv i_7232053(.A(n_5411214), .Z(n_8401122));
	notech_inv i_7242052(.A(i_psram_sub_axi_awaddr[17]), .Z(n_8431121));
	notech_nand2 i_7252051(.A(n_8431121), .B(n_5411214), .Z(n_8441120));
	notech_nand2 i_7262050(.A(i_psram_sub_axi_awaddr[17]), .B(n_8401122), .Z
		(n_8411119));
	notech_nand2 i_7272049(.A(n_8411119), .B(n_8441120), .Z(n_8421118));
	notech_inv i_7282048(.A(n_8421118), .Z(i_psram_sub_function_sub_0[17])
		);
	notech_inv i_7292047(.A(n_5421211), .Z(n_8451117));
	notech_inv i_7302046(.A(i_psram_sub_axi_awaddr[18]), .Z(n_8481116));
	notech_nand2 i_7312045(.A(n_8481116), .B(n_5421211), .Z(n_8491115));
	notech_nand2 i_7322044(.A(i_psram_sub_axi_awaddr[18]), .B(n_8451117), .Z
		(n_8461114));
	notech_nand2 i_7332043(.A(n_8461114), .B(n_8491115), .Z(n_8471113));
	notech_inv i_7342042(.A(n_8471113), .Z(i_psram_sub_function_sub_0[18])
		);
	notech_inv i_7352041(.A(n_5431208), .Z(n_8501112));
	notech_inv i_7362040(.A(i_psram_sub_axi_awaddr[19]), .Z(n_8531111));
	notech_nand2 i_7372039(.A(n_8531111), .B(n_5431208), .Z(n_8541110));
	notech_nand2 i_7382038(.A(i_psram_sub_axi_awaddr[19]), .B(n_8501112), .Z
		(n_8511109));
	notech_nand2 i_7392037(.A(n_8511109), .B(n_8541110), .Z(n_8521108));
	notech_inv i_7402036(.A(n_8521108), .Z(i_psram_sub_function_sub_0[19])
		);
	notech_inv i_7412035(.A(n_5441205), .Z(n_8551107));
	notech_inv i_7422034(.A(i_psram_sub_axi_awaddr[20]), .Z(n_8581106));
	notech_nand2 i_7432033(.A(n_8581106), .B(n_5441205), .Z(n_8591105));
	notech_nand2 i_7442032(.A(i_psram_sub_axi_awaddr[20]), .B(n_8551107), .Z
		(n_8561104));
	notech_nand2 i_7452031(.A(n_8561104), .B(n_8591105), .Z(n_8571103));
	notech_inv i_7462030(.A(n_8571103), .Z(i_psram_sub_function_sub_0[20])
		);
	notech_inv i_7472029(.A(n_5451202), .Z(n_8601102));
	notech_inv i_7482028(.A(i_psram_sub_axi_awaddr[21]), .Z(n_8631101));
	notech_nand2 i_7492027(.A(n_8631101), .B(n_5451202), .Z(n_8641100));
	notech_nand2 i_7502026(.A(i_psram_sub_axi_awaddr[21]), .B(n_8601102), .Z
		(n_8611099));
	notech_nand2 i_7512025(.A(n_8611099), .B(n_8641100), .Z(n_8621098));
	notech_inv i_7522024(.A(n_8621098), .Z(i_psram_sub_function_sub_0[21])
		);
	notech_inv i_7532023(.A(n_5461199), .Z(n_8651097));
	notech_inv i_7542022(.A(i_psram_sub_axi_awaddr[22]), .Z(n_8681096));
	notech_nand2 i_7552021(.A(n_8681096), .B(n_5461199), .Z(n_8691095));
	notech_nand2 i_7562020(.A(i_psram_sub_axi_awaddr[22]), .B(n_8651097), .Z
		(n_8661094));
	notech_nand2 i_7572019(.A(n_8661094), .B(n_8691095), .Z(n_8671093));
	notech_inv i_7582018(.A(n_8671093), .Z(i_psram_sub_function_sub_0[22])
		);
	notech_inv i_7592017(.A(n_5471196), .Z(n_8701092));
	notech_inv i_7602016(.A(i_psram_sub_axi_awaddr[23]), .Z(n_8731091));
	notech_nand2 i_7612015(.A(n_8731091), .B(n_5471196), .Z(n_8741090));
	notech_nand2 i_7622014(.A(i_psram_sub_axi_awaddr[23]), .B(n_8701092), .Z
		(n_8711089));
	notech_nand2 i_7632013(.A(n_8711089), .B(n_8741090), .Z(n_8721088));
	notech_inv i_7642012(.A(n_8721088), .Z(i_psram_sub_function_sub_0[23])
		);
	notech_inv i_02011(.A(i_psram_sub_axi_awaddr[2]), .Z(\i_psram_sub_axi_awaddr_0[2] 
		));
	notech_nand2 i_12010(.A(i_psram_sub_axi_awaddr[2]), .B(i_psram_sub_axi_awaddr
		[3]), .Z(n_1331071));
	notech_nand2 i_22009(.A(i_psram_sub_axi_awaddr[3]), .B(i_psram_sub_axi_awaddr
		[4]), .Z(n_1341070));
	notech_nand2 i_32008(.A(i_psram_sub_axi_awaddr[4]), .B(i_psram_sub_axi_awaddr
		[5]), .Z(n_1351069));
	notech_nand2 i_42007(.A(i_psram_sub_axi_awaddr[5]), .B(i_psram_sub_axi_awaddr
		[6]), .Z(n_1361068));
	notech_nand2 i_52006(.A(i_psram_sub_axi_awaddr[6]), .B(i_psram_sub_axi_awaddr
		[7]), .Z(n_1371067));
	notech_nand2 i_62005(.A(i_psram_sub_axi_awaddr[7]), .B(i_psram_sub_axi_awaddr
		[8]), .Z(n_1381066));
	notech_nand2 i_72004(.A(i_psram_sub_axi_awaddr[8]), .B(i_psram_sub_axi_awaddr
		[9]), .Z(n_1391065));
	notech_nand2 i_82003(.A(i_psram_sub_axi_awaddr[9]), .B(i_psram_sub_axi_awaddr
		[10]), .Z(n_1401064));
	notech_nand2 i_92002(.A(i_psram_sub_axi_awaddr[10]), .B(i_psram_sub_axi_awaddr
		[11]), .Z(n_1411063));
	notech_nand2 i_102001(.A(i_psram_sub_axi_awaddr[11]), .B(i_psram_sub_axi_awaddr
		[12]), .Z(n_1421062));
	notech_nand2 i_112000(.A(i_psram_sub_axi_awaddr[12]), .B(i_psram_sub_axi_awaddr
		[13]), .Z(n_1431061));
	notech_nand2 i_121999(.A(i_psram_sub_axi_awaddr[13]), .B(i_psram_sub_axi_awaddr
		[14]), .Z(n_1441060));
	notech_nand2 i_131998(.A(i_psram_sub_axi_awaddr[14]), .B(i_psram_sub_axi_awaddr
		[15]), .Z(n_1451059));
	notech_nand2 i_141997(.A(i_psram_sub_axi_awaddr[15]), .B(i_psram_sub_axi_awaddr
		[16]), .Z(n_1461058));
	notech_nand2 i_151996(.A(i_psram_sub_axi_awaddr[16]), .B(i_psram_sub_axi_awaddr
		[17]), .Z(n_1471057));
	notech_nand2 i_161995(.A(i_psram_sub_axi_awaddr[17]), .B(i_psram_sub_axi_awaddr
		[18]), .Z(n_1481056));
	notech_nand2 i_171994(.A(i_psram_sub_axi_awaddr[18]), .B(i_psram_sub_axi_awaddr
		[19]), .Z(n_1491055));
	notech_nand2 i_181993(.A(i_psram_sub_axi_awaddr[19]), .B(i_psram_sub_axi_awaddr
		[20]), .Z(n_1501054));
	notech_nand2 i_191992(.A(i_psram_sub_axi_awaddr[20]), .B(i_psram_sub_axi_awaddr
		[21]), .Z(n_1511053));
	notech_nand2 i_201991(.A(i_psram_sub_axi_awaddr[21]), .B(i_psram_sub_axi_awaddr
		[22]), .Z(n_1521052));
	notech_inv i_221990(.A(\i_psram_sub_axi_awaddr_0[2] ), .Z(n_1541051));
	notech_inv i_231989(.A(n_1331071), .Z(n_2651050));
	notech_nor2 i_241988(.A(\i_psram_sub_axi_awaddr_0[2] ), .B(n_1341070), .Z
		(n_1561049));
	notech_nor2 i_251987(.A(n_1331071), .B(n_1351069), .Z(n_1571048));
	notech_nor2 i_261986(.A(n_1341070), .B(n_1361068), .Z(n_1581047));
	notech_nor2 i_271985(.A(n_1351069), .B(n_1371067), .Z(n_1591046));
	notech_nor2 i_281984(.A(n_1361068), .B(n_1381066), .Z(n_1601045));
	notech_nor2 i_291983(.A(n_1371067), .B(n_1391065), .Z(n_1611044));
	notech_nor2 i_301982(.A(n_1381066), .B(n_1401064), .Z(n_1621043));
	notech_nor2 i_311981(.A(n_1391065), .B(n_1411063), .Z(n_1631042));
	notech_nor2 i_321980(.A(n_1401064), .B(n_1421062), .Z(n_1641041));
	notech_nor2 i_331979(.A(n_1411063), .B(n_1431061), .Z(n_1651040));
	notech_nor2 i_341978(.A(n_1421062), .B(n_1441060), .Z(n_1661039));
	notech_nor2 i_351977(.A(n_1431061), .B(n_1451059), .Z(n_1671038));
	notech_nor2 i_361976(.A(n_1441060), .B(n_1461058), .Z(n_1681037));
	notech_nor2 i_371975(.A(n_1451059), .B(n_1471057), .Z(n_1691036));
	notech_nor2 i_381974(.A(n_1461058), .B(n_1481056), .Z(n_1701035));
	notech_nor2 i_391973(.A(n_1471057), .B(n_1491055), .Z(n_1711034));
	notech_nor2 i_401972(.A(n_1481056), .B(n_1501054), .Z(n_1721033));
	notech_nor2 i_411971(.A(n_1491055), .B(n_1511053), .Z(n_1731032));
	notech_nor2 i_421970(.A(n_1501054), .B(n_1521052), .Z(n_1741031));
	notech_inv i_441969(.A(n_1541051), .Z(n_1761030));
	notech_inv i_451968(.A(n_2651050), .Z(n_1771029));
	notech_inv i_461967(.A(n_1561049), .Z(n_1781028));
	notech_inv i_471966(.A(n_1571048), .Z(n_2661027));
	notech_nand2 i_481965(.A(n_1541051), .B(n_1581047), .Z(n_1801026));
	notech_nand2 i_491964(.A(n_2651050), .B(n_1591046), .Z(n_1811025));
	notech_nand2 i_501963(.A(n_1561049), .B(n_1601045), .Z(n_1821024));
	notech_nand2 i_511962(.A(n_1571048), .B(n_1611044), .Z(n_1831023));
	notech_nand2 i_521961(.A(n_1581047), .B(n_1621043), .Z(n_1841022));
	notech_nand2 i_531960(.A(n_1591046), .B(n_1631042), .Z(n_1851021));
	notech_nand2 i_541959(.A(n_1601045), .B(n_1641041), .Z(n_1861020));
	notech_nand2 i_551958(.A(n_1611044), .B(n_1651040), .Z(n_1871019));
	notech_nand2 i_561957(.A(n_1621043), .B(n_1661039), .Z(n_1881018));
	notech_nand2 i_571956(.A(n_1631042), .B(n_1671038), .Z(n_1891017));
	notech_nand2 i_581955(.A(n_1641041), .B(n_1681037), .Z(n_1901016));
	notech_nand2 i_591954(.A(n_1651040), .B(n_1691036), .Z(n_1911015));
	notech_nand2 i_601953(.A(n_1661039), .B(n_1701035), .Z(n_1921014));
	notech_nand2 i_611952(.A(n_1671038), .B(n_1711034), .Z(n_1931013));
	notech_nand2 i_621951(.A(n_1681037), .B(n_1721033), .Z(n_1941012));
	notech_nand2 i_631950(.A(n_1691036), .B(n_1731032), .Z(n_1951011));
	notech_nand2 i_641949(.A(n_1701035), .B(n_1741031), .Z(n_1961010));
	notech_inv i_661948(.A(n_1761030), .Z(n_1981009));
	notech_inv i_671947(.A(n_1771029), .Z(n_1991008));
	notech_inv i_681946(.A(n_1781028), .Z(n_2001007));
	notech_inv i_691945(.A(n_2661027), .Z(n_2011006));
	notech_inv i_701944(.A(n_1801026), .Z(n_2021005));
	notech_nor2 i_741943(.A(n_1761030), .B(n_1841022), .Z(n_2061004));
	notech_nor2 i_751942(.A(n_1771029), .B(n_1851021), .Z(n_2071003));
	notech_nor2 i_761941(.A(n_1781028), .B(n_1861020), .Z(n_2081002));
	notech_nor2 i_771940(.A(n_2661027), .B(n_1871019), .Z(n_2091001));
	notech_nor2 i_781939(.A(n_1801026), .B(n_1881018), .Z(n_2101000));
	notech_nor2 i_791938(.A(n_1811025), .B(n_1891017), .Z(n_211999));
	notech_nor2 i_801937(.A(n_1821024), .B(n_1901016), .Z(n_212998));
	notech_nor2 i_811936(.A(n_1831023), .B(n_1911015), .Z(n_213997));
	notech_nor2 i_821935(.A(n_1841022), .B(n_1921014), .Z(n_214996));
	notech_nor2 i_831934(.A(n_1851021), .B(n_1931013), .Z(n_215995));
	notech_nor2 i_841933(.A(n_1861020), .B(n_1941012), .Z(n_216994));
	notech_nor2 i_851932(.A(n_1871019), .B(n_1951011), .Z(n_217993));
	notech_nor2 i_861931(.A(n_1881018), .B(n_1961010), .Z(n_218992));
	notech_inv i_881930(.A(n_1981009), .Z(n_220991));
	notech_inv i_891929(.A(n_1991008), .Z(n_221990));
	notech_inv i_901928(.A(n_2001007), .Z(n_222989));
	notech_inv i_911927(.A(n_2011006), .Z(n_223988));
	notech_inv i_921926(.A(n_2021005), .Z(n_224987));
	notech_inv i_961925(.A(n_2061004), .Z(n_228986));
	notech_inv i_971924(.A(n_2071003), .Z(n_229985));
	notech_inv i_981923(.A(n_2081002), .Z(n_230984));
	notech_inv i_991922(.A(n_2091001), .Z(n_231983));
	notech_inv i_1001921(.A(n_2101000), .Z(n_232982));
	notech_inv i_1011920(.A(n_211999), .Z(n_233981));
	notech_inv i_1021919(.A(n_212998), .Z(n_234980));
	notech_inv i_1031918(.A(n_213997), .Z(n_272979));
	notech_nand2 i_1041917(.A(n_1981009), .B(n_214996), .Z(n_236978));
	notech_nand2 i_1051916(.A(n_1991008), .B(n_215995), .Z(n_237977));
	notech_nand2 i_1061915(.A(n_2001007), .B(n_216994), .Z(n_238976));
	notech_nand2 i_1071914(.A(n_2011006), .B(n_217993), .Z(n_239975));
	notech_nand2 i_1081913(.A(n_2021005), .B(n_218992), .Z(n_240974));
	notech_inv i_1321912(.A(n_220991), .Z(n_276973));
	notech_inv i_1331911(.A(i_psram_sub_axi_awaddr[3]), .Z(n_279972));
	notech_nand2 i_1341910(.A(n_279972), .B(n_220991), .Z(n_280971));
	notech_nand2 i_1351909(.A(i_psram_sub_axi_awaddr[3]), .B(n_276973), .Z(n_277970
		));
	notech_nand2 i_1361908(.A(n_277970), .B(n_280971), .Z(n_278969));
	notech_inv i_1371907(.A(n_278969), .Z(\i_psram_sub_axi_awaddr_0[3] ));
	notech_inv i_1381906(.A(n_221990), .Z(n_281968));
	notech_inv i_1391905(.A(i_psram_sub_axi_awaddr[4]), .Z(n_284967));
	notech_nand2 i_1401904(.A(n_284967), .B(n_221990), .Z(n_285966));
	notech_nand2 i_1411903(.A(i_psram_sub_axi_awaddr[4]), .B(n_281968), .Z(n_282965
		));
	notech_nand2 i_1421902(.A(n_282965), .B(n_285966), .Z(n_283964));
	notech_inv i_1431901(.A(n_283964), .Z(\i_psram_sub_axi_awaddr_0[4] ));
	notech_inv i_1441900(.A(n_222989), .Z(n_286963));
	notech_inv i_1451899(.A(i_psram_sub_axi_awaddr[5]), .Z(n_289962));
	notech_nand2 i_1461898(.A(n_289962), .B(n_222989), .Z(n_290961));
	notech_nand2 i_1471897(.A(i_psram_sub_axi_awaddr[5]), .B(n_286963), .Z(n_287960
		));
	notech_nand2 i_1481896(.A(n_287960), .B(n_290961), .Z(n_288959));
	notech_inv i_1491895(.A(n_288959), .Z(\i_psram_sub_axi_awaddr_0[5] ));
	notech_inv i_1501894(.A(n_223988), .Z(n_291958));
	notech_inv i_1511893(.A(i_psram_sub_axi_awaddr[6]), .Z(n_294957));
	notech_nand2 i_1521892(.A(n_294957), .B(n_223988), .Z(n_295956));
	notech_nand2 i_1531891(.A(i_psram_sub_axi_awaddr[6]), .B(n_291958), .Z(n_292955
		));
	notech_nand2 i_1541890(.A(n_292955), .B(n_295956), .Z(n_293954));
	notech_inv i_1551889(.A(n_293954), .Z(\i_psram_sub_axi_awaddr_0[6] ));
	notech_inv i_1561888(.A(n_224987), .Z(n_296953));
	notech_inv i_1571887(.A(i_psram_sub_axi_awaddr[7]), .Z(n_299952));
	notech_nand2 i_1581886(.A(n_299952), .B(n_224987), .Z(n_300951));
	notech_nand2 i_1591885(.A(i_psram_sub_axi_awaddr[7]), .B(n_296953), .Z(n_297950
		));
	notech_nand2 i_1601884(.A(n_297950), .B(n_300951), .Z(n_298949));
	notech_inv i_1611883(.A(n_298949), .Z(\i_psram_sub_axi_awaddr_0[7] ));
	notech_inv i_1621882(.A(n_1811025), .Z(n_301948));
	notech_inv i_1631881(.A(i_psram_sub_axi_awaddr[8]), .Z(n_304947));
	notech_nand2 i_1641880(.A(n_304947), .B(n_1811025), .Z(n_305946));
	notech_nand2 i_1651879(.A(i_psram_sub_axi_awaddr[8]), .B(n_301948), .Z(n_302945
		));
	notech_nand2 i_1661878(.A(n_302945), .B(n_305946), .Z(n_303944));
	notech_inv i_1671877(.A(n_303944), .Z(\i_psram_sub_axi_awaddr_0[8] ));
	notech_inv i_1681876(.A(n_1821024), .Z(n_306943));
	notech_inv i_1691875(.A(i_psram_sub_axi_awaddr[9]), .Z(n_309942));
	notech_nand2 i_1701874(.A(n_309942), .B(n_1821024), .Z(n_310941));
	notech_nand2 i_1711873(.A(i_psram_sub_axi_awaddr[9]), .B(n_306943), .Z(n_307940
		));
	notech_nand2 i_1721872(.A(n_307940), .B(n_310941), .Z(n_308939));
	notech_inv i_1731871(.A(n_308939), .Z(\i_psram_sub_axi_awaddr_0[9] ));
	notech_inv i_1741870(.A(n_1831023), .Z(n_311938));
	notech_inv i_1751869(.A(i_psram_sub_axi_awaddr[10]), .Z(n_314937));
	notech_nand2 i_1761868(.A(n_314937), .B(n_1831023), .Z(n_315936));
	notech_nand2 i_1771867(.A(i_psram_sub_axi_awaddr[10]), .B(n_311938), .Z(n_312935
		));
	notech_nand2 i_1781866(.A(n_312935), .B(n_315936), .Z(n_313934));
	notech_inv i_1791865(.A(n_313934), .Z(\i_psram_sub_axi_awaddr_0[10] ));
	notech_inv i_1801864(.A(n_228986), .Z(n_316933));
	notech_inv i_1811863(.A(i_psram_sub_axi_awaddr[11]), .Z(n_319932));
	notech_nand2 i_1821862(.A(n_319932), .B(n_228986), .Z(n_320931));
	notech_nand2 i_1831861(.A(i_psram_sub_axi_awaddr[11]), .B(n_316933), .Z(n_317930
		));
	notech_nand2 i_1841860(.A(n_317930), .B(n_320931), .Z(n_318929));
	notech_inv i_1851859(.A(n_318929), .Z(\i_psram_sub_axi_awaddr_0[11] ));
	notech_inv i_1861858(.A(n_229985), .Z(n_321928));
	notech_inv i_1871857(.A(i_psram_sub_axi_awaddr[12]), .Z(n_324927));
	notech_nand2 i_1881856(.A(n_324927), .B(n_229985), .Z(n_325926));
	notech_nand2 i_1891855(.A(i_psram_sub_axi_awaddr[12]), .B(n_321928), .Z(n_322925
		));
	notech_nand2 i_1901854(.A(n_322925), .B(n_325926), .Z(n_323924));
	notech_inv i_1911853(.A(n_323924), .Z(\i_psram_sub_axi_awaddr_0[12] ));
	notech_inv i_1921852(.A(n_230984), .Z(n_326923));
	notech_inv i_1931851(.A(i_psram_sub_axi_awaddr[13]), .Z(n_329922));
	notech_nand2 i_1941850(.A(n_329922), .B(n_230984), .Z(n_330921));
	notech_nand2 i_1951849(.A(i_psram_sub_axi_awaddr[13]), .B(n_326923), .Z(n_327920
		));
	notech_nand2 i_1961848(.A(n_327920), .B(n_330921), .Z(n_328919));
	notech_inv i_1971847(.A(n_328919), .Z(\i_psram_sub_axi_awaddr_0[13] ));
	notech_inv i_1981846(.A(n_231983), .Z(n_331918));
	notech_inv i_1991845(.A(i_psram_sub_axi_awaddr[14]), .Z(n_334917));
	notech_nand2 i_2001844(.A(n_334917), .B(n_231983), .Z(n_335916));
	notech_nand2 i_2011843(.A(i_psram_sub_axi_awaddr[14]), .B(n_331918), .Z(n_332915
		));
	notech_nand2 i_2021842(.A(n_332915), .B(n_335916), .Z(n_333914));
	notech_inv i_2031841(.A(n_333914), .Z(\i_psram_sub_axi_awaddr_0[14] ));
	notech_inv i_2041840(.A(n_232982), .Z(n_336913));
	notech_inv i_2051839(.A(i_psram_sub_axi_awaddr[15]), .Z(n_339912));
	notech_nand2 i_2061838(.A(n_339912), .B(n_232982), .Z(n_340911));
	notech_nand2 i_2071837(.A(i_psram_sub_axi_awaddr[15]), .B(n_336913), .Z(n_337910
		));
	notech_nand2 i_2081836(.A(n_337910), .B(n_340911), .Z(n_338909));
	notech_inv i_2091835(.A(n_338909), .Z(\i_psram_sub_axi_awaddr_0[15] ));
	notech_inv i_2101834(.A(n_233981), .Z(n_341908));
	notech_inv i_2111833(.A(i_psram_sub_axi_awaddr[16]), .Z(n_344907));
	notech_nand2 i_2121832(.A(n_344907), .B(n_233981), .Z(n_345906));
	notech_nand2 i_2131831(.A(i_psram_sub_axi_awaddr[16]), .B(n_341908), .Z(n_342905
		));
	notech_nand2 i_2141830(.A(n_342905), .B(n_345906), .Z(n_343904));
	notech_inv i_2151829(.A(n_343904), .Z(\i_psram_sub_axi_awaddr_0[16] ));
	notech_inv i_2161828(.A(n_234980), .Z(n_346903));
	notech_inv i_2171827(.A(i_psram_sub_axi_awaddr[17]), .Z(n_349902));
	notech_nand2 i_2181826(.A(n_349902), .B(n_234980), .Z(n_350901));
	notech_nand2 i_2191825(.A(i_psram_sub_axi_awaddr[17]), .B(n_346903), .Z(n_347900
		));
	notech_nand2 i_2201824(.A(n_347900), .B(n_350901), .Z(n_348899));
	notech_inv i_2211823(.A(n_348899), .Z(\i_psram_sub_axi_awaddr_0[17] ));
	notech_inv i_2221822(.A(n_272979), .Z(n_351898));
	notech_inv i_2231821(.A(i_psram_sub_axi_awaddr[18]), .Z(n_354897));
	notech_nand2 i_2241820(.A(n_354897), .B(n_272979), .Z(n_355896));
	notech_nand2 i_2251819(.A(i_psram_sub_axi_awaddr[18]), .B(n_351898), .Z(n_352895
		));
	notech_nand2 i_2261818(.A(n_352895), .B(n_355896), .Z(n_353894));
	notech_inv i_2271817(.A(n_353894), .Z(\i_psram_sub_axi_awaddr_0[18] ));
	notech_inv i_2281816(.A(n_236978), .Z(n_356893));
	notech_inv i_2291815(.A(i_psram_sub_axi_awaddr[19]), .Z(n_359892));
	notech_nand2 i_2301814(.A(n_359892), .B(n_236978), .Z(n_360891));
	notech_nand2 i_2311813(.A(i_psram_sub_axi_awaddr[19]), .B(n_356893), .Z(n_357890
		));
	notech_nand2 i_2321812(.A(n_357890), .B(n_360891), .Z(n_358889));
	notech_inv i_2331811(.A(n_358889), .Z(\i_psram_sub_axi_awaddr_0[19] ));
	notech_inv i_2341810(.A(n_237977), .Z(n_361888));
	notech_inv i_2351809(.A(i_psram_sub_axi_awaddr[20]), .Z(n_364887));
	notech_nand2 i_2361808(.A(n_364887), .B(n_237977), .Z(n_365886));
	notech_nand2 i_2371807(.A(i_psram_sub_axi_awaddr[20]), .B(n_361888), .Z(n_362885
		));
	notech_nand2 i_2381806(.A(n_362885), .B(n_365886), .Z(n_363884));
	notech_inv i_2391805(.A(n_363884), .Z(\i_psram_sub_axi_awaddr_0[20] ));
	notech_inv i_2401804(.A(n_238976), .Z(n_366883));
	notech_inv i_2411803(.A(i_psram_sub_axi_awaddr[21]), .Z(n_369882));
	notech_nand2 i_2421802(.A(n_369882), .B(n_238976), .Z(n_370881));
	notech_nand2 i_2431801(.A(i_psram_sub_axi_awaddr[21]), .B(n_366883), .Z(n_367880
		));
	notech_nand2 i_2441800(.A(n_367880), .B(n_370881), .Z(n_368879));
	notech_inv i_2451799(.A(n_368879), .Z(\i_psram_sub_axi_awaddr_0[21] ));
	notech_inv i_2461798(.A(n_239975), .Z(n_371878));
	notech_inv i_2471797(.A(i_psram_sub_axi_awaddr[22]), .Z(n_374877));
	notech_nand2 i_2481796(.A(n_374877), .B(n_239975), .Z(n_375876));
	notech_nand2 i_2491795(.A(i_psram_sub_axi_awaddr[22]), .B(n_371878), .Z(n_372875
		));
	notech_nand2 i_2501794(.A(n_372875), .B(n_375876), .Z(n_373874));
	notech_inv i_2511793(.A(n_373874), .Z(\i_psram_sub_axi_awaddr_0[22] ));
	notech_inv i_2521792(.A(n_240974), .Z(n_376873));
	notech_inv i_2531791(.A(i_psram_sub_axi_awaddr[23]), .Z(n_379872));
	notech_nand2 i_2541790(.A(n_379872), .B(n_240974), .Z(n_380871));
	notech_nand2 i_2551789(.A(i_psram_sub_axi_awaddr[23]), .B(n_376873), .Z(n_377870
		));
	notech_nand2 i_2561788(.A(n_377870), .B(n_380871), .Z(n_378869));
	notech_inv i_2571787(.A(n_378869), .Z(\i_psram_sub_axi_awaddr_0[23] ));
	notech_inv i_121786(.A(n_249), .Z(n_371801));
	notech_inv i_171785(.A(n_418), .Z(n_469));
	notech_inv i_491784(.A(n_242), .Z(n_363809));
	notech_inv i_591656(.A(n_242), .Z(n_625));
	notech_inv i_591783(.A(i_psram_sub_axi_araddr[1]), .Z(n_265862));
	notech_inv i_601782(.A(i_psram_sub_axi_araddr[10]), .Z(n_274));
	notech_inv i_611655(.A(n_642), .Z(n_690));
	notech_inv i_611781(.A(i_psram_sub_axi_araddr[11]), .Z(n_275));
	notech_inv i_621654(.A(i_psram_sub_axi_araddr[11]), .Z(n_602));
	notech_inv i_621780(.A(i_psram_sub_axi_araddr[12]), .Z(n_276859));
	notech_inv i_631653(.A(n_601), .Z(n_649));
	notech_inv i_631779(.A(i_psram_sub_axi_araddr[13]), .Z(n_277858));
	notech_inv i_641652(.A(i_psram_sub_axi_araddr[13]), .Z(n_606));
	notech_inv i_641778(.A(i_psram_sub_axi_araddr[14]), .Z(n_278857));
	notech_inv i_651651(.A(n_689), .Z(n_737));
	notech_inv i_65(.A(i_psram_sub_axi_araddr[15]), .Z(n_279856));
	notech_inv i_661650(.A(i_psram_sub_axi_araddr[15]), .Z(n_610));
	notech_inv i_661777(.A(i_psram_sub_axi_araddr[16]), .Z(n_280855));
	notech_inv i_671649(.A(n_609), .Z(n_657));
	notech_inv i_671776(.A(i_psram_sub_axi_araddr[17]), .Z(n_281854));
	notech_inv i_681648(.A(i_psram_sub_axi_araddr[17]), .Z(n_614));
	notech_inv i_681775(.A(i_psram_sub_axi_araddr[18]), .Z(n_282853));
	notech_inv i_691647(.A(n_658), .Z(n_706));
	notech_inv i_691774(.A(i_psram_sub_axi_araddr[19]), .Z(n_283852));
	notech_inv i_701646(.A(i_psram_sub_axi_araddr[19]), .Z(n_618));
	notech_inv i_701773(.A(i_psram_sub_axi_araddr[20]), .Z(n_284851));
	notech_inv i_711645(.A(n_617), .Z(n_665));
	notech_inv i_711644(.A(i_psram_sub_axi_araddr[21]), .Z(n_285850));
	notech_inv i_741643(.A(i_psram_sub_axi_araddr[21]), .Z(n_622));
	notech_inv i_741642(.A(i_psram_sub_axi_araddr[22]), .Z(n_286849));
	notech_inv i_741641(.A(n_417), .Z(n_468));
	notech_inv i_761640(.A(n_640), .Z(n_688));
	notech_inv i_761639(.A(i_psram_sub_axi_araddr[10]), .Z(n_600));
	notech_inv i_761638(.A(n_599), .Z(n_647));
	notech_inv i_761637(.A(i_psram_sub_axi_araddr[12]), .Z(n_604));
	notech_inv i_761636(.A(n_687), .Z(n_735));
	notech_inv i_761635(.A(i_psram_sub_axi_araddr[14]), .Z(n_608));
	notech_inv i_761634(.A(n_607), .Z(n_655));
	notech_inv i_761633(.A(i_psram_sub_axi_araddr[16]), .Z(n_612));
	notech_inv i_761632(.A(n_656), .Z(n_704));
	notech_inv i_761631(.A(i_psram_sub_axi_araddr[18]), .Z(n_616));
	notech_inv i_761630(.A(n_615), .Z(n_663));
	notech_inv i_761629(.A(i_psram_sub_axi_araddr[20]), .Z(n_620));
	notech_inv i_741628(.A(n_467), .Z(n_522));
	notech_inv i_761627(.A(n_597), .Z(n_645));
	notech_inv i_761626(.A(n_685), .Z(n_733));
	notech_inv i_761625(.A(n_605), .Z(n_653));
	notech_inv i_761624(.A(n_654), .Z(n_702));
	notech_inv i_761623(.A(n_613), .Z(n_661));
	notech_inv i_741622(.A(n_370802), .Z(n_419));
	notech_inv i_741621(.A(n_466), .Z(n_521));
	notech_inv i_741620(.A(n_364808), .Z(n_411));
	notech_inv i_761619(.A(n_595), .Z(n_643));
	notech_inv i_761618(.A(n_683), .Z(n_731));
	notech_inv i_761617(.A(n_603), .Z(n_651));
	notech_inv i_761616(.A(n_652), .Z(n_700));
	notech_inv i_761615(.A(n_611), .Z(n_659));
	notech_inv i_741614(.A(n_465), .Z(n_520));
	notech_inv i_761613(.A(n_681), .Z(n_729));
	notech_inv i_761612(.A(n_650), .Z(n_698));
	notech_inv i_761611(.A(n_464), .Z(n_744));
	notech_inv i_761610(.A(n_679), .Z(n_727));
	notech_inv i_761609(.A(n_648), .Z(n_696));
	notech_inv i_741608(.A(n_249), .Z(n_471));
	notech_inv i_761607(.A(n_646), .Z(n_694));
	notech_inv i_761772(.A(n_644), .Z(n_692));
	notech_inv i_741606(.A(n_294846), .Z(n_767));
	notech_inv i_741771(.A(i_psram_sub_axi_araddr[1]), .Z(n_762));
	notech_inv i_741605(.A(i_psram_sub_axi_araddr[0]), .Z(n_757));
	notech_inv i_21770(.A(s00_axi_arlen[0]), .Z(n_218868));
	notech_inv i_31769(.A(s00_axi_arlen[1]), .Z(n_219));
	notech_inv i_41768(.A(s00_axi_arlen[2]), .Z(n_220867));
	notech_inv i_51767(.A(s00_axi_arlen[3]), .Z(n_221866));
	notech_inv i_61766(.A(s00_axi_arlen[4]), .Z(n_222865));
	notech_inv i_71765(.A(s00_axi_arlen[5]), .Z(n_223864));
	notech_inv i_81764(.A(s00_axi_arlen[6]), .Z(n_224863));
	notech_inv i_91763(.A(s00_axi_arlen[7]), .Z(n_225));
	notech_nor2 i_261762(.A(i_psram_sub_axi_araddr[2]), .B(n_218868), .Z(n_242
		));
	notech_nor2 i_271761(.A(i_psram_sub_axi_araddr[3]), .B(n_219), .Z(n_243)
		);
	notech_nor2 i_281760(.A(i_psram_sub_axi_araddr[4]), .B(n_220867), .Z(n_244
		));
	notech_nor2 i_291759(.A(i_psram_sub_axi_araddr[5]), .B(n_221866), .Z(n_245
		));
	notech_nor2 i_301758(.A(i_psram_sub_axi_araddr[6]), .B(n_222865), .Z(n_246
		));
	notech_nor2 i_311757(.A(i_psram_sub_axi_araddr[7]), .B(n_223864), .Z(n_247
		));
	notech_nor2 i_321756(.A(i_psram_sub_axi_araddr[8]), .B(n_224863), .Z(n_248
		));
	notech_nor2 i_331755(.A(i_psram_sub_axi_araddr[9]), .B(n_225), .Z(n_249)
		);
	notech_nand2 i_501754(.A(i_psram_sub_axi_araddr[2]), .B(n_218868), .Z(n_266861
		));
	notech_nand2 i_511753(.A(i_psram_sub_axi_araddr[3]), .B(n_219), .Z(n_267
		));
	notech_nand2 i_521752(.A(i_psram_sub_axi_araddr[4]), .B(n_220867), .Z(n_268
		));
	notech_nand2 i_531751(.A(i_psram_sub_axi_araddr[5]), .B(n_221866), .Z(n_269
		));
	notech_nand2 i_541750(.A(i_psram_sub_axi_araddr[6]), .B(n_222865), .Z(n_270
		));
	notech_nand2 i_551749(.A(i_psram_sub_axi_araddr[7]), .B(n_223864), .Z(n_271
		));
	notech_nand2 i_561748(.A(i_psram_sub_axi_araddr[8]), .B(n_224863), .Z(n_272860
		));
	notech_nand2 i_571747(.A(i_psram_sub_axi_araddr[9]), .B(n_225), .Z(n_273
		));
	notech_inv i_72(.A(i_psram_sub_axi_araddr[0]), .Z(n_288848));
	notech_inv i_771746(.A(n_242), .Z(n_293847));
	notech_nand2 i_781745(.A(n_293847), .B(n_266861), .Z(n_294846));
	notech_inv i_791744(.A(n_243), .Z(n_295845));
	notech_nand2 i_801743(.A(n_295845), .B(n_267), .Z(n_296844));
	notech_inv i_811742(.A(n_244), .Z(n_297843));
	notech_nand2 i_821741(.A(n_297843), .B(n_268), .Z(n_298842));
	notech_inv i_831740(.A(n_245), .Z(n_299841));
	notech_nand2 i_841739(.A(n_299841), .B(n_269), .Z(n_300840));
	notech_inv i_851738(.A(n_246), .Z(n_301839));
	notech_nand2 i_861737(.A(n_301839), .B(n_270), .Z(n_302838));
	notech_inv i_87(.A(n_247), .Z(n_303837));
	notech_nand2 i_881736(.A(n_303837), .B(n_271), .Z(n_304836));
	notech_inv i_891735(.A(n_248), .Z(n_305835));
	notech_nand2 i_901734(.A(n_305835), .B(n_272860), .Z(n_306834));
	notech_inv i_911733(.A(n_249), .Z(n_307833));
	notech_nand2 i_921732(.A(n_307833), .B(n_273), .Z(n_308832));
	notech_or2 i_360(.A(n_242), .B(n_265862), .Z(n_582));
	notech_and2 i_361(.A(n_582), .B(n_266861), .Z(n_581));
	notech_inv i_362(.A(n_581), .Z(n_339831));
	notech_or2 i_363(.A(n_243), .B(n_266861), .Z(n_584));
	notech_and2 i_364(.A(n_584), .B(n_267), .Z(n_583));
	notech_inv i_365(.A(n_583), .Z(n_340830));
	notech_or2 i_366(.A(n_244), .B(n_267), .Z(n_586));
	notech_and2 i_367(.A(n_586), .B(n_268), .Z(n_585));
	notech_inv i_368(.A(n_585), .Z(n_341829));
	notech_or2 i_369(.A(n_245), .B(n_268), .Z(n_588));
	notech_and2 i_370(.A(n_588), .B(n_269), .Z(n_587));
	notech_inv i_371(.A(n_587), .Z(n_342828));
	notech_or2 i_372(.A(n_246), .B(n_269), .Z(n_590));
	notech_and2 i_373(.A(n_590), .B(n_270), .Z(n_589));
	notech_inv i_374(.A(n_589), .Z(n_343827));
	notech_or2 i_375(.A(n_247), .B(n_270), .Z(n_592));
	notech_and2 i_376(.A(n_592), .B(n_271), .Z(n_591));
	notech_inv i_377(.A(n_591), .Z(n_344826));
	notech_or2 i_378(.A(n_248), .B(n_271), .Z(n_594));
	notech_and2 i_379(.A(n_594), .B(n_272860), .Z(n_593));
	notech_inv i_380(.A(n_593), .Z(n_345825));
	notech_or2 i_381(.A(n_249), .B(n_272860), .Z(n_596));
	notech_and2 i_382(.A(n_596), .B(n_273), .Z(n_595));
	notech_inv i_383(.A(n_595), .Z(n_346824));
	notech_and2 i_385(.A(n_273), .B(n_274), .Z(n_597));
	notech_inv i_386(.A(n_597), .Z(n_347823));
	notech_and2 i_388(.A(n_600), .B(n_275), .Z(n_599));
	notech_inv i_389(.A(n_599), .Z(n_348822));
	notech_and2 i_391(.A(n_602), .B(n_276859), .Z(n_601));
	notech_inv i_392(.A(n_601), .Z(n_349821));
	notech_and2 i_394(.A(n_604), .B(n_277858), .Z(n_603));
	notech_inv i_395(.A(n_603), .Z(n_350820));
	notech_and2 i_397(.A(n_606), .B(n_278857), .Z(n_605));
	notech_inv i_398(.A(n_605), .Z(n_351819));
	notech_and2 i_400(.A(n_608), .B(n_279856), .Z(n_607));
	notech_inv i_401(.A(n_607), .Z(n_352818));
	notech_and2 i_403(.A(n_610), .B(n_280855), .Z(n_609));
	notech_inv i_404(.A(n_609), .Z(n_353817));
	notech_and2 i_406(.A(n_612), .B(n_281854), .Z(n_611));
	notech_inv i_407(.A(n_611), .Z(n_354816));
	notech_and2 i_409(.A(n_614), .B(n_282853), .Z(n_613));
	notech_inv i_410(.A(n_613), .Z(n_355815));
	notech_and2 i_412(.A(n_616), .B(n_283852), .Z(n_615));
	notech_inv i_413(.A(n_615), .Z(n_356814));
	notech_and2 i_415(.A(n_618), .B(n_284851), .Z(n_617));
	notech_inv i_416(.A(n_617), .Z(n_357813));
	notech_and2 i_418(.A(n_620), .B(n_285850), .Z(n_619));
	notech_inv i_419(.A(n_619), .Z(n_358812));
	notech_and2 i_421(.A(n_622), .B(n_286849), .Z(n_621));
	notech_inv i_422(.A(n_621), .Z(n_359811));
	notech_inv i_1441731(.A(n_288848), .Z(n_360810));
	notech_nor2 i_1481730(.A(n_242), .B(n_243), .Z(n_364808));
	notech_nor2 i_1491729(.A(n_243), .B(n_244), .Z(n_365807));
	notech_nor2 i_1501728(.A(n_244), .B(n_245), .Z(n_366806));
	notech_nor2 i_1511727(.A(n_245), .B(n_246), .Z(n_367805));
	notech_nor2 i_1521726(.A(n_246), .B(n_247), .Z(n_368804));
	notech_nor2 i_1531725(.A(n_247), .B(n_248), .Z(n_369803));
	notech_nor2 i_1541724(.A(n_248), .B(n_249), .Z(n_370802));
	notech_or2 i_427(.A(n_625), .B(n_339831), .Z(n_626));
	notech_inv i_428(.A(n_626), .Z(n_386));
	notech_or2 i_430(.A(n_364808), .B(n_340830), .Z(n_628));
	notech_inv i_431(.A(n_628), .Z(n_387));
	notech_and2 i_432(.A(n_365807), .B(n_339831), .Z(n_629));
	notech_or2 i_433(.A(n_629), .B(n_341829), .Z(n_630));
	notech_inv i_434(.A(n_630), .Z(n_388));
	notech_and2 i_435(.A(n_366806), .B(n_340830), .Z(n_631));
	notech_or2 i_436(.A(n_631), .B(n_342828), .Z(n_632));
	notech_inv i_437(.A(n_632), .Z(n_389));
	notech_and2 i_438(.A(n_367805), .B(n_341829), .Z(n_633));
	notech_or2 i_439(.A(n_633), .B(n_343827), .Z(n_634));
	notech_inv i_440(.A(n_634), .Z(n_390));
	notech_and2 i_441(.A(n_368804), .B(n_342828), .Z(n_635));
	notech_or2 i_442(.A(n_635), .B(n_344826), .Z(n_636));
	notech_inv i_443(.A(n_636), .Z(n_391));
	notech_and2 i_444(.A(n_369803), .B(n_343827), .Z(n_637));
	notech_or2 i_445(.A(n_637), .B(n_345825), .Z(n_638));
	notech_inv i_446(.A(n_638), .Z(n_392));
	notech_and2 i_447(.A(n_370802), .B(n_344826), .Z(n_639));
	notech_or2 i_448(.A(n_639), .B(n_346824), .Z(n_640));
	notech_inv i_449(.A(n_640), .Z(n_393));
	notech_and2 i_450(.A(n_371801), .B(n_345825), .Z(n_641));
	notech_or2 i_451(.A(n_641), .B(n_347823), .Z(n_642));
	notech_inv i_452(.A(n_642), .Z(n_394));
	notech_or2 i_454(.A(n_643), .B(n_348822), .Z(n_644));
	notech_inv i_455(.A(n_644), .Z(n_395));
	notech_or2 i_457(.A(n_645), .B(n_349821), .Z(n_646));
	notech_inv i_458(.A(n_646), .Z(n_396));
	notech_or2 i_460(.A(n_647), .B(n_350820), .Z(n_648));
	notech_inv i_461(.A(n_648), .Z(n_397));
	notech_or2 i_463(.A(n_649), .B(n_351819), .Z(n_650));
	notech_inv i_464(.A(n_650), .Z(n_398));
	notech_or2 i_466(.A(n_651), .B(n_352818), .Z(n_652));
	notech_inv i_467(.A(n_652), .Z(n_399));
	notech_or2 i_469(.A(n_653), .B(n_353817), .Z(n_654));
	notech_inv i_470(.A(n_654), .Z(n_400));
	notech_or2 i_472(.A(n_655), .B(n_354816), .Z(n_656));
	notech_inv i_473(.A(n_656), .Z(n_401));
	notech_or2 i_475(.A(n_657), .B(n_355815), .Z(n_658));
	notech_inv i_476(.A(n_658), .Z(n_402));
	notech_or2 i_478(.A(n_659), .B(n_356814), .Z(n_660));
	notech_inv i_479(.A(n_660), .Z(n_403));
	notech_or2 i_481(.A(n_661), .B(n_357813), .Z(n_662));
	notech_inv i_482(.A(n_662), .Z(n_404));
	notech_or2 i_484(.A(n_663), .B(n_358812), .Z(n_664));
	notech_inv i_485(.A(n_664), .Z(n_405));
	notech_or2 i_487(.A(n_665), .B(n_359811), .Z(n_666));
	notech_inv i_488(.A(n_666), .Z(n_406));
	notech_inv i_1911723(.A(n_360810), .Z(n_407));
	notech_nand2 i_1961722(.A(n_363809), .B(n_365807), .Z(n_412));
	notech_nand2 i_1971721(.A(n_364808), .B(n_366806), .Z(n_413));
	notech_nand2 i_1981720(.A(n_365807), .B(n_367805), .Z(n_414));
	notech_nand2 i_1991719(.A(n_366806), .B(n_368804), .Z(n_415));
	notech_nand2 i_2001718(.A(n_367805), .B(n_369803), .Z(n_416));
	notech_nand2 i_2011717(.A(n_368804), .B(n_370802), .Z(n_417));
	notech_nand2 i_2021716(.A(n_369803), .B(n_371801), .Z(n_418));
	notech_inv i_2171715(.A(n_386), .Z(n_433));
	notech_or2 i_489(.A(n_411), .B(n_407), .Z(n_668));
	notech_and2 i_490(.A(n_668), .B(n_387), .Z(n_667));
	notech_inv i_491(.A(n_667), .Z(n_434));
	notech_and2 i_493(.A(n_412), .B(n_388), .Z(n_669));
	notech_inv i_494(.A(n_669), .Z(n_435));
	notech_and2 i_496(.A(n_413), .B(n_389), .Z(n_671));
	notech_inv i_497(.A(n_671), .Z(n_436));
	notech_or2 i_498(.A(n_414), .B(n_386), .Z(n_674));
	notech_and2 i_499(.A(n_674), .B(n_390), .Z(n_673));
	notech_inv i_500(.A(n_673), .Z(n_437));
	notech_or2 i_501(.A(n_415), .B(n_387), .Z(n_676));
	notech_and2 i_502(.A(n_676), .B(n_391), .Z(n_675));
	notech_inv i_503(.A(n_675), .Z(n_438));
	notech_or2 i_504(.A(n_416), .B(n_388), .Z(n_678));
	notech_and2 i_505(.A(n_678), .B(n_392), .Z(n_677));
	notech_inv i_506(.A(n_677), .Z(n_439));
	notech_or2 i_507(.A(n_417), .B(n_389), .Z(n_680));
	notech_and2 i_508(.A(n_680), .B(n_393), .Z(n_679));
	notech_inv i_509(.A(n_679), .Z(n_440));
	notech_or2 i_510(.A(n_418), .B(n_390), .Z(n_682));
	notech_and2 i_511(.A(n_682), .B(n_394), .Z(n_681));
	notech_inv i_512(.A(n_681), .Z(n_441));
	notech_or2 i_513(.A(n_419), .B(n_391), .Z(n_684));
	notech_and2 i_514(.A(n_684), .B(n_395), .Z(n_683));
	notech_inv i_515(.A(n_683), .Z(n_442));
	notech_or2 i_516(.A(n_249), .B(n_392), .Z(n_686));
	notech_and2 i_517(.A(n_686), .B(n_396), .Z(n_685));
	notech_inv i_518(.A(n_685), .Z(n_443));
	notech_and2 i_520(.A(n_688), .B(n_397), .Z(n_687));
	notech_inv i_521(.A(n_687), .Z(n_444));
	notech_and2 i_523(.A(n_690), .B(n_398), .Z(n_689));
	notech_inv i_524(.A(n_689), .Z(n_445));
	notech_and2 i_526(.A(n_692), .B(n_399), .Z(n_691));
	notech_inv i_527(.A(n_691), .Z(n_446));
	notech_and2 i_529(.A(n_694), .B(n_400), .Z(n_693));
	notech_inv i_530(.A(n_693), .Z(n_447));
	notech_and2 i_532(.A(n_696), .B(n_401), .Z(n_695));
	notech_inv i_533(.A(n_695), .Z(n_448));
	notech_and2 i_535(.A(n_698), .B(n_402), .Z(n_697));
	notech_inv i_536(.A(n_697), .Z(n_449));
	notech_and2 i_538(.A(n_700), .B(n_403), .Z(n_699));
	notech_inv i_539(.A(n_699), .Z(n_450));
	notech_and2 i_541(.A(n_702), .B(n_404), .Z(n_701));
	notech_inv i_542(.A(n_701), .Z(n_451));
	notech_and2 i_544(.A(n_704), .B(n_405), .Z(n_703));
	notech_inv i_545(.A(n_703), .Z(n_452));
	notech_and2 i_547(.A(n_706), .B(n_406), .Z(n_705));
	notech_inv i_548(.A(n_705), .Z(n_453));
	notech_inv i_2381714(.A(n_407), .Z(n_454));
	notech_nor2 i_2461713(.A(n_411), .B(n_415), .Z(n_462));
	notech_nor2 i_2471712(.A(n_412), .B(n_416), .Z(n_463));
	notech_nor2 i_2481711(.A(n_413), .B(n_417), .Z(n_464));
	notech_nor2 i_2491710(.A(n_414), .B(n_418), .Z(n_465));
	notech_nor2 i_2501709(.A(n_415), .B(n_419), .Z(n_466));
	notech_nor2 i_2511708(.A(n_416), .B(n_249), .Z(n_467));
	notech_inv i_264(.A(n_433), .Z(n_480));
	notech_inv i_265(.A(n_434), .Z(n_481));
	notech_inv i_266(.A(n_435), .Z(n_482));
	notech_inv i_267(.A(n_436), .Z(n_483));
	notech_inv i_268(.A(n_437), .Z(n_484));
	notech_and2 i_549(.A(n_462), .B(n_454), .Z(n_707));
	notech_or2 i_550(.A(n_707), .B(n_438), .Z(n_708));
	notech_or2 i_553(.A(n_463), .B(n_439), .Z(n_710));
	notech_or2 i_556(.A(n_464), .B(n_440), .Z(n_712));
	notech_and2 i_558(.A(n_465), .B(n_433), .Z(n_713));
	notech_or2 i_559(.A(n_713), .B(n_441), .Z(n_714));
	notech_and2 i_561(.A(n_466), .B(n_434), .Z(n_715));
	notech_or2 i_562(.A(n_715), .B(n_442), .Z(n_716));
	notech_and2 i_564(.A(n_467), .B(n_435), .Z(n_717));
	notech_or2 i_565(.A(n_717), .B(n_443), .Z(n_718));
	notech_and2 i_567(.A(n_468), .B(n_436), .Z(n_719));
	notech_or2 i_568(.A(n_719), .B(n_444), .Z(n_720));
	notech_and2 i_570(.A(n_469), .B(n_437), .Z(n_721));
	notech_or2 i_571(.A(n_721), .B(n_445), .Z(n_722));
	notech_and2 i_573(.A(n_370802), .B(n_438), .Z(n_723));
	notech_or2 i_574(.A(n_723), .B(n_446), .Z(n_724));
	notech_inv i_575(.A(n_724), .Z(n_493));
	notech_and2 i_576(.A(n_471), .B(n_439), .Z(n_725));
	notech_or2 i_577(.A(n_725), .B(n_447), .Z(n_726));
	notech_inv i_578(.A(n_726), .Z(n_494));
	notech_or2 i_580(.A(n_727), .B(n_448), .Z(n_728));
	notech_inv i_581(.A(n_728), .Z(n_495));
	notech_or2 i_583(.A(n_729), .B(n_449), .Z(n_730));
	notech_inv i_584(.A(n_730), .Z(n_496));
	notech_or2 i_586(.A(n_731), .B(n_450), .Z(n_732));
	notech_inv i_587(.A(n_732), .Z(n_497));
	notech_or2 i_589(.A(n_733), .B(n_451), .Z(n_734));
	notech_inv i_590(.A(n_734), .Z(n_498));
	notech_or2 i_592(.A(n_735), .B(n_452), .Z(n_736));
	notech_inv i_593(.A(n_736), .Z(n_499));
	notech_or2 i_595(.A(n_737), .B(n_453), .Z(n_738));
	notech_inv i_596(.A(n_738), .Z(n_500));
	notech_inv i_285(.A(n_454), .Z(n_501));
	notech_nand2 i_301(.A(n_462), .B(n_370802), .Z(n_517));
	notech_nand2 i_302(.A(n_463), .B(n_471), .Z(n_518));
	notech_inv i_311(.A(n_480), .Z(n_527));
	notech_inv i_312(.A(n_481), .Z(n_528));
	notech_inv i_313(.A(n_482), .Z(n_529));
	notech_inv i_314(.A(n_483), .Z(n_530));
	notech_inv i_315(.A(n_484), .Z(n_531));
	notech_or2 i_597(.A(n_517), .B(n_501), .Z(n_740));
	notech_and2 i_598(.A(n_740), .B(n_493), .Z(n_739));
	notech_inv i_599(.A(n_739), .Z(n_540));
	notech_and2 i_601(.A(n_518), .B(n_494), .Z(n_741));
	notech_inv i_602(.A(n_741), .Z(n_541));
	notech_and2 i_604(.A(n_744), .B(n_495), .Z(n_743));
	notech_inv i_605(.A(n_743), .Z(n_542));
	notech_or2 i_606(.A(n_520), .B(n_480), .Z(n_746));
	notech_and2 i_607(.A(n_746), .B(n_496), .Z(n_745));
	notech_inv i_608(.A(n_745), .Z(n_543));
	notech_or2 i_609(.A(n_521), .B(n_481), .Z(n_748));
	notech_and2 i_610(.A(n_748), .B(n_497), .Z(n_747));
	notech_inv i_611(.A(n_747), .Z(n_544));
	notech_or2 i_612(.A(n_522), .B(n_482), .Z(n_750));
	notech_and2 i_613(.A(n_750), .B(n_498), .Z(n_749));
	notech_inv i_614(.A(n_749), .Z(n_545));
	notech_or2 i_615(.A(n_417), .B(n_483), .Z(n_752));
	notech_and2 i_616(.A(n_752), .B(n_499), .Z(n_751));
	notech_inv i_617(.A(n_751), .Z(n_546));
	notech_or2 i_618(.A(n_418), .B(n_484), .Z(n_754));
	notech_and2 i_619(.A(n_754), .B(n_500), .Z(n_753));
	notech_inv i_620(.A(n_753), .Z(n_547));
	notech_inv i_626(.A(n_757), .Z(i_psram_sub_function_sub[0]));
	notech_inv i_632(.A(n_762), .Z(i_psram_sub_function_sub[1]));
	notech_inv i_638(.A(n_767), .Z(i_psram_sub_function_sub[2]));
	notech_inv i_639(.A(n_527), .Z(n_770));
	notech_inv i_640(.A(n_296844), .Z(n_773));
	notech_nand2 i_641(.A(n_773), .B(n_527), .Z(n_774));
	notech_nand2 i_642(.A(n_296844), .B(n_770), .Z(n_771));
	notech_nand2 i_643(.A(n_771), .B(n_774), .Z(n_772));
	notech_inv i_644(.A(n_772), .Z(i_psram_sub_function_sub[3]));
	notech_inv i_645(.A(n_528), .Z(n_775));
	notech_inv i_646(.A(n_298842), .Z(n_778));
	notech_nand2 i_647(.A(n_778), .B(n_528), .Z(n_779));
	notech_nand2 i_648(.A(n_298842), .B(n_775), .Z(n_776));
	notech_nand2 i_649(.A(n_776), .B(n_779), .Z(n_777));
	notech_inv i_650(.A(n_777), .Z(i_psram_sub_function_sub[4]));
	notech_inv i_651(.A(n_529), .Z(n_780));
	notech_inv i_652(.A(n_300840), .Z(n_783));
	notech_nand2 i_653(.A(n_783), .B(n_529), .Z(n_784));
	notech_nand2 i_654(.A(n_300840), .B(n_780), .Z(n_781));
	notech_nand2 i_655(.A(n_781), .B(n_784), .Z(n_782));
	notech_inv i_656(.A(n_782), .Z(i_psram_sub_function_sub[5]));
	notech_inv i_657(.A(n_530), .Z(n_785));
	notech_inv i_658(.A(n_302838), .Z(n_788));
	notech_nand2 i_659(.A(n_788), .B(n_530), .Z(n_789));
	notech_nand2 i_660(.A(n_302838), .B(n_785), .Z(n_786));
	notech_nand2 i_661(.A(n_786), .B(n_789), .Z(n_787));
	notech_inv i_662(.A(n_787), .Z(i_psram_sub_function_sub[6]));
	notech_inv i_663(.A(n_531), .Z(n_790));
	notech_inv i_664(.A(n_304836), .Z(n_793));
	notech_nand2 i_665(.A(n_793), .B(n_531), .Z(n_794));
	notech_nand2 i_666(.A(n_304836), .B(n_790), .Z(n_791));
	notech_nand2 i_667(.A(n_791), .B(n_794), .Z(n_792));
	notech_inv i_668(.A(n_792), .Z(i_psram_sub_function_sub[7]));
	notech_inv i_669(.A(n_708), .Z(n_795));
	notech_inv i_670(.A(n_306834), .Z(n_798));
	notech_nand2 i_671(.A(n_798), .B(n_708), .Z(n_799));
	notech_nand2 i_672(.A(n_306834), .B(n_795), .Z(n_796));
	notech_nand2 i_673(.A(n_796), .B(n_799), .Z(n_797));
	notech_inv i_674(.A(n_797), .Z(i_psram_sub_function_sub[8]));
	notech_inv i_675(.A(n_710), .Z(n_800));
	notech_inv i_676(.A(n_308832), .Z(n_803));
	notech_nand2 i_677(.A(n_803), .B(n_710), .Z(n_804));
	notech_nand2 i_678(.A(n_308832), .B(n_800), .Z(n_801));
	notech_nand2 i_679(.A(n_801), .B(n_804), .Z(n_802));
	notech_inv i_680(.A(n_802), .Z(i_psram_sub_function_sub[9]));
	notech_inv i_681(.A(n_712), .Z(n_805));
	notech_inv i_682(.A(i_psram_sub_axi_araddr[10]), .Z(n_808));
	notech_nand2 i_683(.A(n_808), .B(n_712), .Z(n_809));
	notech_nand2 i_684(.A(i_psram_sub_axi_araddr[10]), .B(n_805), .Z(n_806)
		);
	notech_nand2 i_685(.A(n_806), .B(n_809), .Z(n_807));
	notech_inv i_686(.A(n_807), .Z(i_psram_sub_function_sub[10]));
	notech_inv i_687(.A(n_714), .Z(n_810));
	notech_inv i_688(.A(i_psram_sub_axi_araddr[11]), .Z(n_813));
	notech_nand2 i_689(.A(n_813), .B(n_714), .Z(n_814));
	notech_nand2 i_690(.A(i_psram_sub_axi_araddr[11]), .B(n_810), .Z(n_811)
		);
	notech_nand2 i_691(.A(n_811), .B(n_814), .Z(n_812));
	notech_inv i_692(.A(n_812), .Z(i_psram_sub_function_sub[11]));
	notech_inv i_693(.A(n_716), .Z(n_815));
	notech_inv i_694(.A(i_psram_sub_axi_araddr[12]), .Z(n_818));
	notech_nand2 i_695(.A(n_818), .B(n_716), .Z(n_819));
	notech_nand2 i_696(.A(i_psram_sub_axi_araddr[12]), .B(n_815), .Z(n_816)
		);
	notech_nand2 i_697(.A(n_816), .B(n_819), .Z(n_817));
	notech_inv i_698(.A(n_817), .Z(i_psram_sub_function_sub[12]));
	notech_inv i_699(.A(n_718), .Z(n_820));
	notech_inv i_700(.A(i_psram_sub_axi_araddr[13]), .Z(n_823));
	notech_nand2 i_701(.A(n_823), .B(n_718), .Z(n_824));
	notech_nand2 i_702(.A(i_psram_sub_axi_araddr[13]), .B(n_820), .Z(n_821)
		);
	notech_nand2 i_703(.A(n_821), .B(n_824), .Z(n_822));
	notech_inv i_704(.A(n_822), .Z(i_psram_sub_function_sub[13]));
	notech_inv i_705(.A(n_720), .Z(n_825));
	notech_inv i_706(.A(i_psram_sub_axi_araddr[14]), .Z(n_828));
	notech_nand2 i_707(.A(n_828), .B(n_720), .Z(n_829));
	notech_nand2 i_708(.A(i_psram_sub_axi_araddr[14]), .B(n_825), .Z(n_826)
		);
	notech_nand2 i_709(.A(n_826), .B(n_829), .Z(n_827));
	notech_inv i_710(.A(n_827), .Z(i_psram_sub_function_sub[14]));
	notech_inv i_711(.A(n_722), .Z(n_830));
	notech_inv i_712(.A(i_psram_sub_axi_araddr[15]), .Z(n_833));
	notech_nand2 i_713(.A(n_833), .B(n_722), .Z(n_834));
	notech_nand2 i_714(.A(i_psram_sub_axi_araddr[15]), .B(n_830), .Z(n_831)
		);
	notech_nand2 i_715(.A(n_831), .B(n_834), .Z(n_832));
	notech_inv i_716(.A(n_832), .Z(i_psram_sub_function_sub[15]));
	notech_inv i_717(.A(n_540), .Z(n_835));
	notech_inv i_718(.A(i_psram_sub_axi_araddr[16]), .Z(n_838));
	notech_nand2 i_719(.A(n_838), .B(n_540), .Z(n_839));
	notech_nand2 i_720(.A(i_psram_sub_axi_araddr[16]), .B(n_835), .Z(n_836)
		);
	notech_nand2 i_721(.A(n_836), .B(n_839), .Z(n_837));
	notech_inv i_722(.A(n_837), .Z(i_psram_sub_function_sub[16]));
	notech_inv i_723(.A(n_541), .Z(n_840));
	notech_inv i_724(.A(i_psram_sub_axi_araddr[17]), .Z(n_843));
	notech_nand2 i_725(.A(n_843), .B(n_541), .Z(n_844));
	notech_nand2 i_726(.A(i_psram_sub_axi_araddr[17]), .B(n_840), .Z(n_841)
		);
	notech_nand2 i_727(.A(n_841), .B(n_844), .Z(n_842));
	notech_inv i_728(.A(n_842), .Z(i_psram_sub_function_sub[17]));
	notech_inv i_729(.A(n_542), .Z(n_845));
	notech_inv i_730(.A(i_psram_sub_axi_araddr[18]), .Z(n_848));
	notech_nand2 i_731(.A(n_848), .B(n_542), .Z(n_849));
	notech_nand2 i_732(.A(i_psram_sub_axi_araddr[18]), .B(n_845), .Z(n_846)
		);
	notech_nand2 i_733(.A(n_846), .B(n_849), .Z(n_847));
	notech_inv i_734(.A(n_847), .Z(i_psram_sub_function_sub[18]));
	notech_inv i_735(.A(n_543), .Z(n_850));
	notech_inv i_736(.A(i_psram_sub_axi_araddr[19]), .Z(n_853));
	notech_nand2 i_737(.A(n_853), .B(n_543), .Z(n_854));
	notech_nand2 i_738(.A(i_psram_sub_axi_araddr[19]), .B(n_850), .Z(n_851)
		);
	notech_nand2 i_739(.A(n_851), .B(n_854), .Z(n_852));
	notech_inv i_740(.A(n_852), .Z(i_psram_sub_function_sub[19]));
	notech_inv i_741(.A(n_544), .Z(n_855));
	notech_inv i_742(.A(i_psram_sub_axi_araddr[20]), .Z(n_858));
	notech_nand2 i_743(.A(n_858), .B(n_544), .Z(n_859));
	notech_nand2 i_744(.A(i_psram_sub_axi_araddr[20]), .B(n_855), .Z(n_856)
		);
	notech_nand2 i_745(.A(n_856), .B(n_859), .Z(n_857));
	notech_inv i_746(.A(n_857), .Z(i_psram_sub_function_sub[20]));
	notech_inv i_747(.A(n_545), .Z(n_860));
	notech_inv i_748(.A(i_psram_sub_axi_araddr[21]), .Z(n_863));
	notech_nand2 i_749(.A(n_863), .B(n_545), .Z(n_864));
	notech_nand2 i_750(.A(i_psram_sub_axi_araddr[21]), .B(n_860), .Z(n_861)
		);
	notech_nand2 i_751(.A(n_861), .B(n_864), .Z(n_862));
	notech_inv i_752(.A(n_862), .Z(i_psram_sub_function_sub[21]));
	notech_inv i_753(.A(n_546), .Z(n_865));
	notech_inv i_754(.A(i_psram_sub_axi_araddr[22]), .Z(n_868));
	notech_nand2 i_755(.A(n_868), .B(n_546), .Z(n_869));
	notech_nand2 i_756(.A(i_psram_sub_axi_araddr[22]), .B(n_865), .Z(n_866)
		);
	notech_nand2 i_757(.A(n_866), .B(n_869), .Z(n_867));
	notech_inv i_758(.A(n_867), .Z(i_psram_sub_function_sub[22]));
	notech_inv i_759(.A(n_547), .Z(n_870));
	notech_inv i_760(.A(i_psram_sub_axi_araddr[23]), .Z(n_873));
	notech_nand2 i_761(.A(n_873), .B(n_547), .Z(n_874));
	notech_nand2 i_762(.A(i_psram_sub_axi_araddr[23]), .B(n_870), .Z(n_871)
		);
	notech_nand2 i_763(.A(n_871), .B(n_874), .Z(n_872));
	notech_inv i_764(.A(n_872), .Z(i_psram_sub_function_sub[23]));
	notech_inv i_0(.A(i_psram_sub_axi_araddr[2]), .Z(\i_psram_sub_axi_araddr_0[2] 
		));
	notech_nand2 i_1(.A(i_psram_sub_axi_araddr[2]), .B(i_psram_sub_axi_araddr
		[3]), .Z(n_133));
	notech_nand2 i_2(.A(i_psram_sub_axi_araddr[3]), .B(i_psram_sub_axi_araddr
		[4]), .Z(n_134));
	notech_nand2 i_3(.A(i_psram_sub_axi_araddr[4]), .B(i_psram_sub_axi_araddr
		[5]), .Z(n_135));
	notech_nand2 i_4(.A(i_psram_sub_axi_araddr[5]), .B(i_psram_sub_axi_araddr
		[6]), .Z(n_136));
	notech_nand2 i_5(.A(i_psram_sub_axi_araddr[6]), .B(i_psram_sub_axi_araddr
		[7]), .Z(n_137));
	notech_nand2 i_6(.A(i_psram_sub_axi_araddr[7]), .B(i_psram_sub_axi_araddr
		[8]), .Z(n_138));
	notech_nand2 i_7(.A(i_psram_sub_axi_araddr[8]), .B(i_psram_sub_axi_araddr
		[9]), .Z(n_139));
	notech_nand2 i_8(.A(i_psram_sub_axi_araddr[9]), .B(i_psram_sub_axi_araddr
		[10]), .Z(n_140));
	notech_nand2 i_9(.A(i_psram_sub_axi_araddr[10]), .B(i_psram_sub_axi_araddr
		[11]), .Z(n_141));
	notech_nand2 i_10(.A(i_psram_sub_axi_araddr[11]), .B(i_psram_sub_axi_araddr
		[12]), .Z(n_142));
	notech_nand2 i_11(.A(i_psram_sub_axi_araddr[12]), .B(i_psram_sub_axi_araddr
		[13]), .Z(n_143));
	notech_nand2 i_12(.A(i_psram_sub_axi_araddr[13]), .B(i_psram_sub_axi_araddr
		[14]), .Z(n_144));
	notech_nand2 i_13(.A(i_psram_sub_axi_araddr[14]), .B(i_psram_sub_axi_araddr
		[15]), .Z(n_145));
	notech_nand2 i_14(.A(i_psram_sub_axi_araddr[15]), .B(i_psram_sub_axi_araddr
		[16]), .Z(n_146));
	notech_nand2 i_15(.A(i_psram_sub_axi_araddr[16]), .B(i_psram_sub_axi_araddr
		[17]), .Z(n_147));
	notech_nand2 i_16(.A(i_psram_sub_axi_araddr[17]), .B(i_psram_sub_axi_araddr
		[18]), .Z(n_148));
	notech_nand2 i_17(.A(i_psram_sub_axi_araddr[18]), .B(i_psram_sub_axi_araddr
		[19]), .Z(n_149));
	notech_nand2 i_18(.A(i_psram_sub_axi_araddr[19]), .B(i_psram_sub_axi_araddr
		[20]), .Z(n_150));
	notech_nand2 i_19(.A(i_psram_sub_axi_araddr[20]), .B(i_psram_sub_axi_araddr
		[21]), .Z(n_151));
	notech_nand2 i_20(.A(i_psram_sub_axi_araddr[21]), .B(i_psram_sub_axi_araddr
		[22]), .Z(n_152));
	notech_inv i_22(.A(\i_psram_sub_axi_araddr_0[2] ), .Z(n_154));
	notech_inv i_23(.A(n_133), .Z(n_265));
	notech_nor2 i_24(.A(\i_psram_sub_axi_araddr_0[2] ), .B(n_134), .Z(n_156)
		);
	notech_nor2 i_25(.A(n_133), .B(n_135), .Z(n_157));
	notech_nor2 i_26(.A(n_134), .B(n_136), .Z(n_158));
	notech_nor2 i_27(.A(n_135), .B(n_137), .Z(n_159));
	notech_nor2 i_28(.A(n_136), .B(n_138), .Z(n_160));
	notech_nor2 i_29(.A(n_137), .B(n_139), .Z(n_161));
	notech_nor2 i_30(.A(n_138), .B(n_140), .Z(n_162));
	notech_nor2 i_31(.A(n_139), .B(n_141), .Z(n_163));
	notech_nor2 i_32(.A(n_140), .B(n_142), .Z(n_164));
	notech_nor2 i_33(.A(n_141), .B(n_143), .Z(n_165));
	notech_nor2 i_34(.A(n_142), .B(n_144), .Z(n_166));
	notech_nor2 i_35(.A(n_143), .B(n_145), .Z(n_167));
	notech_nor2 i_36(.A(n_144), .B(n_146), .Z(n_168));
	notech_nor2 i_37(.A(n_145), .B(n_147), .Z(n_169));
	notech_nor2 i_38(.A(n_146), .B(n_148), .Z(n_170));
	notech_nor2 i_39(.A(n_147), .B(n_149), .Z(n_171));
	notech_nor2 i_40(.A(n_148), .B(n_150), .Z(n_172));
	notech_nor2 i_41(.A(n_149), .B(n_151), .Z(n_173));
	notech_nor2 i_42(.A(n_150), .B(n_152), .Z(n_174));
	notech_inv i_44(.A(n_154), .Z(n_176));
	notech_inv i_45(.A(n_265), .Z(n_177));
	notech_inv i_46(.A(n_156), .Z(n_178));
	notech_inv i_47(.A(n_157), .Z(n_266));
	notech_nand2 i_48(.A(n_154), .B(n_158), .Z(n_180));
	notech_nand2 i_49(.A(n_265), .B(n_159), .Z(n_181));
	notech_nand2 i_50(.A(n_156), .B(n_160), .Z(n_182));
	notech_nand2 i_51(.A(n_157), .B(n_161), .Z(n_183));
	notech_nand2 i_52(.A(n_158), .B(n_162), .Z(n_184));
	notech_nand2 i_53(.A(n_159), .B(n_163), .Z(n_185));
	notech_nand2 i_54(.A(n_160), .B(n_164), .Z(n_186));
	notech_nand2 i_55(.A(n_161), .B(n_165), .Z(n_187));
	notech_nand2 i_56(.A(n_162), .B(n_166), .Z(n_188));
	notech_nand2 i_57(.A(n_163), .B(n_167), .Z(n_189));
	notech_nand2 i_58(.A(n_164), .B(n_168), .Z(n_190));
	notech_nand2 i_59(.A(n_165), .B(n_169), .Z(n_191));
	notech_nand2 i_60(.A(n_166), .B(n_170), .Z(n_192));
	notech_nand2 i_61(.A(n_167), .B(n_171), .Z(n_193));
	notech_nand2 i_62(.A(n_168), .B(n_172), .Z(n_194));
	notech_nand2 i_63(.A(n_169), .B(n_173), .Z(n_195));
	notech_nand2 i_64(.A(n_170), .B(n_174), .Z(n_196));
	notech_inv i_66(.A(n_176), .Z(n_198));
	notech_inv i_67(.A(n_177), .Z(n_199));
	notech_inv i_68(.A(n_178), .Z(n_200));
	notech_inv i_69(.A(n_266), .Z(n_201));
	notech_inv i_70(.A(n_180), .Z(n_202));
	notech_nor2 i_74(.A(n_176), .B(n_184), .Z(n_206));
	notech_nor2 i_75(.A(n_177), .B(n_185), .Z(n_207));
	notech_nor2 i_76(.A(n_178), .B(n_186), .Z(n_208));
	notech_nor2 i_77(.A(n_266), .B(n_187), .Z(n_209));
	notech_nor2 i_78(.A(n_180), .B(n_188), .Z(n_210));
	notech_nor2 i_79(.A(n_181), .B(n_189), .Z(n_211));
	notech_nor2 i_80(.A(n_182), .B(n_190), .Z(n_212));
	notech_nor2 i_81(.A(n_183), .B(n_191), .Z(n_213));
	notech_nor2 i_82(.A(n_184), .B(n_192), .Z(n_214));
	notech_nor2 i_83(.A(n_185), .B(n_193), .Z(n_215));
	notech_nor2 i_84(.A(n_186), .B(n_194), .Z(n_216));
	notech_nor2 i_85(.A(n_187), .B(n_195), .Z(n_217));
	notech_nor2 i_86(.A(n_188), .B(n_196), .Z(n_218));
	notech_inv i_88(.A(n_198), .Z(n_220));
	notech_inv i_89(.A(n_199), .Z(n_221));
	notech_inv i_90(.A(n_200), .Z(n_222));
	notech_inv i_91(.A(n_201), .Z(n_223));
	notech_inv i_92(.A(n_202), .Z(n_224));
	notech_inv i_96(.A(n_206), .Z(n_228));
	notech_inv i_97(.A(n_207), .Z(n_229));
	notech_inv i_98(.A(n_208), .Z(n_230));
	notech_inv i_99(.A(n_209), .Z(n_231));
	notech_inv i_100(.A(n_210), .Z(n_232));
	notech_inv i_101(.A(n_211), .Z(n_233));
	notech_inv i_102(.A(n_212), .Z(n_234));
	notech_inv i_103(.A(n_213), .Z(n_272));
	notech_nand2 i_104(.A(n_198), .B(n_214), .Z(n_236));
	notech_nand2 i_105(.A(n_199), .B(n_215), .Z(n_237));
	notech_nand2 i_106(.A(n_200), .B(n_216), .Z(n_238));
	notech_nand2 i_107(.A(n_201), .B(n_217), .Z(n_239));
	notech_nand2 i_108(.A(n_202), .B(n_218), .Z(n_240));
	notech_inv i_132(.A(n_220), .Z(n_276));
	notech_inv i_133(.A(i_psram_sub_axi_araddr[3]), .Z(n_279));
	notech_nand2 i_134(.A(n_279), .B(n_220), .Z(n_280));
	notech_nand2 i_135(.A(i_psram_sub_axi_araddr[3]), .B(n_276), .Z(n_277)
		);
	notech_nand2 i_136(.A(n_277), .B(n_280), .Z(n_278));
	notech_inv i_137(.A(n_278), .Z(\i_psram_sub_axi_araddr_0[3] ));
	notech_inv i_138(.A(n_221), .Z(n_281));
	notech_inv i_139(.A(i_psram_sub_axi_araddr[4]), .Z(n_284));
	notech_nand2 i_140(.A(n_284), .B(n_221), .Z(n_285));
	notech_nand2 i_141(.A(i_psram_sub_axi_araddr[4]), .B(n_281), .Z(n_282)
		);
	notech_nand2 i_142(.A(n_282), .B(n_285), .Z(n_283));
	notech_inv i_143(.A(n_283), .Z(\i_psram_sub_axi_araddr_0[4] ));
	notech_inv i_144(.A(n_222), .Z(n_286));
	notech_inv i_145(.A(i_psram_sub_axi_araddr[5]), .Z(n_289));
	notech_nand2 i_146(.A(n_289), .B(n_222), .Z(n_290));
	notech_nand2 i_147(.A(i_psram_sub_axi_araddr[5]), .B(n_286), .Z(n_287)
		);
	notech_nand2 i_148(.A(n_287), .B(n_290), .Z(n_288));
	notech_inv i_149(.A(n_288), .Z(\i_psram_sub_axi_araddr_0[5] ));
	notech_inv i_150(.A(n_223), .Z(n_291));
	notech_inv i_151(.A(i_psram_sub_axi_araddr[6]), .Z(n_294));
	notech_nand2 i_152(.A(n_294), .B(n_223), .Z(n_295));
	notech_nand2 i_153(.A(i_psram_sub_axi_araddr[6]), .B(n_291), .Z(n_292)
		);
	notech_nand2 i_154(.A(n_292), .B(n_295), .Z(n_293));
	notech_inv i_155(.A(n_293), .Z(\i_psram_sub_axi_araddr_0[6] ));
	notech_inv i_156(.A(n_224), .Z(n_296));
	notech_inv i_157(.A(i_psram_sub_axi_araddr[7]), .Z(n_299));
	notech_nand2 i_158(.A(n_299), .B(n_224), .Z(n_300));
	notech_nand2 i_159(.A(i_psram_sub_axi_araddr[7]), .B(n_296), .Z(n_297)
		);
	notech_nand2 i_160(.A(n_297), .B(n_300), .Z(n_298));
	notech_inv i_161(.A(n_298), .Z(\i_psram_sub_axi_araddr_0[7] ));
	notech_inv i_162(.A(n_181), .Z(n_301));
	notech_inv i_163(.A(i_psram_sub_axi_araddr[8]), .Z(n_304));
	notech_nand2 i_164(.A(n_304), .B(n_181), .Z(n_305));
	notech_nand2 i_165(.A(i_psram_sub_axi_araddr[8]), .B(n_301), .Z(n_302)
		);
	notech_nand2 i_166(.A(n_302), .B(n_305), .Z(n_303));
	notech_inv i_167(.A(n_303), .Z(\i_psram_sub_axi_araddr_0[8] ));
	notech_inv i_168(.A(n_182), .Z(n_306));
	notech_inv i_169(.A(i_psram_sub_axi_araddr[9]), .Z(n_309));
	notech_nand2 i_170(.A(n_309), .B(n_182), .Z(n_310));
	notech_nand2 i_171(.A(i_psram_sub_axi_araddr[9]), .B(n_306), .Z(n_307)
		);
	notech_nand2 i_172(.A(n_307), .B(n_310), .Z(n_308));
	notech_inv i_173(.A(n_308), .Z(\i_psram_sub_axi_araddr_0[9] ));
	notech_inv i_174(.A(n_183), .Z(n_311));
	notech_inv i_175(.A(i_psram_sub_axi_araddr[10]), .Z(n_314));
	notech_nand2 i_176(.A(n_314), .B(n_183), .Z(n_315));
	notech_nand2 i_177(.A(i_psram_sub_axi_araddr[10]), .B(n_311), .Z(n_312)
		);
	notech_nand2 i_178(.A(n_312), .B(n_315), .Z(n_313));
	notech_inv i_179(.A(n_313), .Z(\i_psram_sub_axi_araddr_0[10] ));
	notech_inv i_180(.A(n_228), .Z(n_316));
	notech_inv i_181(.A(i_psram_sub_axi_araddr[11]), .Z(n_319));
	notech_nand2 i_182(.A(n_319), .B(n_228), .Z(n_320));
	notech_nand2 i_183(.A(i_psram_sub_axi_araddr[11]), .B(n_316), .Z(n_317)
		);
	notech_nand2 i_184(.A(n_317), .B(n_320), .Z(n_318));
	notech_inv i_185(.A(n_318), .Z(\i_psram_sub_axi_araddr_0[11] ));
	notech_inv i_186(.A(n_229), .Z(n_321));
	notech_inv i_187(.A(i_psram_sub_axi_araddr[12]), .Z(n_324));
	notech_nand2 i_188(.A(n_324), .B(n_229), .Z(n_325));
	notech_nand2 i_189(.A(i_psram_sub_axi_araddr[12]), .B(n_321), .Z(n_322)
		);
	notech_nand2 i_190(.A(n_322), .B(n_325), .Z(n_323));
	notech_inv i_191(.A(n_323), .Z(\i_psram_sub_axi_araddr_0[12] ));
	notech_inv i_192(.A(n_230), .Z(n_326));
	notech_inv i_193(.A(i_psram_sub_axi_araddr[13]), .Z(n_329));
	notech_nand2 i_194(.A(n_329), .B(n_230), .Z(n_330));
	notech_nand2 i_195(.A(i_psram_sub_axi_araddr[13]), .B(n_326), .Z(n_327)
		);
	notech_nand2 i_196(.A(n_327), .B(n_330), .Z(n_328));
	notech_inv i_197(.A(n_328), .Z(\i_psram_sub_axi_araddr_0[13] ));
	notech_inv i_198(.A(n_231), .Z(n_331));
	notech_inv i_199(.A(i_psram_sub_axi_araddr[14]), .Z(n_334));
	notech_nand2 i_200(.A(n_334), .B(n_231), .Z(n_335));
	notech_nand2 i_201(.A(i_psram_sub_axi_araddr[14]), .B(n_331), .Z(n_332)
		);
	notech_nand2 i_202(.A(n_332), .B(n_335), .Z(n_333));
	notech_inv i_203(.A(n_333), .Z(\i_psram_sub_axi_araddr_0[14] ));
	notech_inv i_204(.A(n_232), .Z(n_336));
	notech_inv i_205(.A(i_psram_sub_axi_araddr[15]), .Z(n_339));
	notech_nand2 i_206(.A(n_339), .B(n_232), .Z(n_340));
	notech_nand2 i_207(.A(i_psram_sub_axi_araddr[15]), .B(n_336), .Z(n_337)
		);
	notech_nand2 i_208(.A(n_337), .B(n_340), .Z(n_338));
	notech_inv i_209(.A(n_338), .Z(\i_psram_sub_axi_araddr_0[15] ));
	notech_inv i_210(.A(n_233), .Z(n_341));
	notech_inv i_211(.A(i_psram_sub_axi_araddr[16]), .Z(n_344));
	notech_nand2 i_212(.A(n_344), .B(n_233), .Z(n_345));
	notech_nand2 i_213(.A(i_psram_sub_axi_araddr[16]), .B(n_341), .Z(n_342)
		);
	notech_nand2 i_214(.A(n_342), .B(n_345), .Z(n_343));
	notech_inv i_215(.A(n_343), .Z(\i_psram_sub_axi_araddr_0[16] ));
	notech_inv i_216(.A(n_234), .Z(n_346));
	notech_inv i_217(.A(i_psram_sub_axi_araddr[17]), .Z(n_349));
	notech_nand2 i_218(.A(n_349), .B(n_234), .Z(n_350));
	notech_nand2 i_219(.A(i_psram_sub_axi_araddr[17]), .B(n_346), .Z(n_347)
		);
	notech_nand2 i_220(.A(n_347), .B(n_350), .Z(n_348));
	notech_inv i_221(.A(n_348), .Z(\i_psram_sub_axi_araddr_0[17] ));
	notech_inv i_222(.A(n_272), .Z(n_351));
	notech_inv i_223(.A(i_psram_sub_axi_araddr[18]), .Z(n_354));
	notech_nand2 i_224(.A(n_354), .B(n_272), .Z(n_355));
	notech_nand2 i_225(.A(i_psram_sub_axi_araddr[18]), .B(n_351), .Z(n_352)
		);
	notech_nand2 i_226(.A(n_352), .B(n_355), .Z(n_353));
	notech_inv i_227(.A(n_353), .Z(\i_psram_sub_axi_araddr_0[18] ));
	notech_inv i_228(.A(n_236), .Z(n_356));
	notech_inv i_229(.A(i_psram_sub_axi_araddr[19]), .Z(n_359));
	notech_nand2 i_230(.A(n_359), .B(n_236), .Z(n_360));
	notech_nand2 i_231(.A(i_psram_sub_axi_araddr[19]), .B(n_356), .Z(n_357)
		);
	notech_nand2 i_232(.A(n_357), .B(n_360), .Z(n_358));
	notech_inv i_233(.A(n_358), .Z(\i_psram_sub_axi_araddr_0[19] ));
	notech_inv i_234(.A(n_237), .Z(n_361));
	notech_inv i_235(.A(i_psram_sub_axi_araddr[20]), .Z(n_364));
	notech_nand2 i_236(.A(n_364), .B(n_237), .Z(n_365));
	notech_nand2 i_237(.A(i_psram_sub_axi_araddr[20]), .B(n_361), .Z(n_362)
		);
	notech_nand2 i_238(.A(n_362), .B(n_365), .Z(n_363));
	notech_inv i_239(.A(n_363), .Z(\i_psram_sub_axi_araddr_0[20] ));
	notech_inv i_240(.A(n_238), .Z(n_366));
	notech_inv i_241(.A(i_psram_sub_axi_araddr[21]), .Z(n_369));
	notech_nand2 i_242(.A(n_369), .B(n_238), .Z(n_370));
	notech_nand2 i_243(.A(i_psram_sub_axi_araddr[21]), .B(n_366), .Z(n_367)
		);
	notech_nand2 i_244(.A(n_367), .B(n_370), .Z(n_368));
	notech_inv i_245(.A(n_368), .Z(\i_psram_sub_axi_araddr_0[21] ));
	notech_inv i_246(.A(n_239), .Z(n_371));
	notech_inv i_247(.A(i_psram_sub_axi_araddr[22]), .Z(n_374));
	notech_nand2 i_248(.A(n_374), .B(n_239), .Z(n_375));
	notech_nand2 i_249(.A(i_psram_sub_axi_araddr[22]), .B(n_371), .Z(n_372)
		);
	notech_nand2 i_250(.A(n_372), .B(n_375), .Z(n_373));
	notech_inv i_251(.A(n_373), .Z(\i_psram_sub_axi_araddr_0[22] ));
	notech_inv i_252(.A(n_240), .Z(n_376));
	notech_inv i_253(.A(i_psram_sub_axi_araddr[23]), .Z(n_379));
	notech_nand2 i_254(.A(n_379), .B(n_240), .Z(n_380));
	notech_nand2 i_255(.A(i_psram_sub_axi_araddr[23]), .B(n_376), .Z(n_377)
		);
	notech_nand2 i_256(.A(n_377), .B(n_380), .Z(n_378));
	notech_inv i_257(.A(n_378), .Z(\i_psram_sub_axi_araddr_0[23] ));
	notech_inv i_psram_sub_i_5222(.A(s00_axi_awready), .Z(i_psram_sub_n_4399
		));
	notech_inv i_psram_sub_i_5221(.A(i_psram_sub_go), .Z(i_psram_sub_n_4398)
		);
	notech_inv i_psram_sub_i_5220(.A(\i_psram_sub_axi_rdata_0[16] ), .Z(i_psram_sub_n_4397
		));
	notech_inv i_psram_sub_i_5219(.A(\i_psram_sub_axi_rdata_0[17] ), .Z(i_psram_sub_n_4396
		));
	notech_inv i_psram_sub_i_5218(.A(\i_psram_sub_axi_rdata_0[18] ), .Z(i_psram_sub_n_4395
		));
	notech_inv i_psram_sub_i_5217(.A(\i_psram_sub_axi_rdata_0[19] ), .Z(i_psram_sub_n_4394
		));
	notech_inv i_psram_sub_i_5216(.A(\i_psram_sub_axi_rdata_0[20] ), .Z(i_psram_sub_n_4393
		));
	notech_inv i_psram_sub_i_5215(.A(\i_psram_sub_axi_rdata_0[21] ), .Z(i_psram_sub_n_4392
		));
	notech_inv i_psram_sub_i_5214(.A(\i_psram_sub_axi_rdata_0[22] ), .Z(i_psram_sub_n_4391
		));
	notech_inv i_psram_sub_i_5213(.A(\i_psram_sub_axi_rdata_0[23] ), .Z(i_psram_sub_n_4390
		));
	notech_inv i_psram_sub_i_5212(.A(\i_psram_sub_axi_rdata_0[24] ), .Z(i_psram_sub_n_4389
		));
	notech_inv i_psram_sub_i_5211(.A(\i_psram_sub_axi_rdata_0[25] ), .Z(i_psram_sub_n_4388
		));
	notech_inv i_psram_sub_i_5210(.A(\i_psram_sub_axi_rdata_0[26] ), .Z(i_psram_sub_n_4387
		));
	notech_inv i_psram_sub_i_5209(.A(\i_psram_sub_axi_rdata_0[27] ), .Z(i_psram_sub_n_4386
		));
	notech_inv i_psram_sub_i_5208(.A(\i_psram_sub_axi_rdata_0[28] ), .Z(i_psram_sub_n_4385
		));
	notech_inv i_psram_sub_i_5207(.A(\i_psram_sub_axi_rdata_0[29] ), .Z(i_psram_sub_n_4384
		));
	notech_inv i_psram_sub_i_5206(.A(\i_psram_sub_axi_rdata_0[30] ), .Z(i_psram_sub_n_4383
		));
	notech_inv i_psram_sub_i_5205(.A(\i_psram_sub_axi_rdata_0[31] ), .Z(i_psram_sub_n_4382
		));
	notech_inv i_psram_sub_i_5204(.A(\i_psram_sub_axi_awaddr_0[2] ), .Z(i_psram_sub_n_4381
		));
	notech_inv i_psram_sub_i_5203(.A(\i_psram_sub_axi_awaddr_0[3] ), .Z(i_psram_sub_n_4380
		));
	notech_inv i_psram_sub_i_5202(.A(\i_psram_sub_axi_awaddr_0[4] ), .Z(i_psram_sub_n_4379
		));
	notech_inv i_psram_sub_i_5201(.A(\i_psram_sub_axi_awaddr_0[5] ), .Z(i_psram_sub_n_4378
		));
	notech_inv i_psram_sub_i_5200(.A(\i_psram_sub_axi_awaddr_0[6] ), .Z(i_psram_sub_n_4377
		));
	notech_inv i_psram_sub_i_5199(.A(\i_psram_sub_axi_awaddr_0[7] ), .Z(i_psram_sub_n_4376
		));
	notech_inv i_psram_sub_i_5198(.A(\i_psram_sub_axi_awaddr_0[8] ), .Z(i_psram_sub_n_4375
		));
	notech_inv i_psram_sub_i_5197(.A(\i_psram_sub_axi_awaddr_0[9] ), .Z(i_psram_sub_n_4374
		));
	notech_inv i_psram_sub_i_5196(.A(\i_psram_sub_axi_awaddr_0[10] ), .Z(i_psram_sub_n_4373
		));
	notech_inv i_psram_sub_i_5195(.A(\i_psram_sub_axi_awaddr_0[11] ), .Z(i_psram_sub_n_4372
		));
	notech_inv i_psram_sub_i_5194(.A(\i_psram_sub_axi_awaddr_0[12] ), .Z(i_psram_sub_n_4371
		));
	notech_inv i_psram_sub_i_5193(.A(\i_psram_sub_axi_awaddr_0[13] ), .Z(i_psram_sub_n_4370
		));
	notech_inv i_psram_sub_i_5192(.A(\i_psram_sub_axi_awaddr_0[14] ), .Z(i_psram_sub_n_4369
		));
	notech_inv i_psram_sub_i_5191(.A(\i_psram_sub_axi_awaddr_0[15] ), .Z(i_psram_sub_n_4368
		));
	notech_inv i_psram_sub_i_5190(.A(\i_psram_sub_axi_awaddr_0[16] ), .Z(i_psram_sub_n_4367
		));
	notech_inv i_psram_sub_i_5189(.A(\i_psram_sub_axi_awaddr_0[17] ), .Z(i_psram_sub_n_4366
		));
	notech_inv i_psram_sub_i_5188(.A(\i_psram_sub_axi_awaddr_0[18] ), .Z(i_psram_sub_n_4365
		));
	notech_inv i_psram_sub_i_5187(.A(\i_psram_sub_axi_awaddr_0[19] ), .Z(i_psram_sub_n_4364
		));
	notech_inv i_psram_sub_i_5186(.A(\i_psram_sub_axi_awaddr_0[20] ), .Z(i_psram_sub_n_4363
		));
	notech_inv i_psram_sub_i_5185(.A(\i_psram_sub_axi_awaddr_0[21] ), .Z(i_psram_sub_n_4362
		));
	notech_inv i_psram_sub_i_5184(.A(\i_psram_sub_axi_awaddr_0[22] ), .Z(i_psram_sub_n_4361
		));
	notech_inv i_psram_sub_i_5183(.A(\i_psram_sub_axi_awaddr_0[23] ), .Z(i_psram_sub_n_4360
		));
	notech_inv i_psram_sub_i_5182(.A(s00_axi_awlen[0]), .Z(i_psram_sub_n_4359
		));
	notech_inv i_psram_sub_i_5181(.A(s00_axi_awlen[1]), .Z(i_psram_sub_n_4358
		));
	notech_inv i_psram_sub_i_5180(.A(s00_axi_awlen[2]), .Z(i_psram_sub_n_4357
		));
	notech_inv i_psram_sub_i_5179(.A(s00_axi_awlen[3]), .Z(i_psram_sub_n_4356
		));
	notech_inv i_psram_sub_i_5178(.A(s00_axi_awlen[4]), .Z(i_psram_sub_n_4355
		));
	notech_inv i_psram_sub_i_5177(.A(s00_axi_awlen[5]), .Z(i_psram_sub_n_4354
		));
	notech_inv i_psram_sub_i_5176(.A(s00_axi_awlen[6]), .Z(i_psram_sub_n_4353
		));
	notech_inv i_psram_sub_i_5175(.A(s00_axi_awlen[7]), .Z(i_psram_sub_n_4352
		));
	notech_inv i_psram_sub_i_5174(.A(\i_psram_sub_axi_araddr_0[2] ), .Z(i_psram_sub_n_4351
		));
	notech_inv i_psram_sub_i_5173(.A(\i_psram_sub_axi_araddr_0[3] ), .Z(i_psram_sub_n_4350
		));
	notech_inv i_psram_sub_i_5172(.A(\i_psram_sub_axi_araddr_0[4] ), .Z(i_psram_sub_n_4349
		));
	notech_inv i_psram_sub_i_5171(.A(\i_psram_sub_axi_araddr_0[5] ), .Z(i_psram_sub_n_4348
		));
	notech_inv i_psram_sub_i_5170(.A(\i_psram_sub_axi_araddr_0[6] ), .Z(i_psram_sub_n_4347
		));
	notech_inv i_psram_sub_i_5169(.A(\i_psram_sub_axi_araddr_0[7] ), .Z(i_psram_sub_n_4346
		));
	notech_inv i_psram_sub_i_5168(.A(\i_psram_sub_axi_araddr_0[8] ), .Z(i_psram_sub_n_4345
		));
	notech_inv i_psram_sub_i_5167(.A(\i_psram_sub_axi_araddr_0[9] ), .Z(i_psram_sub_n_4344
		));
	notech_inv i_psram_sub_i_5166(.A(\i_psram_sub_axi_araddr_0[10] ), .Z(i_psram_sub_n_4343
		));
	notech_inv i_psram_sub_i_5165(.A(\i_psram_sub_axi_araddr_0[11] ), .Z(i_psram_sub_n_4342
		));
	notech_inv i_psram_sub_i_5164(.A(\i_psram_sub_axi_araddr_0[12] ), .Z(i_psram_sub_n_4341
		));
	notech_inv i_psram_sub_i_5163(.A(\i_psram_sub_axi_araddr_0[13] ), .Z(i_psram_sub_n_4340
		));
	notech_inv i_psram_sub_i_5162(.A(\i_psram_sub_axi_araddr_0[14] ), .Z(i_psram_sub_n_4339
		));
	notech_inv i_psram_sub_i_5161(.A(\i_psram_sub_axi_araddr_0[15] ), .Z(i_psram_sub_n_4338
		));
	notech_inv i_psram_sub_i_5160(.A(\i_psram_sub_axi_araddr_0[16] ), .Z(i_psram_sub_n_4337
		));
	notech_inv i_psram_sub_i_5159(.A(\i_psram_sub_axi_araddr_0[17] ), .Z(i_psram_sub_n_4336
		));
	notech_inv i_psram_sub_i_5158(.A(\i_psram_sub_axi_araddr_0[18] ), .Z(i_psram_sub_n_4335
		));
	notech_inv i_psram_sub_i_5157(.A(\i_psram_sub_axi_araddr_0[19] ), .Z(i_psram_sub_n_4334
		));
	notech_inv i_psram_sub_i_5156(.A(\i_psram_sub_axi_araddr_0[20] ), .Z(i_psram_sub_n_4333
		));
	notech_inv i_psram_sub_i_5155(.A(\i_psram_sub_axi_araddr_0[21] ), .Z(i_psram_sub_n_4332
		));
	notech_inv i_psram_sub_i_5154(.A(\i_psram_sub_axi_araddr_0[22] ), .Z(i_psram_sub_n_4331
		));
	notech_inv i_psram_sub_i_5153(.A(\i_psram_sub_axi_araddr_0[23] ), .Z(i_psram_sub_n_4330
		));
	notech_inv i_psram_sub_i_5152(.A(s00_axi_arlen[0]), .Z(i_psram_sub_n_4329
		));
	notech_inv i_psram_sub_i_5151(.A(s00_axi_arlen[1]), .Z(i_psram_sub_n_4328
		));
	notech_inv i_psram_sub_i_5150(.A(s00_axi_arlen[2]), .Z(i_psram_sub_n_4327
		));
	notech_inv i_psram_sub_i_5149(.A(s00_axi_arlen[3]), .Z(i_psram_sub_n_4326
		));
	notech_inv i_psram_sub_i_5148(.A(s00_axi_arlen[4]), .Z(i_psram_sub_n_4325
		));
	notech_inv i_psram_sub_i_5147(.A(s00_axi_arlen[5]), .Z(i_psram_sub_n_4324
		));
	notech_inv i_psram_sub_i_5146(.A(s00_axi_arlen[6]), .Z(i_psram_sub_n_4323
		));
	notech_inv i_psram_sub_i_5145(.A(s00_axi_arlen[7]), .Z(i_psram_sub_n_4322
		));
	notech_inv i_psram_sub_i_5144(.A(s00_axi_wvalid), .Z(i_psram_sub_n_4321)
		);
	notech_inv i_psram_sub_i_5143(.A(i_psram_sub_mem_idle), .Z(i_psram_sub_n_4320
		));
	notech_inv i_psram_sub_i_5142(.A(s00_axi_aresetn), .Z(i_psram_sub_n_4319
		));
	notech_inv i_psram_sub_i_5141(.A(s00_axi_arburst[1]), .Z(i_psram_sub_n_4318
		));
	notech_inv i_psram_sub_i_5140(.A(s00_axi_awburst[1]), .Z(i_psram_sub_n_4317
		));
	notech_inv i_psram_sub_i_5139(.A(s00_axi_awburst[0]), .Z(i_psram_sub_n_4316
		));
	notech_inv i_psram_sub_i_5138(.A(s00_axi_wstrb[3]), .Z(i_psram_sub_n_4315
		));
	notech_inv i_psram_sub_i_5137(.A(s00_axi_wstrb[2]), .Z(i_psram_sub_n_4314
		));
	notech_inv i_psram_sub_i_5136(.A(s00_axi_rdata[31]), .Z(i_psram_sub_n_4313
		));
	notech_inv i_psram_sub_i_5135(.A(s00_axi_rdata[30]), .Z(i_psram_sub_n_4312
		));
	notech_inv i_psram_sub_i_5134(.A(s00_axi_rdata[29]), .Z(i_psram_sub_n_4311
		));
	notech_inv i_psram_sub_i_5133(.A(s00_axi_rdata[28]), .Z(i_psram_sub_n_4310
		));
	notech_inv i_psram_sub_i_5132(.A(s00_axi_rdata[27]), .Z(i_psram_sub_n_4309
		));
	notech_inv i_psram_sub_i_5131(.A(s00_axi_rdata[26]), .Z(i_psram_sub_n_4308
		));
	notech_inv i_psram_sub_i_5130(.A(s00_axi_rdata[25]), .Z(i_psram_sub_n_4307
		));
	notech_inv i_psram_sub_i_5129(.A(s00_axi_rdata[24]), .Z(i_psram_sub_n_4306
		));
	notech_inv i_psram_sub_i_5128(.A(s00_axi_rdata[23]), .Z(i_psram_sub_n_4305
		));
	notech_inv i_psram_sub_i_5127(.A(s00_axi_rdata[22]), .Z(i_psram_sub_n_4304
		));
	notech_inv i_psram_sub_i_5126(.A(s00_axi_rdata[21]), .Z(i_psram_sub_n_4303
		));
	notech_inv i_psram_sub_i_5125(.A(s00_axi_rdata[20]), .Z(i_psram_sub_n_4302
		));
	notech_inv i_psram_sub_i_5124(.A(s00_axi_rdata[19]), .Z(i_psram_sub_n_4301
		));
	notech_inv i_psram_sub_i_5123(.A(s00_axi_rdata[18]), .Z(i_psram_sub_n_4300
		));
	notech_inv i_psram_sub_i_5122(.A(s00_axi_rdata[17]), .Z(i_psram_sub_n_4299
		));
	notech_inv i_psram_sub_i_5121(.A(s00_axi_rdata[16]), .Z(i_psram_sub_n_4298
		));
	notech_inv i_psram_sub_i_5120(.A(s00_axi_rdata[15]), .Z(i_psram_sub_n_4297
		));
	notech_inv i_psram_sub_i_5119(.A(s00_axi_rdata[14]), .Z(i_psram_sub_n_4296
		));
	notech_inv i_psram_sub_i_5118(.A(s00_axi_rdata[13]), .Z(i_psram_sub_n_4295
		));
	notech_inv i_psram_sub_i_5117(.A(s00_axi_rdata[12]), .Z(i_psram_sub_n_4294
		));
	notech_inv i_psram_sub_i_5116(.A(s00_axi_rdata[11]), .Z(i_psram_sub_n_4293
		));
	notech_inv i_psram_sub_i_5115(.A(s00_axi_rdata[10]), .Z(i_psram_sub_n_4292
		));
	notech_inv i_psram_sub_i_5114(.A(s00_axi_rdata[9]), .Z(i_psram_sub_n_4291
		));
	notech_inv i_psram_sub_i_5113(.A(s00_axi_rdata[8]), .Z(i_psram_sub_n_4290
		));
	notech_inv i_psram_sub_i_5112(.A(s00_axi_rdata[7]), .Z(i_psram_sub_n_4289
		));
	notech_inv i_psram_sub_i_5111(.A(s00_axi_rdata[6]), .Z(i_psram_sub_n_4288
		));
	notech_inv i_psram_sub_i_5110(.A(s00_axi_rdata[5]), .Z(i_psram_sub_n_4287
		));
	notech_inv i_psram_sub_i_5109(.A(s00_axi_rdata[4]), .Z(i_psram_sub_n_4286
		));
	notech_inv i_psram_sub_i_5108(.A(s00_axi_rdata[3]), .Z(i_psram_sub_n_4285
		));
	notech_inv i_psram_sub_i_5107(.A(s00_axi_rdata[2]), .Z(i_psram_sub_n_4284
		));
	notech_inv i_psram_sub_i_5106(.A(s00_axi_rdata[1]), .Z(i_psram_sub_n_4283
		));
	notech_inv i_psram_sub_i_5105(.A(s00_axi_rdata[0]), .Z(i_psram_sub_n_4282
		));
	notech_inv i_psram_sub_i_5104(.A(s00_axi_awaddr[23]), .Z(i_psram_sub_n_4281
		));
	notech_inv i_psram_sub_i_5103(.A(s00_axi_awaddr[22]), .Z(i_psram_sub_n_4280
		));
	notech_inv i_psram_sub_i_5102(.A(s00_axi_awaddr[21]), .Z(i_psram_sub_n_4279
		));
	notech_inv i_psram_sub_i_5101(.A(s00_axi_awaddr[20]), .Z(i_psram_sub_n_4278
		));
	notech_inv i_psram_sub_i_5100(.A(s00_axi_awaddr[19]), .Z(i_psram_sub_n_4277
		));
	notech_inv i_psram_sub_i_5099(.A(s00_axi_awaddr[18]), .Z(i_psram_sub_n_4276
		));
	notech_inv i_psram_sub_i_5098(.A(s00_axi_awaddr[17]), .Z(i_psram_sub_n_4275
		));
	notech_inv i_psram_sub_i_5097(.A(s00_axi_awaddr[16]), .Z(i_psram_sub_n_4274
		));
	notech_inv i_psram_sub_i_5096(.A(s00_axi_awaddr[15]), .Z(i_psram_sub_n_4273
		));
	notech_inv i_psram_sub_i_5095(.A(s00_axi_awaddr[14]), .Z(i_psram_sub_n_4272
		));
	notech_inv i_psram_sub_i_5094(.A(s00_axi_awaddr[13]), .Z(i_psram_sub_n_4271
		));
	notech_inv i_psram_sub_i_5093(.A(s00_axi_awaddr[12]), .Z(i_psram_sub_n_4270
		));
	notech_inv i_psram_sub_i_5092(.A(s00_axi_awaddr[11]), .Z(i_psram_sub_n_4269
		));
	notech_inv i_psram_sub_i_5091(.A(s00_axi_awaddr[10]), .Z(i_psram_sub_n_4268
		));
	notech_inv i_psram_sub_i_5090(.A(s00_axi_awaddr[9]), .Z(i_psram_sub_n_4267
		));
	notech_inv i_psram_sub_i_5089(.A(s00_axi_awaddr[8]), .Z(i_psram_sub_n_4266
		));
	notech_inv i_psram_sub_i_5088(.A(s00_axi_awaddr[7]), .Z(i_psram_sub_n_4265
		));
	notech_inv i_psram_sub_i_5087(.A(s00_axi_awaddr[6]), .Z(i_psram_sub_n_4264
		));
	notech_inv i_psram_sub_i_5086(.A(s00_axi_awaddr[5]), .Z(i_psram_sub_n_4263
		));
	notech_inv i_psram_sub_i_5085(.A(s00_axi_awaddr[4]), .Z(i_psram_sub_n_4262
		));
	notech_inv i_psram_sub_i_5084(.A(s00_axi_awaddr[3]), .Z(i_psram_sub_n_4261
		));
	notech_inv i_psram_sub_i_5083(.A(s00_axi_awaddr[2]), .Z(i_psram_sub_n_4260
		));
	notech_inv i_psram_sub_i_5082(.A(s00_axi_araddr[23]), .Z(i_psram_sub_n_4259
		));
	notech_inv i_psram_sub_i_5081(.A(s00_axi_araddr[22]), .Z(i_psram_sub_n_4258
		));
	notech_inv i_psram_sub_i_5080(.A(s00_axi_araddr[21]), .Z(i_psram_sub_n_4257
		));
	notech_inv i_psram_sub_i_5079(.A(s00_axi_araddr[20]), .Z(i_psram_sub_n_4256
		));
	notech_inv i_psram_sub_i_5078(.A(s00_axi_araddr[19]), .Z(i_psram_sub_n_4255
		));
	notech_inv i_psram_sub_i_5077(.A(s00_axi_araddr[18]), .Z(i_psram_sub_n_4254
		));
	notech_inv i_psram_sub_i_5076(.A(s00_axi_araddr[17]), .Z(i_psram_sub_n_4253
		));
	notech_inv i_psram_sub_i_5075(.A(s00_axi_araddr[16]), .Z(i_psram_sub_n_4252
		));
	notech_inv i_psram_sub_i_5074(.A(s00_axi_araddr[15]), .Z(i_psram_sub_n_4251
		));
	notech_inv i_psram_sub_i_5073(.A(s00_axi_araddr[14]), .Z(i_psram_sub_n_4250
		));
	notech_inv i_psram_sub_i_5072(.A(s00_axi_araddr[13]), .Z(i_psram_sub_n_4249
		));
	notech_inv i_psram_sub_i_5071(.A(s00_axi_araddr[12]), .Z(i_psram_sub_n_4248
		));
	notech_inv i_psram_sub_i_5070(.A(s00_axi_araddr[11]), .Z(i_psram_sub_n_4247
		));
	notech_inv i_psram_sub_i_5069(.A(s00_axi_araddr[10]), .Z(i_psram_sub_n_4246
		));
	notech_inv i_psram_sub_i_5068(.A(s00_axi_araddr[9]), .Z(i_psram_sub_n_4245
		));
	notech_inv i_psram_sub_i_5067(.A(s00_axi_araddr[8]), .Z(i_psram_sub_n_4244
		));
	notech_inv i_psram_sub_i_5066(.A(s00_axi_araddr[7]), .Z(i_psram_sub_n_4243
		));
	notech_inv i_psram_sub_i_5065(.A(s00_axi_araddr[6]), .Z(i_psram_sub_n_4242
		));
	notech_inv i_psram_sub_i_5064(.A(s00_axi_araddr[5]), .Z(i_psram_sub_n_4241
		));
	notech_inv i_psram_sub_i_5063(.A(s00_axi_araddr[4]), .Z(i_psram_sub_n_4240
		));
	notech_inv i_psram_sub_i_5062(.A(s00_axi_araddr[3]), .Z(i_psram_sub_n_4239
		));
	notech_inv i_psram_sub_i_5061(.A(s00_axi_araddr[2]), .Z(i_psram_sub_n_4238
		));
	notech_inv i_psram_sub_i_5060(.A(s00_axi_wdata[15]), .Z(i_psram_sub_n_4237
		));
	notech_inv i_psram_sub_i_5059(.A(s00_axi_wdata[14]), .Z(i_psram_sub_n_4236
		));
	notech_inv i_psram_sub_i_5058(.A(s00_axi_wdata[13]), .Z(i_psram_sub_n_4235
		));
	notech_inv i_psram_sub_i_5057(.A(s00_axi_wdata[12]), .Z(i_psram_sub_n_4234
		));
	notech_inv i_psram_sub_i_5056(.A(s00_axi_wdata[11]), .Z(i_psram_sub_n_4233
		));
	notech_inv i_psram_sub_i_5055(.A(s00_axi_wdata[10]), .Z(i_psram_sub_n_4232
		));
	notech_inv i_psram_sub_i_5054(.A(s00_axi_wdata[9]), .Z(i_psram_sub_n_4231
		));
	notech_inv i_psram_sub_i_5053(.A(s00_axi_wdata[8]), .Z(i_psram_sub_n_4230
		));
	notech_inv i_psram_sub_i_5052(.A(s00_axi_wdata[7]), .Z(i_psram_sub_n_4229
		));
	notech_inv i_psram_sub_i_5051(.A(s00_axi_wdata[6]), .Z(i_psram_sub_n_4228
		));
	notech_inv i_psram_sub_i_5050(.A(s00_axi_wdata[5]), .Z(i_psram_sub_n_4227
		));
	notech_inv i_psram_sub_i_5049(.A(s00_axi_wdata[4]), .Z(i_psram_sub_n_4226
		));
	notech_inv i_psram_sub_i_5048(.A(s00_axi_wdata[3]), .Z(i_psram_sub_n_4225
		));
	notech_inv i_psram_sub_i_5047(.A(s00_axi_wdata[2]), .Z(i_psram_sub_n_4224
		));
	notech_inv i_psram_sub_i_5046(.A(s00_axi_wdata[1]), .Z(i_psram_sub_n_4223
		));
	notech_inv i_psram_sub_i_5045(.A(s00_axi_wdata[0]), .Z(i_psram_sub_n_4222
		));
	notech_inv i_psram_sub_i_5044(.A(i_psram_sub_mem_addr[22]), .Z(i_psram_sub_n_4221
		));
	notech_inv i_psram_sub_i_5043(.A(i_psram_sub_mem_addr[21]), .Z(i_psram_sub_n_4220
		));
	notech_inv i_psram_sub_i_5042(.A(i_psram_sub_mem_addr[20]), .Z(i_psram_sub_n_4219
		));
	notech_inv i_psram_sub_i_5041(.A(i_psram_sub_mem_addr[19]), .Z(i_psram_sub_n_4218
		));
	notech_inv i_psram_sub_i_5040(.A(i_psram_sub_mem_addr[18]), .Z(i_psram_sub_n_4217
		));
	notech_inv i_psram_sub_i_5039(.A(i_psram_sub_mem_addr[17]), .Z(i_psram_sub_n_4216
		));
	notech_inv i_psram_sub_i_5038(.A(i_psram_sub_mem_addr[16]), .Z(i_psram_sub_n_4215
		));
	notech_inv i_psram_sub_i_5037(.A(i_psram_sub_mem_addr[15]), .Z(i_psram_sub_n_4214
		));
	notech_inv i_psram_sub_i_5036(.A(i_psram_sub_mem_addr[14]), .Z(i_psram_sub_n_4213
		));
	notech_inv i_psram_sub_i_5035(.A(i_psram_sub_mem_addr[13]), .Z(i_psram_sub_n_4212
		));
	notech_inv i_psram_sub_i_5034(.A(i_psram_sub_mem_addr[12]), .Z(i_psram_sub_n_4211
		));
	notech_inv i_psram_sub_i_5033(.A(i_psram_sub_mem_addr[11]), .Z(i_psram_sub_n_4210
		));
	notech_inv i_psram_sub_i_5032(.A(i_psram_sub_mem_addr[10]), .Z(i_psram_sub_n_4209
		));
	notech_inv i_psram_sub_i_5031(.A(i_psram_sub_mem_addr[9]), .Z(i_psram_sub_n_4208
		));
	notech_inv i_psram_sub_i_5030(.A(i_psram_sub_mem_addr[8]), .Z(i_psram_sub_n_4207
		));
	notech_inv i_psram_sub_i_5029(.A(i_psram_sub_mem_addr[7]), .Z(i_psram_sub_n_4206
		));
	notech_inv i_psram_sub_i_5028(.A(i_psram_sub_mem_addr[6]), .Z(i_psram_sub_n_4205
		));
	notech_inv i_psram_sub_i_5027(.A(i_psram_sub_mem_addr[5]), .Z(i_psram_sub_n_4204
		));
	notech_inv i_psram_sub_i_5026(.A(i_psram_sub_mem_addr[4]), .Z(i_psram_sub_n_4203
		));
	notech_inv i_psram_sub_i_5025(.A(i_psram_sub_mem_addr[3]), .Z(i_psram_sub_n_4202
		));
	notech_inv i_psram_sub_i_5024(.A(i_psram_sub_mem_addr[2]), .Z(i_psram_sub_n_4201
		));
	notech_inv i_psram_sub_i_5023(.A(i_psram_sub_mem_addr[1]), .Z(i_psram_sub_n_4200
		));
	notech_inv i_psram_sub_i_5022(.A(i_psram_sub_mem_addr[0]), .Z(i_psram_sub_n_4199
		));
	notech_inv i_psram_sub_i_5021(.A(i_psram_sub_function_plus_2[22]), .Z(i_psram_sub_n_4198
		));
	notech_inv i_psram_sub_i_5020(.A(i_psram_sub_function_plus_2[21]), .Z(i_psram_sub_n_4197
		));
	notech_inv i_psram_sub_i_5019(.A(i_psram_sub_function_plus_2[20]), .Z(i_psram_sub_n_4196
		));
	notech_inv i_psram_sub_i_5018(.A(i_psram_sub_function_plus_2[19]), .Z(i_psram_sub_n_4195
		));
	notech_inv i_psram_sub_i_5017(.A(i_psram_sub_function_plus_2[18]), .Z(i_psram_sub_n_4194
		));
	notech_inv i_psram_sub_i_5016(.A(i_psram_sub_function_plus_2[17]), .Z(i_psram_sub_n_4193
		));
	notech_inv i_psram_sub_i_5015(.A(i_psram_sub_function_plus_2[16]), .Z(i_psram_sub_n_4192
		));
	notech_inv i_psram_sub_i_5014(.A(i_psram_sub_function_plus_2[15]), .Z(i_psram_sub_n_4191
		));
	notech_inv i_psram_sub_i_5013(.A(i_psram_sub_function_plus_2[14]), .Z(i_psram_sub_n_4190
		));
	notech_inv i_psram_sub_i_5012(.A(i_psram_sub_function_plus_2[13]), .Z(i_psram_sub_n_4189
		));
	notech_inv i_psram_sub_i_5011(.A(i_psram_sub_function_plus_2[12]), .Z(i_psram_sub_n_4188
		));
	notech_inv i_psram_sub_i_5010(.A(i_psram_sub_function_plus_2[11]), .Z(i_psram_sub_n_4187
		));
	notech_inv i_psram_sub_i_5009(.A(i_psram_sub_function_plus_2[10]), .Z(i_psram_sub_n_4186
		));
	notech_inv i_psram_sub_i_5008(.A(i_psram_sub_function_plus_2[9]), .Z(i_psram_sub_n_4185
		));
	notech_inv i_psram_sub_i_5007(.A(i_psram_sub_function_plus_2[8]), .Z(i_psram_sub_n_4184
		));
	notech_inv i_psram_sub_i_5006(.A(i_psram_sub_function_plus_2[7]), .Z(i_psram_sub_n_4183
		));
	notech_inv i_psram_sub_i_5005(.A(i_psram_sub_function_plus_2[6]), .Z(i_psram_sub_n_4182
		));
	notech_inv i_psram_sub_i_5004(.A(i_psram_sub_function_plus_2[5]), .Z(i_psram_sub_n_4181
		));
	notech_inv i_psram_sub_i_5003(.A(i_psram_sub_function_plus_2[4]), .Z(i_psram_sub_n_4180
		));
	notech_inv i_psram_sub_i_5002(.A(i_psram_sub_function_plus_2[3]), .Z(i_psram_sub_n_4179
		));
	notech_inv i_psram_sub_i_5001(.A(i_psram_sub_function_plus_2[2]), .Z(i_psram_sub_n_4178
		));
	notech_inv i_psram_sub_i_5000(.A(i_psram_sub_function_plus_2[1]), .Z(i_psram_sub_n_4177
		));
	notech_inv i_psram_sub_i_4999(.A(i_psram_sub_function_plus_2[0]), .Z(i_psram_sub_n_4176
		));
	notech_inv i_psram_sub_i_4998(.A(i_psram_sub_axi_awaddr[23]), .Z(i_psram_sub_n_4175
		));
	notech_inv i_psram_sub_i_4997(.A(i_psram_sub_axi_awaddr[22]), .Z(i_psram_sub_n_4174
		));
	notech_inv i_psram_sub_i_4995(.A(i_psram_sub_axi_awaddr[21]), .Z(i_psram_sub_n_4173
		));
	notech_inv i_psram_sub_i_4994(.A(i_psram_sub_axi_awaddr[20]), .Z(i_psram_sub_n_4172
		));
	notech_inv i_psram_sub_i_4993(.A(i_psram_sub_axi_awaddr[19]), .Z(i_psram_sub_n_4171
		));
	notech_inv i_psram_sub_i_4992(.A(i_psram_sub_axi_awaddr[18]), .Z(i_psram_sub_n_4170
		));
	notech_inv i_psram_sub_i_4991(.A(i_psram_sub_axi_awaddr[17]), .Z(i_psram_sub_n_4169
		));
	notech_inv i_psram_sub_i_4990(.A(i_psram_sub_axi_awaddr[16]), .Z(i_psram_sub_n_4168
		));
	notech_inv i_psram_sub_i_4989(.A(i_psram_sub_axi_awaddr[15]), .Z(i_psram_sub_n_4167
		));
	notech_inv i_psram_sub_i_4988(.A(i_psram_sub_axi_awaddr[14]), .Z(i_psram_sub_n_4166
		));
	notech_inv i_psram_sub_i_4987(.A(i_psram_sub_axi_awaddr[13]), .Z(i_psram_sub_n_4165
		));
	notech_inv i_psram_sub_i_4986(.A(i_psram_sub_axi_awaddr[12]), .Z(i_psram_sub_n_4164
		));
	notech_inv i_psram_sub_i_4985(.A(i_psram_sub_axi_awaddr[11]), .Z(i_psram_sub_n_4163
		));
	notech_inv i_psram_sub_i_4984(.A(i_psram_sub_axi_awaddr[10]), .Z(i_psram_sub_n_4162
		));
	notech_inv i_psram_sub_i_4983(.A(i_psram_sub_axi_awaddr[9]), .Z(i_psram_sub_n_4161
		));
	notech_inv i_psram_sub_i_4982(.A(i_psram_sub_axi_awaddr[8]), .Z(i_psram_sub_n_4160
		));
	notech_inv i_psram_sub_i_4981(.A(i_psram_sub_axi_awaddr[7]), .Z(i_psram_sub_n_4159
		));
	notech_inv i_psram_sub_i_4980(.A(i_psram_sub_axi_awaddr[6]), .Z(i_psram_sub_n_4158
		));
	notech_inv i_psram_sub_i_4979(.A(i_psram_sub_axi_awaddr[5]), .Z(i_psram_sub_n_4157
		));
	notech_inv i_psram_sub_i_4978(.A(i_psram_sub_axi_awaddr[4]), .Z(i_psram_sub_n_4156
		));
	notech_inv i_psram_sub_i_4977(.A(i_psram_sub_axi_awaddr[3]), .Z(i_psram_sub_n_4155
		));
	notech_inv i_psram_sub_i_4976(.A(i_psram_sub_axi_awaddr[2]), .Z(i_psram_sub_n_4154
		));
	notech_inv i_psram_sub_i_4975(.A(i_psram_sub_axi_awaddr[1]), .Z(i_psram_sub_n_4153
		));
	notech_inv i_psram_sub_i_4974(.A(i_psram_sub_axi_awaddr[0]), .Z(i_psram_sub_n_4152
		));
	notech_inv i_psram_sub_i_4973(.A(i_psram_sub_function_sub_0[23]), .Z(i_psram_sub_n_4151
		));
	notech_inv i_psram_sub_i_4972(.A(i_psram_sub_function_sub_0[22]), .Z(i_psram_sub_n_4150
		));
	notech_inv i_psram_sub_i_4971(.A(i_psram_sub_function_sub_0[21]), .Z(i_psram_sub_n_4149
		));
	notech_inv i_psram_sub_i_4970(.A(i_psram_sub_function_sub_0[20]), .Z(i_psram_sub_n_4148
		));
	notech_inv i_psram_sub_i_4969(.A(i_psram_sub_function_sub_0[19]), .Z(i_psram_sub_n_4147
		));
	notech_inv i_psram_sub_i_4968(.A(i_psram_sub_function_sub_0[18]), .Z(i_psram_sub_n_4146
		));
	notech_inv i_psram_sub_i_4967(.A(i_psram_sub_function_sub_0[17]), .Z(i_psram_sub_n_4145
		));
	notech_inv i_psram_sub_i_4966(.A(i_psram_sub_function_sub_0[16]), .Z(i_psram_sub_n_4144
		));
	notech_inv i_psram_sub_i_4965(.A(i_psram_sub_function_sub_0[15]), .Z(i_psram_sub_n_4143
		));
	notech_inv i_psram_sub_i_4964(.A(i_psram_sub_function_sub_0[14]), .Z(i_psram_sub_n_4142
		));
	notech_inv i_psram_sub_i_4963(.A(i_psram_sub_function_sub_0[13]), .Z(i_psram_sub_n_4141
		));
	notech_inv i_psram_sub_i_4962(.A(i_psram_sub_function_sub_0[12]), .Z(i_psram_sub_n_4140
		));
	notech_inv i_psram_sub_i_4961(.A(i_psram_sub_function_sub_0[11]), .Z(i_psram_sub_n_4139
		));
	notech_inv i_psram_sub_i_4960(.A(i_psram_sub_function_sub_0[10]), .Z(i_psram_sub_n_4138
		));
	notech_inv i_psram_sub_i_4959(.A(i_psram_sub_function_sub_0[9]), .Z(i_psram_sub_n_4137
		));
	notech_inv i_psram_sub_i_4958(.A(i_psram_sub_function_sub_0[8]), .Z(i_psram_sub_n_4136
		));
	notech_inv i_psram_sub_i_4957(.A(i_psram_sub_function_sub_0[7]), .Z(i_psram_sub_n_4135
		));
	notech_inv i_psram_sub_i_4956(.A(i_psram_sub_function_sub_0[6]), .Z(i_psram_sub_n_4134
		));
	notech_inv i_psram_sub_i_4955(.A(i_psram_sub_function_sub_0[5]), .Z(i_psram_sub_n_4133
		));
	notech_inv i_psram_sub_i_4954(.A(i_psram_sub_function_sub_0[4]), .Z(i_psram_sub_n_4132
		));
	notech_inv i_psram_sub_i_4953(.A(i_psram_sub_function_sub_0[3]), .Z(i_psram_sub_n_4131
		));
	notech_inv i_psram_sub_i_4952(.A(i_psram_sub_function_sub_0[2]), .Z(i_psram_sub_n_4130
		));
	notech_inv i_psram_sub_i_4951(.A(i_psram_sub_function_sub_0[1]), .Z(i_psram_sub_n_4129
		));
	notech_inv i_psram_sub_i_4950(.A(i_psram_sub_function_sub_0[0]), .Z(i_psram_sub_n_4128
		));
	notech_inv i_psram_sub_i_4949(.A(i_psram_sub_axi_araddr[23]), .Z(i_psram_sub_n_4127
		));
	notech_inv i_psram_sub_i_4948(.A(i_psram_sub_axi_araddr[22]), .Z(i_psram_sub_n_4126
		));
	notech_inv i_psram_sub_i_4947(.A(i_psram_sub_axi_araddr[21]), .Z(i_psram_sub_n_4125
		));
	notech_inv i_psram_sub_i_4946(.A(i_psram_sub_axi_araddr[20]), .Z(i_psram_sub_n_4124
		));
	notech_inv i_psram_sub_i_4945(.A(i_psram_sub_axi_araddr[19]), .Z(i_psram_sub_n_4123
		));
	notech_inv i_psram_sub_i_4944(.A(i_psram_sub_axi_araddr[18]), .Z(i_psram_sub_n_4122
		));
	notech_inv i_psram_sub_i_4943(.A(i_psram_sub_axi_araddr[17]), .Z(i_psram_sub_n_4121
		));
	notech_inv i_psram_sub_i_4942(.A(i_psram_sub_axi_araddr[16]), .Z(i_psram_sub_n_4120
		));
	notech_inv i_psram_sub_i_4941(.A(i_psram_sub_axi_araddr[15]), .Z(i_psram_sub_n_4119
		));
	notech_inv i_psram_sub_i_4940(.A(i_psram_sub_axi_araddr[14]), .Z(i_psram_sub_n_4118
		));
	notech_inv i_psram_sub_i_4939(.A(i_psram_sub_axi_araddr[13]), .Z(i_psram_sub_n_4117
		));
	notech_inv i_psram_sub_i_4938(.A(i_psram_sub_axi_araddr[12]), .Z(i_psram_sub_n_4116
		));
	notech_inv i_psram_sub_i_4937(.A(i_psram_sub_axi_araddr[11]), .Z(i_psram_sub_n_4115
		));
	notech_inv i_psram_sub_i_4936(.A(i_psram_sub_axi_araddr[10]), .Z(i_psram_sub_n_4114
		));
	notech_inv i_psram_sub_i_4935(.A(i_psram_sub_axi_araddr[9]), .Z(i_psram_sub_n_4113
		));
	notech_inv i_psram_sub_i_4934(.A(i_psram_sub_axi_araddr[8]), .Z(i_psram_sub_n_4112
		));
	notech_inv i_psram_sub_i_4933(.A(i_psram_sub_axi_araddr[7]), .Z(i_psram_sub_n_4111
		));
	notech_inv i_psram_sub_i_4932(.A(i_psram_sub_axi_araddr[6]), .Z(i_psram_sub_n_4110
		));
	notech_inv i_psram_sub_i_4931(.A(i_psram_sub_axi_araddr[5]), .Z(i_psram_sub_n_4109
		));
	notech_inv i_psram_sub_i_4930(.A(i_psram_sub_axi_araddr[4]), .Z(i_psram_sub_n_4108
		));
	notech_inv i_psram_sub_i_4929(.A(i_psram_sub_axi_araddr[3]), .Z(i_psram_sub_n_4107
		));
	notech_inv i_psram_sub_i_4928(.A(i_psram_sub_axi_araddr[2]), .Z(i_psram_sub_n_4106
		));
	notech_inv i_psram_sub_i_4927(.A(i_psram_sub_axi_araddr[1]), .Z(i_psram_sub_n_4105
		));
	notech_inv i_psram_sub_i_4926(.A(i_psram_sub_axi_araddr[0]), .Z(i_psram_sub_n_4104
		));
	notech_inv i_psram_sub_i_4925(.A(i_psram_sub_function_sub[23]), .Z(i_psram_sub_n_4103
		));
	notech_inv i_psram_sub_i_4924(.A(i_psram_sub_function_sub[22]), .Z(i_psram_sub_n_4102
		));
	notech_inv i_psram_sub_i_4923(.A(i_psram_sub_function_sub[21]), .Z(i_psram_sub_n_4101
		));
	notech_inv i_psram_sub_i_4922(.A(i_psram_sub_function_sub[20]), .Z(i_psram_sub_n_4100
		));
	notech_inv i_psram_sub_i_4921(.A(i_psram_sub_function_sub[19]), .Z(i_psram_sub_n_4099
		));
	notech_inv i_psram_sub_i_4920(.A(i_psram_sub_function_sub[18]), .Z(i_psram_sub_n_4098
		));
	notech_inv i_psram_sub_i_4919(.A(i_psram_sub_function_sub[17]), .Z(i_psram_sub_n_4097
		));
	notech_inv i_psram_sub_i_4918(.A(i_psram_sub_function_sub[16]), .Z(i_psram_sub_n_4096
		));
	notech_inv i_psram_sub_i_4917(.A(i_psram_sub_function_sub[15]), .Z(i_psram_sub_n_4095
		));
	notech_inv i_psram_sub_i_4916(.A(i_psram_sub_function_sub[14]), .Z(i_psram_sub_n_4094
		));
	notech_inv i_psram_sub_i_4915(.A(i_psram_sub_function_sub[13]), .Z(i_psram_sub_n_4093
		));
	notech_inv i_psram_sub_i_4914(.A(i_psram_sub_function_sub[12]), .Z(i_psram_sub_n_4092
		));
	notech_inv i_psram_sub_i_4913(.A(i_psram_sub_function_sub[11]), .Z(i_psram_sub_n_4091
		));
	notech_inv i_psram_sub_i_4912(.A(i_psram_sub_function_sub[10]), .Z(i_psram_sub_n_4090
		));
	notech_inv i_psram_sub_i_4911(.A(i_psram_sub_function_sub[9]), .Z(i_psram_sub_n_4089
		));
	notech_inv i_psram_sub_i_4910(.A(i_psram_sub_function_sub[8]), .Z(i_psram_sub_n_4088
		));
	notech_inv i_psram_sub_i_4909(.A(i_psram_sub_function_sub[7]), .Z(i_psram_sub_n_4087
		));
	notech_inv i_psram_sub_i_4908(.A(i_psram_sub_function_sub[6]), .Z(i_psram_sub_n_4086
		));
	notech_inv i_psram_sub_i_4907(.A(i_psram_sub_function_sub[5]), .Z(i_psram_sub_n_4085
		));
	notech_inv i_psram_sub_i_4906(.A(i_psram_sub_function_sub[4]), .Z(i_psram_sub_n_4084
		));
	notech_inv i_psram_sub_i_4905(.A(i_psram_sub_function_sub[3]), .Z(i_psram_sub_n_4083
		));
	notech_inv i_psram_sub_i_4904(.A(i_psram_sub_function_sub[2]), .Z(i_psram_sub_n_4082
		));
	notech_inv i_psram_sub_i_4903(.A(i_psram_sub_function_sub[1]), .Z(i_psram_sub_n_4081
		));
	notech_inv i_psram_sub_i_4902(.A(i_psram_sub_function_sub[0]), .Z(i_psram_sub_n_4080
		));
	notech_inv i_psram_sub_i_4901(.A(i_psram_sub_mem_data_wr[15]), .Z(i_psram_sub_n_4079
		));
	notech_inv i_psram_sub_i_4900(.A(i_psram_sub_mem_data_wr[14]), .Z(i_psram_sub_n_4078
		));
	notech_inv i_psram_sub_i_4899(.A(i_psram_sub_mem_data_wr[13]), .Z(i_psram_sub_n_4077
		));
	notech_inv i_psram_sub_i_4898(.A(i_psram_sub_mem_data_wr[12]), .Z(i_psram_sub_n_4076
		));
	notech_inv i_psram_sub_i_4897(.A(i_psram_sub_mem_data_wr[11]), .Z(i_psram_sub_n_4075
		));
	notech_inv i_psram_sub_i_4896(.A(i_psram_sub_mem_data_wr[10]), .Z(i_psram_sub_n_4074
		));
	notech_inv i_psram_sub_i_4895(.A(i_psram_sub_mem_data_wr[9]), .Z(i_psram_sub_n_4073
		));
	notech_inv i_psram_sub_i_4894(.A(i_psram_sub_mem_data_wr[8]), .Z(i_psram_sub_n_4072
		));
	notech_inv i_psram_sub_i_4893(.A(i_psram_sub_mem_data_wr[7]), .Z(i_psram_sub_n_4071
		));
	notech_inv i_psram_sub_i_4892(.A(i_psram_sub_mem_data_wr[6]), .Z(i_psram_sub_n_4070
		));
	notech_inv i_psram_sub_i_4891(.A(i_psram_sub_mem_data_wr[5]), .Z(i_psram_sub_n_4069
		));
	notech_inv i_psram_sub_i_4890(.A(i_psram_sub_mem_data_wr[4]), .Z(i_psram_sub_n_4068
		));
	notech_inv i_psram_sub_i_4889(.A(i_psram_sub_mem_data_wr[3]), .Z(i_psram_sub_n_4067
		));
	notech_inv i_psram_sub_i_4888(.A(i_psram_sub_mem_data_wr[2]), .Z(i_psram_sub_n_4066
		));
	notech_inv i_psram_sub_i_4887(.A(i_psram_sub_mem_data_wr[1]), .Z(i_psram_sub_n_4065
		));
	notech_inv i_psram_sub_i_4886(.A(i_psram_sub_mem_data_wr[0]), .Z(i_psram_sub_n_4064
		));
	notech_inv i_psram_sub_i_4885(.A(i_psram_sub_n_1521), .Z(i_psram_sub_n_4063
		));
	notech_inv i_psram_sub_i_4884(.A(i_psram_sub_n_1516), .Z(i_psram_sub_n_4062
		));
	notech_inv i_psram_sub_i_4883(.A(i_psram_sub_n_951), .Z(i_psram_sub_n_4061
		));
	notech_inv i_psram_sub_i_4882(.A(i_psram_sub_n_1511), .Z(i_psram_sub_n_4060
		));
	notech_inv i_psram_sub_i_4881(.A(i_psram_sub_n_1506), .Z(i_psram_sub_n_4059
		));
	notech_inv i_psram_sub_i_4880(.A(i_psram_sub_n_1501), .Z(i_psram_sub_n_4058
		));
	notech_inv i_psram_sub_i_4879(.A(i_psram_sub_n_1496), .Z(i_psram_sub_n_4057
		));
	notech_inv i_psram_sub_i_4878(.A(i_psram_sub_n_1491), .Z(i_psram_sub_n_4056
		));
	notech_inv i_psram_sub_i_4877(.A(i_psram_sub_n_1486), .Z(i_psram_sub_n_4055
		));
	notech_inv i_psram_sub_i_4876(.A(i_psram_sub_n_1481), .Z(i_psram_sub_n_4054
		));
	notech_inv i_psram_sub_i_4875(.A(i_psram_sub_n_1476), .Z(i_psram_sub_n_4053
		));
	notech_inv i_psram_sub_i_4874(.A(i_psram_sub_n_1471), .Z(i_psram_sub_n_4052
		));
	notech_inv i_psram_sub_i_4873(.A(i_psram_sub_n_1466), .Z(i_psram_sub_n_4051
		));
	notech_inv i_psram_sub_i_4872(.A(i_psram_sub_n_1461), .Z(i_psram_sub_n_4050
		));
	notech_inv i_psram_sub_i_4871(.A(i_psram_sub_n_1456), .Z(i_psram_sub_n_4049
		));
	notech_inv i_psram_sub_i_4870(.A(i_psram_sub_n_1451), .Z(i_psram_sub_n_4048
		));
	notech_inv i_psram_sub_i_4869(.A(i_psram_sub_n_1446), .Z(i_psram_sub_n_4047
		));
	notech_inv i_psram_sub_i_4868(.A(i_psram_sub_n_1441), .Z(i_psram_sub_n_4046
		));
	notech_inv i_psram_sub_i_4867(.A(i_psram_sub_n_1436), .Z(i_psram_sub_n_4045
		));
	notech_inv i_psram_sub_i_4866(.A(i_psram_sub_n_1431), .Z(i_psram_sub_n_4044
		));
	notech_inv i_psram_sub_i_4865(.A(i_psram_sub_n_1426), .Z(i_psram_sub_n_4043
		));
	notech_inv i_psram_sub_i_4864(.A(i_psram_sub_n_1421), .Z(i_psram_sub_n_4042
		));
	notech_inv i_psram_sub_i_4863(.A(i_psram_sub_n_1416), .Z(i_psram_sub_n_4041
		));
	notech_inv i_psram_sub_i_4862(.A(i_psram_sub_n_1411), .Z(i_psram_sub_n_4040
		));
	notech_inv i_psram_sub_i_4861(.A(i_psram_sub_n_1406), .Z(i_psram_sub_n_4039
		));
	notech_inv i_psram_sub_i_4860(.A(i_psram_sub_n_1401), .Z(i_psram_sub_n_4038
		));
	notech_inv i_psram_sub_i_4859(.A(i_psram_sub_n_1396), .Z(i_psram_sub_n_4037
		));
	notech_inv i_psram_sub_i_4858(.A(i_psram_sub_n_1391), .Z(i_psram_sub_n_4036
		));
	notech_inv i_psram_sub_i_4857(.A(i_psram_sub_n_1386), .Z(i_psram_sub_n_4035
		));
	notech_inv i_psram_sub_i_4856(.A(i_psram_sub_n_1381), .Z(i_psram_sub_n_4034
		));
	notech_inv i_psram_sub_i_4855(.A(i_psram_sub_n_1376), .Z(i_psram_sub_n_4033
		));
	notech_inv i_psram_sub_i_4854(.A(i_psram_sub_n_1371), .Z(i_psram_sub_n_4032
		));
	notech_inv i_psram_sub_i_4853(.A(i_psram_sub_n_1366), .Z(i_psram_sub_n_4031
		));
	notech_inv i_psram_sub_i_4852(.A(i_psram_sub_n_913), .Z(i_psram_sub_n_4030
		));
	notech_inv i_psram_sub_i_4851(.A(i_psram_sub_axi_awv_awr_flag), .Z(i_psram_sub_n_4029
		));
	notech_inv i_psram_sub_i_4850(.A(i_psram_sub_n_1639), .Z(i_psram_sub_n_4028
		));
	notech_inv i_psram_sub_i_4849(.A(i_psram_sub_state[2]), .Z(i_psram_sub_n_4027
		));
	notech_inv i_psram_sub_i_4848(.A(i_psram_sub_state_5[0]), .Z(i_psram_sub_n_4026
		));
	notech_inv i_psram_sub_i_4847(.A(i_psram_sub_state[0]), .Z(i_psram_sub_n_4025
		));
	notech_inv i_psram_sub_i_4846(.A(i_psram_sub_axi_arv_arr_flag), .Z(i_psram_sub_n_4024
		));
	notech_inv i_psram_sub_i_4845(.A(i_psram_sub_axi_awlen[7]), .Z(i_psram_sub_n_4023
		));
	notech_inv i_psram_sub_i_4844(.A(i_psram_sub_axi_awlen[6]), .Z(i_psram_sub_n_4022
		));
	notech_inv i_psram_sub_i_4843(.A(i_psram_sub_axi_awlen[5]), .Z(i_psram_sub_n_4021
		));
	notech_inv i_psram_sub_i_4842(.A(i_psram_sub_axi_awlen[4]), .Z(i_psram_sub_n_4020
		));
	notech_inv i_psram_sub_i_4841(.A(i_psram_sub_axi_awlen[0]), .Z(i_psram_sub_n_4019
		));
	notech_inv i_psram_sub_i_4839(.A(i_psram_sub_axi_awlen_cntr[3]), .Z(i_psram_sub_n_4018
		));
	notech_inv i_psram_sub_i_4838(.A(i_psram_sub_axi_awlen_cntr[2]), .Z(i_psram_sub_n_4017
		));
	notech_inv i_psram_sub_i_4837(.A(i_psram_sub_n_1931), .Z(i_psram_sub_n_4016
		));
	notech_inv i_psram_sub_i_4836(.A(i_psram_sub_axi_awlen_cntr[1]), .Z(i_psram_sub_n_4015
		));
	notech_inv i_psram_sub_i_4835(.A(i_psram_sub_n_1926), .Z(i_psram_sub_n_4014
		));
	notech_inv i_psram_sub_i_4834(.A(i_psram_sub_axi_arlen[7]), .Z(i_psram_sub_n_4013
		));
	notech_inv i_psram_sub_i_4833(.A(i_psram_sub_n_799775), .Z(i_psram_sub_n_4012
		));
	notech_inv i_psram_sub_i_4832(.A(i_psram_sub_axi_arlen[6]), .Z(i_psram_sub_n_4011
		));
	notech_inv i_psram_sub_i_4831(.A(i_psram_sub_axi_arlen[5]), .Z(i_psram_sub_n_4010
		));
	notech_inv i_psram_sub_i_4830(.A(i_psram_sub_axi_arlen[4]), .Z(i_psram_sub_n_4009
		));
	notech_inv i_psram_sub_i_4829(.A(i_psram_sub_axi_arlen[0]), .Z(i_psram_sub_n_4008
		));
	notech_inv i_psram_sub_i_4828(.A(i_psram_sub_axi_arlen_cntr[3]), .Z(i_psram_sub_n_4007
		));
	notech_inv i_psram_sub_i_4827(.A(i_psram_sub_axi_arlen_cntr[2]), .Z(i_psram_sub_n_4006
		));
	notech_inv i_psram_sub_i_4826(.A(i_psram_sub_n_2072), .Z(i_psram_sub_n_4005
		));
	notech_inv i_psram_sub_i_4825(.A(i_psram_sub_axi_arlen_cntr[1]), .Z(i_psram_sub_n_4004
		));
	notech_inv i_psram_sub_i_4824(.A(i_psram_sub_n_2067), .Z(i_psram_sub_n_4003
		));
	notech_inv i_psram_sub_i_4823(.A(i_psram_sub_go_7), .Z(i_psram_sub_n_4002
		));
	notech_inv i_psram_sub_i_4822(.A(i_psram_sub_n_1015), .Z(i_psram_sub_n_4001
		));
	notech_inv i_psram_sub_i_4821(.A(i_psram_sub_n_1086), .Z(i_psram_sub_n_4000
		));
	notech_inv i_psram_sub_i_4820(.A(i_psram_sub_n_1022), .Z(i_psram_sub_n_3999
		));
	notech_inv i_psram_sub_i_4819(.A(i_psram_sub_n_1094), .Z(i_psram_sub_n_3998
		));
	notech_inv i_psram_sub_i_4818(.A(i_psram_sub_n_588), .Z(i_psram_sub_n_3997
		));
	notech_inv i_psram_sub_i_4817(.A(i_psram_sub_n_965), .Z(i_psram_sub_n_3996
		));
	notech_inv i_psram_sub_i_4816(.A(i_psram_sub_n_968), .Z(i_psram_sub_n_3995
		));
	notech_inv i_psram_sub_i_4815(.A(i_psram_sub_n_960), .Z(i_psram_sub_n_3994
		));
	notech_inv i_psram_sub_i_4814(.A(i_psram_sub_n_458), .Z(i_psram_sub_n_3993
		));
	notech_inv i_psram_sub_i_4813(.A(i_psram_sub_n_1220), .Z(i_psram_sub_n_3992
		));
	notech_inv i_psram_sub_i_4812(.A(i_psram_sub_n_1077), .Z(i_psram_sub_n_3991
		));
	notech_inv i_psram_sub_i_4811(.A(i_psram_sub_n_1006), .Z(i_psram_sub_n_3990
		));
	notech_mux2 i_psram_sub_i_3952(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[31]), .B(i_psram_sub_n_4063), .Z(i_psram_sub_n_3984));
	notech_reg_set i_psram_sub_axi_rdata_reg_31(.CP(s00_axi_aclk), .D(i_psram_sub_n_3984
		), .SD(1'b1), .Q(s00_axi_rdata[31]));
	notech_mux2 i_psram_sub_i_3944(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[30]), .B(i_psram_sub_n_4062), .Z(i_psram_sub_n_3978));
	notech_reg_set i_psram_sub_axi_rdata_reg_30(.CP(s00_axi_aclk), .D(i_psram_sub_n_3978
		), .SD(1'b1), .Q(s00_axi_rdata[30]));
	notech_ao4 i_psram_sub_i_1993(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4282
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4397), .Z(i_psram_sub_n_1366
		));
	notech_mux2 i_psram_sub_i_3936(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[29]), .B(i_psram_sub_n_4060), .Z(i_psram_sub_n_3972));
	notech_reg_set i_psram_sub_axi_rdata_reg_29(.CP(s00_axi_aclk), .D(i_psram_sub_n_3972
		), .SD(1'b1), .Q(s00_axi_rdata[29]));
	notech_ao4 i_psram_sub_i_2994(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4283
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4396), .Z(i_psram_sub_n_1371
		));
	notech_mux2 i_psram_sub_i_3928(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[28]), .B(i_psram_sub_n_4059), .Z(i_psram_sub_n_3966));
	notech_reg_set i_psram_sub_axi_rdata_reg_28(.CP(s00_axi_aclk), .D(i_psram_sub_n_3966
		), .SD(1'b1), .Q(s00_axi_rdata[28]));
	notech_ao4 i_psram_sub_i_3995(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4284
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4395), .Z(i_psram_sub_n_1376
		));
	notech_mux2 i_psram_sub_i_3920(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[27]), .B(i_psram_sub_n_4058), .Z(i_psram_sub_n_3960));
	notech_reg_set i_psram_sub_axi_rdata_reg_27(.CP(s00_axi_aclk), .D(i_psram_sub_n_3960
		), .SD(1'b1), .Q(s00_axi_rdata[27]));
	notech_ao4 i_psram_sub_i_4996(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4285
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4394), .Z(i_psram_sub_n_1381
		));
	notech_mux2 i_psram_sub_i_3912(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[26]), .B(i_psram_sub_n_4057), .Z(i_psram_sub_n_3954));
	notech_reg_set i_psram_sub_axi_rdata_reg_26(.CP(s00_axi_aclk), .D(i_psram_sub_n_3954
		), .SD(1'b1), .Q(s00_axi_rdata[26]));
	notech_ao4 i_psram_sub_i_5997(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4286
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4393), .Z(i_psram_sub_n_1386
		));
	notech_mux2 i_psram_sub_i_3904(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[25]), .B(i_psram_sub_n_4056), .Z(i_psram_sub_n_3948));
	notech_reg_set i_psram_sub_axi_rdata_reg_25(.CP(s00_axi_aclk), .D(i_psram_sub_n_3948
		), .SD(1'b1), .Q(s00_axi_rdata[25]));
	notech_ao4 i_psram_sub_i_6998(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4287
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4392), .Z(i_psram_sub_n_1391
		));
	notech_mux2 i_psram_sub_i_3895(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[24]), .B(i_psram_sub_n_4055), .Z(i_psram_sub_n_3942));
	notech_reg_set i_psram_sub_axi_rdata_reg_24(.CP(s00_axi_aclk), .D(i_psram_sub_n_3942
		), .SD(1'b1), .Q(s00_axi_rdata[24]));
	notech_ao4 i_psram_sub_i_7999(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4288
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4391), .Z(i_psram_sub_n_1396
		));
	notech_mux2 i_psram_sub_i_3887(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[23]), .B(i_psram_sub_n_4054), .Z(i_psram_sub_n_3936));
	notech_reg_set i_psram_sub_axi_rdata_reg_23(.CP(s00_axi_aclk), .D(i_psram_sub_n_3936
		), .SD(1'b1), .Q(s00_axi_rdata[23]));
	notech_ao4 i_psram_sub_i_81000(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4289
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4390), .Z(i_psram_sub_n_1401
		));
	notech_mux2 i_psram_sub_i_3879(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[22]), .B(i_psram_sub_n_4053), .Z(i_psram_sub_n_3930));
	notech_reg_set i_psram_sub_axi_rdata_reg_22(.CP(s00_axi_aclk), .D(i_psram_sub_n_3930
		), .SD(1'b1), .Q(s00_axi_rdata[22]));
	notech_ao4 i_psram_sub_i_91001(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4290
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4389), .Z(i_psram_sub_n_1406
		));
	notech_mux2 i_psram_sub_i_3871(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[21]), .B(i_psram_sub_n_4052), .Z(i_psram_sub_n_3924));
	notech_reg_set i_psram_sub_axi_rdata_reg_21(.CP(s00_axi_aclk), .D(i_psram_sub_n_3924
		), .SD(1'b1), .Q(s00_axi_rdata[21]));
	notech_ao4 i_psram_sub_i_101002(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4291
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4388), .Z(i_psram_sub_n_1411
		));
	notech_mux2 i_psram_sub_i_3863(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[20]), .B(i_psram_sub_n_4051), .Z(i_psram_sub_n_3918));
	notech_reg_set i_psram_sub_axi_rdata_reg_20(.CP(s00_axi_aclk), .D(i_psram_sub_n_3918
		), .SD(1'b1), .Q(s00_axi_rdata[20]));
	notech_ao4 i_psram_sub_i_111003(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4292
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4387), .Z(i_psram_sub_n_1416
		));
	notech_mux2 i_psram_sub_i_3855(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[19]), .B(i_psram_sub_n_4050), .Z(i_psram_sub_n_3912));
	notech_reg_set i_psram_sub_axi_rdata_reg_19(.CP(s00_axi_aclk), .D(i_psram_sub_n_3912
		), .SD(1'b1), .Q(s00_axi_rdata[19]));
	notech_ao4 i_psram_sub_i_121004(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4293
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4386), .Z(i_psram_sub_n_1421
		));
	notech_mux2 i_psram_sub_i_3847(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[18]), .B(i_psram_sub_n_4049), .Z(i_psram_sub_n_3906));
	notech_reg_set i_psram_sub_axi_rdata_reg_18(.CP(s00_axi_aclk), .D(i_psram_sub_n_3906
		), .SD(1'b1), .Q(s00_axi_rdata[18]));
	notech_ao4 i_psram_sub_i_131005(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4294
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4385), .Z(i_psram_sub_n_1426
		));
	notech_mux2 i_psram_sub_i_3838(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[17]), .B(i_psram_sub_n_4048), .Z(i_psram_sub_n_3900));
	notech_reg_set i_psram_sub_axi_rdata_reg_17(.CP(s00_axi_aclk), .D(i_psram_sub_n_3900
		), .SD(1'b1), .Q(s00_axi_rdata[17]));
	notech_ao4 i_psram_sub_i_141006(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4295
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4384), .Z(i_psram_sub_n_1431
		));
	notech_mux2 i_psram_sub_i_3830(.S(\i_psram_sub_nbus_58[16] ), .A(s00_axi_rdata
		[16]), .B(i_psram_sub_n_4047), .Z(i_psram_sub_n_3894));
	notech_reg_set i_psram_sub_axi_rdata_reg_16(.CP(s00_axi_aclk), .D(i_psram_sub_n_3894
		), .SD(1'b1), .Q(s00_axi_rdata[16]));
	notech_ao4 i_psram_sub_i_151007(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4296
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4383), .Z(i_psram_sub_n_1436
		));
	notech_mux2 i_psram_sub_i_3822(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[15]), .B(i_psram_sub_n_4046), .Z(i_psram_sub_n_3888));
	notech_reg_set i_psram_sub_axi_rdata_reg_15(.CP(s00_axi_aclk), .D(i_psram_sub_n_3888
		), .SD(1'b1), .Q(s00_axi_rdata[15]));
	notech_ao4 i_psram_sub_i_161008(.A(i_psram_sub_n_413), .B(i_psram_sub_n_4297
		), .C(i_psram_sub_n_976), .D(i_psram_sub_n_4382), .Z(i_psram_sub_n_1441
		));
	notech_mux2 i_psram_sub_i_3814(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[14]), .B(i_psram_sub_n_4045), .Z(i_psram_sub_n_3882));
	notech_reg_set i_psram_sub_axi_rdata_reg_14(.CP(s00_axi_aclk), .D(i_psram_sub_n_3882
		), .SD(1'b1), .Q(s00_axi_rdata[14]));
	notech_ao4 i_psram_sub_i_171009(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4298
		), .C(i_psram_sub_n_4397), .D(i_psram_sub_n_951), .Z(i_psram_sub_n_1446
		));
	notech_mux2 i_psram_sub_i_3806(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[13]), .B(i_psram_sub_n_4044), .Z(i_psram_sub_n_3876));
	notech_reg_set i_psram_sub_axi_rdata_reg_13(.CP(s00_axi_aclk), .D(i_psram_sub_n_3876
		), .SD(1'b1), .Q(s00_axi_rdata[13]));
	notech_ao4 i_psram_sub_i_181010(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4299
		), .C(i_psram_sub_n_951), .D(i_psram_sub_n_4396), .Z(i_psram_sub_n_1451
		));
	notech_mux2 i_psram_sub_i_3798(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[12]), .B(i_psram_sub_n_4043), .Z(i_psram_sub_n_3870));
	notech_reg_set i_psram_sub_axi_rdata_reg_12(.CP(s00_axi_aclk), .D(i_psram_sub_n_3870
		), .SD(1'b1), .Q(s00_axi_rdata[12]));
	notech_ao4 i_psram_sub_i_191011(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4300
		), .C(i_psram_sub_n_951), .D(i_psram_sub_n_4395), .Z(i_psram_sub_n_1456
		));
	notech_mux2 i_psram_sub_i_3790(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[11]), .B(i_psram_sub_n_4042), .Z(i_psram_sub_n_3864));
	notech_reg_set i_psram_sub_axi_rdata_reg_11(.CP(s00_axi_aclk), .D(i_psram_sub_n_3864
		), .SD(1'b1), .Q(s00_axi_rdata[11]));
	notech_ao4 i_psram_sub_i_201012(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4301
		), .C(i_psram_sub_n_951), .D(i_psram_sub_n_4394), .Z(i_psram_sub_n_1461
		));
	notech_mux2 i_psram_sub_i_3782(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[10]), .B(i_psram_sub_n_4041), .Z(i_psram_sub_n_3858));
	notech_reg_set i_psram_sub_axi_rdata_reg_10(.CP(s00_axi_aclk), .D(i_psram_sub_n_3858
		), .SD(1'b1), .Q(s00_axi_rdata[10]));
	notech_ao4 i_psram_sub_i_211013(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4302
		), .C(i_psram_sub_n_951), .D(i_psram_sub_n_4393), .Z(i_psram_sub_n_1466
		));
	notech_mux2 i_psram_sub_i_3774(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[9]), .B(i_psram_sub_n_4040), .Z(i_psram_sub_n_3852));
	notech_reg_set i_psram_sub_axi_rdata_reg_9(.CP(s00_axi_aclk), .D(i_psram_sub_n_3852
		), .SD(1'b1), .Q(s00_axi_rdata[9]));
	notech_ao4 i_psram_sub_i_221014(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4303
		), .C(i_psram_sub_n_951), .D(i_psram_sub_n_4392), .Z(i_psram_sub_n_1471
		));
	notech_mux2 i_psram_sub_i_3765(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[8]), .B(i_psram_sub_n_4039), .Z(i_psram_sub_n_3846));
	notech_reg_set i_psram_sub_axi_rdata_reg_8(.CP(s00_axi_aclk), .D(i_psram_sub_n_3846
		), .SD(1'b1), .Q(s00_axi_rdata[8]));
	notech_ao4 i_psram_sub_i_231015(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4304
		), .C(i_psram_sub_n_951), .D(i_psram_sub_n_4391), .Z(i_psram_sub_n_1476
		));
	notech_mux2 i_psram_sub_i_3757(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[7]), .B(i_psram_sub_n_4038), .Z(i_psram_sub_n_3840));
	notech_reg_set i_psram_sub_axi_rdata_reg_7(.CP(s00_axi_aclk), .D(i_psram_sub_n_3840
		), .SD(1'b1), .Q(s00_axi_rdata[7]));
	notech_ao4 i_psram_sub_i_241016(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4305
		), .C(i_psram_sub_n_4390), .D(i_psram_sub_n_951), .Z(i_psram_sub_n_1481
		));
	notech_mux2 i_psram_sub_i_3749(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[6]), .B(i_psram_sub_n_4037), .Z(i_psram_sub_n_3834));
	notech_reg_set i_psram_sub_axi_rdata_reg_6(.CP(s00_axi_aclk), .D(i_psram_sub_n_3834
		), .SD(1'b1), .Q(s00_axi_rdata[6]));
	notech_ao4 i_psram_sub_i_251017(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4306
		), .C(i_psram_sub_n_4389), .D(i_psram_sub_n_951), .Z(i_psram_sub_n_1486
		));
	notech_mux2 i_psram_sub_i_3741(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[5]), .B(i_psram_sub_n_4036), .Z(i_psram_sub_n_3828));
	notech_reg_set i_psram_sub_axi_rdata_reg_5(.CP(s00_axi_aclk), .D(i_psram_sub_n_3828
		), .SD(1'b1), .Q(s00_axi_rdata[5]));
	notech_ao4 i_psram_sub_i_261018(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4307
		), .C(i_psram_sub_n_4388), .D(i_psram_sub_n_951), .Z(i_psram_sub_n_1491
		));
	notech_mux2 i_psram_sub_i_3733(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[4]), .B(i_psram_sub_n_4035), .Z(i_psram_sub_n_3822));
	notech_reg_set i_psram_sub_axi_rdata_reg_4(.CP(s00_axi_aclk), .D(i_psram_sub_n_3822
		), .SD(1'b1), .Q(s00_axi_rdata[4]));
	notech_ao4 i_psram_sub_i_271019(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4308
		), .C(i_psram_sub_n_4387), .D(i_psram_sub_n_951), .Z(i_psram_sub_n_1496
		));
	notech_mux2 i_psram_sub_i_3725(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[3]), .B(i_psram_sub_n_4034), .Z(i_psram_sub_n_3816));
	notech_reg_set i_psram_sub_axi_rdata_reg_3(.CP(s00_axi_aclk), .D(i_psram_sub_n_3816
		), .SD(1'b1), .Q(s00_axi_rdata[3]));
	notech_ao4 i_psram_sub_i_281020(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4309
		), .C(i_psram_sub_n_4386), .D(i_psram_sub_n_951), .Z(i_psram_sub_n_1501
		));
	notech_mux2 i_psram_sub_i_3717(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[2]), .B(i_psram_sub_n_4033), .Z(i_psram_sub_n_3810));
	notech_reg_set i_psram_sub_axi_rdata_reg_2(.CP(s00_axi_aclk), .D(i_psram_sub_n_3810
		), .SD(1'b1), .Q(s00_axi_rdata[2]));
	notech_ao4 i_psram_sub_i_291021(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4310
		), .C(i_psram_sub_n_4385), .D(i_psram_sub_n_951), .Z(i_psram_sub_n_1506
		));
	notech_mux2 i_psram_sub_i_3709(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[1]), .B(i_psram_sub_n_4032), .Z(i_psram_sub_n_3804));
	notech_reg_set i_psram_sub_axi_rdata_reg_1(.CP(s00_axi_aclk), .D(i_psram_sub_n_3804
		), .SD(1'b1), .Q(s00_axi_rdata[1]));
	notech_ao4 i_psram_sub_i_301022(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4311
		), .C(i_psram_sub_n_4384), .D(i_psram_sub_n_951), .Z(i_psram_sub_n_1511
		));
	notech_mux2 i_psram_sub_i_3701(.S(\i_psram_sub_nbus_58[0] ), .A(s00_axi_rdata
		[0]), .B(i_psram_sub_n_4031), .Z(i_psram_sub_n_3798));
	notech_reg_set i_psram_sub_axi_rdata_reg_0(.CP(s00_axi_aclk), .D(i_psram_sub_n_3798
		), .SD(1'b1), .Q(s00_axi_rdata[0]));
	notech_ao4 i_psram_sub_i_311023(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4312
		), .C(i_psram_sub_n_4383), .D(i_psram_sub_n_951), .Z(i_psram_sub_n_1516
		));
	notech_and3 i_psram_sub_i_3694(.A(s00_axi_aresetn), .B(i_psram_sub_n_569
		), .C(s00_axi_bresp[1]), .Z(i_psram_sub_n_3795));
	notech_reg_set i_psram_sub_axi_bresp_reg_1(.CP(s00_axi_aclk), .D(i_psram_sub_n_3795
		), .SD(1'b1), .Q(s00_axi_bresp[1]));
	notech_ao4 i_psram_sub_i_321024(.A(i_psram_sub_n_448), .B(i_psram_sub_n_4313
		), .C(i_psram_sub_n_4382), .D(i_psram_sub_n_951), .Z(i_psram_sub_n_1521
		));
	notech_and3 i_psram_sub_i_3686(.A(s00_axi_aresetn), .B(s00_axi_bresp[0])
		, .C(i_psram_sub_n_569), .Z(i_psram_sub_n_3789));
	notech_reg_set i_psram_sub_axi_bresp_reg_0(.CP(s00_axi_aclk), .D(i_psram_sub_n_3789
		), .SD(1'b1), .Q(s00_axi_bresp[0]));
	notech_nand3 i_psram_sub_i_1379(.A(i_psram_sub_n_1198), .B(i_psram_sub_n_1202
		), .C(i_psram_sub_n_593), .Z(i_psram_sub_n_2037));
	notech_nao3 i_psram_sub_i_3678(.A(s00_axi_bvalid), .B(\i_psram_sub_nbus_68[0] 
		), .C(s00_axi_bready), .Z(i_psram_sub_n_3783));
	notech_nao3 i_psram_sub_i_3677(.A(s00_axi_aresetn), .B(i_psram_sub_n_2024
		), .C(s00_axi_bvalid), .Z(i_psram_sub_n_3782));
	notech_nand2 i_psram_sub_i_3676(.A(i_psram_sub_n_3782), .B(i_psram_sub_n_3783
		), .Z(i_psram_sub_n_3780));
	notech_reg_set i_psram_sub_axi_bvalid_reg(.CP(s00_axi_aclk), .D(i_psram_sub_n_3780
		), .SD(1'b1), .Q(s00_axi_bvalid));
	notech_nand3 i_psram_sub_i_2380(.A(i_psram_sub_n_1198), .B(i_psram_sub_n_1196
		), .C(i_psram_sub_n_597), .Z(i_psram_sub_n_2042));
	notech_mux2 i_psram_sub_i_3668(.S(i_psram_sub_n_2173), .A(s00_axi_rlast)
		, .B(i_psram_sub_n_579), .Z(i_psram_sub_n_3774));
	notech_reg_set i_psram_sub_axi_rlast_reg(.CP(s00_axi_aclk), .D(i_psram_sub_n_3774
		), .SD(1'b1), .Q(s00_axi_rlast));
	notech_nand2 i_psram_sub_i_1694(.A(i_psram_sub_n_1194), .B(i_psram_sub_n_1193
		), .Z(i_psram_sub_n_1237));
	notech_and3 i_psram_sub_i_3662(.A(s00_axi_aresetn), .B(i_psram_sub_n_568
		), .C(s00_axi_rresp[1]), .Z(i_psram_sub_n_3771));
	notech_reg_set i_psram_sub_axi_rresp_reg_1(.CP(s00_axi_aclk), .D(i_psram_sub_n_3771
		), .SD(1'b1), .Q(s00_axi_rresp[1]));
	notech_nand2 i_psram_sub_i_2695(.A(i_psram_sub_n_1192), .B(i_psram_sub_n_1191
		), .Z(i_psram_sub_n_1242));
	notech_and3 i_psram_sub_i_3654(.A(s00_axi_aresetn), .B(s00_axi_rresp[0])
		, .C(i_psram_sub_n_568), .Z(i_psram_sub_n_3765));
	notech_reg_set i_psram_sub_axi_rresp_reg_0(.CP(s00_axi_aclk), .D(i_psram_sub_n_3765
		), .SD(1'b1), .Q(s00_axi_rresp[0]));
	notech_nand2 i_psram_sub_i_3696(.A(i_psram_sub_n_1190), .B(i_psram_sub_n_1189
		), .Z(i_psram_sub_n_1247));
	notech_mux2 i_psram_sub_i_3644(.S(i_psram_sub_n_2198), .A(s00_axi_awready
		), .B(i_psram_sub_n_580), .Z(i_psram_sub_n_3756));
	notech_reg_set i_psram_sub_axi_awready_reg(.CP(s00_axi_aclk), .D(i_psram_sub_n_3756
		), .SD(1'b1), .Q(s00_axi_awready));
	notech_nand2 i_psram_sub_i_4697(.A(i_psram_sub_n_1188), .B(i_psram_sub_n_1187
		), .Z(i_psram_sub_n_1252));
	notech_mux2 i_psram_sub_i_3636(.S(i_psram_sub_n_1786), .A(i_psram_sub_axi_awv_awr_flag
		), .B(i_psram_sub_n_580), .Z(i_psram_sub_n_3750));
	notech_reg_set i_psram_sub_axi_awv_awr_flag_reg(.CP(s00_axi_aclk), .D(i_psram_sub_n_3750
		), .SD(1'b1), .Q(i_psram_sub_axi_awv_awr_flag));
	notech_nand2 i_psram_sub_i_5698(.A(i_psram_sub_n_1186), .B(i_psram_sub_n_1185
		), .Z(i_psram_sub_n_1257));
	notech_mux2 i_psram_sub_i_3628(.S(\i_psram_sub_nbus_56[0] ), .A(s00_axi_wready
		), .B(i_psram_sub_n_4028), .Z(i_psram_sub_n_3744));
	notech_reg_set i_psram_sub_axi_wready_reg(.CP(s00_axi_aclk), .D(i_psram_sub_n_3744
		), .SD(1'b1), .Q(s00_axi_wready));
	notech_reg_set i_psram_sub_state_reg_2(.CP(s00_axi_aclk), .D(i_psram_sub_state_5
		[2]), .SD(1'b1), .Q(i_psram_sub_state[2]));
	notech_reg_set i_psram_sub_state_reg_1(.CP(s00_axi_aclk), .D(i_psram_sub_state_5
		[1]), .SD(1'b1), .Q(i_psram_sub_state[1]));
	notech_reg_set i_psram_sub_state_reg_0(.CP(s00_axi_aclk), .D(i_psram_sub_n_4026
		), .SD(1'b1), .Q(i_psram_sub_state[0]));
	notech_nand2 i_psram_sub_i_6699(.A(i_psram_sub_n_1184), .B(i_psram_sub_n_1183
		), .Z(i_psram_sub_n_1262));
	notech_mux2 i_psram_sub_i_3608(.S(i_psram_sub_n_2159), .A(i_psram_sub_axi_arv_arr_flag
		), .B(i_psram_sub_n_581), .Z(i_psram_sub_n_3732));
	notech_reg_set i_psram_sub_axi_arv_arr_flag_reg(.CP(s00_axi_aclk), .D(i_psram_sub_n_3732
		), .SD(1'b1), .Q(i_psram_sub_axi_arv_arr_flag));
	notech_nand2 i_psram_sub_i_7700(.A(i_psram_sub_n_1182), .B(i_psram_sub_n_1181
		), .Z(i_psram_sub_n_1267));
	notech_mux2 i_psram_sub_i_3600(.S(i_psram_sub_n_1970), .A(s00_axi_arready
		), .B(i_psram_sub_n_581), .Z(i_psram_sub_n_3726));
	notech_reg_set i_psram_sub_axi_arready_reg(.CP(s00_axi_aclk), .D(i_psram_sub_n_3726
		), .SD(1'b1), .Q(s00_axi_arready));
	notech_reg_set i_psram_sub_axi_rvalid_reg(.CP(s00_axi_aclk), .D(i_psram_sub_n_4061
		), .SD(1'b1), .Q(s00_axi_rvalid));
	notech_nand2 i_psram_sub_i_8701(.A(i_psram_sub_n_1180), .B(i_psram_sub_n_1179
		), .Z(i_psram_sub_n_1272));
	notech_mux2 i_psram_sub_i_3588(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_command
		), .B(i_psram_sub_n_2054), .Z(i_psram_sub_n_3718));
	notech_reg_set i_psram_sub_command_reg(.CP(s00_axi_aclk), .D(i_psram_sub_n_3718
		), .SD(1'b1), .Q(i_psram_sub_command));
	notech_nand2 i_psram_sub_i_9702(.A(i_psram_sub_n_1178), .B(i_psram_sub_n_1177
		), .Z(i_psram_sub_n_1277));
	notech_mux2 i_psram_sub_i_3580(.S(\i_psram_sub_nbus_64[0] ), .A(i_psram_sub_mem_byte_en
		[1]), .B(i_psram_sub_n_2042), .Z(i_psram_sub_n_3712));
	notech_reg_set i_psram_sub_mem_byte_en_reg_1(.CP(s00_axi_aclk), .D(i_psram_sub_n_3712
		), .SD(1'b1), .Q(i_psram_sub_mem_byte_en[1]));
	notech_nand2 i_psram_sub_i_10703(.A(i_psram_sub_n_1176), .B(i_psram_sub_n_1175
		), .Z(i_psram_sub_n_1282));
	notech_mux2 i_psram_sub_i_3572(.S(\i_psram_sub_nbus_64[0] ), .A(i_psram_sub_mem_byte_en
		[0]), .B(i_psram_sub_n_2037), .Z(i_psram_sub_n_3706));
	notech_reg_set i_psram_sub_mem_byte_en_reg_0(.CP(s00_axi_aclk), .D(i_psram_sub_n_3706
		), .SD(1'b1), .Q(i_psram_sub_mem_byte_en[0]));
	notech_nand2 i_psram_sub_i_11704(.A(i_psram_sub_n_1174), .B(i_psram_sub_n_1173
		), .Z(i_psram_sub_n_1287));
	notech_mux2 i_psram_sub_i_3564(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[22]), .B(i_psram_sub_n_1347), .Z(i_psram_sub_n_3700));
	notech_reg_set i_psram_sub_mem_addr_reg_22(.CP(s00_axi_aclk), .D(i_psram_sub_n_3700
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[22]));
	notech_nand2 i_psram_sub_i_12705(.A(i_psram_sub_n_1172), .B(i_psram_sub_n_1171
		), .Z(i_psram_sub_n_1292));
	notech_mux2 i_psram_sub_i_3556(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[21]), .B(i_psram_sub_n_1342), .Z(i_psram_sub_n_3694));
	notech_reg_set i_psram_sub_mem_addr_reg_21(.CP(s00_axi_aclk), .D(i_psram_sub_n_3694
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[21]));
	notech_nand2 i_psram_sub_i_13706(.A(i_psram_sub_n_1170), .B(i_psram_sub_n_1169
		), .Z(i_psram_sub_n_1297));
	notech_mux2 i_psram_sub_i_3548(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[20]), .B(i_psram_sub_n_1337), .Z(i_psram_sub_n_3688));
	notech_reg_set i_psram_sub_mem_addr_reg_20(.CP(s00_axi_aclk), .D(i_psram_sub_n_3688
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[20]));
	notech_nand2 i_psram_sub_i_14707(.A(i_psram_sub_n_1168), .B(i_psram_sub_n_1167
		), .Z(i_psram_sub_n_1302));
	notech_mux2 i_psram_sub_i_3540(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[19]), .B(i_psram_sub_n_1332), .Z(i_psram_sub_n_3682));
	notech_reg_set i_psram_sub_mem_addr_reg_19(.CP(s00_axi_aclk), .D(i_psram_sub_n_3682
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[19]));
	notech_nand2 i_psram_sub_i_15708(.A(i_psram_sub_n_1166), .B(i_psram_sub_n_1165
		), .Z(i_psram_sub_n_1307));
	notech_mux2 i_psram_sub_i_3532(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[18]), .B(i_psram_sub_n_1327), .Z(i_psram_sub_n_3676));
	notech_reg_set i_psram_sub_mem_addr_reg_18(.CP(s00_axi_aclk), .D(i_psram_sub_n_3676
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[18]));
	notech_nand2 i_psram_sub_i_16709(.A(i_psram_sub_n_1164), .B(i_psram_sub_n_1163
		), .Z(i_psram_sub_n_1312));
	notech_mux2 i_psram_sub_i_3524(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[17]), .B(i_psram_sub_n_1322), .Z(i_psram_sub_n_3670));
	notech_reg_set i_psram_sub_mem_addr_reg_17(.CP(s00_axi_aclk), .D(i_psram_sub_n_3670
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[17]));
	notech_nand2 i_psram_sub_i_17710(.A(i_psram_sub_n_1162), .B(i_psram_sub_n_1161
		), .Z(i_psram_sub_n_1317));
	notech_mux2 i_psram_sub_i_3516(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[16]), .B(i_psram_sub_n_1317), .Z(i_psram_sub_n_3664));
	notech_reg_set i_psram_sub_mem_addr_reg_16(.CP(s00_axi_aclk), .D(i_psram_sub_n_3664
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[16]));
	notech_nand2 i_psram_sub_i_18711(.A(i_psram_sub_n_1160), .B(i_psram_sub_n_1159
		), .Z(i_psram_sub_n_1322));
	notech_mux2 i_psram_sub_i_3508(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[15]), .B(i_psram_sub_n_1312), .Z(i_psram_sub_n_3658));
	notech_reg_set i_psram_sub_mem_addr_reg_15(.CP(s00_axi_aclk), .D(i_psram_sub_n_3658
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[15]));
	notech_nand2 i_psram_sub_i_19712(.A(i_psram_sub_n_1158), .B(i_psram_sub_n_1157
		), .Z(i_psram_sub_n_1327));
	notech_mux2 i_psram_sub_i_3500(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[14]), .B(i_psram_sub_n_1307), .Z(i_psram_sub_n_3652));
	notech_reg_set i_psram_sub_mem_addr_reg_14(.CP(s00_axi_aclk), .D(i_psram_sub_n_3652
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[14]));
	notech_nand2 i_psram_sub_i_20713(.A(i_psram_sub_n_1156), .B(i_psram_sub_n_1155
		), .Z(i_psram_sub_n_1332));
	notech_mux2 i_psram_sub_i_3492(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[13]), .B(i_psram_sub_n_1302), .Z(i_psram_sub_n_3646));
	notech_reg_set i_psram_sub_mem_addr_reg_13(.CP(s00_axi_aclk), .D(i_psram_sub_n_3646
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[13]));
	notech_nand2 i_psram_sub_i_21714(.A(i_psram_sub_n_1154), .B(i_psram_sub_n_1153
		), .Z(i_psram_sub_n_1337));
	notech_mux2 i_psram_sub_i_3484(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[12]), .B(i_psram_sub_n_1297), .Z(i_psram_sub_n_3640));
	notech_reg_set i_psram_sub_mem_addr_reg_12(.CP(s00_axi_aclk), .D(i_psram_sub_n_3640
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[12]));
	notech_nand2 i_psram_sub_i_22715(.A(i_psram_sub_n_1152), .B(i_psram_sub_n_1151
		), .Z(i_psram_sub_n_1342));
	notech_mux2 i_psram_sub_i_3476(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[11]), .B(i_psram_sub_n_1292), .Z(i_psram_sub_n_3634));
	notech_reg_set i_psram_sub_mem_addr_reg_11(.CP(s00_axi_aclk), .D(i_psram_sub_n_3634
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[11]));
	notech_nand2 i_psram_sub_i_23716(.A(i_psram_sub_n_1150), .B(i_psram_sub_n_1148
		), .Z(i_psram_sub_n_1347));
	notech_mux2 i_psram_sub_i_3468(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[10]), .B(i_psram_sub_n_1287), .Z(i_psram_sub_n_3628));
	notech_reg_set i_psram_sub_mem_addr_reg_10(.CP(s00_axi_aclk), .D(i_psram_sub_n_3628
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[10]));
	notech_nand2 i_psram_sub_i_1837(.A(i_psram_sub_n_1147), .B(i_psram_sub_n_460
		), .Z(i_psram_sub_n_1660));
	notech_mux2 i_psram_sub_i_3460(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[9]), .B(i_psram_sub_n_1282), .Z(i_psram_sub_n_3622));
	notech_reg_set i_psram_sub_mem_addr_reg_9(.CP(s00_axi_aclk), .D(i_psram_sub_n_3622
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[9]));
	notech_nand2 i_psram_sub_i_2838(.A(i_psram_sub_n_1146), .B(i_psram_sub_n_461
		), .Z(i_psram_sub_n_1665));
	notech_mux2 i_psram_sub_i_3452(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[8]), .B(i_psram_sub_n_1277), .Z(i_psram_sub_n_3616));
	notech_reg_set i_psram_sub_mem_addr_reg_8(.CP(s00_axi_aclk), .D(i_psram_sub_n_3616
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[8]));
	notech_nand2 i_psram_sub_i_3839(.A(i_psram_sub_n_1145), .B(i_psram_sub_n_1144
		), .Z(i_psram_sub_n_1670));
	notech_mux2 i_psram_sub_i_3444(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[7]), .B(i_psram_sub_n_1272), .Z(i_psram_sub_n_3610));
	notech_reg_set i_psram_sub_mem_addr_reg_7(.CP(s00_axi_aclk), .D(i_psram_sub_n_3610
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[7]));
	notech_nand2 i_psram_sub_i_4840(.A(i_psram_sub_n_1143), .B(i_psram_sub_n_1142
		), .Z(i_psram_sub_n_1675));
	notech_mux2 i_psram_sub_i_3436(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[6]), .B(i_psram_sub_n_1267), .Z(i_psram_sub_n_3604));
	notech_reg_set i_psram_sub_mem_addr_reg_6(.CP(s00_axi_aclk), .D(i_psram_sub_n_3604
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[6]));
	notech_nand2 i_psram_sub_i_5841(.A(i_psram_sub_n_1141), .B(i_psram_sub_n_1140
		), .Z(i_psram_sub_n_1680));
	notech_mux2 i_psram_sub_i_3428(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[5]), .B(i_psram_sub_n_1262), .Z(i_psram_sub_n_3598));
	notech_reg_set i_psram_sub_mem_addr_reg_5(.CP(s00_axi_aclk), .D(i_psram_sub_n_3598
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[5]));
	notech_nand2 i_psram_sub_i_6842(.A(i_psram_sub_n_1139), .B(i_psram_sub_n_1138
		), .Z(i_psram_sub_n_1685));
	notech_mux2 i_psram_sub_i_3420(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[4]), .B(i_psram_sub_n_1257), .Z(i_psram_sub_n_3592));
	notech_reg_set i_psram_sub_mem_addr_reg_4(.CP(s00_axi_aclk), .D(i_psram_sub_n_3592
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[4]));
	notech_nand2 i_psram_sub_i_7843(.A(i_psram_sub_n_1137), .B(i_psram_sub_n_1136
		), .Z(i_psram_sub_n_1690));
	notech_mux2 i_psram_sub_i_3412(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[3]), .B(i_psram_sub_n_1252), .Z(i_psram_sub_n_3586));
	notech_reg_set i_psram_sub_mem_addr_reg_3(.CP(s00_axi_aclk), .D(i_psram_sub_n_3586
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[3]));
	notech_nand2 i_psram_sub_i_8844(.A(i_psram_sub_n_1135), .B(i_psram_sub_n_1134
		), .Z(i_psram_sub_n_1695));
	notech_mux2 i_psram_sub_i_3404(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[2]), .B(i_psram_sub_n_1247), .Z(i_psram_sub_n_3580));
	notech_reg_set i_psram_sub_mem_addr_reg_2(.CP(s00_axi_aclk), .D(i_psram_sub_n_3580
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[2]));
	notech_nand2 i_psram_sub_i_9845(.A(i_psram_sub_n_1133), .B(i_psram_sub_n_1132
		), .Z(i_psram_sub_n_1700));
	notech_mux2 i_psram_sub_i_3396(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[1]), .B(i_psram_sub_n_1242), .Z(i_psram_sub_n_3574));
	notech_reg_set i_psram_sub_mem_addr_reg_1(.CP(s00_axi_aclk), .D(i_psram_sub_n_3574
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[1]));
	notech_nand2 i_psram_sub_i_10846(.A(i_psram_sub_n_1131), .B(i_psram_sub_n_1130
		), .Z(i_psram_sub_n_1705));
	notech_mux2 i_psram_sub_i_3388(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_addr
		[0]), .B(i_psram_sub_n_1237), .Z(i_psram_sub_n_3568));
	notech_reg_set i_psram_sub_mem_addr_reg_0(.CP(s00_axi_aclk), .D(i_psram_sub_n_3568
		), .SD(1'b1), .Q(i_psram_sub_mem_addr[0]));
	notech_nand2 i_psram_sub_i_11847(.A(i_psram_sub_n_1129), .B(i_psram_sub_n_1128
		), .Z(i_psram_sub_n_1710));
	notech_mux2 i_psram_sub_i_3380(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[23]), .B(i_psram_sub_n_1775), .Z(i_psram_sub_n_3562));
	notech_reg_set i_psram_sub_axi_awaddr_reg_23(.CP(s00_axi_aclk), .D(i_psram_sub_n_3562
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[23]));
	notech_nand2 i_psram_sub_i_12848(.A(i_psram_sub_n_1127), .B(i_psram_sub_n_1126
		), .Z(i_psram_sub_n_1715));
	notech_mux2 i_psram_sub_i_3372(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[22]), .B(i_psram_sub_n_1770), .Z(i_psram_sub_n_3556));
	notech_reg_set i_psram_sub_axi_awaddr_reg_22(.CP(s00_axi_aclk), .D(i_psram_sub_n_3556
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[22]));
	notech_nand2 i_psram_sub_i_13849(.A(i_psram_sub_n_1125), .B(i_psram_sub_n_1124
		), .Z(i_psram_sub_n_1720));
	notech_mux2 i_psram_sub_i_3364(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[21]), .B(i_psram_sub_n_1765), .Z(i_psram_sub_n_3550));
	notech_reg_set i_psram_sub_axi_awaddr_reg_21(.CP(s00_axi_aclk), .D(i_psram_sub_n_3550
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[21]));
	notech_nand2 i_psram_sub_i_14850(.A(i_psram_sub_n_1123), .B(i_psram_sub_n_1122
		), .Z(i_psram_sub_n_1725));
	notech_mux2 i_psram_sub_i_3356(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[20]), .B(i_psram_sub_n_1760), .Z(i_psram_sub_n_3544));
	notech_reg_set i_psram_sub_axi_awaddr_reg_20(.CP(s00_axi_aclk), .D(i_psram_sub_n_3544
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[20]));
	notech_nand2 i_psram_sub_i_15851(.A(i_psram_sub_n_1121), .B(i_psram_sub_n_1120
		), .Z(i_psram_sub_n_1730));
	notech_mux2 i_psram_sub_i_3348(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[19]), .B(i_psram_sub_n_1755), .Z(i_psram_sub_n_3538));
	notech_reg_set i_psram_sub_axi_awaddr_reg_19(.CP(s00_axi_aclk), .D(i_psram_sub_n_3538
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[19]));
	notech_nand2 i_psram_sub_i_16852(.A(i_psram_sub_n_1119), .B(i_psram_sub_n_1118
		), .Z(i_psram_sub_n_1735));
	notech_mux2 i_psram_sub_i_3340(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[18]), .B(i_psram_sub_n_1750), .Z(i_psram_sub_n_3532));
	notech_reg_set i_psram_sub_axi_awaddr_reg_18(.CP(s00_axi_aclk), .D(i_psram_sub_n_3532
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[18]));
	notech_nand2 i_psram_sub_i_17853(.A(i_psram_sub_n_1117), .B(i_psram_sub_n_1116
		), .Z(i_psram_sub_n_1740));
	notech_mux2 i_psram_sub_i_3332(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[17]), .B(i_psram_sub_n_1745), .Z(i_psram_sub_n_3526));
	notech_reg_set i_psram_sub_axi_awaddr_reg_17(.CP(s00_axi_aclk), .D(i_psram_sub_n_3526
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[17]));
	notech_nand2 i_psram_sub_i_18854(.A(i_psram_sub_n_1115), .B(i_psram_sub_n_1114
		), .Z(i_psram_sub_n_1745));
	notech_mux2 i_psram_sub_i_3323(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[16]), .B(i_psram_sub_n_1740), .Z(i_psram_sub_n_3520));
	notech_reg_set i_psram_sub_axi_awaddr_reg_16(.CP(s00_axi_aclk), .D(i_psram_sub_n_3520
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[16]));
	notech_nand2 i_psram_sub_i_19855(.A(i_psram_sub_n_1113), .B(i_psram_sub_n_1112
		), .Z(i_psram_sub_n_1750));
	notech_mux2 i_psram_sub_i_3315(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[15]), .B(i_psram_sub_n_1735), .Z(i_psram_sub_n_3514));
	notech_reg_set i_psram_sub_axi_awaddr_reg_15(.CP(s00_axi_aclk), .D(i_psram_sub_n_3514
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[15]));
	notech_nand2 i_psram_sub_i_20856(.A(i_psram_sub_n_1111), .B(i_psram_sub_n_1110
		), .Z(i_psram_sub_n_1755));
	notech_mux2 i_psram_sub_i_3307(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[14]), .B(i_psram_sub_n_1730), .Z(i_psram_sub_n_3508));
	notech_reg_set i_psram_sub_axi_awaddr_reg_14(.CP(s00_axi_aclk), .D(i_psram_sub_n_3508
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[14]));
	notech_nand2 i_psram_sub_i_21857(.A(i_psram_sub_n_1109), .B(i_psram_sub_n_1108
		), .Z(i_psram_sub_n_1760));
	notech_mux2 i_psram_sub_i_3299(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[13]), .B(i_psram_sub_n_1725), .Z(i_psram_sub_n_3502));
	notech_reg_set i_psram_sub_axi_awaddr_reg_13(.CP(s00_axi_aclk), .D(i_psram_sub_n_3502
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[13]));
	notech_nand2 i_psram_sub_i_22858(.A(i_psram_sub_n_1107), .B(i_psram_sub_n_1106
		), .Z(i_psram_sub_n_1765));
	notech_mux2 i_psram_sub_i_3291(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[12]), .B(i_psram_sub_n_1720), .Z(i_psram_sub_n_3496));
	notech_reg_set i_psram_sub_axi_awaddr_reg_12(.CP(s00_axi_aclk), .D(i_psram_sub_n_3496
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[12]));
	notech_nand2 i_psram_sub_i_23859(.A(i_psram_sub_n_1105), .B(i_psram_sub_n_1104
		), .Z(i_psram_sub_n_1770));
	notech_mux2 i_psram_sub_i_3283(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[11]), .B(i_psram_sub_n_1715), .Z(i_psram_sub_n_3490));
	notech_reg_set i_psram_sub_axi_awaddr_reg_11(.CP(s00_axi_aclk), .D(i_psram_sub_n_3490
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[11]));
	notech_nand2 i_psram_sub_i_24860(.A(i_psram_sub_n_1103), .B(i_psram_sub_n_1098
		), .Z(i_psram_sub_n_1775));
	notech_mux2 i_psram_sub_i_3275(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[10]), .B(i_psram_sub_n_1710), .Z(i_psram_sub_n_3484));
	notech_reg_set i_psram_sub_axi_awaddr_reg_10(.CP(s00_axi_aclk), .D(i_psram_sub_n_3484
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[10]));
	notech_ao4 i_psram_sub_i_21066(.A(i_psram_sub_n_4015), .B(i_psram_sub_n_799775
		), .C(\i_psram_sub_nbus_63[0] ), .D(i_psram_sub_n_1084), .Z(i_psram_sub_n_1926
		));
	notech_mux2 i_psram_sub_i_3267(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[9]), .B(i_psram_sub_n_1705), .Z(i_psram_sub_n_3478));
	notech_reg_set i_psram_sub_axi_awaddr_reg_9(.CP(s00_axi_aclk), .D(i_psram_sub_n_3478
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[9]));
	notech_ao4 i_psram_sub_i_31067(.A(i_psram_sub_n_4017), .B(i_psram_sub_n_799775
		), .C(\i_psram_sub_nbus_63[0] ), .D(i_psram_sub_n_494), .Z(i_psram_sub_n_1931
		));
	notech_mux2 i_psram_sub_i_3259(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[8]), .B(i_psram_sub_n_1700), .Z(i_psram_sub_n_3472));
	notech_reg_set i_psram_sub_axi_awaddr_reg_8(.CP(s00_axi_aclk), .D(i_psram_sub_n_3472
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[8]));
	notech_nand2 i_psram_sub_i_1765(.A(i_psram_sub_n_1075), .B(i_psram_sub_n_508
		), .Z(i_psram_sub_n_1797));
	notech_mux2 i_psram_sub_i_3251(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[7]), .B(i_psram_sub_n_1695), .Z(i_psram_sub_n_3466));
	notech_reg_set i_psram_sub_axi_awaddr_reg_7(.CP(s00_axi_aclk), .D(i_psram_sub_n_3466
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[7]));
	notech_nand2 i_psram_sub_i_2766(.A(i_psram_sub_n_1074), .B(i_psram_sub_n_509
		), .Z(i_psram_sub_n_1802));
	notech_mux2 i_psram_sub_i_3243(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[6]), .B(i_psram_sub_n_1690), .Z(i_psram_sub_n_3460));
	notech_reg_set i_psram_sub_axi_awaddr_reg_6(.CP(s00_axi_aclk), .D(i_psram_sub_n_3460
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[6]));
	notech_nand2 i_psram_sub_i_3767(.A(i_psram_sub_n_1073), .B(i_psram_sub_n_1072
		), .Z(i_psram_sub_n_1807));
	notech_mux2 i_psram_sub_i_3235(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[5]), .B(i_psram_sub_n_1685), .Z(i_psram_sub_n_3454));
	notech_reg_set i_psram_sub_axi_awaddr_reg_5(.CP(s00_axi_aclk), .D(i_psram_sub_n_3454
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[5]));
	notech_nand2 i_psram_sub_i_4768(.A(i_psram_sub_n_1071), .B(i_psram_sub_n_1070
		), .Z(i_psram_sub_n_1812));
	notech_mux2 i_psram_sub_i_3227(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[4]), .B(i_psram_sub_n_1680), .Z(i_psram_sub_n_3448));
	notech_reg_set i_psram_sub_axi_awaddr_reg_4(.CP(s00_axi_aclk), .D(i_psram_sub_n_3448
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[4]));
	notech_nand2 i_psram_sub_i_5769(.A(i_psram_sub_n_1069), .B(i_psram_sub_n_1068
		), .Z(i_psram_sub_n_1817));
	notech_mux2 i_psram_sub_i_3219(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[3]), .B(i_psram_sub_n_1675), .Z(i_psram_sub_n_3442));
	notech_reg_set i_psram_sub_axi_awaddr_reg_3(.CP(s00_axi_aclk), .D(i_psram_sub_n_3442
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[3]));
	notech_nand2 i_psram_sub_i_6770(.A(i_psram_sub_n_1067), .B(i_psram_sub_n_1066
		), .Z(i_psram_sub_n_1822));
	notech_mux2 i_psram_sub_i_3211(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[2]), .B(i_psram_sub_n_1670), .Z(i_psram_sub_n_3436));
	notech_reg_set i_psram_sub_axi_awaddr_reg_2(.CP(s00_axi_aclk), .D(i_psram_sub_n_3436
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[2]));
	notech_nand2 i_psram_sub_i_7771(.A(i_psram_sub_n_1065), .B(i_psram_sub_n_1064
		), .Z(i_psram_sub_n_1827));
	notech_mux2 i_psram_sub_i_3203(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[1]), .B(i_psram_sub_n_1665), .Z(i_psram_sub_n_3430));
	notech_reg_set i_psram_sub_axi_awaddr_reg_1(.CP(s00_axi_aclk), .D(i_psram_sub_n_3430
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[1]));
	notech_nand2 i_psram_sub_i_8772(.A(i_psram_sub_n_1063), .B(i_psram_sub_n_1062
		), .Z(i_psram_sub_n_1832));
	notech_mux2 i_psram_sub_i_3195(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awaddr
		[0]), .B(i_psram_sub_n_1660), .Z(i_psram_sub_n_3424));
	notech_reg_set i_psram_sub_axi_awaddr_reg_0(.CP(s00_axi_aclk), .D(i_psram_sub_n_3424
		), .SD(1'b1), .Q(i_psram_sub_axi_awaddr[0]));
	notech_nand2 i_psram_sub_i_9773(.A(i_psram_sub_n_1061), .B(i_psram_sub_n_1060
		), .Z(i_psram_sub_n_1837));
	notech_mux2 i_psram_sub_i_3187(.S(\i_psram_sub_nbus_63[0] ), .A(i_psram_sub_axi_awlen
		[7]), .B(i_psram_sub_n_798774), .Z(i_psram_sub_n_3418));
	notech_reg_set i_psram_sub_axi_awlen_reg_7(.CP(s00_axi_aclk), .D(i_psram_sub_n_3418
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen[7]));
	notech_nand2 i_psram_sub_i_10774(.A(i_psram_sub_n_1059), .B(i_psram_sub_n_1058
		), .Z(i_psram_sub_n_1842));
	notech_mux2 i_psram_sub_i_3179(.S(\i_psram_sub_nbus_63[0] ), .A(i_psram_sub_axi_awlen
		[6]), .B(i_psram_sub_n_797773), .Z(i_psram_sub_n_3412));
	notech_reg_set i_psram_sub_axi_awlen_reg_6(.CP(s00_axi_aclk), .D(i_psram_sub_n_3412
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen[6]));
	notech_nand2 i_psram_sub_i_11775(.A(i_psram_sub_n_1057), .B(i_psram_sub_n_1056
		), .Z(i_psram_sub_n_1847));
	notech_mux2 i_psram_sub_i_3171(.S(\i_psram_sub_nbus_63[0] ), .A(i_psram_sub_axi_awlen
		[5]), .B(i_psram_sub_n_796772), .Z(i_psram_sub_n_3406));
	notech_reg_set i_psram_sub_axi_awlen_reg_5(.CP(s00_axi_aclk), .D(i_psram_sub_n_3406
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen[5]));
	notech_nand2 i_psram_sub_i_12776(.A(i_psram_sub_n_1055), .B(i_psram_sub_n_1054
		), .Z(i_psram_sub_n_1852));
	notech_mux2 i_psram_sub_i_3163(.S(\i_psram_sub_nbus_63[0] ), .A(i_psram_sub_axi_awlen
		[4]), .B(i_psram_sub_n_795771), .Z(i_psram_sub_n_3400));
	notech_reg_set i_psram_sub_axi_awlen_reg_4(.CP(s00_axi_aclk), .D(i_psram_sub_n_3400
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen[4]));
	notech_nand2 i_psram_sub_i_13777(.A(i_psram_sub_n_1053), .B(i_psram_sub_n_1052
		), .Z(i_psram_sub_n_1857));
	notech_mux2 i_psram_sub_i_3155(.S(\i_psram_sub_nbus_63[0] ), .A(i_psram_sub_axi_awlen
		[3]), .B(i_psram_sub_n_794770), .Z(i_psram_sub_n_3394));
	notech_reg_set i_psram_sub_axi_awlen_reg_3(.CP(s00_axi_aclk), .D(i_psram_sub_n_3394
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen[3]));
	notech_nand2 i_psram_sub_i_14778(.A(i_psram_sub_n_1051), .B(i_psram_sub_n_1050
		), .Z(i_psram_sub_n_1862));
	notech_mux2 i_psram_sub_i_3147(.S(\i_psram_sub_nbus_63[0] ), .A(i_psram_sub_axi_awlen
		[2]), .B(i_psram_sub_n_793769), .Z(i_psram_sub_n_3388));
	notech_reg_set i_psram_sub_axi_awlen_reg_2(.CP(s00_axi_aclk), .D(i_psram_sub_n_3388
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen[2]));
	notech_nand2 i_psram_sub_i_15779(.A(i_psram_sub_n_1049), .B(i_psram_sub_n_1048
		), .Z(i_psram_sub_n_1867));
	notech_mux2 i_psram_sub_i_3139(.S(\i_psram_sub_nbus_63[0] ), .A(i_psram_sub_axi_awlen
		[1]), .B(i_psram_sub_n_792768), .Z(i_psram_sub_n_3382));
	notech_reg_set i_psram_sub_axi_awlen_reg_1(.CP(s00_axi_aclk), .D(i_psram_sub_n_3382
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen[1]));
	notech_nand2 i_psram_sub_i_16780(.A(i_psram_sub_n_1047), .B(i_psram_sub_n_1046
		), .Z(i_psram_sub_n_1872));
	notech_mux2 i_psram_sub_i_3131(.S(\i_psram_sub_nbus_63[0] ), .A(i_psram_sub_axi_awlen
		[0]), .B(i_psram_sub_n_791767), .Z(i_psram_sub_n_3376));
	notech_reg_set i_psram_sub_axi_awlen_reg_0(.CP(s00_axi_aclk), .D(i_psram_sub_n_3376
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen[0]));
	notech_nand2 i_psram_sub_i_17781(.A(i_psram_sub_n_1045), .B(i_psram_sub_n_1044
		), .Z(i_psram_sub_n_1877));
	notech_mux2 i_psram_sub_i_3123(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awlen_cntr
		[7]), .B(i_psram_sub_n_804780), .Z(i_psram_sub_n_3370));
	notech_reg_set i_psram_sub_axi_awlen_cntr_reg_7(.CP(s00_axi_aclk), .D(i_psram_sub_n_3370
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen_cntr[7]));
	notech_nand2 i_psram_sub_i_18782(.A(i_psram_sub_n_1043), .B(i_psram_sub_n_1042
		), .Z(i_psram_sub_n_1882));
	notech_mux2 i_psram_sub_i_3115(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awlen_cntr
		[6]), .B(i_psram_sub_n_803779), .Z(i_psram_sub_n_3364));
	notech_reg_set i_psram_sub_axi_awlen_cntr_reg_6(.CP(s00_axi_aclk), .D(i_psram_sub_n_3364
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen_cntr[6]));
	notech_nand2 i_psram_sub_i_19783(.A(i_psram_sub_n_1041), .B(i_psram_sub_n_1040
		), .Z(i_psram_sub_n_1887));
	notech_mux2 i_psram_sub_i_3107(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awlen_cntr
		[5]), .B(i_psram_sub_n_802778), .Z(i_psram_sub_n_3358));
	notech_reg_set i_psram_sub_axi_awlen_cntr_reg_5(.CP(s00_axi_aclk), .D(i_psram_sub_n_3358
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen_cntr[5]));
	notech_nand2 i_psram_sub_i_20784(.A(i_psram_sub_n_1039), .B(i_psram_sub_n_1038
		), .Z(i_psram_sub_n_1892));
	notech_mux2 i_psram_sub_i_3099(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awlen_cntr
		[4]), .B(i_psram_sub_n_801777), .Z(i_psram_sub_n_3352));
	notech_reg_set i_psram_sub_axi_awlen_cntr_reg_4(.CP(s00_axi_aclk), .D(i_psram_sub_n_3352
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen_cntr[4]));
	notech_nand2 i_psram_sub_i_21785(.A(i_psram_sub_n_1037), .B(i_psram_sub_n_1036
		), .Z(i_psram_sub_n_1897));
	notech_mux2 i_psram_sub_i_3091(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awlen_cntr
		[3]), .B(i_psram_sub_n_800776), .Z(i_psram_sub_n_3346));
	notech_reg_set i_psram_sub_axi_awlen_cntr_reg_3(.CP(s00_axi_aclk), .D(i_psram_sub_n_3346
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen_cntr[3]));
	notech_nand2 i_psram_sub_i_22786(.A(i_psram_sub_n_1035), .B(i_psram_sub_n_1034
		), .Z(i_psram_sub_n_1902));
	notech_mux2 i_psram_sub_i_3083(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awlen_cntr
		[2]), .B(i_psram_sub_n_4016), .Z(i_psram_sub_n_3340));
	notech_reg_set i_psram_sub_axi_awlen_cntr_reg_2(.CP(s00_axi_aclk), .D(i_psram_sub_n_3340
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen_cntr[2]));
	notech_nand2 i_psram_sub_i_23787(.A(i_psram_sub_n_1033), .B(i_psram_sub_n_1032
		), .Z(i_psram_sub_n_1907));
	notech_mux2 i_psram_sub_i_3075(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awlen_cntr
		[1]), .B(i_psram_sub_n_4014), .Z(i_psram_sub_n_3334));
	notech_reg_set i_psram_sub_axi_awlen_cntr_reg_1(.CP(s00_axi_aclk), .D(i_psram_sub_n_3334
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen_cntr[1]));
	notech_nand2 i_psram_sub_i_24788(.A(i_psram_sub_n_1031), .B(i_psram_sub_n_1026
		), .Z(i_psram_sub_n_1912));
	notech_mux2 i_psram_sub_i_3067(.S(\i_psram_sub_nbus_60[0] ), .A(i_psram_sub_axi_awlen_cntr
		[0]), .B(i_psram_sub_n_4012), .Z(i_psram_sub_n_3328));
	notech_reg_set i_psram_sub_axi_awlen_cntr_reg_0(.CP(s00_axi_aclk), .D(i_psram_sub_n_3328
		), .SD(1'b1), .Q(i_psram_sub_axi_awlen_cntr[0]));
	notech_ao4 i_psram_sub_i_21050(.A(i_psram_sub_n_913), .B(i_psram_sub_n_4004
		), .C(\i_psram_sub_nbus_67[0] ), .D(i_psram_sub_n_1013), .Z(i_psram_sub_n_2067
		));
	notech_mux2 i_psram_sub_i_3059(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[23]), .B(i_psram_sub_n_1912), .Z(i_psram_sub_n_3322));
	notech_reg_set i_psram_sub_axi_araddr_reg_23(.CP(s00_axi_aclk), .D(i_psram_sub_n_3322
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[23]));
	notech_ao4 i_psram_sub_i_31051(.A(i_psram_sub_n_4006), .B(i_psram_sub_n_913
		), .C(i_psram_sub_n_535), .D(\i_psram_sub_nbus_67[0] ), .Z(i_psram_sub_n_2072
		));
	notech_mux2 i_psram_sub_i_3051(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[22]), .B(i_psram_sub_n_1907), .Z(i_psram_sub_n_3316));
	notech_reg_set i_psram_sub_axi_araddr_reg_22(.CP(s00_axi_aclk), .D(i_psram_sub_n_3316
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[22]));
	notech_nand2 i_psram_sub_i_1329(.A(i_psram_sub_n_1004), .B(i_psram_sub_n_549
		), .Z(i_psram_sub_n_1553));
	notech_mux2 i_psram_sub_i_3043(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[21]), .B(i_psram_sub_n_1902), .Z(i_psram_sub_n_3310));
	notech_reg_set i_psram_sub_axi_araddr_reg_21(.CP(s00_axi_aclk), .D(i_psram_sub_n_3310
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[21]));
	notech_nand2 i_psram_sub_i_2330(.A(i_psram_sub_n_1001), .B(i_psram_sub_n_550
		), .Z(i_psram_sub_n_1558));
	notech_mux2 i_psram_sub_i_3035(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[20]), .B(i_psram_sub_n_1897), .Z(i_psram_sub_n_3304));
	notech_reg_set i_psram_sub_axi_araddr_reg_20(.CP(s00_axi_aclk), .D(i_psram_sub_n_3304
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[20]));
	notech_nand2 i_psram_sub_i_3331(.A(i_psram_sub_n_1000), .B(i_psram_sub_n_551
		), .Z(i_psram_sub_n_1563));
	notech_mux2 i_psram_sub_i_3027(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[19]), .B(i_psram_sub_n_1892), .Z(i_psram_sub_n_3298));
	notech_reg_set i_psram_sub_axi_araddr_reg_19(.CP(s00_axi_aclk), .D(i_psram_sub_n_3298
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[19]));
	notech_nand2 i_psram_sub_i_4332(.A(i_psram_sub_n_999), .B(i_psram_sub_n_552
		), .Z(i_psram_sub_n_1568));
	notech_mux2 i_psram_sub_i_3019(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[18]), .B(i_psram_sub_n_1887), .Z(i_psram_sub_n_3292));
	notech_reg_set i_psram_sub_axi_araddr_reg_18(.CP(s00_axi_aclk), .D(i_psram_sub_n_3292
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[18]));
	notech_nand2 i_psram_sub_i_5333(.A(i_psram_sub_n_998), .B(i_psram_sub_n_553
		), .Z(i_psram_sub_n_1573));
	notech_mux2 i_psram_sub_i_3011(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[17]), .B(i_psram_sub_n_1882), .Z(i_psram_sub_n_3286));
	notech_reg_set i_psram_sub_axi_araddr_reg_17(.CP(s00_axi_aclk), .D(i_psram_sub_n_3286
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[17]));
	notech_nand2 i_psram_sub_i_6334(.A(i_psram_sub_n_997), .B(i_psram_sub_n_554
		), .Z(i_psram_sub_n_1578));
	notech_mux2 i_psram_sub_i_3003(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[16]), .B(i_psram_sub_n_1877), .Z(i_psram_sub_n_3280));
	notech_reg_set i_psram_sub_axi_araddr_reg_16(.CP(s00_axi_aclk), .D(i_psram_sub_n_3280
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[16]));
	notech_nand2 i_psram_sub_i_7335(.A(i_psram_sub_n_996), .B(i_psram_sub_n_555
		), .Z(i_psram_sub_n_1583));
	notech_mux2 i_psram_sub_i_2995(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[15]), .B(i_psram_sub_n_1872), .Z(i_psram_sub_n_3274));
	notech_reg_set i_psram_sub_axi_araddr_reg_15(.CP(s00_axi_aclk), .D(i_psram_sub_n_3274
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[15]));
	notech_nand2 i_psram_sub_i_8336(.A(i_psram_sub_n_995), .B(i_psram_sub_n_556
		), .Z(i_psram_sub_n_1588));
	notech_mux2 i_psram_sub_i_2986(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[14]), .B(i_psram_sub_n_1867), .Z(i_psram_sub_n_3268));
	notech_reg_set i_psram_sub_axi_araddr_reg_14(.CP(s00_axi_aclk), .D(i_psram_sub_n_3268
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[14]));
	notech_nand2 i_psram_sub_i_9337(.A(i_psram_sub_n_994), .B(i_psram_sub_n_557
		), .Z(i_psram_sub_n_1593));
	notech_mux2 i_psram_sub_i_2978(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[13]), .B(i_psram_sub_n_1862), .Z(i_psram_sub_n_3262));
	notech_reg_set i_psram_sub_axi_araddr_reg_13(.CP(s00_axi_aclk), .D(i_psram_sub_n_3262
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[13]));
	notech_nand2 i_psram_sub_i_10338(.A(i_psram_sub_n_993), .B(i_psram_sub_n_558
		), .Z(i_psram_sub_n_1598));
	notech_mux2 i_psram_sub_i_2970(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[12]), .B(i_psram_sub_n_1857), .Z(i_psram_sub_n_3256));
	notech_reg_set i_psram_sub_axi_araddr_reg_12(.CP(s00_axi_aclk), .D(i_psram_sub_n_3256
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[12]));
	notech_nand2 i_psram_sub_i_11339(.A(i_psram_sub_n_992), .B(i_psram_sub_n_559
		), .Z(i_psram_sub_n_1603));
	notech_mux2 i_psram_sub_i_2962(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[11]), .B(i_psram_sub_n_1852), .Z(i_psram_sub_n_3250));
	notech_reg_set i_psram_sub_axi_araddr_reg_11(.CP(s00_axi_aclk), .D(i_psram_sub_n_3250
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[11]));
	notech_nand2 i_psram_sub_i_12340(.A(i_psram_sub_n_991), .B(i_psram_sub_n_560
		), .Z(i_psram_sub_n_1608));
	notech_mux2 i_psram_sub_i_2954(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[10]), .B(i_psram_sub_n_1847), .Z(i_psram_sub_n_3244));
	notech_reg_set i_psram_sub_axi_araddr_reg_10(.CP(s00_axi_aclk), .D(i_psram_sub_n_3244
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[10]));
	notech_nand2 i_psram_sub_i_13341(.A(i_psram_sub_n_990), .B(i_psram_sub_n_561
		), .Z(i_psram_sub_n_1613));
	notech_mux2 i_psram_sub_i_2946(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[9]), .B(i_psram_sub_n_1842), .Z(i_psram_sub_n_3238));
	notech_reg_set i_psram_sub_axi_araddr_reg_9(.CP(s00_axi_aclk), .D(i_psram_sub_n_3238
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[9]));
	notech_nand2 i_psram_sub_i_14342(.A(i_psram_sub_n_989), .B(i_psram_sub_n_562
		), .Z(i_psram_sub_n_1618));
	notech_mux2 i_psram_sub_i_2938(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[8]), .B(i_psram_sub_n_1837), .Z(i_psram_sub_n_3232));
	notech_reg_set i_psram_sub_axi_araddr_reg_8(.CP(s00_axi_aclk), .D(i_psram_sub_n_3232
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[8]));
	notech_nand2 i_psram_sub_i_15343(.A(i_psram_sub_n_988), .B(i_psram_sub_n_563
		), .Z(i_psram_sub_n_1623));
	notech_mux2 i_psram_sub_i_2930(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[7]), .B(i_psram_sub_n_1832), .Z(i_psram_sub_n_3226));
	notech_reg_set i_psram_sub_axi_araddr_reg_7(.CP(s00_axi_aclk), .D(i_psram_sub_n_3226
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[7]));
	notech_nand2 i_psram_sub_i_16344(.A(i_psram_sub_n_987), .B(i_psram_sub_n_565
		), .Z(i_psram_sub_n_1628));
	notech_mux2 i_psram_sub_i_2922(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[6]), .B(i_psram_sub_n_1827), .Z(i_psram_sub_n_3220));
	notech_reg_set i_psram_sub_axi_araddr_reg_6(.CP(s00_axi_aclk), .D(i_psram_sub_n_3220
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[6]));
	notech_ao4 i_psram_sub_i_811(.A(i_psram_sub_n_451), .B(i_psram_sub_n_985
		), .C(i_psram_sub_n_961), .D(i_psram_sub_n_984), .Z(i_psram_sub_n_1639
		));
	notech_mux2 i_psram_sub_i_2914(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[5]), .B(i_psram_sub_n_1822), .Z(i_psram_sub_n_3214));
	notech_reg_set i_psram_sub_axi_araddr_reg_5(.CP(s00_axi_aclk), .D(i_psram_sub_n_3214
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[5]));
	notech_nao3 i_psram_sub_i_798(.A(s00_axi_aresetn), .B(i_psram_sub_n_1205
		), .C(i_psram_sub_n_975), .Z(i_psram_sub_n_2054));
	notech_mux2 i_psram_sub_i_2906(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[4]), .B(i_psram_sub_n_1817), .Z(i_psram_sub_n_3208));
	notech_reg_set i_psram_sub_axi_araddr_reg_4(.CP(s00_axi_aclk), .D(i_psram_sub_n_3208
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[4]));
	notech_nao3 i_psram_sub_i_3896(.A(i_psram_sub_n_570), .B(i_psram_sub_n_372
		), .C(i_psram_sub_n_571), .Z(i_psram_sub_state_5[2]));
	notech_mux2 i_psram_sub_i_2898(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[3]), .B(i_psram_sub_n_1812), .Z(i_psram_sub_n_3202));
	notech_reg_set i_psram_sub_axi_araddr_reg_3(.CP(s00_axi_aclk), .D(i_psram_sub_n_3202
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[3]));
	notech_nao3 i_psram_sub_i_2895(.A(i_psram_sub_n_1235), .B(i_psram_sub_n_574
		), .C(i_psram_sub_n_573), .Z(i_psram_sub_state_5[1]));
	notech_mux2 i_psram_sub_i_2889(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[2]), .B(i_psram_sub_n_1807), .Z(i_psram_sub_n_3196));
	notech_reg_set i_psram_sub_axi_araddr_reg_2(.CP(s00_axi_aclk), .D(i_psram_sub_n_3196
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[2]));
	notech_ao4 i_psram_sub_i_1894(.A(i_psram_sub_n_1231), .B(i_psram_sub_axi_araddr
		[1]), .C(i_psram_sub_n_377), .D(i_psram_sub_mem_idle), .Z(i_psram_sub_state_5
		[0]));
	notech_mux2 i_psram_sub_i_2881(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[1]), .B(i_psram_sub_n_1802), .Z(i_psram_sub_n_3190));
	notech_reg_set i_psram_sub_axi_araddr_reg_1(.CP(s00_axi_aclk), .D(i_psram_sub_n_3190
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[1]));
	notech_nao3 i_psram_sub_i_860(.A(i_psram_sub_n_954), .B(s00_axi_aresetn)
		, .C(i_psram_sub_n_382), .Z(\i_psram_sub_nbus_58[0] ));
	notech_mux2 i_psram_sub_i_2873(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_araddr
		[0]), .B(i_psram_sub_n_1797), .Z(i_psram_sub_n_3184));
	notech_reg_set i_psram_sub_axi_araddr_reg_0(.CP(s00_axi_aclk), .D(i_psram_sub_n_3184
		), .SD(1'b1), .Q(i_psram_sub_axi_araddr[0]));
	notech_nand3 i_psram_sub_i_862(.A(i_psram_sub_n_954), .B(s00_axi_aresetn
		), .C(i_psram_sub_n_416), .Z(\i_psram_sub_nbus_58[16] ));
	notech_mux2 i_psram_sub_i_2865(.S(\i_psram_sub_nbus_67[0] ), .A(i_psram_sub_axi_arlen
		[7]), .B(i_psram_sub_n_912), .Z(i_psram_sub_n_3178));
	notech_reg_set i_psram_sub_axi_arlen_reg_7(.CP(s00_axi_aclk), .D(i_psram_sub_n_3178
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen[7]));
	notech_nand3 i_psram_sub_i_1021(.A(s00_axi_aresetn), .B(i_psram_sub_n_569
		), .C(i_psram_sub_n_449), .Z(i_psram_sub_n_2024));
	notech_mux2 i_psram_sub_i_2857(.S(\i_psram_sub_nbus_67[0] ), .A(i_psram_sub_axi_arlen
		[6]), .B(i_psram_sub_n_911), .Z(i_psram_sub_n_3172));
	notech_reg_set i_psram_sub_axi_arlen_reg_6(.CP(s00_axi_aclk), .D(i_psram_sub_n_3172
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen[6]));
	notech_nand3 i_psram_sub_i_1113(.A(i_psram_sub_n_954), .B(i_psram_sub_n_374
		), .C(s00_axi_aresetn), .Z(i_psram_sub_n_2173));
	notech_mux2 i_psram_sub_i_2849(.S(\i_psram_sub_nbus_67[0] ), .A(i_psram_sub_axi_arlen
		[5]), .B(i_psram_sub_n_910), .Z(i_psram_sub_n_3166));
	notech_reg_set i_psram_sub_axi_arlen_reg_5(.CP(s00_axi_aclk), .D(i_psram_sub_n_3166
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen[5]));
	notech_nao3 i_psram_sub_i_1122(.A(s00_axi_aresetn), .B(i_psram_sub_n_1225
		), .C(i_psram_sub_n_982), .Z(i_psram_sub_n_2198));
	notech_mux2 i_psram_sub_i_2841(.S(\i_psram_sub_nbus_67[0] ), .A(i_psram_sub_axi_arlen
		[4]), .B(i_psram_sub_n_909), .Z(i_psram_sub_n_3160));
	notech_reg_set i_psram_sub_axi_arlen_reg_4(.CP(s00_axi_aclk), .D(i_psram_sub_n_3160
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen[4]));
	notech_nand3 i_psram_sub_i_957(.A(s00_axi_aresetn), .B(i_psram_sub_n_1225
		), .C(i_psram_sub_n_982), .Z(i_psram_sub_n_1786));
	notech_mux2 i_psram_sub_i_2832(.S(\i_psram_sub_nbus_67[0] ), .A(i_psram_sub_axi_arlen
		[3]), .B(i_psram_sub_n_908), .Z(i_psram_sub_n_3154));
	notech_reg_set i_psram_sub_axi_arlen_reg_3(.CP(s00_axi_aclk), .D(i_psram_sub_n_3154
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen[3]));
	notech_or4 i_psram_sub_i_922(.A(i_psram_sub_state[1]), .B(i_psram_sub_n_958
		), .C(i_psram_sub_mem_idle), .D(i_psram_sub_state[2]), .Z(\i_psram_sub_nbus_56[0] 
		));
	notech_mux2 i_psram_sub_i_2824(.S(\i_psram_sub_nbus_67[0] ), .A(i_psram_sub_axi_arlen
		[2]), .B(i_psram_sub_n_907), .Z(i_psram_sub_n_3148));
	notech_reg_set i_psram_sub_axi_arlen_reg_2(.CP(s00_axi_aclk), .D(i_psram_sub_n_3148
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen[2]));
	notech_nao3 i_psram_sub_i_1102(.A(s00_axi_aresetn), .B(i_psram_sub_n_1223
		), .C(i_psram_sub_n_1222), .Z(i_psram_sub_n_2159));
	notech_mux2 i_psram_sub_i_2816(.S(\i_psram_sub_nbus_67[0] ), .A(i_psram_sub_axi_arlen
		[1]), .B(i_psram_sub_n_906), .Z(i_psram_sub_n_3142));
	notech_reg_set i_psram_sub_axi_arlen_reg_1(.CP(s00_axi_aclk), .D(i_psram_sub_n_3142
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen[1]));
	notech_nand3 i_psram_sub_i_1002(.A(s00_axi_aresetn), .B(i_psram_sub_n_1222
		), .C(i_psram_sub_n_1223), .Z(i_psram_sub_n_1970));
	notech_mux2 i_psram_sub_i_2808(.S(\i_psram_sub_nbus_67[0] ), .A(i_psram_sub_axi_arlen
		[0]), .B(i_psram_sub_n_905), .Z(i_psram_sub_n_3136));
	notech_reg_set i_psram_sub_axi_arlen_reg_0(.CP(s00_axi_aclk), .D(i_psram_sub_n_3136
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen[0]));
	notech_nao3 i_psram_sub_i_1029(.A(i_psram_sub_n_985), .B(i_psram_sub_n_596
		), .C(i_psram_sub_n_958), .Z(\i_psram_sub_nbus_64[0] ));
	notech_mux2 i_psram_sub_i_2800(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_arlen_cntr
		[7]), .B(i_psram_sub_n_918), .Z(i_psram_sub_n_3130));
	notech_reg_set i_psram_sub_axi_arlen_cntr_reg_7(.CP(s00_axi_aclk), .D(i_psram_sub_n_3130
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen_cntr[7]));
	notech_nand3 i_psram_sub_i_929(.A(s00_axi_aresetn), .B(i_psram_sub_n_1077
		), .C(i_psram_sub_n_463), .Z(\i_psram_sub_nbus_60[0] ));
	notech_mux2 i_psram_sub_i_2792(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_arlen_cntr
		[6]), .B(i_psram_sub_n_917), .Z(i_psram_sub_n_3124));
	notech_reg_set i_psram_sub_axi_arlen_cntr_reg_6(.CP(s00_axi_aclk), .D(i_psram_sub_n_3124
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen_cntr[6]));
	notech_nand2 i_psram_sub_i_1007(.A(s00_axi_aresetn), .B(i_psram_sub_n_1077
		), .Z(\i_psram_sub_nbus_63[0] ));
	notech_mux2 i_psram_sub_i_2784(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_arlen_cntr
		[5]), .B(i_psram_sub_n_916), .Z(i_psram_sub_n_3118));
	notech_reg_set i_psram_sub_axi_arlen_cntr_reg_5(.CP(s00_axi_aclk), .D(i_psram_sub_n_3118
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen_cntr[5]));
	notech_nand3 i_psram_sub_i_962(.A(s00_axi_aresetn), .B(i_psram_sub_n_1006
		), .C(i_psram_sub_n_511), .Z(\i_psram_sub_nbus_61[0] ));
	notech_mux2 i_psram_sub_i_2776(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_arlen_cntr
		[4]), .B(i_psram_sub_n_915), .Z(i_psram_sub_n_3112));
	notech_reg_set i_psram_sub_axi_arlen_cntr_reg_4(.CP(s00_axi_aclk), .D(i_psram_sub_n_3112
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen_cntr[4]));
	notech_nand2 i_psram_sub_i_1085(.A(s00_axi_aresetn), .B(i_psram_sub_n_1006
		), .Z(\i_psram_sub_nbus_67[0] ));
	notech_mux2 i_psram_sub_i_2768(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_arlen_cntr
		[3]), .B(i_psram_sub_n_914), .Z(i_psram_sub_n_3106));
	notech_reg_set i_psram_sub_axi_arlen_cntr_reg_3(.CP(s00_axi_aclk), .D(i_psram_sub_n_3106
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen_cntr[3]));
	notech_mux2 i_psram_sub_i_2759(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_arlen_cntr
		[2]), .B(i_psram_sub_n_4005), .Z(i_psram_sub_n_3100));
	notech_reg_set i_psram_sub_axi_arlen_cntr_reg_2(.CP(s00_axi_aclk), .D(i_psram_sub_n_3100
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen_cntr[2]));
	notech_and2 i_psram_sub_i_1095(.A(s00_axi_aresetn), .B(i_psram_sub_n_569
		), .Z(\i_psram_sub_nbus_68[0] ));
	notech_mux2 i_psram_sub_i_2751(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_arlen_cntr
		[1]), .B(i_psram_sub_n_4003), .Z(i_psram_sub_n_3094));
	notech_reg_set i_psram_sub_axi_arlen_cntr_reg_1(.CP(s00_axi_aclk), .D(i_psram_sub_n_3094
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen_cntr[1]));
	notech_and4 i_psram_sub_i_765(.A(i_psram_sub_n_976), .B(i_psram_sub_n_972
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_952), .Z(i_psram_sub_go_7
		));
	notech_mux2 i_psram_sub_i_2743(.S(\i_psram_sub_nbus_61[0] ), .A(i_psram_sub_axi_arlen_cntr
		[0]), .B(i_psram_sub_n_4030), .Z(i_psram_sub_n_3088));
	notech_reg_set i_psram_sub_axi_arlen_cntr_reg_0(.CP(s00_axi_aclk), .D(i_psram_sub_n_3088
		), .SD(1'b1), .Q(i_psram_sub_axi_arlen_cntr[0]));
	notech_mux2 i_psram_sub_i_2735(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[15]), .B(i_psram_sub_n_1628), .Z(i_psram_sub_n_3082));
	notech_reg_set i_psram_sub_mem_data_wr_reg_15(.CP(s00_axi_aclk), .D(i_psram_sub_n_3082
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[15]));
	notech_ao4 i_psram_sub_i_651(.A(i_psram_sub_mem_idle), .B(i_psram_sub_n_970
		), .C(i_psram_sub_n_1231), .D(i_psram_sub_axi_araddr[1]), .Z(i_psram_sub_n_1235
		));
	notech_mux2 i_psram_sub_i_2727(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[14]), .B(i_psram_sub_n_1623), .Z(i_psram_sub_n_3076));
	notech_reg_set i_psram_sub_mem_data_wr_reg_14(.CP(s00_axi_aclk), .D(i_psram_sub_n_3076
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[14]));
	notech_mux2 i_psram_sub_i_2719(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[13]), .B(i_psram_sub_n_1618), .Z(i_psram_sub_n_3070));
	notech_reg_set i_psram_sub_mem_data_wr_reg_13(.CP(s00_axi_aclk), .D(i_psram_sub_n_3070
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[13]));
	notech_mux2 i_psram_sub_i_2711(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[12]), .B(i_psram_sub_n_1613), .Z(i_psram_sub_n_3064));
	notech_reg_set i_psram_sub_mem_data_wr_reg_12(.CP(s00_axi_aclk), .D(i_psram_sub_n_3064
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[12]));
	notech_mux2 i_psram_sub_i_2703(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[11]), .B(i_psram_sub_n_1608), .Z(i_psram_sub_n_3058));
	notech_reg_set i_psram_sub_mem_data_wr_reg_11(.CP(s00_axi_aclk), .D(i_psram_sub_n_3058
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[11]));
	notech_or4 i_psram_sub_i_86(.A(i_psram_sub_n_954), .B(i_psram_sub_n_4319
		), .C(i_psram_sub_n_4024), .D(i_psram_sub_mem_idle), .Z(i_psram_sub_n_1231
		));
	notech_mux2 i_psram_sub_i_2694(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[10]), .B(i_psram_sub_n_1603), .Z(i_psram_sub_n_3052));
	notech_reg_set i_psram_sub_mem_data_wr_reg_10(.CP(s00_axi_aclk), .D(i_psram_sub_n_3052
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[10]));
	notech_mux2 i_psram_sub_i_2686(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[9]), .B(i_psram_sub_n_1598), .Z(i_psram_sub_n_3046));
	notech_reg_set i_psram_sub_mem_data_wr_reg_9(.CP(s00_axi_aclk), .D(i_psram_sub_n_3046
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[9]));
	notech_mux2 i_psram_sub_i_2678(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[8]), .B(i_psram_sub_n_1593), .Z(i_psram_sub_n_3040));
	notech_reg_set i_psram_sub_mem_data_wr_reg_8(.CP(s00_axi_aclk), .D(i_psram_sub_n_3040
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[8]));
	notech_ao4 i_psram_sub_i_658(.A(i_psram_sub_n_974), .B(i_psram_sub_n_4319
		), .C(i_psram_sub_n_979), .D(i_psram_sub_n_1227), .Z(i_psram_sub_n_1228
		));
	notech_mux2 i_psram_sub_i_2670(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[7]), .B(i_psram_sub_n_1588), .Z(i_psram_sub_n_3034));
	notech_reg_set i_psram_sub_mem_data_wr_reg_7(.CP(s00_axi_aclk), .D(i_psram_sub_n_3034
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[7]));
	notech_or4 i_psram_sub_i_85(.A(i_psram_sub_state[1]), .B(i_psram_sub_state
		[0]), .C(i_psram_sub_n_4027), .D(i_psram_sub_n_4319), .Z(i_psram_sub_n_1227
		));
	notech_mux2 i_psram_sub_i_2662(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[6]), .B(i_psram_sub_n_1583), .Z(i_psram_sub_n_3028));
	notech_reg_set i_psram_sub_mem_data_wr_reg_6(.CP(s00_axi_aclk), .D(i_psram_sub_n_3028
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[6]));
	notech_mux2 i_psram_sub_i_2654(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[5]), .B(i_psram_sub_n_1578), .Z(i_psram_sub_n_3022));
	notech_reg_set i_psram_sub_mem_data_wr_reg_5(.CP(s00_axi_aclk), .D(i_psram_sub_n_3022
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[5]));
	notech_nand2 i_psram_sub_i_47(.A(i_psram_sub_n_4024), .B(i_psram_sub_n_3991
		), .Z(i_psram_sub_n_1225));
	notech_mux2 i_psram_sub_i_2646(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[4]), .B(i_psram_sub_n_1573), .Z(i_psram_sub_n_3016));
	notech_reg_set i_psram_sub_mem_data_wr_reg_4(.CP(s00_axi_aclk), .D(i_psram_sub_n_3016
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[4]));
	notech_mux2 i_psram_sub_i_2638(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[3]), .B(i_psram_sub_n_1568), .Z(i_psram_sub_n_3010));
	notech_reg_set i_psram_sub_mem_data_wr_reg_3(.CP(s00_axi_aclk), .D(i_psram_sub_n_3010
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[3]));
	notech_or2 i_psram_sub_i_44(.A(i_psram_sub_n_1006), .B(i_psram_sub_axi_awv_awr_flag
		), .Z(i_psram_sub_n_1223));
	notech_mux2 i_psram_sub_i_2630(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[2]), .B(i_psram_sub_n_1563), .Z(i_psram_sub_n_3004));
	notech_reg_set i_psram_sub_mem_data_wr_reg_2(.CP(s00_axi_aclk), .D(i_psram_sub_n_3004
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[2]));
	notech_and4 i_psram_sub_i_77(.A(i_psram_sub_n_1213), .B(s00_axi_rvalid),
		 .C(s00_axi_rready), .D(i_psram_sub_n_3992), .Z(i_psram_sub_n_1222
		));
	notech_mux2 i_psram_sub_i_2622(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[1]), .B(i_psram_sub_n_1558), .Z(i_psram_sub_n_2998));
	notech_reg_set i_psram_sub_mem_data_wr_reg_1(.CP(s00_axi_aclk), .D(i_psram_sub_n_2998
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[1]));
	notech_mux2 i_psram_sub_i_2614(.S(\i_psram_sub_nbus_56[0] ), .A(i_psram_sub_mem_data_wr
		[0]), .B(i_psram_sub_n_1553), .Z(i_psram_sub_n_2992));
	notech_reg_set i_psram_sub_mem_data_wr_reg_0(.CP(s00_axi_aclk), .D(i_psram_sub_n_2992
		), .SD(1'b1), .Q(i_psram_sub_mem_data_wr[0]));
	notech_reg_set i_psram_sub_go_reg(.CP(s00_axi_aclk), .D(i_psram_sub_n_4002
		), .SD(1'b1), .Q(i_psram_sub_go));
	notech_or4 i_psram_sub_i_673(.A(i_psram_sub_n_587), .B(i_psram_sub_n_586
		), .C(i_psram_sub_n_1219), .D(i_psram_sub_n_1214), .Z(i_psram_sub_n_1220
		));
	notech_or4 i_psram_sub_i_669(.A(i_psram_sub_n_583), .B(i_psram_sub_n_582
		), .C(i_psram_sub_n_585), .D(i_psram_sub_n_584), .Z(i_psram_sub_n_1219
		));
	notech_nand2 i_psram_sub_i_671(.A(i_psram_sub_n_589), .B(i_psram_sub_n_588
		), .Z(i_psram_sub_n_1214));
	notech_and4 i_psram_sub_i_680(.A(i_psram_sub_n_1211), .B(i_psram_sub_n_1210
		), .C(i_psram_sub_n_1208), .D(i_psram_sub_n_1207), .Z(i_psram_sub_n_1213
		));
	notech_ao4 i_psram_sub_i_674(.A(i_psram_sub_axi_arlen_cntr[0]), .B(i_psram_sub_n_4008
		), .C(i_psram_sub_axi_arlen[1]), .D(i_psram_sub_n_4004), .Z(i_psram_sub_n_1211
		));
	notech_ao4 i_psram_sub_i_675(.A(i_psram_sub_axi_arlen[2]), .B(i_psram_sub_n_4006
		), .C(i_psram_sub_axi_arlen[3]), .D(i_psram_sub_n_4007), .Z(i_psram_sub_n_1210
		));
	notech_ao4 i_psram_sub_i_677(.A(i_psram_sub_axi_arlen_cntr[4]), .B(i_psram_sub_n_4009
		), .C(i_psram_sub_axi_arlen_cntr[5]), .D(i_psram_sub_n_4010), .Z
		(i_psram_sub_n_1208));
	notech_ao4 i_psram_sub_i_678(.A(i_psram_sub_axi_arlen_cntr[6]), .B(i_psram_sub_n_4011
		), .C(i_psram_sub_axi_arlen_cntr[7]), .D(i_psram_sub_n_4013), .Z
		(i_psram_sub_n_1207));
	notech_ao4 i_psram_sub_i_682(.A(i_psram_sub_n_3995), .B(i_psram_sub_n_954
		), .C(i_psram_sub_n_962), .D(i_psram_sub_n_1204), .Z(i_psram_sub_n_1205
		));
	notech_nand2 i_psram_sub_i_683(.A(i_psram_sub_command), .B(i_psram_sub_n_954
		), .Z(i_psram_sub_n_1204));
	notech_ao4 i_psram_sub_i_685(.A(s00_axi_wstrb[0]), .B(i_psram_sub_n_971)
		, .C(i_psram_sub_n_962), .D(i_psram_sub_n_1201), .Z(i_psram_sub_n_1202
		));
	notech_nand3 i_psram_sub_i_686(.A(s00_axi_aresetn), .B(i_psram_sub_n_954
		), .C(i_psram_sub_mem_byte_en[0]), .Z(i_psram_sub_n_1201));
	notech_ao4 i_psram_sub_i_57(.A(i_psram_sub_n_3994), .B(i_psram_sub_n_980
		), .C(i_psram_sub_n_3995), .D(i_psram_sub_n_1197), .Z(i_psram_sub_n_1198
		));
	notech_nao3 i_psram_sub_i_690(.A(i_psram_sub_n_568), .B(s00_axi_aresetn)
		, .C(i_psram_sub_n_954), .Z(i_psram_sub_n_1197));
	notech_ao4 i_psram_sub_i_689(.A(s00_axi_wstrb[1]), .B(i_psram_sub_n_971)
		, .C(i_psram_sub_n_962), .D(i_psram_sub_n_1195), .Z(i_psram_sub_n_1196
		));
	notech_nand3 i_psram_sub_i_691(.A(s00_axi_aresetn), .B(i_psram_sub_n_954
		), .C(i_psram_sub_mem_byte_en[1]), .Z(i_psram_sub_n_1195));
	notech_ao4 i_psram_sub_i_692(.A(i_psram_sub_n_969), .B(i_psram_sub_n_965
		), .C(i_psram_sub_n_456), .D(i_psram_sub_n_4199), .Z(i_psram_sub_n_1194
		));
	notech_ao4 i_psram_sub_i_693(.A(i_psram_sub_n_455), .B(i_psram_sub_n_4176
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4105), .Z(i_psram_sub_n_1193
		));
	notech_ao4 i_psram_sub_i_694(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4200
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4177), .Z(i_psram_sub_n_1192
		));
	notech_ao4 i_psram_sub_i_695(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4154
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4106), .Z(i_psram_sub_n_1191
		));
	notech_ao4 i_psram_sub_i_696(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4201
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4178), .Z(i_psram_sub_n_1190
		));
	notech_ao4 i_psram_sub_i_697(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4155
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4107), .Z(i_psram_sub_n_1189
		));
	notech_ao4 i_psram_sub_i_698(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4202
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4179), .Z(i_psram_sub_n_1188
		));
	notech_ao4 i_psram_sub_i_699(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4156
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4108), .Z(i_psram_sub_n_1187
		));
	notech_ao4 i_psram_sub_i_700(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4203
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4180), .Z(i_psram_sub_n_1186
		));
	notech_ao4 i_psram_sub_i_701(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4157
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4109), .Z(i_psram_sub_n_1185
		));
	notech_ao4 i_psram_sub_i_702(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4204
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4181), .Z(i_psram_sub_n_1184
		));
	notech_ao4 i_psram_sub_i_703(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4158
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4110), .Z(i_psram_sub_n_1183
		));
	notech_ao4 i_psram_sub_i_704(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4205
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4182), .Z(i_psram_sub_n_1182
		));
	notech_ao4 i_psram_sub_i_705(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4159
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4111), .Z(i_psram_sub_n_1181
		));
	notech_ao4 i_psram_sub_i_706(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4206
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4183), .Z(i_psram_sub_n_1180
		));
	notech_ao4 i_psram_sub_i_707(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4160
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4112), .Z(i_psram_sub_n_1179
		));
	notech_ao4 i_psram_sub_i_708(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4207
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4184), .Z(i_psram_sub_n_1178
		));
	notech_ao4 i_psram_sub_i_709(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4161
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4113), .Z(i_psram_sub_n_1177
		));
	notech_ao4 i_psram_sub_i_710(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4208
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4185), .Z(i_psram_sub_n_1176
		));
	notech_ao4 i_psram_sub_i_711(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4162
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4114), .Z(i_psram_sub_n_1175
		));
	notech_ao4 i_psram_sub_i_712(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4209
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4186), .Z(i_psram_sub_n_1174
		));
	notech_ao4 i_psram_sub_i_713(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4163
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4115), .Z(i_psram_sub_n_1173
		));
	notech_ao4 i_psram_sub_i_714(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4210
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4187), .Z(i_psram_sub_n_1172
		));
	notech_ao4 i_psram_sub_i_715(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4164
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4116), .Z(i_psram_sub_n_1171
		));
	notech_ao4 i_psram_sub_i_716(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4211
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4188), .Z(i_psram_sub_n_1170
		));
	notech_ao4 i_psram_sub_i_717(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4165
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4117), .Z(i_psram_sub_n_1169
		));
	notech_ao4 i_psram_sub_i_718(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4212
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4189), .Z(i_psram_sub_n_1168
		));
	notech_ao4 i_psram_sub_i_719(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4166
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4118), .Z(i_psram_sub_n_1167
		));
	notech_ao4 i_psram_sub_i_720(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4213
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4190), .Z(i_psram_sub_n_1166
		));
	notech_ao4 i_psram_sub_i_721(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4167
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4119), .Z(i_psram_sub_n_1165
		));
	notech_ao4 i_psram_sub_i_722(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4214
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4191), .Z(i_psram_sub_n_1164
		));
	notech_ao4 i_psram_sub_i_723(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4168
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4120), .Z(i_psram_sub_n_1163
		));
	notech_ao4 i_psram_sub_i_724(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4215
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4192), .Z(i_psram_sub_n_1162
		));
	notech_ao4 i_psram_sub_i_725(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4169
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4121), .Z(i_psram_sub_n_1161
		));
	notech_ao4 i_psram_sub_i_726(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4216
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4193), .Z(i_psram_sub_n_1160
		));
	notech_ao4 i_psram_sub_i_727(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4170
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4122), .Z(i_psram_sub_n_1159
		));
	notech_ao4 i_psram_sub_i_728(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4217
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4194), .Z(i_psram_sub_n_1158
		));
	notech_ao4 i_psram_sub_i_729(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4171
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4123), .Z(i_psram_sub_n_1157
		));
	notech_ao4 i_psram_sub_i_730(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4218
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4195), .Z(i_psram_sub_n_1156
		));
	notech_ao4 i_psram_sub_i_731(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4172
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4124), .Z(i_psram_sub_n_1155
		));
	notech_ao4 i_psram_sub_i_732(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4219
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4196), .Z(i_psram_sub_n_1154
		));
	notech_ao4 i_psram_sub_i_733(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4173
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4125), .Z(i_psram_sub_n_1153
		));
	notech_ao4 i_psram_sub_i_734(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4220
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4197), .Z(i_psram_sub_n_1152
		));
	notech_ao4 i_psram_sub_i_735(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4174
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4126), .Z(i_psram_sub_n_1151
		));
	notech_ao4 i_psram_sub_i_736(.A(i_psram_sub_n_456), .B(i_psram_sub_n_4221
		), .C(i_psram_sub_n_455), .D(i_psram_sub_n_4198), .Z(i_psram_sub_n_1150
		));
	notech_and2 i_psram_sub_i_48(.A(i_psram_sub_n_974), .B(i_psram_sub_n_960
		), .Z(i_psram_sub_n_1149));
	notech_ao4 i_psram_sub_i_737(.A(i_psram_sub_n_972), .B(i_psram_sub_n_4175
		), .C(i_psram_sub_n_957), .D(i_psram_sub_n_4127), .Z(i_psram_sub_n_1148
		));
	notech_ao4 i_psram_sub_i_738(.A(i_psram_sub_n_1101), .B(i_psram_sub_n_4128
		), .C(i_psram_sub_n_1097), .D(i_psram_sub_n_4152), .Z(i_psram_sub_n_1147
		));
	notech_ao4 i_psram_sub_i_739(.A(i_psram_sub_n_4129), .B(i_psram_sub_n_1101
		), .C(i_psram_sub_n_1097), .D(i_psram_sub_n_4153), .Z(i_psram_sub_n_1146
		));
	notech_ao4 i_psram_sub_i_740(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4260
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4130), .Z(i_psram_sub_n_1145
		));
	notech_ao4 i_psram_sub_i_741(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4154
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4381), .Z(i_psram_sub_n_1144
		));
	notech_ao4 i_psram_sub_i_742(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4261
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4131), .Z(i_psram_sub_n_1143
		));
	notech_ao4 i_psram_sub_i_743(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4155
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4380), .Z(i_psram_sub_n_1142
		));
	notech_ao4 i_psram_sub_i_744(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4262
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4132), .Z(i_psram_sub_n_1141
		));
	notech_ao4 i_psram_sub_i_745(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4156
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4379), .Z(i_psram_sub_n_1140
		));
	notech_ao4 i_psram_sub_i_746(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4263
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4133), .Z(i_psram_sub_n_1139
		));
	notech_ao4 i_psram_sub_i_747(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4157
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4378), .Z(i_psram_sub_n_1138
		));
	notech_ao4 i_psram_sub_i_749(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4264
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4134), .Z(i_psram_sub_n_1137
		));
	notech_ao4 i_psram_sub_i_750(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4158
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4377), .Z(i_psram_sub_n_1136
		));
	notech_ao4 i_psram_sub_i_751(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4265
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4135), .Z(i_psram_sub_n_1135
		));
	notech_ao4 i_psram_sub_i_752(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4159
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4376), .Z(i_psram_sub_n_1134
		));
	notech_ao4 i_psram_sub_i_753(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4266
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4136), .Z(i_psram_sub_n_1133
		));
	notech_ao4 i_psram_sub_i_754(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4160
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4375), .Z(i_psram_sub_n_1132
		));
	notech_ao4 i_psram_sub_i_755(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4267
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4137), .Z(i_psram_sub_n_1131
		));
	notech_ao4 i_psram_sub_i_756(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4161
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4374), .Z(i_psram_sub_n_1130
		));
	notech_ao4 i_psram_sub_i_757(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4268
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4138), .Z(i_psram_sub_n_1129
		));
	notech_ao4 i_psram_sub_i_758(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4162
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4373), .Z(i_psram_sub_n_1128
		));
	notech_ao4 i_psram_sub_i_759(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4269
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4139), .Z(i_psram_sub_n_1127
		));
	notech_ao4 i_psram_sub_i_760(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4163
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4372), .Z(i_psram_sub_n_1126
		));
	notech_ao4 i_psram_sub_i_761(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4270
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4140), .Z(i_psram_sub_n_1125
		));
	notech_ao4 i_psram_sub_i_762(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4164
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4371), .Z(i_psram_sub_n_1124
		));
	notech_ao4 i_psram_sub_i_763(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4271
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4141), .Z(i_psram_sub_n_1123
		));
	notech_ao4 i_psram_sub_i_764(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4165
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4370), .Z(i_psram_sub_n_1122
		));
	notech_ao4 i_psram_sub_i_766(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4272
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4142), .Z(i_psram_sub_n_1121
		));
	notech_ao4 i_psram_sub_i_767(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4166
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4369), .Z(i_psram_sub_n_1120
		));
	notech_ao4 i_psram_sub_i_768(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4273
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4143), .Z(i_psram_sub_n_1119
		));
	notech_ao4 i_psram_sub_i_769(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4167
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4368), .Z(i_psram_sub_n_1118
		));
	notech_ao4 i_psram_sub_i_770(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4274
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4144), .Z(i_psram_sub_n_1117
		));
	notech_ao4 i_psram_sub_i_771(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4168
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4367), .Z(i_psram_sub_n_1116
		));
	notech_ao4 i_psram_sub_i_772(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4275
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4145), .Z(i_psram_sub_n_1115
		));
	notech_ao4 i_psram_sub_i_773(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4169
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4366), .Z(i_psram_sub_n_1114
		));
	notech_ao4 i_psram_sub_i_774(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4276
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4146), .Z(i_psram_sub_n_1113
		));
	notech_ao4 i_psram_sub_i_775(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4170
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4365), .Z(i_psram_sub_n_1112
		));
	notech_ao4 i_psram_sub_i_776(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4277
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4147), .Z(i_psram_sub_n_1111
		));
	notech_ao4 i_psram_sub_i_777(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4171
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4364), .Z(i_psram_sub_n_1110
		));
	notech_ao4 i_psram_sub_i_778(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4278
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4148), .Z(i_psram_sub_n_1109
		));
	notech_ao4 i_psram_sub_i_779(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4172
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4363), .Z(i_psram_sub_n_1108
		));
	notech_ao4 i_psram_sub_i_780(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4279
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4149), .Z(i_psram_sub_n_1107
		));
	notech_ao4 i_psram_sub_i_781(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4173
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4362), .Z(i_psram_sub_n_1106
		));
	notech_ao4 i_psram_sub_i_782(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4280
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4150), .Z(i_psram_sub_n_1105
		));
	notech_ao4 i_psram_sub_i_783(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4174
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4361), .Z(i_psram_sub_n_1104
		));
	notech_ao4 i_psram_sub_i_784(.A(i_psram_sub_n_1102), .B(i_psram_sub_n_4281
		), .C(i_psram_sub_n_1101), .D(i_psram_sub_n_4151), .Z(i_psram_sub_n_1103
		));
	notech_nand2 i_psram_sub_i_5(.A(s00_axi_aresetn), .B(i_psram_sub_n_3991)
		, .Z(i_psram_sub_n_1102));
	notech_or4 i_psram_sub_i_8(.A(\i_psram_sub_nbus_63[0] ), .B(s00_axi_awburst
		[0]), .C(i_psram_sub_n_3998), .D(i_psram_sub_n_4317), .Z(i_psram_sub_n_1101
		));
	notech_ao4 i_psram_sub_i_785(.A(i_psram_sub_n_1097), .B(i_psram_sub_n_4175
		), .C(i_psram_sub_n_1095), .D(i_psram_sub_n_4360), .Z(i_psram_sub_n_1098
		));
	notech_nao3 i_psram_sub_i_9(.A(i_psram_sub_n_4317), .B(i_psram_sub_n_4316
		), .C(\i_psram_sub_nbus_63[0] ), .Z(i_psram_sub_n_1097));
	notech_nand3 i_psram_sub_i_13(.A(s00_axi_aresetn), .B(i_psram_sub_n_1077
		), .C(i_psram_sub_n_370), .Z(i_psram_sub_n_1095));
	notech_and4 i_psram_sub_i_491563(.A(i_psram_sub_n_1092), .B(i_psram_sub_n_1091
		), .C(i_psram_sub_n_1089), .D(i_psram_sub_n_1088), .Z(i_psram_sub_n_1094
		));
	notech_ao4 i_psram_sub_i_789(.A(i_psram_sub_axi_awaddr[2]), .B(i_psram_sub_n_4359
		), .C(i_psram_sub_axi_awaddr[3]), .D(i_psram_sub_n_4358), .Z(i_psram_sub_n_1092
		));
	notech_ao4 i_psram_sub_i_790(.A(i_psram_sub_axi_awaddr[4]), .B(i_psram_sub_n_4357
		), .C(i_psram_sub_axi_awaddr[5]), .D(i_psram_sub_n_4356), .Z(i_psram_sub_n_1091
		));
	notech_ao4 i_psram_sub_i_792(.A(i_psram_sub_axi_awaddr[6]), .B(i_psram_sub_n_4355
		), .C(i_psram_sub_axi_awaddr[7]), .D(i_psram_sub_n_4354), .Z(i_psram_sub_n_1089
		));
	notech_ao4 i_psram_sub_i_793(.A(i_psram_sub_axi_awaddr[8]), .B(i_psram_sub_n_4353
		), .C(i_psram_sub_axi_awaddr[9]), .D(i_psram_sub_n_4352), .Z(i_psram_sub_n_1088
		));
	notech_ao4 i_psram_sub_i_22(.A(i_psram_sub_axi_awlen[3]), .B(i_psram_sub_n_4018
		), .C(i_psram_sub_n_482), .D(i_psram_sub_n_481), .Z(i_psram_sub_n_1086
		));
	notech_nand2 i_psram_sub_i_806(.A(i_psram_sub_axi_awlen_cntr[0]), .B(i_psram_sub_n_4019
		), .Z(i_psram_sub_n_1085));
	notech_nand2 i_psram_sub_i_807(.A(i_psram_sub_axi_awlen_cntr[0]), .B(i_psram_sub_n_4015
		), .Z(i_psram_sub_n_1084));
	notech_and3 i_psram_sub_i_70(.A(i_psram_sub_axi_awlen_cntr[5]), .B(i_psram_sub_n_1081
		), .C(i_psram_sub_axi_awlen_cntr[6]), .Z(i_psram_sub_n_1083));
	notech_and3 i_psram_sub_i_53(.A(i_psram_sub_axi_awlen_cntr[4]), .B(i_psram_sub_n_1080
		), .C(i_psram_sub_axi_awlen_cntr[5]), .Z(i_psram_sub_n_1082));
	notech_ao3 i_psram_sub_i_46(.A(i_psram_sub_axi_awlen_cntr[4]), .B(i_psram_sub_axi_awlen_cntr
		[3]), .C(i_psram_sub_n_1079), .Z(i_psram_sub_n_1081));
	notech_and4 i_psram_sub_i_40(.A(i_psram_sub_axi_awlen_cntr[0]), .B(i_psram_sub_axi_awlen_cntr
		[1]), .C(i_psram_sub_axi_awlen_cntr[2]), .D(i_psram_sub_axi_awlen_cntr
		[3]), .Z(i_psram_sub_n_1080));
	notech_nand3 i_psram_sub_i_101507(.A(i_psram_sub_axi_awlen_cntr[0]), .B(i_psram_sub_axi_awlen_cntr
		[1]), .C(i_psram_sub_axi_awlen_cntr[2]), .Z(i_psram_sub_n_1079)
		);
	notech_nand2 i_psram_sub_i_818(.A(i_psram_sub_axi_awlen_cntr[0]), .B(i_psram_sub_axi_awlen_cntr
		[1]), .Z(i_psram_sub_n_1078));
	notech_nao3 i_psram_sub_i_472(.A(s00_axi_awvalid), .B(i_psram_sub_n_4399
		), .C(i_psram_sub_axi_awv_awr_flag), .Z(i_psram_sub_n_1077));
	notech_ao4 i_psram_sub_i_826(.A(i_psram_sub_n_4080), .B(i_psram_sub_n_1029
		), .C(i_psram_sub_n_1025), .D(i_psram_sub_n_4104), .Z(i_psram_sub_n_1075
		));
	notech_ao4 i_psram_sub_i_827(.A(i_psram_sub_n_1029), .B(i_psram_sub_n_4081
		), .C(i_psram_sub_n_1025), .D(i_psram_sub_n_4105), .Z(i_psram_sub_n_1074
		));
	notech_ao4 i_psram_sub_i_828(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4238
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4082), .Z(i_psram_sub_n_1073
		));
	notech_ao4 i_psram_sub_i_829(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4106
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4351), .Z(i_psram_sub_n_1072
		));
	notech_ao4 i_psram_sub_i_830(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4239
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4083), .Z(i_psram_sub_n_1071
		));
	notech_ao4 i_psram_sub_i_831(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4107
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4350), .Z(i_psram_sub_n_1070
		));
	notech_ao4 i_psram_sub_i_832(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4240
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4084), .Z(i_psram_sub_n_1069
		));
	notech_ao4 i_psram_sub_i_833(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4108
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4349), .Z(i_psram_sub_n_1068
		));
	notech_ao4 i_psram_sub_i_834(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4241
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4085), .Z(i_psram_sub_n_1067
		));
	notech_ao4 i_psram_sub_i_835(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4109
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4348), .Z(i_psram_sub_n_1066
		));
	notech_ao4 i_psram_sub_i_836(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4242
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4086), .Z(i_psram_sub_n_1065
		));
	notech_ao4 i_psram_sub_i_837(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4110
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4347), .Z(i_psram_sub_n_1064
		));
	notech_ao4 i_psram_sub_i_838(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4243
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4087), .Z(i_psram_sub_n_1063
		));
	notech_ao4 i_psram_sub_i_839(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4111
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4346), .Z(i_psram_sub_n_1062
		));
	notech_ao4 i_psram_sub_i_840(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4244
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4088), .Z(i_psram_sub_n_1061
		));
	notech_ao4 i_psram_sub_i_841(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4112
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4345), .Z(i_psram_sub_n_1060
		));
	notech_ao4 i_psram_sub_i_842(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4245
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4089), .Z(i_psram_sub_n_1059
		));
	notech_ao4 i_psram_sub_i_843(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4113
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4344), .Z(i_psram_sub_n_1058
		));
	notech_ao4 i_psram_sub_i_844(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4246
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4090), .Z(i_psram_sub_n_1057
		));
	notech_ao4 i_psram_sub_i_845(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4114
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4343), .Z(i_psram_sub_n_1056
		));
	notech_ao4 i_psram_sub_i_846(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4247
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4091), .Z(i_psram_sub_n_1055
		));
	notech_ao4 i_psram_sub_i_847(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4115
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4342), .Z(i_psram_sub_n_1054
		));
	notech_ao4 i_psram_sub_i_848(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4248
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4092), .Z(i_psram_sub_n_1053
		));
	notech_ao4 i_psram_sub_i_849(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4116
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4341), .Z(i_psram_sub_n_1052
		));
	notech_ao4 i_psram_sub_i_863(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4249
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4093), .Z(i_psram_sub_n_1051
		));
	notech_ao4 i_psram_sub_i_864(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4117
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4340), .Z(i_psram_sub_n_1050
		));
	notech_ao4 i_psram_sub_i_865(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4250
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4094), .Z(i_psram_sub_n_1049
		));
	notech_ao4 i_psram_sub_i_866(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4118
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4339), .Z(i_psram_sub_n_1048
		));
	notech_ao4 i_psram_sub_i_867(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4251
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4095), .Z(i_psram_sub_n_1047
		));
	notech_ao4 i_psram_sub_i_868(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4119
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4338), .Z(i_psram_sub_n_1046
		));
	notech_ao4 i_psram_sub_i_869(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4252
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4096), .Z(i_psram_sub_n_1045
		));
	notech_ao4 i_psram_sub_i_870(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4120
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4337), .Z(i_psram_sub_n_1044
		));
	notech_ao4 i_psram_sub_i_871(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4253
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4097), .Z(i_psram_sub_n_1043
		));
	notech_ao4 i_psram_sub_i_872(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4121
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4336), .Z(i_psram_sub_n_1042
		));
	notech_ao4 i_psram_sub_i_873(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4254
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4098), .Z(i_psram_sub_n_1041
		));
	notech_ao4 i_psram_sub_i_874(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4122
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4335), .Z(i_psram_sub_n_1040
		));
	notech_ao4 i_psram_sub_i_875(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4255
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4099), .Z(i_psram_sub_n_1039
		));
	notech_ao4 i_psram_sub_i_876(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4123
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4334), .Z(i_psram_sub_n_1038
		));
	notech_ao4 i_psram_sub_i_877(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4256
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4100), .Z(i_psram_sub_n_1037
		));
	notech_ao4 i_psram_sub_i_878(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4124
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4333), .Z(i_psram_sub_n_1036
		));
	notech_ao4 i_psram_sub_i_879(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4257
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4101), .Z(i_psram_sub_n_1035
		));
	notech_ao4 i_psram_sub_i_880(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4125
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4332), .Z(i_psram_sub_n_1034
		));
	notech_ao4 i_psram_sub_i_881(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4258
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4102), .Z(i_psram_sub_n_1033
		));
	notech_ao4 i_psram_sub_i_882(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4126
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4331), .Z(i_psram_sub_n_1032
		));
	notech_ao4 i_psram_sub_i_883(.A(i_psram_sub_n_1030), .B(i_psram_sub_n_4259
		), .C(i_psram_sub_n_1029), .D(i_psram_sub_n_4103), .Z(i_psram_sub_n_1031
		));
	notech_nand2 i_psram_sub_i_6(.A(s00_axi_aresetn), .B(i_psram_sub_n_3990)
		, .Z(i_psram_sub_n_1030));
	notech_or4 i_psram_sub_i_7(.A(\i_psram_sub_nbus_67[0] ), .B(s00_axi_arburst
		[0]), .C(i_psram_sub_n_3999), .D(i_psram_sub_n_4318), .Z(i_psram_sub_n_1029
		));
	notech_ao4 i_psram_sub_i_884(.A(i_psram_sub_n_1025), .B(i_psram_sub_n_4127
		), .C(i_psram_sub_n_1023), .D(i_psram_sub_n_4330), .Z(i_psram_sub_n_1026
		));
	notech_or4 i_psram_sub_i_10(.A(s00_axi_arburst[0]), .B(i_psram_sub_n_4319
		), .C(s00_axi_arburst[1]), .D(i_psram_sub_n_3990), .Z(i_psram_sub_n_1025
		));
	notech_nand3 i_psram_sub_i_15(.A(i_psram_sub_n_1006), .B(s00_axi_aresetn
		), .C(i_psram_sub_n_371), .Z(i_psram_sub_n_1023));
	notech_and4 i_psram_sub_i_49(.A(i_psram_sub_n_1020), .B(i_psram_sub_n_1019
		), .C(i_psram_sub_n_1017), .D(i_psram_sub_n_1016), .Z(i_psram_sub_n_1022
		));
	notech_ao4 i_psram_sub_i_888(.A(i_psram_sub_axi_araddr[2]), .B(i_psram_sub_n_4329
		), .C(i_psram_sub_axi_araddr[3]), .D(i_psram_sub_n_4328), .Z(i_psram_sub_n_1020
		));
	notech_ao4 i_psram_sub_i_889(.A(i_psram_sub_axi_araddr[4]), .B(i_psram_sub_n_4327
		), .C(i_psram_sub_axi_araddr[5]), .D(i_psram_sub_n_4326), .Z(i_psram_sub_n_1019
		));
	notech_ao4 i_psram_sub_i_891(.A(i_psram_sub_axi_araddr[6]), .B(i_psram_sub_n_4325
		), .C(i_psram_sub_axi_araddr[7]), .D(i_psram_sub_n_4324), .Z(i_psram_sub_n_1017
		));
	notech_ao4 i_psram_sub_i_892(.A(i_psram_sub_axi_araddr[8]), .B(i_psram_sub_n_4323
		), .C(i_psram_sub_axi_araddr[9]), .D(i_psram_sub_n_4322), .Z(i_psram_sub_n_1016
		));
	notech_ao4 i_psram_sub_i_21(.A(i_psram_sub_axi_arlen[3]), .B(i_psram_sub_n_4007
		), .C(i_psram_sub_n_525), .D(i_psram_sub_n_584), .Z(i_psram_sub_n_1015
		));
	notech_nand2 i_psram_sub_i_909(.A(i_psram_sub_axi_arlen_cntr[0]), .B(i_psram_sub_n_4004
		), .Z(i_psram_sub_n_1013));
	notech_and3 i_psram_sub_i_69(.A(i_psram_sub_axi_arlen_cntr[5]), .B(i_psram_sub_n_1010
		), .C(i_psram_sub_axi_arlen_cntr[6]), .Z(i_psram_sub_n_1012));
	notech_and3 i_psram_sub_i_52(.A(i_psram_sub_axi_arlen_cntr[4]), .B(i_psram_sub_n_1009
		), .C(i_psram_sub_axi_arlen_cntr[5]), .Z(i_psram_sub_n_1011));
	notech_ao3 i_psram_sub_i_45(.A(i_psram_sub_axi_arlen_cntr[4]), .B(i_psram_sub_axi_arlen_cntr
		[3]), .C(i_psram_sub_n_1008), .Z(i_psram_sub_n_1010));
	notech_and4 i_psram_sub_i_36(.A(i_psram_sub_axi_arlen_cntr[0]), .B(i_psram_sub_axi_arlen_cntr
		[1]), .C(i_psram_sub_axi_arlen_cntr[2]), .D(i_psram_sub_axi_arlen_cntr
		[3]), .Z(i_psram_sub_n_1009));
	notech_nand3 i_psram_sub_i_101456(.A(i_psram_sub_axi_arlen_cntr[0]), .B(i_psram_sub_axi_arlen_cntr
		[1]), .C(i_psram_sub_axi_arlen_cntr[2]), .Z(i_psram_sub_n_1008)
		);
	notech_nand2 i_psram_sub_i_923(.A(i_psram_sub_axi_arlen_cntr[0]), .B(i_psram_sub_axi_arlen_cntr
		[1]), .Z(i_psram_sub_n_1007));
	notech_nao3 i_psram_sub_i_490(.A(s00_axi_arvalid), .B(i_psram_sub_n_4024
		), .C(s00_axi_arready), .Z(i_psram_sub_n_1006));
	notech_ao4 i_psram_sub_i_925(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4064
		), .C(i_psram_sub_n_971), .D(i_psram_sub_n_4222), .Z(i_psram_sub_n_1004
		));
	notech_ao4 i_psram_sub_i_932(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4065
		), .C(i_psram_sub_n_971), .D(i_psram_sub_n_4223), .Z(i_psram_sub_n_1001
		));
	notech_ao4 i_psram_sub_i_933(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4066
		), .C(i_psram_sub_n_971), .D(i_psram_sub_n_4224), .Z(i_psram_sub_n_1000
		));
	notech_ao4 i_psram_sub_i_934(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4067
		), .C(i_psram_sub_n_971), .D(i_psram_sub_n_4225), .Z(i_psram_sub_n_999
		));
	notech_ao4 i_psram_sub_i_935(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4068
		), .C(i_psram_sub_n_971), .D(i_psram_sub_n_4226), .Z(i_psram_sub_n_998
		));
	notech_ao4 i_psram_sub_i_936(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4069
		), .C(i_psram_sub_n_971), .D(i_psram_sub_n_4227), .Z(i_psram_sub_n_997
		));
	notech_ao4 i_psram_sub_i_937(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4070
		), .C(i_psram_sub_n_971), .D(i_psram_sub_n_4228), .Z(i_psram_sub_n_996
		));
	notech_ao4 i_psram_sub_i_938(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4071
		), .C(i_psram_sub_n_971), .D(i_psram_sub_n_4229), .Z(i_psram_sub_n_995
		));
	notech_ao4 i_psram_sub_i_939(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4072
		), .C(i_psram_sub_n_971), .D(i_psram_sub_n_4230), .Z(i_psram_sub_n_994
		));
	notech_ao4 i_psram_sub_i_940(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4073
		), .C(i_psram_sub_n_971), .D(i_psram_sub_n_4231), .Z(i_psram_sub_n_993
		));
	notech_ao4 i_psram_sub_i_941(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4074
		), .C(i_psram_sub_n_971), .D(i_psram_sub_n_4232), .Z(i_psram_sub_n_992
		));
	notech_ao4 i_psram_sub_i_942(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4075
		), .C(i_psram_sub_n_971), .D(i_psram_sub_n_4233), .Z(i_psram_sub_n_991
		));
	notech_ao4 i_psram_sub_i_943(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4076
		), .C(i_psram_sub_n_971), .D(i_psram_sub_n_4234), .Z(i_psram_sub_n_990
		));
	notech_ao4 i_psram_sub_i_944(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4077
		), .C(i_psram_sub_n_971), .D(i_psram_sub_n_4235), .Z(i_psram_sub_n_989
		));
	notech_ao4 i_psram_sub_i_945(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4078
		), .C(i_psram_sub_n_971), .D(i_psram_sub_n_4236), .Z(i_psram_sub_n_988
		));
	notech_ao4 i_psram_sub_i_946(.A(i_psram_sub_n_564), .B(i_psram_sub_n_4079
		), .C(i_psram_sub_n_4237), .D(i_psram_sub_n_971), .Z(i_psram_sub_n_987
		));
	notech_nao3 i_psram_sub_i_947(.A(i_psram_sub_n_954), .B(s00_axi_aresetn)
		, .C(i_psram_sub_n_985), .Z(i_psram_sub_n_986));
	notech_nand2 i_psram_sub_i_61438(.A(i_psram_sub_n_4027), .B(i_psram_sub_n_4025
		), .Z(i_psram_sub_n_985));
	notech_nand3 i_psram_sub_i_83(.A(i_psram_sub_n_954), .B(s00_axi_aresetn)
		, .C(i_psram_sub_n_3994), .Z(i_psram_sub_n_984));
	notech_nand2 i_psram_sub_i_68(.A(s00_axi_wready), .B(s00_axi_wlast), .Z(i_psram_sub_n_982
		));
	notech_nand3 i_psram_sub_i_73(.A(i_psram_sub_n_954), .B(i_psram_sub_n_979
		), .C(s00_axi_aresetn), .Z(i_psram_sub_n_980));
	notech_and2 i_psram_sub_i_35(.A(i_psram_sub_mem_idle), .B(i_psram_sub_n_4398
		), .Z(i_psram_sub_n_979));
	notech_nand3 i_psram_sub_i_87(.A(i_psram_sub_n_954), .B(i_psram_sub_n_975
		), .C(s00_axi_aresetn), .Z(i_psram_sub_n_976));
	notech_and4 i_psram_sub_i_67(.A(i_psram_sub_state[1]), .B(i_psram_sub_n_4027
		), .C(i_psram_sub_state[0]), .D(i_psram_sub_mem_idle), .Z(i_psram_sub_n_975
		));
	notech_nand3 i_psram_sub_i_61441(.A(i_psram_sub_state[1]), .B(i_psram_sub_n_4027
		), .C(i_psram_sub_state[0]), .Z(i_psram_sub_n_974));
	notech_and2 i_psram_sub_i_14(.A(i_psram_sub_n_971), .B(i_psram_sub_n_970
		), .Z(i_psram_sub_n_972));
	notech_or4 i_psram_sub_i_75(.A(i_psram_sub_n_954), .B(i_psram_sub_n_4319
		), .C(i_psram_sub_n_968), .D(i_psram_sub_n_3996), .Z(i_psram_sub_n_971
		));
	notech_or4 i_psram_sub_i_65(.A(i_psram_sub_n_954), .B(i_psram_sub_n_4319
		), .C(i_psram_sub_n_968), .D(i_psram_sub_n_965), .Z(i_psram_sub_n_970
		));
	notech_nao3 i_psram_sub_i_51(.A(s00_axi_aresetn), .B(i_psram_sub_n_3995)
		, .C(i_psram_sub_n_954), .Z(i_psram_sub_n_969));
	notech_or4 i_psram_sub_i_25(.A(s00_axi_wready), .B(i_psram_sub_n_4029), 
		.C(i_psram_sub_axi_arv_arr_flag), .D(i_psram_sub_n_4321), .Z(i_psram_sub_n_968
		));
	notech_or2 i_psram_sub_i_71446(.A(s00_axi_wstrb[0]), .B(s00_axi_wstrb[1]
		), .Z(i_psram_sub_n_965));
	notech_nand3 i_psram_sub_i_88(.A(i_psram_sub_n_954), .B(i_psram_sub_n_962
		), .C(s00_axi_aresetn), .Z(i_psram_sub_n_963));
	notech_ao3 i_psram_sub_i_20(.A(i_psram_sub_n_961), .B(i_psram_sub_state[
		0]), .C(i_psram_sub_n_959), .Z(i_psram_sub_n_962));
	notech_nand2 i_psram_sub_i_74(.A(i_psram_sub_n_4314), .B(i_psram_sub_n_4315
		), .Z(i_psram_sub_n_961));
	notech_nao3 i_psram_sub_i_61435(.A(i_psram_sub_n_4027), .B(i_psram_sub_state
		[0]), .C(i_psram_sub_state[1]), .Z(i_psram_sub_n_960));
	notech_or2 i_psram_sub_i_965(.A(i_psram_sub_state[1]), .B(i_psram_sub_state
		[2]), .Z(i_psram_sub_n_959));
	notech_nand2 i_psram_sub_i_0(.A(i_psram_sub_n_954), .B(s00_axi_aresetn),
		 .Z(i_psram_sub_n_958));
	notech_or4 i_psram_sub_i_89(.A(i_psram_sub_n_954), .B(s00_axi_rvalid), .C
		(i_psram_sub_n_4319), .D(i_psram_sub_n_4024), .Z(i_psram_sub_n_957
		));
	notech_or4 i_psram_sub_i_1(.A(i_psram_sub_state[1]), .B(i_psram_sub_state
		[0]), .C(i_psram_sub_state[2]), .D(i_psram_sub_n_4319), .Z(i_psram_sub_n_955
		));
	notech_nao3 i_psram_sub_i_61588(.A(i_psram_sub_n_4025), .B(i_psram_sub_n_4027
		), .C(i_psram_sub_state[1]), .Z(i_psram_sub_n_954));
	notech_nao3 i_psram_sub_i_649(.A(i_psram_sub_n_962), .B(i_psram_sub_mem_idle
		), .C(i_psram_sub_n_958), .Z(i_psram_sub_n_952));
	notech_or4 i_psram_sub_i_161596(.A(i_psram_sub_state[1]), .B(i_psram_sub_state
		[0]), .C(i_psram_sub_n_980), .D(i_psram_sub_n_4027), .Z(i_psram_sub_n_951
		));
	notech_and3 i_psram_sub_i_81056(.A(s00_axi_aresetn), .B(i_psram_sub_n_1006
		), .C(i_psram_sub_n_360), .Z(i_psram_sub_n_918));
	notech_and3 i_psram_sub_i_71055(.A(s00_axi_aresetn), .B(i_psram_sub_n_1006
		), .C(i_psram_sub_n_361), .Z(i_psram_sub_n_917));
	notech_and3 i_psram_sub_i_61054(.A(s00_axi_aresetn), .B(i_psram_sub_n_1006
		), .C(i_psram_sub_n_362), .Z(i_psram_sub_n_916));
	notech_and3 i_psram_sub_i_51053(.A(s00_axi_aresetn), .B(i_psram_sub_n_1006
		), .C(i_psram_sub_n_363), .Z(i_psram_sub_n_915));
	notech_and3 i_psram_sub_i_41052(.A(s00_axi_aresetn), .B(i_psram_sub_n_1006
		), .C(i_psram_sub_n_364), .Z(i_psram_sub_n_914));
	notech_nao3 i_psram_sub_i_11049(.A(s00_axi_aresetn), .B(i_psram_sub_n_1006
		), .C(i_psram_sub_axi_arlen_cntr[0]), .Z(i_psram_sub_n_913));
	notech_and2 i_psram_sub_i_81032(.A(s00_axi_arlen[7]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_912));
	notech_and2 i_psram_sub_i_71031(.A(s00_axi_arlen[6]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_911));
	notech_and2 i_psram_sub_i_61030(.A(s00_axi_arlen[5]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_910));
	notech_and2 i_psram_sub_i_51029(.A(s00_axi_arlen[4]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_909));
	notech_and2 i_psram_sub_i_41028(.A(s00_axi_arlen[3]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_908));
	notech_and2 i_psram_sub_i_31027(.A(s00_axi_arlen[2]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_907));
	notech_and2 i_psram_sub_i_21026(.A(s00_axi_arlen[1]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_906));
	notech_and2 i_psram_sub_i_11025(.A(s00_axi_arlen[0]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_905));
	notech_xor2 i_psram_sub_i_93(.A(i_psram_sub_axi_arlen_cntr[7]), .B(i_psram_sub_n_1012
		), .Z(i_psram_sub_n_360));
	notech_xor2 i_psram_sub_i_94(.A(i_psram_sub_axi_arlen_cntr[6]), .B(i_psram_sub_n_1011
		), .Z(i_psram_sub_n_361));
	notech_xor2 i_psram_sub_i_95(.A(i_psram_sub_axi_arlen_cntr[5]), .B(i_psram_sub_n_1010
		), .Z(i_psram_sub_n_362));
	notech_xor2 i_psram_sub_i_96(.A(i_psram_sub_axi_arlen_cntr[4]), .B(i_psram_sub_n_1009
		), .Z(i_psram_sub_n_363));
	notech_xor2 i_psram_sub_i_97(.A(i_psram_sub_n_4007), .B(i_psram_sub_n_1008
		), .Z(i_psram_sub_n_364));
	notech_xor2 i_psram_sub_i_99(.A(i_psram_sub_axi_awlen_cntr[7]), .B(i_psram_sub_n_1083
		), .Z(i_psram_sub_n_365));
	notech_xor2 i_psram_sub_i_100(.A(i_psram_sub_axi_awlen_cntr[6]), .B(i_psram_sub_n_1082
		), .Z(i_psram_sub_n_366));
	notech_xor2 i_psram_sub_i_101(.A(i_psram_sub_axi_awlen_cntr[5]), .B(i_psram_sub_n_1081
		), .Z(i_psram_sub_n_367));
	notech_xor2 i_psram_sub_i_102(.A(i_psram_sub_axi_awlen_cntr[4]), .B(i_psram_sub_n_1080
		), .Z(i_psram_sub_n_368));
	notech_xor2 i_psram_sub_i_103(.A(i_psram_sub_n_4018), .B(i_psram_sub_n_1079
		), .Z(i_psram_sub_n_369));
	notech_or2 i_psram_sub_i_106(.A(s00_axi_awburst[0]), .B(i_psram_sub_n_462
		), .Z(i_psram_sub_n_370));
	notech_or2 i_psram_sub_i_107(.A(s00_axi_arburst[0]), .B(i_psram_sub_n_510
		), .Z(i_psram_sub_n_371));
	notech_nao3 i_psram_sub_i_112(.A(i_psram_sub_mem_idle), .B(s00_axi_aresetn
		), .C(i_psram_sub_n_974), .Z(i_psram_sub_n_372));
	notech_nao3 i_psram_sub_i_62(.A(i_psram_sub_n_974), .B(i_psram_sub_n_985
		), .C(i_psram_sub_n_3994), .Z(i_psram_sub_n_374));
	notech_or2 i_psram_sub_i_118(.A(i_psram_sub_state[0]), .B(i_psram_sub_n_4398
		), .Z(i_psram_sub_n_375));
	notech_ao4 i_psram_sub_i_91(.A(i_psram_sub_n_969), .B(i_psram_sub_n_3996
		), .C(i_psram_sub_n_4319), .D(i_psram_sub_n_1149), .Z(i_psram_sub_n_377
		));
	notech_mux2 i_psram_sub_i_124(.S(i_psram_sub_state[0]), .A(i_psram_sub_state
		[2]), .B(i_psram_sub_n_959), .Z(i_psram_sub_n_382));
	notech_and3 i_psram_sub_i_3(.A(i_psram_sub_n_1227), .B(i_psram_sub_n_955
		), .C(i_psram_sub_n_576), .Z(i_psram_sub_n_413));
	notech_nao3 i_psram_sub_i_159(.A(i_psram_sub_n_985), .B(i_psram_sub_n_417
		), .C(i_psram_sub_n_3994), .Z(i_psram_sub_n_416));
	notech_nand2 i_psram_sub_i_76(.A(i_psram_sub_mem_idle), .B(i_psram_sub_n_4027
		), .Z(i_psram_sub_n_417));
	notech_and2 i_psram_sub_i_4(.A(i_psram_sub_n_1228), .B(i_psram_sub_n_955
		), .Z(i_psram_sub_n_448));
	notech_nand2 i_psram_sub_i_192(.A(s00_axi_bvalid), .B(s00_axi_bready), .Z
		(i_psram_sub_n_449));
	notech_and2 i_psram_sub_i_92(.A(i_psram_sub_n_980), .B(i_psram_sub_n_452
		), .Z(i_psram_sub_n_451));
	notech_nand3 i_psram_sub_i_194(.A(i_psram_sub_n_954), .B(s00_axi_wready)
		, .C(s00_axi_aresetn), .Z(i_psram_sub_n_452));
	notech_and2 i_psram_sub_i_12(.A(i_psram_sub_n_976), .B(i_psram_sub_n_963
		), .Z(i_psram_sub_n_455));
	notech_ao4 i_psram_sub_i_11(.A(i_psram_sub_n_958), .B(i_psram_sub_n_3993
		), .C(i_psram_sub_n_961), .D(i_psram_sub_n_984), .Z(i_psram_sub_n_456
		));
	notech_ao4 i_psram_sub_i_105(.A(i_psram_sub_n_959), .B(i_psram_sub_n_4025
		), .C(i_psram_sub_n_974), .D(i_psram_sub_n_4320), .Z(i_psram_sub_n_458
		));
	notech_nao3 i_psram_sub_i_310(.A(s00_axi_aresetn), .B(s00_axi_awaddr[0])
		, .C(i_psram_sub_n_1077), .Z(i_psram_sub_n_460));
	notech_nao3 i_psram_sub_i_313(.A(s00_axi_aresetn), .B(s00_axi_awaddr[1])
		, .C(i_psram_sub_n_1077), .Z(i_psram_sub_n_461));
	notech_and2 i_psram_sub_i_402(.A(s00_axi_awburst[1]), .B(i_psram_sub_n_3998
		), .Z(i_psram_sub_n_462));
	notech_nao3 i_psram_sub_i_416(.A(s00_axi_wvalid), .B(s00_axi_wready), .C
		(i_psram_sub_n_464), .Z(i_psram_sub_n_463));
	notech_ao4 i_psram_sub_i_82(.A(i_psram_sub_axi_awlen_cntr[7]), .B(i_psram_sub_n_4023
		), .C(i_psram_sub_n_467), .D(i_psram_sub_n_466), .Z(i_psram_sub_n_464
		));
	notech_and2 i_psram_sub_i_27(.A(i_psram_sub_axi_awlen_cntr[7]), .B(i_psram_sub_n_4023
		), .Z(i_psram_sub_n_466));
	notech_ao4 i_psram_sub_i_72(.A(i_psram_sub_axi_awlen_cntr[6]), .B(i_psram_sub_n_4022
		), .C(i_psram_sub_n_471), .D(i_psram_sub_n_470), .Z(i_psram_sub_n_467
		));
	notech_and2 i_psram_sub_i_29(.A(i_psram_sub_axi_awlen_cntr[6]), .B(i_psram_sub_n_4022
		), .Z(i_psram_sub_n_470));
	notech_ao4 i_psram_sub_i_64(.A(i_psram_sub_axi_awlen_cntr[5]), .B(i_psram_sub_n_4021
		), .C(i_psram_sub_n_475), .D(i_psram_sub_n_474), .Z(i_psram_sub_n_471
		));
	notech_and2 i_psram_sub_i_33(.A(i_psram_sub_axi_awlen_cntr[5]), .B(i_psram_sub_n_4021
		), .Z(i_psram_sub_n_474));
	notech_ao4 i_psram_sub_i_59(.A(i_psram_sub_axi_awlen_cntr[4]), .B(i_psram_sub_n_4000
		), .C(i_psram_sub_n_478), .D(i_psram_sub_n_4020), .Z(i_psram_sub_n_475
		));
	notech_and2 i_psram_sub_i_55(.A(i_psram_sub_axi_awlen_cntr[4]), .B(i_psram_sub_n_4000
		), .Z(i_psram_sub_n_478));
	notech_and2 i_psram_sub_i_31(.A(i_psram_sub_axi_awlen[3]), .B(i_psram_sub_n_4018
		), .Z(i_psram_sub_n_481));
	notech_ao4 i_psram_sub_i_109(.A(i_psram_sub_axi_awlen[2]), .B(i_psram_sub_n_4017
		), .C(i_psram_sub_n_486), .D(i_psram_sub_n_485), .Z(i_psram_sub_n_482
		));
	notech_and2 i_psram_sub_i_42(.A(i_psram_sub_axi_awlen[2]), .B(i_psram_sub_n_4017
		), .Z(i_psram_sub_n_485));
	notech_ao4 i_psram_sub_i_79(.A(i_psram_sub_axi_awlen[1]), .B(i_psram_sub_n_4015
		), .C(i_psram_sub_n_489), .D(i_psram_sub_n_1085), .Z(i_psram_sub_n_486
		));
	notech_and2 i_psram_sub_i_61(.A(i_psram_sub_axi_awlen[1]), .B(i_psram_sub_n_4015
		), .Z(i_psram_sub_n_489));
	notech_mux2 i_psram_sub_i_104(.S(i_psram_sub_axi_awlen_cntr[2]), .A(i_psram_sub_n_1078
		), .B(i_psram_sub_axi_awlen_cntr[1]), .Z(i_psram_sub_n_494));
	notech_nao3 i_psram_sub_i_457(.A(s00_axi_araddr[0]), .B(s00_axi_aresetn)
		, .C(i_psram_sub_n_1006), .Z(i_psram_sub_n_508));
	notech_nao3 i_psram_sub_i_460(.A(s00_axi_araddr[1]), .B(s00_axi_aresetn)
		, .C(i_psram_sub_n_1006), .Z(i_psram_sub_n_509));
	notech_and2 i_psram_sub_i_558(.A(s00_axi_arburst[1]), .B(i_psram_sub_n_3999
		), .Z(i_psram_sub_n_510));
	notech_nao3 i_psram_sub_i_567(.A(s00_axi_rvalid), .B(s00_axi_rready), .C
		(i_psram_sub_n_512), .Z(i_psram_sub_n_511));
	notech_ao4 i_psram_sub_i_90(.A(i_psram_sub_axi_arlen_cntr[7]), .B(i_psram_sub_n_4013
		), .C(i_psram_sub_n_514), .D(i_psram_sub_n_582), .Z(i_psram_sub_n_512
		));
	notech_ao4 i_psram_sub_i_81(.A(i_psram_sub_axi_arlen_cntr[6]), .B(i_psram_sub_n_4011
		), .C(i_psram_sub_n_517), .D(i_psram_sub_n_583), .Z(i_psram_sub_n_514
		));
	notech_ao4 i_psram_sub_i_71(.A(i_psram_sub_axi_arlen_cntr[5]), .B(i_psram_sub_n_4010
		), .C(i_psram_sub_n_520), .D(i_psram_sub_n_585), .Z(i_psram_sub_n_517
		));
	notech_ao4 i_psram_sub_i_63(.A(i_psram_sub_axi_arlen_cntr[4]), .B(i_psram_sub_n_4009
		), .C(i_psram_sub_n_587), .D(i_psram_sub_n_4001), .Z(i_psram_sub_n_520
		));
	notech_ao4 i_psram_sub_i_108(.A(i_psram_sub_axi_arlen[2]), .B(i_psram_sub_n_4006
		), .C(i_psram_sub_n_528), .D(i_psram_sub_n_586), .Z(i_psram_sub_n_525
		));
	notech_ao4 i_psram_sub_i_78(.A(i_psram_sub_axi_arlen[1]), .B(i_psram_sub_n_4004
		), .C(i_psram_sub_n_3997), .D(i_psram_sub_n_589), .Z(i_psram_sub_n_528
		));
	notech_mux2 i_psram_sub_i_98(.S(i_psram_sub_axi_arlen_cntr[2]), .A(i_psram_sub_n_1007
		), .B(i_psram_sub_axi_arlen_cntr[1]), .Z(i_psram_sub_n_535));
	notech_nand2 i_psram_sub_i_600(.A(s00_axi_wdata[16]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_549));
	notech_nand2 i_psram_sub_i_603(.A(s00_axi_wdata[17]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_550));
	notech_nand2 i_psram_sub_i_606(.A(s00_axi_wdata[18]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_551));
	notech_nand2 i_psram_sub_i_609(.A(s00_axi_wdata[19]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_552));
	notech_nand2 i_psram_sub_i_612(.A(s00_axi_wdata[20]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_553));
	notech_nand2 i_psram_sub_i_615(.A(s00_axi_wdata[21]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_554));
	notech_nand2 i_psram_sub_i_618(.A(s00_axi_wdata[22]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_555));
	notech_nand2 i_psram_sub_i_621(.A(s00_axi_wdata[23]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_556));
	notech_nand2 i_psram_sub_i_624(.A(s00_axi_wdata[24]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_557));
	notech_nand2 i_psram_sub_i_627(.A(s00_axi_wdata[25]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_558));
	notech_nand2 i_psram_sub_i_630(.A(s00_axi_wdata[26]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_559));
	notech_nand2 i_psram_sub_i_633(.A(s00_axi_wdata[27]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_560));
	notech_nand2 i_psram_sub_i_636(.A(s00_axi_wdata[28]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_561));
	notech_nand2 i_psram_sub_i_639(.A(s00_axi_wdata[29]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_562));
	notech_nand2 i_psram_sub_i_642(.A(s00_axi_wdata[30]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_563));
	notech_ao4 i_psram_sub_i_18(.A(i_psram_sub_n_979), .B(i_psram_sub_n_986)
		, .C(i_psram_sub_n_961), .D(i_psram_sub_n_984), .Z(i_psram_sub_n_564
		));
	notech_nand2 i_psram_sub_i_645(.A(s00_axi_wdata[31]), .B(i_psram_sub_n_566
		), .Z(i_psram_sub_n_565));
	notech_nand2 i_psram_sub_i_2(.A(i_psram_sub_n_970), .B(i_psram_sub_n_963
		), .Z(i_psram_sub_n_566));
	notech_or2 i_psram_sub_i_647(.A(s00_axi_rvalid), .B(i_psram_sub_n_4024),
		 .Z(i_psram_sub_n_568));
	notech_or4 i_psram_sub_i_648(.A(s00_axi_bvalid), .B(i_psram_sub_n_982), 
		.C(i_psram_sub_n_4029), .D(i_psram_sub_n_4321), .Z(i_psram_sub_n_569
		));
	notech_or4 i_psram_sub_i_110(.A(i_psram_sub_n_955), .B(i_psram_sub_mem_idle
		), .C(i_psram_sub_n_4024), .D(i_psram_sub_n_4105), .Z(i_psram_sub_n_570
		));
	notech_nor2 i_psram_sub_i_111(.A(i_psram_sub_n_979), .B(i_psram_sub_n_1227
		), .Z(i_psram_sub_n_571));
	notech_and4 i_psram_sub_i_113(.A(i_psram_sub_state[1]), .B(s00_axi_aresetn
		), .C(i_psram_sub_n_575), .D(i_psram_sub_n_374), .Z(i_psram_sub_n_573
		));
	notech_nand3 i_psram_sub_i_114(.A(i_psram_sub_n_962), .B(i_psram_sub_mem_idle
		), .C(s00_axi_aresetn), .Z(i_psram_sub_n_574));
	notech_nand2 i_psram_sub_i_34(.A(i_psram_sub_mem_idle), .B(i_psram_sub_n_375
		), .Z(i_psram_sub_n_575));
	notech_nao3 i_psram_sub_i_155(.A(s00_axi_aresetn), .B(i_psram_sub_n_4320
		), .C(i_psram_sub_n_974), .Z(i_psram_sub_n_576));
	notech_ao3 i_psram_sub_i_748(.A(i_psram_sub_n_1213), .B(i_psram_sub_n_4061
		), .C(i_psram_sub_n_1220), .Z(i_psram_sub_n_579));
	notech_ao3 i_psram_sub_i_813(.A(s00_axi_aresetn), .B(i_psram_sub_n_4024)
		, .C(i_psram_sub_n_1077), .Z(i_psram_sub_n_580));
	notech_ao3 i_psram_sub_i_802(.A(i_psram_sub_n_4029), .B(s00_axi_aresetn)
		, .C(i_psram_sub_n_1006), .Z(i_psram_sub_n_581));
	notech_and2 i_psram_sub_i_26(.A(i_psram_sub_axi_arlen_cntr[7]), .B(i_psram_sub_n_4013
		), .Z(i_psram_sub_n_582));
	notech_and2 i_psram_sub_i_28(.A(i_psram_sub_axi_arlen_cntr[6]), .B(i_psram_sub_n_4011
		), .Z(i_psram_sub_n_583));
	notech_and2 i_psram_sub_i_30(.A(i_psram_sub_axi_arlen[3]), .B(i_psram_sub_n_4007
		), .Z(i_psram_sub_n_584));
	notech_and2 i_psram_sub_i_32(.A(i_psram_sub_axi_arlen_cntr[5]), .B(i_psram_sub_n_4010
		), .Z(i_psram_sub_n_585));
	notech_and2 i_psram_sub_i_41(.A(i_psram_sub_axi_arlen[2]), .B(i_psram_sub_n_4006
		), .Z(i_psram_sub_n_586));
	notech_and2 i_psram_sub_i_54(.A(i_psram_sub_axi_arlen_cntr[4]), .B(i_psram_sub_n_4009
		), .Z(i_psram_sub_n_587));
	notech_nand2 i_psram_sub_i_58(.A(i_psram_sub_axi_arlen[1]), .B(i_psram_sub_n_4004
		), .Z(i_psram_sub_n_588));
	notech_nand2 i_psram_sub_i_203(.A(i_psram_sub_axi_arlen_cntr[0]), .B(i_psram_sub_n_4008
		), .Z(i_psram_sub_n_589));
	notech_nand2 i_psram_sub_i_208(.A(i_psram_sub_n_566), .B(i_psram_sub_n_4314
		), .Z(i_psram_sub_n_593));
	notech_or4 i_psram_sub_i_209(.A(i_psram_sub_state[1]), .B(i_psram_sub_state
		[2]), .C(i_psram_sub_n_4025), .D(i_psram_sub_n_4320), .Z(i_psram_sub_n_596
		));
	notech_nand2 i_psram_sub_i_212(.A(i_psram_sub_n_566), .B(i_psram_sub_n_4315
		), .Z(i_psram_sub_n_597));
	notech_and2 i_psram_sub_i_11033(.A(s00_axi_awlen[0]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_791767));
	notech_and2 i_psram_sub_i_21034(.A(s00_axi_awlen[1]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_792768));
	notech_and2 i_psram_sub_i_31035(.A(s00_axi_awlen[2]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_793769));
	notech_and2 i_psram_sub_i_41036(.A(s00_axi_awlen[3]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_794770));
	notech_and2 i_psram_sub_i_51037(.A(s00_axi_awlen[4]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_795771));
	notech_and2 i_psram_sub_i_61038(.A(s00_axi_awlen[5]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_796772));
	notech_and2 i_psram_sub_i_71039(.A(s00_axi_awlen[6]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_797773));
	notech_and2 i_psram_sub_i_81040(.A(s00_axi_awlen[7]), .B(s00_axi_aresetn
		), .Z(i_psram_sub_n_798774));
	notech_nao3 i_psram_sub_i_11065(.A(s00_axi_aresetn), .B(i_psram_sub_n_1077
		), .C(i_psram_sub_axi_awlen_cntr[0]), .Z(i_psram_sub_n_799775)
		);
	notech_and3 i_psram_sub_i_41068(.A(s00_axi_aresetn), .B(i_psram_sub_n_1077
		), .C(i_psram_sub_n_369), .Z(i_psram_sub_n_800776));
	notech_and3 i_psram_sub_i_51069(.A(s00_axi_aresetn), .B(i_psram_sub_n_1077
		), .C(i_psram_sub_n_368), .Z(i_psram_sub_n_801777));
	notech_and3 i_psram_sub_i_61070(.A(s00_axi_aresetn), .B(i_psram_sub_n_1077
		), .C(i_psram_sub_n_367), .Z(i_psram_sub_n_802778));
	notech_and3 i_psram_sub_i_71071(.A(s00_axi_aresetn), .B(i_psram_sub_n_1077
		), .C(i_psram_sub_n_366), .Z(i_psram_sub_n_803779));
	notech_and3 i_psram_sub_i_81072(.A(s00_axi_aresetn), .B(i_psram_sub_n_1077
		), .C(i_psram_sub_n_365), .Z(i_psram_sub_n_804780));
endmodule
