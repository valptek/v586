
module biu32_axi(rstn, clk, write_req, write_ack, write_data, write_sz, write_msk
		, read_req, read_ack, read_data, read_sz, Daddr, code_req, code_ack
		, code_data, code_addr, code_wreq, code_wack, code_wdata, readio_req
		, writeio_req, readio_ack, writeio_ack, writeio_data, readio_data
		, io_add, axi_AW, axi_AWVALID, axi_AWREADY, axi_AWBURST, axi_AWLEN
		, axi_AWSIZE, axi_W, axi_WVALID, axi_WREADY, axi_WSTRB, axi_WLAST
		, axi_AR, axi_ARVALID, axi_ARREADY, axi_ARBURST, axi_ARLEN, axi_ARSIZE
		, axi_R, axi_RVALID, axi_RREADY, axi_RLAST, axi_io_AW, axi_io_AWVALID
		, axi_io_AWREADY, axi_io_AWBURST, axi_io_AWLEN, axi_io_AWSIZE, axi_io_W
		, axi_io_WVALID, axi_io_WREADY, axi_io_WSTRB, axi_io_WLAST, axi_io_AR
		, axi_io_ARVALID, axi_io_ARREADY, axi_io_ARBURST, axi_io_ARLEN, axi_io_ARSIZE
		, axi_io_R, axi_io_RVALID, axi_io_RREADY, axi_io_RLAST, busy, outstanding
		);

	input rstn;
	input clk;
	input write_req;
	output write_ack;
	input [31:0] write_data;
	input [1:0] write_sz;
	input [3:0] write_msk;
	input read_req;
	output read_ack;
	output [31:0] read_data;
	input [1:0] read_sz;
	input [31:0] Daddr;
	input code_req;
	output code_ack;
	output [127:0] code_data;
	input [31:0] code_addr;
	input code_wreq;
	output code_wack;
	input [31:0] code_wdata;
	input readio_req;
	input writeio_req;
	output readio_ack;
	output writeio_ack;
	input [31:0] writeio_data;
	output [31:0] readio_data;
	input [31:0] io_add;
	output [31:0] axi_AW;
	output axi_AWVALID;
	input axi_AWREADY;
	output [1:0] axi_AWBURST;
	output [7:0] axi_AWLEN;
	output [2:0] axi_AWSIZE;
	output [31:0] axi_W;
	output axi_WVALID;
	input axi_WREADY;
	output [3:0] axi_WSTRB;
	output axi_WLAST;
	output [31:0] axi_AR;
	output axi_ARVALID;
	input axi_ARREADY;
	output [1:0] axi_ARBURST;
	output [7:0] axi_ARLEN;
	output [2:0] axi_ARSIZE;
	input [31:0] axi_R;
	input axi_RVALID;
	output axi_RREADY;
	input axi_RLAST;
	output [31:0] axi_io_AW;
	output axi_io_AWVALID;
	input axi_io_AWREADY;
	output [1:0] axi_io_AWBURST;
	output [7:0] axi_io_AWLEN;
	output [2:0] axi_io_AWSIZE;
	output [31:0] axi_io_W;
	output axi_io_WVALID;
	input axi_io_WREADY;
	output [3:0] axi_io_WSTRB;
	output axi_io_WLAST;
	output [31:0] axi_io_AR;
	output axi_io_ARVALID;
	input axi_io_ARREADY;
	output [1:0] axi_io_ARBURST;
	output [7:0] axi_io_ARLEN;
	output [2:0] axi_io_ARSIZE;
	input [31:0] axi_io_R;
	input axi_io_RVALID;
	output axi_io_RREADY;
	input axi_io_RLAST;
	output busy;
	input outstanding;

	wire [1:0] A4;
	wire [4:0] fsm;
	wire [4:0] burst_idx;
	wire [9:0] cacheA;
	wire [149:0] cacheQ;
	wire [149:0] cacheD;
	wire [15:0] cacheM;



	notech_inv i_15718(.A(n_62052), .Z(n_62053));
	notech_inv i_15717(.A(n_62045), .Z(n_62052));
	notech_inv i_15716(.A(n_62050), .Z(n_62051));
	notech_inv i_15715(.A(n_62037), .Z(n_62050));
	notech_inv i_15714(.A(n_62048), .Z(n_62049));
	notech_inv i_15713(.A(n_62033), .Z(n_62048));
	notech_inv i_15712(.A(n_62046), .Z(n_62047));
	notech_inv i_15711(.A(n_62031), .Z(n_62046));
	notech_inv i_15710(.A(n_62044), .Z(n_62045));
	notech_inv i_15709(.A(n_62029), .Z(n_62044));
	notech_inv i_15708(.A(n_62042), .Z(n_62043));
	notech_inv i_15707(.A(n_62021), .Z(n_62042));
	notech_inv i_15706(.A(n_62040), .Z(n_62041));
	notech_inv i_15705(.A(n_62019), .Z(n_62040));
	notech_inv i_15704(.A(n_62038), .Z(n_62039));
	notech_inv i_15703(.A(n_62017), .Z(n_62038));
	notech_inv i_15702(.A(n_62036), .Z(n_62037));
	notech_inv i_15701(.A(n_62015), .Z(n_62036));
	notech_inv i_15700(.A(n_62034), .Z(n_62035));
	notech_inv i_15699(.A(n_62013), .Z(n_62034));
	notech_inv i_15698(.A(n_62032), .Z(n_62033));
	notech_inv i_15697(.A(n_62011), .Z(n_62032));
	notech_inv i_15696(.A(n_62030), .Z(n_62031));
	notech_inv i_15695(.A(n_62009), .Z(n_62030));
	notech_inv i_15694(.A(n_62028), .Z(n_62029));
	notech_inv i_15693(.A(n_62047), .Z(n_62028));
	notech_inv i_15692(.A(n_62026), .Z(n_62027));
	notech_inv i_15691(.A(n_62003), .Z(n_62026));
	notech_inv i_15690(.A(n_62024), .Z(n_62025));
	notech_inv i_15689(.A(n_61999), .Z(n_62024));
	notech_inv i_15688(.A(n_62022), .Z(n_62023));
	notech_inv i_15687(.A(n_61997), .Z(n_62022));
	notech_inv i_15686(.A(n_62020), .Z(n_62021));
	notech_inv i_15685(.A(n_62023), .Z(n_62020));
	notech_inv i_15684(.A(n_62018), .Z(n_62019));
	notech_inv i_15683(.A(n_61993), .Z(n_62018));
	notech_inv i_15682(.A(n_62016), .Z(n_62017));
	notech_inv i_15681(.A(n_61991), .Z(n_62016));
	notech_inv i_15680(.A(n_62014), .Z(n_62015));
	notech_inv i_15679(.A(n_62039), .Z(n_62014));
	notech_inv i_15678(.A(n_62012), .Z(n_62013));
	notech_inv i_15677(.A(n_61989), .Z(n_62012));
	notech_inv i_15676(.A(n_62010), .Z(n_62011));
	notech_inv i_15675(.A(n_62035), .Z(n_62010));
	notech_inv i_15674(.A(n_62008), .Z(n_62009));
	notech_inv i_15673(.A(n_62049), .Z(n_62008));
	notech_inv i_15672(.A(n_62006), .Z(n_62007));
	notech_inv i_15671(.A(n_61985), .Z(n_62006));
	notech_inv i_15670(.A(n_62004), .Z(n_62005));
	notech_inv i_15669(.A(n_61983), .Z(n_62004));
	notech_inv i_15668(.A(n_62002), .Z(n_62003));
	notech_inv i_15667(.A(n_62005), .Z(n_62002));
	notech_inv i_15666(.A(n_62000), .Z(n_62001));
	notech_inv i_15665(.A(n_61981), .Z(n_62000));
	notech_inv i_15664(.A(n_61998), .Z(n_61999));
	notech_inv i_15663(.A(n_62001), .Z(n_61998));
	notech_inv i_15662(.A(n_61996), .Z(n_61997));
	notech_inv i_15661(.A(n_62025), .Z(n_61996));
	notech_inv i_15660(.A(n_61994), .Z(n_61995));
	notech_inv i_15659(.A(n_61979), .Z(n_61994));
	notech_inv i_15658(.A(n_61992), .Z(n_61993));
	notech_inv i_15657(.A(n_61995), .Z(n_61992));
	notech_inv i_15656(.A(n_61990), .Z(n_61991));
	notech_inv i_15655(.A(n_62041), .Z(n_61990));
	notech_inv i_15654(.A(n_61988), .Z(n_61989));
	notech_inv i_15653(.A(n_62051), .Z(n_61988));
	notech_inv i_15652(.A(n_61986), .Z(n_61987));
	notech_inv i_15651(.A(clk), .Z(n_61986));
	notech_inv i_15650(.A(n_61984), .Z(n_61985));
	notech_inv i_15649(.A(n_61987), .Z(n_61984));
	notech_inv i_15648(.A(n_61982), .Z(n_61983));
	notech_inv i_15647(.A(n_62007), .Z(n_61982));
	notech_inv i_15646(.A(n_61980), .Z(n_61981));
	notech_inv i_15645(.A(n_62027), .Z(n_61980));
	notech_inv i_15644(.A(n_61978), .Z(n_61979));
	notech_inv i_15643(.A(n_62043), .Z(n_61978));
	notech_inv i_15194(.A(n_61517), .Z(n_61529));
	notech_inv i_15193(.A(n_61517), .Z(n_61528));
	notech_inv i_15188(.A(n_61517), .Z(n_61523));
	notech_inv i_15183(.A(n_61517), .Z(n_61518));
	notech_inv i_15182(.A(n_2008), .Z(n_61517));
	notech_inv i_15179(.A(n_61501), .Z(n_61513));
	notech_inv i_15178(.A(n_61501), .Z(n_61512));
	notech_inv i_15173(.A(n_61501), .Z(n_61507));
	notech_inv i_15168(.A(n_61501), .Z(n_61502));
	notech_inv i_15167(.A(n_1996), .Z(n_61501));
	notech_inv i_15163(.A(n_61490), .Z(n_61496));
	notech_inv i_15158(.A(n_61490), .Z(n_61491));
	notech_inv i_15157(.A(n_968), .Z(n_61490));
	notech_inv i_15154(.A(n_61474), .Z(n_61486));
	notech_inv i_15153(.A(n_61474), .Z(n_61485));
	notech_inv i_15148(.A(n_61474), .Z(n_61480));
	notech_inv i_15143(.A(n_61474), .Z(n_61475));
	notech_inv i_15142(.A(n_972), .Z(n_61474));
	notech_inv i_14795(.A(n_61436), .Z(n_61442));
	notech_inv i_14790(.A(n_61436), .Z(n_61437));
	notech_inv i_14789(.A(n_2004), .Z(n_61436));
	notech_inv i_14788(.A(n_61414), .Z(n_61434));
	notech_inv i_14787(.A(n_61414), .Z(n_61433));
	notech_inv i_14786(.A(n_61414), .Z(n_61432));
	notech_inv i_14785(.A(n_61414), .Z(n_61431));
	notech_inv i_14784(.A(n_61414), .Z(n_61430));
	notech_inv i_14783(.A(n_61414), .Z(n_61429));
	notech_inv i_14781(.A(n_61414), .Z(n_61427));
	notech_inv i_14780(.A(n_61414), .Z(n_61426));
	notech_inv i_14779(.A(n_61414), .Z(n_61425));
	notech_inv i_14778(.A(n_61414), .Z(n_61424));
	notech_inv i_14777(.A(n_61414), .Z(n_61423));
	notech_inv i_14776(.A(n_61414), .Z(n_61422));
	notech_inv i_14774(.A(n_61414), .Z(n_61420));
	notech_inv i_14773(.A(n_61414), .Z(n_61419));
	notech_inv i_14772(.A(n_61414), .Z(n_61418));
	notech_inv i_14771(.A(n_61414), .Z(n_61417));
	notech_inv i_14770(.A(n_61414), .Z(n_61416));
	notech_inv i_14769(.A(n_61414), .Z(n_61415));
	notech_inv i_14768(.A(rstn), .Z(n_61414));
	notech_inv i_14233(.A(n_60872), .Z(n_60873));
	notech_inv i_14232(.A(n_2033), .Z(n_60872));
	notech_inv i_14225(.A(n_60863), .Z(n_60864));
	notech_inv i_14224(.A(n_2010), .Z(n_60863));
	notech_inv i_14215(.A(n_60852), .Z(n_60853));
	notech_inv i_14214(.A(n_1067), .Z(n_60852));
	notech_inv i_14207(.A(n_60843), .Z(n_60844));
	notech_inv i_14206(.A(n_1061), .Z(n_60843));
	notech_inv i_14199(.A(n_60834), .Z(n_60835));
	notech_inv i_14198(.A(n_2023), .Z(n_60834));
	notech_inv i_14191(.A(n_60825), .Z(n_60826));
	notech_inv i_14190(.A(n_6652), .Z(n_60825));
	notech_inv i_14183(.A(n_60816), .Z(n_60817));
	notech_inv i_14182(.A(n_6673), .Z(n_60816));
	notech_inv i_14175(.A(n_60803), .Z(n_60808));
	notech_inv i_14171(.A(n_60803), .Z(n_60804));
	notech_inv i_14170(.A(\nbus_11662[0] ), .Z(n_60803));
	notech_inv i_13822(.A(n_60427), .Z(n_60429));
	notech_inv i_13821(.A(n_60427), .Z(code_data[0]));
	notech_inv i_13820(.A(\nbus_14528[0] ), .Z(n_60427));
	notech_inv i_13047(.A(n_59556), .Z(n_59557));
	notech_inv i_13046(.A(n_1277), .Z(n_59556));
	notech_inv i_13037(.A(n_59545), .Z(n_59546));
	notech_inv i_13036(.A(n_1375), .Z(n_59545));
	notech_inv i_13029(.A(n_59532), .Z(n_59537));
	notech_inv i_13025(.A(n_59532), .Z(n_59533));
	notech_inv i_13024(.A(A4[1]), .Z(n_59532));
	notech_inv i_13020(.A(n_59513), .Z(n_59527));
	notech_inv i_13019(.A(n_59513), .Z(n_59526));
	notech_inv i_13013(.A(n_59513), .Z(n_59520));
	notech_inv i_13007(.A(n_59513), .Z(n_59514));
	notech_inv i_13006(.A(n_2072), .Z(n_59513));
	notech_inv i_13004(.A(n_59497), .Z(n_59510));
	notech_inv i_13002(.A(n_59497), .Z(n_59508));
	notech_inv i_12998(.A(n_59497), .Z(n_59504));
	notech_inv i_12997(.A(n_59497), .Z(n_59503));
	notech_inv i_12992(.A(n_59497), .Z(n_59498));
	notech_inv i_12991(.A(A4[0]), .Z(n_59497));
	notech_inv i_12987(.A(n_59478), .Z(n_59492));
	notech_inv i_12986(.A(n_59478), .Z(n_59491));
	notech_inv i_12980(.A(n_59478), .Z(n_59485));
	notech_inv i_12974(.A(n_59478), .Z(n_59479));
	notech_inv i_12973(.A(n_2074), .Z(n_59478));
	notech_inv i_12971(.A(n_59503), .Z(n_59475));
	notech_inv i_12969(.A(n_59503), .Z(n_59473));
	notech_inv i_12966(.A(n_59503), .Z(n_59470));
	notech_inv i_12964(.A(n_59503), .Z(n_59468));
	notech_inv i_12961(.A(n_59503), .Z(n_59465));
	notech_inv i_12959(.A(n_59503), .Z(n_59463));
	notech_inv i_12949(.A(n_59451), .Z(n_59452));
	notech_inv i_12948(.A(n_1377), .Z(n_59451));
	notech_inv i_12939(.A(n_59440), .Z(n_59441));
	notech_inv i_12938(.A(n_1474), .Z(n_59440));
	notech_inv i_12929(.A(n_59429), .Z(n_59430));
	notech_inv i_12928(.A(n_1476), .Z(n_59429));
	notech_inv i_12919(.A(n_59418), .Z(n_59419));
	notech_inv i_12918(.A(n_1573), .Z(n_59418));
	notech_inv i_12909(.A(n_59407), .Z(n_59408));
	notech_inv i_12908(.A(n_1575), .Z(n_59407));
	notech_inv i_12899(.A(n_59396), .Z(n_59397));
	notech_inv i_12898(.A(n_1703), .Z(n_59396));
	notech_inv i_12889(.A(n_59385), .Z(n_59386));
	notech_inv i_12888(.A(n_1705), .Z(n_59385));
	notech_inv i_10340(.A(n_56597), .Z(n_56598));
	notech_inv i_10339(.A(\nbus_11667[0] ), .Z(n_56597));
	notech_inv i_7961(.A(n_53872), .Z(n_53873));
	notech_inv i_7960(.A(\nbus_11671[0] ), .Z(n_53872));
	notech_inv i_7839(.A(n_53693), .Z(n_53694));
	notech_inv i_7838(.A(\nbus_11667[96] ), .Z(n_53693));
	notech_inv i_7829(.A(n_53682), .Z(n_53683));
	notech_inv i_7828(.A(\nbus_11667[64] ), .Z(n_53682));
	notech_inv i_7819(.A(n_53671), .Z(n_53672));
	notech_inv i_7818(.A(\nbus_11667[32] ), .Z(n_53671));
	notech_inv i_7738(.A(n_53547), .Z(n_53548));
	notech_inv i_7737(.A(n_2244), .Z(n_53547));
	notech_inv i_7728(.A(n_53536), .Z(n_53537));
	notech_inv i_7727(.A(n_2239), .Z(n_53536));
	notech_inv i_7720(.A(n_53483), .Z(n_53484));
	notech_inv i_7719(.A(n_2237), .Z(n_53483));
	notech_ao4 i_56395(.A(n_1061), .B(n_6834), .C(n_2010), .D(n_6872), .Z(n_986
		));
	notech_ao4 i_56401(.A(n_1061), .B(n_6835), .C(n_2010), .D(n_6873), .Z(n_983
		));
	notech_ao4 i_56407(.A(n_1061), .B(n_6836), .C(n_2010), .D(n_6874), .Z(n_980
		));
	notech_and4 i_57641(.A(n_61528), .B(n_61442), .C(n_973), .D(n_976), .Z(n_977
		));
	notech_nand3 i_151(.A(axi_RVALID), .B(axi_RLAST), .C(n_22749), .Z(n_976)
		);
	notech_ao3 i_58570(.A(n_61485), .B(n_973), .C(n_974), .Z(n_975));
	notech_and2 i_147(.A(axi_WREADY), .B(n_25082), .Z(n_974));
	notech_and2 i_45(.A(n_1215), .B(n_2010), .Z(n_973));
	notech_and3 i_50(.A(n_61528), .B(n_61496), .C(n_6763), .Z(n_972));
	notech_nor2 i_137(.A(code_ack), .B(n_7004), .Z(n_971));
	notech_nor2 i_136(.A(read_ack), .B(n_7005), .Z(n_970));
	notech_nao3 i_64(.A(n_6765), .B(n_6768), .C(n_2000), .Z(busy));
	notech_and2 i_11(.A(n_61512), .B(n_6665), .Z(n_968));
	notech_xor2 i_132(.A(burst_idx[4]), .B(n_2027), .Z(n_967));
	notech_xor2 i_131(.A(burst_idx[3]), .B(n_2026), .Z(n_966));
	notech_xor2 i_130(.A(burst_idx[2]), .B(n_2025), .Z(n_965));
	notech_nand2 i_127(.A(n_1215), .B(n_6763), .Z(n_963));
	notech_xor2 i_1879479(.A(axi_AR[14]), .B(cacheQ[128]), .Z(n_960));
	notech_xor2 i_1979480(.A(axi_AR[15]), .B(cacheQ[129]), .Z(n_959));
	notech_xor2 i_20(.A(axi_AR[16]), .B(cacheQ[130]), .Z(n_958));
	notech_xor2 i_2179481(.A(axi_AR[17]), .B(cacheQ[131]), .Z(n_957));
	notech_xor2 i_2279482(.A(axi_AR[18]), .B(cacheQ[132]), .Z(n_956));
	notech_xor2 i_2379483(.A(axi_AR[19]), .B(cacheQ[133]), .Z(n_955));
	notech_xor2 i_24(.A(axi_AR[20]), .B(cacheQ[134]), .Z(n_954));
	notech_xor2 i_25(.A(axi_AR[21]), .B(cacheQ[135]), .Z(n_953));
	notech_xor2 i_2679484(.A(axi_AR[22]), .B(cacheQ[136]), .Z(n_952));
	notech_xor2 i_2779485(.A(axi_AR[23]), .B(cacheQ[137]), .Z(n_951));
	notech_xor2 i_28(.A(axi_AR[24]), .B(cacheQ[138]), .Z(n_950));
	notech_xor2 i_2979486(.A(axi_AR[25]), .B(cacheQ[139]), .Z(n_949));
	notech_xor2 i_3079487(.A(axi_AR[26]), .B(cacheQ[140]), .Z(n_948));
	notech_xor2 i_3179488(.A(axi_AR[27]), .B(cacheQ[141]), .Z(n_947));
	notech_xor2 i_3279489(.A(axi_AR[28]), .B(cacheQ[142]), .Z(n_946));
	notech_xor2 i_3379490(.A(axi_AR[29]), .B(cacheQ[143]), .Z(n_945));
	notech_xor2 i_3479491(.A(axi_AR[30]), .B(cacheQ[144]), .Z(n_944));
	notech_xor2 i_3579492(.A(axi_AR[31]), .B(cacheQ[145]), .Z(n_943));
	notech_or4 i_4779502(.A(n_960), .B(n_959), .C(n_958), .D(n_957), .Z(n_934
		));
	notech_or4 i_4879503(.A(n_956), .B(n_955), .C(n_954), .D(n_953), .Z(n_933
		));
	notech_or4 i_4979504(.A(n_952), .B(n_951), .C(n_950), .D(n_949), .Z(n_932
		));
	notech_or4 i_5079505(.A(n_948), .B(n_947), .C(n_946), .D(n_945), .Z(n_931
		));
	notech_or4 i_5579508(.A(n_934), .B(n_933), .C(n_932), .D(n_931), .Z(n_928
		));
	notech_xor2 i_1879528(.A(cacheQ[128]), .B(axi_AW[14]), .Z(n_926));
	notech_xor2 i_1979529(.A(cacheQ[129]), .B(axi_AW[15]), .Z(n_925));
	notech_xor2 i_2079530(.A(cacheQ[130]), .B(axi_AW[16]), .Z(n_924));
	notech_xor2 i_2179531(.A(cacheQ[131]), .B(axi_AW[17]), .Z(n_923));
	notech_xor2 i_2279532(.A(cacheQ[132]), .B(axi_AW[18]), .Z(n_922));
	notech_xor2 i_2379533(.A(cacheQ[133]), .B(axi_AW[19]), .Z(n_921));
	notech_xor2 i_2479534(.A(cacheQ[134]), .B(axi_AW[20]), .Z(n_920));
	notech_xor2 i_2579535(.A(cacheQ[135]), .B(axi_AW[21]), .Z(n_919));
	notech_xor2 i_2679536(.A(cacheQ[136]), .B(axi_AW[22]), .Z(n_918));
	notech_xor2 i_2779537(.A(cacheQ[137]), .B(axi_AW[23]), .Z(n_917));
	notech_xor2 i_2879538(.A(cacheQ[138]), .B(axi_AW[24]), .Z(n_916));
	notech_xor2 i_2979539(.A(cacheQ[139]), .B(axi_AW[25]), .Z(n_915));
	notech_xor2 i_3079540(.A(cacheQ[140]), .B(axi_AW[26]), .Z(n_914));
	notech_xor2 i_3179541(.A(cacheQ[141]), .B(axi_AW[27]), .Z(n_913));
	notech_xor2 i_3279542(.A(cacheQ[142]), .B(axi_AW[28]), .Z(n_912));
	notech_xor2 i_3379543(.A(cacheQ[143]), .B(axi_AW[29]), .Z(n_911));
	notech_xor2 i_3479544(.A(n_6995), .B(axi_AW[30]), .Z(n_910));
	notech_xor2 i_3579545(.A(n_6996), .B(axi_AW[31]), .Z(n_909));
	notech_or4 i_4779555(.A(n_926), .B(n_925), .C(n_924), .D(n_923), .Z(n_900
		));
	notech_or4 i_4879556(.A(n_922), .B(n_921), .C(n_920), .D(n_919), .Z(n_899
		));
	notech_or4 i_4979557(.A(n_918), .B(n_917), .C(n_916), .D(n_915), .Z(n_898
		));
	notech_or4 i_5079558(.A(n_914), .B(n_913), .C(n_912), .D(n_911), .Z(n_897
		));
	notech_or4 i_5579561(.A(n_900), .B(n_899), .C(n_898), .D(n_897), .Z(n_894
		));
	notech_ao4 i_56389(.A(n_1061), .B(n_6833), .C(n_2010), .D(n_6871), .Z(n_989
		));
	notech_ao4 i_56383(.A(n_1061), .B(n_6832), .C(n_2010), .D(n_6870), .Z(n_992
		));
	notech_ao4 i_56377(.A(n_1061), .B(n_6831), .C(n_2010), .D(n_6869), .Z(n_995
		));
	notech_ao4 i_56371(.A(n_1061), .B(n_6830), .C(n_2010), .D(n_6868), .Z(n_998
		));
	notech_ao4 i_56365(.A(n_1061), .B(n_6829), .C(n_2010), .D(n_6867), .Z(n_1001
		));
	notech_ao4 i_56359(.A(n_1061), .B(n_6828), .C(n_2010), .D(n_6866), .Z(n_1004
		));
	notech_ao4 i_56353(.A(n_1061), .B(n_6827), .C(n_2010), .D(n_6865), .Z(n_1007
		));
	notech_ao4 i_56347(.A(n_1061), .B(n_6826), .C(n_2010), .D(n_6864), .Z(n_1010
		));
	notech_ao4 i_56341(.A(n_1061), .B(n_6825), .C(n_2010), .D(n_6863), .Z(n_1013
		));
	notech_ao4 i_56335(.A(n_1061), .B(n_6824), .C(n_2010), .D(n_6862), .Z(n_1016
		));
	notech_ao4 i_56329(.A(n_1061), .B(n_6823), .C(n_2010), .D(n_6861), .Z(n_1019
		));
	notech_ao4 i_56323(.A(n_60844), .B(n_6822), .C(n_2010), .D(n_6860), .Z(n_1022
		));
	notech_ao4 i_56317(.A(n_60844), .B(n_6821), .C(n_2010), .D(n_6859), .Z(n_1025
		));
	notech_ao4 i_56311(.A(n_60844), .B(n_6820), .C(n_2010), .D(n_6858), .Z(n_1028
		));
	notech_ao4 i_56305(.A(n_60844), .B(n_6819), .C(n_60864), .D(n_6857), .Z(n_1031
		));
	notech_ao4 i_56299(.A(n_60844), .B(n_6809), .C(n_60864), .D(n_6856), .Z(n_1034
		));
	notech_ao4 i_56293(.A(n_60844), .B(n_6810), .C(n_60864), .D(n_6855), .Z(n_1037
		));
	notech_ao4 i_56287(.A(n_60844), .B(n_6811), .C(n_60864), .D(n_6854), .Z(n_1040
		));
	notech_ao4 i_56281(.A(n_60844), .B(n_6812), .C(n_60864), .D(n_6853), .Z(n_1043
		));
	notech_ao4 i_56275(.A(n_60844), .B(n_6813), .C(n_60864), .D(n_6852), .Z(n_1046
		));
	notech_ao4 i_56269(.A(n_1061), .B(n_6814), .C(n_60864), .D(n_6851), .Z(n_1049
		));
	notech_ao4 i_56263(.A(n_60844), .B(n_6815), .C(n_60864), .D(n_6850), .Z(n_1052
		));
	notech_ao4 i_56257(.A(n_60844), .B(n_6816), .C(n_60864), .D(n_6849), .Z(n_1055
		));
	notech_ao4 i_56251(.A(n_60844), .B(n_6817), .C(n_60864), .D(n_6848), .Z(n_1058
		));
	notech_and3 i_32(.A(n_2019), .B(n_1215), .C(n_61496), .Z(n_1061));
	notech_ao4 i_56245(.A(n_60844), .B(n_6818), .C(n_60864), .D(n_6847), .Z(n_1062
		));
	notech_ao4 i_56239(.A(n_2020), .B(n_6808), .C(n_60864), .D(n_6846), .Z(n_1065
		));
	notech_nao3 i_242(.A(axi_AR[30]), .B(n_6999), .C(n_2019), .Z(n_1066));
	notech_and4 i_58500(.A(n_1215), .B(n_60864), .C(n_1066), .D(n_61496), .Z
		(n_1067));
	notech_ao4 i_56234(.A(n_2020), .B(n_6807), .C(n_60864), .D(n_6845), .Z(n_1070
		));
	notech_ao4 i_56558(.A(n_61528), .B(n_6874), .C(n_61442), .D(n_6836), .Z(n_1073
		));
	notech_ao4 i_56553(.A(n_61528), .B(n_6873), .C(n_61442), .D(n_6835), .Z(n_1076
		));
	notech_ao4 i_56548(.A(n_61528), .B(n_6872), .C(n_61442), .D(n_6834), .Z(n_1079
		));
	notech_ao4 i_56543(.A(n_61528), .B(n_6871), .C(n_61442), .D(n_6833), .Z(n_1082
		));
	notech_ao4 i_56538(.A(n_61528), .B(n_6870), .C(n_61442), .D(n_6832), .Z(n_1085
		));
	notech_ao4 i_56533(.A(n_61528), .B(n_6869), .C(n_61442), .D(n_6831), .Z(n_1088
		));
	notech_ao4 i_56528(.A(n_61528), .B(n_6868), .C(n_61442), .D(n_6830), .Z(n_1091
		));
	notech_ao4 i_56523(.A(n_61528), .B(n_6867), .C(n_61442), .D(n_6829), .Z(n_1094
		));
	notech_ao4 i_56518(.A(n_61528), .B(n_6866), .C(n_61442), .D(n_6828), .Z(n_1097
		));
	notech_ao4 i_56513(.A(n_61528), .B(n_6865), .C(n_61442), .D(n_6827), .Z(n_1100
		));
	notech_ao4 i_56508(.A(n_61528), .B(n_6864), .C(n_61442), .D(n_6826), .Z(n_1103
		));
	notech_ao4 i_56503(.A(n_61528), .B(n_6863), .C(n_61442), .D(n_6825), .Z(n_1106
		));
	notech_ao4 i_56498(.A(n_61528), .B(n_6862), .C(n_61442), .D(n_6824), .Z(n_1109
		));
	notech_ao4 i_56493(.A(n_61528), .B(n_6861), .C(n_61442), .D(n_6823), .Z(n_1112
		));
	notech_ao4 i_56488(.A(n_61528), .B(n_6860), .C(n_61442), .D(n_6822), .Z(n_1115
		));
	notech_ao4 i_56483(.A(n_61528), .B(n_6859), .C(n_61442), .D(n_6821), .Z(n_1118
		));
	notech_ao4 i_56478(.A(n_61529), .B(n_6858), .C(n_61442), .D(n_6820), .Z(n_1121
		));
	notech_ao4 i_56473(.A(n_61529), .B(n_6857), .C(n_61442), .D(n_6819), .Z(n_1124
		));
	notech_ao4 i_56468(.A(n_61529), .B(n_6856), .C(n_61442), .D(n_6809), .Z(n_1127
		));
	notech_ao4 i_56463(.A(n_61529), .B(n_6855), .C(n_61437), .D(n_6810), .Z(n_1130
		));
	notech_ao4 i_56458(.A(n_61529), .B(n_6854), .C(n_61437), .D(n_6811), .Z(n_1133
		));
	notech_ao4 i_56453(.A(n_61529), .B(n_6853), .C(n_61437), .D(n_6812), .Z(n_1136
		));
	notech_ao4 i_56448(.A(n_61529), .B(n_6852), .C(n_61437), .D(n_6813), .Z(n_1139
		));
	notech_ao4 i_56443(.A(n_61529), .B(n_6851), .C(n_61437), .D(n_6814), .Z(n_1142
		));
	notech_ao4 i_56438(.A(n_61529), .B(n_6850), .C(n_61437), .D(n_6815), .Z(n_1145
		));
	notech_ao4 i_56433(.A(n_61529), .B(n_6849), .C(n_61437), .D(n_6816), .Z(n_1148
		));
	notech_ao4 i_56428(.A(n_61529), .B(n_6848), .C(n_61437), .D(n_6817), .Z(n_1151
		));
	notech_ao4 i_56423(.A(n_61529), .B(n_6847), .C(n_61437), .D(n_6818), .Z(n_1154
		));
	notech_ao4 i_56418(.A(n_61529), .B(n_6846), .C(n_61437), .D(n_6808), .Z(n_1157
		));
	notech_ao4 i_56413(.A(n_61529), .B(n_6845), .C(n_61437), .D(n_6807), .Z(n_1160
		));
	notech_nao3 i_348(.A(n_2033), .B(n_2035), .C(n_2040), .Z(n_1167));
	notech_and3 i_126(.A(n_6763), .B(n_973), .C(n_1167), .Z(n_1170));
	notech_ao4 i_58875(.A(n_1170), .B(n_7001), .C(n_2024), .D(n_2030), .Z(n_1171
		));
	notech_ao4 i_56563(.A(n_2024), .B(burst_idx[0]), .C(n_2032), .D(n_2000),
		 .Z(n_1173));
	notech_nand2 i_354(.A(axi_AWREADY), .B(n_6669), .Z(n_1174));
	notech_and4 i_57295(.A(n_61529), .B(n_61496), .C(n_6763), .D(n_1174), .Z
		(n_1175));
	notech_nand2 i_105(.A(n_61529), .B(n_6763), .Z(n_1176));
	notech_ao4 i_56627(.A(n_61529), .B(n_6844), .C(n_61437), .D(n_6882), .Z(n_1179
		));
	notech_ao4 i_56622(.A(n_61529), .B(n_6843), .C(n_61437), .D(n_6881), .Z(n_1182
		));
	notech_ao4 i_56617(.A(n_61518), .B(n_6842), .C(n_61437), .D(n_6880), .Z(n_1185
		));
	notech_ao4 i_56612(.A(n_61518), .B(n_6841), .C(n_61437), .D(n_6879), .Z(n_1188
		));
	notech_ao4 i_56607(.A(n_61518), .B(n_6840), .C(n_61437), .D(n_6878), .Z(n_1191
		));
	notech_ao4 i_56602(.A(n_61518), .B(n_6839), .C(n_61437), .D(n_6877), .Z(n_1194
		));
	notech_ao4 i_56597(.A(n_61518), .B(n_6838), .C(n_61437), .D(n_6876), .Z(n_1197
		));
	notech_ao4 i_56592(.A(n_61518), .B(n_6837), .C(n_61437), .D(n_6875), .Z(n_1200
		));
	notech_and4 i_59042(.A(n_2046), .B(n_61496), .C(n_6763), .D(n_973), .Z(n_1203
		));
	notech_nand2 i_56726(.A(n_2045), .B(n_6705), .Z(n_1204));
	notech_or2 i_389(.A(n_1995), .B(n_2017), .Z(n_1205));
	notech_nao3 i_391(.A(read_req), .B(n_2052), .C(n_2045), .Z(n_1207));
	notech_and4 i_57932(.A(n_61485), .B(n_2051), .C(n_973), .D(n_1207), .Z(n_1208
		));
	notech_or2 i_396(.A(abort), .B(n_2045), .Z(n_1209));
	notech_nand3 i_56729(.A(n_2019), .B(n_1205), .C(n_1209), .Z(n_1210));
	notech_ao3 i_57886(.A(n_61485), .B(n_973), .C(n_2033), .Z(n_1211));
	notech_nand3 i_56741(.A(n_60864), .B(n_2058), .C(n_61518), .Z(n_1212));
	notech_and4 i_56739(.A(n_2061), .B(n_61518), .C(n_2024), .D(n_2056), .Z(n_1213
		));
	notech_nand2 i_56738(.A(n_1066), .B(n_2058), .Z(n_1214));
	notech_or4 i_60(.A(read_ack), .B(n_2003), .C(busy), .D(n_7005), .Z(n_1215
		));
	notech_nao3 i_56736(.A(n_1215), .B(n_2058), .C(n_1221), .Z(n_1216));
	notech_nand2 i_410(.A(axi_WREADY), .B(n_6669), .Z(n_1217));
	notech_and4 i_57916(.A(n_61518), .B(n_1217), .C(n_61496), .D(n_6763), .Z
		(n_1218));
	notech_ao3 i_61(.A(fsm[3]), .B(fsm[0]), .C(n_2000), .Z(n_1221));
	notech_and4 i_58102(.A(n_61485), .B(n_2064), .C(n_2066), .D(n_1217), .Z(n_1222
		));
	notech_and4 i_56734(.A(n_2024), .B(n_6763), .C(n_2057), .D(n_973), .Z(n_1223
		));
	notech_nand2 i_57210(.A(n_6652), .B(n_6661), .Z(n_1224));
	notech_ao4 i_57204(.A(n_6652), .B(n_6836), .C(n_6996), .D(n_6661), .Z(n_1227
		));
	notech_ao4 i_57201(.A(n_6652), .B(n_6835), .C(n_6995), .D(n_6661), .Z(n_1230
		));
	notech_ao4 i_57198(.A(n_6652), .B(n_6834), .C(n_6661), .D(n_6994), .Z(n_1233
		));
	notech_ao4 i_57195(.A(n_6652), .B(n_6833), .C(n_6661), .D(n_6993), .Z(n_1236
		));
	notech_ao4 i_57192(.A(n_6652), .B(n_6832), .C(n_6661), .D(n_6992), .Z(n_1239
		));
	notech_ao4 i_57189(.A(n_6652), .B(n_6831), .C(n_6661), .D(n_6991), .Z(n_1242
		));
	notech_ao4 i_57186(.A(n_6652), .B(n_6830), .C(n_6661), .D(n_6990), .Z(n_1245
		));
	notech_ao4 i_57183(.A(n_6652), .B(n_6829), .C(n_6661), .D(n_6989), .Z(n_1248
		));
	notech_ao4 i_57180(.A(n_6652), .B(n_6828), .C(n_6661), .D(n_6988), .Z(n_1251
		));
	notech_ao4 i_57177(.A(n_6652), .B(n_6827), .C(n_6661), .D(n_6987), .Z(n_1254
		));
	notech_ao4 i_57174(.A(n_6652), .B(n_6826), .C(n_6661), .D(n_6986), .Z(n_1257
		));
	notech_ao4 i_57171(.A(n_60826), .B(n_6825), .C(n_6661), .D(n_6985), .Z(n_1260
		));
	notech_ao4 i_57168(.A(n_60826), .B(n_6824), .C(n_6661), .D(n_6984), .Z(n_1263
		));
	notech_ao4 i_57165(.A(n_60826), .B(n_6823), .C(n_6661), .D(n_6983), .Z(n_1266
		));
	notech_ao4 i_57162(.A(n_60826), .B(n_6822), .C(n_6661), .D(n_6982), .Z(n_1269
		));
	notech_ao4 i_57159(.A(n_60826), .B(n_6821), .C(n_6661), .D(n_6981), .Z(n_1272
		));
	notech_ao4 i_57156(.A(n_60826), .B(n_6820), .C(n_6661), .D(n_6980), .Z(n_1275
		));
	notech_ao4 i_57714(.A(n_60826), .B(n_2071), .C(n_2070), .D(n_7001), .Z(n_1277
		));
	notech_ao4 i_57153(.A(n_60826), .B(n_6819), .C(n_6661), .D(n_6979), .Z(n_1280
		));
	notech_nand2 i_480(.A(cacheQ[127]), .B(n_1377), .Z(n_1281));
	notech_nand3 i_479(.A(n_59526), .B(axi_W[31]), .C(n_59508), .Z(n_1282)
		);
	notech_nand3 i_57150(.A(n_1282), .B(n_1579), .C(n_1281), .Z(n_1283));
	notech_nand2 i_484(.A(n_1377), .B(cacheQ[126]), .Z(n_1284));
	notech_nand3 i_483(.A(n_59526), .B(axi_W[30]), .C(n_59508), .Z(n_1285)
		);
	notech_nand3 i_57147(.A(n_1285), .B(n_1583), .C(n_1284), .Z(n_1286));
	notech_nand2 i_488(.A(n_1377), .B(cacheQ[125]), .Z(n_1287));
	notech_nand3 i_487(.A(n_59526), .B(axi_W[29]), .C(n_59504), .Z(n_1288)
		);
	notech_nand3 i_57144(.A(n_1288), .B(n_1587), .C(n_1287), .Z(n_1289));
	notech_nand2 i_492(.A(n_1377), .B(cacheQ[124]), .Z(n_1290));
	notech_nand3 i_491(.A(n_59526), .B(axi_W[28]), .C(n_59508), .Z(n_1291)
		);
	notech_nand3 i_57141(.A(n_1291), .B(n_1591), .C(n_1290), .Z(n_1292));
	notech_nand2 i_496(.A(n_1377), .B(cacheQ[123]), .Z(n_1293));
	notech_nand3 i_495(.A(n_59526), .B(axi_W[27]), .C(n_59508), .Z(n_1294)
		);
	notech_nand3 i_57138(.A(n_1294), .B(n_1595), .C(n_1293), .Z(n_1295));
	notech_nand2 i_500(.A(n_1377), .B(cacheQ[122]), .Z(n_1296));
	notech_nand3 i_499(.A(n_59527), .B(axi_W[26]), .C(n_59508), .Z(n_1297)
		);
	notech_nand3 i_57135(.A(n_1297), .B(n_1599), .C(n_1296), .Z(n_1298));
	notech_nand2 i_504(.A(n_1377), .B(cacheQ[121]), .Z(n_1299));
	notech_nand3 i_503(.A(n_59527), .B(axi_W[25]), .C(n_59508), .Z(n_1300)
		);
	notech_nand3 i_57132(.A(n_1300), .B(n_1603), .C(n_1299), .Z(n_1301));
	notech_nand2 i_508(.A(n_1377), .B(cacheQ[120]), .Z(n_1302));
	notech_nand3 i_507(.A(n_59526), .B(axi_W[24]), .C(n_59508), .Z(n_1303)
		);
	notech_nand3 i_57129(.A(n_1303), .B(n_1607), .C(n_1302), .Z(n_1304));
	notech_nand2 i_512(.A(n_1377), .B(cacheQ[119]), .Z(n_1305));
	notech_nand3 i_511(.A(n_59526), .B(axi_W[23]), .C(n_59508), .Z(n_1306)
		);
	notech_nand3 i_57126(.A(n_1306), .B(n_1611), .C(n_1305), .Z(n_1307));
	notech_nand2 i_516(.A(n_1377), .B(cacheQ[118]), .Z(n_1308));
	notech_nand3 i_515(.A(n_59526), .B(axi_W[22]), .C(n_59504), .Z(n_1309)
		);
	notech_nand3 i_57123(.A(n_1309), .B(n_1615), .C(n_1308), .Z(n_1310));
	notech_nand2 i_520(.A(n_1377), .B(cacheQ[117]), .Z(n_1311));
	notech_nand3 i_519(.A(n_59526), .B(axi_W[21]), .C(n_59504), .Z(n_1312)
		);
	notech_nand3 i_57120(.A(n_1312), .B(n_1619), .C(n_1311), .Z(n_1313));
	notech_nand2 i_524(.A(n_1377), .B(cacheQ[116]), .Z(n_1314));
	notech_nand3 i_523(.A(n_59526), .B(axi_W[20]), .C(n_59504), .Z(n_1315)
		);
	notech_nand3 i_57117(.A(n_1315), .B(n_1623), .C(n_1314), .Z(n_1316));
	notech_nand2 i_528(.A(n_1377), .B(cacheQ[115]), .Z(n_1317));
	notech_nand3 i_527(.A(n_59526), .B(axi_W[19]), .C(n_59504), .Z(n_1318)
		);
	notech_nand3 i_57114(.A(n_1318), .B(n_1627), .C(n_1317), .Z(n_1319));
	notech_nand2 i_532(.A(n_1377), .B(cacheQ[114]), .Z(n_1320));
	notech_nand3 i_531(.A(n_59526), .B(axi_W[18]), .C(n_59504), .Z(n_1321)
		);
	notech_nand3 i_57111(.A(n_1321), .B(n_1631), .C(n_1320), .Z(n_1322));
	notech_nand2 i_536(.A(n_1377), .B(cacheQ[113]), .Z(n_1323));
	notech_nand3 i_535(.A(n_59526), .B(axi_W[17]), .C(n_59504), .Z(n_1324)
		);
	notech_nand3 i_57108(.A(n_1324), .B(n_1635), .C(n_1323), .Z(n_1325));
	notech_nand2 i_540(.A(n_1377), .B(cacheQ[112]), .Z(n_1326));
	notech_nand3 i_539(.A(n_59526), .B(axi_W[16]), .C(n_59504), .Z(n_1327)
		);
	notech_nand3 i_57105(.A(n_1327), .B(n_1639), .C(n_1326), .Z(n_1328));
	notech_nand2 i_544(.A(n_59452), .B(cacheQ[111]), .Z(n_1329));
	notech_nand3 i_543(.A(n_59526), .B(axi_W[15]), .C(n_59504), .Z(n_1330)
		);
	notech_nand3 i_57102(.A(n_1330), .B(n_1643), .C(n_1329), .Z(n_1331));
	notech_nand2 i_548(.A(n_59452), .B(cacheQ[110]), .Z(n_1332));
	notech_nand3 i_547(.A(n_59526), .B(axi_W[14]), .C(n_59504), .Z(n_1333)
		);
	notech_nand3 i_57099(.A(n_1333), .B(n_1647), .C(n_1332), .Z(n_1334));
	notech_nand2 i_552(.A(n_59452), .B(cacheQ[109]), .Z(n_1335));
	notech_nand3 i_551(.A(n_59527), .B(axi_W[13]), .C(n_59504), .Z(n_1336)
		);
	notech_nand3 i_57096(.A(n_1336), .B(n_1651), .C(n_1335), .Z(n_1337));
	notech_nand2 i_556(.A(n_59452), .B(cacheQ[108]), .Z(n_1338));
	notech_nand3 i_555(.A(n_59527), .B(axi_W[12]), .C(n_59508), .Z(n_1339)
		);
	notech_nand3 i_57093(.A(n_1339), .B(n_1655), .C(n_1338), .Z(n_1340));
	notech_nand2 i_560(.A(n_59452), .B(cacheQ[107]), .Z(n_1341));
	notech_nand3 i_559(.A(n_59527), .B(axi_W[11]), .C(n_59510), .Z(n_1342)
		);
	notech_nand3 i_57090(.A(n_1342), .B(n_1659), .C(n_1341), .Z(n_1343));
	notech_nand2 i_564(.A(n_59452), .B(cacheQ[106]), .Z(n_1344));
	notech_nand3 i_563(.A(n_59527), .B(axi_W[10]), .C(n_59510), .Z(n_1345)
		);
	notech_nand3 i_57087(.A(n_1345), .B(n_1663), .C(n_1344), .Z(n_1346));
	notech_nand2 i_568(.A(n_59452), .B(cacheQ[105]), .Z(n_1347));
	notech_nand3 i_567(.A(n_59527), .B(axi_W[9]), .C(n_59510), .Z(n_1348));
	notech_nand3 i_57084(.A(n_1348), .B(n_1667), .C(n_1347), .Z(n_1349));
	notech_nand2 i_572(.A(n_59452), .B(cacheQ[104]), .Z(n_1350));
	notech_nand3 i_571(.A(n_59527), .B(axi_W[8]), .C(n_59510), .Z(n_1351));
	notech_nand3 i_57081(.A(n_1351), .B(n_1671), .C(n_1350), .Z(n_1352));
	notech_nand2 i_576(.A(n_59452), .B(cacheQ[103]), .Z(n_1353));
	notech_nand3 i_575(.A(n_59527), .B(axi_W[7]), .C(n_59510), .Z(n_1354));
	notech_nand3 i_57078(.A(n_1354), .B(n_1675), .C(n_1353), .Z(n_1355));
	notech_nand2 i_580(.A(n_59452), .B(cacheQ[102]), .Z(n_1356));
	notech_nand3 i_579(.A(n_59527), .B(axi_W[6]), .C(n_59510), .Z(n_1357));
	notech_nand3 i_57075(.A(n_1357), .B(n_1679), .C(n_1356), .Z(n_1358));
	notech_nand2 i_584(.A(n_59452), .B(cacheQ[101]), .Z(n_1359));
	notech_nand3 i_583(.A(n_59527), .B(axi_W[5]), .C(n_59510), .Z(n_1360));
	notech_nand3 i_57072(.A(n_1360), .B(n_1683), .C(n_1359), .Z(n_1361));
	notech_nand2 i_588(.A(n_59452), .B(cacheQ[100]), .Z(n_1362));
	notech_nand3 i_587(.A(n_59527), .B(axi_W[4]), .C(n_59510), .Z(n_1363));
	notech_nand3 i_57069(.A(n_1363), .B(n_1687), .C(n_1362), .Z(n_1364));
	notech_nand2 i_592(.A(n_59452), .B(cacheQ[99]), .Z(n_1365));
	notech_nand3 i_591(.A(n_59527), .B(axi_W[3]), .C(n_59510), .Z(n_1366));
	notech_nand3 i_57066(.A(n_1366), .B(n_1691), .C(n_1365), .Z(n_1367));
	notech_nand2 i_596(.A(n_59452), .B(cacheQ[98]), .Z(n_1368));
	notech_nand3 i_595(.A(n_59527), .B(axi_W[2]), .C(n_59510), .Z(n_1369));
	notech_nand3 i_57063(.A(n_1369), .B(n_1695), .C(n_1368), .Z(n_1370));
	notech_nand2 i_600(.A(n_59452), .B(cacheQ[97]), .Z(n_1371));
	notech_nand3 i_599(.A(n_59527), .B(axi_W[1]), .C(n_59508), .Z(n_1372));
	notech_nand3 i_57060(.A(n_1372), .B(n_1699), .C(n_1371), .Z(n_1373));
	notech_ao4 i_57713(.A(n_210855939), .B(n_2025), .C(n_2070), .D(n_7001), 
		.Z(n_1375));
	notech_nand2 i_606(.A(n_59452), .B(cacheQ[96]), .Z(n_1376));
	notech_nand2 i_19(.A(n_59491), .B(n_2073), .Z(n_1377));
	notech_nand3 i_605(.A(n_59527), .B(axi_W[0]), .C(n_59508), .Z(n_1378));
	notech_nand3 i_57057(.A(n_1378), .B(n_1706), .C(n_1376), .Z(n_1379));
	notech_nand2 i_610(.A(cacheQ[95]), .B(n_1476), .Z(n_1380));
	notech_nand3 i_609(.A(n_59527), .B(axi_W[31]), .C(n_59470), .Z(n_1381)
		);
	notech_nand3 i_57054(.A(n_1579), .B(n_1381), .C(n_1380), .Z(n_1382));
	notech_nand2 i_614(.A(n_1476), .B(cacheQ[94]), .Z(n_1383));
	notech_nand3 i_613(.A(n_59527), .B(axi_W[30]), .C(n_59473), .Z(n_1384)
		);
	notech_nand3 i_57051(.A(n_1583), .B(n_1384), .C(n_1383), .Z(n_1385));
	notech_nand2 i_618(.A(n_1476), .B(cacheQ[93]), .Z(n_1386));
	notech_nand3 i_617(.A(n_59527), .B(axi_W[29]), .C(n_59473), .Z(n_1387)
		);
	notech_nand3 i_57048(.A(n_1587), .B(n_1387), .C(n_1386), .Z(n_1388));
	notech_nand2 i_622(.A(n_1476), .B(cacheQ[92]), .Z(n_1389));
	notech_nand3 i_621(.A(n_59527), .B(axi_W[28]), .C(n_59470), .Z(n_1390)
		);
	notech_nand3 i_57045(.A(n_1591), .B(n_1390), .C(n_1389), .Z(n_1391));
	notech_nand2 i_626(.A(n_1476), .B(cacheQ[91]), .Z(n_1392));
	notech_nand3 i_625(.A(n_59526), .B(axi_W[27]), .C(n_59470), .Z(n_1393)
		);
	notech_nand3 i_57042(.A(n_1595), .B(n_1393), .C(n_1392), .Z(n_1394));
	notech_nand2 i_630(.A(n_1476), .B(cacheQ[90]), .Z(n_1395));
	notech_nand3 i_629(.A(n_59514), .B(axi_W[26]), .C(n_59470), .Z(n_1396)
		);
	notech_nand3 i_57039(.A(n_1599), .B(n_1396), .C(n_1395), .Z(n_1397));
	notech_nand2 i_634(.A(n_1476), .B(cacheQ[89]), .Z(n_1398));
	notech_nand3 i_633(.A(n_59514), .B(axi_W[25]), .C(n_59473), .Z(n_1399)
		);
	notech_nand3 i_57036(.A(n_1603), .B(n_1399), .C(n_1398), .Z(n_1400));
	notech_nand2 i_638(.A(n_1476), .B(cacheQ[88]), .Z(n_1401));
	notech_nand3 i_637(.A(n_59514), .B(axi_W[24]), .C(n_59473), .Z(n_1402)
		);
	notech_nand3 i_57033(.A(n_1607), .B(n_1402), .C(n_1401), .Z(n_1403));
	notech_nand2 i_642(.A(n_1476), .B(cacheQ[87]), .Z(n_1404));
	notech_nand3 i_641(.A(n_59514), .B(axi_W[23]), .C(n_59473), .Z(n_1405)
		);
	notech_nand3 i_57030(.A(n_1611), .B(n_1405), .C(n_1404), .Z(n_1406));
	notech_nand2 i_646(.A(n_1476), .B(cacheQ[86]), .Z(n_1407));
	notech_nand3 i_645(.A(n_59520), .B(axi_W[22]), .C(n_59473), .Z(n_1408)
		);
	notech_nand3 i_57027(.A(n_1615), .B(n_1408), .C(n_1407), .Z(n_1409));
	notech_nand2 i_650(.A(n_1476), .B(cacheQ[85]), .Z(n_1410));
	notech_nand3 i_649(.A(n_59520), .B(axi_W[21]), .C(n_59473), .Z(n_1411)
		);
	notech_nand3 i_57024(.A(n_1619), .B(n_1411), .C(n_1410), .Z(n_1412));
	notech_nand2 i_654(.A(n_1476), .B(cacheQ[84]), .Z(n_1413));
	notech_nand3 i_653(.A(n_59520), .B(axi_W[20]), .C(n_59473), .Z(n_1414)
		);
	notech_nand3 i_57021(.A(n_1623), .B(n_1414), .C(n_1413), .Z(n_1415));
	notech_nand2 i_658(.A(n_1476), .B(cacheQ[83]), .Z(n_1416));
	notech_nand3 i_657(.A(n_59520), .B(axi_W[19]), .C(n_59473), .Z(n_1417)
		);
	notech_nand3 i_57018(.A(n_1627), .B(n_1417), .C(n_1416), .Z(n_1418));
	notech_nand2 i_662(.A(n_1476), .B(cacheQ[82]), .Z(n_1419));
	notech_nand3 i_661(.A(n_59520), .B(axi_W[18]), .C(n_59470), .Z(n_1420)
		);
	notech_nand3 i_57015(.A(n_1631), .B(n_1420), .C(n_1419), .Z(n_1421));
	notech_nand2 i_666(.A(n_1476), .B(cacheQ[81]), .Z(n_1422));
	notech_nand3 i_665(.A(n_59514), .B(axi_W[17]), .C(n_59470), .Z(n_1423)
		);
	notech_nand3 i_57012(.A(n_1635), .B(n_1423), .C(n_1422), .Z(n_1424));
	notech_nand2 i_670(.A(n_1476), .B(cacheQ[80]), .Z(n_1425));
	notech_nand3 i_669(.A(n_59514), .B(axi_W[16]), .C(n_59470), .Z(n_1426)
		);
	notech_nand3 i_57009(.A(n_1639), .B(n_1426), .C(n_1425), .Z(n_1427));
	notech_nand2 i_674(.A(n_59430), .B(cacheQ[79]), .Z(n_1428));
	notech_nand3 i_673(.A(n_59514), .B(axi_W[15]), .C(n_59470), .Z(n_1429)
		);
	notech_nand3 i_57006(.A(n_1643), .B(n_1429), .C(n_1428), .Z(n_1430));
	notech_nand2 i_678(.A(n_59430), .B(cacheQ[78]), .Z(n_1431));
	notech_nand3 i_677(.A(n_59514), .B(axi_W[14]), .C(n_59470), .Z(n_1432)
		);
	notech_nand3 i_57003(.A(n_1647), .B(n_1432), .C(n_1431), .Z(n_1433));
	notech_nand2 i_682(.A(n_59430), .B(cacheQ[77]), .Z(n_1434));
	notech_nand3 i_681(.A(n_59514), .B(axi_W[13]), .C(n_59470), .Z(n_1435)
		);
	notech_nand3 i_57000(.A(n_1651), .B(n_1435), .C(n_1434), .Z(n_1436));
	notech_nand2 i_686(.A(n_59430), .B(cacheQ[76]), .Z(n_1437));
	notech_nand3 i_685(.A(n_59514), .B(axi_W[12]), .C(n_59470), .Z(n_1438)
		);
	notech_nand3 i_56997(.A(n_1655), .B(n_1438), .C(n_1437), .Z(n_1439));
	notech_nand2 i_690(.A(n_59430), .B(cacheQ[75]), .Z(n_1440));
	notech_nand3 i_689(.A(n_59514), .B(axi_W[11]), .C(n_59470), .Z(n_1441)
		);
	notech_nand3 i_56994(.A(n_1659), .B(n_1441), .C(n_1440), .Z(n_1442));
	notech_nand2 i_694(.A(n_59430), .B(cacheQ[74]), .Z(n_1443));
	notech_nand3 i_693(.A(n_59514), .B(axi_W[10]), .C(n_59470), .Z(n_1444)
		);
	notech_nand3 i_56991(.A(n_1663), .B(n_1444), .C(n_1443), .Z(n_1445));
	notech_nand2 i_698(.A(n_59430), .B(cacheQ[73]), .Z(n_1446));
	notech_nand3 i_697(.A(n_59514), .B(axi_W[9]), .C(n_59470), .Z(n_1447));
	notech_nand3 i_56988(.A(n_1667), .B(n_1447), .C(n_1446), .Z(n_1448));
	notech_nand2 i_702(.A(n_59430), .B(cacheQ[72]), .Z(n_1449));
	notech_nand3 i_701(.A(n_59520), .B(axi_W[8]), .C(n_59470), .Z(n_1450));
	notech_nand3 i_56985(.A(n_1671), .B(n_1450), .C(n_1449), .Z(n_1451));
	notech_nand2 i_706(.A(n_59430), .B(cacheQ[71]), .Z(n_1452));
	notech_nand3 i_705(.A(n_59520), .B(axi_W[7]), .C(n_59470), .Z(n_1453));
	notech_nand3 i_56982(.A(n_1675), .B(n_1453), .C(n_1452), .Z(n_1454));
	notech_nand2 i_710(.A(n_59430), .B(cacheQ[70]), .Z(n_1455));
	notech_nand3 i_709(.A(n_59520), .B(axi_W[6]), .C(n_59470), .Z(n_1456));
	notech_nand3 i_56979(.A(n_1679), .B(n_1456), .C(n_1455), .Z(n_1457));
	notech_nand2 i_714(.A(n_59430), .B(cacheQ[69]), .Z(n_1458));
	notech_nand3 i_713(.A(n_59520), .B(axi_W[5]), .C(n_59473), .Z(n_1459));
	notech_nand3 i_56976(.A(n_1683), .B(n_1459), .C(n_1458), .Z(n_1460));
	notech_nand2 i_718(.A(n_59430), .B(cacheQ[68]), .Z(n_1461));
	notech_nand3 i_717(.A(n_59520), .B(axi_W[4]), .C(n_59475), .Z(n_1462));
	notech_nand3 i_56973(.A(n_1687), .B(n_1462), .C(n_1461), .Z(n_1463));
	notech_nand2 i_722(.A(n_59430), .B(cacheQ[67]), .Z(n_1464));
	notech_nand3 i_721(.A(n_59526), .B(axi_W[3]), .C(n_59475), .Z(n_1465));
	notech_nand3 i_56970(.A(n_1691), .B(n_1465), .C(n_1464), .Z(n_1466));
	notech_nand2 i_726(.A(n_59430), .B(cacheQ[66]), .Z(n_1467));
	notech_nand3 i_725(.A(n_59526), .B(axi_W[2]), .C(n_59475), .Z(n_1468));
	notech_nand3 i_56967(.A(n_1695), .B(n_1468), .C(n_1467), .Z(n_1469));
	notech_nand2 i_730(.A(n_59430), .B(cacheQ[65]), .Z(n_1470));
	notech_nand3 i_729(.A(n_59520), .B(axi_W[1]), .C(n_59475), .Z(n_1471));
	notech_nand3 i_56964(.A(n_1699), .B(n_1471), .C(n_1470), .Z(n_1472));
	notech_ao4 i_57712(.A(n_210855939), .B(n_6663), .C(n_2070), .D(n_7001), 
		.Z(n_1474));
	notech_nand2 i_736(.A(n_59430), .B(cacheQ[64]), .Z(n_1475));
	notech_nand2 i_18(.A(n_59491), .B(n_2075), .Z(n_1476));
	notech_nand3 i_735(.A(n_59526), .B(axi_W[0]), .C(n_59475), .Z(n_1477));
	notech_nand3 i_56961(.A(n_1706), .B(n_1477), .C(n_1475), .Z(n_1478));
	notech_nand2 i_740(.A(cacheQ[63]), .B(n_1575), .Z(n_1479));
	notech_nao3 i_739(.A(axi_W[31]), .B(n_59508), .C(n_59491), .Z(n_1480));
	notech_nand3 i_56958(.A(n_1579), .B(n_1480), .C(n_1479), .Z(n_1481));
	notech_nand2 i_744(.A(n_1575), .B(cacheQ[62]), .Z(n_1482));
	notech_nao3 i_743(.A(axi_W[30]), .B(n_59508), .C(n_59491), .Z(n_1483));
	notech_nand3 i_56955(.A(n_1583), .B(n_1483), .C(n_1482), .Z(n_1484));
	notech_nand2 i_748(.A(n_1575), .B(cacheQ[61]), .Z(n_1485));
	notech_nao3 i_747(.A(axi_W[29]), .B(n_59508), .C(n_59491), .Z(n_1486));
	notech_nand3 i_56952(.A(n_1587), .B(n_1486), .C(n_1485), .Z(n_1487));
	notech_nand2 i_752(.A(n_1575), .B(cacheQ[60]), .Z(n_1488));
	notech_nao3 i_751(.A(axi_W[28]), .B(n_59510), .C(n_59491), .Z(n_1489));
	notech_nand3 i_56949(.A(n_1591), .B(n_1489), .C(n_1488), .Z(n_1490));
	notech_nand2 i_756(.A(n_1575), .B(cacheQ[59]), .Z(n_1491));
	notech_nao3 i_755(.A(axi_W[27]), .B(n_59510), .C(n_59492), .Z(n_1492));
	notech_nand3 i_56946(.A(n_1595), .B(n_1492), .C(n_1491), .Z(n_1493));
	notech_nand2 i_760(.A(n_1575), .B(cacheQ[58]), .Z(n_1494));
	notech_nao3 i_759(.A(axi_W[26]), .B(n_59510), .C(n_59491), .Z(n_1495));
	notech_nand3 i_56943(.A(n_1599), .B(n_1495), .C(n_1494), .Z(n_1496));
	notech_nand2 i_764(.A(n_1575), .B(cacheQ[57]), .Z(n_1497));
	notech_nao3 i_763(.A(axi_W[25]), .B(n_59510), .C(n_59491), .Z(n_1498));
	notech_nand3 i_56940(.A(n_1603), .B(n_1498), .C(n_1497), .Z(n_1499));
	notech_nand2 i_768(.A(n_1575), .B(cacheQ[56]), .Z(n_1500));
	notech_nao3 i_767(.A(axi_W[24]), .B(n_59510), .C(n_59491), .Z(n_1501));
	notech_nand3 i_56937(.A(n_1607), .B(n_1501), .C(n_1500), .Z(n_1502));
	notech_nand2 i_772(.A(n_1575), .B(cacheQ[55]), .Z(n_1503));
	notech_nao3 i_771(.A(axi_W[23]), .B(n_59510), .C(n_59491), .Z(n_1504));
	notech_nand3 i_56934(.A(n_1611), .B(n_1504), .C(n_1503), .Z(n_1505));
	notech_nand2 i_776(.A(n_1575), .B(cacheQ[54]), .Z(n_1506));
	notech_nao3 i_775(.A(axi_W[22]), .B(n_59503), .C(n_59491), .Z(n_1507));
	notech_nand3 i_56931(.A(n_1615), .B(n_1507), .C(n_1506), .Z(n_1508));
	notech_nand2 i_780(.A(n_1575), .B(cacheQ[53]), .Z(n_1509));
	notech_nao3 i_779(.A(axi_W[21]), .B(n_59503), .C(n_59491), .Z(n_1510));
	notech_nand3 i_56928(.A(n_1619), .B(n_1510), .C(n_1509), .Z(n_1511));
	notech_nand2 i_784(.A(n_1575), .B(cacheQ[52]), .Z(n_1512));
	notech_nao3 i_783(.A(axi_W[20]), .B(n_59510), .C(n_59491), .Z(n_1513));
	notech_nand3 i_56925(.A(n_1623), .B(n_1513), .C(n_1512), .Z(n_1514));
	notech_nand2 i_788(.A(n_1575), .B(cacheQ[51]), .Z(n_1515));
	notech_nao3 i_787(.A(axi_W[19]), .B(n_59510), .C(n_59491), .Z(n_1516));
	notech_nand3 i_56922(.A(n_1627), .B(n_1516), .C(n_1515), .Z(n_1517));
	notech_nand2 i_792(.A(n_1575), .B(cacheQ[50]), .Z(n_1518));
	notech_nao3 i_791(.A(axi_W[18]), .B(n_59508), .C(n_59491), .Z(n_1519));
	notech_nand3 i_56919(.A(n_1631), .B(n_1519), .C(n_1518), .Z(n_1520));
	notech_nand2 i_796(.A(n_1575), .B(cacheQ[49]), .Z(n_1521));
	notech_nao3 i_795(.A(axi_W[17]), .B(n_59510), .C(n_59491), .Z(n_1522));
	notech_nand3 i_56916(.A(n_1635), .B(n_1522), .C(n_1521), .Z(n_1523));
	notech_nand2 i_800(.A(n_1575), .B(cacheQ[48]), .Z(n_1524));
	notech_nao3 i_799(.A(axi_W[16]), .B(n_59510), .C(n_59491), .Z(n_1525));
	notech_nand3 i_56913(.A(n_1639), .B(n_1525), .C(n_1524), .Z(n_1526));
	notech_nand2 i_804(.A(n_59408), .B(cacheQ[47]), .Z(n_1527));
	notech_nao3 i_803(.A(axi_W[15]), .B(n_59503), .C(n_59492), .Z(n_1528));
	notech_nand3 i_56910(.A(n_1643), .B(n_1528), .C(n_1527), .Z(n_1529));
	notech_nand2 i_808(.A(n_59408), .B(cacheQ[46]), .Z(n_1530));
	notech_nao3 i_807(.A(axi_W[14]), .B(n_59498), .C(n_59492), .Z(n_1531));
	notech_nand3 i_56907(.A(n_1647), .B(n_1531), .C(n_1530), .Z(n_1532));
	notech_nand2 i_812(.A(n_59408), .B(cacheQ[45]), .Z(n_1533));
	notech_nao3 i_811(.A(axi_W[13]), .B(n_59498), .C(n_59492), .Z(n_1534));
	notech_nand3 i_56904(.A(n_1651), .B(n_1534), .C(n_1533), .Z(n_1535));
	notech_nand2 i_816(.A(n_59408), .B(cacheQ[44]), .Z(n_1536));
	notech_nao3 i_815(.A(axi_W[12]), .B(n_59498), .C(n_59492), .Z(n_1537));
	notech_nand3 i_56901(.A(n_1655), .B(n_1537), .C(n_1536), .Z(n_1538));
	notech_nand2 i_820(.A(n_59408), .B(cacheQ[43]), .Z(n_1539));
	notech_nao3 i_819(.A(axi_W[11]), .B(n_59498), .C(n_59492), .Z(n_1540));
	notech_nand3 i_56898(.A(n_1659), .B(n_1540), .C(n_1539), .Z(n_1541));
	notech_nand2 i_824(.A(n_59408), .B(cacheQ[42]), .Z(n_1542));
	notech_nao3 i_823(.A(axi_W[10]), .B(n_59498), .C(n_59492), .Z(n_1543));
	notech_nand3 i_56895(.A(n_1663), .B(n_1543), .C(n_1542), .Z(n_1544));
	notech_nand2 i_828(.A(n_59408), .B(cacheQ[41]), .Z(n_1545));
	notech_nao3 i_827(.A(axi_W[9]), .B(n_59503), .C(n_59492), .Z(n_1546));
	notech_nand3 i_56892(.A(n_1667), .B(n_1546), .C(n_1545), .Z(n_1547));
	notech_nand2 i_832(.A(n_59408), .B(cacheQ[40]), .Z(n_1548));
	notech_nao3 i_831(.A(axi_W[8]), .B(n_59503), .C(n_59492), .Z(n_1549));
	notech_nand3 i_56889(.A(n_1671), .B(n_1549), .C(n_1548), .Z(n_1550));
	notech_nand2 i_836(.A(n_59408), .B(cacheQ[39]), .Z(n_1551));
	notech_nao3 i_835(.A(axi_W[7]), .B(n_59498), .C(n_59492), .Z(n_1552));
	notech_nand3 i_56886(.A(n_1675), .B(n_1552), .C(n_1551), .Z(n_1553));
	notech_nand2 i_840(.A(n_59408), .B(cacheQ[38]), .Z(n_1554));
	notech_nao3 i_839(.A(axi_W[6]), .B(n_59503), .C(n_59492), .Z(n_1555));
	notech_nand3 i_56883(.A(n_1679), .B(n_1555), .C(n_1554), .Z(n_1556));
	notech_nand2 i_844(.A(n_59408), .B(cacheQ[37]), .Z(n_1557));
	notech_nao3 i_843(.A(axi_W[5]), .B(n_59508), .C(n_59492), .Z(n_1558));
	notech_nand3 i_56880(.A(n_1683), .B(n_1558), .C(n_1557), .Z(n_1559));
	notech_nand2 i_848(.A(n_59408), .B(cacheQ[36]), .Z(n_1560));
	notech_nao3 i_847(.A(axi_W[4]), .B(n_59504), .C(n_59492), .Z(n_1561));
	notech_nand3 i_56877(.A(n_1687), .B(n_1561), .C(n_1560), .Z(n_1562));
	notech_nand2 i_852(.A(n_59408), .B(cacheQ[35]), .Z(n_1563));
	notech_nao3 i_851(.A(axi_W[3]), .B(n_59504), .C(n_59492), .Z(n_1564));
	notech_nand3 i_56874(.A(n_1691), .B(n_1564), .C(n_1563), .Z(n_1565));
	notech_nand2 i_856(.A(n_59408), .B(cacheQ[34]), .Z(n_1566));
	notech_nao3 i_855(.A(axi_W[2]), .B(n_59504), .C(n_59492), .Z(n_1567));
	notech_nand3 i_56871(.A(n_1695), .B(n_1567), .C(n_1566), .Z(n_1568));
	notech_nand2 i_860(.A(n_59408), .B(cacheQ[33]), .Z(n_1569));
	notech_nao3 i_859(.A(axi_W[1]), .B(n_59504), .C(n_59492), .Z(n_1570));
	notech_nand3 i_56868(.A(n_1699), .B(n_1570), .C(n_1569), .Z(n_1571));
	notech_ao4 i_57711(.A(n_210855939), .B(n_6662), .C(n_2070), .D(n_7001), 
		.Z(n_1573));
	notech_nand2 i_866(.A(n_59408), .B(cacheQ[32]), .Z(n_1574));
	notech_or2 i_17(.A(n_59520), .B(n_214255973), .Z(n_1575));
	notech_nao3 i_865(.A(axi_W[0]), .B(n_59504), .C(n_59492), .Z(n_1576));
	notech_nand3 i_56865(.A(n_1706), .B(n_1576), .C(n_1574), .Z(n_1577));
	notech_nand2 i_870(.A(cacheQ[31]), .B(n_1705), .Z(n_1578));
	notech_nand2 i_104(.A(axi_R[31]), .B(n_2023), .Z(n_1579));
	notech_nao3 i_869(.A(axi_W[31]), .B(n_59475), .C(n_59492), .Z(n_1580));
	notech_nand3 i_56862(.A(n_1579), .B(n_1580), .C(n_1578), .Z(n_1581));
	notech_nand2 i_874(.A(n_1705), .B(cacheQ[30]), .Z(n_1582));
	notech_nand2 i_102(.A(axi_R[30]), .B(n_2023), .Z(n_1583));
	notech_nao3 i_873(.A(axi_W[30]), .B(n_59475), .C(n_59492), .Z(n_1584));
	notech_nand3 i_56859(.A(n_1583), .B(n_1584), .C(n_1582), .Z(n_1585));
	notech_nand2 i_878(.A(n_1705), .B(cacheQ[29]), .Z(n_1586));
	notech_nand2 i_101(.A(axi_R[29]), .B(n_2023), .Z(n_1587));
	notech_nao3 i_877(.A(axi_W[29]), .B(n_59475), .C(n_59492), .Z(n_1588));
	notech_nand3 i_56856(.A(n_1587), .B(n_1588), .C(n_1586), .Z(n_1589));
	notech_nand2 i_882(.A(n_1705), .B(cacheQ[28]), .Z(n_1590));
	notech_nand2 i_106(.A(axi_R[28]), .B(n_2023), .Z(n_1591));
	notech_nao3 i_881(.A(axi_W[28]), .B(n_59475), .C(n_59479), .Z(n_1592));
	notech_nand3 i_56853(.A(n_1591), .B(n_1592), .C(n_1590), .Z(n_1593));
	notech_nand2 i_886(.A(n_1705), .B(cacheQ[27]), .Z(n_1594));
	notech_nand2 i_99(.A(axi_R[27]), .B(n_2023), .Z(n_1595));
	notech_nao3 i_885(.A(axi_W[27]), .B(n_59475), .C(n_59479), .Z(n_1596));
	notech_nand3 i_56850(.A(n_1595), .B(n_1596), .C(n_1594), .Z(n_1597));
	notech_nand2 i_890(.A(n_1705), .B(cacheQ[26]), .Z(n_1598));
	notech_nand2 i_97(.A(axi_R[26]), .B(n_2023), .Z(n_1599));
	notech_nao3 i_889(.A(axi_W[26]), .B(n_59475), .C(n_59479), .Z(n_1600));
	notech_nand3 i_56847(.A(n_1599), .B(n_1600), .C(n_1598), .Z(n_1601));
	notech_nand2 i_901(.A(n_1705), .B(cacheQ[25]), .Z(n_1602));
	notech_nand2 i_76(.A(axi_R[25]), .B(n_2023), .Z(n_1603));
	notech_nao3 i_897(.A(axi_W[25]), .B(n_59475), .C(n_59479), .Z(n_1604));
	notech_nand3 i_56844(.A(n_1603), .B(n_1604), .C(n_1602), .Z(n_1605));
	notech_nand2 i_905(.A(n_1705), .B(cacheQ[24]), .Z(n_1606));
	notech_nand2 i_108(.A(axi_R[24]), .B(n_2023), .Z(n_1607));
	notech_nao3 i_904(.A(axi_W[24]), .B(n_59475), .C(n_59479), .Z(n_1608));
	notech_nand3 i_56841(.A(n_1607), .B(n_1608), .C(n_1606), .Z(n_1609));
	notech_nand2 i_909(.A(n_1705), .B(cacheQ[23]), .Z(n_1610));
	notech_nand2 i_96(.A(axi_R[23]), .B(n_2023), .Z(n_1611));
	notech_nao3 i_908(.A(axi_W[23]), .B(n_59473), .C(n_59485), .Z(n_1612));
	notech_nand3 i_56838(.A(n_1611), .B(n_1612), .C(n_1610), .Z(n_1613));
	notech_nand2 i_913(.A(n_1705), .B(cacheQ[22]), .Z(n_1614));
	notech_nand2 i_95(.A(axi_R[22]), .B(n_2023), .Z(n_1615));
	notech_nao3 i_912(.A(axi_W[22]), .B(n_59473), .C(n_59485), .Z(n_1616));
	notech_nand3 i_56835(.A(n_1615), .B(n_1616), .C(n_1614), .Z(n_1617));
	notech_nand2 i_917(.A(n_1705), .B(cacheQ[21]), .Z(n_1618));
	notech_nand2 i_94(.A(axi_R[21]), .B(n_2023), .Z(n_1619));
	notech_nao3 i_916(.A(axi_W[21]), .B(n_59473), .C(n_59485), .Z(n_1620));
	notech_nand3 i_56832(.A(n_1619), .B(n_1620), .C(n_1618), .Z(n_1621));
	notech_nand2 i_924(.A(n_1705), .B(cacheQ[20]), .Z(n_1622));
	notech_nand2 i_86(.A(axi_R[20]), .B(n_2023), .Z(n_1623));
	notech_nao3 i_923(.A(axi_W[20]), .B(n_59473), .C(n_59485), .Z(n_1624));
	notech_nand3 i_56829(.A(n_1623), .B(n_1624), .C(n_1622), .Z(n_1625));
	notech_nand2 i_928(.A(n_1705), .B(cacheQ[19]), .Z(n_1626));
	notech_nand2 i_88(.A(axi_R[19]), .B(n_2023), .Z(n_1627));
	notech_nao3 i_927(.A(axi_W[19]), .B(n_59473), .C(n_59479), .Z(n_1628));
	notech_nand3 i_56826(.A(n_1627), .B(n_1628), .C(n_1626), .Z(n_1629));
	notech_nand2 i_932(.A(n_1705), .B(cacheQ[18]), .Z(n_1630));
	notech_nand2 i_89(.A(axi_R[18]), .B(n_2023), .Z(n_1631));
	notech_nao3 i_931(.A(axi_W[18]), .B(n_59473), .C(n_59479), .Z(n_1632));
	notech_nand3 i_56823(.A(n_1631), .B(n_1632), .C(n_1630), .Z(n_1633));
	notech_nand2 i_936(.A(n_1705), .B(cacheQ[17]), .Z(n_1634));
	notech_nand2 i_90(.A(axi_R[17]), .B(n_2023), .Z(n_1635));
	notech_nao3 i_935(.A(axi_W[17]), .B(n_59473), .C(n_59479), .Z(n_1636));
	notech_nand3 i_56820(.A(n_1635), .B(n_1636), .C(n_1634), .Z(n_1637));
	notech_nand2 i_940(.A(n_1705), .B(cacheQ[16]), .Z(n_1638));
	notech_nand2 i_91(.A(axi_R[16]), .B(n_2023), .Z(n_1639));
	notech_nao3 i_939(.A(axi_W[16]), .B(n_59475), .C(n_59479), .Z(n_1640));
	notech_nand3 i_56817(.A(n_1639), .B(n_1640), .C(n_1638), .Z(n_1641));
	notech_nand2 i_944(.A(n_59386), .B(cacheQ[15]), .Z(n_1642));
	notech_nand2 i_92(.A(axi_R[15]), .B(n_2023), .Z(n_1643));
	notech_nao3 i_943(.A(axi_W[15]), .B(n_59475), .C(n_59479), .Z(n_1644));
	notech_nand3 i_56814(.A(n_1643), .B(n_1644), .C(n_1642), .Z(n_1645));
	notech_nand2 i_948(.A(n_59386), .B(cacheQ[14]), .Z(n_1646));
	notech_nand2 i_93(.A(axi_R[14]), .B(n_2023), .Z(n_1647));
	notech_nao3 i_947(.A(axi_W[14]), .B(n_59475), .C(n_59479), .Z(n_1648));
	notech_nand3 i_56811(.A(n_1647), .B(n_1648), .C(n_1646), .Z(n_1649));
	notech_nand2 i_952(.A(n_59386), .B(cacheQ[13]), .Z(n_1650));
	notech_nand2 i_87(.A(axi_R[13]), .B(n_60835), .Z(n_1651));
	notech_nao3 i_951(.A(axi_W[13]), .B(n_59473), .C(n_59479), .Z(n_1652));
	notech_nand3 i_56808(.A(n_1651), .B(n_1652), .C(n_1650), .Z(n_1653));
	notech_nand2 i_956(.A(n_59386), .B(cacheQ[12]), .Z(n_1654));
	notech_nand2 i_103(.A(axi_R[12]), .B(n_60835), .Z(n_1655));
	notech_nao3 i_955(.A(axi_W[12]), .B(n_59475), .C(n_59479), .Z(n_1656));
	notech_nand3 i_56805(.A(n_1655), .B(n_1656), .C(n_1654), .Z(n_1657));
	notech_nand2 i_960(.A(n_59386), .B(cacheQ[11]), .Z(n_1658));
	notech_nand2 i_85(.A(axi_R[11]), .B(n_60835), .Z(n_1659));
	notech_nao3 i_959(.A(axi_W[11]), .B(n_59475), .C(n_59479), .Z(n_1660));
	notech_nand3 i_56802(.A(n_1659), .B(n_1660), .C(n_1658), .Z(n_1661));
	notech_nand2 i_964(.A(n_59386), .B(cacheQ[10]), .Z(n_1662));
	notech_nand2 i_84(.A(axi_R[10]), .B(n_60835), .Z(n_1663));
	notech_nao3 i_963(.A(axi_W[10]), .B(n_59470), .C(n_59485), .Z(n_1664));
	notech_nand3 i_56799(.A(n_1663), .B(n_1664), .C(n_1662), .Z(n_1665));
	notech_nand2 i_968(.A(n_59386), .B(cacheQ[9]), .Z(n_1666));
	notech_nand2 i_83(.A(axi_R[9]), .B(n_60835), .Z(n_1667));
	notech_nao3 i_967(.A(axi_W[9]), .B(n_59463), .C(n_59485), .Z(n_1668));
	notech_nand3 i_56796(.A(n_1667), .B(n_1668), .C(n_1666), .Z(n_1669));
	notech_nand2 i_972(.A(n_59386), .B(cacheQ[8]), .Z(n_1670));
	notech_nand2 i_82(.A(axi_R[8]), .B(n_60835), .Z(n_1671));
	notech_nao3 i_971(.A(axi_W[8]), .B(n_59465), .C(n_59485), .Z(n_1672));
	notech_nand3 i_56793(.A(n_1671), .B(n_1672), .C(n_1670), .Z(n_1673));
	notech_nand2 i_976(.A(n_59386), .B(cacheQ[7]), .Z(n_1674));
	notech_nand2 i_81(.A(axi_R[7]), .B(n_60835), .Z(n_1675));
	notech_nao3 i_975(.A(axi_W[7]), .B(n_59465), .C(n_59485), .Z(n_1676));
	notech_nand3 i_56790(.A(n_1675), .B(n_1676), .C(n_1674), .Z(n_1677));
	notech_nand2 i_980(.A(n_59386), .B(cacheQ[6]), .Z(n_1678));
	notech_nand2 i_80(.A(axi_R[6]), .B(n_60835), .Z(n_1679));
	notech_nao3 i_979(.A(axi_W[6]), .B(n_59463), .C(n_59485), .Z(n_1680));
	notech_nand3 i_56787(.A(n_1679), .B(n_1680), .C(n_1678), .Z(n_1681));
	notech_nand2 i_984(.A(n_59386), .B(cacheQ[5]), .Z(n_1682));
	notech_nand2 i_79(.A(axi_R[5]), .B(n_60835), .Z(n_1683));
	notech_nao3 i_983(.A(axi_W[5]), .B(n_59463), .C(n_59485), .Z(n_1684));
	notech_nand3 i_56784(.A(n_1683), .B(n_1684), .C(n_1682), .Z(n_1685));
	notech_nand2 i_988(.A(n_59386), .B(cacheQ[4]), .Z(n_1686));
	notech_nand2 i_107(.A(axi_R[4]), .B(n_60835), .Z(n_1687));
	notech_nao3 i_987(.A(axi_W[4]), .B(n_59463), .C(n_59491), .Z(n_1688));
	notech_nand3 i_56781(.A(n_1687), .B(n_1688), .C(n_1686), .Z(n_1689));
	notech_nand2 i_992(.A(n_59386), .B(cacheQ[3]), .Z(n_1690));
	notech_nand2 i_100(.A(axi_R[3]), .B(n_60835), .Z(n_1691));
	notech_nao3 i_991(.A(axi_W[3]), .B(n_59465), .C(n_59491), .Z(n_1692));
	notech_nand3 i_56778(.A(n_1691), .B(n_1692), .C(n_1690), .Z(n_1693));
	notech_nand2 i_996(.A(n_59386), .B(cacheQ[2]), .Z(n_1694));
	notech_nand2 i_77(.A(axi_R[2]), .B(n_60835), .Z(n_1695));
	notech_nao3 i_995(.A(axi_W[2]), .B(n_59465), .C(n_59485), .Z(n_1696));
	notech_nand3 i_56775(.A(n_1695), .B(n_1696), .C(n_1694), .Z(n_1697));
	notech_nand2 i_1000(.A(n_59386), .B(cacheQ[1]), .Z(n_1698));
	notech_nand2 i_74(.A(axi_R[1]), .B(n_60835), .Z(n_1699));
	notech_nao3 i_999(.A(axi_W[1]), .B(n_59465), .C(n_59491), .Z(n_1700));
	notech_nand3 i_56772(.A(n_1699), .B(n_1700), .C(n_1698), .Z(n_1701));
	notech_ao4 i_57710(.A(n_210855939), .B(n_2036), .C(n_2070), .D(n_7001), 
		.Z(n_1703));
	notech_nand2 i_1006(.A(n_59386), .B(cacheQ[0]), .Z(n_1704));
	notech_or2 i_16(.A(n_59520), .B(n_214355974), .Z(n_1705));
	notech_nand2 i_98(.A(axi_R[0]), .B(n_60835), .Z(n_1706));
	notech_nao3 i_1005(.A(axi_W[0]), .B(n_59465), .C(n_59485), .Z(n_1707));
	notech_nand3 i_56769(.A(n_1706), .B(n_1707), .C(n_1704), .Z(n_1708));
	notech_ao4 i_56182(.A(n_6763), .B(n_6998), .C(n_2002), .D(n_2007), .Z(n_1710
		));
	notech_nand2 i_1011(.A(n_2033), .B(n_21501), .Z(n_1711));
	notech_nand3 i_1014(.A(n_59520), .B(axi_WSTRB[3]), .C(n_59504), .Z(n_1712
		));
	notech_nand3 i_57246(.A(n_61518), .B(n_220956040), .C(n_1712), .Z(n_1713
		));
	notech_nand3 i_1016(.A(n_59520), .B(axi_WSTRB[2]), .C(n_59504), .Z(n_1714
		));
	notech_nand3 i_57244(.A(n_61518), .B(n_220956040), .C(n_1714), .Z(n_1715
		));
	notech_nand3 i_1018(.A(n_59520), .B(axi_WSTRB[1]), .C(n_59504), .Z(n_1716
		));
	notech_nand3 i_57242(.A(n_61518), .B(n_220956040), .C(n_1716), .Z(n_1717
		));
	notech_and4 i_1020(.A(A4[1]), .B(n_59504), .C(axi_WSTRB[0]), .D(n_2069),
		 .Z(n_1718));
	notech_nao3 i_57240(.A(n_61518), .B(n_220956040), .C(n_1718), .Z(n_1719)
		);
	notech_nand3 i_1022(.A(n_59520), .B(axi_WSTRB[3]), .C(n_59465), .Z(n_1720
		));
	notech_nand3 i_57238(.A(n_61518), .B(n_220956040), .C(n_1720), .Z(n_1721
		));
	notech_nand3 i_1024(.A(n_59520), .B(axi_WSTRB[2]), .C(n_59465), .Z(n_1722
		));
	notech_nand3 i_57236(.A(n_61518), .B(n_220956040), .C(n_1722), .Z(n_1723
		));
	notech_nand3 i_1026(.A(n_59520), .B(axi_WSTRB[1]), .C(n_59465), .Z(n_1724
		));
	notech_nand3 i_57234(.A(n_61518), .B(n_220956040), .C(n_1724), .Z(n_1725
		));
	notech_nand3 i_1028(.A(axi_WSTRB[0]), .B(n_59463), .C(n_59520), .Z(n_1726
		));
	notech_nand3 i_57232(.A(n_61518), .B(n_220956040), .C(n_1726), .Z(n_1727
		));
	notech_nao3 i_1030(.A(axi_WSTRB[3]), .B(n_59503), .C(n_59485), .Z(n_1728
		));
	notech_nand3 i_57230(.A(n_61518), .B(n_220956040), .C(n_1728), .Z(n_1729
		));
	notech_nao3 i_1032(.A(axi_WSTRB[2]), .B(n_59508), .C(n_59485), .Z(n_1730
		));
	notech_nand3 i_57228(.A(n_61523), .B(n_220956040), .C(n_1730), .Z(n_1731
		));
	notech_nao3 i_1034(.A(axi_WSTRB[1]), .B(n_59508), .C(n_59485), .Z(n_1732
		));
	notech_nand3 i_57226(.A(n_61523), .B(n_220956040), .C(n_1732), .Z(n_1733
		));
	notech_nao3 i_1036(.A(axi_WSTRB[0]), .B(n_59508), .C(n_59485), .Z(n_1734
		));
	notech_nand3 i_57224(.A(n_61523), .B(n_220956040), .C(n_1734), .Z(n_1735
		));
	notech_nao3 i_1038(.A(axi_WSTRB[3]), .B(n_59463), .C(n_59485), .Z(n_1736
		));
	notech_nand3 i_57222(.A(n_61523), .B(n_220956040), .C(n_1736), .Z(n_1737
		));
	notech_nao3 i_1040(.A(axi_WSTRB[2]), .B(n_59463), .C(n_59485), .Z(n_1738
		));
	notech_nand3 i_57220(.A(n_61523), .B(n_220956040), .C(n_1738), .Z(n_1739
		));
	notech_nao3 i_1042(.A(axi_WSTRB[1]), .B(n_59463), .C(n_59485), .Z(n_1740
		));
	notech_nand3 i_57218(.A(n_61523), .B(n_220956040), .C(n_1740), .Z(n_1741
		));
	notech_ao3 i_123(.A(fsm[4]), .B(fsm[2]), .C(n_1998), .Z(n_1742));
	notech_nand2 i_1044(.A(n_2049), .B(n_2050), .Z(n_1743));
	notech_ao3 i_58742(.A(n_2070), .B(n_1743), .C(n_1742), .Z(n_1744));
	notech_nao3 i_1047(.A(axi_WSTRB[0]), .B(n_59463), .C(n_59485), .Z(n_1745
		));
	notech_nand3 i_57216(.A(n_61523), .B(n_220956040), .C(n_1745), .Z(n_1746
		));
	notech_nand3 i_1050(.A(axi_RVALID), .B(axi_RLAST), .C(n_60835), .Z(n_1747
		));
	notech_and4 i_1051(.A(axi_AWREADY), .B(axi_AWVALID), .C(n_2037), .D(n_25082
		), .Z(n_1748));
	notech_ao3 i_57875(.A(n_61496), .B(n_1747), .C(n_221656047), .Z(n_1749)
		);
	notech_and2 i_1061(.A(n_2041), .B(n_2033), .Z(n_1750));
	notech_or4 i_57251(.A(n_1221), .B(n_974), .C(n_1750), .D(n_6664), .Z(n_1751
		));
	notech_nand2 i_1066(.A(axi_ARREADY), .B(n_6655), .Z(n_1754));
	notech_and4 i_59064(.A(n_2064), .B(n_61496), .C(n_973), .D(n_1754), .Z(n_1755
		));
	notech_nand2 i_57256(.A(n_60864), .B(n_221956050), .Z(n_1756));
	notech_nand2 i_1072(.A(axi_ARREADY), .B(n_1758), .Z(n_1757));
	notech_nand3 i_128(.A(n_2045), .B(n_6705), .C(n_60826), .Z(n_1758));
	notech_and4 i_59030(.A(n_60864), .B(n_1743), .C(n_2022), .D(n_1757), .Z(n_1759
		));
	notech_nand2 i_56192(.A(n_60864), .B(n_2019), .Z(n_1760));
	notech_ao4 i_69(.A(n_222656057), .B(n_222556056), .C(n_222456055), .D(n_6773
		), .Z(n_1763));
	notech_ao4 i_57653(.A(n_223056061), .B(n_223356064), .C(n_222756058), .D
		(n_6770), .Z(n_1765));
	notech_ao4 i_57895(.A(n_6659), .B(n_6658), .C(n_222756058), .D(n_6770), 
		.Z(n_1766));
	notech_ao4 i_58560(.A(readio_ack), .B(n_7000), .C(n_222656057), .D(n_222556056
		), .Z(n_1769));
	notech_ao4 i_59015(.A(n_223056061), .B(n_223156062), .C(n_6773), .D(n_222456055
		), .Z(n_1770));
	notech_mux2 i_1(.S(n_2033), .A(Daddr[4]), .B(axi_AW[4]), .Z(cacheA[0])
		);
	notech_mux2 i_211493(.S(n_2033), .A(Daddr[5]), .B(axi_AW[5]), .Z(cacheA[
		1]));
	notech_mux2 i_3(.S(n_2033), .A(Daddr[6]), .B(axi_AW[6]), .Z(cacheA[2])
		);
	notech_mux2 i_4(.S(n_2033), .A(Daddr[7]), .B(axi_AW[7]), .Z(cacheA[3])
		);
	notech_mux2 i_5(.S(n_2033), .A(Daddr[8]), .B(axi_AW[8]), .Z(cacheA[4])
		);
	notech_mux2 i_6(.S(n_2033), .A(Daddr[9]), .B(axi_AW[9]), .Z(cacheA[5])
		);
	notech_mux2 i_7(.S(n_2033), .A(Daddr[10]), .B(axi_AW[10]), .Z(cacheA[6])
		);
	notech_mux2 i_8(.S(n_60873), .A(Daddr[11]), .B(axi_AW[11]), .Z(cacheA[7]
		));
	notech_mux2 i_9(.S(n_60873), .A(Daddr[12]), .B(axi_AW[12]), .Z(cacheA[8]
		));
	notech_mux2 i_10(.S(n_60873), .A(Daddr[13]), .B(axi_AW[13]), .Z(cacheA[9
		]));
	notech_and4 i_1161(.A(n_59537), .B(n_61512), .C(cacheQ[64]), .D(n_59463)
		, .Z(n_1805));
	notech_nao3 i_122028(.A(n_2245), .B(n_2240), .C(n_1805), .Z(read_data[0]
		));
	notech_reg code_wack_reg(.CP(n_61979), .D(n_3180), .CD(n_61429), .Q(code_wack
		));
	notech_mux2 i_2330(.S(n_975), .A(n_25082), .B(code_wack), .Z(n_3180));
	notech_and4 i_1170(.A(A4[1]), .B(n_61512), .C(cacheQ[65]), .D(n_59463), 
		.Z(n_1811));
	notech_reg code_ack_slow_reg(.CP(n_61979), .D(n_3186), .CD(n_61429), .Q(code_ack
		));
	notech_mux2 i_2338(.S(n_977), .A(n_22749), .B(code_ack), .Z(n_3186));
	notech_nao3 i_222029(.A(n_2248), .B(n_2247), .C(n_1811), .Z(read_data[1]
		));
	notech_reg axi_AR_reg_0(.CP(n_61979), .D(n_3195), .CD(n_61429), .Q(axi_AR
		[0]));
	notech_and4 i_2348(.A(n_1066), .B(n_973), .C(axi_AR[0]), .D(n_61496), .Z
		(n_3195));
	notech_reg axi_AR_reg_1(.CP(n_61979), .D(n_3201), .CD(n_61429), .Q(axi_AR
		[1]));
	notech_and4 i_2356(.A(n_61496), .B(n_1066), .C(n_973), .D(axi_AR[1]), .Z
		(n_3201));
	notech_reg axi_AR_reg_2(.CP(n_61979), .D(n_3204), .CD(n_61429), .Q(axi_AR
		[2]));
	notech_mux2 i_2362(.S(n_1067), .A(n_6698), .B(axi_AR[2]), .Z(n_3204));
	notech_reg axi_AR_reg_3(.CP(n_61979), .D(n_3210), .CD(n_61429), .Q(axi_AR
		[3]));
	notech_mux2 i_2370(.S(n_1067), .A(n_6697), .B(axi_AR[3]), .Z(n_3210));
	notech_reg axi_AR_reg_4(.CP(n_61979), .D(n_3216), .CD(n_61429), .Q(axi_AR
		[4]));
	notech_mux2 i_2378(.S(n_1067), .A(n_6696), .B(axi_AR[4]), .Z(n_3216));
	notech_and4 i_1179(.A(A4[1]), .B(n_61512), .C(cacheQ[66]), .D(n_59463), 
		.Z(n_1817));
	notech_reg axi_AR_reg_5(.CP(n_61979), .D(n_3222), .CD(n_61429), .Q(axi_AR
		[5]));
	notech_mux2 i_2386(.S(n_1067), .A(n_6695), .B(axi_AR[5]), .Z(n_3222));
	notech_nao3 i_322030(.A(n_2251), .B(n_2250), .C(n_1817), .Z(read_data[2]
		));
	notech_reg axi_AR_reg_6(.CP(n_61979), .D(n_3228), .CD(n_61427), .Q(axi_AR
		[6]));
	notech_mux2 i_2394(.S(n_1067), .A(n_6694), .B(axi_AR[6]), .Z(n_3228));
	notech_reg axi_AR_reg_7(.CP(n_61979), .D(n_3234), .CD(n_61427), .Q(axi_AR
		[7]));
	notech_mux2 i_2402(.S(n_1067), .A(n_6693), .B(axi_AR[7]), .Z(n_3234));
	notech_reg axi_AR_reg_8(.CP(n_61979), .D(n_3240), .CD(n_61427), .Q(axi_AR
		[8]));
	notech_mux2 i_2410(.S(n_1067), .A(n_6692), .B(axi_AR[8]), .Z(n_3240));
	notech_reg axi_AR_reg_9(.CP(n_61979), .D(n_3246), .CD(n_61427), .Q(axi_AR
		[9]));
	notech_mux2 i_2418(.S(n_1067), .A(n_6691), .B(axi_AR[9]), .Z(n_3246));
	notech_reg axi_AR_reg_10(.CP(n_61979), .D(n_3252), .CD(n_61427), .Q(axi_AR
		[10]));
	notech_mux2 i_2426(.S(n_1067), .A(n_6690), .B(axi_AR[10]), .Z(n_3252));
	notech_and4 i_1188(.A(A4[1]), .B(n_61512), .C(cacheQ[67]), .D(n_59463), 
		.Z(n_1823));
	notech_reg axi_AR_reg_11(.CP(n_61979), .D(n_3258), .CD(n_61427), .Q(axi_AR
		[11]));
	notech_mux2 i_2434(.S(n_1067), .A(n_6689), .B(axi_AR[11]), .Z(n_3258));
	notech_nao3 i_422031(.A(n_2254), .B(n_2253), .C(n_1823), .Z(read_data[3]
		));
	notech_reg axi_AR_reg_12(.CP(n_61979), .D(n_3264), .CD(n_61427), .Q(axi_AR
		[12]));
	notech_mux2 i_2442(.S(n_1067), .A(n_6688), .B(axi_AR[12]), .Z(n_3264));
	notech_reg axi_AR_reg_13(.CP(n_61979), .D(n_3270), .CD(n_61427), .Q(axi_AR
		[13]));
	notech_mux2 i_2450(.S(n_1067), .A(n_6687), .B(axi_AR[13]), .Z(n_3270));
	notech_reg axi_AR_reg_14(.CP(n_61979), .D(n_3276), .CD(n_61429), .Q(axi_AR
		[14]));
	notech_mux2 i_2458(.S(n_1067), .A(n_6686), .B(axi_AR[14]), .Z(n_3276));
	notech_reg axi_AR_reg_15(.CP(n_61979), .D(n_3282), .CD(n_61430), .Q(axi_AR
		[15]));
	notech_mux2 i_2466(.S(n_1067), .A(n_6685), .B(axi_AR[15]), .Z(n_3282));
	notech_reg axi_AR_reg_16(.CP(n_61979), .D(n_3288), .CD(n_61430), .Q(axi_AR
		[16]));
	notech_mux2 i_2474(.S(n_1067), .A(n_6684), .B(axi_AR[16]), .Z(n_3288));
	notech_and4 i_1197(.A(n_59537), .B(n_61512), .C(cacheQ[68]), .D(n_59463)
		, .Z(n_1829));
	notech_reg axi_AR_reg_17(.CP(n_61995), .D(n_3294), .CD(n_61430), .Q(axi_AR
		[17]));
	notech_mux2 i_2482(.S(n_1067), .A(n_6683), .B(axi_AR[17]), .Z(n_3294));
	notech_nao3 i_522032(.A(n_2257), .B(n_2256), .C(n_1829), .Z(read_data[4]
		));
	notech_reg axi_AR_reg_18(.CP(n_61995), .D(n_3300), .CD(n_61430), .Q(axi_AR
		[18]));
	notech_mux2 i_2490(.S(n_60853), .A(n_6682), .B(axi_AR[18]), .Z(n_3300)
		);
	notech_reg axi_AR_reg_19(.CP(n_61995), .D(n_3306), .CD(n_61430), .Q(axi_AR
		[19]));
	notech_mux2 i_2498(.S(n_60853), .A(n_6681), .B(axi_AR[19]), .Z(n_3306)
		);
	notech_reg axi_AR_reg_20(.CP(n_61995), .D(n_3312), .CD(n_61430), .Q(axi_AR
		[20]));
	notech_mux2 i_2506(.S(n_60853), .A(n_6680), .B(axi_AR[20]), .Z(n_3312)
		);
	notech_reg axi_AR_reg_21(.CP(n_61995), .D(n_3318), .CD(n_61430), .Q(axi_AR
		[21]));
	notech_mux2 i_2514(.S(n_60853), .A(n_6679), .B(axi_AR[21]), .Z(n_3318)
		);
	notech_reg axi_AR_reg_22(.CP(n_61995), .D(n_3324), .CD(n_61430), .Q(axi_AR
		[22]));
	notech_mux2 i_2522(.S(n_60853), .A(n_6678), .B(axi_AR[22]), .Z(n_3324)
		);
	notech_and4 i_1206(.A(n_59537), .B(n_61512), .C(cacheQ[69]), .D(n_59463)
		, .Z(n_1835));
	notech_reg axi_AR_reg_23(.CP(n_61995), .D(n_3330), .CD(n_61429), .Q(axi_AR
		[23]));
	notech_mux2 i_2530(.S(n_60853), .A(n_6677), .B(axi_AR[23]), .Z(n_3330)
		);
	notech_nao3 i_622033(.A(n_2260), .B(n_2259), .C(n_1835), .Z(read_data[5]
		));
	notech_reg axi_AR_reg_24(.CP(n_61995), .D(n_3336), .CD(n_61429), .Q(axi_AR
		[24]));
	notech_mux2 i_2538(.S(n_60853), .A(n_6676), .B(axi_AR[24]), .Z(n_3336)
		);
	notech_reg axi_AR_reg_25(.CP(n_61995), .D(n_3342), .CD(n_61429), .Q(axi_AR
		[25]));
	notech_mux2 i_2546(.S(n_60853), .A(n_6675), .B(axi_AR[25]), .Z(n_3342)
		);
	notech_reg axi_AR_reg_26(.CP(n_61995), .D(n_3348), .CD(n_61429), .Q(axi_AR
		[26]));
	notech_mux2 i_2554(.S(n_60853), .A(n_6674), .B(axi_AR[26]), .Z(n_3348)
		);
	notech_reg axi_AR_reg_27(.CP(n_61995), .D(n_3354), .CD(n_61430), .Q(axi_AR
		[27]));
	notech_mux2 i_2562(.S(n_60853), .A(n_6672), .B(axi_AR[27]), .Z(n_3354)
		);
	notech_reg axi_AR_reg_28(.CP(n_61995), .D(n_3360), .CD(n_61430), .Q(axi_AR
		[28]));
	notech_mux2 i_2570(.S(n_60853), .A(n_6671), .B(axi_AR[28]), .Z(n_3360)
		);
	notech_and4 i_1215(.A(n_59537), .B(n_61512), .C(cacheQ[70]), .D(n_59463)
		, .Z(n_1841));
	notech_reg axi_AR_reg_29(.CP(n_61995), .D(n_3366), .CD(n_61429), .Q(axi_AR
		[29]));
	notech_mux2 i_2578(.S(n_60853), .A(n_6670), .B(axi_AR[29]), .Z(n_3366)
		);
	notech_nao3 i_722034(.A(n_2263), .B(n_2262), .C(n_1841), .Z(read_data[6]
		));
	notech_reg axi_AR_reg_30(.CP(n_61995), .D(n_3372), .CD(n_61429), .Q(axi_AR
		[30]));
	notech_mux2 i_2586(.S(n_60853), .A(n_6668), .B(axi_AR[30]), .Z(n_3372)
		);
	notech_reg axi_AR_reg_31(.CP(n_61995), .D(n_3378), .CD(n_61427), .Q(axi_AR
		[31]));
	notech_mux2 i_2594(.S(n_60853), .A(n_6667), .B(axi_AR[31]), .Z(n_3378)
		);
	notech_reg axi_AW_reg_0(.CP(n_61995), .D(n_3387), .CD(n_61425), .Q(axi_AW
		[0]));
	notech_and4 i_2604(.A(n_61496), .B(n_6763), .C(n_61523), .D(axi_AW[0]), 
		.Z(n_3387));
	notech_reg axi_AW_reg_1(.CP(n_61995), .D(n_3393), .CD(n_61425), .Q(axi_AW
		[1]));
	notech_and4 i_2612(.A(n_61496), .B(n_6763), .C(n_61523), .D(axi_AW[1]), 
		.Z(n_3393));
	notech_reg axi_AW_reg_2(.CP(n_61995), .D(n_3396), .CD(n_61425), .Q(axi_AW
		[2]));
	notech_mux2 i_2618(.S(n_61485), .A(n_6729), .B(axi_AW[2]), .Z(n_3396));
	notech_and4 i_1224(.A(n_59537), .B(n_61512), .C(cacheQ[71]), .D(n_59463)
		, .Z(n_1847));
	notech_reg axi_AW_reg_3(.CP(n_61995), .D(n_3402), .CD(n_61425), .Q(axi_AW
		[3]));
	notech_mux2 i_2626(.S(n_61485), .A(n_6728), .B(axi_AW[3]), .Z(n_3402));
	notech_nao3 i_822035(.A(n_2266), .B(n_2265), .C(n_1847), .Z(read_data[7]
		));
	notech_reg axi_AW_reg_4(.CP(n_62041), .D(n_3408), .CD(n_61426), .Q(axi_AW
		[4]));
	notech_mux2 i_2634(.S(n_61485), .A(n_6727), .B(axi_AW[4]), .Z(n_3408));
	notech_reg axi_AW_reg_5(.CP(n_61993), .D(n_3414), .CD(n_61426), .Q(axi_AW
		[5]));
	notech_mux2 i_2642(.S(n_61485), .A(n_6726), .B(axi_AW[5]), .Z(n_3414));
	notech_reg axi_AW_reg_6(.CP(n_62041), .D(n_3420), .CD(n_61426), .Q(axi_AW
		[6]));
	notech_mux2 i_2650(.S(n_61485), .A(n_6725), .B(axi_AW[6]), .Z(n_3420));
	notech_reg axi_AW_reg_7(.CP(n_62041), .D(n_3426), .CD(n_61426), .Q(axi_AW
		[7]));
	notech_mux2 i_2658(.S(n_61485), .A(n_6724), .B(axi_AW[7]), .Z(n_3426));
	notech_reg axi_AW_reg_8(.CP(n_62041), .D(n_3432), .CD(n_61425), .Q(axi_AW
		[8]));
	notech_mux2 i_2666(.S(n_61485), .A(n_6723), .B(axi_AW[8]), .Z(n_3432));
	notech_and4 i_1233(.A(n_59537), .B(n_61512), .C(cacheQ[72]), .D(n_59465)
		, .Z(n_1853));
	notech_reg axi_AW_reg_9(.CP(n_62041), .D(n_3438), .CD(n_61425), .Q(axi_AW
		[9]));
	notech_mux2 i_2674(.S(n_61485), .A(n_6722), .B(axi_AW[9]), .Z(n_3438));
	notech_nao3 i_922036(.A(n_2269), .B(n_2268), .C(n_1853), .Z(read_data[8]
		));
	notech_reg axi_AW_reg_10(.CP(n_62041), .D(n_3444), .CD(n_61425), .Q(axi_AW
		[10]));
	notech_mux2 i_2682(.S(n_61485), .A(n_6721), .B(axi_AW[10]), .Z(n_3444)
		);
	notech_reg axi_AW_reg_11(.CP(n_62041), .D(n_3450), .CD(n_61425), .Q(axi_AW
		[11]));
	notech_mux2 i_2690(.S(n_61485), .A(n_6720), .B(axi_AW[11]), .Z(n_3450)
		);
	notech_reg axi_AW_reg_12(.CP(n_62041), .D(n_3456), .CD(n_61425), .Q(axi_AW
		[12]));
	notech_mux2 i_2698(.S(n_61485), .A(n_6719), .B(axi_AW[12]), .Z(n_3456)
		);
	notech_reg axi_AW_reg_13(.CP(n_62041), .D(n_3462), .CD(n_61425), .Q(axi_AW
		[13]));
	notech_mux2 i_2706(.S(n_61485), .A(n_6718), .B(axi_AW[13]), .Z(n_3462)
		);
	notech_reg axi_AW_reg_14(.CP(n_62041), .D(n_3468), .CD(n_61425), .Q(axi_AW
		[14]));
	notech_mux2 i_2714(.S(n_61485), .A(n_6717), .B(axi_AW[14]), .Z(n_3468)
		);
	notech_and4 i_1242(.A(A4[1]), .B(n_61512), .C(cacheQ[73]), .D(n_59468), 
		.Z(n_1859));
	notech_reg axi_AW_reg_15(.CP(n_62041), .D(n_3474), .CD(n_61425), .Q(axi_AW
		[15]));
	notech_mux2 i_2722(.S(n_61486), .A(n_6716), .B(axi_AW[15]), .Z(n_3474)
		);
	notech_nao3 i_1022037(.A(n_2272), .B(n_2271), .C(n_1859), .Z(read_data[9
		]));
	notech_reg axi_AW_reg_16(.CP(n_62041), .D(n_3480), .CD(n_61426), .Q(axi_AW
		[16]));
	notech_mux2 i_2730(.S(n_61486), .A(n_6715), .B(axi_AW[16]), .Z(n_3480)
		);
	notech_reg axi_AW_reg_17(.CP(n_62041), .D(n_3486), .CD(n_61427), .Q(axi_AW
		[17]));
	notech_mux2 i_2738(.S(n_61486), .A(n_6714), .B(axi_AW[17]), .Z(n_3486)
		);
	notech_reg axi_AW_reg_18(.CP(n_62041), .D(n_3492), .CD(n_61427), .Q(axi_AW
		[18]));
	notech_mux2 i_2746(.S(n_61486), .A(n_6713), .B(axi_AW[18]), .Z(n_3492)
		);
	notech_reg axi_AW_reg_19(.CP(n_62041), .D(n_3498), .CD(n_61426), .Q(axi_AW
		[19]));
	notech_mux2 i_2754(.S(n_61486), .A(n_6712), .B(axi_AW[19]), .Z(n_3498)
		);
	notech_reg axi_AW_reg_20(.CP(n_62041), .D(n_3504), .CD(n_61426), .Q(axi_AW
		[20]));
	notech_mux2 i_2762(.S(n_61486), .A(n_6711), .B(axi_AW[20]), .Z(n_3504)
		);
	notech_and4 i_1251(.A(A4[1]), .B(n_61512), .C(cacheQ[74]), .D(n_59468), 
		.Z(n_1865));
	notech_reg axi_AW_reg_21(.CP(n_62041), .D(n_3510), .CD(n_61427), .Q(axi_AW
		[21]));
	notech_mux2 i_2770(.S(n_61486), .A(n_6710), .B(axi_AW[21]), .Z(n_3510)
		);
	notech_nao3 i_1122038(.A(n_2275), .B(n_2274), .C(n_1865), .Z(read_data[
		10]));
	notech_reg axi_AW_reg_22(.CP(n_62041), .D(n_3516), .CD(n_61427), .Q(axi_AW
		[22]));
	notech_mux2 i_2778(.S(n_61486), .A(n_6709), .B(axi_AW[22]), .Z(n_3516)
		);
	notech_reg axi_AW_reg_23(.CP(n_62019), .D(n_3522), .CD(n_61427), .Q(axi_AW
		[23]));
	notech_mux2 i_2786(.S(n_61486), .A(n_6708), .B(axi_AW[23]), .Z(n_3522)
		);
	notech_reg axi_AW_reg_24(.CP(n_61993), .D(n_3528), .CD(n_61427), .Q(axi_AW
		[24]));
	notech_mux2 i_2794(.S(n_61486), .A(n_6707), .B(axi_AW[24]), .Z(n_3528)
		);
	notech_reg axi_AW_reg_25(.CP(n_61993), .D(n_3534), .CD(n_61426), .Q(axi_AW
		[25]));
	notech_mux2 i_2802(.S(n_61486), .A(n_6706), .B(axi_AW[25]), .Z(n_3534)
		);
	notech_reg axi_AW_reg_26(.CP(n_61993), .D(n_3540), .CD(n_61426), .Q(axi_AW
		[26]));
	notech_mux2 i_2810(.S(n_61486), .A(n_6704), .B(axi_AW[26]), .Z(n_3540)
		);
	notech_and4 i_1260(.A(A4[1]), .B(n_61512), .C(cacheQ[75]), .D(n_59468), 
		.Z(n_1871));
	notech_reg axi_AW_reg_27(.CP(n_61993), .D(n_3546), .CD(n_61426), .Q(axi_AW
		[27]));
	notech_mux2 i_2818(.S(n_61486), .A(n_6703), .B(axi_AW[27]), .Z(n_3546)
		);
	notech_nao3 i_1222039(.A(n_2278), .B(n_2277), .C(n_1871), .Z(read_data[
		11]));
	notech_reg axi_AW_reg_28(.CP(n_61993), .D(n_3552), .CD(n_61426), .Q(axi_AW
		[28]));
	notech_mux2 i_2826(.S(n_61486), .A(n_6702), .B(axi_AW[28]), .Z(n_3552)
		);
	notech_reg axi_AW_reg_29(.CP(n_61993), .D(n_3558), .CD(n_61426), .Q(axi_AW
		[29]));
	notech_mux2 i_2834(.S(n_61486), .A(n_6701), .B(axi_AW[29]), .Z(n_3558)
		);
	notech_reg axi_AW_reg_30(.CP(n_61993), .D(n_3564), .CD(n_61426), .Q(axi_AW
		[30]));
	notech_mux2 i_2842(.S(n_61486), .A(n_6700), .B(axi_AW[30]), .Z(n_3564)
		);
	notech_reg axi_AW_reg_31(.CP(n_61993), .D(n_3570), .CD(n_61426), .Q(axi_AW
		[31]));
	notech_mux2 i_2850(.S(n_61486), .A(n_6699), .B(axi_AW[31]), .Z(n_3570)
		);
	notech_reg_set burst_idx_reg_0(.CP(n_61993), .D(n_3576), .SD(1'b1), .Q(burst_idx
		[0]));
	notech_mux2 i_2858(.S(n_1171), .A(n_6730), .B(burst_idx[0]), .Z(n_3576)
		);
	notech_and4 i_1269(.A(A4[1]), .B(n_61512), .C(cacheQ[76]), .D(n_59468), 
		.Z(n_1877));
	notech_reg_set burst_idx_reg_1(.CP(n_61993), .D(n_3582), .SD(1'b1), .Q(burst_idx
		[1]));
	notech_mux2 i_2866(.S(n_1171), .A(n_25530), .B(burst_idx[1]), .Z(n_3582)
		);
	notech_nao3 i_1322040(.A(n_2281), .B(n_2280), .C(n_1877), .Z(read_data[
		12]));
	notech_reg_set burst_idx_reg_2(.CP(n_61993), .D(n_3588), .SD(1'b1), .Q(burst_idx
		[2]));
	notech_mux2 i_2874(.S(n_1171), .A(n_25535), .B(burst_idx[2]), .Z(n_3588)
		);
	notech_reg_set burst_idx_reg_3(.CP(n_61993), .D(n_3594), .SD(1'b1), .Q(burst_idx
		[3]));
	notech_mux2 i_2882(.S(n_1171), .A(n_25540), .B(burst_idx[3]), .Z(n_3594)
		);
	notech_reg_set burst_idx_reg_4(.CP(n_61993), .D(n_3600), .SD(1'b1), .Q(burst_idx
		[4]));
	notech_mux2 i_2890(.S(n_1171), .A(n_25545), .B(burst_idx[4]), .Z(n_3600)
		);
	notech_reg axi_AWVALID_reg(.CP(n_61993), .D(n_3606), .CD(n_61426), .Q(axi_AWVALID
		));
	notech_mux2 i_2898(.S(n_1175), .A(n_1176), .B(axi_AWVALID), .Z(n_3606)
		);
	notech_reg_set A4_reg_0(.CP(n_61993), .D(n_3612), .SD(1'b1), .Q(A4[0])
		);
	notech_mux2 i_2906(.S(\nbus_11672[0] ), .A(n_59508), .B(Daddr[2]), .Z(n_3612
		));
	notech_and4 i_1278(.A(A4[1]), .B(n_61512), .C(cacheQ[77]), .D(n_59468), 
		.Z(n_1883));
	notech_reg_set A4_reg_1(.CP(n_61993), .D(n_3618), .SD(1'b1), .Q(A4[1])
		);
	notech_mux2 i_2914(.S(\nbus_11672[0] ), .A(A4[1]), .B(Daddr[3]), .Z(n_3618
		));
	notech_nao3 i_1422041(.A(n_2284), .B(n_2283), .C(n_1883), .Z(read_data[
		13]));
	notech_reg axi_W_reg_0(.CP(n_61993), .D(n_3624), .CD(n_61433), .Q(axi_W[
		0]));
	notech_mux2 i_2922(.S(n_61486), .A(n_6738), .B(axi_W[0]), .Z(n_3624));
	notech_reg axi_W_reg_1(.CP(n_61993), .D(n_3630), .CD(n_61433), .Q(axi_W[
		1]));
	notech_mux2 i_2930(.S(n_61485), .A(n_6737), .B(axi_W[1]), .Z(n_3630));
	notech_reg axi_W_reg_2(.CP(n_62041), .D(n_3636), .CD(n_61433), .Q(axi_W[
		2]));
	notech_mux2 i_2938(.S(n_61475), .A(n_6736), .B(axi_W[2]), .Z(n_3636));
	notech_reg axi_W_reg_3(.CP(n_62015), .D(n_3642), .CD(n_61433), .Q(axi_W[
		3]));
	notech_mux2 i_2946(.S(n_61475), .A(n_6735), .B(axi_W[3]), .Z(n_3642));
	notech_reg axi_W_reg_4(.CP(n_61991), .D(n_3648), .CD(n_61433), .Q(axi_W[
		4]));
	notech_mux2 i_2954(.S(n_61475), .A(n_6734), .B(axi_W[4]), .Z(n_3648));
	notech_and4 i_1287(.A(A4[1]), .B(n_61512), .C(cacheQ[78]), .D(n_59468), 
		.Z(n_1889));
	notech_reg axi_W_reg_5(.CP(n_62015), .D(n_3654), .CD(n_61433), .Q(axi_W[
		5]));
	notech_mux2 i_2962(.S(n_61475), .A(n_6733), .B(axi_W[5]), .Z(n_3654));
	notech_nao3 i_1522042(.A(n_2287), .B(n_2286), .C(n_1889), .Z(read_data[
		14]));
	notech_reg axi_W_reg_6(.CP(n_62015), .D(n_3660), .CD(n_61433), .Q(axi_W[
		6]));
	notech_mux2 i_2970(.S(n_61475), .A(n_6732), .B(axi_W[6]), .Z(n_3660));
	notech_reg axi_W_reg_7(.CP(n_62015), .D(n_3666), .CD(n_61433), .Q(axi_W[
		7]));
	notech_mux2 i_2978(.S(n_61475), .A(n_6731), .B(axi_W[7]), .Z(n_3666));
	notech_reg axi_W_reg_8(.CP(n_62015), .D(n_3672), .CD(n_61433), .Q(axi_W[
		8]));
	notech_mux2 i_2986(.S(n_61475), .A(n_24863), .B(axi_W[8]), .Z(n_3672));
	notech_reg axi_W_reg_9(.CP(n_62015), .D(n_3678), .CD(n_61433), .Q(axi_W[
		9]));
	notech_mux2 i_2994(.S(n_61475), .A(n_24869), .B(axi_W[9]), .Z(n_3678));
	notech_reg axi_W_reg_10(.CP(n_62015), .D(n_3684), .CD(n_61432), .Q(axi_W
		[10]));
	notech_mux2 i_3002(.S(n_61475), .A(n_24875), .B(axi_W[10]), .Z(n_3684)
		);
	notech_and4 i_1296(.A(A4[1]), .B(n_61512), .C(cacheQ[79]), .D(n_59468), 
		.Z(n_1895));
	notech_reg axi_W_reg_11(.CP(n_62015), .D(n_3690), .CD(n_61433), .Q(axi_W
		[11]));
	notech_mux2 i_3010(.S(n_61475), .A(n_24881), .B(axi_W[11]), .Z(n_3690)
		);
	notech_nao3 i_1622043(.A(n_2290), .B(n_2289), .C(n_1895), .Z(read_data[
		15]));
	notech_reg axi_W_reg_12(.CP(n_62015), .D(n_3696), .CD(n_61433), .Q(axi_W
		[12]));
	notech_mux2 i_3018(.S(n_61475), .A(n_24887), .B(axi_W[12]), .Z(n_3696)
		);
	notech_reg axi_W_reg_13(.CP(n_62015), .D(n_3702), .CD(n_61433), .Q(axi_W
		[13]));
	notech_mux2 i_3026(.S(n_61475), .A(n_24893), .B(axi_W[13]), .Z(n_3702)
		);
	notech_reg axi_W_reg_14(.CP(n_62015), .D(n_3708), .CD(n_61433), .Q(axi_W
		[14]));
	notech_mux2 i_3034(.S(n_61475), .A(n_24899), .B(axi_W[14]), .Z(n_3708)
		);
	notech_reg axi_W_reg_15(.CP(n_62015), .D(n_3714), .CD(n_61433), .Q(axi_W
		[15]));
	notech_mux2 i_3042(.S(n_61475), .A(n_24905), .B(axi_W[15]), .Z(n_3714)
		);
	notech_reg axi_W_reg_16(.CP(n_62015), .D(n_3720), .CD(n_61433), .Q(axi_W
		[16]));
	notech_mux2 i_3050(.S(n_61475), .A(n_24911), .B(axi_W[16]), .Z(n_3720)
		);
	notech_and4 i_1305(.A(A4[1]), .B(n_61513), .C(cacheQ[80]), .D(n_59468), 
		.Z(n_1901));
	notech_reg axi_W_reg_17(.CP(n_62015), .D(n_3726), .CD(n_61434), .Q(axi_W
		[17]));
	notech_mux2 i_3058(.S(n_61475), .A(n_24917), .B(axi_W[17]), .Z(n_3726)
		);
	notech_nao3 i_1722044(.A(n_2293), .B(n_2292), .C(n_1901), .Z(read_data[
		16]));
	notech_reg axi_W_reg_18(.CP(n_62015), .D(n_3732), .CD(n_61434), .Q(axi_W
		[18]));
	notech_mux2 i_3066(.S(n_61475), .A(n_24923), .B(axi_W[18]), .Z(n_3732)
		);
	notech_reg axi_W_reg_19(.CP(n_62015), .D(n_3738), .CD(n_61434), .Q(axi_W
		[19]));
	notech_mux2 i_3074(.S(n_61480), .A(n_24929), .B(axi_W[19]), .Z(n_3738)
		);
	notech_reg axi_W_reg_20(.CP(n_62015), .D(n_3744), .CD(n_61434), .Q(axi_W
		[20]));
	notech_mux2 i_3082(.S(n_61480), .A(n_24935), .B(axi_W[20]), .Z(n_3744)
		);
	notech_reg axi_W_reg_21(.CP(n_62015), .D(n_3750), .CD(n_61434), .Q(axi_W
		[21]));
	notech_mux2 i_3090(.S(n_61480), .A(n_24941), .B(axi_W[21]), .Z(n_3750)
		);
	notech_reg axi_W_reg_22(.CP(n_62051), .D(n_3756), .CD(n_61434), .Q(axi_W
		[22]));
	notech_mux2 i_3098(.S(n_61480), .A(n_24947), .B(axi_W[22]), .Z(n_3756)
		);
	notech_and4 i_1314(.A(A4[1]), .B(n_61513), .C(cacheQ[81]), .D(n_59468), 
		.Z(n_1907));
	notech_reg axi_W_reg_23(.CP(n_62037), .D(n_3762), .CD(n_61434), .Q(axi_W
		[23]));
	notech_mux2 i_3106(.S(n_61480), .A(n_24953), .B(axi_W[23]), .Z(n_3762)
		);
	notech_nao3 i_1822045(.A(n_2296), .B(n_2295), .C(n_1907), .Z(read_data[
		17]));
	notech_reg axi_W_reg_24(.CP(n_62051), .D(n_3768), .CD(n_61434), .Q(axi_W
		[24]));
	notech_mux2 i_3114(.S(n_61480), .A(n_24959), .B(axi_W[24]), .Z(n_3768)
		);
	notech_reg axi_W_reg_25(.CP(n_62051), .D(n_3774), .CD(n_61434), .Q(axi_W
		[25]));
	notech_mux2 i_3122(.S(n_61480), .A(n_24965), .B(axi_W[25]), .Z(n_3774)
		);
	notech_reg axi_W_reg_26(.CP(n_62051), .D(n_3780), .CD(n_61434), .Q(axi_W
		[26]));
	notech_mux2 i_3130(.S(n_61480), .A(n_24971), .B(axi_W[26]), .Z(n_3780)
		);
	notech_reg axi_W_reg_27(.CP(n_62051), .D(n_3786), .CD(n_61434), .Q(axi_W
		[27]));
	notech_mux2 i_3138(.S(n_61480), .A(n_24977), .B(axi_W[27]), .Z(n_3786)
		);
	notech_reg axi_W_reg_28(.CP(n_62051), .D(n_3792), .CD(n_61434), .Q(axi_W
		[28]));
	notech_mux2 i_3146(.S(n_61480), .A(n_24983), .B(axi_W[28]), .Z(n_3792)
		);
	notech_and4 i_1323(.A(A4[1]), .B(n_61513), .C(cacheQ[82]), .D(n_59468), 
		.Z(n_1913));
	notech_reg axi_W_reg_29(.CP(n_62051), .D(n_3798), .CD(n_61434), .Q(axi_W
		[29]));
	notech_mux2 i_3154(.S(n_61480), .A(n_24989), .B(axi_W[29]), .Z(n_3798)
		);
	notech_nao3 i_1922046(.A(n_2299), .B(n_2298), .C(n_1913), .Z(read_data[
		18]));
	notech_reg axi_W_reg_30(.CP(n_62051), .D(n_3804), .CD(n_61434), .Q(axi_W
		[30]));
	notech_mux2 i_3162(.S(n_61480), .A(n_24995), .B(axi_W[30]), .Z(n_3804)
		);
	notech_reg axi_W_reg_31(.CP(n_62051), .D(n_3810), .CD(n_61434), .Q(axi_W
		[31]));
	notech_mux2 i_3170(.S(n_61480), .A(n_25001), .B(axi_W[31]), .Z(n_3810)
		);
	notech_reg abort_reg(.CP(n_62051), .D(n_3816), .CD(n_61434), .Q(abort)
		);
	notech_mux2 i_3178(.S(n_1203), .A(n_1204), .B(abort), .Z(n_3816));
	notech_reg read_ack_slow_reg(.CP(n_62051), .D(n_3822), .CD(n_61432), .Q(read_ack
		));
	notech_mux2 i_3186(.S(n_1208), .A(n_1210), .B(read_ack), .Z(n_3822));
	notech_reg wrint_ack_reg(.CP(n_62051), .D(n_3828), .CD(n_61431), .Q(write_ack
		));
	notech_mux2 i_3194(.S(n_1211), .A(n_23592), .B(write_ack), .Z(n_3828));
	notech_and4 i_1332(.A(n_59537), .B(n_61513), .C(cacheQ[83]), .D(n_59468)
		, .Z(n_1919));
	notech_reg fsm_reg_0(.CP(n_62051), .D(n_3834), .CD(n_61431), .Q(fsm[0])
		);
	notech_mux2 i_3202(.S(n_1222), .A(n_6741), .B(fsm[0]), .Z(n_3834));
	notech_nao3 i_2022047(.A(n_2302), .B(n_2301), .C(n_1919), .Z(read_data[
		19]));
	notech_reg fsm_reg_1(.CP(n_62051), .D(n_3840), .CD(n_61431), .Q(fsm[1])
		);
	notech_mux2 i_3210(.S(n_1222), .A(n_1216), .B(fsm[1]), .Z(n_3840));
	notech_reg fsm_reg_2(.CP(n_62051), .D(n_3846), .CD(n_61431), .Q(fsm[2])
		);
	notech_mux2 i_3218(.S(n_1222), .A(n_1214), .B(fsm[2]), .Z(n_3846));
	notech_reg fsm_reg_3(.CP(n_62051), .D(n_3852), .CD(n_61431), .Q(fsm[3])
		);
	notech_mux2 i_3226(.S(n_1222), .A(n_6739), .B(fsm[3]), .Z(n_3852));
	notech_reg fsm_reg_4(.CP(n_62051), .D(n_3858), .CD(n_61431), .Q(fsm[4])
		);
	notech_mux2 i_3234(.S(n_1222), .A(n_1212), .B(fsm[4]), .Z(n_3858));
	notech_reg_set cacheD_reg_0(.CP(n_62051), .D(n_3864), .SD(1'b1), .Q(cacheD
		[0]));
	notech_mux2 i_3242(.S(n_1703), .A(n_1708), .B(cacheD[0]), .Z(n_3864));
	notech_and4 i_1341(.A(n_59533), .B(n_61513), .C(cacheQ[84]), .D(n_59468)
		, .Z(n_1925));
	notech_reg_set cacheD_reg_1(.CP(n_62015), .D(n_3870), .SD(1'b1), .Q(cacheD
		[1]));
	notech_mux2 i_3250(.S(n_1703), .A(n_1701), .B(cacheD[1]), .Z(n_3870));
	notech_nao3 i_2122048(.A(n_2305), .B(n_2304), .C(n_1925), .Z(read_data[
		20]));
	notech_reg_set cacheD_reg_2(.CP(n_62051), .D(n_3876), .SD(1'b1), .Q(cacheD
		[2]));
	notech_mux2 i_3258(.S(n_1703), .A(n_1697), .B(cacheD[2]), .Z(n_3876));
	notech_reg_set cacheD_reg_3(.CP(n_62039), .D(n_3882), .SD(1'b1), .Q(cacheD
		[3]));
	notech_mux2 i_3266(.S(n_1703), .A(n_1693), .B(cacheD[3]), .Z(n_3882));
	notech_reg_set cacheD_reg_4(.CP(n_62039), .D(n_3888), .SD(1'b1), .Q(cacheD
		[4]));
	notech_mux2 i_3274(.S(n_1703), .A(n_1689), .B(cacheD[4]), .Z(n_3888));
	notech_reg_set cacheD_reg_5(.CP(n_62039), .D(n_3894), .SD(1'b1), .Q(cacheD
		[5]));
	notech_mux2 i_3282(.S(n_1703), .A(n_1685), .B(cacheD[5]), .Z(n_3894));
	notech_reg_set cacheD_reg_6(.CP(n_62039), .D(n_3900), .SD(1'b1), .Q(cacheD
		[6]));
	notech_mux2 i_3290(.S(n_1703), .A(n_1681), .B(cacheD[6]), .Z(n_3900));
	notech_and4 i_1350(.A(n_59533), .B(n_61513), .C(cacheQ[85]), .D(n_59468)
		, .Z(n_1931));
	notech_reg_set cacheD_reg_7(.CP(n_62039), .D(n_3906), .SD(1'b1), .Q(cacheD
		[7]));
	notech_mux2 i_3298(.S(n_1703), .A(n_1677), .B(cacheD[7]), .Z(n_3906));
	notech_nao3 i_2222049(.A(n_2308), .B(n_2307), .C(n_1931), .Z(read_data[
		21]));
	notech_reg_set cacheD_reg_8(.CP(n_62039), .D(n_3912), .SD(1'b1), .Q(cacheD
		[8]));
	notech_mux2 i_3306(.S(n_1703), .A(n_1673), .B(cacheD[8]), .Z(n_3912));
	notech_reg_set cacheD_reg_9(.CP(n_62039), .D(n_3918), .SD(1'b1), .Q(cacheD
		[9]));
	notech_mux2 i_3314(.S(n_1703), .A(n_1669), .B(cacheD[9]), .Z(n_3918));
	notech_reg_set cacheD_reg_10(.CP(n_62039), .D(n_3924), .SD(1'b1), .Q(cacheD
		[10]));
	notech_mux2 i_3322(.S(n_1703), .A(n_1665), .B(cacheD[10]), .Z(n_3924));
	notech_reg_set cacheD_reg_11(.CP(n_62039), .D(n_3930), .SD(1'b1), .Q(cacheD
		[11]));
	notech_mux2 i_3330(.S(n_1703), .A(n_1661), .B(cacheD[11]), .Z(n_3930));
	notech_reg_set cacheD_reg_12(.CP(n_62039), .D(n_3936), .SD(1'b1), .Q(cacheD
		[12]));
	notech_mux2 i_3338(.S(n_1703), .A(n_1657), .B(cacheD[12]), .Z(n_3936));
	notech_and4 i_1359(.A(n_59533), .B(n_61513), .C(cacheQ[86]), .D(n_59465)
		, .Z(n_1937));
	notech_reg_set cacheD_reg_13(.CP(n_62039), .D(n_3942), .SD(1'b1), .Q(cacheD
		[13]));
	notech_mux2 i_3346(.S(n_1703), .A(n_1653), .B(cacheD[13]), .Z(n_3942));
	notech_nao3 i_2322050(.A(n_2311), .B(n_2310), .C(n_1937), .Z(read_data[
		22]));
	notech_reg_set cacheD_reg_14(.CP(n_62039), .D(n_3948), .SD(1'b1), .Q(cacheD
		[14]));
	notech_mux2 i_3354(.S(n_1703), .A(n_1649), .B(cacheD[14]), .Z(n_3948));
	notech_reg_set cacheD_reg_15(.CP(n_62039), .D(n_3954), .SD(1'b1), .Q(cacheD
		[15]));
	notech_mux2 i_3362(.S(n_1703), .A(n_1645), .B(cacheD[15]), .Z(n_3954));
	notech_reg_set cacheD_reg_16(.CP(n_62039), .D(n_3960), .SD(1'b1), .Q(cacheD
		[16]));
	notech_mux2 i_3370(.S(n_59397), .A(n_1641), .B(cacheD[16]), .Z(n_3960)
		);
	notech_reg_set cacheD_reg_17(.CP(n_62039), .D(n_3966), .SD(1'b1), .Q(cacheD
		[17]));
	notech_mux2 i_3378(.S(n_59397), .A(n_1637), .B(cacheD[17]), .Z(n_3966)
		);
	notech_reg_set cacheD_reg_18(.CP(n_62039), .D(n_3972), .SD(1'b1), .Q(cacheD
		[18]));
	notech_mux2 i_3386(.S(n_59397), .A(n_1633), .B(cacheD[18]), .Z(n_3972)
		);
	notech_and4 i_1368(.A(n_59537), .B(n_61513), .C(cacheQ[87]), .D(n_59465)
		, .Z(n_1943));
	notech_reg_set cacheD_reg_19(.CP(n_62039), .D(n_3978), .SD(1'b1), .Q(cacheD
		[19]));
	notech_mux2 i_3394(.S(n_59397), .A(n_1629), .B(cacheD[19]), .Z(n_3978)
		);
	notech_nao3 i_2422051(.A(n_2314), .B(n_2313), .C(n_1943), .Z(read_data[
		23]));
	notech_reg_set cacheD_reg_20(.CP(n_62039), .D(n_3984), .SD(1'b1), .Q(cacheD
		[20]));
	notech_mux2 i_3402(.S(n_59397), .A(n_1625), .B(cacheD[20]), .Z(n_3984)
		);
	notech_reg_set cacheD_reg_21(.CP(n_62017), .D(n_3990), .SD(1'b1), .Q(cacheD
		[21]));
	notech_mux2 i_3410(.S(n_59397), .A(n_1621), .B(cacheD[21]), .Z(n_3990)
		);
	notech_reg_set cacheD_reg_22(.CP(n_61991), .D(n_3996), .SD(1'b1), .Q(cacheD
		[22]));
	notech_mux2 i_3418(.S(n_59397), .A(n_1617), .B(cacheD[22]), .Z(n_3996)
		);
	notech_reg_set cacheD_reg_23(.CP(n_61991), .D(n_4002), .SD(1'b1), .Q(cacheD
		[23]));
	notech_mux2 i_3426(.S(n_59397), .A(n_1613), .B(cacheD[23]), .Z(n_4002)
		);
	notech_reg_set cacheD_reg_24(.CP(n_61991), .D(n_4008), .SD(1'b1), .Q(cacheD
		[24]));
	notech_mux2 i_3434(.S(n_59397), .A(n_1609), .B(cacheD[24]), .Z(n_4008)
		);
	notech_and4 i_1377(.A(n_59537), .B(n_61513), .C(cacheQ[88]), .D(n_59465)
		, .Z(n_1949));
	notech_reg_set cacheD_reg_25(.CP(n_61991), .D(n_4014), .SD(1'b1), .Q(cacheD
		[25]));
	notech_mux2 i_3442(.S(n_59397), .A(n_1605), .B(cacheD[25]), .Z(n_4014)
		);
	notech_nao3 i_2522052(.A(n_2317), .B(n_2316), .C(n_1949), .Z(read_data[
		24]));
	notech_reg_set cacheD_reg_26(.CP(n_61991), .D(n_4020), .SD(1'b1), .Q(cacheD
		[26]));
	notech_mux2 i_3450(.S(n_59397), .A(n_1601), .B(cacheD[26]), .Z(n_4020)
		);
	notech_reg_set cacheD_reg_27(.CP(n_61991), .D(n_4026), .SD(1'b1), .Q(cacheD
		[27]));
	notech_mux2 i_3458(.S(n_59397), .A(n_1597), .B(cacheD[27]), .Z(n_4026)
		);
	notech_reg_set cacheD_reg_28(.CP(n_61991), .D(n_4032), .SD(1'b1), .Q(cacheD
		[28]));
	notech_mux2 i_3466(.S(n_59397), .A(n_1593), .B(cacheD[28]), .Z(n_4032)
		);
	notech_reg_set cacheD_reg_29(.CP(n_61991), .D(n_4038), .SD(1'b1), .Q(cacheD
		[29]));
	notech_mux2 i_3474(.S(n_59397), .A(n_1589), .B(cacheD[29]), .Z(n_4038)
		);
	notech_reg_set cacheD_reg_30(.CP(n_61991), .D(n_4044), .SD(1'b1), .Q(cacheD
		[30]));
	notech_mux2 i_3482(.S(n_59397), .A(n_1585), .B(cacheD[30]), .Z(n_4044)
		);
	notech_and4 i_1386(.A(n_59533), .B(n_61513), .C(cacheQ[89]), .D(n_59465)
		, .Z(n_1955));
	notech_reg_set cacheD_reg_31(.CP(n_61991), .D(n_4050), .SD(1'b1), .Q(cacheD
		[31]));
	notech_mux2 i_3490(.S(n_59397), .A(n_1581), .B(cacheD[31]), .Z(n_4050)
		);
	notech_nao3 i_2622053(.A(n_2320), .B(n_2319), .C(n_1955), .Z(read_data[
		25]));
	notech_reg_set cacheD_reg_32(.CP(n_61991), .D(n_4056), .SD(1'b1), .Q(cacheD
		[32]));
	notech_mux2 i_3498(.S(n_1573), .A(n_1577), .B(cacheD[32]), .Z(n_4056));
	notech_reg_set cacheD_reg_33(.CP(n_61991), .D(n_4062), .SD(1'b1), .Q(cacheD
		[33]));
	notech_mux2 i_3506(.S(n_1573), .A(n_1571), .B(cacheD[33]), .Z(n_4062));
	notech_reg_set cacheD_reg_34(.CP(n_61991), .D(n_4068), .SD(1'b1), .Q(cacheD
		[34]));
	notech_mux2 i_3514(.S(n_1573), .A(n_1568), .B(cacheD[34]), .Z(n_4068));
	notech_reg_set cacheD_reg_35(.CP(n_61991), .D(n_4074), .SD(1'b1), .Q(cacheD
		[35]));
	notech_mux2 i_3522(.S(n_1573), .A(n_1565), .B(cacheD[35]), .Z(n_4074));
	notech_reg_set cacheD_reg_36(.CP(n_61991), .D(n_4080), .SD(1'b1), .Q(cacheD
		[36]));
	notech_mux2 i_3530(.S(n_1573), .A(n_1562), .B(cacheD[36]), .Z(n_4080));
	notech_and4 i_1395(.A(n_59533), .B(n_61513), .C(cacheQ[90]), .D(n_59465)
		, .Z(n_1961));
	notech_reg_set cacheD_reg_37(.CP(n_61991), .D(n_4086), .SD(1'b1), .Q(cacheD
		[37]));
	notech_mux2 i_3538(.S(n_1573), .A(n_1559), .B(cacheD[37]), .Z(n_4086));
	notech_nao3 i_2722054(.A(n_2323), .B(n_2322), .C(n_1961), .Z(read_data[
		26]));
	notech_reg_set cacheD_reg_38(.CP(n_61991), .D(n_4092), .SD(1'b1), .Q(cacheD
		[38]));
	notech_mux2 i_3546(.S(n_1573), .A(n_1556), .B(cacheD[38]), .Z(n_4092));
	notech_reg_set cacheD_reg_39(.CP(n_61991), .D(n_4098), .SD(1'b1), .Q(cacheD
		[39]));
	notech_mux2 i_3554(.S(n_1573), .A(n_1553), .B(cacheD[39]), .Z(n_4098));
	notech_reg_set cacheD_reg_40(.CP(n_62039), .D(n_4104), .SD(1'b1), .Q(cacheD
		[40]));
	notech_mux2 i_3562(.S(n_1573), .A(n_1550), .B(cacheD[40]), .Z(n_4104));
	notech_reg_set cacheD_reg_41(.CP(n_62009), .D(n_4110), .SD(1'b1), .Q(cacheD
		[41]));
	notech_mux2 i_3570(.S(n_1573), .A(n_1547), .B(cacheD[41]), .Z(n_4110));
	notech_reg_set cacheD_reg_42(.CP(n_62009), .D(n_4116), .SD(1'b1), .Q(cacheD
		[42]));
	notech_mux2 i_3578(.S(n_1573), .A(n_1544), .B(cacheD[42]), .Z(n_4116));
	notech_and4 i_1404(.A(n_59533), .B(n_61513), .C(cacheQ[91]), .D(n_59465)
		, .Z(n_1967));
	notech_reg_set cacheD_reg_43(.CP(n_62009), .D(n_4122), .SD(1'b1), .Q(cacheD
		[43]));
	notech_mux2 i_3586(.S(n_1573), .A(n_1541), .B(cacheD[43]), .Z(n_4122));
	notech_nao3 i_2822055(.A(n_2326), .B(n_2325), .C(n_1967), .Z(read_data[
		27]));
	notech_reg_set cacheD_reg_44(.CP(n_62009), .D(n_4128), .SD(1'b1), .Q(cacheD
		[44]));
	notech_mux2 i_3594(.S(n_1573), .A(n_1538), .B(cacheD[44]), .Z(n_4128));
	notech_reg_set cacheD_reg_45(.CP(n_62009), .D(n_4134), .SD(1'b1), .Q(cacheD
		[45]));
	notech_mux2 i_3602(.S(n_1573), .A(n_1535), .B(cacheD[45]), .Z(n_4134));
	notech_reg_set cacheD_reg_46(.CP(n_62009), .D(n_4140), .SD(1'b1), .Q(cacheD
		[46]));
	notech_mux2 i_3610(.S(n_1573), .A(n_1532), .B(cacheD[46]), .Z(n_4140));
	notech_reg_set cacheD_reg_47(.CP(n_62009), .D(n_4146), .SD(1'b1), .Q(cacheD
		[47]));
	notech_mux2 i_3618(.S(n_1573), .A(n_1529), .B(cacheD[47]), .Z(n_4146));
	notech_reg_set cacheD_reg_48(.CP(n_62009), .D(n_4152), .SD(1'b1), .Q(cacheD
		[48]));
	notech_mux2 i_3626(.S(n_59419), .A(n_1526), .B(cacheD[48]), .Z(n_4152)
		);
	notech_and4 i_1413(.A(n_59533), .B(n_61513), .C(cacheQ[92]), .D(n_59465)
		, .Z(n_1973));
	notech_reg_set cacheD_reg_49(.CP(n_62009), .D(n_4158), .SD(1'b1), .Q(cacheD
		[49]));
	notech_mux2 i_3634(.S(n_59419), .A(n_1523), .B(cacheD[49]), .Z(n_4158)
		);
	notech_nao3 i_2922056(.A(n_2329), .B(n_2328), .C(n_1973), .Z(read_data[
		28]));
	notech_reg_set cacheD_reg_50(.CP(n_62009), .D(n_4164), .SD(1'b1), .Q(cacheD
		[50]));
	notech_mux2 i_3642(.S(n_59419), .A(n_1520), .B(cacheD[50]), .Z(n_4164)
		);
	notech_reg_set cacheD_reg_51(.CP(n_62009), .D(n_4170), .SD(1'b1), .Q(cacheD
		[51]));
	notech_mux2 i_3650(.S(n_59419), .A(n_1517), .B(cacheD[51]), .Z(n_4170)
		);
	notech_reg_set cacheD_reg_52(.CP(n_62009), .D(n_4176), .SD(1'b1), .Q(cacheD
		[52]));
	notech_mux2 i_3658(.S(n_59419), .A(n_1514), .B(cacheD[52]), .Z(n_4176)
		);
	notech_reg_set cacheD_reg_53(.CP(n_62009), .D(n_4182), .SD(1'b1), .Q(cacheD
		[53]));
	notech_mux2 i_3666(.S(n_59419), .A(n_1511), .B(cacheD[53]), .Z(n_4182)
		);
	notech_reg_set cacheD_reg_54(.CP(n_62009), .D(n_4188), .SD(1'b1), .Q(cacheD
		[54]));
	notech_mux2 i_3674(.S(n_59419), .A(n_1508), .B(cacheD[54]), .Z(n_4188)
		);
	notech_and4 i_1422(.A(n_59533), .B(n_61513), .C(cacheQ[93]), .D(n_59468)
		, .Z(n_1979));
	notech_reg_set cacheD_reg_55(.CP(n_62009), .D(n_4194), .SD(1'b1), .Q(cacheD
		[55]));
	notech_mux2 i_3682(.S(n_59419), .A(n_1505), .B(cacheD[55]), .Z(n_4194)
		);
	notech_nao3 i_3022057(.A(n_2332), .B(n_2331), .C(n_1979), .Z(read_data[
		29]));
	notech_reg_set cacheD_reg_56(.CP(n_62009), .D(n_4200), .SD(1'b1), .Q(cacheD
		[56]));
	notech_mux2 i_3690(.S(n_59419), .A(n_1502), .B(cacheD[56]), .Z(n_4200)
		);
	notech_reg_set cacheD_reg_57(.CP(n_62009), .D(n_4206), .SD(1'b1), .Q(cacheD
		[57]));
	notech_mux2 i_3698(.S(n_59419), .A(n_1499), .B(cacheD[57]), .Z(n_4206)
		);
	notech_reg_set cacheD_reg_58(.CP(n_62009), .D(n_4212), .SD(1'b1), .Q(cacheD
		[58]));
	notech_mux2 i_3706(.S(n_59419), .A(n_1496), .B(cacheD[58]), .Z(n_4212)
		);
	notech_reg_set cacheD_reg_59(.CP(n_62009), .D(n_4218), .SD(1'b1), .Q(cacheD
		[59]));
	notech_mux2 i_3714(.S(n_59419), .A(n_1493), .B(cacheD[59]), .Z(n_4218)
		);
	notech_reg_set cacheD_reg_60(.CP(n_62047), .D(n_4224), .SD(1'b1), .Q(cacheD
		[60]));
	notech_mux2 i_3722(.S(n_59419), .A(n_1490), .B(cacheD[60]), .Z(n_4224)
		);
	notech_and4 i_1431(.A(n_59537), .B(n_61513), .C(cacheQ[94]), .D(n_59468)
		, .Z(n_1985));
	notech_reg_set cacheD_reg_61(.CP(n_62031), .D(n_4230), .SD(1'b1), .Q(cacheD
		[61]));
	notech_mux2 i_3730(.S(n_59419), .A(n_1487), .B(cacheD[61]), .Z(n_4230)
		);
	notech_nao3 i_3122058(.A(n_2335), .B(n_2334), .C(n_1985), .Z(read_data[
		30]));
	notech_reg_set cacheD_reg_62(.CP(n_62047), .D(n_4236), .SD(1'b1), .Q(cacheD
		[62]));
	notech_mux2 i_3738(.S(n_59419), .A(n_1484), .B(cacheD[62]), .Z(n_4236)
		);
	notech_reg_set cacheD_reg_63(.CP(n_62047), .D(n_4242), .SD(1'b1), .Q(cacheD
		[63]));
	notech_mux2 i_3746(.S(n_59419), .A(n_1481), .B(cacheD[63]), .Z(n_4242)
		);
	notech_reg_set cacheD_reg_64(.CP(n_62047), .D(n_4248), .SD(1'b1), .Q(cacheD
		[64]));
	notech_mux2 i_3754(.S(n_1474), .A(n_1478), .B(cacheD[64]), .Z(n_4248));
	notech_reg_set cacheD_reg_65(.CP(n_62047), .D(n_4254), .SD(1'b1), .Q(cacheD
		[65]));
	notech_mux2 i_3762(.S(n_1474), .A(n_1472), .B(cacheD[65]), .Z(n_4254));
	notech_reg_set cacheD_reg_66(.CP(n_62047), .D(n_4260), .SD(1'b1), .Q(cacheD
		[66]));
	notech_mux2 i_3770(.S(n_1474), .A(n_1469), .B(cacheD[66]), .Z(n_4260));
	notech_and4 i_1440(.A(n_59537), .B(n_61513), .C(cacheQ[95]), .D(n_59468)
		, .Z(n_1991));
	notech_reg_set cacheD_reg_67(.CP(n_62047), .D(n_4266), .SD(1'b1), .Q(cacheD
		[67]));
	notech_mux2 i_3778(.S(n_1474), .A(n_1466), .B(cacheD[67]), .Z(n_4266));
	notech_nao3 i_3222059(.A(n_2338), .B(n_2337), .C(n_1991), .Z(read_data[
		31]));
	notech_reg_set cacheD_reg_68(.CP(n_62047), .D(n_4272), .SD(1'b1), .Q(cacheD
		[68]));
	notech_mux2 i_3786(.S(n_1474), .A(n_1463), .B(cacheD[68]), .Z(n_4272));
	notech_reg_set cacheD_reg_69(.CP(n_62047), .D(n_4278), .SD(1'b1), .Q(cacheD
		[69]));
	notech_mux2 i_3794(.S(n_1474), .A(n_1460), .B(cacheD[69]), .Z(n_4278));
	notech_nand2 i_49(.A(n_6765), .B(fsm[3]), .Z(n_1994));
	notech_reg_set cacheD_reg_70(.CP(n_62047), .D(n_4284), .SD(1'b1), .Q(cacheD
		[70]));
	notech_mux2 i_3802(.S(n_1474), .A(n_1457), .B(cacheD[70]), .Z(n_4284));
	notech_nao3 i_117(.A(fsm[1]), .B(fsm[3]), .C(fsm[0]), .Z(n_1995));
	notech_reg_set cacheD_reg_71(.CP(n_62047), .D(n_4290), .SD(1'b1), .Q(cacheD
		[71]));
	notech_mux2 i_3810(.S(n_1474), .A(n_1454), .B(cacheD[71]), .Z(n_4290));
	notech_nao3 i_1329957(.A(fsm[4]), .B(fsm[2]), .C(n_1995), .Z(n_1996));
	notech_reg_set cacheD_reg_72(.CP(n_62047), .D(n_4296), .SD(1'b1), .Q(cacheD
		[72]));
	notech_mux2 i_3818(.S(n_1474), .A(n_1451), .B(cacheD[72]), .Z(n_4296));
	notech_reg_set cacheD_reg_73(.CP(n_62047), .D(n_4302), .SD(1'b1), .Q(cacheD
		[73]));
	notech_mux2 i_3826(.S(n_1474), .A(n_1448), .B(cacheD[73]), .Z(n_4302));
	notech_nand3 i_68(.A(fsm[1]), .B(fsm[3]), .C(fsm[0]), .Z(n_1998));
	notech_reg_set cacheD_reg_74(.CP(n_62047), .D(n_4308), .SD(1'b1), .Q(cacheD
		[74]));
	notech_mux2 i_3834(.S(n_1474), .A(n_1445), .B(cacheD[74]), .Z(n_4308));
	notech_and2 i_48(.A(n_6767), .B(n_6766), .Z(n_1999));
	notech_reg_set cacheD_reg_75(.CP(n_62047), .D(n_4314), .SD(1'b1), .Q(cacheD
		[75]));
	notech_mux2 i_3842(.S(n_1474), .A(n_1442), .B(cacheD[75]), .Z(n_4314));
	notech_nao3 i_31(.A(n_6767), .B(n_6766), .C(fsm[4]), .Z(n_2000));
	notech_reg_set cacheD_reg_76(.CP(n_62047), .D(n_4320), .SD(1'b1), .Q(cacheD
		[76]));
	notech_mux2 i_3850(.S(n_1474), .A(n_1439), .B(cacheD[76]), .Z(n_4320));
	notech_reg_set cacheD_reg_77(.CP(n_62047), .D(n_4326), .SD(1'b1), .Q(cacheD
		[77]));
	notech_mux2 i_3858(.S(n_1474), .A(n_1436), .B(cacheD[77]), .Z(n_4326));
	notech_or4 i_113(.A(fsm[0]), .B(fsm[3]), .C(n_2000), .D(n_970), .Z(n_2002
		));
	notech_reg_set cacheD_reg_78(.CP(n_62047), .D(n_4332), .SD(1'b1), .Q(cacheD
		[78]));
	notech_mux2 i_3866(.S(n_1474), .A(n_1433), .B(cacheD[78]), .Z(n_4332));
	notech_and2 i_56059(.A(write_req), .B(n_7003), .Z(n_2003));
	notech_reg_set cacheD_reg_79(.CP(n_62047), .D(n_4338), .SD(1'b1), .Q(cacheD
		[79]));
	notech_mux2 i_3874(.S(n_1474), .A(n_1430), .B(cacheD[79]), .Z(n_4338));
	notech_ao3 i_14(.A(n_61513), .B(n_6763), .C(n_1742), .Z(n_2004));
	notech_reg_set cacheD_reg_80(.CP(n_62045), .D(n_4344), .SD(1'b1), .Q(cacheD
		[80]));
	notech_mux2 i_3882(.S(n_59441), .A(n_1427), .B(cacheD[80]), .Z(n_4344)
		);
	notech_reg_set cacheD_reg_81(.CP(n_62053), .D(n_4350), .SD(1'b1), .Q(cacheD
		[81]));
	notech_mux2 i_3890(.S(n_59441), .A(n_1424), .B(cacheD[81]), .Z(n_4350)
		);
	notech_reg_set cacheD_reg_82(.CP(n_62053), .D(n_4356), .SD(1'b1), .Q(cacheD
		[82]));
	notech_mux2 i_3898(.S(n_59441), .A(n_1421), .B(cacheD[82]), .Z(n_4356)
		);
	notech_or4 i_140(.A(code_wack), .B(n_971), .C(n_2003), .D(n_7006), .Z(n_2007
		));
	notech_reg_set cacheD_reg_83(.CP(n_62053), .D(n_4362), .SD(1'b1), .Q(cacheD
		[83]));
	notech_mux2 i_3906(.S(n_59441), .A(n_1418), .B(cacheD[83]), .Z(n_4362)
		);
	notech_or2 i_56170(.A(n_2002), .B(n_2007), .Z(n_2008));
	notech_reg_set cacheD_reg_84(.CP(n_62053), .D(n_4368), .SD(1'b1), .Q(cacheD
		[84]));
	notech_mux2 i_3914(.S(n_59441), .A(n_1415), .B(cacheD[84]), .Z(n_4368)
		);
	notech_reg_set cacheD_reg_85(.CP(n_62053), .D(n_4374), .SD(1'b1), .Q(cacheD
		[85]));
	notech_mux2 i_3922(.S(n_59441), .A(n_1412), .B(cacheD[85]), .Z(n_4374)
		);
	notech_or4 i_56157(.A(code_ack), .B(n_2003), .C(n_2002), .D(n_7004), .Z(n_2010
		));
	notech_reg_set cacheD_reg_86(.CP(n_62053), .D(n_4380), .SD(1'b1), .Q(cacheD
		[86]));
	notech_mux2 i_3930(.S(n_59441), .A(n_1409), .B(cacheD[86]), .Z(n_4380)
		);
	notech_reg_set cacheD_reg_87(.CP(n_62053), .D(n_4386), .SD(1'b1), .Q(cacheD
		[87]));
	notech_mux2 i_3938(.S(n_59441), .A(n_1406), .B(cacheD[87]), .Z(n_4386)
		);
	notech_reg_set cacheD_reg_88(.CP(n_62053), .D(n_4392), .SD(1'b1), .Q(cacheD
		[88]));
	notech_mux2 i_3946(.S(n_59441), .A(n_1403), .B(cacheD[88]), .Z(n_4392)
		);
	notech_reg_set cacheD_reg_89(.CP(n_62053), .D(n_4398), .SD(1'b1), .Q(cacheD
		[89]));
	notech_mux2 i_3954(.S(n_59441), .A(n_1400), .B(cacheD[89]), .Z(n_4398)
		);
	notech_reg_set cacheD_reg_90(.CP(n_62053), .D(n_4404), .SD(1'b1), .Q(cacheD
		[90]));
	notech_mux2 i_3962(.S(n_59441), .A(n_1397), .B(cacheD[90]), .Z(n_4404)
		);
	notech_reg_set cacheD_reg_91(.CP(n_62053), .D(n_4410), .SD(1'b1), .Q(cacheD
		[91]));
	notech_mux2 i_3970(.S(n_59441), .A(n_1394), .B(cacheD[91]), .Z(n_4410)
		);
	notech_and2 i_27(.A(axi_RVALID), .B(axi_RLAST), .Z(n_2016));
	notech_reg_set cacheD_reg_92(.CP(n_62053), .D(n_4416), .SD(1'b1), .Q(cacheD
		[92]));
	notech_mux2 i_3978(.S(n_59441), .A(n_1391), .B(cacheD[92]), .Z(n_4416)
		);
	notech_or2 i_116(.A(fsm[4]), .B(fsm[2]), .Z(n_2017));
	notech_reg_set cacheD_reg_93(.CP(n_62053), .D(n_4422), .SD(1'b1), .Q(cacheD
		[93]));
	notech_mux2 i_3986(.S(n_59441), .A(n_1388), .B(cacheD[93]), .Z(n_4422)
		);
	notech_reg_set cacheD_reg_94(.CP(n_62053), .D(n_4428), .SD(1'b1), .Q(cacheD
		[94]));
	notech_mux2 i_3994(.S(n_59441), .A(n_1385), .B(cacheD[94]), .Z(n_4428)
		);
	notech_or4 i_56132(.A(n_2017), .B(n_2003), .C(n_1998), .D(n_6657), .Z(n_2019
		));
	notech_reg_set cacheD_reg_95(.CP(n_62053), .D(n_4434), .SD(1'b1), .Q(cacheD
		[95]));
	notech_mux2 i_4002(.S(n_59441), .A(n_1382), .B(cacheD[95]), .Z(n_4434)
		);
	notech_ao3 i_52(.A(n_61513), .B(n_2019), .C(n_1742), .Z(n_2020));
	notech_reg_set cacheD_reg_96(.CP(n_62053), .D(n_4440), .SD(1'b1), .Q(cacheD
		[96]));
	notech_mux2 i_4010(.S(n_1375), .A(n_1379), .B(cacheD[96]), .Z(n_4440));
	notech_and2 i_12(.A(axi_AR[30]), .B(n_6999), .Z(n_2021));
	notech_reg_set cacheD_reg_97(.CP(n_62053), .D(n_4446), .SD(1'b1), .Q(cacheD
		[97]));
	notech_mux2 i_4018(.S(n_1375), .A(n_1373), .B(cacheD[97]), .Z(n_4446));
	notech_and2 i_110(.A(n_1066), .B(n_61496), .Z(n_2022));
	notech_reg_set cacheD_reg_98(.CP(n_62053), .D(n_4452), .SD(1'b1), .Q(cacheD
		[98]));
	notech_mux2 i_4026(.S(n_1375), .A(n_1370), .B(cacheD[98]), .Z(n_4452));
	notech_ao3 i_56137(.A(n_6765), .B(fsm[3]), .C(n_2000), .Z(n_2023));
	notech_reg_set cacheD_reg_99(.CP(n_62053), .D(n_4458), .SD(1'b1), .Q(cacheD
		[99]));
	notech_mux2 i_4034(.S(n_1375), .A(n_1367), .B(cacheD[99]), .Z(n_4458));
	notech_and2 i_33(.A(n_6705), .B(n_60826), .Z(n_2024));
	notech_reg_set cacheD_reg_100(.CP(n_62053), .D(n_4464), .SD(1'b1), .Q(cacheD
		[100]));
	notech_mux2 i_4042(.S(n_1375), .A(n_1364), .B(cacheD[100]), .Z(n_4464)
		);
	notech_nand2 i_13(.A(burst_idx[0]), .B(burst_idx[1]), .Z(n_2025));
	notech_reg_set cacheD_reg_101(.CP(n_62029), .D(n_4470), .SD(1'b1), .Q(cacheD
		[101]));
	notech_mux2 i_4050(.S(n_1375), .A(n_1361), .B(cacheD[101]), .Z(n_4470)
		);
	notech_nand3 i_42(.A(burst_idx[0]), .B(burst_idx[1]), .C(burst_idx[2]), 
		.Z(n_2026));
	notech_reg_set cacheD_reg_102(.CP(n_62029), .D(n_4476), .SD(1'b1), .Q(cacheD
		[102]));
	notech_mux2 i_4058(.S(n_1375), .A(n_1358), .B(cacheD[102]), .Z(n_4476)
		);
	notech_nao3 i_72(.A(burst_idx[2]), .B(burst_idx[3]), .C(n_2025), .Z(n_2027
		));
	notech_reg_set cacheD_reg_103(.CP(n_62029), .D(n_4482), .SD(1'b1), .Q(cacheD
		[103]));
	notech_mux2 i_4066(.S(n_1375), .A(n_1355), .B(cacheD[103]), .Z(n_4482)
		);
	notech_nor2 i_120(.A(burst_idx[0]), .B(n_6742), .Z(n_2028));
	notech_reg_set cacheD_reg_104(.CP(n_62029), .D(n_4488), .SD(1'b1), .Q(cacheD
		[104]));
	notech_mux2 i_4074(.S(n_1375), .A(n_1352), .B(cacheD[104]), .Z(n_4488)
		);
	notech_and2 i_124(.A(burst_idx[0]), .B(n_6742), .Z(n_2029));
	notech_reg_set cacheD_reg_105(.CP(n_62029), .D(n_4494), .SD(1'b1), .Q(cacheD
		[105]));
	notech_mux2 i_4082(.S(n_1375), .A(n_1349), .B(cacheD[105]), .Z(n_4494)
		);
	notech_nand2 i_53(.A(axi_RVALID), .B(n_61431), .Z(n_2030));
	notech_reg_set cacheD_reg_106(.CP(n_62029), .D(n_4500), .SD(1'b1), .Q(cacheD
		[106]));
	notech_mux2 i_4090(.S(n_1375), .A(n_1346), .B(cacheD[106]), .Z(n_4500)
		);
	notech_reg_set cacheD_reg_107(.CP(n_62029), .D(n_4506), .SD(1'b1), .Q(cacheD
		[107]));
	notech_mux2 i_4098(.S(n_1375), .A(n_1343), .B(cacheD[107]), .Z(n_4506)
		);
	notech_nand2 i_343(.A(n_6768), .B(fsm[0]), .Z(n_2032));
	notech_reg_set cacheD_reg_108(.CP(n_62029), .D(n_4512), .SD(1'b1), .Q(cacheD
		[108]));
	notech_mux2 i_4106(.S(n_1375), .A(n_1340), .B(cacheD[108]), .Z(n_4512)
		);
	notech_ao3 i_1129948(.A(n_6768), .B(fsm[0]), .C(n_2000), .Z(n_2033));
	notech_reg_set cacheD_reg_109(.CP(n_62029), .D(n_4518), .SD(1'b1), .Q(cacheD
		[109]));
	notech_mux2 i_4114(.S(n_1375), .A(n_1337), .B(cacheD[109]), .Z(n_4518)
		);
	notech_reg_set cacheD_reg_110(.CP(n_62029), .D(n_4524), .SD(1'b1), .Q(cacheD
		[110]));
	notech_mux2 i_4122(.S(n_1375), .A(n_1334), .B(cacheD[110]), .Z(n_4524)
		);
	notech_ao3 i_56(.A(n_6743), .B(n_6744), .C(burst_idx[4]), .Z(n_2035));
	notech_reg_set cacheD_reg_111(.CP(n_62029), .D(n_4530), .SD(1'b1), .Q(cacheD
		[111]));
	notech_mux2 i_4130(.S(n_1375), .A(n_1331), .B(cacheD[111]), .Z(n_4530)
		);
	notech_or2 i_114(.A(burst_idx[0]), .B(burst_idx[1]), .Z(n_2036));
	notech_reg_set cacheD_reg_112(.CP(n_62029), .D(n_4536), .SD(1'b1), .Q(cacheD
		[112]));
	notech_mux2 i_4138(.S(n_59546), .A(n_1328), .B(cacheD[112]), .Z(n_4536)
		);
	notech_ao3 i_5779562(.A(n_910), .B(n_909), .C(n_894), .Z(n_2037));
	notech_reg_set cacheD_reg_113(.CP(n_62029), .D(n_4542), .SD(1'b1), .Q(cacheD
		[113]));
	notech_mux2 i_4146(.S(n_59546), .A(n_1325), .B(cacheD[113]), .Z(n_4542)
		);
	notech_reg_set cacheD_reg_114(.CP(n_62029), .D(n_4548), .SD(1'b1), .Q(cacheD
		[114]));
	notech_mux2 i_4154(.S(n_59546), .A(n_1322), .B(cacheD[114]), .Z(n_4548)
		);
	notech_reg_set cacheD_reg_115(.CP(n_62029), .D(n_4554), .SD(1'b1), .Q(cacheD
		[115]));
	notech_mux2 i_4162(.S(n_59546), .A(n_1319), .B(cacheD[115]), .Z(n_4554)
		);
	notech_or4 i_347(.A(axi_AWVALID), .B(n_2036), .C(n_6660), .D(n_6997), .Z
		(n_2040));
	notech_reg_set cacheD_reg_116(.CP(n_62029), .D(n_4560), .SD(1'b1), .Q(cacheD
		[116]));
	notech_mux2 i_4170(.S(n_59546), .A(n_1316), .B(cacheD[116]), .Z(n_4560)
		);
	notech_or4 i_21(.A(burst_idx[2]), .B(burst_idx[3]), .C(burst_idx[4]), .D
		(n_2040), .Z(n_2041));
	notech_reg_set cacheD_reg_117(.CP(n_62029), .D(n_4566), .SD(1'b1), .Q(cacheD
		[117]));
	notech_mux2 i_4178(.S(n_59546), .A(n_1313), .B(cacheD[117]), .Z(n_4566)
		);
	notech_nor2 i_15(.A(n_25082), .B(n_60873), .Z(n_2042));
	notech_reg_set cacheD_reg_118(.CP(n_62029), .D(n_4572), .SD(1'b1), .Q(cacheD
		[118]));
	notech_mux2 i_4186(.S(n_59546), .A(n_1310), .B(cacheD[118]), .Z(n_4572)
		);
	notech_reg_set cacheD_reg_119(.CP(n_62029), .D(n_4578), .SD(1'b1), .Q(cacheD
		[119]));
	notech_mux2 i_4194(.S(n_59546), .A(n_1307), .B(cacheD[119]), .Z(n_4578)
		);
	notech_reg_set cacheD_reg_120(.CP(n_62049), .D(n_4584), .SD(1'b1), .Q(cacheD
		[120]));
	notech_mux2 i_4202(.S(n_59546), .A(n_1304), .B(cacheD[120]), .Z(n_4584)
		);
	notech_or4 i_56149(.A(fsm[4]), .B(fsm[1]), .C(n_1994), .D(n_6767), .Z(n_2045
		));
	notech_reg_set cacheD_reg_121(.CP(n_62011), .D(n_4590), .SD(1'b1), .Q(cacheD
		[121]));
	notech_mux2 i_4210(.S(n_59546), .A(n_1301), .B(cacheD[121]), .Z(n_4590)
		);
	notech_ao4 i_385(.A(code_req), .B(n_6705), .C(n_2045), .D(read_req), .Z(n_2046
		));
	notech_reg_set cacheD_reg_122(.CP(n_62011), .D(n_4596), .SD(1'b1), .Q(cacheD
		[122]));
	notech_mux2 i_4218(.S(n_59546), .A(n_1298), .B(cacheD[122]), .Z(n_4596)
		);
	notech_reg_set cacheD_reg_123(.CP(n_62011), .D(n_4602), .SD(1'b1), .Q(cacheD
		[123]));
	notech_mux2 i_4226(.S(n_59546), .A(n_1295), .B(cacheD[123]), .Z(n_4602)
		);
	notech_reg_set cacheD_reg_124(.CP(n_62011), .D(n_4608), .SD(1'b1), .Q(cacheD
		[124]));
	notech_mux2 i_4234(.S(n_59546), .A(n_1292), .B(cacheD[124]), .Z(n_4608)
		);
	notech_or4 i_47(.A(n_928), .B(n_944), .C(n_943), .D(n_6997), .Z(n_2049)
		);
	notech_reg_set cacheD_reg_125(.CP(n_62011), .D(n_4614), .SD(1'b1), .Q(cacheD
		[125]));
	notech_mux2 i_4242(.S(n_59546), .A(n_1289), .B(cacheD[125]), .Z(n_4614)
		);
	notech_nor2 i_125(.A(n_2019), .B(n_2021), .Z(n_2050));
	notech_reg_set cacheD_reg_126(.CP(n_62011), .D(n_4620), .SD(1'b1), .Q(cacheD
		[126]));
	notech_mux2 i_4250(.S(n_59546), .A(n_1286), .B(cacheD[126]), .Z(n_4620)
		);
	notech_ao4 i_46(.A(n_2049), .B(n_6656), .C(n_1995), .D(n_2017), .Z(n_2051
		));
	notech_reg_set cacheD_reg_127(.CP(n_62011), .D(n_4626), .SD(1'b1), .Q(cacheD
		[127]));
	notech_mux2 i_4258(.S(n_59546), .A(n_1283), .B(cacheD[127]), .Z(n_4626)
		);
	notech_and2 i_30(.A(axi_RREADY), .B(axi_RVALID), .Z(n_2052));
	notech_reg_set cacheD_reg_128(.CP(n_62011), .D(n_4632), .SD(1'b1), .Q(cacheD
		[128]));
	notech_mux2 i_4266(.S(n_1277), .A(n_6764), .B(cacheD[128]), .Z(n_4632)
		);
	notech_reg_set cacheD_reg_129(.CP(n_62011), .D(n_4638), .SD(1'b1), .Q(cacheD
		[129]));
	notech_mux2 i_4274(.S(n_1277), .A(n_6762), .B(cacheD[129]), .Z(n_4638)
		);
	notech_reg_set cacheD_reg_130(.CP(n_62011), .D(n_4644), .SD(1'b1), .Q(cacheD
		[130]));
	notech_mux2 i_4282(.S(n_1277), .A(n_6761), .B(cacheD[130]), .Z(n_4644)
		);
	notech_reg_set cacheD_reg_131(.CP(n_62011), .D(n_4650), .SD(1'b1), .Q(cacheD
		[131]));
	notech_mux2 i_4290(.S(n_1277), .A(n_6760), .B(cacheD[131]), .Z(n_4650)
		);
	notech_and2 i_57(.A(n_2045), .B(n_2042), .Z(n_2056));
	notech_reg_set cacheD_reg_132(.CP(n_62011), .D(n_4656), .SD(1'b1), .Q(cacheD
		[132]));
	notech_mux2 i_4298(.S(n_1277), .A(n_6759), .B(cacheD[132]), .Z(n_4656)
		);
	notech_and3 i_73(.A(n_2045), .B(n_2051), .C(n_2042), .Z(n_2057));
	notech_reg_set cacheD_reg_133(.CP(n_62011), .D(n_4662), .SD(1'b1), .Q(cacheD
		[133]));
	notech_mux2 i_4306(.S(n_1277), .A(n_6758), .B(cacheD[133]), .Z(n_4662)
		);
	notech_and2 i_119(.A(n_2057), .B(n_6705), .Z(n_2058));
	notech_reg_set cacheD_reg_134(.CP(n_62011), .D(n_4668), .SD(1'b1), .Q(cacheD
		[134]));
	notech_mux2 i_4314(.S(n_1277), .A(n_6757), .B(cacheD[134]), .Z(n_4668)
		);
	notech_reg_set cacheD_reg_135(.CP(n_62011), .D(n_4674), .SD(1'b1), .Q(cacheD
		[135]));
	notech_mux2 i_4322(.S(n_1277), .A(n_6756), .B(cacheD[135]), .Z(n_4674)
		);
	notech_reg_set cacheD_reg_136(.CP(n_62011), .D(n_4680), .SD(1'b1), .Q(cacheD
		[136]));
	notech_mux2 i_4330(.S(n_1277), .A(n_6755), .B(cacheD[136]), .Z(n_4680)
		);
	notech_and4 i_402(.A(n_2019), .B(n_1205), .C(n_1215), .D(n_6740), .Z(n_2061
		));
	notech_reg_set cacheD_reg_137(.CP(n_62011), .D(n_4686), .SD(1'b1), .Q(cacheD
		[137]));
	notech_mux2 i_4338(.S(n_1277), .A(n_6754), .B(cacheD[137]), .Z(n_4686)
		);
	notech_reg_set cacheD_reg_138(.CP(n_62049), .D(n_4692), .SD(1'b1), .Q(cacheD
		[138]));
	notech_mux2 i_4346(.S(n_1277), .A(n_6753), .B(cacheD[138]), .Z(n_4692)
		);
	notech_reg_set cacheD_reg_139(.CP(n_62033), .D(n_4698), .SD(1'b1), .Q(cacheD
		[139]));
	notech_mux2 i_4354(.S(n_59557), .A(n_6752), .B(cacheD[139]), .Z(n_4698)
		);
	notech_ao4 i_71(.A(n_2045), .B(n_6653), .C(n_2024), .D(n_6654), .Z(n_2064
		));
	notech_reg_set cacheD_reg_140(.CP(n_62049), .D(n_4704), .SD(1'b1), .Q(cacheD
		[140]));
	notech_mux2 i_4362(.S(n_59557), .A(n_6751), .B(cacheD[140]), .Z(n_4704)
		);
	notech_reg_set cacheD_reg_141(.CP(n_62049), .D(n_4710), .SD(1'b1), .Q(cacheD
		[141]));
	notech_mux2 i_4370(.S(n_59557), .A(n_6750), .B(cacheD[141]), .Z(n_4710)
		);
	notech_and4 i_415(.A(n_2019), .B(n_1205), .C(n_973), .D(n_6740), .Z(n_2066
		));
	notech_reg_set cacheD_reg_142(.CP(n_62049), .D(n_4716), .SD(1'b1), .Q(cacheD
		[142]));
	notech_mux2 i_4378(.S(n_59557), .A(n_6749), .B(cacheD[142]), .Z(n_4716)
		);
	notech_reg_set cacheD_reg_143(.CP(n_62049), .D(n_4722), .SD(1'b1), .Q(cacheD
		[143]));
	notech_mux2 i_4386(.S(n_59557), .A(n_6748), .B(cacheD[143]), .Z(n_4722)
		);
	notech_reg_set cacheD_reg_144(.CP(n_62049), .D(n_4728), .SD(1'b1), .Q(cacheD
		[144]));
	notech_mux2 i_4394(.S(n_59557), .A(n_6746), .B(cacheD[144]), .Z(n_4728)
		);
	notech_and2 i_0(.A(n_60873), .B(n_7002), .Z(n_2069));
	notech_reg_set cacheD_reg_145(.CP(n_62049), .D(n_4734), .SD(1'b1), .Q(cacheD
		[145]));
	notech_mux2 i_4402(.S(n_59557), .A(n_6745), .B(cacheD[145]), .Z(n_4734)
		);
	notech_and2 i_51(.A(n_61523), .B(n_1167), .Z(n_2070));
	notech_reg_set cacheD_reg_146(.CP(n_62049), .D(n_4740), .SD(1'b1), .Q(cacheD
		[146]));
	notech_mux2 i_4410(.S(n_1277), .A(n_23547), .B(cacheD[146]), .Z(n_4740)
		);
	notech_nand3 i_474(.A(axi_RVALID), .B(axi_RLAST), .C(n_61431), .Z(n_2071
		));
	notech_reg_set cacheD_reg_147(.CP(n_62049), .D(n_4746), .SD(1'b1), .Q(cacheD
		[147]));
	notech_mux2 i_4418(.S(n_59557), .A(n_23552), .B(cacheD[147]), .Z(n_4746)
		);
	notech_ao3 i_67(.A(n_60873), .B(n_59537), .C(n_21501), .Z(n_2072));
	notech_reg_set cacheD_reg_148(.CP(n_62049), .D(n_4752), .SD(1'b1), .Q(cacheD
		[148]));
	notech_mux2 i_4426(.S(n_59557), .A(n_1224), .B(cacheD[148]), .Z(n_4752)
		);
	notech_nand3 i_37(.A(n_59537), .B(n_2069), .C(n_59465), .Z(n_2073));
	notech_reg_set cacheD_reg_149(.CP(n_62049), .D(n_4758), .SD(1'b1), .Q(cacheD
		[149]));
	notech_mux2 i_4434(.S(n_59557), .A(n_23562), .B(cacheD[149]), .Z(n_4758)
		);
	notech_or4 i_65(.A(n_21501), .B(n_59537), .C(n_2032), .D(n_2000), .Z(n_2074
		));
	notech_reg axi_WSTRB_reg_0(.CP(n_62049), .D(n_4764), .CD(n_61430), .Q(axi_WSTRB
		[0]));
	notech_mux2 i_4442(.S(n_61480), .A(n_6772), .B(axi_WSTRB[0]), .Z(n_4764)
		);
	notech_nand3 i_35(.A(n_59537), .B(n_2069), .C(n_59503), .Z(n_2075));
	notech_reg axi_WSTRB_reg_1(.CP(n_62049), .D(n_4770), .CD(n_61430), .Q(axi_WSTRB
		[1]));
	notech_mux2 i_4450(.S(n_61480), .A(n_25361), .B(axi_WSTRB[1]), .Z(n_4770
		));
	notech_reg axi_WSTRB_reg_2(.CP(n_62049), .D(n_4776), .CD(n_61430), .Q(axi_WSTRB
		[2]));
	notech_mux2 i_4458(.S(n_61480), .A(n_25367), .B(axi_WSTRB[2]), .Z(n_4776
		));
	notech_reg axi_WSTRB_reg_3(.CP(n_62049), .D(n_4782), .CD(n_61430), .Q(axi_WSTRB
		[3]));
	notech_mux2 i_4466(.S(n_61480), .A(n_25373), .B(axi_WSTRB[3]), .Z(n_4782
		));
	notech_reg_set cacheM_reg_0(.CP(n_62049), .D(n_4788), .SD(n_61431), .Q(cacheM
		[0]));
	notech_mux2 i_4474(.S(n_1744), .A(n_1746), .B(cacheM[0]), .Z(n_4788));
	notech_reg_set cacheM_reg_1(.CP(n_62049), .D(n_4794), .SD(n_61431), .Q(cacheM
		[1]));
	notech_mux2 i_4482(.S(n_1744), .A(n_1741), .B(cacheM[1]), .Z(n_4794));
	notech_reg_set cacheM_reg_2(.CP(n_62049), .D(n_4800), .SD(n_61430), .Q(cacheM
		[2]));
	notech_mux2 i_4490(.S(n_1744), .A(n_1739), .B(cacheM[2]), .Z(n_4800));
	notech_reg_set cacheM_reg_3(.CP(n_62011), .D(n_4806), .SD(n_61431), .Q(cacheM
		[3]));
	notech_mux2 i_4498(.S(n_1744), .A(n_1737), .B(cacheM[3]), .Z(n_4806));
	notech_reg_set cacheM_reg_4(.CP(n_62011), .D(n_4812), .SD(n_61431), .Q(cacheM
		[4]));
	notech_mux2 i_4506(.S(n_1744), .A(n_1735), .B(cacheM[4]), .Z(n_4812));
	notech_reg_set cacheM_reg_5(.CP(n_62035), .D(n_4818), .SD(n_61432), .Q(cacheM
		[5]));
	notech_mux2 i_4514(.S(n_1744), .A(n_1733), .B(cacheM[5]), .Z(n_4818));
	notech_reg_set cacheM_reg_6(.CP(n_62035), .D(n_4824), .SD(n_61432), .Q(cacheM
		[6]));
	notech_mux2 i_4522(.S(n_1744), .A(n_1731), .B(cacheM[6]), .Z(n_4824));
	notech_reg_set cacheM_reg_7(.CP(n_62035), .D(n_4830), .SD(n_61432), .Q(cacheM
		[7]));
	notech_mux2 i_4530(.S(n_1744), .A(n_1729), .B(cacheM[7]), .Z(n_4830));
	notech_reg_set cacheM_reg_8(.CP(n_62035), .D(n_4836), .SD(n_61432), .Q(cacheM
		[8]));
	notech_mux2 i_4538(.S(n_1744), .A(n_1727), .B(cacheM[8]), .Z(n_4836));
	notech_reg_set cacheM_reg_9(.CP(n_62035), .D(n_4842), .SD(n_61432), .Q(cacheM
		[9]));
	notech_mux2 i_4546(.S(n_1744), .A(n_1725), .B(cacheM[9]), .Z(n_4842));
	notech_reg_set cacheM_reg_10(.CP(n_62035), .D(n_4848), .SD(n_61432), .Q(cacheM
		[10]));
	notech_mux2 i_4554(.S(n_1744), .A(n_1723), .B(cacheM[10]), .Z(n_4848));
	notech_reg_set cacheM_reg_11(.CP(n_62035), .D(n_4854), .SD(n_61432), .Q(cacheM
		[11]));
	notech_mux2 i_4562(.S(n_1744), .A(n_1721), .B(cacheM[11]), .Z(n_4854));
	notech_reg_set cacheM_reg_12(.CP(n_62035), .D(n_4860), .SD(n_61432), .Q(cacheM
		[12]));
	notech_mux2 i_4570(.S(n_1744), .A(n_1719), .B(cacheM[12]), .Z(n_4860));
	notech_reg_set cacheM_reg_13(.CP(n_62035), .D(n_4866), .SD(n_61432), .Q(cacheM
		[13]));
	notech_mux2 i_4578(.S(n_1744), .A(n_1717), .B(cacheM[13]), .Z(n_4866));
	notech_reg_set cacheM_reg_14(.CP(n_62035), .D(n_4872), .SD(n_61432), .Q(cacheM
		[14]));
	notech_mux2 i_4586(.S(n_1744), .A(n_1715), .B(cacheM[14]), .Z(n_4872));
	notech_reg_set cacheM_reg_15(.CP(n_62035), .D(n_4878), .SD(n_61431), .Q(cacheM
		[15]));
	notech_mux2 i_4594(.S(n_1744), .A(n_1713), .B(cacheM[15]), .Z(n_4878));
	notech_reg_set cacheWEN_reg(.CP(n_62035), .D(n_4884), .SD(n_61431), .Q(cacheWEN
		));
	notech_mux2 i_4602(.S(n_1749), .A(n_1751), .B(cacheWEN), .Z(n_4884));
	notech_reg axi_RREADY_reg(.CP(n_62035), .D(n_4890), .CD(n_61432), .Q(axi_RREADY
		));
	notech_mux2 i_4610(.S(n_1755), .A(n_1756), .B(axi_RREADY), .Z(n_4890));
	notech_reg axi_ARVALID_reg(.CP(n_62035), .D(n_4896), .CD(n_61432), .Q(axi_ARVALID
		));
	notech_mux2 i_4618(.S(n_1759), .A(n_1760), .B(axi_ARVALID), .Z(n_4896)
		);
	notech_reg axi_io_WVALID_reg(.CP(n_62035), .D(n_4902), .CD(n_61432), .Q(axi_io_WVALID
		));
	notech_mux2 i_4626(.S(n_1763), .A(n_23659), .B(axi_io_WVALID), .Z(n_4902
		));
	notech_reg wf_reg(.CP(n_62035), .D(writeio_req), .CD(n_61432), .Q(wf));
	notech_reg rf_reg(.CP(n_62035), .D(readio_req), .CD(n_61425), .Q(rf));
	notech_reg axi_io_ARVALID_reg(.CP(n_62035), .D(n_4912), .CD(n_61418), .Q
		(axi_io_ARVALID));
	notech_mux2 i_4642(.S(n_1765), .A(n_6770), .B(axi_io_ARVALID), .Z(n_4912
		));
	notech_reg axi_io_RREADY_reg(.CP(n_62013), .D(n_4918), .CD(n_61418), .Q(axi_io_RREADY
		));
	notech_mux2 i_4650(.S(n_1766), .A(n_23604), .B(axi_io_RREADY), .Z(n_4918
		));
	notech_reg readio_ack_reg(.CP(n_62035), .D(n_4926), .CD(n_61417), .Q(readio_ack
		));
	notech_ao3 i_4659(.A(n_222956060), .B(n_222856059), .C(readio_ack), .Z(n_4926
		));
	notech_reg writeio_ack_reg(.CP(n_61989), .D(n_4930), .CD(n_61417), .Q(writeio_ack
		));
	notech_xor2 i_4666(.A(n_7000), .B(n_1769), .Z(n_4930));
	notech_reg axi_io_AWVALID_reg(.CP(n_61989), .D(n_4936), .CD(n_61418), .Q
		(axi_io_AWVALID));
	notech_mux2 i_4674(.S(n_1770), .A(n_6773), .B(axi_io_AWVALID), .Z(n_4936
		));
	notech_reg axi_ARSIZE_reg_0(.CP(n_61989), .D(n_4945), .CD(n_61418), .Q(axi_ARSIZE
		[0]));
	notech_and2 i_4684(.A(n_61496), .B(axi_ARSIZE[0]), .Z(n_4945));
	notech_reg_set axi_ARSIZE_reg_1(.CP(n_61989), .D(n_4953), .SD(n_61418), 
		.Q(axi_ARSIZE[1]));
	notech_nao3 i_4695(.A(n_61496), .B(1'b1), .C(axi_ARSIZE[1]), .Z(n_4953)
		);
	notech_reg axi_ARSIZE_reg_2(.CP(n_61989), .D(n_4957), .CD(n_61418), .Q(axi_ARSIZE
		[2]));
	notech_and2 i_4700(.A(n_61496), .B(axi_ARSIZE[2]), .Z(n_4957));
	notech_reg axi_AWLEN_reg_0(.CP(n_61989), .D(n_4963), .CD(n_61417), .Q(axi_AWLEN
		[0]));
	notech_and4 i_4708(.A(n_61496), .B(n_6763), .C(n_61523), .D(axi_AWLEN[0]
		), .Z(n_4963));
	notech_and3 i_44(.A(axi_RVALID), .B(n_2035), .C(n_61417), .Z(n_210755938
		));
	notech_reg axi_AWLEN_reg_1(.CP(n_61989), .D(n_4969), .CD(n_61417), .Q(axi_AWLEN
		[1]));
	notech_and4 i_4716(.A(n_61496), .B(n_6763), .C(n_61523), .D(axi_AWLEN[1]
		), .Z(n_4969));
	notech_nao3 i_109(.A(n_2035), .B(n_60835), .C(n_2030), .Z(n_210855939)
		);
	notech_reg axi_AWLEN_reg_2(.CP(n_61989), .D(n_4975), .CD(n_61417), .Q(axi_AWLEN
		[2]));
	notech_and4 i_4724(.A(n_61496), .B(n_6763), .C(n_61523), .D(axi_AWLEN[2]
		), .Z(n_4975));
	notech_reg axi_AWLEN_reg_3(.CP(n_61989), .D(n_4981), .CD(n_61417), .Q(axi_AWLEN
		[3]));
	notech_and4 i_4732(.A(n_61491), .B(n_6763), .C(n_61523), .D(axi_AWLEN[3]
		), .Z(n_4981));
	notech_reg axi_AWLEN_reg_4(.CP(n_61989), .D(n_4987), .CD(n_61417), .Q(axi_AWLEN
		[4]));
	notech_and4 i_4740(.A(n_61491), .B(n_6763), .C(n_61523), .D(axi_AWLEN[4]
		), .Z(n_4987));
	notech_reg axi_AWLEN_reg_5(.CP(n_61989), .D(n_4993), .CD(n_61417), .Q(axi_AWLEN
		[5]));
	notech_and4 i_4748(.A(n_61491), .B(n_6763), .C(n_61523), .D(axi_AWLEN[5]
		), .Z(n_4993));
	notech_reg axi_AWLEN_reg_6(.CP(n_61989), .D(n_4999), .CD(n_61417), .Q(axi_AWLEN
		[6]));
	notech_and4 i_4756(.A(n_61491), .B(n_6763), .C(n_61523), .D(axi_AWLEN[6]
		), .Z(n_4999));
	notech_reg axi_AWLEN_reg_7(.CP(n_61989), .D(n_5005), .CD(n_61418), .Q(axi_AWLEN
		[7]));
	notech_and4 i_4764(.A(n_61491), .B(n_6763), .C(n_61523), .D(axi_AWLEN[7]
		), .Z(n_5005));
	notech_reg axi_WLAST_reg(.CP(n_61989), .D(n_5008), .CD(n_61419), .Q(axi_WLAST
		));
	notech_mux2 i_4770(.S(n_61480), .A(n_1176), .B(axi_WLAST), .Z(n_5008));
	notech_reg axi_ARLEN_reg_0(.CP(n_61989), .D(n_5014), .CD(n_61419), .Q(axi_ARLEN
		[0]));
	notech_mux2 i_4778(.S(n_60853), .A(n_6666), .B(axi_ARLEN[0]), .Z(n_5014)
		);
	notech_reg axi_ARLEN_reg_1(.CP(n_61989), .D(n_5020), .CD(n_61419), .Q(axi_ARLEN
		[1]));
	notech_mux2 i_4786(.S(n_60853), .A(n_6666), .B(axi_ARLEN[1]), .Z(n_5020)
		);
	notech_reg axi_ARLEN_reg_2(.CP(n_61989), .D(n_5029), .CD(n_61419), .Q(axi_ARLEN
		[2]));
	notech_and4 i_4796(.A(n_61491), .B(n_1066), .C(axi_ARLEN[2]), .D(n_973),
		 .Z(n_5029));
	notech_reg axi_ARLEN_reg_3(.CP(n_61989), .D(n_5035), .CD(n_61419), .Q(axi_ARLEN
		[3]));
	notech_and4 i_4804(.A(n_61491), .B(n_1066), .C(axi_ARLEN[3]), .D(n_973),
		 .Z(n_5035));
	notech_reg axi_ARLEN_reg_4(.CP(n_61989), .D(n_5041), .CD(n_61419), .Q(axi_ARLEN
		[4]));
	notech_and4 i_4812(.A(n_61491), .B(n_1066), .C(axi_ARLEN[4]), .D(n_973),
		 .Z(n_5041));
	notech_reg axi_ARLEN_reg_5(.CP(n_61997), .D(n_5047), .CD(n_61419), .Q(axi_ARLEN
		[5]));
	notech_and4 i_4820(.A(n_61491), .B(n_1066), .C(axi_ARLEN[5]), .D(n_973),
		 .Z(n_5047));
	notech_reg axi_ARLEN_reg_6(.CP(n_61981), .D(n_5053), .CD(n_61419), .Q(axi_ARLEN
		[6]));
	notech_and4 i_4828(.A(n_61491), .B(n_1066), .C(axi_ARLEN[6]), .D(n_973),
		 .Z(n_5053));
	notech_reg axi_ARLEN_reg_7(.CP(n_61981), .D(n_5059), .CD(n_61418), .Q(axi_ARLEN
		[7]));
	notech_and4 i_4836(.A(n_61491), .B(n_1066), .C(axi_ARLEN[7]), .D(n_973),
		 .Z(n_5059));
	notech_reg axi_io_AR_reg_0(.CP(n_61981), .D(n_5065), .CD(n_61418), .Q(axi_io_AR
		[0]));
	notech_and2 i_4844(.A(axi_io_AR[0]), .B(n_6771), .Z(n_5065));
	notech_reg axi_io_AR_reg_1(.CP(n_61981), .D(n_5071), .CD(n_61418), .Q(axi_io_AR
		[1]));
	notech_and2 i_4852(.A(n_6771), .B(axi_io_AR[1]), .Z(n_5071));
	notech_reg axi_io_AR_reg_2(.CP(n_61981), .D(n_5074), .CD(n_61418), .Q(axi_io_AR
		[2]));
	notech_mux2 i_4858(.S(\nbus_11673[0] ), .A(axi_io_AR[2]), .B(io_add[0]),
		 .Z(n_5074));
	notech_reg axi_io_AR_reg_3(.CP(n_61981), .D(n_5080), .CD(n_61418), .Q(axi_io_AR
		[3]));
	notech_mux2 i_4866(.S(\nbus_11673[0] ), .A(axi_io_AR[3]), .B(io_add[1]),
		 .Z(n_5080));
	notech_reg axi_io_AR_reg_4(.CP(n_61981), .D(n_5086), .CD(n_61418), .Q(axi_io_AR
		[4]));
	notech_mux2 i_4874(.S(\nbus_11673[0] ), .A(axi_io_AR[4]), .B(io_add[2]),
		 .Z(n_5086));
	notech_reg axi_io_AR_reg_5(.CP(n_61981), .D(n_5092), .CD(n_61418), .Q(axi_io_AR
		[5]));
	notech_mux2 i_4882(.S(\nbus_11673[0] ), .A(axi_io_AR[5]), .B(io_add[3]),
		 .Z(n_5092));
	notech_reg axi_io_AR_reg_6(.CP(n_61981), .D(n_5098), .CD(n_61418), .Q(axi_io_AR
		[6]));
	notech_mux2 i_4890(.S(\nbus_11673[0] ), .A(axi_io_AR[6]), .B(io_add[4]),
		 .Z(n_5098));
	notech_reg axi_io_AR_reg_7(.CP(n_61981), .D(n_5104), .CD(n_61417), .Q(axi_io_AR
		[7]));
	notech_mux2 i_4898(.S(\nbus_11673[0] ), .A(axi_io_AR[7]), .B(io_add[5]),
		 .Z(n_5104));
	notech_reg axi_io_AR_reg_8(.CP(n_61981), .D(n_5110), .CD(n_61415), .Q(axi_io_AR
		[8]));
	notech_mux2 i_4906(.S(\nbus_11673[0] ), .A(axi_io_AR[8]), .B(io_add[6]),
		 .Z(n_5110));
	notech_reg axi_io_AR_reg_9(.CP(n_61981), .D(n_5116), .CD(n_61415), .Q(axi_io_AR
		[9]));
	notech_mux2 i_4914(.S(\nbus_11673[0] ), .A(axi_io_AR[9]), .B(io_add[7]),
		 .Z(n_5116));
	notech_reg axi_io_AR_reg_10(.CP(n_61981), .D(n_5122), .CD(n_61415), .Q(axi_io_AR
		[10]));
	notech_mux2 i_4922(.S(\nbus_11673[0] ), .A(axi_io_AR[10]), .B(io_add[8])
		, .Z(n_5122));
	notech_reg axi_io_AR_reg_11(.CP(n_61981), .D(n_5128), .CD(n_61415), .Q(axi_io_AR
		[11]));
	notech_mux2 i_4930(.S(\nbus_11673[0] ), .A(axi_io_AR[11]), .B(io_add[9])
		, .Z(n_5128));
	notech_reg axi_io_AR_reg_12(.CP(n_61981), .D(n_5134), .CD(n_61416), .Q(axi_io_AR
		[12]));
	notech_mux2 i_4938(.S(\nbus_11673[0] ), .A(axi_io_AR[12]), .B(io_add[10]
		), .Z(n_5134));
	notech_reg axi_io_AR_reg_13(.CP(n_62001), .D(n_5140), .CD(n_61416), .Q(axi_io_AR
		[13]));
	notech_mux2 i_4946(.S(\nbus_11673[0] ), .A(axi_io_AR[13]), .B(io_add[11]
		), .Z(n_5140));
	notech_reg axi_io_AR_reg_14(.CP(n_62001), .D(n_5146), .CD(n_61415), .Q(axi_io_AR
		[14]));
	notech_mux2 i_4954(.S(\nbus_11673[0] ), .A(axi_io_AR[14]), .B(io_add[12]
		), .Z(n_5146));
	notech_reg axi_io_AR_reg_15(.CP(n_62001), .D(n_5152), .CD(n_61415), .Q(axi_io_AR
		[15]));
	notech_mux2 i_4962(.S(\nbus_11673[0] ), .A(axi_io_AR[15]), .B(io_add[13]
		), .Z(n_5152));
	notech_reg axi_io_AR_reg_16(.CP(n_62001), .D(n_5158), .CD(n_61415), .Q(axi_io_AR
		[16]));
	notech_mux2 i_4970(.S(\nbus_11673[0] ), .A(axi_io_AR[16]), .B(io_add[14]
		), .Z(n_5158));
	notech_reg axi_io_AR_reg_17(.CP(n_62001), .D(n_5164), .CD(n_61415), .Q(axi_io_AR
		[17]));
	notech_mux2 i_4978(.S(\nbus_11673[0] ), .A(axi_io_AR[17]), .B(io_add[15]
		), .Z(n_5164));
	notech_reg axi_io_AR_reg_18(.CP(n_62001), .D(n_5173), .CD(n_61415), .Q(axi_io_AR
		[18]));
	notech_and2 i_4988(.A(axi_io_AR[18]), .B(n_6771), .Z(n_5173));
	notech_ao3 i_36(.A(n_2069), .B(n_59468), .C(n_59537), .Z(n_214255973));
	notech_reg axi_io_AR_reg_19(.CP(n_62001), .D(n_5179), .CD(n_61415), .Q(axi_io_AR
		[19]));
	notech_and2 i_4996(.A(axi_io_AR[19]), .B(n_6771), .Z(n_5179));
	notech_ao3 i_34(.A(n_2069), .B(n_59503), .C(n_59537), .Z(n_214355974));
	notech_reg axi_io_AR_reg_20(.CP(n_62001), .D(n_5185), .CD(n_61415), .Q(axi_io_AR
		[20]));
	notech_and2 i_5004(.A(axi_io_AR[20]), .B(n_6771), .Z(n_5185));
	notech_reg axi_io_AR_reg_21(.CP(n_62001), .D(n_5191), .CD(n_61415), .Q(axi_io_AR
		[21]));
	notech_and2 i_5012(.A(axi_io_AR[21]), .B(n_6771), .Z(n_5191));
	notech_reg axi_io_AR_reg_22(.CP(n_62001), .D(n_5197), .CD(n_61415), .Q(axi_io_AR
		[22]));
	notech_and2 i_5020(.A(axi_io_AR[22]), .B(n_6771), .Z(n_5197));
	notech_reg axi_io_AR_reg_23(.CP(n_62001), .D(n_5203), .CD(n_61415), .Q(axi_io_AR
		[23]));
	notech_and2 i_5028(.A(axi_io_AR[23]), .B(n_6771), .Z(n_5203));
	notech_reg axi_io_AR_reg_24(.CP(n_62001), .D(n_5209), .CD(n_61416), .Q(axi_io_AR
		[24]));
	notech_and2 i_5036(.A(axi_io_AR[24]), .B(n_6771), .Z(n_5209));
	notech_reg axi_io_AR_reg_25(.CP(n_62001), .D(n_5215), .CD(n_61416), .Q(axi_io_AR
		[25]));
	notech_and2 i_5044(.A(axi_io_AR[25]), .B(n_6771), .Z(n_5215));
	notech_reg axi_io_AR_reg_26(.CP(n_62001), .D(n_5221), .CD(n_61416), .Q(axi_io_AR
		[26]));
	notech_and2 i_5052(.A(axi_io_AR[26]), .B(n_6771), .Z(n_5221));
	notech_reg axi_io_AR_reg_27(.CP(n_62001), .D(n_5227), .CD(n_61416), .Q(axi_io_AR
		[27]));
	notech_and2 i_5060(.A(axi_io_AR[27]), .B(n_6771), .Z(n_5227));
	notech_reg axi_io_AR_reg_28(.CP(n_62001), .D(n_5233), .CD(n_61416), .Q(axi_io_AR
		[28]));
	notech_and2 i_5068(.A(axi_io_AR[28]), .B(n_6771), .Z(n_5233));
	notech_reg axi_io_AR_reg_29(.CP(n_62001), .D(n_5239), .CD(n_61417), .Q(axi_io_AR
		[29]));
	notech_and2 i_5076(.A(axi_io_AR[29]), .B(n_6771), .Z(n_5239));
	notech_reg axi_io_AR_reg_30(.CP(n_62001), .D(n_5245), .CD(n_61417), .Q(axi_io_AR
		[30]));
	notech_and2 i_5084(.A(axi_io_AR[30]), .B(n_6771), .Z(n_5245));
	notech_reg axi_io_AR_reg_31(.CP(n_62001), .D(n_5251), .CD(n_61417), .Q(axi_io_AR
		[31]));
	notech_and2 i_5092(.A(axi_io_AR[31]), .B(n_6771), .Z(n_5251));
	notech_reg_set readio_data_reg_0(.CP(n_61999), .D(n_5254), .SD(1'b1), .Q
		(readio_data[0]));
	notech_mux2 i_5098(.S(\nbus_11671[0] ), .A(readio_data[0]), .B(axi_io_R[
		0]), .Z(n_5254));
	notech_reg_set readio_data_reg_1(.CP(n_61999), .D(n_5260), .SD(1'b1), .Q
		(readio_data[1]));
	notech_mux2 i_5106(.S(\nbus_11671[0] ), .A(readio_data[1]), .B(axi_io_R[
		1]), .Z(n_5260));
	notech_reg_set readio_data_reg_2(.CP(n_62025), .D(n_5266), .SD(1'b1), .Q
		(readio_data[2]));
	notech_mux2 i_5114(.S(\nbus_11671[0] ), .A(readio_data[2]), .B(axi_io_R[
		2]), .Z(n_5266));
	notech_reg_set readio_data_reg_3(.CP(n_62025), .D(n_5272), .SD(1'b1), .Q
		(readio_data[3]));
	notech_mux2 i_5122(.S(\nbus_11671[0] ), .A(readio_data[3]), .B(axi_io_R[
		3]), .Z(n_5272));
	notech_reg_set readio_data_reg_4(.CP(n_62025), .D(n_5278), .SD(1'b1), .Q
		(readio_data[4]));
	notech_mux2 i_5130(.S(\nbus_11671[0] ), .A(readio_data[4]), .B(axi_io_R[
		4]), .Z(n_5278));
	notech_reg_set readio_data_reg_5(.CP(n_62025), .D(n_5284), .SD(1'b1), .Q
		(readio_data[5]));
	notech_mux2 i_5138(.S(\nbus_11671[0] ), .A(readio_data[5]), .B(axi_io_R[
		5]), .Z(n_5284));
	notech_reg_set readio_data_reg_6(.CP(n_62025), .D(n_5290), .SD(1'b1), .Q
		(readio_data[6]));
	notech_mux2 i_5146(.S(\nbus_11671[0] ), .A(readio_data[6]), .B(axi_io_R[
		6]), .Z(n_5290));
	notech_reg_set readio_data_reg_7(.CP(n_62025), .D(n_5296), .SD(1'b1), .Q
		(readio_data[7]));
	notech_mux2 i_5154(.S(\nbus_11671[0] ), .A(readio_data[7]), .B(axi_io_R[
		7]), .Z(n_5296));
	notech_reg_set readio_data_reg_8(.CP(n_62025), .D(n_5302), .SD(1'b1), .Q
		(readio_data[8]));
	notech_mux2 i_5162(.S(\nbus_11671[0] ), .A(readio_data[8]), .B(axi_io_R[
		8]), .Z(n_5302));
	notech_reg_set readio_data_reg_9(.CP(n_62025), .D(n_5308), .SD(1'b1), .Q
		(readio_data[9]));
	notech_mux2 i_5170(.S(\nbus_11671[0] ), .A(readio_data[9]), .B(axi_io_R[
		9]), .Z(n_5308));
	notech_reg_set readio_data_reg_10(.CP(n_62025), .D(n_5314), .SD(1'b1), .Q
		(readio_data[10]));
	notech_mux2 i_5178(.S(\nbus_11671[0] ), .A(readio_data[10]), .B(axi_io_R
		[10]), .Z(n_5314));
	notech_reg_set readio_data_reg_11(.CP(n_62025), .D(n_5320), .SD(1'b1), .Q
		(readio_data[11]));
	notech_mux2 i_5186(.S(\nbus_11671[0] ), .A(readio_data[11]), .B(axi_io_R
		[11]), .Z(n_5320));
	notech_reg_set readio_data_reg_12(.CP(n_62025), .D(n_5326), .SD(1'b1), .Q
		(readio_data[12]));
	notech_mux2 i_5194(.S(\nbus_11671[0] ), .A(readio_data[12]), .B(axi_io_R
		[12]), .Z(n_5326));
	notech_reg_set readio_data_reg_13(.CP(n_62025), .D(n_5332), .SD(1'b1), .Q
		(readio_data[13]));
	notech_mux2 i_5202(.S(\nbus_11671[0] ), .A(readio_data[13]), .B(axi_io_R
		[13]), .Z(n_5332));
	notech_reg_set readio_data_reg_14(.CP(n_62025), .D(n_5338), .SD(1'b1), .Q
		(readio_data[14]));
	notech_mux2 i_5210(.S(\nbus_11671[0] ), .A(readio_data[14]), .B(axi_io_R
		[14]), .Z(n_5338));
	notech_reg_set readio_data_reg_15(.CP(n_62025), .D(n_5344), .SD(1'b1), .Q
		(readio_data[15]));
	notech_mux2 i_5218(.S(\nbus_11671[0] ), .A(readio_data[15]), .B(axi_io_R
		[15]), .Z(n_5344));
	notech_reg_set readio_data_reg_16(.CP(n_62025), .D(n_5350), .SD(1'b1), .Q
		(readio_data[16]));
	notech_mux2 i_5226(.S(n_53873), .A(readio_data[16]), .B(axi_io_R[16]), .Z
		(n_5350));
	notech_reg_set readio_data_reg_17(.CP(n_62025), .D(n_5356), .SD(1'b1), .Q
		(readio_data[17]));
	notech_mux2 i_5234(.S(n_53873), .A(readio_data[17]), .B(axi_io_R[17]), .Z
		(n_5356));
	notech_reg_set readio_data_reg_18(.CP(n_62025), .D(n_5362), .SD(1'b1), .Q
		(readio_data[18]));
	notech_mux2 i_5242(.S(n_53873), .A(readio_data[18]), .B(axi_io_R[18]), .Z
		(n_5362));
	notech_reg_set readio_data_reg_19(.CP(n_62025), .D(n_5368), .SD(1'b1), .Q
		(readio_data[19]));
	notech_mux2 i_5250(.S(n_53873), .A(readio_data[19]), .B(axi_io_R[19]), .Z
		(n_5368));
	notech_reg_set readio_data_reg_20(.CP(n_61999), .D(n_5374), .SD(1'b1), .Q
		(readio_data[20]));
	notech_mux2 i_5258(.S(n_53873), .A(readio_data[20]), .B(axi_io_R[20]), .Z
		(n_5374));
	notech_reg_set readio_data_reg_21(.CP(n_61999), .D(n_5380), .SD(1'b1), .Q
		(readio_data[21]));
	notech_mux2 i_5266(.S(n_53873), .A(readio_data[21]), .B(axi_io_R[21]), .Z
		(n_5380));
	notech_reg_set readio_data_reg_22(.CP(n_61999), .D(n_5386), .SD(1'b1), .Q
		(readio_data[22]));
	notech_mux2 i_5274(.S(n_53873), .A(readio_data[22]), .B(axi_io_R[22]), .Z
		(n_5386));
	notech_reg_set readio_data_reg_23(.CP(n_61999), .D(n_5392), .SD(1'b1), .Q
		(readio_data[23]));
	notech_mux2 i_5282(.S(n_53873), .A(readio_data[23]), .B(axi_io_R[23]), .Z
		(n_5392));
	notech_reg_set readio_data_reg_24(.CP(n_61999), .D(n_5398), .SD(1'b1), .Q
		(readio_data[24]));
	notech_mux2 i_5290(.S(n_53873), .A(readio_data[24]), .B(axi_io_R[24]), .Z
		(n_5398));
	notech_reg_set readio_data_reg_25(.CP(n_61999), .D(n_5404), .SD(1'b1), .Q
		(readio_data[25]));
	notech_mux2 i_5298(.S(n_53873), .A(readio_data[25]), .B(axi_io_R[25]), .Z
		(n_5404));
	notech_reg_set readio_data_reg_26(.CP(n_61999), .D(n_5410), .SD(1'b1), .Q
		(readio_data[26]));
	notech_mux2 i_5306(.S(n_53873), .A(readio_data[26]), .B(axi_io_R[26]), .Z
		(n_5410));
	notech_reg_set readio_data_reg_27(.CP(n_61999), .D(n_5416), .SD(1'b1), .Q
		(readio_data[27]));
	notech_mux2 i_5314(.S(n_53873), .A(readio_data[27]), .B(axi_io_R[27]), .Z
		(n_5416));
	notech_reg_set readio_data_reg_28(.CP(n_61999), .D(n_5422), .SD(1'b1), .Q
		(readio_data[28]));
	notech_mux2 i_5322(.S(n_53873), .A(readio_data[28]), .B(axi_io_R[28]), .Z
		(n_5422));
	notech_reg_set readio_data_reg_29(.CP(n_61999), .D(n_5428), .SD(1'b1), .Q
		(readio_data[29]));
	notech_mux2 i_5330(.S(n_53873), .A(readio_data[29]), .B(axi_io_R[29]), .Z
		(n_5428));
	notech_reg_set readio_data_reg_30(.CP(n_61999), .D(n_5434), .SD(1'b1), .Q
		(readio_data[30]));
	notech_mux2 i_5338(.S(n_53873), .A(readio_data[30]), .B(axi_io_R[30]), .Z
		(n_5434));
	notech_reg_set readio_data_reg_31(.CP(n_61999), .D(n_5440), .SD(1'b1), .Q
		(readio_data[31]));
	notech_mux2 i_5346(.S(n_53873), .A(readio_data[31]), .B(axi_io_R[31]), .Z
		(n_5440));
	notech_reg axi_AWSIZE_reg_0(.CP(n_61999), .D(n_5449), .CD(n_61417), .Q(axi_AWSIZE
		[0]));
	notech_and2 i_5356(.A(n_61496), .B(axi_AWSIZE[0]), .Z(n_5449));
	notech_reg_set axi_AWSIZE_reg_1(.CP(n_61999), .D(n_5457), .SD(n_61416), 
		.Q(axi_AWSIZE[1]));
	notech_nao3 i_5367(.A(n_61491), .B(1'b1), .C(axi_AWSIZE[1]), .Z(n_5457)
		);
	notech_reg axi_AWSIZE_reg_2(.CP(n_61999), .D(n_5461), .CD(n_61416), .Q(axi_AWSIZE
		[2]));
	notech_and2 i_5372(.A(n_61491), .B(axi_AWSIZE[2]), .Z(n_5461));
	notech_reg_set axi_AWBURST_reg_0(.CP(n_62025), .D(n_5469), .SD(n_61416),
		 .Q(axi_AWBURST[0]));
	notech_nao3 i_5383(.A(n_61491), .B(1'b1), .C(axi_AWBURST[0]), .Z(n_5469)
		);
	notech_reg axi_AWBURST_reg_1(.CP(n_62021), .D(n_5473), .CD(n_61416), .Q(axi_AWBURST
		[1]));
	notech_and2 i_5388(.A(n_61491), .B(axi_AWBURST[1]), .Z(n_5473));
	notech_reg_set code_data_reg_0(.CP(n_61997), .D(n_5476), .SD(1'b1), .Q(\nbus_14528[0] 
		));
	notech_mux2 i_5394(.S(\nbus_11667[0] ), .A(n_60429), .B(axi_R[0]), .Z(n_5476
		));
	notech_reg_set code_data_reg_1(.CP(n_62021), .D(n_5482), .SD(1'b1), .Q(code_data
		[1]));
	notech_mux2 i_5402(.S(\nbus_11667[0] ), .A(code_data[1]), .B(axi_R[1]), 
		.Z(n_5482));
	notech_reg_set code_data_reg_2(.CP(n_62021), .D(n_5488), .SD(1'b1), .Q(code_data
		[2]));
	notech_mux2 i_5410(.S(\nbus_11667[0] ), .A(code_data[2]), .B(axi_R[2]), 
		.Z(n_5488));
	notech_reg_set code_data_reg_3(.CP(n_62021), .D(n_5494), .SD(1'b1), .Q(code_data
		[3]));
	notech_mux2 i_5418(.S(\nbus_11667[0] ), .A(code_data[3]), .B(axi_R[3]), 
		.Z(n_5494));
	notech_reg_set code_data_reg_4(.CP(n_62021), .D(n_5500), .SD(1'b1), .Q(code_data
		[4]));
	notech_mux2 i_5426(.S(\nbus_11667[0] ), .A(code_data[4]), .B(axi_R[4]), 
		.Z(n_5500));
	notech_reg_set code_data_reg_5(.CP(n_62021), .D(n_5506), .SD(1'b1), .Q(code_data
		[5]));
	notech_mux2 i_5434(.S(\nbus_11667[0] ), .A(code_data[5]), .B(axi_R[5]), 
		.Z(n_5506));
	notech_reg_set code_data_reg_6(.CP(n_62021), .D(n_5512), .SD(1'b1), .Q(code_data
		[6]));
	notech_mux2 i_5442(.S(\nbus_11667[0] ), .A(code_data[6]), .B(axi_R[6]), 
		.Z(n_5512));
	notech_reg_set code_data_reg_7(.CP(n_62021), .D(n_5518), .SD(1'b1), .Q(code_data
		[7]));
	notech_mux2 i_5450(.S(\nbus_11667[0] ), .A(code_data[7]), .B(axi_R[7]), 
		.Z(n_5518));
	notech_reg_set code_data_reg_8(.CP(n_62021), .D(n_5524), .SD(1'b1), .Q(code_data
		[8]));
	notech_mux2 i_5458(.S(\nbus_11667[0] ), .A(code_data[8]), .B(axi_R[8]), 
		.Z(n_5524));
	notech_reg_set code_data_reg_9(.CP(n_62021), .D(n_5530), .SD(1'b1), .Q(code_data
		[9]));
	notech_mux2 i_5466(.S(\nbus_11667[0] ), .A(code_data[9]), .B(axi_R[9]), 
		.Z(n_5530));
	notech_reg_set code_data_reg_10(.CP(n_62021), .D(n_5536), .SD(1'b1), .Q(code_data
		[10]));
	notech_mux2 i_5474(.S(\nbus_11667[0] ), .A(code_data[10]), .B(axi_R[10])
		, .Z(n_5536));
	notech_reg_set code_data_reg_11(.CP(n_62021), .D(n_5542), .SD(1'b1), .Q(code_data
		[11]));
	notech_mux2 i_5482(.S(\nbus_11667[0] ), .A(code_data[11]), .B(axi_R[11])
		, .Z(n_5542));
	notech_reg_set code_data_reg_12(.CP(n_62021), .D(n_5548), .SD(1'b1), .Q(code_data
		[12]));
	notech_mux2 i_5490(.S(\nbus_11667[0] ), .A(code_data[12]), .B(axi_R[12])
		, .Z(n_5548));
	notech_reg_set code_data_reg_13(.CP(n_62021), .D(n_5554), .SD(1'b1), .Q(code_data
		[13]));
	notech_mux2 i_5498(.S(\nbus_11667[0] ), .A(code_data[13]), .B(axi_R[13])
		, .Z(n_5554));
	notech_reg_set code_data_reg_14(.CP(n_62021), .D(n_5560), .SD(1'b1), .Q(code_data
		[14]));
	notech_mux2 i_5506(.S(\nbus_11667[0] ), .A(code_data[14]), .B(axi_R[14])
		, .Z(n_5560));
	notech_reg_set code_data_reg_15(.CP(n_62021), .D(n_5566), .SD(1'b1), .Q(code_data
		[15]));
	notech_mux2 i_5514(.S(\nbus_11667[0] ), .A(code_data[15]), .B(axi_R[15])
		, .Z(n_5566));
	notech_reg_set code_data_reg_16(.CP(n_62043), .D(n_5572), .SD(1'b1), .Q(code_data
		[16]));
	notech_mux2 i_5522(.S(n_56598), .A(code_data[16]), .B(axi_R[16]), .Z(n_5572
		));
	notech_ao3 i_1013(.A(n_2019), .B(n_1711), .C(n_1742), .Z(n_220956040));
	notech_reg_set code_data_reg_17(.CP(n_62043), .D(n_5578), .SD(1'b1), .Q(code_data
		[17]));
	notech_mux2 i_5530(.S(n_56598), .A(code_data[17]), .B(axi_R[17]), .Z(n_5578
		));
	notech_reg_set code_data_reg_18(.CP(n_62043), .D(n_5584), .SD(1'b1), .Q(code_data
		[18]));
	notech_mux2 i_5538(.S(n_56598), .A(code_data[18]), .B(axi_R[18]), .Z(n_5584
		));
	notech_reg_set code_data_reg_19(.CP(n_62043), .D(n_5590), .SD(1'b1), .Q(code_data
		[19]));
	notech_mux2 i_5546(.S(n_56598), .A(code_data[19]), .B(axi_R[19]), .Z(n_5590
		));
	notech_reg_set code_data_reg_20(.CP(n_62043), .D(n_5596), .SD(1'b1), .Q(code_data
		[20]));
	notech_mux2 i_5554(.S(n_56598), .A(code_data[20]), .B(axi_R[20]), .Z(n_5596
		));
	notech_reg_set code_data_reg_21(.CP(n_62043), .D(n_5602), .SD(1'b1), .Q(code_data
		[21]));
	notech_mux2 i_5562(.S(n_56598), .A(code_data[21]), .B(axi_R[21]), .Z(n_5602
		));
	notech_reg_set code_data_reg_22(.CP(n_62043), .D(n_5608), .SD(1'b1), .Q(code_data
		[22]));
	notech_mux2 i_5570(.S(n_56598), .A(code_data[22]), .B(axi_R[22]), .Z(n_5608
		));
	notech_reg_set code_data_reg_23(.CP(n_62043), .D(n_5614), .SD(1'b1), .Q(code_data
		[23]));
	notech_mux2 i_5578(.S(n_56598), .A(code_data[23]), .B(axi_R[23]), .Z(n_5614
		));
	notech_or4 i_1058(.A(n_1221), .B(n_974), .C(n_1748), .D(n_2033), .Z(n_221656047
		));
	notech_reg_set code_data_reg_24(.CP(n_62043), .D(n_5620), .SD(1'b1), .Q(code_data
		[24]));
	notech_mux2 i_5586(.S(n_56598), .A(code_data[24]), .B(axi_R[24]), .Z(n_5620
		));
	notech_reg_set code_data_reg_25(.CP(n_62043), .D(n_5626), .SD(1'b1), .Q(code_data
		[25]));
	notech_mux2 i_5594(.S(n_56598), .A(code_data[25]), .B(axi_R[25]), .Z(n_5626
		));
	notech_reg_set code_data_reg_26(.CP(n_62043), .D(n_5632), .SD(1'b1), .Q(code_data
		[26]));
	notech_mux2 i_5602(.S(n_56598), .A(code_data[26]), .B(axi_R[26]), .Z(n_5632
		));
	notech_ao4 i_58(.A(n_2045), .B(n_2052), .C(n_60826), .D(n_2016), .Z(n_221956050
		));
	notech_reg_set code_data_reg_27(.CP(n_62043), .D(n_5638), .SD(1'b1), .Q(code_data
		[27]));
	notech_mux2 i_5610(.S(n_56598), .A(code_data[27]), .B(axi_R[27]), .Z(n_5638
		));
	notech_reg_set code_data_reg_28(.CP(n_62043), .D(n_5644), .SD(1'b1), .Q(code_data
		[28]));
	notech_mux2 i_5618(.S(n_56598), .A(code_data[28]), .B(axi_R[28]), .Z(n_5644
		));
	notech_reg_set code_data_reg_29(.CP(n_62043), .D(n_5650), .SD(1'b1), .Q(code_data
		[29]));
	notech_mux2 i_5626(.S(n_56598), .A(code_data[29]), .B(axi_R[29]), .Z(n_5650
		));
	notech_reg_set code_data_reg_30(.CP(n_62043), .D(n_5656), .SD(1'b1), .Q(code_data
		[30]));
	notech_mux2 i_5634(.S(n_56598), .A(code_data[30]), .B(axi_R[30]), .Z(n_5656
		));
	notech_reg_set code_data_reg_31(.CP(n_62043), .D(n_5662), .SD(1'b1), .Q(code_data
		[31]));
	notech_mux2 i_5642(.S(n_56598), .A(code_data[31]), .B(axi_R[31]), .Z(n_5662
		));
	notech_or2 i_55(.A(readio_ack), .B(writeio_ack), .Z(n_222456055));
	notech_reg_set code_data_reg_32(.CP(n_62043), .D(n_5668), .SD(1'b1), .Q(code_data
		[32]));
	notech_mux2 i_5650(.S(\nbus_11667[32] ), .A(code_data[32]), .B(axi_R[0])
		, .Z(n_5668));
	notech_nao3 i_118(.A(n_7000), .B(n_6773), .C(readio_ack), .Z(n_222556056
		));
	notech_reg_set code_data_reg_33(.CP(n_62043), .D(n_5674), .SD(1'b1), .Q(code_data
		[33]));
	notech_mux2 i_5658(.S(\nbus_11667[32] ), .A(code_data[33]), .B(axi_R[1])
		, .Z(n_5674));
	notech_nand2 i_122(.A(axi_io_WVALID), .B(axi_io_WREADY), .Z(n_222656057)
		);
	notech_reg_set code_data_reg_34(.CP(n_62021), .D(n_5680), .SD(1'b1), .Q(code_data
		[34]));
	notech_mux2 i_5666(.S(\nbus_11667[32] ), .A(code_data[34]), .B(axi_R[2])
		, .Z(n_5680));
	notech_nao3 i_54(.A(n_222656057), .B(n_6773), .C(n_222456055), .Z(n_222756058
		));
	notech_reg_set code_data_reg_35(.CP(n_62043), .D(n_5686), .SD(1'b1), .Q(code_data
		[35]));
	notech_mux2 i_5674(.S(\nbus_11667[32] ), .A(code_data[35]), .B(axi_R[3])
		, .Z(n_5686));
	notech_ao3 i_63(.A(n_222656057), .B(n_6770), .C(n_222556056), .Z(n_222856059
		));
	notech_reg_set code_data_reg_36(.CP(n_62023), .D(n_5692), .SD(1'b1), .Q(code_data
		[36]));
	notech_mux2 i_5682(.S(\nbus_11667[32] ), .A(code_data[36]), .B(axi_R[4])
		, .Z(n_5692));
	notech_and2 i_75(.A(axi_io_RREADY), .B(axi_io_RVALID), .Z(n_222956060)
		);
	notech_reg_set code_data_reg_37(.CP(n_62023), .D(n_5698), .SD(1'b1), .Q(code_data
		[37]));
	notech_mux2 i_5690(.S(\nbus_11667[32] ), .A(code_data[37]), .B(axi_R[5])
		, .Z(n_5698));
	notech_nao3 i_66(.A(n_6770), .B(n_6659), .C(n_222756058), .Z(n_223056061
		));
	notech_reg_set code_data_reg_38(.CP(n_62023), .D(n_5704), .SD(1'b1), .Q(code_data
		[38]));
	notech_mux2 i_5698(.S(\nbus_11667[32] ), .A(code_data[38]), .B(axi_R[6])
		, .Z(n_5704));
	notech_nand2 i_23(.A(writeio_req), .B(n_6769), .Z(n_223156062));
	notech_reg_set code_data_reg_39(.CP(n_62023), .D(n_5710), .SD(1'b1), .Q(code_data
		[39]));
	notech_mux2 i_5706(.S(\nbus_11667[32] ), .A(code_data[39]), .B(axi_R[7])
		, .Z(n_5710));
	notech_reg_set code_data_reg_40(.CP(n_62023), .D(n_5716), .SD(1'b1), .Q(code_data
		[40]));
	notech_mux2 i_5714(.S(\nbus_11667[32] ), .A(code_data[40]), .B(axi_R[8])
		, .Z(n_5716));
	notech_nao3 i_1112(.A(readio_req), .B(n_223156062), .C(rf), .Z(n_223356064
		));
	notech_reg_set code_data_reg_41(.CP(n_62023), .D(n_5722), .SD(1'b1), .Q(code_data
		[41]));
	notech_mux2 i_5722(.S(\nbus_11667[32] ), .A(code_data[41]), .B(axi_R[9])
		, .Z(n_5722));
	notech_reg_set code_data_reg_42(.CP(n_62023), .D(n_5728), .SD(1'b1), .Q(code_data
		[42]));
	notech_mux2 i_5730(.S(\nbus_11667[32] ), .A(code_data[42]), .B(axi_R[10]
		), .Z(n_5728));
	notech_reg_set code_data_reg_43(.CP(n_62023), .D(n_5734), .SD(1'b1), .Q(code_data
		[43]));
	notech_mux2 i_5738(.S(\nbus_11667[32] ), .A(code_data[43]), .B(axi_R[11]
		), .Z(n_5734));
	notech_reg_set code_data_reg_44(.CP(n_62023), .D(n_5740), .SD(1'b1), .Q(code_data
		[44]));
	notech_mux2 i_5746(.S(\nbus_11667[32] ), .A(code_data[44]), .B(axi_R[12]
		), .Z(n_5740));
	notech_nand3 i_40(.A(n_59537), .B(n_61502), .C(n_59503), .Z(n_2237));
	notech_reg_set code_data_reg_45(.CP(n_62023), .D(n_5746), .SD(1'b1), .Q(code_data
		[45]));
	notech_mux2 i_5754(.S(\nbus_11667[32] ), .A(code_data[45]), .B(axi_R[13]
		), .Z(n_5746));
	notech_reg_set code_data_reg_46(.CP(n_62023), .D(n_5752), .SD(1'b1), .Q(code_data
		[46]));
	notech_mux2 i_5762(.S(\nbus_11667[32] ), .A(code_data[46]), .B(axi_R[14]
		), .Z(n_5752));
	notech_nao3 i_41(.A(n_61502), .B(n_59503), .C(n_59537), .Z(n_2239));
	notech_reg_set code_data_reg_47(.CP(n_62023), .D(n_5758), .SD(1'b1), .Q(code_data
		[47]));
	notech_mux2 i_5770(.S(\nbus_11667[32] ), .A(code_data[47]), .B(axi_R[15]
		), .Z(n_5758));
	notech_ao4 i_1164(.A(n_2239), .B(n_6915), .C(n_2237), .D(n_6947), .Z(n_2240
		));
	notech_reg_set code_data_reg_48(.CP(n_62023), .D(n_5764), .SD(1'b1), .Q(code_data
		[48]));
	notech_mux2 i_5778(.S(n_53672), .A(code_data[48]), .B(axi_R[16]), .Z(n_5764
		));
	notech_reg_set code_data_reg_49(.CP(n_62023), .D(n_5770), .SD(1'b1), .Q(code_data
		[49]));
	notech_mux2 i_5786(.S(n_53672), .A(code_data[49]), .B(axi_R[17]), .Z(n_5770
		));
	notech_reg_set code_data_reg_50(.CP(n_62023), .D(n_5776), .SD(1'b1), .Q(code_data
		[50]));
	notech_mux2 i_5794(.S(n_53672), .A(code_data[50]), .B(axi_R[18]), .Z(n_5776
		));
	notech_reg_set code_data_reg_51(.CP(n_62023), .D(n_5782), .SD(1'b1), .Q(code_data
		[51]));
	notech_mux2 i_5802(.S(n_53672), .A(code_data[51]), .B(axi_R[19]), .Z(n_5782
		));
	notech_nao3 i_38(.A(n_61502), .B(n_59468), .C(n_59537), .Z(n_2244));
	notech_reg_set code_data_reg_52(.CP(n_62023), .D(n_5788), .SD(1'b1), .Q(code_data
		[52]));
	notech_mux2 i_5810(.S(n_53672), .A(code_data[52]), .B(axi_R[20]), .Z(n_5788
		));
	notech_ao4 i_1163(.A(n_61502), .B(n_6775), .C(n_2244), .D(n_6883), .Z(n_2245
		));
	notech_reg_set code_data_reg_53(.CP(n_62023), .D(n_5794), .SD(1'b1), .Q(code_data
		[53]));
	notech_mux2 i_5818(.S(n_53672), .A(code_data[53]), .B(axi_R[21]), .Z(n_5794
		));
	notech_reg_set code_data_reg_54(.CP(n_62023), .D(n_5800), .SD(1'b1), .Q(code_data
		[54]));
	notech_mux2 i_5826(.S(n_53672), .A(code_data[54]), .B(axi_R[22]), .Z(n_5800
		));
	notech_ao4 i_1173(.A(n_2239), .B(n_6916), .C(n_2237), .D(n_6948), .Z(n_2247
		));
	notech_reg_set code_data_reg_55(.CP(n_61997), .D(n_5806), .SD(1'b1), .Q(code_data
		[55]));
	notech_mux2 i_5834(.S(n_53672), .A(code_data[55]), .B(axi_R[23]), .Z(n_5806
		));
	notech_ao4 i_1172(.A(n_61502), .B(n_6776), .C(n_2244), .D(n_6884), .Z(n_2248
		));
	notech_reg_set code_data_reg_56(.CP(n_61997), .D(n_5812), .SD(1'b1), .Q(code_data
		[56]));
	notech_mux2 i_5842(.S(n_53672), .A(code_data[56]), .B(axi_R[24]), .Z(n_5812
		));
	notech_reg_set code_data_reg_57(.CP(n_61997), .D(n_5818), .SD(1'b1), .Q(code_data
		[57]));
	notech_mux2 i_5850(.S(n_53672), .A(code_data[57]), .B(axi_R[25]), .Z(n_5818
		));
	notech_ao4 i_1182(.A(n_2239), .B(n_6917), .C(n_2237), .D(n_6949), .Z(n_2250
		));
	notech_reg_set code_data_reg_58(.CP(n_61997), .D(n_5824), .SD(1'b1), .Q(code_data
		[58]));
	notech_mux2 i_5858(.S(n_53672), .A(code_data[58]), .B(axi_R[26]), .Z(n_5824
		));
	notech_ao4 i_1181(.A(n_61507), .B(n_6777), .C(n_2244), .D(n_6885), .Z(n_2251
		));
	notech_reg_set code_data_reg_59(.CP(n_61997), .D(n_5830), .SD(1'b1), .Q(code_data
		[59]));
	notech_mux2 i_5866(.S(n_53672), .A(code_data[59]), .B(axi_R[27]), .Z(n_5830
		));
	notech_reg_set code_data_reg_60(.CP(n_61997), .D(n_5836), .SD(1'b1), .Q(code_data
		[60]));
	notech_mux2 i_5874(.S(n_53672), .A(code_data[60]), .B(axi_R[28]), .Z(n_5836
		));
	notech_ao4 i_1191(.A(n_2239), .B(n_6918), .C(n_2237), .D(n_6950), .Z(n_2253
		));
	notech_reg_set code_data_reg_61(.CP(n_61981), .D(n_5842), .SD(1'b1), .Q(code_data
		[61]));
	notech_mux2 i_5882(.S(n_53672), .A(code_data[61]), .B(axi_R[29]), .Z(n_5842
		));
	notech_ao4 i_1190(.A(n_61502), .B(n_6778), .C(n_2244), .D(n_6886), .Z(n_2254
		));
	notech_reg_set code_data_reg_62(.CP(n_61997), .D(n_5848), .SD(1'b1), .Q(code_data
		[62]));
	notech_mux2 i_5890(.S(n_53672), .A(code_data[62]), .B(axi_R[30]), .Z(n_5848
		));
	notech_reg_set code_data_reg_63(.CP(n_61997), .D(n_5854), .SD(1'b1), .Q(code_data
		[63]));
	notech_mux2 i_5898(.S(n_53672), .A(code_data[63]), .B(axi_R[31]), .Z(n_5854
		));
	notech_ao4 i_1200(.A(n_2239), .B(n_6919), .C(n_2237), .D(n_6951), .Z(n_2256
		));
	notech_reg_set code_data_reg_64(.CP(n_61997), .D(n_5860), .SD(1'b1), .Q(code_data
		[64]));
	notech_mux2 i_5906(.S(\nbus_11667[64] ), .A(code_data[64]), .B(axi_R[0])
		, .Z(n_5860));
	notech_ao4 i_1199(.A(n_61502), .B(n_6779), .C(n_2244), .D(n_6887), .Z(n_2257
		));
	notech_reg_set code_data_reg_65(.CP(n_61997), .D(n_5866), .SD(1'b1), .Q(code_data
		[65]));
	notech_mux2 i_5914(.S(\nbus_11667[64] ), .A(code_data[65]), .B(axi_R[1])
		, .Z(n_5866));
	notech_reg_set code_data_reg_66(.CP(n_61997), .D(n_5872), .SD(1'b1), .Q(code_data
		[66]));
	notech_mux2 i_5922(.S(\nbus_11667[64] ), .A(code_data[66]), .B(axi_R[2])
		, .Z(n_5872));
	notech_ao4 i_1209(.A(n_2239), .B(n_6920), .C(n_2237), .D(n_6952), .Z(n_2259
		));
	notech_reg_set code_data_reg_67(.CP(n_61997), .D(n_5878), .SD(1'b1), .Q(code_data
		[67]));
	notech_mux2 i_5930(.S(\nbus_11667[64] ), .A(code_data[67]), .B(axi_R[3])
		, .Z(n_5878));
	notech_ao4 i_1208(.A(n_61502), .B(n_6780), .C(n_2244), .D(n_6888), .Z(n_2260
		));
	notech_reg_set code_data_reg_68(.CP(n_61997), .D(n_5884), .SD(1'b1), .Q(code_data
		[68]));
	notech_mux2 i_5938(.S(\nbus_11667[64] ), .A(code_data[68]), .B(axi_R[4])
		, .Z(n_5884));
	notech_reg_set code_data_reg_69(.CP(n_61997), .D(n_5890), .SD(1'b1), .Q(code_data
		[69]));
	notech_mux2 i_5946(.S(\nbus_11667[64] ), .A(code_data[69]), .B(axi_R[5])
		, .Z(n_5890));
	notech_ao4 i_1218(.A(n_2239), .B(n_6921), .C(n_2237), .D(n_6953), .Z(n_2262
		));
	notech_reg_set code_data_reg_70(.CP(n_61981), .D(n_5896), .SD(1'b1), .Q(code_data
		[70]));
	notech_mux2 i_5954(.S(\nbus_11667[64] ), .A(code_data[70]), .B(axi_R[6])
		, .Z(n_5896));
	notech_ao4 i_1217(.A(n_61502), .B(n_6781), .C(n_2244), .D(n_6889), .Z(n_2263
		));
	notech_reg_set code_data_reg_71(.CP(n_61997), .D(n_5902), .SD(1'b1), .Q(code_data
		[71]));
	notech_mux2 i_5962(.S(\nbus_11667[64] ), .A(code_data[71]), .B(axi_R[7])
		, .Z(n_5902));
	notech_reg_set code_data_reg_72(.CP(n_62003), .D(n_5908), .SD(1'b1), .Q(code_data
		[72]));
	notech_mux2 i_5970(.S(\nbus_11667[64] ), .A(code_data[72]), .B(axi_R[8])
		, .Z(n_5908));
	notech_ao4 i_1227(.A(n_2239), .B(n_6922), .C(n_2237), .D(n_6954), .Z(n_2265
		));
	notech_reg_set code_data_reg_73(.CP(n_61983), .D(n_5914), .SD(1'b1), .Q(code_data
		[73]));
	notech_mux2 i_5978(.S(\nbus_11667[64] ), .A(code_data[73]), .B(axi_R[9])
		, .Z(n_5914));
	notech_ao4 i_1226(.A(n_61502), .B(n_6782), .C(n_2244), .D(n_6890), .Z(n_2266
		));
	notech_reg_set code_data_reg_74(.CP(n_61983), .D(n_5920), .SD(1'b1), .Q(code_data
		[74]));
	notech_mux2 i_5986(.S(\nbus_11667[64] ), .A(code_data[74]), .B(axi_R[10]
		), .Z(n_5920));
	notech_reg_set code_data_reg_75(.CP(n_61983), .D(n_5926), .SD(1'b1), .Q(code_data
		[75]));
	notech_mux2 i_5994(.S(\nbus_11667[64] ), .A(code_data[75]), .B(axi_R[11]
		), .Z(n_5926));
	notech_ao4 i_1236(.A(n_2239), .B(n_6923), .C(n_2237), .D(n_6955), .Z(n_2268
		));
	notech_reg_set code_data_reg_76(.CP(n_61983), .D(n_5932), .SD(1'b1), .Q(code_data
		[76]));
	notech_mux2 i_6002(.S(\nbus_11667[64] ), .A(code_data[76]), .B(axi_R[12]
		), .Z(n_5932));
	notech_ao4 i_1235(.A(n_61502), .B(n_6783), .C(n_2244), .D(n_6891), .Z(n_2269
		));
	notech_reg_set code_data_reg_77(.CP(n_61983), .D(n_5938), .SD(1'b1), .Q(code_data
		[77]));
	notech_mux2 i_6010(.S(\nbus_11667[64] ), .A(code_data[77]), .B(axi_R[13]
		), .Z(n_5938));
	notech_reg_set code_data_reg_78(.CP(n_61983), .D(n_5944), .SD(1'b1), .Q(code_data
		[78]));
	notech_mux2 i_6018(.S(\nbus_11667[64] ), .A(code_data[78]), .B(axi_R[14]
		), .Z(n_5944));
	notech_ao4 i_1245(.A(n_2239), .B(n_6924), .C(n_2237), .D(n_6956), .Z(n_2271
		));
	notech_reg_set code_data_reg_79(.CP(n_61983), .D(n_5950), .SD(1'b1), .Q(code_data
		[79]));
	notech_mux2 i_6026(.S(\nbus_11667[64] ), .A(code_data[79]), .B(axi_R[15]
		), .Z(n_5950));
	notech_ao4 i_1244(.A(n_61502), .B(n_6784), .C(n_2244), .D(n_6892), .Z(n_2272
		));
	notech_reg_set code_data_reg_80(.CP(n_61983), .D(n_5956), .SD(1'b1), .Q(code_data
		[80]));
	notech_mux2 i_6034(.S(n_53683), .A(code_data[80]), .B(axi_R[16]), .Z(n_5956
		));
	notech_reg_set code_data_reg_81(.CP(n_61983), .D(n_5962), .SD(1'b1), .Q(code_data
		[81]));
	notech_mux2 i_6042(.S(n_53683), .A(code_data[81]), .B(axi_R[17]), .Z(n_5962
		));
	notech_ao4 i_1254(.A(n_2239), .B(n_6925), .C(n_2237), .D(n_6957), .Z(n_2274
		));
	notech_reg_set code_data_reg_82(.CP(n_61983), .D(n_5968), .SD(1'b1), .Q(code_data
		[82]));
	notech_mux2 i_6050(.S(n_53683), .A(code_data[82]), .B(axi_R[18]), .Z(n_5968
		));
	notech_ao4 i_1253(.A(n_61502), .B(n_6785), .C(n_2244), .D(n_6893), .Z(n_2275
		));
	notech_reg_set code_data_reg_83(.CP(n_62005), .D(n_5974), .SD(1'b1), .Q(code_data
		[83]));
	notech_mux2 i_6058(.S(n_53683), .A(code_data[83]), .B(axi_R[19]), .Z(n_5974
		));
	notech_reg_set code_data_reg_84(.CP(n_62005), .D(n_5980), .SD(1'b1), .Q(code_data
		[84]));
	notech_mux2 i_6066(.S(n_53683), .A(code_data[84]), .B(axi_R[20]), .Z(n_5980
		));
	notech_ao4 i_1263(.A(n_2239), .B(n_6926), .C(n_2237), .D(n_6958), .Z(n_2277
		));
	notech_reg_set code_data_reg_85(.CP(n_62005), .D(n_5986), .SD(1'b1), .Q(code_data
		[85]));
	notech_mux2 i_6074(.S(n_53683), .A(code_data[85]), .B(axi_R[21]), .Z(n_5986
		));
	notech_ao4 i_1262(.A(n_61502), .B(n_6786), .C(n_2244), .D(n_6894), .Z(n_2278
		));
	notech_reg_set code_data_reg_86(.CP(n_62005), .D(n_5992), .SD(1'b1), .Q(code_data
		[86]));
	notech_mux2 i_6082(.S(n_53683), .A(code_data[86]), .B(axi_R[22]), .Z(n_5992
		));
	notech_reg_set code_data_reg_87(.CP(n_62005), .D(n_5998), .SD(1'b1), .Q(code_data
		[87]));
	notech_mux2 i_6090(.S(n_53683), .A(code_data[87]), .B(axi_R[23]), .Z(n_5998
		));
	notech_ao4 i_1272(.A(n_2239), .B(n_6927), .C(n_2237), .D(n_6959), .Z(n_2280
		));
	notech_reg_set code_data_reg_88(.CP(n_62005), .D(n_6004), .SD(1'b1), .Q(code_data
		[88]));
	notech_mux2 i_6098(.S(n_53683), .A(code_data[88]), .B(axi_R[24]), .Z(n_6004
		));
	notech_ao4 i_1271(.A(n_61502), .B(n_6787), .C(n_2244), .D(n_6895), .Z(n_2281
		));
	notech_reg_set code_data_reg_89(.CP(n_62005), .D(n_6010), .SD(1'b1), .Q(code_data
		[89]));
	notech_mux2 i_6106(.S(n_53683), .A(code_data[89]), .B(axi_R[25]), .Z(n_6010
		));
	notech_reg_set code_data_reg_90(.CP(n_62005), .D(n_6016), .SD(1'b1), .Q(code_data
		[90]));
	notech_mux2 i_6114(.S(n_53683), .A(code_data[90]), .B(axi_R[26]), .Z(n_6016
		));
	notech_ao4 i_1281(.A(n_2239), .B(n_6928), .C(n_2237), .D(n_6960), .Z(n_2283
		));
	notech_reg_set code_data_reg_91(.CP(n_62005), .D(n_6022), .SD(1'b1), .Q(code_data
		[91]));
	notech_mux2 i_6122(.S(n_53683), .A(code_data[91]), .B(axi_R[27]), .Z(n_6022
		));
	notech_ao4 i_1280(.A(n_61502), .B(n_6788), .C(n_2244), .D(n_6896), .Z(n_2284
		));
	notech_reg_set code_data_reg_92(.CP(n_62005), .D(n_6028), .SD(1'b1), .Q(code_data
		[92]));
	notech_mux2 i_6130(.S(n_53683), .A(code_data[92]), .B(axi_R[28]), .Z(n_6028
		));
	notech_reg_set code_data_reg_93(.CP(n_62005), .D(n_6034), .SD(1'b1), .Q(code_data
		[93]));
	notech_mux2 i_6138(.S(n_53683), .A(code_data[93]), .B(axi_R[29]), .Z(n_6034
		));
	notech_ao4 i_1290(.A(n_2239), .B(n_6929), .C(n_2237), .D(n_6961), .Z(n_2286
		));
	notech_reg_set code_data_reg_94(.CP(n_62005), .D(n_6040), .SD(1'b1), .Q(code_data
		[94]));
	notech_mux2 i_6146(.S(n_53683), .A(code_data[94]), .B(axi_R[30]), .Z(n_6040
		));
	notech_ao4 i_1289(.A(n_61507), .B(n_6789), .C(n_2244), .D(n_6897), .Z(n_2287
		));
	notech_reg_set code_data_reg_95(.CP(n_62005), .D(n_6046), .SD(1'b1), .Q(code_data
		[95]));
	notech_mux2 i_6154(.S(n_53683), .A(code_data[95]), .B(axi_R[31]), .Z(n_6046
		));
	notech_reg_set code_data_reg_96(.CP(n_62005), .D(n_6052), .SD(1'b1), .Q(code_data
		[96]));
	notech_mux2 i_6162(.S(\nbus_11667[96] ), .A(code_data[96]), .B(axi_R[0])
		, .Z(n_6052));
	notech_ao4 i_1299(.A(n_2239), .B(n_6930), .C(n_2237), .D(n_6962), .Z(n_2289
		));
	notech_reg_set code_data_reg_97(.CP(n_62005), .D(n_6058), .SD(1'b1), .Q(code_data
		[97]));
	notech_mux2 i_6170(.S(\nbus_11667[96] ), .A(code_data[97]), .B(axi_R[1])
		, .Z(n_6058));
	notech_ao4 i_1298(.A(n_61507), .B(n_6790), .C(n_2244), .D(n_6898), .Z(n_2290
		));
	notech_reg_set code_data_reg_98(.CP(n_62005), .D(n_6064), .SD(1'b1), .Q(code_data
		[98]));
	notech_mux2 i_6178(.S(\nbus_11667[96] ), .A(code_data[98]), .B(axi_R[2])
		, .Z(n_6064));
	notech_reg_set code_data_reg_99(.CP(n_62005), .D(n_6070), .SD(1'b1), .Q(code_data
		[99]));
	notech_mux2 i_6186(.S(\nbus_11667[96] ), .A(code_data[99]), .B(axi_R[3])
		, .Z(n_6070));
	notech_ao4 i_1308(.A(n_53537), .B(n_6931), .C(n_53484), .D(n_6963), .Z(n_2292
		));
	notech_reg_set code_data_reg_100(.CP(n_62005), .D(n_6076), .SD(1'b1), .Q
		(code_data[100]));
	notech_mux2 i_6194(.S(\nbus_11667[96] ), .A(code_data[100]), .B(axi_R[4]
		), .Z(n_6076));
	notech_ao4 i_1307(.A(n_61507), .B(n_6791), .C(n_53548), .D(n_6899), .Z(n_2293
		));
	notech_reg_set code_data_reg_101(.CP(n_62005), .D(n_6082), .SD(1'b1), .Q
		(code_data[101]));
	notech_mux2 i_6202(.S(\nbus_11667[96] ), .A(code_data[101]), .B(axi_R[5]
		), .Z(n_6082));
	notech_reg_set code_data_reg_102(.CP(n_62027), .D(n_6088), .SD(1'b1), .Q
		(code_data[102]));
	notech_mux2 i_6210(.S(\nbus_11667[96] ), .A(code_data[102]), .B(axi_R[6]
		), .Z(n_6088));
	notech_ao4 i_1317(.A(n_53537), .B(n_6932), .C(n_53484), .D(n_6964), .Z(n_2295
		));
	notech_reg_set code_data_reg_103(.CP(n_62003), .D(n_6094), .SD(1'b1), .Q
		(code_data[103]));
	notech_mux2 i_6218(.S(\nbus_11667[96] ), .A(code_data[103]), .B(axi_R[7]
		), .Z(n_6094));
	notech_ao4 i_1316(.A(n_61507), .B(n_6792), .C(n_53548), .D(n_6900), .Z(n_2296
		));
	notech_reg_set code_data_reg_104(.CP(n_62027), .D(n_6100), .SD(1'b1), .Q
		(code_data[104]));
	notech_mux2 i_6226(.S(\nbus_11667[96] ), .A(code_data[104]), .B(axi_R[8]
		), .Z(n_6100));
	notech_reg_set code_data_reg_105(.CP(n_62027), .D(n_6106), .SD(1'b1), .Q
		(code_data[105]));
	notech_mux2 i_6234(.S(\nbus_11667[96] ), .A(code_data[105]), .B(axi_R[9]
		), .Z(n_6106));
	notech_ao4 i_1326(.A(n_53537), .B(n_6933), .C(n_53484), .D(n_6965), .Z(n_2298
		));
	notech_reg_set code_data_reg_106(.CP(n_62027), .D(n_6112), .SD(1'b1), .Q
		(code_data[106]));
	notech_mux2 i_6242(.S(\nbus_11667[96] ), .A(code_data[106]), .B(axi_R[10
		]), .Z(n_6112));
	notech_ao4 i_1325(.A(n_61507), .B(n_6793), .C(n_53548), .D(n_6901), .Z(n_2299
		));
	notech_reg_set code_data_reg_107(.CP(n_62027), .D(n_6118), .SD(1'b1), .Q
		(code_data[107]));
	notech_mux2 i_6250(.S(\nbus_11667[96] ), .A(code_data[107]), .B(axi_R[11
		]), .Z(n_6118));
	notech_reg_set code_data_reg_108(.CP(n_62027), .D(n_6124), .SD(1'b1), .Q
		(code_data[108]));
	notech_mux2 i_6258(.S(\nbus_11667[96] ), .A(code_data[108]), .B(axi_R[12
		]), .Z(n_6124));
	notech_ao4 i_1335(.A(n_53537), .B(n_6934), .C(n_53484), .D(n_6966), .Z(n_2301
		));
	notech_reg_set code_data_reg_109(.CP(n_62027), .D(n_6130), .SD(1'b1), .Q
		(code_data[109]));
	notech_mux2 i_6266(.S(\nbus_11667[96] ), .A(code_data[109]), .B(axi_R[13
		]), .Z(n_6130));
	notech_ao4 i_1334(.A(n_61507), .B(n_6794), .C(n_53548), .D(n_6902), .Z(n_2302
		));
	notech_reg_set code_data_reg_110(.CP(n_62027), .D(n_6136), .SD(1'b1), .Q
		(code_data[110]));
	notech_mux2 i_6274(.S(\nbus_11667[96] ), .A(code_data[110]), .B(axi_R[14
		]), .Z(n_6136));
	notech_reg_set code_data_reg_111(.CP(n_62027), .D(n_6142), .SD(1'b1), .Q
		(code_data[111]));
	notech_mux2 i_6282(.S(\nbus_11667[96] ), .A(code_data[111]), .B(axi_R[15
		]), .Z(n_6142));
	notech_ao4 i_1344(.A(n_53537), .B(n_6935), .C(n_53484), .D(n_6967), .Z(n_2304
		));
	notech_reg_set code_data_reg_112(.CP(n_62027), .D(n_6148), .SD(1'b1), .Q
		(code_data[112]));
	notech_mux2 i_6290(.S(n_53694), .A(code_data[112]), .B(axi_R[16]), .Z(n_6148
		));
	notech_ao4 i_1343(.A(n_61512), .B(n_6795), .C(n_53548), .D(n_6903), .Z(n_2305
		));
	notech_reg_set code_data_reg_113(.CP(n_62027), .D(n_6154), .SD(1'b1), .Q
		(code_data[113]));
	notech_mux2 i_6298(.S(n_53694), .A(code_data[113]), .B(axi_R[17]), .Z(n_6154
		));
	notech_reg_set code_data_reg_114(.CP(n_62027), .D(n_6160), .SD(1'b1), .Q
		(code_data[114]));
	notech_mux2 i_6306(.S(n_53694), .A(code_data[114]), .B(axi_R[18]), .Z(n_6160
		));
	notech_ao4 i_1353(.A(n_53537), .B(n_6936), .C(n_53484), .D(n_6968), .Z(n_2307
		));
	notech_reg_set code_data_reg_115(.CP(n_62027), .D(n_6166), .SD(1'b1), .Q
		(code_data[115]));
	notech_mux2 i_6314(.S(n_53694), .A(code_data[115]), .B(axi_R[19]), .Z(n_6166
		));
	notech_ao4 i_1352(.A(n_61507), .B(n_6796), .C(n_53548), .D(n_6904), .Z(n_2308
		));
	notech_reg_set code_data_reg_116(.CP(n_62027), .D(n_6172), .SD(1'b1), .Q
		(code_data[116]));
	notech_mux2 i_6322(.S(n_53694), .A(code_data[116]), .B(axi_R[20]), .Z(n_6172
		));
	notech_reg_set code_data_reg_117(.CP(n_62027), .D(n_6178), .SD(1'b1), .Q
		(code_data[117]));
	notech_mux2 i_6330(.S(n_53694), .A(code_data[117]), .B(axi_R[21]), .Z(n_6178
		));
	notech_ao4 i_1362(.A(n_53537), .B(n_6937), .C(n_53484), .D(n_6969), .Z(n_2310
		));
	notech_reg_set code_data_reg_118(.CP(n_62027), .D(n_6184), .SD(1'b1), .Q
		(code_data[118]));
	notech_mux2 i_6338(.S(n_53694), .A(code_data[118]), .B(axi_R[22]), .Z(n_6184
		));
	notech_ao4 i_1361(.A(n_61507), .B(n_6797), .C(n_53548), .D(n_6905), .Z(n_2311
		));
	notech_reg_set code_data_reg_119(.CP(n_62027), .D(n_6190), .SD(1'b1), .Q
		(code_data[119]));
	notech_mux2 i_6346(.S(n_53694), .A(code_data[119]), .B(axi_R[23]), .Z(n_6190
		));
	notech_reg_set code_data_reg_120(.CP(n_62027), .D(n_6196), .SD(1'b1), .Q
		(code_data[120]));
	notech_mux2 i_6354(.S(n_53694), .A(code_data[120]), .B(axi_R[24]), .Z(n_6196
		));
	notech_ao4 i_1371(.A(n_53537), .B(n_6938), .C(n_53484), .D(n_6970), .Z(n_2313
		));
	notech_reg_set code_data_reg_121(.CP(n_62027), .D(n_6202), .SD(1'b1), .Q
		(code_data[121]));
	notech_mux2 i_6362(.S(n_53694), .A(code_data[121]), .B(axi_R[25]), .Z(n_6202
		));
	notech_ao4 i_1370(.A(n_61507), .B(n_6798), .C(n_53548), .D(n_6906), .Z(n_2314
		));
	notech_reg_set code_data_reg_122(.CP(n_62003), .D(n_6208), .SD(1'b1), .Q
		(code_data[122]));
	notech_mux2 i_6370(.S(n_53694), .A(code_data[122]), .B(axi_R[26]), .Z(n_6208
		));
	notech_reg_set code_data_reg_123(.CP(n_62003), .D(n_6214), .SD(1'b1), .Q
		(code_data[123]));
	notech_mux2 i_6378(.S(n_53694), .A(code_data[123]), .B(axi_R[27]), .Z(n_6214
		));
	notech_ao4 i_1380(.A(n_53537), .B(n_6939), .C(n_53484), .D(n_6971), .Z(n_2316
		));
	notech_reg_set code_data_reg_124(.CP(n_62003), .D(n_6220), .SD(1'b1), .Q
		(code_data[124]));
	notech_mux2 i_6386(.S(n_53694), .A(code_data[124]), .B(axi_R[28]), .Z(n_6220
		));
	notech_ao4 i_1379(.A(n_61507), .B(n_6799), .C(n_53548), .D(n_6907), .Z(n_2317
		));
	notech_reg_set code_data_reg_125(.CP(n_62003), .D(n_6226), .SD(1'b1), .Q
		(code_data[125]));
	notech_mux2 i_6394(.S(n_53694), .A(code_data[125]), .B(axi_R[29]), .Z(n_6226
		));
	notech_reg_set code_data_reg_126(.CP(n_62003), .D(n_6232), .SD(1'b1), .Q
		(code_data[126]));
	notech_mux2 i_6402(.S(n_53694), .A(code_data[126]), .B(axi_R[30]), .Z(n_6232
		));
	notech_ao4 i_1389(.A(n_53537), .B(n_6940), .C(n_53484), .D(n_6972), .Z(n_2319
		));
	notech_reg_set code_data_reg_127(.CP(n_62003), .D(n_6238), .SD(1'b1), .Q
		(code_data[127]));
	notech_mux2 i_6410(.S(n_53694), .A(code_data[127]), .B(axi_R[31]), .Z(n_6238
		));
	notech_ao4 i_1388(.A(n_61507), .B(n_6800), .C(n_53548), .D(n_6908), .Z(n_2320
		));
	notech_reg axi_io_WLAST_reg(.CP(n_62003), .D(n_6244), .CD(n_61416), .Q(axi_io_WLAST
		));
	notech_mux2 i_6418(.S(n_1763), .A(n_23659), .B(axi_io_WLAST), .Z(n_6244)
		);
	notech_reg axi_WVALID_reg(.CP(n_62003), .D(n_6250), .CD(n_61416), .Q(axi_WVALID
		));
	notech_mux2 i_6426(.S(n_1218), .A(n_1176), .B(axi_WVALID), .Z(n_6250));
	notech_ao4 i_1398(.A(n_53537), .B(n_6941), .C(n_2237), .D(n_6973), .Z(n_2322
		));
	notech_reg_set axi_ARBURST_reg_0(.CP(n_62003), .D(n_6256), .SD(n_61416),
		 .Q(axi_ARBURST[0]));
	notech_or2 i_6434(.A(axi_ARBURST[0]), .B(n_6664), .Z(n_6256));
	notech_ao4 i_1397(.A(n_61507), .B(n_6801), .C(n_2244), .D(n_6909), .Z(n_2323
		));
	notech_reg axi_ARBURST_reg_1(.CP(n_62003), .D(n_6265), .CD(n_61416), .Q(axi_ARBURST
		[1]));
	notech_and2 i_6444(.A(axi_ARBURST[1]), .B(n_61491), .Z(n_6265));
	notech_reg axi_io_AW_reg_0(.CP(n_61983), .D(n_6271), .CD(n_61423), .Q(axi_io_AW
		[0]));
	notech_and2 i_6452(.A(n_6774), .B(axi_io_AW[0]), .Z(n_6271));
	notech_ao4 i_1407(.A(n_53537), .B(n_6942), .C(n_53484), .D(n_6974), .Z(n_2325
		));
	notech_reg axi_io_AW_reg_1(.CP(n_61983), .D(n_6277), .CD(n_61423), .Q(axi_io_AW
		[1]));
	notech_and2 i_6460(.A(n_6774), .B(axi_io_AW[1]), .Z(n_6277));
	notech_ao4 i_1406(.A(n_61507), .B(n_6802), .C(n_53548), .D(n_6910), .Z(n_2326
		));
	notech_reg axi_io_AW_reg_2(.CP(n_62007), .D(n_6280), .CD(n_61423), .Q(axi_io_AW
		[2]));
	notech_mux2 i_6466(.S(\nbus_11662[0] ), .A(axi_io_AW[2]), .B(io_add[0]),
		 .Z(n_6280));
	notech_reg axi_io_AW_reg_3(.CP(n_61985), .D(n_6286), .CD(n_61423), .Q(axi_io_AW
		[3]));
	notech_mux2 i_6474(.S(\nbus_11662[0] ), .A(axi_io_AW[3]), .B(io_add[1]),
		 .Z(n_6286));
	notech_ao4 i_1416(.A(n_53537), .B(n_6943), .C(n_53484), .D(n_6975), .Z(n_2328
		));
	notech_reg axi_io_AW_reg_4(.CP(n_61985), .D(n_6292), .CD(n_61423), .Q(axi_io_AW
		[4]));
	notech_mux2 i_6482(.S(\nbus_11662[0] ), .A(axi_io_AW[4]), .B(io_add[2]),
		 .Z(n_6292));
	notech_ao4 i_1415(.A(n_61507), .B(n_6803), .C(n_53548), .D(n_6911), .Z(n_2329
		));
	notech_reg axi_io_AW_reg_5(.CP(n_61985), .D(n_6298), .CD(n_61423), .Q(axi_io_AW
		[5]));
	notech_mux2 i_6490(.S(\nbus_11662[0] ), .A(axi_io_AW[5]), .B(io_add[3]),
		 .Z(n_6298));
	notech_reg axi_io_AW_reg_6(.CP(n_61985), .D(n_6304), .CD(n_61423), .Q(axi_io_AW
		[6]));
	notech_mux2 i_6498(.S(\nbus_11662[0] ), .A(axi_io_AW[6]), .B(io_add[4]),
		 .Z(n_6304));
	notech_ao4 i_1425(.A(n_53537), .B(n_6944), .C(n_53484), .D(n_6976), .Z(n_2331
		));
	notech_reg axi_io_AW_reg_7(.CP(n_61985), .D(n_6310), .CD(n_61423), .Q(axi_io_AW
		[7]));
	notech_mux2 i_6506(.S(\nbus_11662[0] ), .A(axi_io_AW[7]), .B(io_add[5]),
		 .Z(n_6310));
	notech_ao4 i_1424(.A(n_61507), .B(n_6804), .C(n_53548), .D(n_6912), .Z(n_2332
		));
	notech_reg axi_io_AW_reg_8(.CP(n_61985), .D(n_6316), .CD(n_61423), .Q(axi_io_AW
		[8]));
	notech_mux2 i_6514(.S(n_60808), .A(axi_io_AW[8]), .B(io_add[6]), .Z(n_6316
		));
	notech_reg axi_io_AW_reg_9(.CP(n_61985), .D(n_6322), .CD(n_61423), .Q(axi_io_AW
		[9]));
	notech_mux2 i_6522(.S(n_60808), .A(axi_io_AW[9]), .B(io_add[7]), .Z(n_6322
		));
	notech_ao4 i_1434(.A(n_53537), .B(n_6945), .C(n_53484), .D(n_6977), .Z(n_2334
		));
	notech_reg axi_io_AW_reg_10(.CP(n_61985), .D(n_6328), .CD(n_61422), .Q(axi_io_AW
		[10]));
	notech_mux2 i_6530(.S(n_60808), .A(axi_io_AW[10]), .B(io_add[8]), .Z(n_6328
		));
	notech_ao4 i_1433(.A(n_61507), .B(n_6805), .C(n_53548), .D(n_6913), .Z(n_2335
		));
	notech_reg axi_io_AW_reg_11(.CP(n_61985), .D(n_6334), .CD(n_61422), .Q(axi_io_AW
		[11]));
	notech_mux2 i_6538(.S(n_60808), .A(axi_io_AW[11]), .B(io_add[9]), .Z(n_6334
		));
	notech_reg axi_io_AW_reg_12(.CP(n_61985), .D(n_6340), .CD(n_61423), .Q(axi_io_AW
		[12]));
	notech_mux2 i_6546(.S(n_60808), .A(axi_io_AW[12]), .B(io_add[10]), .Z(n_6340
		));
	notech_ao4 i_1443(.A(n_53537), .B(n_6946), .C(n_53484), .D(n_6978), .Z(n_2337
		));
	notech_reg axi_io_AW_reg_13(.CP(n_62007), .D(n_6346), .CD(n_61423), .Q(axi_io_AW
		[13]));
	notech_mux2 i_6554(.S(n_60808), .A(axi_io_AW[13]), .B(io_add[11]), .Z(n_6346
		));
	notech_ao4 i_1442(.A(n_61507), .B(n_6806), .C(n_53548), .D(n_6914), .Z(n_2338
		));
	notech_reg axi_io_AW_reg_14(.CP(n_62007), .D(n_6352), .CD(n_61423), .Q(axi_io_AW
		[14]));
	notech_mux2 i_6562(.S(\nbus_11662[0] ), .A(axi_io_AW[14]), .B(io_add[12]
		), .Z(n_6352));
	notech_reg axi_io_AW_reg_15(.CP(n_62007), .D(n_6358), .CD(n_61423), .Q(axi_io_AW
		[15]));
	notech_mux2 i_6570(.S(\nbus_11662[0] ), .A(axi_io_AW[15]), .B(io_add[13]
		), .Z(n_6358));
	notech_and2 i_1098(.A(n_61423), .B(n_963), .Z(\nbus_11672[0] ));
	notech_reg axi_io_AW_reg_16(.CP(n_62007), .D(n_6364), .CD(n_61424), .Q(axi_io_AW
		[16]));
	notech_mux2 i_6578(.S(\nbus_11662[0] ), .A(axi_io_AW[16]), .B(io_add[14]
		), .Z(n_6364));
	notech_nor2 i_900(.A(n_223056061), .B(n_223356064), .Z(\nbus_11673[0] )
		);
	notech_reg axi_io_AW_reg_17(.CP(n_62007), .D(n_6370), .CD(n_61424), .Q(axi_io_AW
		[17]));
	notech_mux2 i_6586(.S(\nbus_11662[0] ), .A(axi_io_AW[17]), .B(io_add[15]
		), .Z(n_6370));
	notech_nor2 i_899(.A(n_223156062), .B(n_223056061), .Z(\nbus_11662[0] )
		);
	notech_reg axi_io_AW_reg_18(.CP(n_62007), .D(n_6379), .CD(n_61424), .Q(axi_io_AW
		[18]));
	notech_and2 i_6596(.A(axi_io_AW[18]), .B(n_6774), .Z(n_6379));
	notech_and4 i_898(.A(axi_io_RREADY), .B(axi_io_RVALID), .C(n_222856059),
		 .D(n_61424), .Z(\nbus_11671[0] ));
	notech_reg axi_io_AW_reg_19(.CP(n_62007), .D(n_6385), .CD(n_61425), .Q(axi_io_AW
		[19]));
	notech_and2 i_6604(.A(axi_io_AW[19]), .B(n_6774), .Z(n_6385));
	notech_and4 i_896(.A(burst_idx[0]), .B(burst_idx[1]), .C(n_22749), .D(n_210755938
		), .Z(\nbus_11667[96] ));
	notech_reg axi_io_AW_reg_20(.CP(n_62007), .D(n_6391), .CD(n_61425), .Q(axi_io_AW
		[20]));
	notech_and2 i_6612(.A(axi_io_AW[20]), .B(n_6774), .Z(n_6391));
	notech_and3 i_894(.A(n_210755938), .B(n_22749), .C(n_2028), .Z(\nbus_11667[64] 
		));
	notech_reg axi_io_AW_reg_21(.CP(n_62007), .D(n_6397), .CD(n_61424), .Q(axi_io_AW
		[21]));
	notech_and2 i_6620(.A(axi_io_AW[21]), .B(n_6774), .Z(n_6397));
	notech_and3 i_893(.A(n_210755938), .B(n_22749), .C(n_2029), .Z(\nbus_11667[32] 
		));
	notech_reg axi_io_AW_reg_22(.CP(n_62007), .D(n_6403), .CD(n_61424), .Q(axi_io_AW
		[22]));
	notech_and2 i_6628(.A(axi_io_AW[22]), .B(n_6774), .Z(n_6403));
	notech_ao3 i_891(.A(n_210755938), .B(n_22749), .C(n_2036), .Z(\nbus_11667[0] 
		));
	notech_reg axi_io_AW_reg_23(.CP(n_62007), .D(n_6409), .CD(n_61424), .Q(axi_io_AW
		[23]));
	notech_and2 i_6636(.A(axi_io_AW[23]), .B(n_6774), .Z(n_6409));
	notech_ao3 i_26(.A(n_6657), .B(n_2003), .C(busy), .Z(n_23592));
	notech_reg axi_io_AW_reg_24(.CP(n_62007), .D(n_6415), .CD(n_61424), .Q(axi_io_AW
		[24]));
	notech_and2 i_6644(.A(axi_io_AW[24]), .B(n_6774), .Z(n_6415));
	notech_and2 i_211(.A(axi_io_AWVALID), .B(axi_io_AWREADY), .Z(n_23659));
	notech_reg axi_io_AW_reg_25(.CP(n_62007), .D(n_6421), .CD(n_61424), .Q(axi_io_AW
		[25]));
	notech_and2 i_6652(.A(axi_io_AW[25]), .B(n_6774), .Z(n_6421));
	notech_and2 i_29(.A(axi_io_ARVALID), .B(axi_io_ARREADY), .Z(n_23604));
	notech_reg axi_io_AW_reg_26(.CP(n_62007), .D(n_6427), .CD(n_61424), .Q(axi_io_AW
		[26]));
	notech_and2 i_6660(.A(axi_io_AW[26]), .B(n_6774), .Z(n_6427));
	notech_ao3 i_918(.A(n_2003), .B(write_msk[1]), .C(n_2002), .Z(n_25361)
		);
	notech_reg axi_io_AW_reg_27(.CP(n_62007), .D(n_6433), .CD(n_61424), .Q(axi_io_AW
		[27]));
	notech_and2 i_6668(.A(axi_io_AW[27]), .B(n_6774), .Z(n_6433));
	notech_ao3 i_919(.A(n_2003), .B(write_msk[2]), .C(n_2002), .Z(n_25367)
		);
	notech_reg axi_io_AW_reg_28(.CP(n_62007), .D(n_6439), .CD(n_61424), .Q(axi_io_AW
		[28]));
	notech_and2 i_6676(.A(axi_io_AW[28]), .B(n_6774), .Z(n_6439));
	notech_ao3 i_920(.A(n_2003), .B(write_msk[3]), .C(n_2002), .Z(n_25373)
		);
	notech_reg axi_io_AW_reg_29(.CP(n_62007), .D(n_6445), .CD(n_61424), .Q(axi_io_AW
		[29]));
	notech_and2 i_6684(.A(axi_io_AW[29]), .B(n_6774), .Z(n_6445));
	notech_ao3 i_1053(.A(n_60873), .B(cacheQ[146]), .C(n_21501), .Z(n_23547)
		);
	notech_reg axi_io_AW_reg_30(.CP(n_62007), .D(n_6451), .CD(n_61424), .Q(axi_io_AW
		[30]));
	notech_and2 i_6692(.A(axi_io_AW[30]), .B(n_6774), .Z(n_6451));
	notech_ao3 i_1054(.A(n_60873), .B(cacheQ[147]), .C(n_21501), .Z(n_23552)
		);
	notech_reg axi_io_AW_reg_31(.CP(n_61985), .D(n_6457), .CD(n_61422), .Q(axi_io_AW
		[31]));
	notech_and2 i_6700(.A(axi_io_AW[31]), .B(n_6774), .Z(n_6457));
	notech_ao3 i_1055(.A(n_60873), .B(cacheQ[149]), .C(n_21501), .Z(n_23562)
		);
	notech_reg axi_io_W_reg_0(.CP(n_61985), .D(n_6460), .CD(n_61420), .Q(axi_io_W
		[0]));
	notech_mux2 i_6706(.S(\nbus_11662[0] ), .A(axi_io_W[0]), .B(writeio_data
		[0]), .Z(n_6460));
	notech_and4 i_56161(.A(fsm[4]), .B(fsm[0]), .C(n_1999), .D(n_6768), .Z(n_22749
		));
	notech_reg axi_io_W_reg_1(.CP(n_61987), .D(n_6466), .CD(n_61420), .Q(axi_io_W
		[1]));
	notech_mux2 i_6714(.S(\nbus_11662[0] ), .A(axi_io_W[1]), .B(writeio_data
		[1]), .Z(n_6466));
	notech_and2 i_1074(.A(write_data[8]), .B(n_6673), .Z(n_24863));
	notech_reg axi_io_W_reg_2(.CP(n_61987), .D(n_6472), .CD(n_61420), .Q(axi_io_W
		[2]));
	notech_mux2 i_6722(.S(\nbus_11662[0] ), .A(axi_io_W[2]), .B(writeio_data
		[2]), .Z(n_6472));
	notech_and2 i_1075(.A(write_data[9]), .B(n_6673), .Z(n_24869));
	notech_reg axi_io_W_reg_3(.CP(n_61987), .D(n_6478), .CD(n_61420), .Q(axi_io_W
		[3]));
	notech_mux2 i_6730(.S(\nbus_11662[0] ), .A(axi_io_W[3]), .B(writeio_data
		[3]), .Z(n_6478));
	notech_and2 i_1076(.A(write_data[10]), .B(n_6673), .Z(n_24875));
	notech_reg axi_io_W_reg_4(.CP(n_61987), .D(n_6484), .CD(n_61420), .Q(axi_io_W
		[4]));
	notech_mux2 i_6738(.S(\nbus_11662[0] ), .A(axi_io_W[4]), .B(writeio_data
		[4]), .Z(n_6484));
	notech_and2 i_1077(.A(write_data[11]), .B(n_6673), .Z(n_24881));
	notech_reg axi_io_W_reg_5(.CP(n_61987), .D(n_6490), .CD(n_61420), .Q(axi_io_W
		[5]));
	notech_mux2 i_6746(.S(\nbus_11662[0] ), .A(axi_io_W[5]), .B(writeio_data
		[5]), .Z(n_6490));
	notech_and2 i_1078(.A(write_data[12]), .B(n_6673), .Z(n_24887));
	notech_reg axi_io_W_reg_6(.CP(n_61987), .D(n_6496), .CD(n_61420), .Q(axi_io_W
		[6]));
	notech_mux2 i_6754(.S(\nbus_11662[0] ), .A(axi_io_W[6]), .B(writeio_data
		[6]), .Z(n_6496));
	notech_and2 i_1079(.A(write_data[13]), .B(n_6673), .Z(n_24893));
	notech_reg axi_io_W_reg_7(.CP(n_61987), .D(n_6502), .CD(n_61420), .Q(axi_io_W
		[7]));
	notech_mux2 i_6762(.S(\nbus_11662[0] ), .A(axi_io_W[7]), .B(writeio_data
		[7]), .Z(n_6502));
	notech_and2 i_1080(.A(write_data[14]), .B(n_6673), .Z(n_24899));
	notech_reg axi_io_W_reg_8(.CP(n_61987), .D(n_6508), .CD(n_61419), .Q(axi_io_W
		[8]));
	notech_mux2 i_6770(.S(n_60808), .A(axi_io_W[8]), .B(writeio_data[8]), .Z
		(n_6508));
	notech_and2 i_1081(.A(write_data[15]), .B(n_6673), .Z(n_24905));
	notech_reg axi_io_W_reg_9(.CP(n_61987), .D(n_6514), .CD(n_61419), .Q(axi_io_W
		[9]));
	notech_mux2 i_6778(.S(n_60804), .A(axi_io_W[9]), .B(writeio_data[9]), .Z
		(n_6514));
	notech_and2 i_1082(.A(write_data[16]), .B(n_6673), .Z(n_24911));
	notech_reg axi_io_W_reg_10(.CP(n_61987), .D(n_6520), .CD(n_61419), .Q(axi_io_W
		[10]));
	notech_mux2 i_6786(.S(n_60804), .A(axi_io_W[10]), .B(writeio_data[10]), 
		.Z(n_6520));
	notech_and2 i_1083(.A(write_data[17]), .B(n_6673), .Z(n_24917));
	notech_reg axi_io_W_reg_11(.CP(n_61987), .D(n_6526), .CD(n_61419), .Q(axi_io_W
		[11]));
	notech_mux2 i_6794(.S(n_60804), .A(axi_io_W[11]), .B(writeio_data[11]), 
		.Z(n_6526));
	notech_and2 i_1084(.A(write_data[18]), .B(n_6673), .Z(n_24923));
	notech_reg axi_io_W_reg_12(.CP(n_61987), .D(n_6532), .CD(n_61419), .Q(axi_io_W
		[12]));
	notech_mux2 i_6802(.S(n_60804), .A(axi_io_W[12]), .B(writeio_data[12]), 
		.Z(n_6532));
	notech_and2 i_1085(.A(write_data[19]), .B(n_6673), .Z(n_24929));
	notech_reg axi_io_W_reg_13(.CP(n_61987), .D(n_6538), .CD(n_61420), .Q(axi_io_W
		[13]));
	notech_mux2 i_6810(.S(n_60804), .A(axi_io_W[13]), .B(writeio_data[13]), 
		.Z(n_6538));
	notech_and2 i_1086(.A(write_data[20]), .B(n_60817), .Z(n_24935));
	notech_reg axi_io_W_reg_14(.CP(n_61987), .D(n_6544), .CD(n_61419), .Q(axi_io_W
		[14]));
	notech_mux2 i_6818(.S(n_60804), .A(axi_io_W[14]), .B(writeio_data[14]), 
		.Z(n_6544));
	notech_and2 i_1087(.A(write_data[21]), .B(n_60817), .Z(n_24941));
	notech_reg axi_io_W_reg_15(.CP(n_61987), .D(n_6550), .CD(n_61419), .Q(axi_io_W
		[15]));
	notech_mux2 i_6826(.S(n_60804), .A(axi_io_W[15]), .B(writeio_data[15]), 
		.Z(n_6550));
	notech_and2 i_1088(.A(write_data[22]), .B(n_60817), .Z(n_24947));
	notech_reg axi_io_W_reg_16(.CP(n_61987), .D(n_6556), .CD(n_61420), .Q(axi_io_W
		[16]));
	notech_mux2 i_6834(.S(n_60804), .A(axi_io_W[16]), .B(writeio_data[16]), 
		.Z(n_6556));
	notech_and2 i_1089(.A(write_data[23]), .B(n_60817), .Z(n_24953));
	notech_reg axi_io_W_reg_17(.CP(n_61987), .D(n_6562), .CD(n_61422), .Q(axi_io_W
		[17]));
	notech_mux2 i_6842(.S(n_60804), .A(axi_io_W[17]), .B(writeio_data[17]), 
		.Z(n_6562));
	notech_and2 i_1090(.A(write_data[24]), .B(n_60817), .Z(n_24959));
	notech_reg axi_io_W_reg_18(.CP(n_61987), .D(n_6568), .CD(n_61422), .Q(axi_io_W
		[18]));
	notech_mux2 i_6850(.S(n_60804), .A(axi_io_W[18]), .B(writeio_data[18]), 
		.Z(n_6568));
	notech_and2 i_1091(.A(write_data[25]), .B(n_60817), .Z(n_24965));
	notech_reg axi_io_W_reg_19(.CP(n_61987), .D(n_6574), .CD(n_61422), .Q(axi_io_W
		[19]));
	notech_mux2 i_6858(.S(n_60804), .A(axi_io_W[19]), .B(writeio_data[19]), 
		.Z(n_6574));
	notech_and2 i_1092(.A(write_data[26]), .B(n_60817), .Z(n_24971));
	notech_reg axi_io_W_reg_20(.CP(clk), .D(n_6580), .CD(n_61422), .Q(axi_io_W
		[20]));
	notech_mux2 i_6866(.S(n_60804), .A(axi_io_W[20]), .B(writeio_data[20]), 
		.Z(n_6580));
	notech_and2 i_1093(.A(write_data[27]), .B(n_60817), .Z(n_24977));
	notech_reg axi_io_W_reg_21(.CP(clk), .D(n_6586), .CD(n_61422), .Q(axi_io_W
		[21]));
	notech_mux2 i_6874(.S(n_60808), .A(axi_io_W[21]), .B(writeio_data[21]), 
		.Z(n_6586));
	notech_and2 i_1094(.A(write_data[28]), .B(n_60817), .Z(n_24983));
	notech_reg axi_io_W_reg_22(.CP(clk), .D(n_6592), .CD(n_61422), .Q(axi_io_W
		[22]));
	notech_mux2 i_6882(.S(n_60808), .A(axi_io_W[22]), .B(writeio_data[22]), 
		.Z(n_6592));
	notech_and2 i_1095(.A(write_data[29]), .B(n_60817), .Z(n_24989));
	notech_reg axi_io_W_reg_23(.CP(clk), .D(n_6598), .CD(n_61422), .Q(axi_io_W
		[23]));
	notech_mux2 i_6890(.S(n_60808), .A(axi_io_W[23]), .B(writeio_data[23]), 
		.Z(n_6598));
	notech_and2 i_1096(.A(write_data[30]), .B(n_60817), .Z(n_24995));
	notech_reg axi_io_W_reg_24(.CP(clk), .D(n_6604), .CD(n_61422), .Q(axi_io_W
		[24]));
	notech_mux2 i_6898(.S(n_60808), .A(axi_io_W[24]), .B(writeio_data[24]), 
		.Z(n_6604));
	notech_and2 i_1097(.A(write_data[31]), .B(n_60817), .Z(n_25001));
	notech_reg axi_io_W_reg_25(.CP(clk), .D(n_6610), .CD(n_61420), .Q(axi_io_W
		[25]));
	notech_mux2 i_6906(.S(n_60808), .A(axi_io_W[25]), .B(writeio_data[25]), 
		.Z(n_6610));
	notech_ao4 i_1104(.A(n_2029), .B(n_2028), .C(n_22749), .D(n_60835), .Z(n_25530
		));
	notech_reg axi_io_W_reg_26(.CP(clk), .D(n_6616), .CD(n_61420), .Q(axi_io_W
		[26]));
	notech_mux2 i_6914(.S(n_60808), .A(axi_io_W[26]), .B(writeio_data[26]), 
		.Z(n_6616));
	notech_nor2 i_1105(.A(n_965), .B(n_2024), .Z(n_25535));
	notech_reg axi_io_W_reg_27(.CP(clk), .D(n_6622), .CD(n_61420), .Q(axi_io_W
		[27]));
	notech_mux2 i_6922(.S(n_60804), .A(axi_io_W[27]), .B(writeio_data[27]), 
		.Z(n_6622));
	notech_nor2 i_1106(.A(n_2024), .B(n_966), .Z(n_25540));
	notech_reg axi_io_W_reg_28(.CP(clk), .D(n_6628), .CD(n_61420), .Q(axi_io_W
		[28]));
	notech_mux2 i_6930(.S(n_60804), .A(axi_io_W[28]), .B(writeio_data[28]), 
		.Z(n_6628));
	notech_nor2 i_1107(.A(n_2024), .B(n_967), .Z(n_25545));
	notech_reg axi_io_W_reg_29(.CP(clk), .D(n_6634), .CD(n_61422), .Q(axi_io_W
		[29]));
	notech_mux2 i_6938(.S(n_60804), .A(axi_io_W[29]), .B(writeio_data[29]), 
		.Z(n_6634));
	notech_and4 i_56174(.A(fsm[4]), .B(n_1999), .C(fsm[3]), .D(n_6765), .Z(n_25082
		));
	notech_reg axi_io_W_reg_30(.CP(clk), .D(n_6640), .CD(n_61422), .Q(axi_io_W
		[30]));
	notech_mux2 i_6946(.S(n_60808), .A(axi_io_W[30]), .B(writeio_data[30]), 
		.Z(n_6640));
	notech_reg axi_io_W_reg_31(.CP(clk), .D(n_6646), .CD(n_61420), .Q(axi_io_W
		[31]));
	notech_mux2 i_6954(.S(n_60808), .A(axi_io_W[31]), .B(writeio_data[31]), 
		.Z(n_6646));
	notech_inv i_9031(.A(n_60835), .Z(n_6652));
	notech_inv i_9032(.A(n_2052), .Z(n_6653));
	notech_inv i_9033(.A(n_2016), .Z(n_6654));
	notech_inv i_9034(.A(n_221956050), .Z(n_6655));
	notech_inv i_9035(.A(n_2050), .Z(n_6656));
	notech_inv i_9036(.A(n_970), .Z(n_6657));
	notech_inv i_9037(.A(n_222856059), .Z(n_6658));
	notech_inv i_9038(.A(n_222956060), .Z(n_6659));
	notech_inv i_9039(.A(n_2037), .Z(n_6660));
	notech_inv i_9040(.A(n_2069), .Z(n_6661));
	notech_inv i_9041(.A(n_2029), .Z(n_6662));
	notech_inv i_9042(.A(n_2028), .Z(n_6663));
	notech_inv i_9043(.A(n_61491), .Z(n_6664));
	notech_inv i_9044(.A(n_1742), .Z(n_6665));
	notech_inv i_9045(.A(n_973), .Z(n_6666));
	notech_inv i_9046(.A(n_980), .Z(n_6667));
	notech_inv i_9047(.A(n_983), .Z(n_6668));
	notech_inv i_9048(.A(n_2042), .Z(n_6669));
	notech_inv i_9049(.A(n_986), .Z(n_6670));
	notech_inv i_9050(.A(n_989), .Z(n_6671));
	notech_inv i_9051(.A(n_992), .Z(n_6672));
	notech_inv i_9052(.A(n_61437), .Z(n_6673));
	notech_inv i_9053(.A(n_995), .Z(n_6674));
	notech_inv i_9054(.A(n_998), .Z(n_6675));
	notech_inv i_9055(.A(n_1001), .Z(n_6676));
	notech_inv i_9056(.A(n_1004), .Z(n_6677));
	notech_inv i_9057(.A(n_1007), .Z(n_6678));
	notech_inv i_9058(.A(n_1010), .Z(n_6679));
	notech_inv i_9059(.A(n_1013), .Z(n_6680));
	notech_inv i_9060(.A(n_1016), .Z(n_6681));
	notech_inv i_9061(.A(n_1019), .Z(n_6682));
	notech_inv i_9062(.A(n_1022), .Z(n_6683));
	notech_inv i_9063(.A(n_1025), .Z(n_6684));
	notech_inv i_9064(.A(n_1028), .Z(n_6685));
	notech_inv i_9065(.A(n_1031), .Z(n_6686));
	notech_inv i_9066(.A(n_1034), .Z(n_6687));
	notech_inv i_9067(.A(n_1037), .Z(n_6688));
	notech_inv i_9068(.A(n_1040), .Z(n_6689));
	notech_inv i_9069(.A(n_1043), .Z(n_6690));
	notech_inv i_9070(.A(n_1046), .Z(n_6691));
	notech_inv i_9071(.A(n_1049), .Z(n_6692));
	notech_inv i_9072(.A(n_1052), .Z(n_6693));
	notech_inv i_9073(.A(n_1055), .Z(n_6694));
	notech_inv i_9074(.A(n_1058), .Z(n_6695));
	notech_inv i_9075(.A(n_1062), .Z(n_6696));
	notech_inv i_9076(.A(n_1065), .Z(n_6697));
	notech_inv i_9077(.A(n_1070), .Z(n_6698));
	notech_inv i_9078(.A(n_1073), .Z(n_6699));
	notech_inv i_9079(.A(n_1076), .Z(n_6700));
	notech_inv i_9080(.A(n_1079), .Z(n_6701));
	notech_inv i_9081(.A(n_1082), .Z(n_6702));
	notech_inv i_9082(.A(n_1085), .Z(n_6703));
	notech_inv i_9083(.A(n_1088), .Z(n_6704));
	notech_inv i_9084(.A(n_22749), .Z(n_6705));
	notech_inv i_9085(.A(n_1091), .Z(n_6706));
	notech_inv i_9086(.A(n_1094), .Z(n_6707));
	notech_inv i_9087(.A(n_1097), .Z(n_6708));
	notech_inv i_9088(.A(n_1100), .Z(n_6709));
	notech_inv i_9089(.A(n_1103), .Z(n_6710));
	notech_inv i_9090(.A(n_1106), .Z(n_6711));
	notech_inv i_9091(.A(n_1109), .Z(n_6712));
	notech_inv i_9092(.A(n_1112), .Z(n_6713));
	notech_inv i_9093(.A(n_1115), .Z(n_6714));
	notech_inv i_9094(.A(n_1118), .Z(n_6715));
	notech_inv i_9095(.A(n_1121), .Z(n_6716));
	notech_inv i_9096(.A(n_1124), .Z(n_6717));
	notech_inv i_9097(.A(n_1127), .Z(n_6718));
	notech_inv i_9098(.A(n_1130), .Z(n_6719));
	notech_inv i_9099(.A(n_1133), .Z(n_6720));
	notech_inv i_9100(.A(n_1136), .Z(n_6721));
	notech_inv i_9101(.A(n_1139), .Z(n_6722));
	notech_inv i_9102(.A(n_1142), .Z(n_6723));
	notech_inv i_9103(.A(n_1145), .Z(n_6724));
	notech_inv i_9104(.A(n_1148), .Z(n_6725));
	notech_inv i_9105(.A(n_1151), .Z(n_6726));
	notech_inv i_9106(.A(n_1154), .Z(n_6727));
	notech_inv i_9107(.A(n_1157), .Z(n_6728));
	notech_inv i_9108(.A(n_1160), .Z(n_6729));
	notech_inv i_9109(.A(n_1173), .Z(n_6730));
	notech_inv i_9110(.A(n_1179), .Z(n_6731));
	notech_inv i_9111(.A(n_1182), .Z(n_6732));
	notech_inv i_9112(.A(n_1185), .Z(n_6733));
	notech_inv i_9113(.A(n_1188), .Z(n_6734));
	notech_inv i_9114(.A(n_1191), .Z(n_6735));
	notech_inv i_9115(.A(n_1194), .Z(n_6736));
	notech_inv i_9116(.A(n_1197), .Z(n_6737));
	notech_inv i_9117(.A(n_1200), .Z(n_6738));
	notech_inv i_9118(.A(n_1213), .Z(n_6739));
	notech_inv i_9119(.A(n_1221), .Z(n_6740));
	notech_inv i_9120(.A(n_1223), .Z(n_6741));
	notech_inv i_9121(.A(burst_idx[1]), .Z(n_6742));
	notech_inv i_9122(.A(burst_idx[2]), .Z(n_6743));
	notech_inv i_9123(.A(burst_idx[3]), .Z(n_6744));
	notech_inv i_9124(.A(n_1227), .Z(n_6745));
	notech_inv i_9125(.A(n_1230), .Z(n_6746));
	notech_inv i_9127(.A(n_1233), .Z(n_6748));
	notech_inv i_9128(.A(n_1236), .Z(n_6749));
	notech_inv i_9129(.A(n_1239), .Z(n_6750));
	notech_inv i_9130(.A(n_1242), .Z(n_6751));
	notech_inv i_9131(.A(n_1245), .Z(n_6752));
	notech_inv i_9132(.A(n_1248), .Z(n_6753));
	notech_inv i_9133(.A(n_1251), .Z(n_6754));
	notech_inv i_9134(.A(n_1254), .Z(n_6755));
	notech_inv i_9135(.A(n_1257), .Z(n_6756));
	notech_inv i_9136(.A(n_1260), .Z(n_6757));
	notech_inv i_9137(.A(n_1263), .Z(n_6758));
	notech_inv i_9138(.A(n_1266), .Z(n_6759));
	notech_inv i_9139(.A(n_1269), .Z(n_6760));
	notech_inv i_9140(.A(n_1272), .Z(n_6761));
	notech_inv i_9141(.A(n_1275), .Z(n_6762));
	notech_inv i_9142(.A(n_23592), .Z(n_6763));
	notech_inv i_9143(.A(n_1280), .Z(n_6764));
	notech_inv i_9144(.A(fsm[0]), .Z(n_6765));
	notech_inv i_9145(.A(fsm[1]), .Z(n_6766));
	notech_inv i_9146(.A(fsm[2]), .Z(n_6767));
	notech_inv i_9147(.A(fsm[3]), .Z(n_6768));
	notech_inv i_9148(.A(wf), .Z(n_6769));
	notech_inv i_9149(.A(n_23604), .Z(n_6770));
	notech_inv i_9150(.A(\nbus_11673[0] ), .Z(n_6771));
	notech_inv i_9151(.A(n_1710), .Z(n_6772));
	notech_inv i_9152(.A(n_23659), .Z(n_6773));
	notech_inv i_9153(.A(n_60808), .Z(n_6774));
	notech_inv i_9154(.A(axi_R[0]), .Z(n_6775));
	notech_inv i_9155(.A(axi_R[1]), .Z(n_6776));
	notech_inv i_9156(.A(axi_R[2]), .Z(n_6777));
	notech_inv i_9157(.A(axi_R[3]), .Z(n_6778));
	notech_inv i_9158(.A(axi_R[4]), .Z(n_6779));
	notech_inv i_9159(.A(axi_R[5]), .Z(n_6780));
	notech_inv i_9160(.A(axi_R[6]), .Z(n_6781));
	notech_inv i_9161(.A(axi_R[7]), .Z(n_6782));
	notech_inv i_9162(.A(axi_R[8]), .Z(n_6783));
	notech_inv i_9163(.A(axi_R[9]), .Z(n_6784));
	notech_inv i_9164(.A(axi_R[10]), .Z(n_6785));
	notech_inv i_9165(.A(axi_R[11]), .Z(n_6786));
	notech_inv i_9166(.A(axi_R[12]), .Z(n_6787));
	notech_inv i_9167(.A(axi_R[13]), .Z(n_6788));
	notech_inv i_9168(.A(axi_R[14]), .Z(n_6789));
	notech_inv i_9169(.A(axi_R[15]), .Z(n_6790));
	notech_inv i_9170(.A(axi_R[16]), .Z(n_6791));
	notech_inv i_9171(.A(axi_R[17]), .Z(n_6792));
	notech_inv i_9172(.A(axi_R[18]), .Z(n_6793));
	notech_inv i_9173(.A(axi_R[19]), .Z(n_6794));
	notech_inv i_9174(.A(axi_R[20]), .Z(n_6795));
	notech_inv i_9175(.A(axi_R[21]), .Z(n_6796));
	notech_inv i_9176(.A(axi_R[22]), .Z(n_6797));
	notech_inv i_9177(.A(axi_R[23]), .Z(n_6798));
	notech_inv i_9178(.A(axi_R[24]), .Z(n_6799));
	notech_inv i_9179(.A(axi_R[25]), .Z(n_6800));
	notech_inv i_9180(.A(axi_R[26]), .Z(n_6801));
	notech_inv i_9181(.A(axi_R[27]), .Z(n_6802));
	notech_inv i_9182(.A(axi_R[28]), .Z(n_6803));
	notech_inv i_9183(.A(axi_R[29]), .Z(n_6804));
	notech_inv i_9184(.A(axi_R[30]), .Z(n_6805));
	notech_inv i_9185(.A(axi_R[31]), .Z(n_6806));
	notech_inv i_9186(.A(Daddr[2]), .Z(n_6807));
	notech_inv i_9187(.A(Daddr[3]), .Z(n_6808));
	notech_inv i_9188(.A(Daddr[13]), .Z(n_6809));
	notech_inv i_9189(.A(Daddr[12]), .Z(n_6810));
	notech_inv i_9190(.A(Daddr[11]), .Z(n_6811));
	notech_inv i_9191(.A(Daddr[10]), .Z(n_6812));
	notech_inv i_9192(.A(Daddr[9]), .Z(n_6813));
	notech_inv i_9193(.A(Daddr[8]), .Z(n_6814));
	notech_inv i_9194(.A(Daddr[7]), .Z(n_6815));
	notech_inv i_9195(.A(Daddr[6]), .Z(n_6816));
	notech_inv i_9196(.A(Daddr[5]), .Z(n_6817));
	notech_inv i_9197(.A(Daddr[4]), .Z(n_6818));
	notech_inv i_9198(.A(Daddr[14]), .Z(n_6819));
	notech_inv i_9199(.A(Daddr[15]), .Z(n_6820));
	notech_inv i_9200(.A(Daddr[16]), .Z(n_6821));
	notech_inv i_9201(.A(Daddr[17]), .Z(n_6822));
	notech_inv i_9202(.A(Daddr[18]), .Z(n_6823));
	notech_inv i_9203(.A(Daddr[19]), .Z(n_6824));
	notech_inv i_9204(.A(Daddr[20]), .Z(n_6825));
	notech_inv i_9205(.A(Daddr[21]), .Z(n_6826));
	notech_inv i_9206(.A(Daddr[22]), .Z(n_6827));
	notech_inv i_9207(.A(Daddr[23]), .Z(n_6828));
	notech_inv i_9208(.A(Daddr[24]), .Z(n_6829));
	notech_inv i_9209(.A(Daddr[25]), .Z(n_6830));
	notech_inv i_9210(.A(Daddr[26]), .Z(n_6831));
	notech_inv i_9211(.A(Daddr[27]), .Z(n_6832));
	notech_inv i_9212(.A(Daddr[28]), .Z(n_6833));
	notech_inv i_9213(.A(Daddr[29]), .Z(n_6834));
	notech_inv i_9214(.A(Daddr[30]), .Z(n_6835));
	notech_inv i_9215(.A(Daddr[31]), .Z(n_6836));
	notech_inv i_9216(.A(code_wdata[0]), .Z(n_6837));
	notech_inv i_9217(.A(code_wdata[1]), .Z(n_6838));
	notech_inv i_9218(.A(code_wdata[2]), .Z(n_6839));
	notech_inv i_9219(.A(code_wdata[3]), .Z(n_6840));
	notech_inv i_9220(.A(code_wdata[4]), .Z(n_6841));
	notech_inv i_9221(.A(code_wdata[5]), .Z(n_6842));
	notech_inv i_9222(.A(code_wdata[6]), .Z(n_6843));
	notech_inv i_9223(.A(code_wdata[7]), .Z(n_6844));
	notech_inv i_9224(.A(code_addr[2]), .Z(n_6845));
	notech_inv i_9225(.A(code_addr[3]), .Z(n_6846));
	notech_inv i_9226(.A(code_addr[4]), .Z(n_6847));
	notech_inv i_9227(.A(code_addr[5]), .Z(n_6848));
	notech_inv i_9228(.A(code_addr[6]), .Z(n_6849));
	notech_inv i_9229(.A(code_addr[7]), .Z(n_6850));
	notech_inv i_9230(.A(code_addr[8]), .Z(n_6851));
	notech_inv i_9231(.A(code_addr[9]), .Z(n_6852));
	notech_inv i_9232(.A(code_addr[10]), .Z(n_6853));
	notech_inv i_9233(.A(code_addr[11]), .Z(n_6854));
	notech_inv i_9234(.A(code_addr[12]), .Z(n_6855));
	notech_inv i_9235(.A(code_addr[13]), .Z(n_6856));
	notech_inv i_9236(.A(code_addr[14]), .Z(n_6857));
	notech_inv i_9237(.A(code_addr[15]), .Z(n_6858));
	notech_inv i_9238(.A(code_addr[16]), .Z(n_6859));
	notech_inv i_9239(.A(code_addr[17]), .Z(n_6860));
	notech_inv i_9240(.A(code_addr[18]), .Z(n_6861));
	notech_inv i_9241(.A(code_addr[19]), .Z(n_6862));
	notech_inv i_9242(.A(code_addr[20]), .Z(n_6863));
	notech_inv i_9243(.A(code_addr[21]), .Z(n_6864));
	notech_inv i_9244(.A(code_addr[22]), .Z(n_6865));
	notech_inv i_9245(.A(code_addr[23]), .Z(n_6866));
	notech_inv i_9246(.A(code_addr[24]), .Z(n_6867));
	notech_inv i_9247(.A(code_addr[25]), .Z(n_6868));
	notech_inv i_9248(.A(code_addr[26]), .Z(n_6869));
	notech_inv i_9249(.A(code_addr[27]), .Z(n_6870));
	notech_inv i_9250(.A(code_addr[28]), .Z(n_6871));
	notech_inv i_9251(.A(code_addr[29]), .Z(n_6872));
	notech_inv i_9252(.A(code_addr[30]), .Z(n_6873));
	notech_inv i_9253(.A(code_addr[31]), .Z(n_6874));
	notech_inv i_9254(.A(write_data[0]), .Z(n_6875));
	notech_inv i_9255(.A(write_data[1]), .Z(n_6876));
	notech_inv i_9256(.A(write_data[2]), .Z(n_6877));
	notech_inv i_9257(.A(write_data[3]), .Z(n_6878));
	notech_inv i_9258(.A(write_data[4]), .Z(n_6879));
	notech_inv i_9259(.A(write_data[5]), .Z(n_6880));
	notech_inv i_9260(.A(write_data[6]), .Z(n_6881));
	notech_inv i_9261(.A(write_data[7]), .Z(n_6882));
	notech_inv i_9262(.A(cacheQ[0]), .Z(n_6883));
	notech_inv i_9263(.A(cacheQ[1]), .Z(n_6884));
	notech_inv i_9264(.A(cacheQ[2]), .Z(n_6885));
	notech_inv i_9265(.A(cacheQ[3]), .Z(n_6886));
	notech_inv i_9266(.A(cacheQ[4]), .Z(n_6887));
	notech_inv i_9267(.A(cacheQ[5]), .Z(n_6888));
	notech_inv i_9268(.A(cacheQ[6]), .Z(n_6889));
	notech_inv i_9269(.A(cacheQ[7]), .Z(n_6890));
	notech_inv i_9270(.A(cacheQ[8]), .Z(n_6891));
	notech_inv i_9271(.A(cacheQ[9]), .Z(n_6892));
	notech_inv i_9272(.A(cacheQ[10]), .Z(n_6893));
	notech_inv i_9273(.A(cacheQ[11]), .Z(n_6894));
	notech_inv i_9274(.A(cacheQ[12]), .Z(n_6895));
	notech_inv i_9275(.A(cacheQ[13]), .Z(n_6896));
	notech_inv i_9276(.A(cacheQ[14]), .Z(n_6897));
	notech_inv i_9277(.A(cacheQ[15]), .Z(n_6898));
	notech_inv i_9278(.A(cacheQ[16]), .Z(n_6899));
	notech_inv i_9279(.A(cacheQ[17]), .Z(n_6900));
	notech_inv i_9280(.A(cacheQ[18]), .Z(n_6901));
	notech_inv i_9281(.A(cacheQ[19]), .Z(n_6902));
	notech_inv i_9282(.A(cacheQ[20]), .Z(n_6903));
	notech_inv i_9283(.A(cacheQ[21]), .Z(n_6904));
	notech_inv i_9284(.A(cacheQ[22]), .Z(n_6905));
	notech_inv i_9285(.A(cacheQ[23]), .Z(n_6906));
	notech_inv i_9286(.A(cacheQ[24]), .Z(n_6907));
	notech_inv i_9287(.A(cacheQ[25]), .Z(n_6908));
	notech_inv i_9288(.A(cacheQ[26]), .Z(n_6909));
	notech_inv i_9289(.A(cacheQ[27]), .Z(n_6910));
	notech_inv i_9290(.A(cacheQ[28]), .Z(n_6911));
	notech_inv i_9291(.A(cacheQ[29]), .Z(n_6912));
	notech_inv i_9292(.A(cacheQ[30]), .Z(n_6913));
	notech_inv i_9293(.A(cacheQ[31]), .Z(n_6914));
	notech_inv i_9294(.A(cacheQ[32]), .Z(n_6915));
	notech_inv i_9295(.A(cacheQ[33]), .Z(n_6916));
	notech_inv i_9296(.A(cacheQ[34]), .Z(n_6917));
	notech_inv i_9297(.A(cacheQ[35]), .Z(n_6918));
	notech_inv i_9298(.A(cacheQ[36]), .Z(n_6919));
	notech_inv i_9299(.A(cacheQ[37]), .Z(n_6920));
	notech_inv i_9300(.A(cacheQ[38]), .Z(n_6921));
	notech_inv i_9301(.A(cacheQ[39]), .Z(n_6922));
	notech_inv i_9302(.A(cacheQ[40]), .Z(n_6923));
	notech_inv i_9303(.A(cacheQ[41]), .Z(n_6924));
	notech_inv i_9304(.A(cacheQ[42]), .Z(n_6925));
	notech_inv i_9305(.A(cacheQ[43]), .Z(n_6926));
	notech_inv i_9306(.A(cacheQ[44]), .Z(n_6927));
	notech_inv i_9307(.A(cacheQ[45]), .Z(n_6928));
	notech_inv i_9308(.A(cacheQ[46]), .Z(n_6929));
	notech_inv i_9309(.A(cacheQ[47]), .Z(n_6930));
	notech_inv i_9310(.A(cacheQ[48]), .Z(n_6931));
	notech_inv i_9311(.A(cacheQ[49]), .Z(n_6932));
	notech_inv i_9312(.A(cacheQ[50]), .Z(n_6933));
	notech_inv i_9313(.A(cacheQ[51]), .Z(n_6934));
	notech_inv i_9314(.A(cacheQ[52]), .Z(n_6935));
	notech_inv i_9315(.A(cacheQ[53]), .Z(n_6936));
	notech_inv i_9316(.A(cacheQ[54]), .Z(n_6937));
	notech_inv i_9317(.A(cacheQ[55]), .Z(n_6938));
	notech_inv i_9318(.A(cacheQ[56]), .Z(n_6939));
	notech_inv i_9319(.A(cacheQ[57]), .Z(n_6940));
	notech_inv i_9320(.A(cacheQ[58]), .Z(n_6941));
	notech_inv i_9321(.A(cacheQ[59]), .Z(n_6942));
	notech_inv i_9322(.A(cacheQ[60]), .Z(n_6943));
	notech_inv i_9323(.A(cacheQ[61]), .Z(n_6944));
	notech_inv i_9324(.A(cacheQ[62]), .Z(n_6945));
	notech_inv i_9325(.A(cacheQ[63]), .Z(n_6946));
	notech_inv i_9326(.A(cacheQ[96]), .Z(n_6947));
	notech_inv i_9327(.A(cacheQ[97]), .Z(n_6948));
	notech_inv i_9328(.A(cacheQ[98]), .Z(n_6949));
	notech_inv i_9329(.A(cacheQ[99]), .Z(n_6950));
	notech_inv i_9330(.A(cacheQ[100]), .Z(n_6951));
	notech_inv i_9331(.A(cacheQ[101]), .Z(n_6952));
	notech_inv i_9332(.A(cacheQ[102]), .Z(n_6953));
	notech_inv i_9333(.A(cacheQ[103]), .Z(n_6954));
	notech_inv i_9334(.A(cacheQ[104]), .Z(n_6955));
	notech_inv i_9335(.A(cacheQ[105]), .Z(n_6956));
	notech_inv i_9336(.A(cacheQ[106]), .Z(n_6957));
	notech_inv i_9337(.A(cacheQ[107]), .Z(n_6958));
	notech_inv i_9338(.A(cacheQ[108]), .Z(n_6959));
	notech_inv i_9339(.A(cacheQ[109]), .Z(n_6960));
	notech_inv i_9340(.A(cacheQ[110]), .Z(n_6961));
	notech_inv i_9341(.A(cacheQ[111]), .Z(n_6962));
	notech_inv i_9342(.A(cacheQ[112]), .Z(n_6963));
	notech_inv i_9343(.A(cacheQ[113]), .Z(n_6964));
	notech_inv i_9344(.A(cacheQ[114]), .Z(n_6965));
	notech_inv i_9345(.A(cacheQ[115]), .Z(n_6966));
	notech_inv i_9346(.A(cacheQ[116]), .Z(n_6967));
	notech_inv i_9347(.A(cacheQ[117]), .Z(n_6968));
	notech_inv i_9348(.A(cacheQ[118]), .Z(n_6969));
	notech_inv i_9349(.A(cacheQ[119]), .Z(n_6970));
	notech_inv i_9350(.A(cacheQ[120]), .Z(n_6971));
	notech_inv i_9351(.A(cacheQ[121]), .Z(n_6972));
	notech_inv i_9352(.A(cacheQ[122]), .Z(n_6973));
	notech_inv i_9353(.A(cacheQ[123]), .Z(n_6974));
	notech_inv i_9354(.A(cacheQ[124]), .Z(n_6975));
	notech_inv i_9355(.A(cacheQ[125]), .Z(n_6976));
	notech_inv i_9356(.A(cacheQ[126]), .Z(n_6977));
	notech_inv i_9357(.A(cacheQ[127]), .Z(n_6978));
	notech_inv i_9358(.A(cacheQ[128]), .Z(n_6979));
	notech_inv i_9359(.A(cacheQ[129]), .Z(n_6980));
	notech_inv i_9360(.A(cacheQ[130]), .Z(n_6981));
	notech_inv i_9361(.A(cacheQ[131]), .Z(n_6982));
	notech_inv i_9362(.A(cacheQ[132]), .Z(n_6983));
	notech_inv i_9363(.A(cacheQ[133]), .Z(n_6984));
	notech_inv i_9364(.A(cacheQ[134]), .Z(n_6985));
	notech_inv i_9365(.A(cacheQ[135]), .Z(n_6986));
	notech_inv i_9366(.A(cacheQ[136]), .Z(n_6987));
	notech_inv i_9367(.A(cacheQ[137]), .Z(n_6988));
	notech_inv i_9368(.A(cacheQ[138]), .Z(n_6989));
	notech_inv i_9369(.A(cacheQ[139]), .Z(n_6990));
	notech_inv i_9370(.A(cacheQ[140]), .Z(n_6991));
	notech_inv i_9371(.A(cacheQ[141]), .Z(n_6992));
	notech_inv i_9372(.A(cacheQ[142]), .Z(n_6993));
	notech_inv i_9373(.A(cacheQ[143]), .Z(n_6994));
	notech_inv i_9374(.A(cacheQ[144]), .Z(n_6995));
	notech_inv i_9375(.A(cacheQ[145]), .Z(n_6996));
	notech_inv i_9376(.A(cacheQ[148]), .Z(n_6997));
	notech_inv i_9377(.A(write_msk[0]), .Z(n_6998));
	notech_inv i_9378(.A(axi_AR[31]), .Z(n_6999));
	notech_inv i_9379(.A(writeio_ack), .Z(n_7000));
	notech_inv i_9380(.A(n_61422), .Z(n_7001));
	notech_inv i_9381(.A(n_21501), .Z(n_7002));
	notech_inv i_9382(.A(write_ack), .Z(n_7003));
	notech_inv i_9383(.A(code_req), .Z(n_7004));
	notech_inv i_9384(.A(read_req), .Z(n_7005));
	notech_inv i_9385(.A(code_wreq), .Z(n_7006));
	datacache datacache1(.A(cacheA), .D(cacheD), .Q(cacheQ), .M(cacheM), .WEN
		(cacheWEN), .clk(clk));
endmodule
module AWDP_INC_34(O0, fsm5_cnt);

	output [8:0] O0;
	input [8:0] fsm5_cnt;




	notech_ha2 i_8(.A(fsm5_cnt[8]), .B(n_86), .Z(O0[8]));
	notech_ha2 i_7(.A(fsm5_cnt[7]), .B(n_84), .Z(O0[7]), .CO(n_86));
	notech_ha2 i_6(.A(fsm5_cnt[6]), .B(n_82), .Z(O0[6]), .CO(n_84));
	notech_ha2 i_5(.A(fsm5_cnt[5]), .B(n_80), .Z(O0[5]), .CO(n_82));
	notech_ha2 i_4(.A(fsm5_cnt[4]), .B(n_78), .Z(O0[4]), .CO(n_80));
	notech_ha2 i_3(.A(fsm5_cnt[3]), .B(n_76), .Z(O0[3]), .CO(n_78));
	notech_ha2 i_2(.A(fsm5_cnt[2]), .B(n_74), .Z(O0[2]), .CO(n_76));
	notech_ha2 i_1(.A(fsm5_cnt[1]), .B(fsm5_cnt[0]), .Z(O0[1]), .CO(n_74));
	notech_inv i_0(.A(fsm5_cnt[0]), .Z(O0[0]));
endmodule
module cmp14_0(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_10(.A(inb[2]), .B(ina[2]), .Z(n_34));
	notech_xor2 i_9(.A(inb[4]), .B(ina[4]), .Z(n_33));
	notech_xor2 i_8(.A(inb[6]), .B(ina[6]), .Z(n_32));
	notech_xor2 i_6(.A(inb[3]), .B(ina[3]), .Z(n_31));
	notech_xor2 i_5(.A(inb[5]), .B(ina[5]), .Z(n_30));
	notech_xor2 i_4(.A(inb[7]), .B(ina[7]), .Z(n_29));
	notech_xor2 i_0(.A(inb[9]), .B(ina[9]), .Z(n_55));
	notech_xor2 i_1(.A(inb[8]), .B(ina[8]), .Z(n_56));
	notech_xor2 i_3(.A(inb[1]), .B(ina[1]), .Z(n_57));
	notech_xor2 i_7(.A(inb[0]), .B(ina[0]), .Z(n_58));
	notech_or4 i_38(.A(n_57), .B(n_56), .C(n_55), .D(ina[13]), .Z(n_61));
	notech_or4 i_37(.A(n_34), .B(n_31), .C(n_33), .D(n_30), .Z(n_66));
	notech_or4 i_39(.A(n_32), .B(n_29), .C(n_58), .D(n_66), .Z(n_67));
	notech_nor2 i_2(.A(n_67), .B(n_61), .Z(out));
endmodule
module cmp14_1(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_10(.A(inb[2]), .B(ina[2]), .Z(n_34));
	notech_xor2 i_9(.A(inb[4]), .B(ina[4]), .Z(n_33));
	notech_xor2 i_8(.A(inb[6]), .B(ina[6]), .Z(n_32));
	notech_xor2 i_6(.A(inb[3]), .B(ina[3]), .Z(n_31));
	notech_xor2 i_5(.A(inb[5]), .B(ina[5]), .Z(n_30));
	notech_xor2 i_4(.A(inb[7]), .B(ina[7]), .Z(n_29));
	notech_xor2 i_0(.A(inb[9]), .B(ina[9]), .Z(n_55));
	notech_xor2 i_1(.A(inb[8]), .B(ina[8]), .Z(n_56));
	notech_xor2 i_3(.A(inb[1]), .B(ina[1]), .Z(n_57));
	notech_xor2 i_7(.A(inb[0]), .B(ina[0]), .Z(n_58));
	notech_or4 i_38(.A(n_57), .B(n_56), .C(n_55), .D(ina[13]), .Z(n_61));
	notech_or4 i_37(.A(n_34), .B(n_31), .C(n_33), .D(n_30), .Z(n_66));
	notech_or4 i_39(.A(n_32), .B(n_29), .C(n_58), .D(n_66), .Z(n_67));
	notech_nor2 i_2(.A(n_67), .B(n_61), .Z(out));
endmodule
module cmp14_2(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out297031));
	notech_inv i_15292(.A(out297031), .Z(out2));
endmodule
module cmp14_3(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out297030));
	notech_inv i_15273(.A(out297030), .Z(out2));
endmodule
module cmp14_4(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out297029));
	notech_inv i_15254(.A(out297029), .Z(out2));
endmodule
module cmp14_5(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out297028));
	notech_inv i_15235(.A(out297028), .Z(out2));
endmodule
module cmp14_6(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out297027));
	notech_inv i_15216(.A(out297027), .Z(out2));
endmodule
module cmp14_7(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out297026));
	notech_inv i_15197(.A(out297026), .Z(out2));
endmodule
module cmp14_8(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out297025));
	notech_inv i_15178(.A(out297025), .Z(out2));
endmodule
module cmp14_9(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_nand2 i_41(.A(ina[10]), .B(n_63), .Z(n_62));
	notech_or2 i_0(.A(ina[12]), .B(inb[12]), .Z(n_63));
	notech_nand2 i_1(.A(inb[10]), .B(n_62), .Z(n_64));
	notech_xor2 i_26(.A(inb[5]), .B(ina[5]), .Z(n_65));
	notech_xor2 i_27(.A(inb[4]), .B(ina[4]), .Z(n_66));
	notech_xor2 i_28(.A(inb[3]), .B(ina[3]), .Z(n_68));
	notech_xor2 i_29(.A(inb[2]), .B(ina[2]), .Z(n_69));
	notech_or4 i_39(.A(n_69), .B(n_68), .C(n_66), .D(n_65), .Z(n_71));
	notech_xor2 i_30(.A(inb[1]), .B(ina[1]), .Z(n_72));
	notech_xor2 i_31(.A(inb[0]), .B(ina[0]), .Z(n_73));
	notech_xor2 i_22(.A(inb[9]), .B(ina[9]), .Z(n_75));
	notech_xor2 i_23(.A(inb[8]), .B(ina[8]), .Z(n_76));
	notech_xor2 i_24(.A(inb[7]), .B(ina[7]), .Z(n_78));
	notech_xor2 i_25(.A(inb[6]), .B(ina[6]), .Z(n_79));
	notech_or4 i_38(.A(n_79), .B(n_78), .C(n_76), .D(n_75), .Z(n_81));
	notech_ao3 i_216(.A(n_64), .B(out2), .C(ina[13]), .Z(out));
	notech_or4 i_32(.A(n_73), .B(n_72), .C(n_81), .D(n_71), .Z(out297024));
	notech_inv i_15159(.A(out297024), .Z(out2));
endmodule
module Dtlb(clk, rstn, addr_phys, cr3, cr0, data_miss, iDaddr, pg_en, iwrite_data
		, owrite_data, iread_req, iread_ack, iwrite_req, iwrite_ack, iread_sz
		, oread_sz, iwrite_sz, owrite_sz, oread_req, oread_ack, owrite_req
		, owrite_ack, pg_fault, wr_fault, cr2, flush_tlb, cs, pt_fault, busy_ram
		, outstanding);

	input clk;
	input rstn;
	output [31:0] addr_phys;
	input [31:0] cr3;
	input [31:0] cr0;
	input [31:0] data_miss;
	input [31:0] iDaddr;
	input pg_en;
	input [31:0] iwrite_data;
	output [31:0] owrite_data;
	input iread_req;
	input iread_ack;
	input iwrite_req;
	input iwrite_ack;
	input [1:0] iread_sz;
	output [1:0] oread_sz;
	input [1:0] iwrite_sz;
	output [1:0] owrite_sz;
	output oread_req;
	output oread_ack;
	output owrite_req;
	output owrite_ack;
	output pg_fault;
	output wr_fault;
	output [31:0] cr2;
	input flush_tlb;
	input [31:0] cs;
	output pt_fault;
	input busy_ram;
	output outstanding;

	wire [3:0] fsm;
	wire [31:0] addr_miss;
	wire [31:0] wrA;
	wire [31:0] iDaddr_f;
	wire [31:0] wrD;
	wire [1:0] nx_dir;
	wire [8:0] fsm5_cnt_0;
	wire [8:0] fsm5_cnt;



	notech_inv i_15444(.A(n_61750), .Z(n_61777));
	notech_inv i_15443(.A(n_61750), .Z(n_61776));
	notech_inv i_15442(.A(n_61750), .Z(n_61775));
	notech_inv i_15440(.A(n_61750), .Z(n_61773));
	notech_inv i_15439(.A(n_61750), .Z(n_61772));
	notech_inv i_15438(.A(n_61750), .Z(n_61771));
	notech_inv i_15435(.A(n_61750), .Z(n_61768));
	notech_inv i_15434(.A(n_61750), .Z(n_61767));
	notech_inv i_15433(.A(n_61750), .Z(n_61766));
	notech_inv i_15431(.A(n_61750), .Z(n_61764));
	notech_inv i_15429(.A(n_61750), .Z(n_61763));
	notech_inv i_15428(.A(n_61750), .Z(n_61762));
	notech_inv i_15425(.A(n_61750), .Z(n_61759));
	notech_inv i_15424(.A(n_61750), .Z(n_61758));
	notech_inv i_15423(.A(n_61750), .Z(n_61757));
	notech_inv i_15420(.A(n_61750), .Z(n_61755));
	notech_inv i_15419(.A(n_61750), .Z(n_61754));
	notech_inv i_15418(.A(n_61750), .Z(n_61753));
	notech_inv i_15415(.A(clk), .Z(n_61750));
	notech_inv i_15413(.A(n_61722), .Z(n_61749));
	notech_inv i_15412(.A(n_61722), .Z(n_61748));
	notech_inv i_15411(.A(n_61722), .Z(n_61747));
	notech_inv i_15409(.A(n_61722), .Z(n_61745));
	notech_inv i_15408(.A(n_61722), .Z(n_61744));
	notech_inv i_15407(.A(n_61722), .Z(n_61743));
	notech_inv i_15403(.A(n_61722), .Z(n_61740));
	notech_inv i_15402(.A(n_61722), .Z(n_61739));
	notech_inv i_15401(.A(n_61722), .Z(n_61738));
	notech_inv i_15399(.A(n_61722), .Z(n_61736));
	notech_inv i_15397(.A(n_61722), .Z(n_61735));
	notech_inv i_15396(.A(n_61722), .Z(n_61734));
	notech_inv i_15393(.A(n_61722), .Z(n_61731));
	notech_inv i_15392(.A(n_61722), .Z(n_61730));
	notech_inv i_15391(.A(n_61722), .Z(n_61729));
	notech_inv i_15388(.A(n_61722), .Z(n_61727));
	notech_inv i_15387(.A(n_61722), .Z(n_61726));
	notech_inv i_15386(.A(n_61722), .Z(n_61725));
	notech_inv i_15383(.A(clk), .Z(n_61722));
	notech_inv i_15381(.A(n_61694), .Z(n_61721));
	notech_inv i_15380(.A(n_61694), .Z(n_61720));
	notech_inv i_15379(.A(n_61694), .Z(n_61719));
	notech_inv i_15377(.A(n_61694), .Z(n_61717));
	notech_inv i_15376(.A(n_61694), .Z(n_61716));
	notech_inv i_15375(.A(n_61694), .Z(n_61715));
	notech_inv i_15371(.A(n_61694), .Z(n_61712));
	notech_inv i_15370(.A(n_61694), .Z(n_61711));
	notech_inv i_15369(.A(n_61694), .Z(n_61710));
	notech_inv i_15367(.A(n_61694), .Z(n_61708));
	notech_inv i_15365(.A(n_61694), .Z(n_61707));
	notech_inv i_15364(.A(n_61694), .Z(n_61706));
	notech_inv i_15361(.A(n_61694), .Z(n_61703));
	notech_inv i_15359(.A(n_61694), .Z(n_61701));
	notech_inv i_15355(.A(n_61694), .Z(n_61698));
	notech_inv i_15354(.A(n_61694), .Z(n_61697));
	notech_inv i_15351(.A(clk), .Z(n_61694));
	notech_inv i_15263(.A(n_61598), .Z(n_61605));
	notech_inv i_15262(.A(n_61598), .Z(n_61604));
	notech_inv i_15257(.A(n_61598), .Z(n_61599));
	notech_inv i_15256(.A(pg_en), .Z(n_61598));
	notech_inv i_14437(.A(n_61053), .Z(n_61080));
	notech_inv i_14436(.A(n_61053), .Z(n_61079));
	notech_inv i_14435(.A(n_61053), .Z(n_61078));
	notech_inv i_14433(.A(n_61053), .Z(n_61076));
	notech_inv i_14432(.A(n_61053), .Z(n_61075));
	notech_inv i_14431(.A(n_61053), .Z(n_61074));
	notech_inv i_14428(.A(n_61053), .Z(n_61071));
	notech_inv i_14427(.A(n_61053), .Z(n_61070));
	notech_inv i_14426(.A(n_61053), .Z(n_61069));
	notech_inv i_14424(.A(n_61053), .Z(n_61067));
	notech_inv i_14423(.A(n_61053), .Z(n_61066));
	notech_inv i_14422(.A(n_61053), .Z(n_61065));
	notech_inv i_14419(.A(n_61053), .Z(n_61062));
	notech_inv i_14418(.A(n_61053), .Z(n_61061));
	notech_inv i_14417(.A(n_61053), .Z(n_61060));
	notech_inv i_14415(.A(n_61053), .Z(n_61058));
	notech_inv i_14414(.A(n_61053), .Z(n_61057));
	notech_inv i_14413(.A(n_61053), .Z(n_61056));
	notech_inv i_14410(.A(rstn), .Z(n_61053));
	notech_inv i_14409(.A(n_61025), .Z(n_61052));
	notech_inv i_14408(.A(n_61025), .Z(n_61051));
	notech_inv i_14407(.A(n_61025), .Z(n_61050));
	notech_inv i_14405(.A(n_61025), .Z(n_61048));
	notech_inv i_14404(.A(n_61025), .Z(n_61047));
	notech_inv i_14403(.A(n_61025), .Z(n_61046));
	notech_inv i_14400(.A(n_61025), .Z(n_61043));
	notech_inv i_14399(.A(n_61025), .Z(n_61042));
	notech_inv i_14398(.A(n_61025), .Z(n_61041));
	notech_inv i_14396(.A(n_61025), .Z(n_61039));
	notech_inv i_14395(.A(n_61025), .Z(n_61038));
	notech_inv i_14394(.A(n_61025), .Z(n_61037));
	notech_inv i_14391(.A(n_61025), .Z(n_61034));
	notech_inv i_14390(.A(n_61025), .Z(n_61033));
	notech_inv i_14389(.A(n_61025), .Z(n_61032));
	notech_inv i_14387(.A(n_61025), .Z(n_61030));
	notech_inv i_14386(.A(n_61025), .Z(n_61029));
	notech_inv i_14385(.A(n_61025), .Z(n_61028));
	notech_inv i_14382(.A(rstn), .Z(n_61025));
	notech_inv i_14381(.A(n_60997), .Z(n_61024));
	notech_inv i_14380(.A(n_60997), .Z(n_61023));
	notech_inv i_14379(.A(n_60997), .Z(n_61022));
	notech_inv i_14377(.A(n_60997), .Z(n_61020));
	notech_inv i_14376(.A(n_60997), .Z(n_61019));
	notech_inv i_14375(.A(n_60997), .Z(n_61018));
	notech_inv i_14372(.A(n_60997), .Z(n_61015));
	notech_inv i_14371(.A(n_60997), .Z(n_61014));
	notech_inv i_14370(.A(n_60997), .Z(n_61013));
	notech_inv i_14368(.A(n_60997), .Z(n_61011));
	notech_inv i_14367(.A(n_60997), .Z(n_61010));
	notech_inv i_14366(.A(n_60997), .Z(n_61009));
	notech_inv i_14363(.A(n_60997), .Z(n_61006));
	notech_inv i_14361(.A(n_60997), .Z(n_61004));
	notech_inv i_14358(.A(n_60997), .Z(n_61001));
	notech_inv i_14357(.A(n_60997), .Z(n_61000));
	notech_inv i_14354(.A(rstn), .Z(n_60997));
	notech_inv i_12124(.A(n_58635), .Z(n_58636));
	notech_inv i_12123(.A(fsm[0]), .Z(n_58635));
	notech_inv i_12116(.A(n_58626), .Z(n_58627));
	notech_inv i_12115(.A(n_948), .Z(n_58626));
	notech_inv i_12108(.A(n_58617), .Z(n_58618));
	notech_inv i_12107(.A(hit_tab21), .Z(n_58617));
	notech_inv i_12100(.A(n_58608), .Z(n_58609));
	notech_inv i_12099(.A(\hit_dir1[7] ), .Z(n_58608));
	notech_inv i_12092(.A(n_58599), .Z(n_58600));
	notech_inv i_12091(.A(hit_tab11), .Z(n_58599));
	notech_inv i_8840(.A(n_54824), .Z(n_54825));
	notech_inv i_8839(.A(\nbus_14033[0] ), .Z(n_54824));
	notech_inv i_8832(.A(n_54815), .Z(n_54816));
	notech_inv i_8831(.A(n_1043), .Z(n_54815));
	notech_inv i_8824(.A(n_54806), .Z(n_54807));
	notech_inv i_8823(.A(n_13460), .Z(n_54806));
	notech_inv i_8814(.A(n_54795), .Z(n_54796));
	notech_inv i_8813(.A(n_1040), .Z(n_54795));
	notech_inv i_8697(.A(n_54647), .Z(n_54648));
	notech_inv i_8696(.A(\nbus_14043[0] ), .Z(n_54647));
	notech_inv i_8678(.A(n_54627), .Z(n_54628));
	notech_inv i_8677(.A(n_13488), .Z(n_54627));
	notech_inv i_8670(.A(n_54618), .Z(n_54619));
	notech_inv i_8669(.A(\nbus_14037[0] ), .Z(n_54618));
	notech_inv i_8665(.A(n_54607), .Z(n_54613));
	notech_inv i_8660(.A(n_54607), .Z(n_54608));
	notech_inv i_8659(.A(n_52575), .Z(n_54607));
	notech_inv i_8652(.A(n_54598), .Z(n_54599));
	notech_inv i_8651(.A(\nbus_14028[0] ), .Z(n_54598));
	notech_inv i_8644(.A(n_54589), .Z(n_54590));
	notech_inv i_8643(.A(\nbus_14036[0] ), .Z(n_54589));
	notech_inv i_8636(.A(n_54580), .Z(n_54581));
	notech_inv i_8635(.A(\nbus_14017[0] ), .Z(n_54580));
	notech_inv i_8626(.A(n_54569), .Z(n_54570));
	notech_inv i_8625(.A(\nbus_14042[0] ), .Z(n_54569));
	notech_inv i_8618(.A(n_54560), .Z(n_54561));
	notech_inv i_8617(.A(\nbus_14035[0] ), .Z(n_54560));
	notech_inv i_8610(.A(n_54551), .Z(n_54552));
	notech_inv i_8609(.A(\nbus_14034[0] ), .Z(n_54551));
	notech_inv i_8602(.A(n_54542), .Z(n_54543));
	notech_inv i_8601(.A(\nbus_14015[0] ), .Z(n_54542));
	notech_inv i_8594(.A(n_54533), .Z(n_54534));
	notech_inv i_8593(.A(\nbus_14016[0] ), .Z(n_54533));
	notech_inv i_7767(.A(n_53620), .Z(n_53621));
	notech_inv i_7766(.A(n_656), .Z(n_53620));
	notech_inv i_7715(.A(n_53472), .Z(n_53478));
	notech_inv i_7710(.A(n_53472), .Z(n_53473));
	notech_inv i_7709(.A(n_1042), .Z(n_53472));
	notech_inv i_7707(.A(n_1085), .Z(n_53469));
	notech_inv i_7706(.A(n_1085), .Z(n_53468));
	notech_inv i_7702(.A(n_1085), .Z(n_53464));
	notech_inv i_7694(.A(n_53454), .Z(n_53455));
	notech_inv i_7693(.A(n_1098), .Z(n_53454));
	notech_inv i_7686(.A(n_53445), .Z(n_53446));
	notech_inv i_7685(.A(n_1081), .Z(n_53445));
	notech_inv i_7683(.A(\nbus_14013[0] ), .Z(n_53369));
	notech_inv i_7681(.A(\nbus_14013[0] ), .Z(n_53367));
	notech_inv i_7678(.A(\nbus_14013[0] ), .Z(n_53364));
	notech_inv i_7676(.A(\nbus_14013[0] ), .Z(n_53362));
	notech_xor2 i_149(.A(n_13608), .B(\nnx_tab2[0] ), .Z(n_573));
	notech_or4 i_139(.A(hit_adr23), .B(hit_adr24), .C(hit_adr22), .D(hit_adr21
		), .Z(n_571));
	notech_ao4 i_148(.A(hit_adr22), .B(n_1024), .C(n_13613), .D(n_1025), .Z(n_564
		));
	notech_nor2 i_96(.A(hit_adr24), .B(\nx_tab2[0] ), .Z(n_562));
	notech_nor2 i_607(.A(hit_adr23), .B(n_562), .Z(n_561));
	notech_nor2 i_147(.A(hit_adr22), .B(n_561), .Z(n_559));
	notech_nand3 i_604(.A(n_13466), .B(n_13538), .C(n_13536), .Z(n_557));
	notech_or2 i_79(.A(fsm5_cnt[2]), .B(fsm5_cnt[3]), .Z(n_556));
	notech_and3 i_603(.A(fsm5_cnt[4]), .B(fsm5_cnt[5]), .C(n_556), .Z(n_555)
		);
	notech_or2 i_153(.A(fsm5_cnt[6]), .B(n_555), .Z(n_554));
	notech_and2 i_602(.A(fsm5_cnt[7]), .B(n_554), .Z(n_553));
	notech_or4 i_601(.A(fsm5_cnt[8]), .B(n_1028), .C(n_553), .D(n_13783), .Z
		(n_552));
	notech_ao3 i_75612(.A(data_miss[5]), .B(n_960), .C(n_972), .Z(n_550));
	notech_ao3 i_596(.A(n_995), .B(n_13464), .C(n_550), .Z(n_549));
	notech_or4 i_145(.A(hit_dir2), .B(\hit_dir1[7] ), .C(n_972), .D(busy_ram
		), .Z(n_547));
	notech_ao4 i_144(.A(n_13617), .B(n_13616), .C(fsm[0]), .D(n_13618), .Z(n_546
		));
	notech_or4 i_589(.A(fsm[2]), .B(fsm[1]), .C(n_1015), .D(n_13783), .Z(n_545
		));
	notech_xor2 i_143(.A(fsm[0]), .B(iwrite_ack), .Z(n_541));
	notech_nao3 i_142(.A(n_1043), .B(n_947), .C(n_946), .Z(n_538));
	notech_ao4 i_141(.A(iwrite_req), .B(n_61605), .C(n_946), .D(n_1053), .Z(n_536
		));
	notech_nao3 i_575(.A(n_13460), .B(\dir2[29] ), .C(\hit_dir1[7] ), .Z(n_534
		));
	notech_nao3 i_572(.A(n_13460), .B(\dir2[28] ), .C(\hit_dir1[7] ), .Z(n_533
		));
	notech_nao3 i_568(.A(n_13460), .B(\dir2[27] ), .C(\hit_dir1[7] ), .Z(n_532
		));
	notech_nao3 i_565(.A(n_13460), .B(\dir2[26] ), .C(\hit_dir1[7] ), .Z(n_531
		));
	notech_nao3 i_562(.A(n_13460), .B(\dir2[25] ), .C(\hit_dir1[7] ), .Z(n_530
		));
	notech_nao3 i_559(.A(n_13460), .B(\dir2[24] ), .C(\hit_dir1[7] ), .Z(n_529
		));
	notech_nao3 i_556(.A(n_13460), .B(\dir2[23] ), .C(\hit_dir1[7] ), .Z(n_528
		));
	notech_nao3 i_553(.A(n_13460), .B(\dir2[22] ), .C(\hit_dir1[7] ), .Z(n_527
		));
	notech_nao3 i_550(.A(n_13460), .B(\dir2[21] ), .C(\hit_dir1[7] ), .Z(n_526
		));
	notech_nao3 i_547(.A(n_13460), .B(\dir2[20] ), .C(\hit_dir1[7] ), .Z(n_525
		));
	notech_nao3 i_544(.A(n_13460), .B(\dir2[19] ), .C(\hit_dir1[7] ), .Z(n_524
		));
	notech_nao3 i_541(.A(n_54807), .B(\dir2[18] ), .C(\hit_dir1[7] ), .Z(n_523
		));
	notech_nao3 i_538(.A(n_54807), .B(\dir2[17] ), .C(\hit_dir1[7] ), .Z(n_522
		));
	notech_nao3 i_535(.A(n_54807), .B(\dir2[16] ), .C(n_58609), .Z(n_521));
	notech_nao3 i_532(.A(n_54807), .B(\dir2[15] ), .C(n_58609), .Z(n_520));
	notech_nao3 i_529(.A(n_54807), .B(\dir2[14] ), .C(n_58609), .Z(n_519));
	notech_nao3 i_526(.A(n_54807), .B(\dir2[13] ), .C(n_58609), .Z(n_518));
	notech_nao3 i_523(.A(n_54807), .B(\dir2[12] ), .C(n_58609), .Z(n_517));
	notech_nao3 i_520(.A(n_13460), .B(\dir2[11] ), .C(n_58609), .Z(n_516));
	notech_nao3 i_517(.A(\dir2[10] ), .B(n_54807), .C(n_58609), .Z(n_515));
	notech_nand3 i_494(.A(n_52185), .B(iread_ack), .C(n_61605), .Z(n_494));
	notech_nao3 i_491(.A(n_406), .B(n_13461), .C(req_miss), .Z(n_491));
	notech_xor2 i_140(.A(iread_req), .B(iread_ack), .Z(n_490));
	notech_nand3 i_257(.A(n_61605), .B(n_13463), .C(wrA[11]), .Z(n_487));
	notech_and2 i_18(.A(n_61605), .B(n_1080), .Z(n_486));
	notech_nand3 i_254(.A(n_61605), .B(n_13463), .C(wrA[10]), .Z(n_485));
	notech_nand3 i_251(.A(n_61605), .B(n_13463), .C(wrA[9]), .Z(n_484));
	notech_nand3 i_248(.A(n_61604), .B(n_13463), .C(wrA[8]), .Z(n_483));
	notech_nand3 i_245(.A(n_61604), .B(n_13463), .C(wrA[7]), .Z(n_482));
	notech_nand3 i_242(.A(n_61604), .B(n_13463), .C(wrA[6]), .Z(n_481));
	notech_nand3 i_239(.A(n_61604), .B(n_13463), .C(wrA[5]), .Z(n_480));
	notech_nand3 i_236(.A(n_61604), .B(n_13463), .C(wrA[4]), .Z(n_479));
	notech_nand3 i_233(.A(n_61604), .B(n_13463), .C(wrA[3]), .Z(n_478));
	notech_nand3 i_230(.A(n_61605), .B(n_13463), .C(wrA[2]), .Z(n_477));
	notech_nand3 i_227(.A(n_61605), .B(n_13463), .C(wrA[1]), .Z(n_476));
	notech_nand3 i_224(.A(n_61605), .B(wrA[0]), .C(n_13463), .Z(n_475));
	notech_and4 i_221(.A(n_995), .B(n_13464), .C(iread_ack), .D(n_61605), .Z
		(n_474));
	notech_ao3 i_220(.A(n_61605), .B(n_1030), .C(n_1028), .Z(n_473));
	notech_nand2 i_146(.A(n_1032), .B(n_13618), .Z(n_408));
	notech_nand2 i_137(.A(n_986), .B(n_61605), .Z(n_407));
	notech_nand3 i_82(.A(n_983), .B(iread_req), .C(n_13513), .Z(n_406));
	notech_or4 i_619(.A(n_1001), .B(n_1002), .C(n_13611), .D(n_13613), .Z(n_577
		));
	notech_or4 i_620(.A(n_1001), .B(n_1002), .C(n_13613), .D(\nx_tab2[0] ), 
		.Z(n_578));
	notech_or4 i_621(.A(n_1001), .B(n_1002), .C(n_13611), .D(\nx_tab2[1] ), 
		.Z(n_579));
	notech_or4 i_138(.A(hit_adr13), .B(hit_adr14), .C(hit_adr12), .D(hit_adr11
		), .Z(n_583));
	notech_xor2 i_150(.A(n_13542), .B(\nnx_tab1[0] ), .Z(n_585));
	notech_nor2 i_151(.A(hit_adr12), .B(n_592), .Z(n_590));
	notech_nor2 i_631(.A(hit_adr13), .B(n_593), .Z(n_592));
	notech_nor2 i_128(.A(hit_adr14), .B(\nx_tab1[0] ), .Z(n_593));
	notech_ao4 i_152(.A(hit_adr12), .B(n_1018), .C(n_13538), .D(n_1019), .Z(n_595
		));
	notech_nand3 i_636(.A(n_13466), .B(\nx_tab1[1] ), .C(\nx_tab1[0] ), .Z(n_599
		));
	notech_nand3 i_637(.A(n_13466), .B(\nx_tab1[1] ), .C(n_13536), .Z(n_600)
		);
	notech_nand3 i_638(.A(\nx_tab1[0] ), .B(n_13538), .C(n_13466), .Z(n_601)
		);
	notech_or4 i_641(.A(n_1001), .B(n_1002), .C(\nx_tab2[1] ), .D(\nx_tab2[0] 
		), .Z(n_604));
	notech_nao3 i_642(.A(iwrite_req), .B(n_606), .C(data_miss[1]), .Z(n_605)
		);
	notech_nao3 i_92(.A(n_13755), .B(n_13756), .C(cs[0]), .Z(n_606));
	notech_or4 i_661(.A(data_miss[0]), .B(n_989), .C(n_13784), .D(n_13783), 
		.Z(n_625));
	notech_nor2 i_70(.A(nx_dir[0]), .B(nx_dir[1]), .Z(n_627));
	notech_and3 i_663(.A(n_61605), .B(n_13513), .C(flush_tlb), .Z(n_628));
	notech_nand2 i_667(.A(n_627), .B(n_13757), .Z(n_631));
	notech_and2 i_689(.A(n_58609), .B(n_653), .Z(n_652));
	notech_or4 i_154(.A(hit_tab12), .B(hit_tab11), .C(hit_tab13), .D(hit_tab14
		), .Z(n_653));
	notech_and2 i_690(.A(hit_dir2), .B(n_655), .Z(n_654));
	notech_or4 i_155(.A(hit_tab22), .B(hit_tab24), .C(hit_tab21), .D(hit_tab23
		), .Z(n_655));
	notech_nand3 i_90(.A(iread_ack), .B(n_61605), .C(n_13614), .Z(n_656));
	notech_ao3 i_789(.A(n_974), .B(n_999), .C(data_miss[1]), .Z(n_657));
	notech_nand3 i_271(.A(n_53469), .B(\tab13[10] ), .C(n_1096), .Z(n_686)
		);
	notech_nand3 i_264(.A(hit_tab11), .B(\tab11[10] ), .C(n_53468), .Z(n_689
		));
	notech_nao3 i_260(.A(hit_tab21), .B(\tab21[10] ), .C(n_1081), .Z(n_692)
		);
	notech_nand3 i_286(.A(n_53469), .B(n_1096), .C(\tab13[11] ), .Z(n_697)
		);
	notech_nand3 i_283(.A(hit_tab11), .B(n_53469), .C(\tab11[11] ), .Z(n_700
		));
	notech_nao3 i_280(.A(hit_tab21), .B(\tab21[11] ), .C(n_1081), .Z(n_703)
		);
	notech_nand3 i_297(.A(n_53469), .B(n_1096), .C(\tab13[12] ), .Z(n_708)
		);
	notech_nand3 i_294(.A(hit_tab11), .B(n_53468), .C(\tab11[12] ), .Z(n_711
		));
	notech_nao3 i_291(.A(hit_tab21), .B(\tab21[12] ), .C(n_1081), .Z(n_714)
		);
	notech_nand3 i_308(.A(n_53468), .B(n_1096), .C(\tab13[13] ), .Z(n_719)
		);
	notech_nand3 i_305(.A(hit_tab11), .B(n_53468), .C(\tab11[13] ), .Z(n_722
		));
	notech_nao3 i_302(.A(hit_tab21), .B(\tab21[13] ), .C(n_1081), .Z(n_725)
		);
	notech_nand3 i_319(.A(n_53468), .B(n_1096), .C(\tab13[14] ), .Z(n_730)
		);
	notech_nand3 i_316(.A(hit_tab11), .B(n_53468), .C(\tab11[14] ), .Z(n_733
		));
	notech_nao3 i_313(.A(hit_tab21), .B(\tab21[14] ), .C(n_1081), .Z(n_736)
		);
	notech_nand3 i_330(.A(n_53469), .B(n_1096), .C(\tab13[15] ), .Z(n_741)
		);
	notech_nand3 i_327(.A(hit_tab11), .B(n_53469), .C(\tab11[15] ), .Z(n_744
		));
	notech_nao3 i_324(.A(hit_tab21), .B(\tab21[15] ), .C(n_1081), .Z(n_747)
		);
	notech_nand3 i_341(.A(n_53469), .B(n_1096), .C(\tab13[16] ), .Z(n_752)
		);
	notech_nand3 i_338(.A(hit_tab11), .B(n_53469), .C(\tab11[16] ), .Z(n_755
		));
	notech_nao3 i_335(.A(hit_tab21), .B(\tab21[16] ), .C(n_1081), .Z(n_758)
		);
	notech_nand3 i_352(.A(n_53469), .B(n_1096), .C(\tab13[17] ), .Z(n_763)
		);
	notech_nand3 i_349(.A(hit_tab11), .B(n_53469), .C(\tab11[17] ), .Z(n_766
		));
	notech_nao3 i_346(.A(hit_tab21), .B(\tab21[17] ), .C(n_1081), .Z(n_769)
		);
	notech_nand3 i_363(.A(n_53469), .B(n_1096), .C(\tab13[18] ), .Z(n_774)
		);
	notech_nand3 i_360(.A(hit_tab11), .B(n_53469), .C(\tab11[18] ), .Z(n_777
		));
	notech_nao3 i_357(.A(hit_tab21), .B(\tab21[18] ), .C(n_1081), .Z(n_780)
		);
	notech_nand3 i_374(.A(n_53469), .B(n_1096), .C(\tab13[19] ), .Z(n_785)
		);
	notech_nand3 i_371(.A(hit_tab11), .B(n_53469), .C(\tab11[19] ), .Z(n_788
		));
	notech_nao3 i_368(.A(hit_tab21), .B(\tab21[19] ), .C(n_1081), .Z(n_791)
		);
	notech_nand3 i_385(.A(n_53468), .B(n_1096), .C(\tab13[20] ), .Z(n_796)
		);
	notech_nand3 i_382(.A(hit_tab11), .B(n_53464), .C(\tab11[20] ), .Z(n_799
		));
	notech_nao3 i_379(.A(hit_tab21), .B(\tab21[20] ), .C(n_1081), .Z(n_802)
		);
	notech_nand3 i_396(.A(n_53464), .B(n_1096), .C(\tab13[21] ), .Z(n_807)
		);
	notech_nand3 i_393(.A(n_58600), .B(n_53464), .C(\tab11[21] ), .Z(n_810)
		);
	notech_nao3 i_390(.A(n_58618), .B(\tab21[21] ), .C(n_1081), .Z(n_813));
	notech_nand3 i_407(.A(n_53464), .B(n_1096), .C(\tab13[22] ), .Z(n_818)
		);
	notech_nand3 i_404(.A(n_58600), .B(n_53464), .C(\tab11[22] ), .Z(n_821)
		);
	notech_nao3 i_401(.A(n_58618), .B(\tab21[22] ), .C(n_53446), .Z(n_824)
		);
	notech_nand3 i_418(.A(n_53464), .B(n_1096), .C(\tab13[23] ), .Z(n_829)
		);
	notech_nand3 i_415(.A(n_58600), .B(n_53464), .C(\tab11[23] ), .Z(n_832)
		);
	notech_nao3 i_412(.A(n_58618), .B(\tab21[23] ), .C(n_53446), .Z(n_835)
		);
	notech_nand3 i_429(.A(n_53464), .B(n_1096), .C(\tab13[24] ), .Z(n_840)
		);
	notech_nand3 i_426(.A(n_58600), .B(n_53464), .C(\tab11[24] ), .Z(n_843)
		);
	notech_nao3 i_423(.A(n_58618), .B(\tab21[24] ), .C(n_53446), .Z(n_846)
		);
	notech_nand3 i_440(.A(n_53464), .B(n_1096), .C(\tab13[25] ), .Z(n_851)
		);
	notech_nand3 i_437(.A(n_58600), .B(n_53468), .C(\tab11[25] ), .Z(n_854)
		);
	notech_nao3 i_434(.A(n_58618), .B(\tab21[25] ), .C(n_53446), .Z(n_857)
		);
	notech_nand3 i_451(.A(n_53468), .B(n_1096), .C(\tab13[26] ), .Z(n_862)
		);
	notech_nand3 i_448(.A(n_58600), .B(n_53468), .C(\tab11[26] ), .Z(n_865)
		);
	notech_nao3 i_445(.A(n_58618), .B(\tab21[26] ), .C(n_53446), .Z(n_868)
		);
	notech_nand3 i_462(.A(n_53468), .B(n_1096), .C(\tab13[27] ), .Z(n_873)
		);
	notech_nand3 i_459(.A(n_58600), .B(n_53468), .C(\tab11[27] ), .Z(n_876)
		);
	notech_nao3 i_456(.A(n_58618), .B(\tab21[27] ), .C(n_53446), .Z(n_879)
		);
	notech_nand3 i_473(.A(n_53464), .B(n_1096), .C(\tab13[28] ), .Z(n_884)
		);
	notech_nand3 i_470(.A(n_58600), .B(n_53464), .C(\tab11[28] ), .Z(n_887)
		);
	notech_nao3 i_467(.A(n_58618), .B(\tab21[28] ), .C(n_53446), .Z(n_890)
		);
	notech_nand3 i_484(.A(n_53464), .B(n_1096), .C(\tab13[29] ), .Z(n_895)
		);
	notech_nand3 i_481(.A(n_58600), .B(n_53468), .C(\tab11[29] ), .Z(n_898)
		);
	notech_nao3 i_478(.A(n_58618), .B(\tab21[29] ), .C(n_53446), .Z(n_901)
		);
	notech_and2 i_983(.A(iwrite_sz[0]), .B(n_53478), .Z(n_902));
	notech_and2 i_984(.A(iwrite_sz[1]), .B(n_53478), .Z(n_903));
	notech_nao3 i_489(.A(n_61605), .B(n_1077), .C(iread_ack), .Z(n_904));
	notech_nand2 i_490(.A(n_490), .B(n_13783), .Z(n_905));
	notech_and3 i_84(.A(n_983), .B(iwrite_req), .C(n_13513), .Z(n_946));
	notech_nand2 i_580(.A(iwrite_req), .B(n_1053), .Z(n_947));
	notech_or4 i_91(.A(fsm[0]), .B(fsm[2]), .C(fsm[1]), .D(fsm[3]), .Z(n_948
		));
	notech_and4 i_583(.A(n_13464), .B(n_988), .C(data_miss[0]), .D(data_miss
		[5]), .Z(n_951));
	notech_or4 i_586(.A(n_954), .B(n_992), .C(n_972), .D(n_1005), .Z(n_952)
		);
	notech_or4 i_587(.A(fsm[2]), .B(fsm[1]), .C(n_13618), .D(n_13783), .Z(n_953
		));
	notech_ao4 i_67(.A(hit_dir2), .B(n_58609), .C(pg_fault), .D(n_983), .Z(n_954
		));
	notech_nao3 i_592(.A(n_547), .B(n_13464), .C(n_984), .Z(n_957));
	notech_or2 i_597(.A(iread_req), .B(data_miss[6]), .Z(n_960));
	notech_and2 i_1021(.A(iwrite_ack), .B(n_408), .Z(n_961));
	notech_and4 i_1022(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[0]), .D(n_13618)
		, .Z(n_962));
	notech_and4 i_1024(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[1]), .D(n_13618)
		, .Z(n_963));
	notech_and4 i_1025(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[2]), .D(n_13618)
		, .Z(n_964));
	notech_and4 i_1026(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[3]), .D(n_13618)
		, .Z(n_965));
	notech_and4 i_1027(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[4]), .D(n_13618)
		, .Z(n_966));
	notech_and4 i_1028(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[5]), .D(n_13618)
		, .Z(n_967));
	notech_and4 i_1029(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[6]), .D(n_13618)
		, .Z(n_968));
	notech_and4 i_1030(.A(fsm[0]), .B(n_995), .C(fsm5_cnt_0[7]), .D(n_13618)
		, .Z(n_969));
	notech_and4 i_1031(.A(n_58636), .B(n_995), .C(fsm5_cnt_0[8]), .D(n_13618
		), .Z(n_970));
	notech_or4 i_1053(.A(n_972), .B(n_992), .C(n_1006), .D(n_1007), .Z(n_971
		));
	notech_nor2 i_4(.A(iwrite_req), .B(iread_req), .Z(n_972));
	notech_and3 i_1063(.A(n_13464), .B(n_995), .C(\tab11_0[4] ), .Z(n_973)
		);
	notech_and3 i_136(.A(n_995), .B(iwrite_req), .C(n_13464), .Z(n_974));
	notech_and3 i_1065(.A(n_995), .B(data_miss[1]), .C(n_13464), .Z(n_975)
		);
	notech_and4 i_1066(.A(n_13464), .B(data_miss[0]), .C(n_988), .D(\dir1_0[4] 
		), .Z(n_976));
	notech_nao3 i_94(.A(data_miss[0]), .B(n_13461), .C(n_989), .Z(n_977));
	notech_and2 i_1069(.A(iwrite_ack), .B(n_407), .Z(owrite_ack));
	notech_reg nx_dir_reg_0(.CP(n_61753), .D(n_10194), .CD(n_61056), .Q(nx_dir
		[0]));
	notech_mux2 i_15326(.S(n_977), .A(n_627), .B(nx_dir[0]), .Z(n_10194));
	notech_or2 i_75629(.A(n_654), .B(n_652), .Z(n_983));
	notech_reg nx_dir_reg_1(.CP(n_61753), .D(n_10204), .CD(n_61056), .Q(nx_dir
		[1]));
	notech_nand2 i_129(.A(n_13617), .B(n_13616), .Z(n_984));
	notech_ao3 i_15338(.A(nx_dir[1]), .B(1'b1), .C(n_13757), .Z(n_10204));
	notech_reg iDaddr_f_reg_0(.CP(n_61753), .D(n_10206), .CD(n_61056), .Q(iDaddr_f
		[0]));
	notech_mux2 i_15342(.S(n_948), .A(iDaddr[0]), .B(iDaddr_f[0]), .Z(n_10206
		));
	notech_or2 i_130(.A(n_58636), .B(fsm[3]), .Z(n_985));
	notech_reg iDaddr_f_reg_1(.CP(n_61753), .D(n_10212), .CD(n_61056), .Q(iDaddr_f
		[1]));
	notech_mux2 i_15350(.S(n_948), .A(iDaddr[1]), .B(iDaddr_f[1]), .Z(n_10212
		));
	notech_nao3 i_7(.A(n_983), .B(n_13464), .C(n_984), .Z(n_986));
	notech_reg iDaddr_f_reg_2(.CP(n_61753), .D(n_10218), .CD(n_61056), .Q(iDaddr_f
		[2]));
	notech_mux2 i_15358(.S(n_948), .A(iDaddr[2]), .B(iDaddr_f[2]), .Z(n_10218
		));
	notech_nand2 i_11(.A(iread_ack), .B(n_61605), .Z(n_987));
	notech_reg iDaddr_f_reg_3(.CP(n_61749), .D(n_10224), .CD(n_61052), .Q(iDaddr_f
		[3]));
	notech_mux2 i_15366(.S(n_948), .A(iDaddr[3]), .B(iDaddr_f[3]), .Z(n_10224
		));
	notech_and2 i_969(.A(fsm[1]), .B(n_13617), .Z(n_988));
	notech_reg iDaddr_f_reg_4(.CP(n_61749), .D(n_10230), .CD(n_61052), .Q(iDaddr_f
		[4]));
	notech_mux2 i_15374(.S(n_948), .A(iDaddr[4]), .B(iDaddr_f[4]), .Z(n_10230
		));
	notech_nao3 i_89(.A(n_988), .B(n_13618), .C(n_58636), .Z(n_989));
	notech_reg iDaddr_f_reg_5(.CP(n_61749), .D(n_10236), .CD(n_61052), .Q(iDaddr_f
		[5]));
	notech_mux2 i_15382(.S(n_948), .A(iDaddr[5]), .B(iDaddr_f[5]), .Z(n_10236
		));
	notech_nand3 i_10(.A(n_988), .B(data_miss[0]), .C(n_13464), .Z(n_990));
	notech_reg iDaddr_f_reg_6(.CP(n_61749), .D(n_10242), .CD(n_61052), .Q(iDaddr_f
		[6]));
	notech_mux2 i_15390(.S(n_948), .A(iDaddr[6]), .B(iDaddr_f[6]), .Z(n_10242
		));
	notech_reg iDaddr_f_reg_7(.CP(n_61754), .D(n_10248), .CD(n_61057), .Q(iDaddr_f
		[7]));
	notech_mux2 i_15398(.S(n_948), .A(iDaddr[7]), .B(iDaddr_f[7]), .Z(n_10248
		));
	notech_or4 i_72(.A(n_58636), .B(n_984), .C(fsm[3]), .D(n_13783), .Z(n_992
		));
	notech_reg iDaddr_f_reg_8(.CP(n_61753), .D(n_10254), .CD(n_61056), .Q(iDaddr_f
		[8]));
	notech_mux2 i_15406(.S(n_948), .A(iDaddr[8]), .B(iDaddr_f[8]), .Z(n_10254
		));
	notech_reg iDaddr_f_reg_9(.CP(n_61754), .D(n_10260), .CD(n_61057), .Q(iDaddr_f
		[9]));
	notech_mux2 i_15414(.S(n_948), .A(iDaddr[9]), .B(iDaddr_f[9]), .Z(n_10260
		));
	notech_ao4 i_20(.A(n_992), .B(n_13785), .C(n_627), .D(n_977), .Z(n_994)
		);
	notech_reg iDaddr_f_reg_10(.CP(n_61754), .D(n_10266), .CD(n_61057), .Q(iDaddr_f
		[10]));
	notech_mux2 i_15422(.S(n_948), .A(iDaddr[10]), .B(iDaddr_f[10]), .Z(n_10266
		));
	notech_and2 i_966(.A(fsm[2]), .B(n_13616), .Z(n_995));
	notech_reg iDaddr_f_reg_11(.CP(n_61753), .D(n_10272), .CD(n_61056), .Q(iDaddr_f
		[11]));
	notech_mux2 i_15430(.S(n_948), .A(iDaddr[11]), .B(iDaddr_f[11]), .Z(n_10272
		));
	notech_nao3 i_88(.A(n_995), .B(n_13618), .C(n_58636), .Z(n_996));
	notech_reg iDaddr_f_reg_12(.CP(n_61753), .D(\tab11_0[0] ), .CD(n_61056),
		 .Q(iDaddr_f[12]));
	notech_reg iDaddr_f_reg_13(.CP(n_61753), .D(\tab11_0[1] ), .CD(n_61056),
		 .Q(iDaddr_f[13]));
	notech_reg iDaddr_f_reg_14(.CP(n_61753), .D(\tab11_0[2] ), .CD(n_61056),
		 .Q(iDaddr_f[14]));
	notech_nand2 i_75673(.A(data_miss[0]), .B(n_605), .Z(n_999));
	notech_reg iDaddr_f_reg_15(.CP(n_61753), .D(\tab11_0[3] ), .CD(n_61056),
		 .Q(iDaddr_f[15]));
	notech_nand3 i_961(.A(n_995), .B(n_13464), .C(n_13462), .Z(n_1000));
	notech_reg iDaddr_f_reg_16(.CP(n_61748), .D(\tab11_0[4] ), .CD(n_61051),
		 .Q(iDaddr_f[16]));
	notech_nao3 i_17(.A(iread_ack), .B(n_61605), .C(n_1000), .Z(n_1001));
	notech_reg iDaddr_f_reg_17(.CP(n_61748), .D(\tab11_0[5] ), .CD(n_61051),
		 .Q(iDaddr_f[17]));
	notech_nand2 i_98(.A(hit_dir2), .B(n_13781), .Z(n_1002));
	notech_reg iDaddr_f_reg_18(.CP(n_61748), .D(\tab11_0[6] ), .CD(n_61051),
		 .Q(iDaddr_f[18]));
	notech_or4 i_12(.A(n_1000), .B(n_1002), .C(n_13784), .D(n_13783), .Z(n_1003
		));
	notech_reg iDaddr_f_reg_19(.CP(n_61748), .D(\tab11_0[7] ), .CD(n_61051),
		 .Q(iDaddr_f[19]));
	notech_reg iDaddr_f_reg_20(.CP(n_61748), .D(\tab11_0[8] ), .CD(n_61051),
		 .Q(iDaddr_f[20]));
	notech_or2 i_958(.A(busy_ram), .B(flush_tlb), .Z(n_1005));
	notech_reg iDaddr_f_reg_21(.CP(n_61748), .D(\tab11_0[9] ), .CD(n_61051),
		 .Q(iDaddr_f[21]));
	notech_or4 i_959(.A(pg_fault), .B(n_1005), .C(n_654), .D(n_652), .Z(n_1006
		));
	notech_reg iDaddr_f_reg_22(.CP(n_61748), .D(\dir1_0[0] ), .CD(n_61051), 
		.Q(iDaddr_f[22]));
	notech_nor2 i_6(.A(hit_dir2), .B(\hit_dir1[7] ), .Z(n_1007));
	notech_reg iDaddr_f_reg_23(.CP(n_61748), .D(\dir1_0[1] ), .CD(n_61051), 
		.Q(iDaddr_f[23]));
	notech_reg iDaddr_f_reg_24(.CP(n_61748), .D(\dir1_0[2] ), .CD(n_61051), 
		.Q(iDaddr_f[24]));
	notech_reg iDaddr_f_reg_25(.CP(n_61749), .D(\dir1_0[3] ), .CD(n_61052), 
		.Q(iDaddr_f[25]));
	notech_or2 i_97(.A(hit_dir2), .B(n_13781), .Z(n_1010));
	notech_reg iDaddr_f_reg_26(.CP(n_61749), .D(\dir1_0[4] ), .CD(n_61052), 
		.Q(iDaddr_f[26]));
	notech_or4 i_13(.A(n_1000), .B(n_1010), .C(n_13784), .D(n_13783), .Z(n_1011
		));
	notech_reg iDaddr_f_reg_27(.CP(n_61749), .D(\dir1_0[5] ), .CD(n_61052), 
		.Q(iDaddr_f[27]));
	notech_reg iDaddr_f_reg_28(.CP(n_61749), .D(\dir1_0[6] ), .CD(n_61052), 
		.Q(iDaddr_f[28]));
	notech_reg iDaddr_f_reg_29(.CP(n_61749), .D(\dir1_0[7] ), .CD(n_61052), 
		.Q(iDaddr_f[29]));
	notech_reg iDaddr_f_reg_30(.CP(n_61748), .D(\dir1_0[8] ), .CD(n_61051), 
		.Q(iDaddr_f[30]));
	notech_nand2 i_78(.A(n_58636), .B(n_13618), .Z(n_1015));
	notech_reg iDaddr_f_reg_31(.CP(n_61748), .D(\dir1_0[9] ), .CD(n_61051), 
		.Q(iDaddr_f[31]));
	notech_nand3 i_75725(.A(fsm[0]), .B(n_988), .C(n_13618), .Z(n_1016));
	notech_reg_set dir1_reg_0(.CP(n_61749), .D(n_10398), .SD(n_61052), .Q(\dir1[0] 
		));
	notech_mux2 i_15598(.S(\nbus_14042[0] ), .A(\dir1[0] ), .B(n_55516), .Z(n_10398
		));
	notech_or2 i_71(.A(hit_adr11), .B(n_1016), .Z(n_1017));
	notech_reg_set dir1_reg_1(.CP(n_61749), .D(n_10404), .SD(n_61052), .Q(\dir1[1] 
		));
	notech_mux2 i_15606(.S(\nbus_14042[0] ), .A(\dir1[1] ), .B(n_55522), .Z(n_10404
		));
	notech_nor2 i_16(.A(hit_adr13), .B(hit_adr14), .Z(n_1018));
	notech_reg_set dir1_reg_2(.CP(n_61754), .D(n_10410), .SD(n_61057), .Q(\dir1[2] 
		));
	notech_mux2 i_15614(.S(\nbus_14042[0] ), .A(\dir1[2] ), .B(n_55528), .Z(n_10410
		));
	notech_nand2 i_131(.A(n_1018), .B(n_13512), .Z(n_1019));
	notech_reg_set dir1_reg_3(.CP(n_61757), .D(n_10416), .SD(n_61060), .Q(\dir1[3] 
		));
	notech_mux2 i_15622(.S(\nbus_14042[0] ), .A(\dir1[3] ), .B(n_55534), .Z(n_10416
		));
	notech_nao3 i_9(.A(n_988), .B(n_61605), .C(n_1015), .Z(n_1020));
	notech_reg dir1_reg_4(.CP(n_61757), .D(n_10422), .CD(n_61060), .Q(\dir1[4] 
		));
	notech_mux2 i_15630(.S(\nbus_14042[0] ), .A(\dir1[4] ), .B(n_976), .Z(n_10422
		));
	notech_reg_set dir1_reg_5(.CP(n_61757), .D(n_10428), .SD(n_61060), .Q(\dir1[5] 
		));
	notech_mux2 i_15638(.S(\nbus_14042[0] ), .A(\dir1[5] ), .B(n_55546), .Z(n_10428
		));
	notech_reg_set dir1_reg_6(.CP(n_61757), .D(n_10434), .SD(n_61060), .Q(\dir1[6] 
		));
	notech_mux2 i_15646(.S(\nbus_14042[0] ), .A(\dir1[6] ), .B(n_55552), .Z(n_10434
		));
	notech_reg_set dir1_reg_7(.CP(n_61757), .D(n_10440), .SD(n_61060), .Q(\dir1[7] 
		));
	notech_mux2 i_15654(.S(\nbus_14042[0] ), .A(\dir1[7] ), .B(n_55558), .Z(n_10440
		));
	notech_nor2 i_31(.A(hit_adr23), .B(hit_adr24), .Z(n_1024));
	notech_reg_set dir1_reg_8(.CP(n_61757), .D(n_10446), .SD(n_61060), .Q(\dir1[8] 
		));
	notech_mux2 i_15662(.S(\nbus_14042[0] ), .A(\dir1[8] ), .B(n_55564), .Z(n_10446
		));
	notech_nand2 i_132(.A(n_1024), .B(n_13564), .Z(n_1025));
	notech_reg_set dir1_reg_9(.CP(n_61757), .D(n_10452), .SD(n_61060), .Q(\dir1[9] 
		));
	notech_mux2 i_15670(.S(\nbus_14042[0] ), .A(\dir1[9] ), .B(n_55570), .Z(n_10452
		));
	notech_or2 i_73(.A(hit_adr21), .B(n_1016), .Z(n_1026));
	notech_reg_set dir1_reg_10(.CP(n_61757), .D(n_10458), .SD(n_61060), .Q(\dir1[10] 
		));
	notech_mux2 i_15678(.S(\nbus_14042[0] ), .A(\dir1[10] ), .B(n_55576), .Z
		(n_10458));
	notech_reg_set dir1_reg_11(.CP(n_61757), .D(n_10464), .SD(n_61060), .Q(\dir1[11] 
		));
	notech_mux2 i_15686(.S(\nbus_14042[0] ), .A(\dir1[11] ), .B(n_55582), .Z
		(n_10464));
	notech_nand3 i_75732(.A(n_58636), .B(n_995), .C(n_13618), .Z(n_1028));
	notech_reg_set dir1_reg_12(.CP(n_61758), .D(n_10470), .SD(n_61061), .Q(\dir1[12] 
		));
	notech_mux2 i_15694(.S(\nbus_14042[0] ), .A(\dir1[12] ), .B(n_55588), .Z
		(n_10470));
	notech_reg_set dir1_reg_13(.CP(n_61758), .D(n_10476), .SD(n_61061), .Q(\dir1[13] 
		));
	notech_mux2 i_15702(.S(\nbus_14042[0] ), .A(\dir1[13] ), .B(n_55594), .Z
		(n_10476));
	notech_or2 i_50(.A(n_553), .B(fsm5_cnt[8]), .Z(n_1030));
	notech_reg_set dir1_reg_14(.CP(n_61758), .D(n_10482), .SD(n_61061), .Q(\dir1[14] 
		));
	notech_mux2 i_15710(.S(\nbus_14042[0] ), .A(\dir1[14] ), .B(n_55600), .Z
		(n_10482));
	notech_reg_set dir1_reg_15(.CP(n_61758), .D(n_10488), .SD(n_61061), .Q(\dir1[15] 
		));
	notech_mux2 i_15718(.S(\nbus_14042[0] ), .A(\dir1[15] ), .B(n_55606), .Z
		(n_10488));
	notech_nand2 i_69(.A(fsm[2]), .B(fsm[1]), .Z(n_1032));
	notech_reg_set dir1_reg_16(.CP(n_61758), .D(n_10494), .SD(n_61061), .Q(\dir1[16] 
		));
	notech_mux2 i_15726(.S(n_54570), .A(\dir1[16] ), .B(n_55612), .Z(n_10494
		));
	notech_ao4 i_932(.A(n_990), .B(data_miss[5]), .C(iwrite_ack), .D(n_1032)
		, .Z(n_1033));
	notech_reg_set dir1_reg_17(.CP(n_61757), .D(n_10500), .SD(n_61060), .Q(\dir1[17] 
		));
	notech_mux2 i_15734(.S(n_54570), .A(\dir1[17] ), .B(n_55618), .Z(n_10500
		));
	notech_reg_set dir1_reg_18(.CP(n_61757), .D(n_10506), .SD(n_61060), .Q(\dir1[18] 
		));
	notech_mux2 i_15742(.S(n_54570), .A(\dir1[18] ), .B(n_55624), .Z(n_10506
		));
	notech_or2 i_95(.A(n_549), .B(n_13614), .Z(n_1035));
	notech_reg_set dir1_reg_19(.CP(n_61758), .D(n_10512), .SD(n_61061), .Q(\dir1[19] 
		));
	notech_mux2 i_15750(.S(n_54570), .A(\dir1[19] ), .B(n_55630), .Z(n_10512
		));
	notech_reg_set dir1_reg_20(.CP(n_61758), .D(n_10518), .SD(n_61061), .Q(\dir1[20] 
		));
	notech_mux2 i_15758(.S(n_54570), .A(\dir1[20] ), .B(n_55636), .Z(n_10518
		));
	notech_reg_set dir1_reg_21(.CP(n_61754), .D(n_10524), .SD(n_61057), .Q(\dir1[21] 
		));
	notech_mux2 i_15766(.S(n_54570), .A(\dir1[21] ), .B(n_55642), .Z(n_10524
		));
	notech_ao4 i_927(.A(n_546), .B(iwrite_ack), .C(n_550), .D(n_1000), .Z(n_1038
		));
	notech_reg_set dir1_reg_22(.CP(n_61754), .D(n_10530), .SD(n_61057), .Q(\dir1[22] 
		));
	notech_mux2 i_15774(.S(n_54570), .A(\dir1[22] ), .B(n_55648), .Z(n_10530
		));
	notech_reg_set dir1_reg_23(.CP(n_61755), .D(n_10536), .SD(n_61058), .Q(\dir1[23] 
		));
	notech_mux2 i_15782(.S(n_54570), .A(\dir1[23] ), .B(n_55654), .Z(n_10536
		));
	notech_nao3 i_75718(.A(n_58636), .B(n_13618), .C(n_984), .Z(n_1040));
	notech_reg_set dir1_reg_24(.CP(n_61755), .D(n_10542), .SD(n_61058), .Q(\dir1[24] 
		));
	notech_mux2 i_15790(.S(n_54570), .A(\dir1[24] ), .B(n_55660), .Z(n_10542
		));
	notech_reg_set dir1_reg_25(.CP(n_61754), .D(n_10548), .SD(n_61057), .Q(\dir1[25] 
		));
	notech_mux2 i_15798(.S(n_54570), .A(\dir1[25] ), .B(n_55666), .Z(n_10548
		));
	notech_nand3 i_81(.A(fsm[2]), .B(fsm[1]), .C(n_13618), .Z(n_1042));
	notech_reg_set dir1_reg_26(.CP(n_61754), .D(n_10554), .SD(n_61057), .Q(\dir1[26] 
		));
	notech_mux2 i_15806(.S(n_54570), .A(\dir1[26] ), .B(n_55672), .Z(n_10554
		));
	notech_or4 i_14(.A(n_13617), .B(n_13616), .C(fsm[3]), .D(n_13783), .Z(n_1043
		));
	notech_reg_set dir1_reg_27(.CP(n_61754), .D(n_10560), .SD(n_61057), .Q(\dir1[27] 
		));
	notech_mux2 i_15814(.S(n_54570), .A(\dir1[27] ), .B(n_55678), .Z(n_10560
		));
	notech_reg_set dir1_reg_28(.CP(n_61754), .D(n_10566), .SD(n_61057), .Q(\dir1[28] 
		));
	notech_mux2 i_15822(.S(n_54570), .A(\dir1[28] ), .B(n_55684), .Z(n_10566
		));
	notech_reg_set dir1_reg_29(.CP(n_61754), .D(n_10572), .SD(n_61057), .Q(\dir1[29] 
		));
	notech_mux2 i_15830(.S(n_54570), .A(\dir1[29] ), .B(n_55690), .Z(n_10572
		));
	notech_reg_set dir1_reg_33(.CP(n_61755), .D(n_10578), .SD(n_61058), .Q(\dir1[33] 
		));
	notech_mux2 i_15838(.S(n_54570), .A(\dir1[33] ), .B(n_13488), .Z(n_10578
		));
	notech_reg_set dir2_reg_0(.CP(n_61755), .D(n_10584), .SD(n_61058), .Q(\dir2[0] 
		));
	notech_mux2 i_15846(.S(\nbus_14043[0] ), .A(\dir2[0] ), .B(n_55516), .Z(n_10584
		));
	notech_nand3 i_921(.A(n_952), .B(n_1043), .C(n_953), .Z(n_1048));
	notech_reg_set dir2_reg_1(.CP(n_61755), .D(n_10590), .SD(n_61058), .Q(\dir2[1] 
		));
	notech_mux2 i_15854(.S(\nbus_14043[0] ), .A(\dir2[1] ), .B(n_55522), .Z(n_10590
		));
	notech_reg_set dir2_reg_2(.CP(n_61755), .D(n_10596), .SD(n_61058), .Q(\dir2[2] 
		));
	notech_mux2 i_15862(.S(\nbus_14043[0] ), .A(\dir2[2] ), .B(n_55528), .Z(n_10596
		));
	notech_ao4 i_917(.A(n_1032), .B(n_1015), .C(n_541), .D(n_13618), .Z(n_1050
		));
	notech_reg_set dir2_reg_3(.CP(n_61755), .D(n_10602), .SD(n_61058), .Q(\dir2[3] 
		));
	notech_mux2 i_15870(.S(\nbus_14043[0] ), .A(\dir2[3] ), .B(n_55534), .Z(n_10602
		));
	notech_reg dir2_reg_4(.CP(n_61755), .D(n_10608), .CD(n_61058), .Q(\dir2[4] 
		));
	notech_mux2 i_15878(.S(\nbus_14043[0] ), .A(\dir2[4] ), .B(n_976), .Z(n_10608
		));
	notech_reg_set dir2_reg_5(.CP(n_61755), .D(n_10614), .SD(n_61058), .Q(\dir2[5] 
		));
	notech_mux2 i_15886(.S(\nbus_14043[0] ), .A(\dir2[5] ), .B(n_55546), .Z(n_10614
		));
	notech_nand2 i_44(.A(n_61599), .B(n_53478), .Z(n_1053));
	notech_reg_set dir2_reg_6(.CP(n_61755), .D(n_10620), .SD(n_61058), .Q(\dir2[6] 
		));
	notech_mux2 i_15894(.S(\nbus_14043[0] ), .A(\dir2[6] ), .B(n_55552), .Z(n_10620
		));
	notech_reg_set dir2_reg_7(.CP(n_61755), .D(n_10626), .SD(n_61058), .Q(\dir2[7] 
		));
	notech_mux2 i_15902(.S(\nbus_14043[0] ), .A(\dir2[7] ), .B(n_55558), .Z(n_10626
		));
	notech_reg_set dir2_reg_8(.CP(n_61747), .D(n_10632), .SD(n_61050), .Q(\dir2[8] 
		));
	notech_mux2 i_15910(.S(\nbus_14043[0] ), .A(\dir2[8] ), .B(n_55564), .Z(n_10632
		));
	notech_nao3 i_29(.A(n_988), .B(n_58609), .C(n_1015), .Z(n_1056));
	notech_reg_set dir2_reg_9(.CP(n_61740), .D(n_10638), .SD(n_61043), .Q(\dir2[9] 
		));
	notech_mux2 i_15918(.S(\nbus_14043[0] ), .A(\dir2[9] ), .B(n_55570), .Z(n_10638
		));
	notech_ao4 i_914(.A(n_1056), .B(n_13487), .C(n_1040), .D(n_13703), .Z(n_1057
		));
	notech_reg_set dir2_reg_10(.CP(n_61740), .D(n_10644), .SD(n_61043), .Q(\dir2[10] 
		));
	notech_mux2 i_15926(.S(\nbus_14043[0] ), .A(\dir2[10] ), .B(n_55576), .Z
		(n_10644));
	notech_ao4 i_913(.A(n_1056), .B(n_13486), .C(n_1040), .D(n_13704), .Z(n_1058
		));
	notech_reg_set dir2_reg_11(.CP(n_61740), .D(n_10650), .SD(n_61043), .Q(\dir2[11] 
		));
	notech_mux2 i_15934(.S(\nbus_14043[0] ), .A(\dir2[11] ), .B(n_55582), .Z
		(n_10650));
	notech_ao4 i_912(.A(n_1056), .B(n_13485), .C(n_1040), .D(n_13705), .Z(n_1059
		));
	notech_reg_set dir2_reg_12(.CP(n_61740), .D(n_10656), .SD(n_61043), .Q(\dir2[12] 
		));
	notech_mux2 i_15942(.S(\nbus_14043[0] ), .A(\dir2[12] ), .B(n_55588), .Z
		(n_10656));
	notech_ao4 i_911(.A(n_1056), .B(n_13483), .C(n_1040), .D(n_13706), .Z(n_1060
		));
	notech_reg_set dir2_reg_13(.CP(n_61740), .D(n_10662), .SD(n_61043), .Q(\dir2[13] 
		));
	notech_mux2 i_15950(.S(\nbus_14043[0] ), .A(\dir2[13] ), .B(n_55594), .Z
		(n_10662));
	notech_ao4 i_910(.A(n_1056), .B(n_13482), .C(n_1040), .D(n_13707), .Z(n_1061
		));
	notech_reg_set dir2_reg_14(.CP(n_61740), .D(n_10668), .SD(n_61043), .Q(\dir2[14] 
		));
	notech_mux2 i_15958(.S(\nbus_14043[0] ), .A(\dir2[14] ), .B(n_55600), .Z
		(n_10668));
	notech_ao4 i_909(.A(n_1056), .B(n_13481), .C(n_1040), .D(n_13708), .Z(n_1062
		));
	notech_reg_set dir2_reg_15(.CP(n_61739), .D(n_10674), .SD(n_61042), .Q(\dir2[15] 
		));
	notech_mux2 i_15966(.S(\nbus_14043[0] ), .A(\dir2[15] ), .B(n_55606), .Z
		(n_10674));
	notech_ao4 i_908(.A(n_1056), .B(n_13480), .C(n_1040), .D(n_13709), .Z(n_1063
		));
	notech_reg_set dir2_reg_16(.CP(n_61740), .D(n_10680), .SD(n_61043), .Q(\dir2[16] 
		));
	notech_mux2 i_15974(.S(n_54648), .A(\dir2[16] ), .B(n_55612), .Z(n_10680
		));
	notech_ao4 i_907(.A(n_1056), .B(n_13479), .C(n_1040), .D(n_13710), .Z(n_1064
		));
	notech_reg_set dir2_reg_17(.CP(n_61740), .D(n_10686), .SD(n_61043), .Q(\dir2[17] 
		));
	notech_mux2 i_15982(.S(n_54648), .A(\dir2[17] ), .B(n_55618), .Z(n_10686
		));
	notech_ao4 i_906(.A(n_1056), .B(n_13478), .C(n_1040), .D(n_13711), .Z(n_1065
		));
	notech_reg_set dir2_reg_18(.CP(n_61743), .D(n_10692), .SD(n_61046), .Q(\dir2[18] 
		));
	notech_mux2 i_15990(.S(n_54648), .A(\dir2[18] ), .B(n_55624), .Z(n_10692
		));
	notech_ao4 i_905(.A(n_1056), .B(n_13477), .C(n_1040), .D(n_13712), .Z(n_1066
		));
	notech_reg_set dir2_reg_19(.CP(n_61743), .D(n_10698), .SD(n_61046), .Q(\dir2[19] 
		));
	notech_mux2 i_15998(.S(n_54648), .A(\dir2[19] ), .B(n_55630), .Z(n_10698
		));
	notech_ao4 i_904(.A(n_1056), .B(n_13476), .C(n_1040), .D(n_13713), .Z(n_1067
		));
	notech_reg_set dir2_reg_20(.CP(n_61743), .D(n_10704), .SD(n_61046), .Q(\dir2[20] 
		));
	notech_mux2 i_16006(.S(n_54648), .A(\dir2[20] ), .B(n_55636), .Z(n_10704
		));
	notech_ao4 i_903(.A(n_1056), .B(n_13475), .C(n_1040), .D(n_13714), .Z(n_1068
		));
	notech_reg_set dir2_reg_21(.CP(n_61743), .D(n_10710), .SD(n_61046), .Q(\dir2[21] 
		));
	notech_mux2 i_16014(.S(n_54648), .A(\dir2[21] ), .B(n_55642), .Z(n_10710
		));
	notech_ao4 i_902(.A(n_1056), .B(n_13474), .C(n_1040), .D(n_13715), .Z(n_1069
		));
	notech_reg_set dir2_reg_22(.CP(n_61743), .D(n_10716), .SD(n_61046), .Q(\dir2[22] 
		));
	notech_mux2 i_16022(.S(n_54648), .A(\dir2[22] ), .B(n_55648), .Z(n_10716
		));
	notech_ao4 i_901(.A(n_1056), .B(n_13473), .C(n_1040), .D(n_13716), .Z(n_1070
		));
	notech_reg_set dir2_reg_23(.CP(n_61740), .D(n_10722), .SD(n_61043), .Q(\dir2[23] 
		));
	notech_mux2 i_16030(.S(n_54648), .A(\dir2[23] ), .B(n_55654), .Z(n_10722
		));
	notech_ao4 i_900(.A(n_1056), .B(n_13472), .C(n_1040), .D(n_13717), .Z(n_1071
		));
	notech_reg_set dir2_reg_24(.CP(n_61740), .D(n_10728), .SD(n_61043), .Q(\dir2[24] 
		));
	notech_mux2 i_16038(.S(n_54648), .A(\dir2[24] ), .B(n_55660), .Z(n_10728
		));
	notech_ao4 i_899(.A(n_1056), .B(n_13471), .C(n_1040), .D(n_13718), .Z(n_1072
		));
	notech_reg_set dir2_reg_25(.CP(n_61743), .D(n_10734), .SD(n_61046), .Q(\dir2[25] 
		));
	notech_mux2 i_16046(.S(n_54648), .A(\dir2[25] ), .B(n_55666), .Z(n_10734
		));
	notech_ao4 i_898(.A(n_1056), .B(n_13470), .C(n_54796), .D(n_13719), .Z(n_1073
		));
	notech_reg_set dir2_reg_26(.CP(n_61740), .D(n_10740), .SD(n_61043), .Q(\dir2[26] 
		));
	notech_mux2 i_16054(.S(n_54648), .A(\dir2[26] ), .B(n_55672), .Z(n_10740
		));
	notech_ao4 i_897(.A(n_1056), .B(n_13469), .C(n_54796), .D(n_13720), .Z(n_1074
		));
	notech_reg_set dir2_reg_27(.CP(n_61738), .D(n_10746), .SD(n_61041), .Q(\dir2[27] 
		));
	notech_mux2 i_16062(.S(n_54648), .A(\dir2[27] ), .B(n_55678), .Z(n_10746
		));
	notech_ao4 i_896(.A(n_1056), .B(n_13468), .C(n_54796), .D(n_13721), .Z(n_1075
		));
	notech_reg_set dir2_reg_28(.CP(n_61738), .D(n_10752), .SD(n_61041), .Q(\dir2[28] 
		));
	notech_mux2 i_16070(.S(n_54648), .A(\dir2[28] ), .B(n_55684), .Z(n_10752
		));
	notech_ao4 i_895(.A(n_1056), .B(n_13467), .C(n_54796), .D(n_13722), .Z(n_1076
		));
	notech_reg_set dir2_reg_29(.CP(n_61739), .D(n_10758), .SD(n_61042), .Q(\dir2[29] 
		));
	notech_mux2 i_16078(.S(n_54648), .A(\dir2[29] ), .B(n_55690), .Z(n_10758
		));
	notech_nand2 i_83(.A(n_406), .B(n_13629), .Z(n_1077));
	notech_reg_set dir2_reg_33(.CP(n_61738), .D(n_10764), .SD(n_61041), .Q(\dir2[33] 
		));
	notech_mux2 i_16086(.S(n_54648), .A(\dir2[33] ), .B(n_13488), .Z(n_10764
		));
	notech_reg_set tab21_reg_0(.CP(n_61738), .D(n_10770), .SD(n_61041), .Q(\tab21[0] 
		));
	notech_mux2 i_16094(.S(\nbus_14036[0] ), .A(\tab21[0] ), .B(n_52377), .Z
		(n_10770));
	notech_reg_set tab21_reg_1(.CP(n_61738), .D(n_10776), .SD(n_61041), .Q(\tab21[1] 
		));
	notech_mux2 i_16102(.S(\nbus_14036[0] ), .A(\tab21[1] ), .B(n_52383), .Z
		(n_10776));
	notech_nand3 i_1(.A(n_61599), .B(n_53478), .C(n_983), .Z(n_1080));
	notech_reg_set tab21_reg_2(.CP(n_61738), .D(n_10782), .SD(n_61041), .Q(\tab21[2] 
		));
	notech_mux2 i_16110(.S(\nbus_14036[0] ), .A(\tab21[2] ), .B(n_52389), .Z
		(n_10782));
	notech_or4 i_77(.A(n_58609), .B(n_13783), .C(n_13463), .D(n_13465), .Z(n_1081
		));
	notech_reg_set tab21_reg_3(.CP(n_61738), .D(n_10788), .SD(n_61041), .Q(\tab21[3] 
		));
	notech_mux2 i_16118(.S(\nbus_14036[0] ), .A(\tab21[3] ), .B(n_52395), .Z
		(n_10788));
	notech_reg tab21_reg_4(.CP(n_61738), .D(n_10794), .CD(n_61041), .Q(\tab21[4] 
		));
	notech_mux2 i_16126(.S(\nbus_14036[0] ), .A(\tab21[4] ), .B(n_973), .Z(n_10794
		));
	notech_reg_set tab21_reg_5(.CP(n_61739), .D(n_10800), .SD(n_61042), .Q(\tab21[5] 
		));
	notech_mux2 i_16134(.S(\nbus_14036[0] ), .A(\tab21[5] ), .B(n_52407), .Z
		(n_10800));
	notech_nao3 i_27(.A(hit_tab22), .B(n_13782), .C(n_53446), .Z(n_1084));
	notech_reg_set tab21_reg_6(.CP(n_61739), .D(n_10806), .SD(n_61042), .Q(\tab21[6] 
		));
	notech_mux2 i_16142(.S(\nbus_14036[0] ), .A(\tab21[6] ), .B(n_52413), .Z
		(n_10806));
	notech_nao3 i_75(.A(n_58609), .B(n_983), .C(n_1053), .Z(n_1085));
	notech_reg_set tab21_reg_7(.CP(n_61739), .D(n_10812), .SD(n_61042), .Q(\tab21[7] 
		));
	notech_mux2 i_16150(.S(\nbus_14036[0] ), .A(\tab21[7] ), .B(n_52419), .Z
		(n_10812));
	notech_or4 i_30(.A(hit_tab12), .B(n_58600), .C(hit_tab13), .D(n_1085), .Z
		(n_1086));
	notech_reg_set tab21_reg_8(.CP(n_61739), .D(n_10818), .SD(n_61042), .Q(\tab21[8] 
		));
	notech_mux2 i_16158(.S(\nbus_14036[0] ), .A(\tab21[8] ), .B(n_52425), .Z
		(n_10818));
	notech_ao4 i_884(.A(n_1086), .B(n_13534), .C(n_1084), .D(n_13563), .Z(n_1087
		));
	notech_reg_set tab21_reg_9(.CP(n_61739), .D(n_10824), .SD(n_61042), .Q(\tab21[9] 
		));
	notech_mux2 i_16166(.S(\nbus_14036[0] ), .A(\tab21[9] ), .B(n_52431), .Z
		(n_10824));
	notech_reg_set tab21_reg_10(.CP(n_61739), .D(n_10830), .SD(n_61042), .Q(\tab21[10] 
		));
	notech_mux2 i_16174(.S(\nbus_14036[0] ), .A(\tab21[10] ), .B(n_52437), .Z
		(n_10830));
	notech_reg_set tab21_reg_11(.CP(n_61739), .D(n_10836), .SD(n_61042), .Q(\tab21[11] 
		));
	notech_mux2 i_16182(.S(\nbus_14036[0] ), .A(\tab21[11] ), .B(n_52443), .Z
		(n_10836));
	notech_or4 i_24(.A(hit_tab22), .B(n_58618), .C(n_53446), .D(hit_tab23), 
		.Z(n_1090));
	notech_reg_set tab21_reg_12(.CP(n_61739), .D(n_10842), .SD(n_61042), .Q(\tab21[12] 
		));
	notech_mux2 i_16190(.S(\nbus_14036[0] ), .A(\tab21[12] ), .B(n_52449), .Z
		(n_10842));
	notech_reg_set tab21_reg_13(.CP(n_61739), .D(n_10848), .SD(n_61042), .Q(\tab21[13] 
		));
	notech_mux2 i_16198(.S(\nbus_14036[0] ), .A(\tab21[13] ), .B(n_52455), .Z
		(n_10848));
	notech_or4 i_26(.A(hit_tab22), .B(n_58618), .C(n_53446), .D(n_13780), .Z
		(n_1092));
	notech_reg_set tab21_reg_14(.CP(n_61743), .D(n_10854), .SD(n_61046), .Q(\tab21[14] 
		));
	notech_mux2 i_16206(.S(\nbus_14036[0] ), .A(\tab21[14] ), .B(n_52461), .Z
		(n_10854));
	notech_ao4 i_882(.A(n_1092), .B(n_13584), .C(n_1090), .D(n_13604), .Z(n_1093
		));
	notech_reg_set tab21_reg_15(.CP(n_61745), .D(n_10860), .SD(n_61048), .Q(\tab21[15] 
		));
	notech_mux2 i_16214(.S(\nbus_14036[0] ), .A(\tab21[15] ), .B(n_52467), .Z
		(n_10860));
	notech_reg_set tab21_reg_16(.CP(n_61745), .D(n_10866), .SD(n_61048), .Q(\tab21[16] 
		));
	notech_mux2 i_16222(.S(\nbus_14036[0] ), .A(\tab21[16] ), .B(n_52473), .Z
		(n_10866));
	notech_and4 i_886(.A(n_1093), .B(n_1087), .C(n_898), .D(n_901), .Z(n_1095
		));
	notech_reg_set tab21_reg_17(.CP(n_61747), .D(n_10872), .SD(n_61050), .Q(\tab21[17] 
		));
	notech_mux2 i_16230(.S(n_54590), .A(\tab21[17] ), .B(n_52479), .Z(n_10872
		));
	notech_ao3 i_887(.A(hit_tab13), .B(n_13779), .C(n_58600), .Z(n_1096));
	notech_reg_set tab21_reg_18(.CP(n_61745), .D(n_10878), .SD(n_61048), .Q(\tab21[18] 
		));
	notech_mux2 i_16238(.S(n_54590), .A(\tab21[18] ), .B(n_52485), .Z(n_10878
		));
	notech_reg_set tab21_reg_19(.CP(n_61745), .D(n_10884), .SD(n_61048), .Q(\tab21[19] 
		));
	notech_mux2 i_16246(.S(n_54590), .A(\tab21[19] ), .B(n_52491), .Z(n_10884
		));
	notech_or4 i_15(.A(n_654), .B(n_652), .C(n_13783), .D(n_13463), .Z(n_1098
		));
	notech_reg_set tab21_reg_20(.CP(n_61745), .D(n_10890), .SD(n_61048), .Q(\tab21[20] 
		));
	notech_mux2 i_16254(.S(n_54590), .A(\tab21[20] ), .B(n_52497), .Z(n_10890
		));
	notech_reg_set tab21_reg_21(.CP(n_61745), .D(n_10896), .SD(n_61048), .Q(\tab21[21] 
		));
	notech_mux2 i_16262(.S(n_54590), .A(\tab21[21] ), .B(n_52503), .Z(n_10896
		));
	notech_nao3 i_23(.A(hit_tab12), .B(n_53468), .C(n_58600), .Z(n_1100));
	notech_reg_set tab21_reg_22(.CP(n_61745), .D(n_10902), .SD(n_61048), .Q(\tab21[22] 
		));
	notech_mux2 i_16270(.S(n_54590), .A(\tab21[22] ), .B(n_52509), .Z(n_10902
		));
	notech_ao4 i_879(.A(n_1100), .B(n_13511), .C(n_1098), .D(n_13680), .Z(n_1101
		));
	notech_reg_set tab21_reg_23(.CP(n_61745), .D(n_10908), .SD(n_61048), .Q(\tab21[23] 
		));
	notech_mux2 i_16278(.S(n_54590), .A(\tab21[23] ), .B(n_52515), .Z(n_10908
		));
	notech_reg_set tab21_reg_24(.CP(n_61747), .D(n_10914), .SD(n_61050), .Q(\tab21[24] 
		));
	notech_mux2 i_16286(.S(n_54590), .A(\tab21[24] ), .B(n_52521), .Z(n_10914
		));
	notech_ao4 i_878(.A(n_61599), .B(n_13754), .C(n_1043), .D(n_13681), .Z(n_1103
		));
	notech_reg_set tab21_reg_25(.CP(n_61747), .D(n_10920), .SD(n_61050), .Q(\tab21[25] 
		));
	notech_mux2 i_16294(.S(n_54590), .A(\tab21[25] ), .B(n_52527), .Z(n_10920
		));
	notech_reg_set tab21_reg_26(.CP(n_61747), .D(n_10926), .SD(n_61050), .Q(\tab21[26] 
		));
	notech_mux2 i_16302(.S(n_54590), .A(\tab21[26] ), .B(n_52533), .Z(n_10926
		));
	notech_ao4 i_875(.A(n_1086), .B(n_13533), .C(n_1084), .D(n_13562), .Z(n_1105
		));
	notech_reg_set tab21_reg_27(.CP(n_61747), .D(n_10932), .SD(n_61050), .Q(\tab21[27] 
		));
	notech_mux2 i_16310(.S(\nbus_14036[0] ), .A(\tab21[27] ), .B(n_52539), .Z
		(n_10932));
	notech_reg_set tab21_reg_28(.CP(n_61747), .D(n_10938), .SD(n_61050), .Q(\tab21[28] 
		));
	notech_mux2 i_16318(.S(n_54590), .A(\tab21[28] ), .B(n_52545), .Z(n_10938
		));
	notech_ao4 i_873(.A(n_1092), .B(n_13583), .C(n_1090), .D(n_13603), .Z(n_1107
		));
	notech_reg_set tab21_reg_29(.CP(n_61747), .D(n_10944), .SD(n_61050), .Q(\tab21[29] 
		));
	notech_mux2 i_16326(.S(n_54590), .A(\tab21[29] ), .B(n_52551), .Z(n_10944
		));
	notech_reg tab21_reg_30(.CP(n_61747), .D(n_10950), .CD(n_61050), .Q(\tab21[30] 
		));
	notech_mux2 i_16334(.S(n_54590), .A(\tab21[30] ), .B(n_974), .Z(n_10950)
		);
	notech_and4 i_877(.A(n_1107), .B(n_1105), .C(n_887), .D(n_890), .Z(n_1109
		));
	notech_reg tab21_reg_32(.CP(n_61747), .D(n_10956), .CD(n_61050), .Q(\tab21[32] 
		));
	notech_mux2 i_16342(.S(n_54590), .A(\tab21[32] ), .B(n_975), .Z(n_10956)
		);
	notech_ao4 i_870(.A(n_1100), .B(n_13510), .C(n_1098), .D(n_13678), .Z(n_1110
		));
	notech_reg_set tab21_reg_33(.CP(n_61747), .D(n_10962), .SD(n_61050), .Q(\tab21[33] 
		));
	notech_mux2 i_16350(.S(n_54590), .A(\tab21[33] ), .B(n_54613), .Z(n_10962
		));
	notech_reg hit_adr11_reg(.CP(n_61744), .D(n_10968), .CD(n_61047), .Q(hit_adr11
		));
	notech_mux2 i_16358(.S(n_971), .A(hit_add11), .B(hit_adr11), .Z(n_10968)
		);
	notech_ao4 i_869(.A(n_61599), .B(n_13753), .C(n_1043), .D(n_13679), .Z(n_1112
		));
	notech_reg_set tab12_reg_0(.CP(n_61744), .D(n_10974), .SD(n_61047), .Q(\tab12[0] 
		));
	notech_mux2 i_16366(.S(\nbus_14035[0] ), .A(\tab12[0] ), .B(n_52377), .Z
		(n_10974));
	notech_reg_set tab12_reg_1(.CP(n_61744), .D(n_10980), .SD(n_61047), .Q(\tab12[1] 
		));
	notech_mux2 i_16374(.S(\nbus_14035[0] ), .A(\tab12[1] ), .B(n_52383), .Z
		(n_10980));
	notech_ao4 i_866(.A(n_1086), .B(n_13532), .C(n_1084), .D(n_13561), .Z(n_1114
		));
	notech_reg_set tab12_reg_2(.CP(n_61744), .D(n_10986), .SD(n_61047), .Q(\tab12[2] 
		));
	notech_mux2 i_16382(.S(\nbus_14035[0] ), .A(\tab12[2] ), .B(n_52389), .Z
		(n_10986));
	notech_reg_set tab12_reg_3(.CP(n_61744), .D(n_10992), .SD(n_61047), .Q(\tab12[3] 
		));
	notech_mux2 i_16390(.S(\nbus_14035[0] ), .A(\tab12[3] ), .B(n_52395), .Z
		(n_10992));
	notech_ao4 i_864(.A(n_1092), .B(n_13582), .C(n_1090), .D(n_13602), .Z(n_1116
		));
	notech_reg tab12_reg_4(.CP(n_61743), .D(n_10998), .CD(n_61046), .Q(\tab12[4] 
		));
	notech_mux2 i_16398(.S(\nbus_14035[0] ), .A(\tab12[4] ), .B(n_973), .Z(n_10998
		));
	notech_reg_set tab12_reg_5(.CP(n_61743), .D(n_11004), .SD(n_61046), .Q(\tab12[5] 
		));
	notech_mux2 i_16406(.S(\nbus_14035[0] ), .A(\tab12[5] ), .B(n_52407), .Z
		(n_11004));
	notech_and4 i_868(.A(n_1116), .B(n_1114), .C(n_876), .D(n_879), .Z(n_1118
		));
	notech_reg_set tab12_reg_6(.CP(n_61743), .D(n_11010), .SD(n_61046), .Q(\tab12[6] 
		));
	notech_mux2 i_16414(.S(\nbus_14035[0] ), .A(\tab12[6] ), .B(n_52413), .Z
		(n_11010));
	notech_ao4 i_861(.A(n_1100), .B(n_13509), .C(n_1098), .D(n_13676), .Z(n_1119
		));
	notech_reg_set tab12_reg_7(.CP(n_61743), .D(n_11016), .SD(n_61046), .Q(\tab12[7] 
		));
	notech_mux2 i_16422(.S(\nbus_14035[0] ), .A(\tab12[7] ), .B(n_52419), .Z
		(n_11016));
	notech_reg_set tab12_reg_8(.CP(n_61745), .D(n_11022), .SD(n_61048), .Q(\tab12[8] 
		));
	notech_mux2 i_16430(.S(\nbus_14035[0] ), .A(\tab12[8] ), .B(n_52425), .Z
		(n_11022));
	notech_ao4 i_860(.A(n_61599), .B(n_13752), .C(n_1043), .D(n_13677), .Z(n_1121
		));
	notech_reg_set tab12_reg_9(.CP(n_61744), .D(n_11028), .SD(n_61047), .Q(\tab12[9] 
		));
	notech_mux2 i_16438(.S(\nbus_14035[0] ), .A(\tab12[9] ), .B(n_52431), .Z
		(n_11028));
	notech_reg_set tab12_reg_10(.CP(n_61745), .D(n_11034), .SD(n_61048), .Q(\tab12[10] 
		));
	notech_mux2 i_16446(.S(\nbus_14035[0] ), .A(\tab12[10] ), .B(n_52437), .Z
		(n_11034));
	notech_ao4 i_857(.A(n_1086), .B(n_13531), .C(n_1084), .D(n_13560), .Z(n_1123
		));
	notech_reg_set tab12_reg_11(.CP(n_61745), .D(n_11040), .SD(n_61048), .Q(\tab12[11] 
		));
	notech_mux2 i_16454(.S(\nbus_14035[0] ), .A(\tab12[11] ), .B(n_52443), .Z
		(n_11040));
	notech_reg_set tab12_reg_12(.CP(n_61744), .D(n_11046), .SD(n_61047), .Q(\tab12[12] 
		));
	notech_mux2 i_16462(.S(\nbus_14035[0] ), .A(\tab12[12] ), .B(n_52449), .Z
		(n_11046));
	notech_ao4 i_855(.A(n_1092), .B(n_13581), .C(n_1090), .D(n_13601), .Z(n_1125
		));
	notech_reg_set tab12_reg_13(.CP(n_61744), .D(n_11052), .SD(n_61047), .Q(\tab12[13] 
		));
	notech_mux2 i_16470(.S(\nbus_14035[0] ), .A(\tab12[13] ), .B(n_52455), .Z
		(n_11052));
	notech_reg_set tab12_reg_14(.CP(n_61744), .D(n_11058), .SD(n_61047), .Q(\tab12[14] 
		));
	notech_mux2 i_16478(.S(\nbus_14035[0] ), .A(\tab12[14] ), .B(n_52461), .Z
		(n_11058));
	notech_and4 i_859(.A(n_1125), .B(n_1123), .C(n_865), .D(n_868), .Z(n_1127
		));
	notech_reg_set tab12_reg_15(.CP(n_61744), .D(n_11064), .SD(n_61047), .Q(\tab12[15] 
		));
	notech_mux2 i_16486(.S(\nbus_14035[0] ), .A(\tab12[15] ), .B(n_52467), .Z
		(n_11064));
	notech_ao4 i_852(.A(n_1100), .B(n_13508), .C(n_1098), .D(n_13674), .Z(n_1128
		));
	notech_reg_set tab12_reg_16(.CP(n_61744), .D(n_11070), .SD(n_61047), .Q(\tab12[16] 
		));
	notech_mux2 i_16494(.S(\nbus_14035[0] ), .A(\tab12[16] ), .B(n_52473), .Z
		(n_11070));
	notech_reg_set tab12_reg_17(.CP(n_61772), .D(n_11076), .SD(n_61075), .Q(\tab12[17] 
		));
	notech_mux2 i_16502(.S(n_54561), .A(\tab12[17] ), .B(n_52479), .Z(n_11076
		));
	notech_ao4 i_851(.A(n_61599), .B(n_13751), .C(n_1043), .D(n_13675), .Z(n_1130
		));
	notech_reg_set tab12_reg_18(.CP(n_61772), .D(n_11082), .SD(n_61075), .Q(\tab12[18] 
		));
	notech_mux2 i_16510(.S(n_54561), .A(\tab12[18] ), .B(n_52485), .Z(n_11082
		));
	notech_reg_set tab12_reg_19(.CP(n_61772), .D(n_11088), .SD(n_61075), .Q(\tab12[19] 
		));
	notech_mux2 i_16518(.S(n_54561), .A(\tab12[19] ), .B(n_52491), .Z(n_11088
		));
	notech_ao4 i_848(.A(n_1086), .B(n_13530), .C(n_1084), .D(n_13559), .Z(n_1132
		));
	notech_reg_set tab12_reg_20(.CP(n_61772), .D(n_11094), .SD(n_61075), .Q(\tab12[20] 
		));
	notech_mux2 i_16526(.S(n_54561), .A(\tab12[20] ), .B(n_52497), .Z(n_11094
		));
	notech_reg_set tab12_reg_21(.CP(n_61772), .D(n_11100), .SD(n_61075), .Q(\tab12[21] 
		));
	notech_mux2 i_16534(.S(n_54561), .A(\tab12[21] ), .B(n_52503), .Z(n_11100
		));
	notech_ao4 i_846(.A(n_1092), .B(n_13580), .C(n_1090), .D(n_13600), .Z(n_1134
		));
	notech_reg_set tab12_reg_22(.CP(n_61772), .D(n_11106), .SD(n_61075), .Q(\tab12[22] 
		));
	notech_mux2 i_16542(.S(n_54561), .A(\tab12[22] ), .B(n_52509), .Z(n_11106
		));
	notech_reg_set tab12_reg_23(.CP(n_61772), .D(n_11112), .SD(n_61075), .Q(\tab12[23] 
		));
	notech_mux2 i_16550(.S(n_54561), .A(\tab12[23] ), .B(n_52515), .Z(n_11112
		));
	notech_and4 i_850(.A(n_1134), .B(n_1132), .C(n_854), .D(n_857), .Z(n_1136
		));
	notech_reg_set tab12_reg_24(.CP(n_61772), .D(n_11118), .SD(n_61075), .Q(\tab12[24] 
		));
	notech_mux2 i_16558(.S(n_54561), .A(\tab12[24] ), .B(n_52521), .Z(n_11118
		));
	notech_ao4 i_843(.A(n_1100), .B(n_13507), .C(n_1098), .D(n_13672), .Z(n_1137
		));
	notech_reg_set tab12_reg_25(.CP(n_61772), .D(n_11124), .SD(n_61075), .Q(\tab12[25] 
		));
	notech_mux2 i_16566(.S(n_54561), .A(\tab12[25] ), .B(n_52527), .Z(n_11124
		));
	notech_reg_set tab12_reg_26(.CP(n_61773), .D(n_11130), .SD(n_61076), .Q(\tab12[26] 
		));
	notech_mux2 i_16574(.S(n_54561), .A(\tab12[26] ), .B(n_52533), .Z(n_11130
		));
	notech_ao4 i_842(.A(n_61599), .B(n_13750), .C(n_1043), .D(n_13673), .Z(n_1139
		));
	notech_reg_set tab12_reg_27(.CP(n_61773), .D(n_11136), .SD(n_61076), .Q(\tab12[27] 
		));
	notech_mux2 i_16582(.S(\nbus_14035[0] ), .A(\tab12[27] ), .B(n_52539), .Z
		(n_11136));
	notech_reg_set tab12_reg_28(.CP(n_61773), .D(n_11142), .SD(n_61076), .Q(\tab12[28] 
		));
	notech_mux2 i_16590(.S(n_54561), .A(\tab12[28] ), .B(n_52545), .Z(n_11142
		));
	notech_ao4 i_839(.A(n_1086), .B(n_13529), .C(n_1084), .D(n_13558), .Z(n_1141
		));
	notech_reg_set tab12_reg_29(.CP(n_61773), .D(n_11148), .SD(n_61076), .Q(\tab12[29] 
		));
	notech_mux2 i_16598(.S(n_54561), .A(\tab12[29] ), .B(n_52551), .Z(n_11148
		));
	notech_reg tab12_reg_30(.CP(n_61773), .D(n_11154), .CD(n_61076), .Q(\tab12[30] 
		));
	notech_mux2 i_16606(.S(n_54561), .A(\tab12[30] ), .B(n_974), .Z(n_11154)
		);
	notech_ao4 i_837(.A(n_1092), .B(n_13579), .C(n_1090), .D(n_13599), .Z(n_1143
		));
	notech_reg tab12_reg_32(.CP(n_61772), .D(n_11160), .CD(n_61075), .Q(\tab12[32] 
		));
	notech_mux2 i_16614(.S(n_54561), .A(\tab12[32] ), .B(n_975), .Z(n_11160)
		);
	notech_reg_set tab12_reg_33(.CP(n_61772), .D(n_11166), .SD(n_61075), .Q(\tab12[33] 
		));
	notech_mux2 i_16622(.S(n_54561), .A(\tab12[33] ), .B(n_54613), .Z(n_11166
		));
	notech_and4 i_841(.A(n_1143), .B(n_1141), .C(n_843), .D(n_846), .Z(n_1145
		));
	notech_reg hit_adr12_reg(.CP(n_61773), .D(n_11172), .CD(n_61076), .Q(hit_adr12
		));
	notech_mux2 i_16630(.S(n_971), .A(hit_add12), .B(hit_adr12), .Z(n_11172)
		);
	notech_ao4 i_834(.A(n_1100), .B(n_13506), .C(n_1098), .D(n_13670), .Z(n_1146
		));
	notech_reg_set tab13_reg_0(.CP(n_61773), .D(n_11178), .SD(n_61076), .Q(\tab13[0] 
		));
	notech_mux2 i_16638(.S(\nbus_14015[0] ), .A(\tab13[0] ), .B(n_52377), .Z
		(n_11178));
	notech_reg_set tab13_reg_1(.CP(n_61768), .D(n_11184), .SD(n_61071), .Q(\tab13[1] 
		));
	notech_mux2 i_16646(.S(\nbus_14015[0] ), .A(\tab13[1] ), .B(n_52383), .Z
		(n_11184));
	notech_ao4 i_833(.A(n_61599), .B(n_13749), .C(n_1043), .D(n_13671), .Z(n_1148
		));
	notech_reg_set tab13_reg_2(.CP(n_61768), .D(n_11190), .SD(n_61071), .Q(\tab13[2] 
		));
	notech_mux2 i_16654(.S(\nbus_14015[0] ), .A(\tab13[2] ), .B(n_52389), .Z
		(n_11190));
	notech_reg_set tab13_reg_3(.CP(n_61771), .D(n_11196), .SD(n_61074), .Q(\tab13[3] 
		));
	notech_mux2 i_16662(.S(\nbus_14015[0] ), .A(\tab13[3] ), .B(n_52395), .Z
		(n_11196));
	notech_ao4 i_830(.A(n_1086), .B(n_13528), .C(n_1084), .D(n_13557), .Z(n_1150
		));
	notech_reg tab13_reg_4(.CP(n_61771), .D(n_11202), .CD(n_61074), .Q(\tab13[4] 
		));
	notech_mux2 i_16670(.S(\nbus_14015[0] ), .A(\tab13[4] ), .B(n_973), .Z(n_11202
		));
	notech_reg_set tab13_reg_5(.CP(n_61768), .D(n_11208), .SD(n_61071), .Q(\tab13[5] 
		));
	notech_mux2 i_16678(.S(\nbus_14015[0] ), .A(\tab13[5] ), .B(n_52407), .Z
		(n_11208));
	notech_ao4 i_828(.A(n_1092), .B(n_13578), .C(n_1090), .D(n_13598), .Z(n_1152
		));
	notech_reg_set tab13_reg_6(.CP(n_61768), .D(n_11214), .SD(n_61071), .Q(\tab13[6] 
		));
	notech_mux2 i_16686(.S(\nbus_14015[0] ), .A(\tab13[6] ), .B(n_52413), .Z
		(n_11214));
	notech_reg_set tab13_reg_7(.CP(n_61768), .D(n_11220), .SD(n_61071), .Q(\tab13[7] 
		));
	notech_mux2 i_16694(.S(\nbus_14015[0] ), .A(\tab13[7] ), .B(n_52419), .Z
		(n_11220));
	notech_and4 i_832(.A(n_1152), .B(n_1150), .C(n_832), .D(n_835), .Z(n_1154
		));
	notech_reg_set tab13_reg_8(.CP(n_61768), .D(n_11226), .SD(n_61071), .Q(\tab13[8] 
		));
	notech_mux2 i_16702(.S(\nbus_14015[0] ), .A(\tab13[8] ), .B(n_52425), .Z
		(n_11226));
	notech_ao4 i_825(.A(n_1100), .B(n_13505), .C(n_1098), .D(n_13668), .Z(n_1155
		));
	notech_reg_set tab13_reg_9(.CP(n_61768), .D(n_11232), .SD(n_61071), .Q(\tab13[9] 
		));
	notech_mux2 i_16710(.S(\nbus_14015[0] ), .A(\tab13[9] ), .B(n_52431), .Z
		(n_11232));
	notech_reg_set tab13_reg_10(.CP(n_61771), .D(n_11238), .SD(n_61074), .Q(\tab13[10] 
		));
	notech_mux2 i_16718(.S(\nbus_14015[0] ), .A(\tab13[10] ), .B(n_52437), .Z
		(n_11238));
	notech_ao4 i_824(.A(n_61599), .B(n_13748), .C(n_1043), .D(n_13669), .Z(n_1157
		));
	notech_reg_set tab13_reg_11(.CP(n_61771), .D(n_11244), .SD(n_61074), .Q(\tab13[11] 
		));
	notech_mux2 i_16726(.S(\nbus_14015[0] ), .A(\tab13[11] ), .B(n_52443), .Z
		(n_11244));
	notech_reg_set tab13_reg_12(.CP(n_61771), .D(n_11250), .SD(n_61074), .Q(\tab13[12] 
		));
	notech_mux2 i_16734(.S(\nbus_14015[0] ), .A(\tab13[12] ), .B(n_52449), .Z
		(n_11250));
	notech_ao4 i_821(.A(n_1086), .B(n_13527), .C(n_1084), .D(n_13556), .Z(n_1159
		));
	notech_reg_set tab13_reg_13(.CP(n_61771), .D(n_11256), .SD(n_61074), .Q(\tab13[13] 
		));
	notech_mux2 i_16742(.S(\nbus_14015[0] ), .A(\tab13[13] ), .B(n_52455), .Z
		(n_11256));
	notech_reg_set tab13_reg_14(.CP(n_61771), .D(n_11262), .SD(n_61074), .Q(\tab13[14] 
		));
	notech_mux2 i_16750(.S(\nbus_14015[0] ), .A(\tab13[14] ), .B(n_52461), .Z
		(n_11262));
	notech_ao4 i_819(.A(n_1092), .B(n_13577), .C(n_1090), .D(n_13597), .Z(n_1161
		));
	notech_reg_set tab13_reg_15(.CP(n_61771), .D(n_11268), .SD(n_61074), .Q(\tab13[15] 
		));
	notech_mux2 i_16758(.S(\nbus_14015[0] ), .A(\tab13[15] ), .B(n_52467), .Z
		(n_11268));
	notech_reg_set tab13_reg_16(.CP(n_61771), .D(n_11274), .SD(n_61074), .Q(\tab13[16] 
		));
	notech_mux2 i_16766(.S(\nbus_14015[0] ), .A(\tab13[16] ), .B(n_52473), .Z
		(n_11274));
	notech_and4 i_823(.A(n_1161), .B(n_1159), .C(n_821), .D(n_824), .Z(n_1163
		));
	notech_reg_set tab13_reg_17(.CP(n_61771), .D(n_11280), .SD(n_61074), .Q(\tab13[17] 
		));
	notech_mux2 i_16774(.S(n_54543), .A(\tab13[17] ), .B(n_52479), .Z(n_11280
		));
	notech_ao4 i_816(.A(n_1100), .B(n_13504), .C(n_1098), .D(n_13666), .Z(n_1164
		));
	notech_reg_set tab13_reg_18(.CP(n_61771), .D(n_11286), .SD(n_61074), .Q(\tab13[18] 
		));
	notech_mux2 i_16782(.S(n_54543), .A(\tab13[18] ), .B(n_52485), .Z(n_11286
		));
	notech_reg_set tab13_reg_19(.CP(n_61773), .D(n_11292), .SD(n_61076), .Q(\tab13[19] 
		));
	notech_mux2 i_16790(.S(n_54543), .A(\tab13[19] ), .B(n_52491), .Z(n_11292
		));
	notech_ao4 i_815(.A(n_61599), .B(n_13747), .C(n_1043), .D(n_13667), .Z(n_1166
		));
	notech_reg_set tab13_reg_20(.CP(n_61776), .D(n_11298), .SD(n_61079), .Q(\tab13[20] 
		));
	notech_mux2 i_16798(.S(n_54543), .A(\tab13[20] ), .B(n_52497), .Z(n_11298
		));
	notech_reg_set tab13_reg_21(.CP(n_61776), .D(n_11304), .SD(n_61079), .Q(\tab13[21] 
		));
	notech_mux2 i_16806(.S(n_54543), .A(\tab13[21] ), .B(n_52503), .Z(n_11304
		));
	notech_ao4 i_812(.A(n_1086), .B(n_13526), .C(n_1084), .D(n_13555), .Z(n_1168
		));
	notech_reg_set tab13_reg_22(.CP(n_61777), .D(n_11310), .SD(n_61080), .Q(\tab13[22] 
		));
	notech_mux2 i_16814(.S(n_54543), .A(\tab13[22] ), .B(n_52509), .Z(n_11310
		));
	notech_reg_set tab13_reg_23(.CP(n_61777), .D(n_11316), .SD(n_61080), .Q(\tab13[23] 
		));
	notech_mux2 i_16822(.S(n_54543), .A(\tab13[23] ), .B(n_52515), .Z(n_11316
		));
	notech_ao4 i_810(.A(n_1092), .B(n_13576), .C(n_1090), .D(n_13596), .Z(n_1170
		));
	notech_reg_set tab13_reg_24(.CP(n_61776), .D(n_11322), .SD(n_61079), .Q(\tab13[24] 
		));
	notech_mux2 i_16830(.S(n_54543), .A(\tab13[24] ), .B(n_52521), .Z(n_11322
		));
	notech_reg_set tab13_reg_25(.CP(n_61776), .D(n_11328), .SD(n_61079), .Q(\tab13[25] 
		));
	notech_mux2 i_16838(.S(n_54543), .A(\tab13[25] ), .B(n_52527), .Z(n_11328
		));
	notech_and4 i_814(.A(n_1170), .B(n_1168), .C(n_810), .D(n_813), .Z(n_1172
		));
	notech_reg_set tab13_reg_26(.CP(n_61776), .D(n_11334), .SD(n_61079), .Q(\tab13[26] 
		));
	notech_mux2 i_16846(.S(n_54543), .A(\tab13[26] ), .B(n_52533), .Z(n_11334
		));
	notech_ao4 i_807(.A(n_1100), .B(n_13503), .C(n_1098), .D(n_13664), .Z(n_1173
		));
	notech_reg_set tab13_reg_27(.CP(n_61776), .D(n_11340), .SD(n_61079), .Q(\tab13[27] 
		));
	notech_mux2 i_16854(.S(\nbus_14015[0] ), .A(\tab13[27] ), .B(n_52539), .Z
		(n_11340));
	notech_reg_set tab13_reg_28(.CP(n_61776), .D(n_11346), .SD(n_61079), .Q(\tab13[28] 
		));
	notech_mux2 i_16862(.S(n_54543), .A(\tab13[28] ), .B(n_52545), .Z(n_11346
		));
	notech_ao4 i_806(.A(n_61599), .B(n_13746), .C(n_1043), .D(n_13665), .Z(n_1175
		));
	notech_reg_set tab13_reg_29(.CP(n_61777), .D(n_11352), .SD(n_61080), .Q(\tab13[29] 
		));
	notech_mux2 i_16870(.S(n_54543), .A(\tab13[29] ), .B(n_52551), .Z(n_11352
		));
	notech_reg tab13_reg_30(.CP(n_61777), .D(n_11358), .CD(n_61080), .Q(\tab13[30] 
		));
	notech_mux2 i_16878(.S(n_54543), .A(\tab13[30] ), .B(n_974), .Z(n_11358)
		);
	notech_ao4 i_803(.A(n_1086), .B(n_13525), .C(n_1084), .D(n_13554), .Z(n_1177
		));
	notech_reg tab13_reg_32(.CP(n_61777), .D(n_11364), .CD(n_61080), .Q(\tab13[32] 
		));
	notech_mux2 i_16886(.S(n_54543), .A(\tab13[32] ), .B(n_975), .Z(n_11364)
		);
	notech_reg_set tab13_reg_33(.CP(n_61777), .D(n_11370), .SD(n_61080), .Q(\tab13[33] 
		));
	notech_mux2 i_16894(.S(n_54543), .A(\tab13[33] ), .B(n_54613), .Z(n_11370
		));
	notech_ao4 i_801(.A(n_1092), .B(n_13575), .C(n_1090), .D(n_13595), .Z(n_1179
		));
	notech_reg hit_adr13_reg(.CP(n_61777), .D(n_11376), .CD(n_61080), .Q(hit_adr13
		));
	notech_mux2 i_16902(.S(n_971), .A(hit_add13), .B(hit_adr13), .Z(n_11376)
		);
	notech_reg_set tab14_reg_0(.CP(n_61777), .D(n_11382), .SD(n_61080), .Q(\tab14[0] 
		));
	notech_mux2 i_16910(.S(\nbus_14016[0] ), .A(\tab14[0] ), .B(n_52377), .Z
		(n_11382));
	notech_and4 i_805(.A(n_1179), .B(n_1177), .C(n_799), .D(n_802), .Z(n_1181
		));
	notech_reg_set tab14_reg_1(.CP(n_61777), .D(n_11388), .SD(n_61080), .Q(\tab14[1] 
		));
	notech_mux2 i_16918(.S(\nbus_14016[0] ), .A(\tab14[1] ), .B(n_52383), .Z
		(n_11388));
	notech_ao4 i_798(.A(n_1100), .B(n_13502), .C(n_1098), .D(n_13662), .Z(n_1182
		));
	notech_reg_set tab14_reg_2(.CP(n_61777), .D(n_11394), .SD(n_61080), .Q(\tab14[2] 
		));
	notech_mux2 i_16926(.S(\nbus_14016[0] ), .A(\tab14[2] ), .B(n_52389), .Z
		(n_11394));
	notech_reg_set tab14_reg_3(.CP(n_61777), .D(n_11400), .SD(n_61080), .Q(\tab14[3] 
		));
	notech_mux2 i_16934(.S(\nbus_14016[0] ), .A(\tab14[3] ), .B(n_52395), .Z
		(n_11400));
	notech_ao4 i_797(.A(n_61599), .B(n_13745), .C(n_54816), .D(n_13663), .Z(n_1184
		));
	notech_reg tab14_reg_4(.CP(n_61775), .D(n_11406), .CD(n_61078), .Q(\tab14[4] 
		));
	notech_mux2 i_16942(.S(\nbus_14016[0] ), .A(\tab14[4] ), .B(n_973), .Z(n_11406
		));
	notech_reg_set tab14_reg_5(.CP(n_61775), .D(n_11412), .SD(n_61078), .Q(\tab14[5] 
		));
	notech_mux2 i_16950(.S(\nbus_14016[0] ), .A(\tab14[5] ), .B(n_52407), .Z
		(n_11412));
	notech_ao4 i_794(.A(n_1086), .B(n_13524), .C(n_1084), .D(n_13553), .Z(n_1186
		));
	notech_reg_set tab14_reg_6(.CP(n_61775), .D(n_11418), .SD(n_61078), .Q(\tab14[6] 
		));
	notech_mux2 i_16958(.S(\nbus_14016[0] ), .A(\tab14[6] ), .B(n_52413), .Z
		(n_11418));
	notech_reg_set tab14_reg_7(.CP(n_61775), .D(n_11424), .SD(n_61078), .Q(\tab14[7] 
		));
	notech_mux2 i_16966(.S(\nbus_14016[0] ), .A(\tab14[7] ), .B(n_52419), .Z
		(n_11424));
	notech_ao4 i_792(.A(n_1092), .B(n_13574), .C(n_1090), .D(n_13594), .Z(n_1188
		));
	notech_reg_set tab14_reg_8(.CP(n_61775), .D(n_11430), .SD(n_61078), .Q(\tab14[8] 
		));
	notech_mux2 i_16974(.S(\nbus_14016[0] ), .A(\tab14[8] ), .B(n_52425), .Z
		(n_11430));
	notech_reg_set tab14_reg_9(.CP(n_61773), .D(n_11436), .SD(n_61076), .Q(\tab14[9] 
		));
	notech_mux2 i_16982(.S(\nbus_14016[0] ), .A(\tab14[9] ), .B(n_52431), .Z
		(n_11436));
	notech_and4 i_796(.A(n_1188), .B(n_1186), .C(n_788), .D(n_791), .Z(n_1190
		));
	notech_reg_set tab14_reg_10(.CP(n_61773), .D(n_11442), .SD(n_61076), .Q(\tab14[10] 
		));
	notech_mux2 i_16990(.S(\nbus_14016[0] ), .A(\tab14[10] ), .B(n_52437), .Z
		(n_11442));
	notech_ao4 i_788(.A(n_1100), .B(n_13501), .C(n_1098), .D(n_13660), .Z(n_1191
		));
	notech_reg_set tab14_reg_11(.CP(n_61775), .D(n_11448), .SD(n_61078), .Q(\tab14[11] 
		));
	notech_mux2 i_16998(.S(\nbus_14016[0] ), .A(\tab14[11] ), .B(n_52443), .Z
		(n_11448));
	notech_reg_set tab14_reg_12(.CP(n_61773), .D(n_11454), .SD(n_61076), .Q(\tab14[12] 
		));
	notech_mux2 i_17006(.S(\nbus_14016[0] ), .A(\tab14[12] ), .B(n_52449), .Z
		(n_11454));
	notech_ao4 i_787(.A(n_61604), .B(n_13744), .C(n_54816), .D(n_13661), .Z(n_1193
		));
	notech_reg_set tab14_reg_13(.CP(n_61776), .D(n_11460), .SD(n_61079), .Q(\tab14[13] 
		));
	notech_mux2 i_17014(.S(\nbus_14016[0] ), .A(\tab14[13] ), .B(n_52455), .Z
		(n_11460));
	notech_reg_set tab14_reg_14(.CP(n_61776), .D(n_11466), .SD(n_61079), .Q(\tab14[14] 
		));
	notech_mux2 i_17022(.S(\nbus_14016[0] ), .A(\tab14[14] ), .B(n_52461), .Z
		(n_11466));
	notech_ao4 i_784(.A(n_1086), .B(n_13523), .C(n_1084), .D(n_13552), .Z(n_1195
		));
	notech_reg_set tab14_reg_15(.CP(n_61776), .D(n_11472), .SD(n_61079), .Q(\tab14[15] 
		));
	notech_mux2 i_17030(.S(\nbus_14016[0] ), .A(\tab14[15] ), .B(n_52467), .Z
		(n_11472));
	notech_reg_set tab14_reg_16(.CP(n_61776), .D(n_11478), .SD(n_61079), .Q(\tab14[16] 
		));
	notech_mux2 i_17038(.S(\nbus_14016[0] ), .A(\tab14[16] ), .B(n_52473), .Z
		(n_11478));
	notech_ao4 i_782(.A(n_1092), .B(n_13573), .C(n_1090), .D(n_13593), .Z(n_1197
		));
	notech_reg_set tab14_reg_17(.CP(n_61775), .D(n_11484), .SD(n_61078), .Q(\tab14[17] 
		));
	notech_mux2 i_17046(.S(n_54534), .A(\tab14[17] ), .B(n_52479), .Z(n_11484
		));
	notech_reg_set tab14_reg_18(.CP(n_61775), .D(n_11490), .SD(n_61078), .Q(\tab14[18] 
		));
	notech_mux2 i_17054(.S(n_54534), .A(\tab14[18] ), .B(n_52485), .Z(n_11490
		));
	notech_and4 i_786(.A(n_1197), .B(n_1195), .C(n_777), .D(n_780), .Z(n_1199
		));
	notech_reg_set tab14_reg_19(.CP(n_61775), .D(n_11496), .SD(n_61078), .Q(\tab14[19] 
		));
	notech_mux2 i_17062(.S(n_54534), .A(\tab14[19] ), .B(n_52491), .Z(n_11496
		));
	notech_ao4 i_779(.A(n_1100), .B(n_13500), .C(n_1098), .D(n_13658), .Z(n_1200
		));
	notech_reg_set tab14_reg_20(.CP(n_61775), .D(n_11502), .SD(n_61078), .Q(\tab14[20] 
		));
	notech_mux2 i_17070(.S(n_54534), .A(\tab14[20] ), .B(n_52497), .Z(n_11502
		));
	notech_reg_set tab14_reg_21(.CP(n_61775), .D(n_11508), .SD(n_61078), .Q(\tab14[21] 
		));
	notech_mux2 i_17078(.S(n_54534), .A(\tab14[21] ), .B(n_52503), .Z(n_11508
		));
	notech_ao4 i_778(.A(n_61604), .B(n_13743), .C(n_54816), .D(n_13659), .Z(n_1202
		));
	notech_reg_set tab14_reg_22(.CP(n_61768), .D(n_11514), .SD(n_61071), .Q(\tab14[22] 
		));
	notech_mux2 i_17086(.S(n_54534), .A(\tab14[22] ), .B(n_52509), .Z(n_11514
		));
	notech_reg_set tab14_reg_23(.CP(n_61762), .D(n_11520), .SD(n_61065), .Q(\tab14[23] 
		));
	notech_mux2 i_17094(.S(n_54534), .A(\tab14[23] ), .B(n_52515), .Z(n_11520
		));
	notech_ao4 i_775(.A(n_1086), .B(n_13522), .C(n_1084), .D(n_13551), .Z(n_1204
		));
	notech_reg_set tab14_reg_24(.CP(n_61762), .D(n_11526), .SD(n_61065), .Q(\tab14[24] 
		));
	notech_mux2 i_17102(.S(n_54534), .A(\tab14[24] ), .B(n_52521), .Z(n_11526
		));
	notech_reg_set tab14_reg_25(.CP(n_61763), .D(n_11532), .SD(n_61066), .Q(\tab14[25] 
		));
	notech_mux2 i_17110(.S(n_54534), .A(\tab14[25] ), .B(n_52527), .Z(n_11532
		));
	notech_ao4 i_773(.A(n_1092), .B(n_13572), .C(n_1090), .D(n_13592), .Z(n_1206
		));
	notech_reg_set tab14_reg_26(.CP(n_61762), .D(n_11538), .SD(n_61065), .Q(\tab14[26] 
		));
	notech_mux2 i_17118(.S(n_54534), .A(\tab14[26] ), .B(n_52533), .Z(n_11538
		));
	notech_reg_set tab14_reg_27(.CP(n_61762), .D(n_11544), .SD(n_61065), .Q(\tab14[27] 
		));
	notech_mux2 i_17126(.S(\nbus_14016[0] ), .A(\tab14[27] ), .B(n_52539), .Z
		(n_11544));
	notech_and4 i_777(.A(n_1206), .B(n_1204), .C(n_766), .D(n_769), .Z(n_1208
		));
	notech_reg_set tab14_reg_28(.CP(n_61762), .D(n_11550), .SD(n_61065), .Q(\tab14[28] 
		));
	notech_mux2 i_17134(.S(n_54534), .A(\tab14[28] ), .B(n_52545), .Z(n_11550
		));
	notech_ao4 i_770(.A(n_1100), .B(n_13498), .C(n_1098), .D(n_13656), .Z(n_1209
		));
	notech_reg_set tab14_reg_29(.CP(n_61762), .D(n_11556), .SD(n_61065), .Q(\tab14[29] 
		));
	notech_mux2 i_17142(.S(n_54534), .A(\tab14[29] ), .B(n_52551), .Z(n_11556
		));
	notech_reg tab14_reg_30(.CP(n_61762), .D(n_11562), .CD(n_61065), .Q(\tab14[30] 
		));
	notech_mux2 i_17150(.S(n_54534), .A(\tab14[30] ), .B(n_974), .Z(n_11562)
		);
	notech_ao4 i_769(.A(n_61604), .B(n_13742), .C(n_54816), .D(n_13657), .Z(n_1211
		));
	notech_reg tab14_reg_32(.CP(n_61762), .D(n_11568), .CD(n_61065), .Q(\tab14[32] 
		));
	notech_mux2 i_17158(.S(n_54534), .A(\tab14[32] ), .B(n_975), .Z(n_11568)
		);
	notech_reg_set tab14_reg_33(.CP(n_61763), .D(n_11574), .SD(n_61066), .Q(\tab14[33] 
		));
	notech_mux2 i_17166(.S(n_54534), .A(\tab14[33] ), .B(n_54613), .Z(n_11574
		));
	notech_ao4 i_766(.A(n_1086), .B(n_13521), .C(n_1084), .D(n_13550), .Z(n_1213
		));
	notech_reg hit_adr14_reg(.CP(n_61763), .D(n_11580), .CD(n_61066), .Q(hit_adr14
		));
	notech_mux2 i_17174(.S(n_971), .A(hit_add14), .B(hit_adr14), .Z(n_11580)
		);
	notech_reg nx_tab1_reg_0(.CP(n_61763), .D(n_11586), .CD(n_61066), .Q(\nx_tab1[0] 
		));
	notech_mux2 i_17182(.S(\nbus_14041[0] ), .A(\nx_tab1[0] ), .B(n_13535), 
		.Z(n_11586));
	notech_ao4 i_764(.A(n_1092), .B(n_13571), .C(n_1090), .D(n_13591), .Z(n_1215
		));
	notech_reg nx_tab1_reg_1(.CP(n_61763), .D(n_11592), .CD(n_61066), .Q(\nx_tab1[1] 
		));
	notech_mux2 i_17190(.S(\nbus_14041[0] ), .A(\nx_tab1[1] ), .B(n_13537), 
		.Z(n_11592));
	notech_reg_set nnx_tab1_reg_0(.CP(n_61763), .D(n_11598), .SD(n_61066), .Q
		(\nnx_tab1[0] ));
	notech_mux2 i_17198(.S(n_13543), .A(\nnx_tab1[0] ), .B(n_13539), .Z(n_11598
		));
	notech_and4 i_768(.A(n_1215), .B(n_1213), .C(n_755), .D(n_758), .Z(n_1217
		));
	notech_reg nnx_tab1_reg_1(.CP(n_61763), .D(n_11604), .CD(n_61066), .Q(\nnx_tab1[1] 
		));
	notech_mux2 i_17206(.S(n_13543), .A(\nnx_tab1[1] ), .B(n_13541), .Z(n_11604
		));
	notech_ao4 i_761(.A(n_1100), .B(n_13497), .C(n_1098), .D(n_13654), .Z(n_1218
		));
	notech_reg hit_adr21_reg(.CP(n_61763), .D(n_11610), .CD(n_61066), .Q(hit_adr21
		));
	notech_mux2 i_17214(.S(n_971), .A(hit_add21), .B(hit_adr21), .Z(n_11610)
		);
	notech_reg_set tab22_reg_0(.CP(n_61763), .D(n_11616), .SD(n_61066), .Q(\tab22[0] 
		));
	notech_mux2 i_17222(.S(\nbus_14037[0] ), .A(\tab22[0] ), .B(n_52377), .Z
		(n_11616));
	notech_ao4 i_760(.A(n_61604), .B(n_13741), .C(n_54816), .D(n_13655), .Z(n_1220
		));
	notech_reg_set tab22_reg_1(.CP(n_61763), .D(n_11622), .SD(n_61066), .Q(\tab22[1] 
		));
	notech_mux2 i_17230(.S(\nbus_14037[0] ), .A(\tab22[1] ), .B(n_52383), .Z
		(n_11622));
	notech_reg_set tab22_reg_2(.CP(n_61759), .D(n_11628), .SD(n_61062), .Q(\tab22[2] 
		));
	notech_mux2 i_17238(.S(\nbus_14037[0] ), .A(\tab22[2] ), .B(n_52389), .Z
		(n_11628));
	notech_ao4 i_757(.A(n_1086), .B(n_13520), .C(n_1084), .D(n_13549), .Z(n_1222
		));
	notech_reg_set tab22_reg_3(.CP(n_61759), .D(n_11634), .SD(n_61062), .Q(\tab22[3] 
		));
	notech_mux2 i_17246(.S(\nbus_14037[0] ), .A(\tab22[3] ), .B(n_52395), .Z
		(n_11634));
	notech_reg tab22_reg_4(.CP(n_61759), .D(n_11640), .CD(n_61062), .Q(\tab22[4] 
		));
	notech_mux2 i_17254(.S(\nbus_14037[0] ), .A(\tab22[4] ), .B(n_973), .Z(n_11640
		));
	notech_ao4 i_755(.A(n_1092), .B(n_13570), .C(n_1090), .D(n_13590), .Z(n_1224
		));
	notech_reg_set tab22_reg_5(.CP(n_61759), .D(n_11646), .SD(n_61062), .Q(\tab22[5] 
		));
	notech_mux2 i_17262(.S(\nbus_14037[0] ), .A(\tab22[5] ), .B(n_52407), .Z
		(n_11646));
	notech_reg_set tab22_reg_6(.CP(n_61759), .D(n_11652), .SD(n_61062), .Q(\tab22[6] 
		));
	notech_mux2 i_17270(.S(\nbus_14037[0] ), .A(\tab22[6] ), .B(n_52413), .Z
		(n_11652));
	notech_and4 i_759(.A(n_1224), .B(n_1222), .C(n_744), .D(n_747), .Z(n_1226
		));
	notech_reg_set tab22_reg_7(.CP(n_61758), .D(n_11658), .SD(n_61061), .Q(\tab22[7] 
		));
	notech_mux2 i_17278(.S(\nbus_14037[0] ), .A(\tab22[7] ), .B(n_52419), .Z
		(n_11658));
	notech_ao4 i_752(.A(n_1100), .B(n_13496), .C(n_1098), .D(n_13652), .Z(n_1227
		));
	notech_reg_set tab22_reg_8(.CP(n_61758), .D(n_11664), .SD(n_61061), .Q(\tab22[8] 
		));
	notech_mux2 i_17286(.S(\nbus_14037[0] ), .A(\tab22[8] ), .B(n_52425), .Z
		(n_11664));
	notech_reg_set tab22_reg_9(.CP(n_61758), .D(n_11670), .SD(n_61061), .Q(\tab22[9] 
		));
	notech_mux2 i_17294(.S(\nbus_14037[0] ), .A(\tab22[9] ), .B(n_52431), .Z
		(n_11670));
	notech_ao4 i_751(.A(n_61604), .B(n_13740), .C(n_54816), .D(n_13653), .Z(n_1229
		));
	notech_reg_set tab22_reg_10(.CP(n_61758), .D(n_11676), .SD(n_61061), .Q(\tab22[10] 
		));
	notech_mux2 i_17302(.S(\nbus_14037[0] ), .A(\tab22[10] ), .B(n_52437), .Z
		(n_11676));
	notech_reg_set tab22_reg_11(.CP(n_61762), .D(n_11682), .SD(n_61065), .Q(\tab22[11] 
		));
	notech_mux2 i_17310(.S(\nbus_14037[0] ), .A(\tab22[11] ), .B(n_52443), .Z
		(n_11682));
	notech_ao4 i_748(.A(n_1086), .B(n_13519), .C(n_1084), .D(n_13548), .Z(n_1231
		));
	notech_reg_set tab22_reg_12(.CP(n_61759), .D(n_11688), .SD(n_61062), .Q(\tab22[12] 
		));
	notech_mux2 i_17318(.S(\nbus_14037[0] ), .A(\tab22[12] ), .B(n_52449), .Z
		(n_11688));
	notech_reg_set tab22_reg_13(.CP(n_61762), .D(n_11694), .SD(n_61065), .Q(\tab22[13] 
		));
	notech_mux2 i_17326(.S(\nbus_14037[0] ), .A(\tab22[13] ), .B(n_52455), .Z
		(n_11694));
	notech_ao4 i_746(.A(n_1092), .B(n_13569), .C(n_1090), .D(n_13589), .Z(n_1233
		));
	notech_reg_set tab22_reg_14(.CP(n_61762), .D(n_11700), .SD(n_61065), .Q(\tab22[14] 
		));
	notech_mux2 i_17334(.S(\nbus_14037[0] ), .A(\tab22[14] ), .B(n_52461), .Z
		(n_11700));
	notech_reg_set tab22_reg_15(.CP(n_61759), .D(n_11706), .SD(n_61062), .Q(\tab22[15] 
		));
	notech_mux2 i_17342(.S(\nbus_14037[0] ), .A(\tab22[15] ), .B(n_52467), .Z
		(n_11706));
	notech_and4 i_750(.A(n_1233), .B(n_1231), .C(n_733), .D(n_736), .Z(n_1235
		));
	notech_reg_set tab22_reg_16(.CP(n_61759), .D(n_11712), .SD(n_61062), .Q(\tab22[16] 
		));
	notech_mux2 i_17350(.S(\nbus_14037[0] ), .A(\tab22[16] ), .B(n_52473), .Z
		(n_11712));
	notech_ao4 i_743(.A(n_1100), .B(n_13495), .C(n_1098), .D(n_13650), .Z(n_1236
		));
	notech_reg_set tab22_reg_17(.CP(n_61759), .D(n_11718), .SD(n_61062), .Q(\tab22[17] 
		));
	notech_mux2 i_17358(.S(n_54619), .A(\tab22[17] ), .B(n_52479), .Z(n_11718
		));
	notech_reg_set tab22_reg_18(.CP(n_61759), .D(n_11724), .SD(n_61062), .Q(\tab22[18] 
		));
	notech_mux2 i_17366(.S(n_54619), .A(\tab22[18] ), .B(n_52485), .Z(n_11724
		));
	notech_ao4 i_742(.A(n_61604), .B(n_13739), .C(n_54816), .D(n_13651), .Z(n_1238
		));
	notech_reg_set tab22_reg_19(.CP(n_61759), .D(n_11730), .SD(n_61062), .Q(\tab22[19] 
		));
	notech_mux2 i_17374(.S(n_54619), .A(\tab22[19] ), .B(n_52491), .Z(n_11730
		));
	notech_reg_set tab22_reg_20(.CP(n_61763), .D(n_11736), .SD(n_61066), .Q(\tab22[20] 
		));
	notech_mux2 i_17382(.S(n_54619), .A(\tab22[20] ), .B(n_52497), .Z(n_11736
		));
	notech_ao4 i_739(.A(n_1086), .B(n_13518), .C(n_1084), .D(n_13547), .Z(n_1240
		));
	notech_reg_set tab22_reg_21(.CP(n_61767), .D(n_11742), .SD(n_61070), .Q(\tab22[21] 
		));
	notech_mux2 i_17390(.S(n_54619), .A(\tab22[21] ), .B(n_52503), .Z(n_11742
		));
	notech_reg_set tab22_reg_22(.CP(n_61767), .D(n_11748), .SD(n_61070), .Q(\tab22[22] 
		));
	notech_mux2 i_17398(.S(n_54619), .A(\tab22[22] ), .B(n_52509), .Z(n_11748
		));
	notech_ao4 i_737(.A(n_1092), .B(n_13568), .C(n_1090), .D(n_13588), .Z(n_1242
		));
	notech_reg_set tab22_reg_23(.CP(n_61767), .D(n_11754), .SD(n_61070), .Q(\tab22[23] 
		));
	notech_mux2 i_17406(.S(n_54619), .A(\tab22[23] ), .B(n_52515), .Z(n_11754
		));
	notech_reg_set tab22_reg_24(.CP(n_61767), .D(n_11760), .SD(n_61070), .Q(\tab22[24] 
		));
	notech_mux2 i_17414(.S(n_54619), .A(\tab22[24] ), .B(n_52521), .Z(n_11760
		));
	notech_and4 i_741(.A(n_1242), .B(n_1240), .C(n_722), .D(n_725), .Z(n_1244
		));
	notech_reg_set tab22_reg_25(.CP(n_61767), .D(n_11766), .SD(n_61070), .Q(\tab22[25] 
		));
	notech_mux2 i_17422(.S(n_54619), .A(\tab22[25] ), .B(n_52527), .Z(n_11766
		));
	notech_ao4 i_734(.A(n_1100), .B(n_13494), .C(n_53455), .D(n_13648), .Z(n_1245
		));
	notech_reg_set tab22_reg_26(.CP(n_61766), .D(n_11772), .SD(n_61069), .Q(\tab22[26] 
		));
	notech_mux2 i_17430(.S(n_54619), .A(\tab22[26] ), .B(n_52533), .Z(n_11772
		));
	notech_reg_set tab22_reg_27(.CP(n_61766), .D(n_11778), .SD(n_61069), .Q(\tab22[27] 
		));
	notech_mux2 i_17438(.S(\nbus_14037[0] ), .A(\tab22[27] ), .B(n_52539), .Z
		(n_11778));
	notech_ao4 i_733(.A(n_61604), .B(n_13738), .C(n_1043), .D(n_13649), .Z(n_1247
		));
	notech_reg_set tab22_reg_28(.CP(n_61766), .D(n_11784), .SD(n_61069), .Q(\tab22[28] 
		));
	notech_mux2 i_17446(.S(n_54619), .A(\tab22[28] ), .B(n_52545), .Z(n_11784
		));
	notech_reg_set tab22_reg_29(.CP(n_61766), .D(n_11790), .SD(n_61069), .Q(\tab22[29] 
		));
	notech_mux2 i_17454(.S(n_54619), .A(\tab22[29] ), .B(n_52551), .Z(n_11790
		));
	notech_ao4 i_730(.A(n_1086), .B(n_13517), .C(n_1084), .D(n_13546), .Z(n_1249
		));
	notech_reg tab22_reg_30(.CP(n_61768), .D(n_11796), .CD(n_61071), .Q(\tab22[30] 
		));
	notech_mux2 i_17462(.S(n_54619), .A(\tab22[30] ), .B(n_974), .Z(n_11796)
		);
	notech_reg tab22_reg_32(.CP(n_61767), .D(n_11802), .CD(n_61070), .Q(\tab22[32] 
		));
	notech_mux2 i_17470(.S(n_54619), .A(\tab22[32] ), .B(n_975), .Z(n_11802)
		);
	notech_ao4 i_728(.A(n_1092), .B(n_13567), .C(n_1090), .D(n_13587), .Z(n_1251
		));
	notech_reg_set tab22_reg_33(.CP(n_61768), .D(n_11808), .SD(n_61071), .Q(\tab22[33] 
		));
	notech_mux2 i_17478(.S(n_54619), .A(\tab22[33] ), .B(n_54613), .Z(n_11808
		));
	notech_reg hit_adr22_reg(.CP(n_61768), .D(n_11814), .CD(n_61071), .Q(hit_adr22
		));
	notech_mux2 i_17486(.S(n_971), .A(hit_add22), .B(hit_adr22), .Z(n_11814)
		);
	notech_and4 i_732(.A(n_1251), .B(n_1249), .C(n_711), .D(n_714), .Z(n_1253
		));
	notech_reg_set tab23_reg_0(.CP(n_61767), .D(n_11820), .SD(n_61070), .Q(\tab23[0] 
		));
	notech_mux2 i_17494(.S(\nbus_14017[0] ), .A(\tab23[0] ), .B(n_52377), .Z
		(n_11820));
	notech_ao4 i_725(.A(n_1100), .B(n_13493), .C(n_53455), .D(n_13646), .Z(n_1254
		));
	notech_reg_set tab23_reg_1(.CP(n_61767), .D(n_11826), .SD(n_61070), .Q(\tab23[1] 
		));
	notech_mux2 i_17502(.S(\nbus_14017[0] ), .A(\tab23[1] ), .B(n_52383), .Z
		(n_11826));
	notech_reg_set tab23_reg_2(.CP(n_61767), .D(n_11832), .SD(n_61070), .Q(\tab23[2] 
		));
	notech_mux2 i_17510(.S(\nbus_14017[0] ), .A(\tab23[2] ), .B(n_52389), .Z
		(n_11832));
	notech_ao4 i_724(.A(n_61604), .B(n_13737), .C(n_54816), .D(n_13647), .Z(n_1256
		));
	notech_reg_set tab23_reg_3(.CP(n_61767), .D(n_11838), .SD(n_61070), .Q(\tab23[3] 
		));
	notech_mux2 i_17518(.S(\nbus_14017[0] ), .A(\tab23[3] ), .B(n_52395), .Z
		(n_11838));
	notech_reg tab23_reg_4(.CP(n_61767), .D(n_11844), .CD(n_61070), .Q(\tab23[4] 
		));
	notech_mux2 i_17526(.S(\nbus_14017[0] ), .A(\tab23[4] ), .B(n_973), .Z(n_11844
		));
	notech_ao4 i_721(.A(n_1086), .B(n_13516), .C(n_1084), .D(n_13545), .Z(n_1258
		));
	notech_reg_set tab23_reg_5(.CP(n_61764), .D(n_11850), .SD(n_61067), .Q(\tab23[5] 
		));
	notech_mux2 i_17534(.S(\nbus_14017[0] ), .A(\tab23[5] ), .B(n_52407), .Z
		(n_11850));
	notech_reg_set tab23_reg_6(.CP(n_61764), .D(n_11856), .SD(n_61067), .Q(\tab23[6] 
		));
	notech_mux2 i_17542(.S(\nbus_14017[0] ), .A(\tab23[6] ), .B(n_52413), .Z
		(n_11856));
	notech_ao4 i_719(.A(n_1092), .B(n_13566), .C(n_1090), .D(n_13586), .Z(n_1260
		));
	notech_reg_set tab23_reg_7(.CP(n_61764), .D(n_11862), .SD(n_61067), .Q(\tab23[7] 
		));
	notech_mux2 i_17550(.S(\nbus_14017[0] ), .A(\tab23[7] ), .B(n_52419), .Z
		(n_11862));
	notech_reg_set tab23_reg_8(.CP(n_61764), .D(n_11868), .SD(n_61067), .Q(\tab23[8] 
		));
	notech_mux2 i_17558(.S(\nbus_14017[0] ), .A(\tab23[8] ), .B(n_52425), .Z
		(n_11868));
	notech_and4 i_723(.A(n_1260), .B(n_1258), .C(n_700), .D(n_703), .Z(n_1262
		));
	notech_reg_set tab23_reg_9(.CP(n_61764), .D(n_11874), .SD(n_61067), .Q(\tab23[9] 
		));
	notech_mux2 i_17566(.S(\nbus_14017[0] ), .A(\tab23[9] ), .B(n_52431), .Z
		(n_11874));
	notech_ao4 i_716(.A(n_1100), .B(n_13492), .C(n_53455), .D(n_13644), .Z(n_1263
		));
	notech_reg_set tab23_reg_10(.CP(n_61764), .D(n_11880), .SD(n_61067), .Q(\tab23[10] 
		));
	notech_mux2 i_17574(.S(\nbus_14017[0] ), .A(\tab23[10] ), .B(n_52437), .Z
		(n_11880));
	notech_reg_set tab23_reg_11(.CP(n_61764), .D(n_11886), .SD(n_61067), .Q(\tab23[11] 
		));
	notech_mux2 i_17582(.S(\nbus_14017[0] ), .A(\tab23[11] ), .B(n_52443), .Z
		(n_11886));
	notech_ao4 i_715(.A(n_61604), .B(n_13736), .C(n_54816), .D(n_13645), .Z(n_1265
		));
	notech_reg_set tab23_reg_12(.CP(n_61764), .D(n_11892), .SD(n_61067), .Q(\tab23[12] 
		));
	notech_mux2 i_17590(.S(\nbus_14017[0] ), .A(\tab23[12] ), .B(n_52449), .Z
		(n_11892));
	notech_reg_set tab23_reg_13(.CP(n_61764), .D(n_11898), .SD(n_61067), .Q(\tab23[13] 
		));
	notech_mux2 i_17598(.S(\nbus_14017[0] ), .A(\tab23[13] ), .B(n_52455), .Z
		(n_11898));
	notech_ao4 i_712(.A(n_1086), .B(n_13515), .C(n_1084), .D(n_13544), .Z(n_1267
		));
	notech_reg_set tab23_reg_14(.CP(n_61766), .D(n_11904), .SD(n_61069), .Q(\tab23[14] 
		));
	notech_mux2 i_17606(.S(\nbus_14017[0] ), .A(\tab23[14] ), .B(n_52461), .Z
		(n_11904));
	notech_reg_set tab23_reg_15(.CP(n_61766), .D(n_11910), .SD(n_61069), .Q(\tab23[15] 
		));
	notech_mux2 i_17614(.S(\nbus_14017[0] ), .A(\tab23[15] ), .B(n_52467), .Z
		(n_11910));
	notech_ao4 i_710(.A(n_1092), .B(n_13565), .C(n_1090), .D(n_13585), .Z(n_1269
		));
	notech_reg_set tab23_reg_16(.CP(n_61766), .D(n_11916), .SD(n_61069), .Q(\tab23[16] 
		));
	notech_mux2 i_17622(.S(\nbus_14017[0] ), .A(\tab23[16] ), .B(n_52473), .Z
		(n_11916));
	notech_reg_set tab23_reg_17(.CP(n_61766), .D(n_11922), .SD(n_61069), .Q(\tab23[17] 
		));
	notech_mux2 i_17630(.S(n_54581), .A(\tab23[17] ), .B(n_52479), .Z(n_11922
		));
	notech_and4 i_714(.A(n_1269), .B(n_1267), .C(n_692), .D(n_689), .Z(n_1271
		));
	notech_reg_set tab23_reg_18(.CP(n_61766), .D(n_11928), .SD(n_61069), .Q(\tab23[18] 
		));
	notech_mux2 i_17638(.S(n_54581), .A(\tab23[18] ), .B(n_52485), .Z(n_11928
		));
	notech_ao4 i_707(.A(n_1100), .B(n_13491), .C(n_53455), .D(n_13642), .Z(n_1272
		));
	notech_reg_set tab23_reg_19(.CP(n_61764), .D(n_11934), .SD(n_61067), .Q(\tab23[19] 
		));
	notech_mux2 i_17646(.S(n_54581), .A(\tab23[19] ), .B(n_52491), .Z(n_11934
		));
	notech_reg_set tab23_reg_20(.CP(n_61764), .D(n_11940), .SD(n_61067), .Q(\tab23[20] 
		));
	notech_mux2 i_17654(.S(n_54581), .A(\tab23[20] ), .B(n_52497), .Z(n_11940
		));
	notech_ao4 i_706(.A(n_61604), .B(n_13735), .C(n_54816), .D(n_13643), .Z(n_1274
		));
	notech_reg_set tab23_reg_21(.CP(n_61766), .D(n_11946), .SD(n_61069), .Q(\tab23[21] 
		));
	notech_mux2 i_17662(.S(n_54581), .A(\tab23[21] ), .B(n_52503), .Z(n_11946
		));
	notech_reg_set tab23_reg_22(.CP(n_61766), .D(n_11952), .SD(n_61069), .Q(\tab23[22] 
		));
	notech_mux2 i_17670(.S(n_54581), .A(\tab23[22] ), .B(n_52509), .Z(n_11952
		));
	notech_ao4 i_705(.A(n_53455), .B(n_13641), .C(n_486), .D(n_13734), .Z(n_1276
		));
	notech_reg_set tab23_reg_23(.CP(n_61738), .D(n_11958), .SD(n_61041), .Q(\tab23[23] 
		));
	notech_mux2 i_17678(.S(n_54581), .A(\tab23[23] ), .B(n_52515), .Z(n_11958
		));
	notech_ao4 i_704(.A(n_53455), .B(n_13640), .C(n_486), .D(n_13733), .Z(n_1277
		));
	notech_reg_set tab23_reg_24(.CP(n_61710), .D(n_11964), .SD(n_61013), .Q(\tab23[24] 
		));
	notech_mux2 i_17686(.S(n_54581), .A(\tab23[24] ), .B(n_52521), .Z(n_11964
		));
	notech_ao4 i_703(.A(n_53455), .B(n_13639), .C(n_486), .D(n_13732), .Z(n_1278
		));
	notech_reg_set tab23_reg_25(.CP(n_61710), .D(n_11970), .SD(n_61013), .Q(\tab23[25] 
		));
	notech_mux2 i_17694(.S(n_54581), .A(\tab23[25] ), .B(n_52527), .Z(n_11970
		));
	notech_ao4 i_702(.A(n_53455), .B(n_13638), .C(n_486), .D(n_13731), .Z(n_1279
		));
	notech_reg_set tab23_reg_26(.CP(n_61710), .D(n_11976), .SD(n_61013), .Q(\tab23[26] 
		));
	notech_mux2 i_17702(.S(n_54581), .A(\tab23[26] ), .B(n_52533), .Z(n_11976
		));
	notech_ao4 i_701(.A(n_53455), .B(n_13637), .C(n_486), .D(n_13730), .Z(n_1280
		));
	notech_reg_set tab23_reg_27(.CP(n_61710), .D(n_11982), .SD(n_61013), .Q(\tab23[27] 
		));
	notech_mux2 i_17710(.S(\nbus_14017[0] ), .A(\tab23[27] ), .B(n_52539), .Z
		(n_11982));
	notech_ao4 i_700(.A(n_53455), .B(n_13636), .C(n_486), .D(n_13729), .Z(n_1281
		));
	notech_reg_set tab23_reg_28(.CP(n_61710), .D(n_11988), .SD(n_61013), .Q(\tab23[28] 
		));
	notech_mux2 i_17718(.S(n_54581), .A(\tab23[28] ), .B(n_52545), .Z(n_11988
		));
	notech_ao4 i_699(.A(n_1098), .B(n_13635), .C(n_486), .D(n_13728), .Z(n_1282
		));
	notech_reg_set tab23_reg_29(.CP(n_61708), .D(n_11994), .SD(n_61011), .Q(\tab23[29] 
		));
	notech_mux2 i_17726(.S(n_54581), .A(\tab23[29] ), .B(n_52551), .Z(n_11994
		));
	notech_ao4 i_698(.A(n_53455), .B(n_13634), .C(n_486), .D(n_13727), .Z(n_1283
		));
	notech_reg tab23_reg_30(.CP(n_61708), .D(n_12000), .CD(n_61011), .Q(\tab23[30] 
		));
	notech_mux2 i_17734(.S(n_54581), .A(\tab23[30] ), .B(n_974), .Z(n_12000)
		);
	notech_ao4 i_697(.A(n_53455), .B(n_13633), .C(n_486), .D(n_13726), .Z(n_1284
		));
	notech_reg tab23_reg_32(.CP(n_61710), .D(n_12006), .CD(n_61013), .Q(\tab23[32] 
		));
	notech_mux2 i_17742(.S(n_54581), .A(\tab23[32] ), .B(n_975), .Z(n_12006)
		);
	notech_ao4 i_696(.A(n_53455), .B(n_13632), .C(n_486), .D(n_13725), .Z(n_1285
		));
	notech_reg_set tab23_reg_33(.CP(n_61710), .D(n_12012), .SD(n_61013), .Q(\tab23[33] 
		));
	notech_mux2 i_17750(.S(n_54581), .A(\tab23[33] ), .B(n_54613), .Z(n_12012
		));
	notech_ao4 i_695(.A(n_53455), .B(n_13631), .C(n_486), .D(n_13724), .Z(n_1286
		));
	notech_reg hit_adr23_reg(.CP(n_61711), .D(n_12018), .CD(n_61014), .Q(hit_adr23
		));
	notech_mux2 i_17758(.S(n_971), .A(hit_add23), .B(hit_adr23), .Z(n_12018)
		);
	notech_ao4 i_694(.A(n_53455), .B(n_13630), .C(n_486), .D(n_13723), .Z(n_1287
		));
	notech_reg_set tab24_reg_0(.CP(n_61711), .D(n_12024), .SD(n_61014), .Q(\tab24[0] 
		));
	notech_mux2 i_17766(.S(\nbus_14028[0] ), .A(\tab24[0] ), .B(n_52377), .Z
		(n_12024));
	notech_reg_set tab24_reg_1(.CP(n_61711), .D(n_12030), .SD(n_61014), .Q(\tab24[1] 
		));
	notech_mux2 i_17774(.S(\nbus_14028[0] ), .A(\tab24[1] ), .B(n_52383), .Z
		(n_12030));
	notech_ao4 i_76262(.A(n_61604), .B(n_13784), .C(n_986), .D(n_987), .Z(oread_ack97032
		));
	notech_reg_set tab24_reg_2(.CP(n_61711), .D(n_12036), .SD(n_61014), .Q(\tab24[2] 
		));
	notech_mux2 i_17782(.S(\nbus_14028[0] ), .A(\tab24[2] ), .B(n_52389), .Z
		(n_12036));
	notech_nao3 i_78751(.A(n_631), .B(n_625), .C(n_628), .Z(\nbus_14042[0] )
		);
	notech_reg_set tab24_reg_3(.CP(n_61711), .D(n_12042), .SD(n_61014), .Q(\tab24[3] 
		));
	notech_mux2 i_17790(.S(\nbus_14028[0] ), .A(\tab24[3] ), .B(n_52395), .Z
		(n_12042));
	notech_nand2 i_78860(.A(n_625), .B(n_994), .Z(\nbus_14043[0] ));
	notech_reg tab24_reg_4(.CP(n_61710), .D(n_12048), .CD(n_61013), .Q(\tab24[4] 
		));
	notech_mux2 i_17798(.S(\nbus_14028[0] ), .A(\tab24[4] ), .B(n_973), .Z(n_12048
		));
	notech_nand2 i_78386(.A(n_604), .B(n_994), .Z(\nbus_14036[0] ));
	notech_reg_set tab24_reg_5(.CP(n_61710), .D(n_12054), .SD(n_61013), .Q(\tab24[5] 
		));
	notech_mux2 i_17806(.S(\nbus_14028[0] ), .A(\tab24[5] ), .B(n_52407), .Z
		(n_12054));
	notech_nao3 i_78274(.A(n_631), .B(n_601), .C(n_628), .Z(\nbus_14035[0] )
		);
	notech_reg_set tab24_reg_6(.CP(n_61710), .D(n_12060), .SD(n_61013), .Q(\tab24[6] 
		));
	notech_mux2 i_17814(.S(\nbus_14028[0] ), .A(\tab24[6] ), .B(n_52413), .Z
		(n_12060));
	notech_nao3 i_77064(.A(n_631), .B(n_600), .C(n_628), .Z(\nbus_14015[0] )
		);
	notech_reg_set tab24_reg_7(.CP(n_61710), .D(n_12066), .SD(n_61013), .Q(\tab24[7] 
		));
	notech_mux2 i_17822(.S(\nbus_14028[0] ), .A(\tab24[7] ), .B(n_52419), .Z
		(n_12066));
	notech_nao3 i_77176(.A(n_631), .B(n_599), .C(n_628), .Z(\nbus_14016[0] )
		);
	notech_reg_set tab24_reg_8(.CP(n_61707), .D(n_12072), .SD(n_61010), .Q(\tab24[8] 
		));
	notech_mux2 i_17830(.S(\nbus_14028[0] ), .A(\tab24[8] ), .B(n_52425), .Z
		(n_12072));
	notech_nand2 i_78728(.A(n_1020), .B(n_1011), .Z(\nbus_14041[0] ));
	notech_reg_set tab24_reg_9(.CP(n_61707), .D(n_12078), .SD(n_61010), .Q(\tab24[9] 
		));
	notech_mux2 i_17838(.S(\nbus_14028[0] ), .A(\tab24[9] ), .B(n_52431), .Z
		(n_12078));
	notech_ao4 i_78006(.A(n_1001), .B(n_1010), .C(n_1020), .D(n_13499), .Z(\nbus_14031[0] 
		));
	notech_reg_set tab24_reg_10(.CP(n_61707), .D(n_12084), .SD(n_61010), .Q(\tab24[10] 
		));
	notech_mux2 i_17846(.S(\nbus_14028[0] ), .A(\tab24[10] ), .B(n_52437), .Z
		(n_12084));
	notech_nand2 i_78498(.A(n_994), .B(n_579), .Z(\nbus_14037[0] ));
	notech_reg_set tab24_reg_11(.CP(n_61707), .D(n_12090), .SD(n_61010), .Q(\tab24[11] 
		));
	notech_mux2 i_17854(.S(\nbus_14028[0] ), .A(\tab24[11] ), .B(n_52443), .Z
		(n_12090));
	notech_nand2 i_77288(.A(n_994), .B(n_578), .Z(\nbus_14017[0] ));
	notech_reg_set tab24_reg_12(.CP(n_61707), .D(n_12096), .SD(n_61010), .Q(\tab24[12] 
		));
	notech_mux2 i_17862(.S(\nbus_14028[0] ), .A(\tab24[12] ), .B(n_52449), .Z
		(n_12096));
	notech_nand2 i_77719(.A(n_994), .B(n_577), .Z(\nbus_14028[0] ));
	notech_reg_set tab24_reg_13(.CP(n_61707), .D(n_12102), .SD(n_61010), .Q(\tab24[13] 
		));
	notech_mux2 i_17870(.S(\nbus_14028[0] ), .A(\tab24[13] ), .B(n_52455), .Z
		(n_12102));
	notech_ao4 i_77982(.A(n_1002), .B(n_1001), .C(n_1020), .D(n_13490), .Z(\nbus_14030[0] 
		));
	notech_reg_set tab24_reg_14(.CP(n_61707), .D(n_12108), .SD(n_61010), .Q(\tab24[14] 
		));
	notech_mux2 i_17878(.S(\nbus_14028[0] ), .A(\tab24[14] ), .B(n_52461), .Z
		(n_12108));
	notech_nand2 i_78711(.A(n_1020), .B(n_1003), .Z(\nbus_14040[0] ));
	notech_reg_set tab24_reg_15(.CP(n_61707), .D(n_12114), .SD(n_61010), .Q(\tab24[15] 
		));
	notech_mux2 i_17886(.S(\nbus_14028[0] ), .A(\tab24[15] ), .B(n_52467), .Z
		(n_12114));
	notech_nao3 i_78162(.A(n_631), .B(n_557), .C(n_628), .Z(\nbus_14034[0] )
		);
	notech_reg_set tab24_reg_16(.CP(n_61707), .D(n_12120), .SD(n_61010), .Q(\tab24[16] 
		));
	notech_mux2 i_17894(.S(\nbus_14028[0] ), .A(\tab24[16] ), .B(n_52473), .Z
		(n_12120));
	notech_nand2 i_77499(.A(n_992), .B(n_552), .Z(\nbus_14018[0] ));
	notech_reg_set tab24_reg_17(.CP(n_61708), .D(n_12126), .SD(n_61011), .Q(\tab24[17] 
		));
	notech_mux2 i_17902(.S(n_54599), .A(\tab24[17] ), .B(n_52479), .Z(n_12126
		));
	notech_or2 i_85(.A(n_473), .B(n_13484), .Z(n_53238));
	notech_reg_set tab24_reg_18(.CP(n_61708), .D(n_12132), .SD(n_61011), .Q(\tab24[18] 
		));
	notech_mux2 i_17910(.S(n_54599), .A(\tab24[18] ), .B(n_52485), .Z(n_12132
		));
	notech_or4 i_78035(.A(n_473), .B(\nbus_14033[0] ), .C(n_1048), .D(n_13484
		), .Z(\nbus_14032[0] ));
	notech_reg_set tab24_reg_19(.CP(n_61708), .D(n_12138), .SD(n_61011), .Q(\tab24[19] 
		));
	notech_mux2 i_17918(.S(n_54599), .A(\tab24[19] ), .B(n_52491), .Z(n_12138
		));
	notech_nand2 i_87(.A(n_1020), .B(n_545), .Z(\nbus_14033[0] ));
	notech_reg_set tab24_reg_20(.CP(n_61708), .D(n_12144), .SD(n_61011), .Q(\tab24[20] 
		));
	notech_mux2 i_17926(.S(n_54599), .A(\tab24[20] ), .B(n_52497), .Z(n_12144
		));
	notech_reg_set tab24_reg_21(.CP(n_61708), .D(n_12150), .SD(n_61011), .Q(\tab24[21] 
		));
	notech_mux2 i_17934(.S(n_54599), .A(\tab24[21] ), .B(n_52503), .Z(n_12150
		));
	notech_ao4 i_86(.A(n_1001), .B(n_550), .C(data_miss[5]), .D(n_977), .Z(\nbus_14013[0] 
		));
	notech_reg_set tab24_reg_22(.CP(n_61708), .D(n_12156), .SD(n_61011), .Q(\tab24[22] 
		));
	notech_mux2 i_17942(.S(n_54599), .A(\tab24[22] ), .B(n_52509), .Z(n_12156
		));
	notech_or2 i_77832(.A(n_473), .B(n_474), .Z(n_53749));
	notech_reg_set tab24_reg_23(.CP(n_61708), .D(n_12162), .SD(n_61011), .Q(\tab24[23] 
		));
	notech_mux2 i_17950(.S(n_54599), .A(\tab24[23] ), .B(n_52515), .Z(n_12162
		));
	notech_ao4 i_68(.A(data_miss[0]), .B(n_989), .C(n_996), .D(n_13462), .Z(n_53241
		));
	notech_reg_set tab24_reg_24(.CP(n_61708), .D(n_12168), .SD(n_61011), .Q(\tab24[24] 
		));
	notech_mux2 i_17958(.S(n_54599), .A(\tab24[24] ), .B(n_52521), .Z(n_12168
		));
	notech_mux2 i_122741(.S(n_948), .A(iDaddr[12]), .B(iDaddr_f[12]), .Z(\tab11_0[0] 
		));
	notech_reg_set tab24_reg_25(.CP(n_61708), .D(n_12174), .SD(n_61011), .Q(\tab24[25] 
		));
	notech_mux2 i_17966(.S(n_54599), .A(\tab24[25] ), .B(n_52527), .Z(n_12174
		));
	notech_mux2 i_222742(.S(n_948), .A(iDaddr[13]), .B(iDaddr_f[13]), .Z(\tab11_0[1] 
		));
	notech_reg_set tab24_reg_26(.CP(n_61711), .D(n_12180), .SD(n_61014), .Q(\tab24[26] 
		));
	notech_mux2 i_17974(.S(n_54599), .A(\tab24[26] ), .B(n_52533), .Z(n_12180
		));
	notech_mux2 i_322743(.S(n_948), .A(iDaddr[14]), .B(iDaddr_f[14]), .Z(\tab11_0[2] 
		));
	notech_reg_set tab24_reg_27(.CP(n_61715), .D(n_12186), .SD(n_61018), .Q(\tab24[27] 
		));
	notech_mux2 i_17982(.S(\nbus_14028[0] ), .A(\tab24[27] ), .B(n_52539), .Z
		(n_12186));
	notech_mux2 i_422744(.S(n_948), .A(iDaddr[15]), .B(iDaddr_f[15]), .Z(\tab11_0[3] 
		));
	notech_reg_set tab24_reg_28(.CP(n_61715), .D(n_12192), .SD(n_61018), .Q(\tab24[28] 
		));
	notech_mux2 i_17990(.S(n_54599), .A(\tab24[28] ), .B(n_52545), .Z(n_12192
		));
	notech_mux2 i_522745(.S(n_948), .A(iDaddr[16]), .B(iDaddr_f[16]), .Z(\tab11_0[4] 
		));
	notech_reg_set tab24_reg_29(.CP(n_61715), .D(n_12198), .SD(n_61018), .Q(\tab24[29] 
		));
	notech_mux2 i_17998(.S(n_54599), .A(\tab24[29] ), .B(n_52551), .Z(n_12198
		));
	notech_mux2 i_622746(.S(n_58627), .A(iDaddr[17]), .B(iDaddr_f[17]), .Z(\tab11_0[5] 
		));
	notech_reg tab24_reg_30(.CP(n_61715), .D(n_12204), .CD(n_61018), .Q(\tab24[30] 
		));
	notech_mux2 i_18006(.S(n_54599), .A(\tab24[30] ), .B(n_974), .Z(n_12204)
		);
	notech_mux2 i_722747(.S(n_58627), .A(iDaddr[18]), .B(iDaddr_f[18]), .Z(\tab11_0[6] 
		));
	notech_reg tab24_reg_32(.CP(n_61715), .D(n_12210), .CD(n_61018), .Q(\tab24[32] 
		));
	notech_mux2 i_18014(.S(n_54599), .A(\tab24[32] ), .B(n_975), .Z(n_12210)
		);
	notech_mux2 i_822748(.S(n_58627), .A(iDaddr[19]), .B(iDaddr_f[19]), .Z(\tab11_0[7] 
		));
	notech_reg_set tab24_reg_33(.CP(n_61715), .D(n_12216), .SD(n_61018), .Q(\tab24[33] 
		));
	notech_mux2 i_18022(.S(n_54599), .A(\tab24[33] ), .B(n_54613), .Z(n_12216
		));
	notech_mux2 i_922749(.S(n_58627), .A(iDaddr[20]), .B(iDaddr_f[20]), .Z(\tab11_0[8] 
		));
	notech_reg hit_adr24_reg(.CP(n_61715), .D(n_12222), .CD(n_61018), .Q(hit_adr24
		));
	notech_mux2 i_18030(.S(n_971), .A(hit_add24), .B(hit_adr24), .Z(n_12222)
		);
	notech_mux2 i_1022750(.S(n_58627), .A(iDaddr[21]), .B(iDaddr_f[21]), .Z(\tab11_0[9] 
		));
	notech_reg_set nnx_tab2_reg_0(.CP(n_61715), .D(n_12228), .SD(n_61018), .Q
		(\nnx_tab2[0] ));
	notech_mux2 i_18038(.S(n_13609), .A(\nnx_tab2[0] ), .B(n_13605), .Z(n_12228
		));
	notech_mux2 i_1122751(.S(n_58627), .A(iDaddr[22]), .B(iDaddr_f[22]), .Z(\dir1_0[0] 
		));
	notech_reg nnx_tab2_reg_1(.CP(n_61715), .D(n_12234), .CD(n_61018), .Q(\nnx_tab2[1] 
		));
	notech_mux2 i_18046(.S(n_13609), .A(\nnx_tab2[1] ), .B(n_13607), .Z(n_12234
		));
	notech_mux2 i_1222752(.S(n_58627), .A(iDaddr[23]), .B(iDaddr_f[23]), .Z(\dir1_0[1] 
		));
	notech_reg nx_tab2_reg_0(.CP(n_61716), .D(n_12240), .CD(n_61019), .Q(\nx_tab2[0] 
		));
	notech_mux2 i_18054(.S(\nbus_14040[0] ), .A(\nx_tab2[0] ), .B(n_13610), 
		.Z(n_12240));
	notech_mux2 i_1322753(.S(n_58627), .A(iDaddr[24]), .B(iDaddr_f[24]), .Z(\dir1_0[2] 
		));
	notech_reg nx_tab2_reg_1(.CP(n_61716), .D(n_12246), .CD(n_61019), .Q(\nx_tab2[1] 
		));
	notech_mux2 i_18062(.S(\nbus_14040[0] ), .A(\nx_tab2[1] ), .B(n_13612), 
		.Z(n_12246));
	notech_mux2 i_1422754(.S(n_58627), .A(iDaddr[25]), .B(iDaddr_f[25]), .Z(\dir1_0[3] 
		));
	notech_reg_set tab11_reg_0(.CP(n_61716), .D(n_12252), .SD(n_61019), .Q(\tab11[0] 
		));
	notech_mux2 i_18070(.S(\nbus_14034[0] ), .A(\tab11[0] ), .B(n_52377), .Z
		(n_12252));
	notech_mux2 i_1522755(.S(n_58627), .A(iDaddr[26]), .B(iDaddr_f[26]), .Z(\dir1_0[4] 
		));
	notech_reg_set tab11_reg_1(.CP(n_61716), .D(n_12258), .SD(n_61019), .Q(\tab11[1] 
		));
	notech_mux2 i_18078(.S(\nbus_14034[0] ), .A(\tab11[1] ), .B(n_52383), .Z
		(n_12258));
	notech_mux2 i_1622756(.S(n_58627), .A(iDaddr[27]), .B(iDaddr_f[27]), .Z(\dir1_0[5] 
		));
	notech_reg_set tab11_reg_2(.CP(n_61716), .D(n_12264), .SD(n_61019), .Q(\tab11[2] 
		));
	notech_mux2 i_18086(.S(\nbus_14034[0] ), .A(\tab11[2] ), .B(n_52389), .Z
		(n_12264));
	notech_mux2 i_1722757(.S(n_948), .A(iDaddr[28]), .B(iDaddr_f[28]), .Z(\dir1_0[6] 
		));
	notech_reg_set tab11_reg_3(.CP(n_61716), .D(n_12270), .SD(n_61019), .Q(\tab11[3] 
		));
	notech_mux2 i_18094(.S(\nbus_14034[0] ), .A(\tab11[3] ), .B(n_52395), .Z
		(n_12270));
	notech_mux2 i_1822758(.S(n_58627), .A(iDaddr[29]), .B(iDaddr_f[29]), .Z(\dir1_0[7] 
		));
	notech_reg tab11_reg_4(.CP(n_61716), .D(n_12276), .CD(n_61019), .Q(\tab11[4] 
		));
	notech_mux2 i_18102(.S(\nbus_14034[0] ), .A(\tab11[4] ), .B(n_973), .Z(n_12276
		));
	notech_mux2 i_1922759(.S(n_58627), .A(iDaddr[30]), .B(iDaddr_f[30]), .Z(\dir1_0[8] 
		));
	notech_reg_set tab11_reg_5(.CP(n_61716), .D(n_12282), .SD(n_61019), .Q(\tab11[5] 
		));
	notech_mux2 i_18110(.S(\nbus_14034[0] ), .A(\tab11[5] ), .B(n_52407), .Z
		(n_12282));
	notech_mux2 i_2022760(.S(n_58627), .A(iDaddr[31]), .B(iDaddr_f[31]), .Z(\dir1_0[9] 
		));
	notech_reg_set tab11_reg_6(.CP(n_61716), .D(n_12288), .SD(n_61019), .Q(\tab11[6] 
		));
	notech_mux2 i_18118(.S(\nbus_14034[0] ), .A(\tab11[6] ), .B(n_52413), .Z
		(n_12288));
	notech_mux2 i_122280(.S(n_53478), .A(wrD[0]), .B(iwrite_data[0]), .Z(n_53009
		));
	notech_reg_set tab11_reg_7(.CP(n_61712), .D(n_12294), .SD(n_61015), .Q(\tab11[7] 
		));
	notech_mux2 i_18126(.S(\nbus_14034[0] ), .A(\tab11[7] ), .B(n_52419), .Z
		(n_12294));
	notech_mux2 i_222281(.S(n_53478), .A(wrD[1]), .B(iwrite_data[1]), .Z(n_53016
		));
	notech_reg_set tab11_reg_8(.CP(n_61712), .D(n_12300), .SD(n_61015), .Q(\tab11[8] 
		));
	notech_mux2 i_18134(.S(\nbus_14034[0] ), .A(\tab11[8] ), .B(n_52425), .Z
		(n_12300));
	notech_mux2 i_322282(.S(n_53478), .A(wrD[2]), .B(iwrite_data[2]), .Z(n_53023
		));
	notech_reg_set tab11_reg_9(.CP(n_61712), .D(n_12306), .SD(n_61015), .Q(\tab11[9] 
		));
	notech_mux2 i_18142(.S(\nbus_14034[0] ), .A(\tab11[9] ), .B(n_52431), .Z
		(n_12306));
	notech_mux2 i_422283(.S(n_53478), .A(wrD[3]), .B(iwrite_data[3]), .Z(n_53030
		));
	notech_reg_set tab11_reg_10(.CP(n_61712), .D(n_12312), .SD(n_61015), .Q(\tab11[10] 
		));
	notech_mux2 i_18150(.S(\nbus_14034[0] ), .A(\tab11[10] ), .B(n_52437), .Z
		(n_12312));
	notech_mux2 i_522284(.S(n_53478), .A(wrD[4]), .B(iwrite_data[4]), .Z(n_53037
		));
	notech_reg_set tab11_reg_11(.CP(n_61711), .D(n_12318), .SD(n_61014), .Q(\tab11[11] 
		));
	notech_mux2 i_18158(.S(\nbus_14034[0] ), .A(\tab11[11] ), .B(n_52443), .Z
		(n_12318));
	notech_mux2 i_622285(.S(n_53478), .A(wrD[5]), .B(iwrite_data[5]), .Z(n_53044
		));
	notech_reg_set tab11_reg_12(.CP(n_61711), .D(n_12324), .SD(n_61014), .Q(\tab11[12] 
		));
	notech_mux2 i_18166(.S(\nbus_14034[0] ), .A(\tab11[12] ), .B(n_52449), .Z
		(n_12324));
	notech_mux2 i_722286(.S(n_53478), .A(wrD[6]), .B(iwrite_data[6]), .Z(n_53051
		));
	notech_reg_set tab11_reg_13(.CP(n_61711), .D(n_12330), .SD(n_61014), .Q(\tab11[13] 
		));
	notech_mux2 i_18174(.S(\nbus_14034[0] ), .A(\tab11[13] ), .B(n_52455), .Z
		(n_12330));
	notech_mux2 i_822287(.S(n_53478), .A(wrD[7]), .B(iwrite_data[7]), .Z(n_53058
		));
	notech_reg_set tab11_reg_14(.CP(n_61711), .D(n_12336), .SD(n_61014), .Q(\tab11[14] 
		));
	notech_mux2 i_18182(.S(\nbus_14034[0] ), .A(\tab11[14] ), .B(n_52461), .Z
		(n_12336));
	notech_mux2 i_922288(.S(n_53478), .A(wrD[8]), .B(iwrite_data[8]), .Z(n_53065
		));
	notech_reg_set tab11_reg_15(.CP(n_61711), .D(n_12342), .SD(n_61014), .Q(\tab11[15] 
		));
	notech_mux2 i_18190(.S(\nbus_14034[0] ), .A(\tab11[15] ), .B(n_52467), .Z
		(n_12342));
	notech_mux2 i_1022289(.S(n_53478), .A(wrD[9]), .B(iwrite_data[9]), .Z(n_53072
		));
	notech_reg_set tab11_reg_16(.CP(n_61712), .D(n_12348), .SD(n_61015), .Q(\tab11[16] 
		));
	notech_mux2 i_18198(.S(\nbus_14034[0] ), .A(\tab11[16] ), .B(n_52473), .Z
		(n_12348));
	notech_mux2 i_1122290(.S(n_53478), .A(wrD[10]), .B(iwrite_data[10]), .Z(n_53079
		));
	notech_reg_set tab11_reg_17(.CP(n_61712), .D(n_12354), .SD(n_61015), .Q(\tab11[17] 
		));
	notech_mux2 i_18206(.S(n_54552), .A(\tab11[17] ), .B(n_52479), .Z(n_12354
		));
	notech_mux2 i_1222291(.S(n_53478), .A(wrD[11]), .B(iwrite_data[11]), .Z(n_53086
		));
	notech_reg_set tab11_reg_18(.CP(n_61715), .D(n_12360), .SD(n_61018), .Q(\tab11[18] 
		));
	notech_mux2 i_18214(.S(n_54552), .A(\tab11[18] ), .B(n_52485), .Z(n_12360
		));
	notech_mux2 i_1322292(.S(n_53478), .A(wrD[12]), .B(iwrite_data[12]), .Z(n_53093
		));
	notech_reg_set tab11_reg_19(.CP(n_61715), .D(n_12366), .SD(n_61018), .Q(\tab11[19] 
		));
	notech_mux2 i_18222(.S(n_54552), .A(\tab11[19] ), .B(n_52491), .Z(n_12366
		));
	notech_mux2 i_1422293(.S(n_53478), .A(wrD[13]), .B(iwrite_data[13]), .Z(n_53100
		));
	notech_reg_set tab11_reg_20(.CP(n_61712), .D(n_12372), .SD(n_61015), .Q(\tab11[20] 
		));
	notech_mux2 i_18230(.S(n_54552), .A(\tab11[20] ), .B(n_52497), .Z(n_12372
		));
	notech_mux2 i_1522294(.S(n_53478), .A(wrD[14]), .B(iwrite_data[14]), .Z(n_53107
		));
	notech_reg_set tab11_reg_21(.CP(n_61712), .D(n_12378), .SD(n_61015), .Q(\tab11[21] 
		));
	notech_mux2 i_18238(.S(n_54552), .A(\tab11[21] ), .B(n_52503), .Z(n_12378
		));
	notech_mux2 i_1622295(.S(n_53473), .A(wrD[15]), .B(iwrite_data[15]), .Z(n_53114
		));
	notech_reg_set tab11_reg_22(.CP(n_61712), .D(n_12384), .SD(n_61015), .Q(\tab11[22] 
		));
	notech_mux2 i_18246(.S(n_54552), .A(\tab11[22] ), .B(n_52509), .Z(n_12384
		));
	notech_mux2 i_1722296(.S(n_53473), .A(wrD[16]), .B(iwrite_data[16]), .Z(n_53121
		));
	notech_reg_set tab11_reg_23(.CP(n_61712), .D(n_12390), .SD(n_61015), .Q(\tab11[23] 
		));
	notech_mux2 i_18254(.S(n_54552), .A(\tab11[23] ), .B(n_52515), .Z(n_12390
		));
	notech_mux2 i_1822297(.S(n_53473), .A(wrD[17]), .B(iwrite_data[17]), .Z(n_53128
		));
	notech_reg_set tab11_reg_24(.CP(n_61712), .D(n_12396), .SD(n_61015), .Q(\tab11[24] 
		));
	notech_mux2 i_18262(.S(n_54552), .A(\tab11[24] ), .B(n_52521), .Z(n_12396
		));
	notech_mux2 i_1922298(.S(n_53473), .A(wrD[18]), .B(iwrite_data[18]), .Z(n_53135
		));
	notech_reg_set tab11_reg_25(.CP(n_61707), .D(n_12402), .SD(n_61010), .Q(\tab11[25] 
		));
	notech_mux2 i_18270(.S(n_54552), .A(\tab11[25] ), .B(n_52527), .Z(n_12402
		));
	notech_mux2 i_2022299(.S(n_53473), .A(wrD[19]), .B(iwrite_data[19]), .Z(n_53142
		));
	notech_reg_set tab11_reg_26(.CP(n_61698), .D(n_12408), .SD(n_61001), .Q(\tab11[26] 
		));
	notech_mux2 i_18278(.S(n_54552), .A(\tab11[26] ), .B(n_52533), .Z(n_12408
		));
	notech_mux2 i_2122300(.S(n_53473), .A(wrD[20]), .B(iwrite_data[20]), .Z(n_53149
		));
	notech_reg_set tab11_reg_27(.CP(n_61698), .D(n_12414), .SD(n_61001), .Q(\tab11[27] 
		));
	notech_mux2 i_18286(.S(\nbus_14034[0] ), .A(\tab11[27] ), .B(n_52539), .Z
		(n_12414));
	notech_mux2 i_2222301(.S(n_53473), .A(wrD[21]), .B(iwrite_data[21]), .Z(n_53156
		));
	notech_reg_set tab11_reg_28(.CP(n_61698), .D(n_12420), .SD(n_61001), .Q(\tab11[28] 
		));
	notech_mux2 i_18294(.S(n_54552), .A(\tab11[28] ), .B(n_52545), .Z(n_12420
		));
	notech_mux2 i_2322302(.S(n_53473), .A(wrD[22]), .B(iwrite_data[22]), .Z(n_53163
		));
	notech_reg_set tab11_reg_29(.CP(n_61698), .D(n_12426), .SD(n_61001), .Q(\tab11[29] 
		));
	notech_mux2 i_18302(.S(n_54552), .A(\tab11[29] ), .B(n_52551), .Z(n_12426
		));
	notech_mux2 i_2422303(.S(n_53473), .A(wrD[23]), .B(iwrite_data[23]), .Z(n_53170
		));
	notech_reg tab11_reg_30(.CP(n_61698), .D(n_12432), .CD(n_61001), .Q(\tab11[30] 
		));
	notech_mux2 i_18310(.S(n_54552), .A(\tab11[30] ), .B(n_974), .Z(n_12432)
		);
	notech_mux2 i_2522304(.S(n_53473), .A(wrD[24]), .B(iwrite_data[24]), .Z(n_53177
		));
	notech_reg tab11_reg_32(.CP(n_61698), .D(n_12438), .CD(n_61001), .Q(\tab11[32] 
		));
	notech_mux2 i_18318(.S(n_54552), .A(\tab11[32] ), .B(n_975), .Z(n_12438)
		);
	notech_mux2 i_2622305(.S(n_53473), .A(wrD[25]), .B(iwrite_data[25]), .Z(n_53184
		));
	notech_reg_set tab11_reg_33(.CP(n_61698), .D(n_12444), .SD(n_61001), .Q(\tab11[33] 
		));
	notech_mux2 i_18326(.S(n_54552), .A(\tab11[33] ), .B(n_54613), .Z(n_12444
		));
	notech_mux2 i_2722306(.S(n_53478), .A(wrD[26]), .B(iwrite_data[26]), .Z(n_53191
		));
	notech_reg fsm5_cnt_reg_0(.CP(n_61698), .D(n_12450), .CD(n_61001), .Q(fsm5_cnt
		[0]));
	notech_mux2 i_18334(.S(\nbus_14018[0] ), .A(fsm5_cnt[0]), .B(n_962), .Z(n_12450
		));
	notech_mux2 i_2822307(.S(n_53473), .A(wrD[27]), .B(iwrite_data[27]), .Z(n_53198
		));
	notech_reg fsm5_cnt_reg_1(.CP(n_61698), .D(n_12456), .CD(n_61001), .Q(fsm5_cnt
		[1]));
	notech_mux2 i_18342(.S(\nbus_14018[0] ), .A(fsm5_cnt[1]), .B(n_963), .Z(n_12456
		));
	notech_mux2 i_2922308(.S(n_53473), .A(wrD[28]), .B(iwrite_data[28]), .Z(n_53205
		));
	notech_reg fsm5_cnt_reg_2(.CP(n_61701), .D(n_12462), .CD(n_61004), .Q(fsm5_cnt
		[2]));
	notech_mux2 i_18350(.S(\nbus_14018[0] ), .A(fsm5_cnt[2]), .B(n_964), .Z(n_12462
		));
	notech_mux2 i_3022309(.S(n_53473), .A(wrD[29]), .B(iwrite_data[29]), .Z(n_53212
		));
	notech_reg fsm5_cnt_reg_3(.CP(n_61701), .D(n_12468), .CD(n_61004), .Q(fsm5_cnt
		[3]));
	notech_mux2 i_18358(.S(\nbus_14018[0] ), .A(fsm5_cnt[3]), .B(n_965), .Z(n_12468
		));
	notech_mux2 i_3122310(.S(n_53473), .A(wrD[30]), .B(iwrite_data[30]), .Z(n_53219
		));
	notech_reg fsm5_cnt_reg_4(.CP(n_61701), .D(n_12474), .CD(n_61004), .Q(fsm5_cnt
		[4]));
	notech_mux2 i_18366(.S(\nbus_14018[0] ), .A(fsm5_cnt[4]), .B(n_966), .Z(n_12474
		));
	notech_mux2 i_3222311(.S(n_53473), .A(wrD[31]), .B(iwrite_data[31]), .Z(n_53226
		));
	notech_reg fsm5_cnt_reg_5(.CP(n_61701), .D(n_12480), .CD(n_61004), .Q(fsm5_cnt
		[5]));
	notech_mux2 i_18374(.S(\nbus_14018[0] ), .A(fsm5_cnt[5]), .B(n_967), .Z(n_12480
		));
	notech_nand2 i_8(.A(n_996), .B(n_989), .Z(n_52185));
	notech_reg fsm5_cnt_reg_6(.CP(n_61701), .D(n_12486), .CD(n_61004), .Q(fsm5_cnt
		[6]));
	notech_mux2 i_18382(.S(\nbus_14018[0] ), .A(fsm5_cnt[6]), .B(n_968), .Z(n_12486
		));
	notech_or2 i_76179(.A(n_974), .B(data_miss[6]), .Z(n_52191));
	notech_reg fsm5_cnt_reg_7(.CP(n_61698), .D(n_12492), .CD(n_61001), .Q(fsm5_cnt
		[7]));
	notech_mux2 i_18390(.S(\nbus_14018[0] ), .A(fsm5_cnt[7]), .B(n_969), .Z(n_12492
		));
	notech_nand2 i_122248(.A(n_1287), .B(n_475), .Z(n_53761));
	notech_reg fsm5_cnt_reg_8(.CP(n_61698), .D(n_12498), .CD(n_61001), .Q(fsm5_cnt
		[8]));
	notech_mux2 i_18398(.S(\nbus_14018[0] ), .A(fsm5_cnt[8]), .B(n_970), .Z(n_12498
		));
	notech_nand2 i_222249(.A(n_1286), .B(n_476), .Z(n_53768));
	notech_reg pg_fault_reg(.CP(n_61701), .D(n_12504), .CD(n_61004), .Q(pg_fault
		));
	notech_mux2 i_18406(.S(n_53238), .A(pg_fault), .B(n_13614), .Z(n_12504)
		);
	notech_nand2 i_322250(.A(n_1285), .B(n_477), .Z(n_53775));
	notech_reg fsm_reg_0(.CP(n_61698), .D(n_12510), .CD(n_61001), .Q(fsm[0])
		);
	notech_mux2 i_18414(.S(\nbus_14032[0] ), .A(n_58636), .B(n_54148), .Z(n_12510
		));
	notech_nand2 i_422251(.A(n_1284), .B(n_478), .Z(n_53782));
	notech_reg fsm_reg_1(.CP(n_61697), .D(n_12516), .CD(n_61000), .Q(fsm[1])
		);
	notech_mux2 i_18422(.S(\nbus_14032[0] ), .A(fsm[1]), .B(n_13615), .Z(n_12516
		));
	notech_nand2 i_522252(.A(n_1283), .B(n_479), .Z(n_53789));
	notech_reg fsm_reg_2(.CP(n_61697), .D(n_12522), .CD(n_61000), .Q(fsm[2])
		);
	notech_mux2 i_18430(.S(\nbus_14032[0] ), .A(fsm[2]), .B(n_54160), .Z(n_12522
		));
	notech_nand2 i_622253(.A(n_1282), .B(n_480), .Z(n_53796));
	notech_reg fsm_reg_3(.CP(n_61697), .D(n_12528), .CD(n_61000), .Q(fsm[3])
		);
	notech_mux2 i_18438(.S(\nbus_14032[0] ), .A(fsm[3]), .B(n_961), .Z(n_12528
		));
	notech_nand2 i_722254(.A(n_1281), .B(n_481), .Z(n_53803));
	notech_reg owrite_req_reg(.CP(n_61697), .D(n_55943), .CD(n_61000), .Q(owrite_req
		));
	notech_reg addr_miss_reg_0(.CP(n_61697), .D(n_12539), .CD(n_61000), .Q(addr_miss
		[0]));
	notech_and3 i_18452(.A(n_1020), .B(n_545), .C(addr_miss[0]), .Z(n_12539)
		);
	notech_nand2 i_822255(.A(n_1280), .B(n_482), .Z(n_53810));
	notech_reg addr_miss_reg_1(.CP(n_61697), .D(n_12545), .CD(n_61000), .Q(addr_miss
		[1]));
	notech_and3 i_18460(.A(n_1020), .B(n_545), .C(addr_miss[1]), .Z(n_12545)
		);
	notech_nand2 i_922256(.A(n_1279), .B(n_483), .Z(n_53817));
	notech_reg addr_miss_reg_2(.CP(n_61697), .D(n_12548), .CD(n_61000), .Q(addr_miss
		[2]));
	notech_mux2 i_18466(.S(\nbus_14033[0] ), .A(addr_miss[2]), .B(n_13619), 
		.Z(n_12548));
	notech_nand2 i_1022257(.A(n_1278), .B(n_484), .Z(n_53824));
	notech_reg addr_miss_reg_3(.CP(n_61697), .D(n_12554), .CD(n_61000), .Q(addr_miss
		[3]));
	notech_mux2 i_18474(.S(\nbus_14033[0] ), .A(addr_miss[3]), .B(n_13620), 
		.Z(n_12554));
	notech_nand2 i_1122258(.A(n_1277), .B(n_485), .Z(n_53831));
	notech_reg addr_miss_reg_4(.CP(n_61697), .D(n_12560), .CD(n_61000), .Q(addr_miss
		[4]));
	notech_mux2 i_18482(.S(\nbus_14033[0] ), .A(addr_miss[4]), .B(n_13621), 
		.Z(n_12560));
	notech_nand2 i_1222259(.A(n_1276), .B(n_487), .Z(n_53838));
	notech_reg addr_miss_reg_5(.CP(n_61698), .D(n_12566), .CD(n_61001), .Q(addr_miss
		[5]));
	notech_mux2 i_18490(.S(\nbus_14033[0] ), .A(addr_miss[5]), .B(n_13622), 
		.Z(n_12566));
	notech_and4 i_1322260(.A(n_1272), .B(n_1274), .C(n_1271), .D(n_686), .Z(n_53845
		));
	notech_reg addr_miss_reg_6(.CP(n_61698), .D(n_12572), .CD(n_61001), .Q(addr_miss
		[6]));
	notech_mux2 i_18498(.S(\nbus_14033[0] ), .A(addr_miss[6]), .B(n_13623), 
		.Z(n_12572));
	notech_and4 i_1422261(.A(n_1263), .B(n_1265), .C(n_1262), .D(n_697), .Z(n_53852
		));
	notech_reg addr_miss_reg_7(.CP(n_61698), .D(n_12578), .CD(n_61001), .Q(addr_miss
		[7]));
	notech_mux2 i_18506(.S(\nbus_14033[0] ), .A(addr_miss[7]), .B(n_13624), 
		.Z(n_12578));
	notech_and4 i_1522262(.A(n_1254), .B(n_1256), .C(n_1253), .D(n_708), .Z(n_53859
		));
	notech_reg addr_miss_reg_8(.CP(n_61698), .D(n_12584), .CD(n_61001), .Q(addr_miss
		[8]));
	notech_mux2 i_18514(.S(\nbus_14033[0] ), .A(addr_miss[8]), .B(n_13625), 
		.Z(n_12584));
	notech_and4 i_1622263(.A(n_1245), .B(n_1247), .C(n_1244), .D(n_719), .Z(n_53866
		));
	notech_reg addr_miss_reg_9(.CP(n_61698), .D(n_12590), .CD(n_61001), .Q(addr_miss
		[9]));
	notech_mux2 i_18522(.S(\nbus_14033[0] ), .A(addr_miss[9]), .B(n_13626), 
		.Z(n_12590));
	notech_and4 i_1722264(.A(n_1236), .B(n_1238), .C(n_1235), .D(n_730), .Z(n_53873
		));
	notech_reg addr_miss_reg_10(.CP(n_61698), .D(n_12596), .CD(n_61001), .Q(addr_miss
		[10]));
	notech_mux2 i_18530(.S(\nbus_14033[0] ), .A(addr_miss[10]), .B(n_13627),
		 .Z(n_12596));
	notech_and4 i_1822265(.A(n_1227), .B(n_1229), .C(n_1226), .D(n_741), .Z(n_53880
		));
	notech_reg addr_miss_reg_11(.CP(n_61697), .D(n_12602), .CD(n_61000), .Q(addr_miss
		[11]));
	notech_mux2 i_18538(.S(\nbus_14033[0] ), .A(addr_miss[11]), .B(n_13628),
		 .Z(n_12602));
	notech_and4 i_1922266(.A(n_1218), .B(n_1220), .C(n_1217), .D(n_752), .Z(n_53887
		));
	notech_reg addr_miss_reg_12(.CP(n_61698), .D(n_12608), .CD(n_61001), .Q(addr_miss
		[12]));
	notech_mux2 i_18546(.S(\nbus_14033[0] ), .A(addr_miss[12]), .B(n_54249),
		 .Z(n_12608));
	notech_and4 i_2022267(.A(n_1209), .B(n_1211), .C(n_1208), .D(n_763), .Z(n_53894
		));
	notech_reg addr_miss_reg_13(.CP(n_61698), .D(n_12614), .CD(n_61001), .Q(addr_miss
		[13]));
	notech_mux2 i_18554(.S(\nbus_14033[0] ), .A(addr_miss[13]), .B(n_54255),
		 .Z(n_12614));
	notech_and4 i_2122268(.A(n_1200), .B(n_1202), .C(n_1199), .D(n_774), .Z(n_53901
		));
	notech_reg addr_miss_reg_14(.CP(n_61701), .D(n_12620), .CD(n_61004), .Q(addr_miss
		[14]));
	notech_mux2 i_18562(.S(\nbus_14033[0] ), .A(addr_miss[14]), .B(n_54261),
		 .Z(n_12620));
	notech_and4 i_2222269(.A(n_1191), .B(n_1193), .C(n_1190), .D(n_785), .Z(n_53908
		));
	notech_reg addr_miss_reg_15(.CP(n_61706), .D(n_12626), .CD(n_61009), .Q(addr_miss
		[15]));
	notech_mux2 i_18570(.S(\nbus_14033[0] ), .A(addr_miss[15]), .B(n_54267),
		 .Z(n_12626));
	notech_and4 i_2322270(.A(n_1182), .B(n_1184), .C(n_1181), .D(n_796), .Z(n_53915
		));
	notech_reg addr_miss_reg_16(.CP(n_61703), .D(n_12632), .CD(n_61006), .Q(addr_miss
		[16]));
	notech_mux2 i_18578(.S(\nbus_14033[0] ), .A(addr_miss[16]), .B(n_54273),
		 .Z(n_12632));
	notech_and4 i_2422271(.A(n_1173), .B(n_1175), .C(n_1172), .D(n_807), .Z(n_53922
		));
	notech_reg addr_miss_reg_17(.CP(n_61706), .D(n_12638), .CD(n_61009), .Q(addr_miss
		[17]));
	notech_mux2 i_18586(.S(n_54825), .A(addr_miss[17]), .B(n_54279), .Z(n_12638
		));
	notech_and4 i_2522272(.A(n_1164), .B(n_1166), .C(n_1163), .D(n_818), .Z(n_53929
		));
	notech_reg addr_miss_reg_18(.CP(n_61706), .D(n_12644), .CD(n_61009), .Q(addr_miss
		[18]));
	notech_mux2 i_18594(.S(n_54825), .A(addr_miss[18]), .B(n_54285), .Z(n_12644
		));
	notech_and4 i_2622273(.A(n_1155), .B(n_1157), .C(n_1154), .D(n_829), .Z(n_53936
		));
	notech_reg addr_miss_reg_19(.CP(n_61703), .D(n_12650), .CD(n_61006), .Q(addr_miss
		[19]));
	notech_mux2 i_18602(.S(n_54825), .A(addr_miss[19]), .B(n_54291), .Z(n_12650
		));
	notech_and4 i_2722274(.A(n_1146), .B(n_1148), .C(n_1145), .D(n_840), .Z(n_53943
		));
	notech_reg addr_miss_reg_20(.CP(n_61703), .D(n_12656), .CD(n_61006), .Q(addr_miss
		[20]));
	notech_mux2 i_18610(.S(n_54825), .A(addr_miss[20]), .B(n_54297), .Z(n_12656
		));
	notech_and4 i_2822275(.A(n_1137), .B(n_1139), .C(n_1136), .D(n_851), .Z(n_53950
		));
	notech_reg addr_miss_reg_21(.CP(n_61703), .D(n_12662), .CD(n_61006), .Q(addr_miss
		[21]));
	notech_mux2 i_18618(.S(n_54825), .A(addr_miss[21]), .B(n_54303), .Z(n_12662
		));
	notech_and4 i_2922276(.A(n_1128), .B(n_1130), .C(n_1127), .D(n_862), .Z(n_53957
		));
	notech_reg addr_miss_reg_22(.CP(n_61703), .D(n_12668), .CD(n_61006), .Q(addr_miss
		[22]));
	notech_mux2 i_18626(.S(n_54825), .A(addr_miss[22]), .B(n_54309), .Z(n_12668
		));
	notech_and4 i_3022277(.A(n_1119), .B(n_1121), .C(n_1118), .D(n_873), .Z(n_53964
		));
	notech_reg addr_miss_reg_23(.CP(n_61703), .D(n_12674), .CD(n_61006), .Q(addr_miss
		[23]));
	notech_mux2 i_18634(.S(n_54825), .A(addr_miss[23]), .B(n_54315), .Z(n_12674
		));
	notech_and4 i_3122278(.A(n_1110), .B(n_1112), .C(n_1109), .D(n_884), .Z(n_53971
		));
	notech_reg addr_miss_reg_24(.CP(n_61706), .D(n_12680), .CD(n_61009), .Q(addr_miss
		[24]));
	notech_mux2 i_18642(.S(n_54825), .A(addr_miss[24]), .B(n_54321), .Z(n_12680
		));
	notech_and4 i_3222279(.A(n_1101), .B(n_1103), .C(n_1095), .D(n_895), .Z(n_53978
		));
	notech_reg addr_miss_reg_25(.CP(n_61706), .D(n_12686), .CD(n_61009), .Q(addr_miss
		[25]));
	notech_mux2 i_18650(.S(n_54825), .A(addr_miss[25]), .B(n_54327), .Z(n_12686
		));
	notech_nand3 i_76120(.A(n_905), .B(n_904), .C(n_491), .Z(n_54124));
	notech_reg addr_miss_reg_26(.CP(n_61707), .D(n_12692), .CD(n_61010), .Q(addr_miss
		[26]));
	notech_mux2 i_18658(.S(n_54825), .A(addr_miss[26]), .B(n_54333), .Z(n_12692
		));
	notech_reg addr_miss_reg_27(.CP(n_61706), .D(n_12698), .CD(n_61009), .Q(addr_miss
		[27]));
	notech_mux2 i_18666(.S(n_54825), .A(addr_miss[27]), .B(n_54339), .Z(n_12698
		));
	notech_ao4 i_76027(.A(n_54796), .B(n_13767), .C(n_13777), .D(n_1016), .Z
		(n_54189));
	notech_reg addr_miss_reg_28(.CP(n_61706), .D(n_12704), .CD(n_61009), .Q(addr_miss
		[28]));
	notech_mux2 i_18674(.S(n_54825), .A(addr_miss[28]), .B(n_54345), .Z(n_12704
		));
	notech_ao4 i_76030(.A(n_54796), .B(n_13766), .C(n_1016), .D(n_13776), .Z
		(n_54195));
	notech_reg addr_miss_reg_29(.CP(n_61706), .D(n_12710), .CD(n_61009), .Q(addr_miss
		[29]));
	notech_mux2 i_18682(.S(n_54825), .A(addr_miss[29]), .B(n_54351), .Z(n_12710
		));
	notech_ao4 i_76033(.A(n_54796), .B(n_13765), .C(n_1016), .D(n_13775), .Z
		(n_54201));
	notech_reg addr_miss_reg_30(.CP(n_61706), .D(n_12716), .CD(n_61009), .Q(addr_miss
		[30]));
	notech_mux2 i_18690(.S(n_54825), .A(addr_miss[30]), .B(n_54357), .Z(n_12716
		));
	notech_ao4 i_76036(.A(n_54796), .B(n_13764), .C(n_1016), .D(n_13774), .Z
		(n_54207));
	notech_reg addr_miss_reg_31(.CP(n_61706), .D(n_12722), .CD(n_61009), .Q(addr_miss
		[31]));
	notech_mux2 i_18698(.S(n_54825), .A(addr_miss[31]), .B(n_54363), .Z(n_12722
		));
	notech_ao4 i_76039(.A(n_54796), .B(n_13763), .C(n_1016), .D(n_13773), .Z
		(n_54213));
	notech_reg req_miss_reg(.CP(n_61706), .D(n_12728), .CD(n_61009), .Q(req_miss
		));
	notech_or2 i_18706(.A(n_12730), .B(n_12731), .Z(n_12728));
	notech_ao4 i_18707(.A(n_54807), .B(n_13458), .C(n_54825), .D(n_13484), .Z
		(n_12730));
	notech_and4 i_18708(.A(req_miss), .B(n_1020), .C(n_545), .D(n_494), .Z(n_12731
		));
	notech_ao4 i_76042(.A(n_54796), .B(n_13762), .C(n_1016), .D(n_13772), .Z
		(n_54219));
	notech_reg oread_req_reg(.CP(n_61701), .D(n_54124), .CD(n_61004), .Q(oread_req
		));
	notech_reg owrite_sz_reg_0(.CP(n_61701), .D(n_902), .CD(n_61004), .Q(owrite_sz
		[0]));
	notech_reg owrite_sz_reg_1(.CP(n_61701), .D(n_903), .CD(n_61004), .Q(owrite_sz
		[1]));
	notech_reg wrA_reg_0(.CP(n_61701), .D(n_12740), .CD(n_61004), .Q(wrA[0])
		);
	notech_mux2 i_18726(.S(n_53367), .A(wrA[0]), .B(addr_miss[0]), .Z(n_12740
		));
	notech_ao4 i_76045(.A(n_54796), .B(n_13761), .C(n_1016), .D(n_13771), .Z
		(n_54225));
	notech_reg wrA_reg_1(.CP(n_61701), .D(n_12746), .CD(n_61004), .Q(wrA[1])
		);
	notech_mux2 i_18734(.S(n_53367), .A(wrA[1]), .B(addr_miss[1]), .Z(n_12746
		));
	notech_ao4 i_76048(.A(n_54796), .B(n_13760), .C(n_1016), .D(n_13770), .Z
		(n_54231));
	notech_reg wrA_reg_2(.CP(n_61701), .D(n_12752), .CD(n_61004), .Q(wrA[2])
		);
	notech_mux2 i_18742(.S(n_53367), .A(wrA[2]), .B(addr_miss[2]), .Z(n_12752
		));
	notech_ao4 i_76051(.A(n_54796), .B(n_13759), .C(n_1016), .D(n_13769), .Z
		(n_54237));
	notech_reg wrA_reg_3(.CP(n_61701), .D(n_12758), .CD(n_61004), .Q(wrA[3])
		);
	notech_mux2 i_18750(.S(n_53367), .A(wrA[3]), .B(addr_miss[3]), .Z(n_12758
		));
	notech_ao4 i_76054(.A(n_54796), .B(n_13758), .C(n_1016), .D(n_13768), .Z
		(n_54243));
	notech_reg wrA_reg_4(.CP(n_61701), .D(n_12764), .CD(n_61004), .Q(wrA[4])
		);
	notech_mux2 i_18758(.S(n_53367), .A(wrA[4]), .B(addr_miss[4]), .Z(n_12764
		));
	notech_nand2 i_76057(.A(n_1076), .B(n_515), .Z(n_54249));
	notech_reg wrA_reg_5(.CP(n_61701), .D(n_12770), .CD(n_61004), .Q(wrA[5])
		);
	notech_mux2 i_18766(.S(n_53367), .A(wrA[5]), .B(addr_miss[5]), .Z(n_12770
		));
	notech_nand2 i_76060(.A(n_1075), .B(n_516), .Z(n_54255));
	notech_reg wrA_reg_6(.CP(n_61703), .D(n_12776), .CD(n_61006), .Q(wrA[6])
		);
	notech_mux2 i_18774(.S(n_53367), .A(wrA[6]), .B(addr_miss[6]), .Z(n_12776
		));
	notech_nand2 i_76063(.A(n_1074), .B(n_517), .Z(n_54261));
	notech_reg wrA_reg_7(.CP(n_61703), .D(n_12782), .CD(n_61006), .Q(wrA[7])
		);
	notech_mux2 i_18782(.S(n_53367), .A(wrA[7]), .B(addr_miss[7]), .Z(n_12782
		));
	notech_nand2 i_76066(.A(n_1073), .B(n_518), .Z(n_54267));
	notech_reg wrA_reg_8(.CP(n_61703), .D(n_12788), .CD(n_61006), .Q(wrA[8])
		);
	notech_mux2 i_18790(.S(n_53367), .A(wrA[8]), .B(addr_miss[8]), .Z(n_12788
		));
	notech_nand2 i_76069(.A(n_1072), .B(n_519), .Z(n_54273));
	notech_reg wrA_reg_9(.CP(n_61703), .D(n_12794), .CD(n_61006), .Q(wrA[9])
		);
	notech_mux2 i_18798(.S(n_53367), .A(wrA[9]), .B(addr_miss[9]), .Z(n_12794
		));
	notech_nand2 i_76072(.A(n_1071), .B(n_520), .Z(n_54279));
	notech_reg wrA_reg_10(.CP(n_61703), .D(n_12800), .CD(n_61006), .Q(wrA[10
		]));
	notech_mux2 i_18806(.S(n_53367), .A(wrA[10]), .B(addr_miss[10]), .Z(n_12800
		));
	notech_nand2 i_76075(.A(n_1070), .B(n_521), .Z(n_54285));
	notech_reg wrA_reg_11(.CP(n_61701), .D(n_12806), .CD(n_61004), .Q(wrA[11
		]));
	notech_mux2 i_18814(.S(n_53367), .A(wrA[11]), .B(addr_miss[11]), .Z(n_12806
		));
	notech_nand2 i_76078(.A(n_1069), .B(n_522), .Z(n_54291));
	notech_reg wrA_reg_12(.CP(n_61701), .D(n_12812), .CD(n_61004), .Q(wrA[12
		]));
	notech_mux2 i_18822(.S(n_53367), .A(wrA[12]), .B(addr_miss[12]), .Z(n_12812
		));
	notech_nand2 i_76081(.A(n_1068), .B(n_523), .Z(n_54297));
	notech_reg wrA_reg_13(.CP(n_61701), .D(n_12818), .CD(n_61004), .Q(wrA[13
		]));
	notech_mux2 i_18830(.S(n_53367), .A(wrA[13]), .B(addr_miss[13]), .Z(n_12818
		));
	notech_nand2 i_76084(.A(n_1067), .B(n_524), .Z(n_54303));
	notech_reg wrA_reg_14(.CP(n_61701), .D(n_12824), .CD(n_61004), .Q(wrA[14
		]));
	notech_mux2 i_18838(.S(n_53367), .A(wrA[14]), .B(addr_miss[14]), .Z(n_12824
		));
	notech_nand2 i_76087(.A(n_1066), .B(n_525), .Z(n_54309));
	notech_reg wrA_reg_15(.CP(n_61730), .D(n_12830), .CD(n_61033), .Q(wrA[15
		]));
	notech_mux2 i_18846(.S(n_53367), .A(wrA[15]), .B(addr_miss[15]), .Z(n_12830
		));
	notech_nand2 i_76090(.A(n_1065), .B(n_526), .Z(n_54315));
	notech_reg wrA_reg_16(.CP(n_61730), .D(n_12836), .CD(n_61033), .Q(wrA[16
		]));
	notech_mux2 i_18854(.S(n_53369), .A(wrA[16]), .B(addr_miss[16]), .Z(n_12836
		));
	notech_nand2 i_76093(.A(n_1064), .B(n_527), .Z(n_54321));
	notech_reg wrA_reg_17(.CP(n_61730), .D(n_12842), .CD(n_61033), .Q(wrA[17
		]));
	notech_mux2 i_18862(.S(n_53369), .A(wrA[17]), .B(addr_miss[17]), .Z(n_12842
		));
	notech_nand2 i_76096(.A(n_1063), .B(n_528), .Z(n_54327));
	notech_reg wrA_reg_18(.CP(n_61730), .D(n_12848), .CD(n_61033), .Q(wrA[18
		]));
	notech_mux2 i_18870(.S(n_53369), .A(wrA[18]), .B(addr_miss[18]), .Z(n_12848
		));
	notech_nand2 i_76099(.A(n_1062), .B(n_529), .Z(n_54333));
	notech_reg wrA_reg_19(.CP(n_61730), .D(n_12854), .CD(n_61033), .Q(wrA[19
		]));
	notech_mux2 i_18878(.S(n_53369), .A(wrA[19]), .B(addr_miss[19]), .Z(n_12854
		));
	notech_nand2 i_76102(.A(n_1061), .B(n_530), .Z(n_54339));
	notech_reg wrA_reg_20(.CP(n_61730), .D(n_12860), .CD(n_61033), .Q(wrA[20
		]));
	notech_mux2 i_18886(.S(n_53369), .A(wrA[20]), .B(addr_miss[20]), .Z(n_12860
		));
	notech_nand2 i_76105(.A(n_1060), .B(n_531), .Z(n_54345));
	notech_reg wrA_reg_21(.CP(n_61730), .D(n_12866), .CD(n_61033), .Q(wrA[21
		]));
	notech_mux2 i_18894(.S(n_53369), .A(wrA[21]), .B(addr_miss[21]), .Z(n_12866
		));
	notech_nand2 i_76108(.A(n_1059), .B(n_532), .Z(n_54351));
	notech_reg wrA_reg_22(.CP(n_61730), .D(n_12872), .CD(n_61033), .Q(wrA[22
		]));
	notech_mux2 i_18902(.S(n_53369), .A(wrA[22]), .B(addr_miss[22]), .Z(n_12872
		));
	notech_nand2 i_76111(.A(n_1058), .B(n_533), .Z(n_54357));
	notech_reg wrA_reg_23(.CP(n_61730), .D(n_12878), .CD(n_61033), .Q(wrA[23
		]));
	notech_mux2 i_18910(.S(n_53369), .A(wrA[23]), .B(addr_miss[23]), .Z(n_12878
		));
	notech_nand2 i_76114(.A(n_1057), .B(n_534), .Z(n_54363));
	notech_reg wrA_reg_24(.CP(n_61731), .D(n_12884), .CD(n_61034), .Q(wrA[24
		]));
	notech_mux2 i_18918(.S(n_53369), .A(wrA[24]), .B(addr_miss[24]), .Z(n_12884
		));
	notech_mux2 i_76015(.S(iwrite_ack), .A(n_538), .B(n_13489), .Z(n_55943)
		);
	notech_reg wrA_reg_25(.CP(n_61731), .D(n_12890), .CD(n_61034), .Q(wrA[25
		]));
	notech_mux2 i_18926(.S(n_53369), .A(wrA[25]), .B(addr_miss[25]), .Z(n_12890
		));
	notech_or4 i_41(.A(n_951), .B(n_1035), .C(n_13513), .D(n_13457), .Z(n_54148
		));
	notech_reg wrA_reg_26(.CP(n_61731), .D(n_12896), .CD(n_61034), .Q(wrA[26
		]));
	notech_mux2 i_18934(.S(n_53369), .A(wrA[26]), .B(addr_miss[26]), .Z(n_12896
		));
	notech_and4 i_42(.A(n_54796), .B(n_1038), .C(n_990), .D(n_957), .Z(n_54154
		));
	notech_reg wrA_reg_27(.CP(n_61731), .D(n_12902), .CD(n_61034), .Q(wrA[27
		]));
	notech_mux2 i_18942(.S(n_53369), .A(wrA[27]), .B(addr_miss[27]), .Z(n_12902
		));
	notech_or4 i_43(.A(n_549), .B(n_13614), .C(n_54807), .D(n_13459), .Z(n_54160
		));
	notech_reg wrA_reg_28(.CP(n_61731), .D(n_12908), .CD(n_61034), .Q(wrA[28
		]));
	notech_mux2 i_18950(.S(n_53369), .A(wrA[28]), .B(addr_miss[28]), .Z(n_12908
		));
	notech_or2 i_32(.A(n_54613), .B(\tab11_0[0] ), .Z(n_52377));
	notech_reg wrA_reg_29(.CP(n_61731), .D(n_12914), .CD(n_61034), .Q(wrA[29
		]));
	notech_mux2 i_18958(.S(n_53369), .A(wrA[29]), .B(addr_miss[29]), .Z(n_12914
		));
	notech_or2 i_33(.A(n_54613), .B(\tab11_0[1] ), .Z(n_52383));
	notech_reg wrA_reg_30(.CP(n_61731), .D(n_12920), .CD(n_61034), .Q(wrA[30
		]));
	notech_mux2 i_18966(.S(n_53369), .A(wrA[30]), .B(addr_miss[30]), .Z(n_12920
		));
	notech_or2 i_34(.A(n_54613), .B(\tab11_0[2] ), .Z(n_52389));
	notech_reg wrA_reg_31(.CP(n_61731), .D(n_12926), .CD(n_61034), .Q(wrA[31
		]));
	notech_mux2 i_18974(.S(n_53369), .A(wrA[31]), .B(addr_miss[31]), .Z(n_12926
		));
	notech_or2 i_35(.A(n_54613), .B(\tab11_0[3] ), .Z(n_52395));
	notech_reg addr_phys_reg_0(.CP(n_61731), .D(n_53761), .CD(n_61034), .Q(addr_phys
		[0]));
	notech_reg addr_phys_reg_1(.CP(n_61729), .D(n_53768), .CD(n_61032), .Q(addr_phys
		[1]));
	notech_reg addr_phys_reg_2(.CP(n_61729), .D(n_53775), .CD(n_61032), .Q(addr_phys
		[2]));
	notech_reg addr_phys_reg_3(.CP(n_61729), .D(n_53782), .CD(n_61032), .Q(addr_phys
		[3]));
	notech_reg addr_phys_reg_4(.CP(n_61729), .D(n_53789), .CD(n_61032), .Q(addr_phys
		[4]));
	notech_reg addr_phys_reg_5(.CP(n_61727), .D(n_53796), .CD(n_61030), .Q(addr_phys
		[5]));
	notech_reg addr_phys_reg_6(.CP(n_61727), .D(n_53803), .CD(n_61030), .Q(addr_phys
		[6]));
	notech_reg addr_phys_reg_7(.CP(n_61727), .D(n_53810), .CD(n_61030), .Q(addr_phys
		[7]));
	notech_reg addr_phys_reg_8(.CP(n_61727), .D(n_53817), .CD(n_61030), .Q(addr_phys
		[8]));
	notech_reg addr_phys_reg_9(.CP(n_61727), .D(n_53824), .CD(n_61030), .Q(addr_phys
		[9]));
	notech_reg addr_phys_reg_10(.CP(n_61729), .D(n_53831), .CD(n_61032), .Q(addr_phys
		[10]));
	notech_reg addr_phys_reg_11(.CP(n_61729), .D(n_53838), .CD(n_61032), .Q(addr_phys
		[11]));
	notech_reg addr_phys_reg_12(.CP(n_61730), .D(n_13682), .CD(n_61033), .Q(addr_phys
		[12]));
	notech_reg addr_phys_reg_13(.CP(n_61730), .D(n_13683), .CD(n_61033), .Q(addr_phys
		[13]));
	notech_reg addr_phys_reg_14(.CP(n_61729), .D(n_13684), .CD(n_61032), .Q(addr_phys
		[14]));
	notech_reg addr_phys_reg_15(.CP(n_61729), .D(n_13685), .CD(n_61032), .Q(addr_phys
		[15]));
	notech_reg addr_phys_reg_16(.CP(n_61729), .D(n_13686), .CD(n_61032), .Q(addr_phys
		[16]));
	notech_reg addr_phys_reg_17(.CP(n_61729), .D(n_13687), .CD(n_61032), .Q(addr_phys
		[17]));
	notech_reg addr_phys_reg_18(.CP(n_61729), .D(n_13688), .CD(n_61032), .Q(addr_phys
		[18]));
	notech_reg addr_phys_reg_19(.CP(n_61731), .D(n_13689), .CD(n_61034), .Q(addr_phys
		[19]));
	notech_reg addr_phys_reg_20(.CP(n_61736), .D(n_13690), .CD(n_61039), .Q(addr_phys
		[20]));
	notech_reg addr_phys_reg_21(.CP(n_61736), .D(n_13691), .CD(n_61039), .Q(addr_phys
		[21]));
	notech_reg addr_phys_reg_22(.CP(n_61736), .D(n_13692), .CD(n_61039), .Q(addr_phys
		[22]));
	notech_reg addr_phys_reg_23(.CP(n_61736), .D(n_13693), .CD(n_61039), .Q(addr_phys
		[23]));
	notech_reg addr_phys_reg_24(.CP(n_61735), .D(n_13694), .CD(n_61038), .Q(addr_phys
		[24]));
	notech_reg addr_phys_reg_25(.CP(n_61735), .D(n_13695), .CD(n_61038), .Q(addr_phys
		[25]));
	notech_reg addr_phys_reg_26(.CP(n_61735), .D(n_13696), .CD(n_61038), .Q(addr_phys
		[26]));
	notech_reg addr_phys_reg_27(.CP(n_61735), .D(n_13697), .CD(n_61038), .Q(addr_phys
		[27]));
	notech_reg addr_phys_reg_28(.CP(n_61735), .D(n_13698), .CD(n_61038), .Q(addr_phys
		[28]));
	notech_reg addr_phys_reg_29(.CP(n_61736), .D(n_13699), .CD(n_61039), .Q(addr_phys
		[29]));
	notech_reg addr_phys_reg_30(.CP(n_61736), .D(n_13700), .CD(n_61039), .Q(addr_phys
		[30]));
	notech_reg addr_phys_reg_31(.CP(n_61738), .D(n_13701), .CD(n_61041), .Q(addr_phys
		[31]));
	notech_reg wr_fault_reg(.CP(n_61738), .D(n_12996), .CD(n_61041), .Q(wr_fault
		));
	notech_mux2 i_19110(.S(n_53749), .A(wr_fault), .B(n_657), .Z(n_12996));
	notech_or2 i_36(.A(n_54613), .B(\tab11_0[5] ), .Z(n_52407));
	notech_reg pt_fault_reg(.CP(n_61736), .D(n_13002), .CD(n_61039), .Q(pt_fault
		));
	notech_mux2 i_19118(.S(n_656), .A(data_miss[0]), .B(pt_fault), .Z(n_13002
		));
	notech_or2 i_37(.A(n_54613), .B(\tab11_0[6] ), .Z(n_52413));
	notech_reg cr2_reg_0(.CP(n_61736), .D(n_13008), .CD(n_61039), .Q(cr2[0])
		);
	notech_mux2 i_19126(.S(n_656), .A(iDaddr_f[0]), .B(cr2[0]), .Z(n_13008)
		);
	notech_or2 i_38(.A(n_54613), .B(\tab11_0[7] ), .Z(n_52419));
	notech_reg cr2_reg_1(.CP(n_61736), .D(n_13014), .CD(n_61039), .Q(cr2[1])
		);
	notech_mux2 i_19134(.S(n_656), .A(iDaddr_f[1]), .B(cr2[1]), .Z(n_13014)
		);
	notech_or2 i_39(.A(n_54613), .B(\tab11_0[8] ), .Z(n_52425));
	notech_reg cr2_reg_2(.CP(n_61736), .D(n_13020), .CD(n_61039), .Q(cr2[2])
		);
	notech_mux2 i_19142(.S(n_656), .A(iDaddr_f[2]), .B(cr2[2]), .Z(n_13020)
		);
	notech_or2 i_40(.A(n_54613), .B(\tab11_0[9] ), .Z(n_52431));
	notech_reg cr2_reg_3(.CP(n_61736), .D(n_13026), .CD(n_61039), .Q(cr2[3])
		);
	notech_mux2 i_19150(.S(n_656), .A(iDaddr_f[3]), .B(cr2[3]), .Z(n_13026)
		);
	notech_or2 i_45(.A(data_miss[12]), .B(n_54613), .Z(n_52437));
	notech_reg cr2_reg_4(.CP(n_61734), .D(n_13032), .CD(n_61037), .Q(cr2[4])
		);
	notech_mux2 i_19158(.S(n_656), .A(iDaddr_f[4]), .B(cr2[4]), .Z(n_13032)
		);
	notech_or2 i_47(.A(data_miss[13]), .B(n_54613), .Z(n_52443));
	notech_reg cr2_reg_5(.CP(n_61734), .D(n_13038), .CD(n_61037), .Q(cr2[5])
		);
	notech_mux2 i_19166(.S(n_656), .A(iDaddr_f[5]), .B(cr2[5]), .Z(n_13038)
		);
	notech_or2 i_48(.A(data_miss[14]), .B(n_54608), .Z(n_52449));
	notech_reg cr2_reg_6(.CP(n_61734), .D(n_13044), .CD(n_61037), .Q(cr2[6])
		);
	notech_mux2 i_19174(.S(n_656), .A(iDaddr_f[6]), .B(cr2[6]), .Z(n_13044)
		);
	notech_or2 i_49(.A(data_miss[15]), .B(n_54608), .Z(n_52455));
	notech_reg cr2_reg_7(.CP(n_61734), .D(n_13050), .CD(n_61037), .Q(cr2[7])
		);
	notech_mux2 i_19182(.S(n_656), .A(iDaddr_f[7]), .B(cr2[7]), .Z(n_13050)
		);
	notech_or2 i_51(.A(data_miss[16]), .B(n_54608), .Z(n_52461));
	notech_reg cr2_reg_8(.CP(n_61734), .D(n_13056), .CD(n_61037), .Q(cr2[8])
		);
	notech_mux2 i_19190(.S(n_656), .A(iDaddr_f[8]), .B(cr2[8]), .Z(n_13056)
		);
	notech_or2 i_52(.A(data_miss[17]), .B(n_54608), .Z(n_52467));
	notech_reg cr2_reg_9(.CP(n_61734), .D(n_13062), .CD(n_61037), .Q(cr2[9])
		);
	notech_mux2 i_19198(.S(n_656), .A(iDaddr_f[9]), .B(cr2[9]), .Z(n_13062)
		);
	notech_or2 i_53(.A(data_miss[18]), .B(n_54608), .Z(n_52473));
	notech_reg cr2_reg_10(.CP(n_61731), .D(n_13068), .CD(n_61034), .Q(cr2[10
		]));
	notech_mux2 i_19206(.S(n_656), .A(iDaddr_f[10]), .B(cr2[10]), .Z(n_13068
		));
	notech_or2 i_54(.A(data_miss[19]), .B(n_54608), .Z(n_52479));
	notech_reg cr2_reg_11(.CP(n_61734), .D(n_13074), .CD(n_61037), .Q(cr2[11
		]));
	notech_mux2 i_19214(.S(n_656), .A(iDaddr_f[11]), .B(cr2[11]), .Z(n_13074
		));
	notech_or2 i_55(.A(data_miss[20]), .B(n_54608), .Z(n_52485));
	notech_reg cr2_reg_12(.CP(n_61734), .D(n_13080), .CD(n_61037), .Q(cr2[12
		]));
	notech_mux2 i_19222(.S(n_656), .A(iDaddr_f[12]), .B(cr2[12]), .Z(n_13080
		));
	notech_or2 i_56(.A(data_miss[21]), .B(n_54608), .Z(n_52491));
	notech_reg cr2_reg_13(.CP(n_61735), .D(n_13086), .CD(n_61038), .Q(cr2[13
		]));
	notech_mux2 i_19230(.S(n_656), .A(iDaddr_f[13]), .B(cr2[13]), .Z(n_13086
		));
	notech_or2 i_57(.A(data_miss[22]), .B(n_54608), .Z(n_52497));
	notech_reg cr2_reg_14(.CP(n_61735), .D(n_13092), .CD(n_61038), .Q(cr2[14
		]));
	notech_mux2 i_19238(.S(n_656), .A(iDaddr_f[14]), .B(cr2[14]), .Z(n_13092
		));
	notech_or2 i_58(.A(data_miss[23]), .B(n_54608), .Z(n_52503));
	notech_reg cr2_reg_15(.CP(n_61735), .D(n_13098), .CD(n_61038), .Q(cr2[15
		]));
	notech_mux2 i_19246(.S(n_656), .A(iDaddr_f[15]), .B(cr2[15]), .Z(n_13098
		));
	notech_or2 i_59(.A(data_miss[24]), .B(n_54608), .Z(n_52509));
	notech_reg cr2_reg_16(.CP(n_61735), .D(n_13104), .CD(n_61038), .Q(cr2[16
		]));
	notech_mux2 i_19254(.S(n_53621), .A(iDaddr_f[16]), .B(cr2[16]), .Z(n_13104
		));
	notech_or2 i_60(.A(data_miss[25]), .B(n_54613), .Z(n_52515));
	notech_reg cr2_reg_17(.CP(n_61735), .D(n_13110), .CD(n_61038), .Q(cr2[17
		]));
	notech_mux2 i_19262(.S(n_53621), .A(iDaddr_f[17]), .B(cr2[17]), .Z(n_13110
		));
	notech_or2 i_61(.A(data_miss[26]), .B(n_54608), .Z(n_52521));
	notech_reg cr2_reg_18(.CP(n_61734), .D(n_13116), .CD(n_61037), .Q(cr2[18
		]));
	notech_mux2 i_19270(.S(n_53621), .A(iDaddr_f[18]), .B(cr2[18]), .Z(n_13116
		));
	notech_or2 i_62(.A(data_miss[27]), .B(n_54608), .Z(n_52527));
	notech_reg cr2_reg_19(.CP(n_61734), .D(n_13122), .CD(n_61037), .Q(cr2[19
		]));
	notech_mux2 i_19278(.S(n_53621), .A(iDaddr_f[19]), .B(cr2[19]), .Z(n_13122
		));
	notech_or2 i_63(.A(data_miss[28]), .B(n_54608), .Z(n_52533));
	notech_reg cr2_reg_20(.CP(n_61735), .D(n_13128), .CD(n_61038), .Q(cr2[20
		]));
	notech_mux2 i_19286(.S(n_53621), .A(iDaddr_f[20]), .B(cr2[20]), .Z(n_13128
		));
	notech_or2 i_64(.A(data_miss[29]), .B(n_54608), .Z(n_52539));
	notech_reg cr2_reg_21(.CP(n_61734), .D(n_13134), .CD(n_61037), .Q(cr2[21
		]));
	notech_mux2 i_19294(.S(n_53621), .A(iDaddr_f[21]), .B(cr2[21]), .Z(n_13134
		));
	notech_or2 i_65(.A(data_miss[30]), .B(n_54608), .Z(n_52545));
	notech_reg cr2_reg_22(.CP(n_61727), .D(n_13140), .CD(n_61030), .Q(cr2[22
		]));
	notech_mux2 i_19302(.S(n_53621), .A(iDaddr_f[22]), .B(cr2[22]), .Z(n_13140
		));
	notech_or2 i_66(.A(data_miss[31]), .B(n_54608), .Z(n_52551));
	notech_reg cr2_reg_23(.CP(n_61720), .D(n_13146), .CD(n_61023), .Q(cr2[23
		]));
	notech_mux2 i_19310(.S(n_53621), .A(iDaddr_f[23]), .B(cr2[23]), .Z(n_13146
		));
	notech_nand2 i_031214(.A(n_989), .B(n_58627), .Z(n_52575));
	notech_reg cr2_reg_24(.CP(n_61719), .D(n_13152), .CD(n_61022), .Q(cr2[24
		]));
	notech_mux2 i_19318(.S(n_53621), .A(iDaddr_f[24]), .B(cr2[24]), .Z(n_13152
		));
	notech_ao4 i_76771(.A(n_996), .B(n_13606), .C(n_559), .D(n_1026), .Z(n_55457
		));
	notech_reg cr2_reg_25(.CP(n_61720), .D(n_13158), .CD(n_61023), .Q(cr2[25
		]));
	notech_mux2 i_19326(.S(n_53621), .A(iDaddr_f[25]), .B(cr2[25]), .Z(n_13158
		));
	notech_ao4 i_76774(.A(n_996), .B(n_13608), .C(n_564), .D(n_1026), .Z(n_55463
		));
	notech_reg cr2_reg_26(.CP(n_61720), .D(n_13164), .CD(n_61023), .Q(cr2[26
		]));
	notech_mux2 i_19334(.S(n_656), .A(iDaddr_f[26]), .B(cr2[26]), .Z(n_13164
		));
	notech_ao4 i_76761(.A(n_1016), .B(n_13611), .C(n_996), .D(\nnx_tab2[0] )
		, .Z(n_54069));
	notech_reg cr2_reg_27(.CP(n_61719), .D(n_13170), .CD(n_61022), .Q(cr2[27
		]));
	notech_mux2 i_19342(.S(n_53621), .A(iDaddr_f[27]), .B(cr2[27]), .Z(n_13170
		));
	notech_ao4 i_76764(.A(n_1016), .B(n_13613), .C(n_996), .D(n_573), .Z(n_54075
		));
	notech_reg cr2_reg_28(.CP(n_61719), .D(n_13176), .CD(n_61022), .Q(cr2[28
		]));
	notech_mux2 i_19350(.S(n_53621), .A(iDaddr_f[28]), .B(cr2[28]), .Z(n_13176
		));
	notech_ao4 i_76542(.A(n_1016), .B(n_13536), .C(n_996), .D(\nnx_tab1[0] )
		, .Z(n_54104));
	notech_reg cr2_reg_29(.CP(n_61719), .D(n_13182), .CD(n_61022), .Q(cr2[29
		]));
	notech_mux2 i_19358(.S(n_53621), .A(iDaddr_f[29]), .B(cr2[29]), .Z(n_13182
		));
	notech_ao4 i_76545(.A(n_1016), .B(n_13538), .C(n_996), .D(n_585), .Z(n_54110
		));
	notech_reg cr2_reg_30(.CP(n_61719), .D(n_13188), .CD(n_61022), .Q(cr2[30
		]));
	notech_mux2 i_19366(.S(n_53621), .A(iDaddr_f[30]), .B(cr2[30]), .Z(n_13188
		));
	notech_ao4 i_76791(.A(n_996), .B(n_13540), .C(n_590), .D(n_1017), .Z(n_55482
		));
	notech_reg cr2_reg_31(.CP(n_61719), .D(n_13194), .CD(n_61022), .Q(cr2[31
		]));
	notech_mux2 i_19374(.S(n_53621), .A(iDaddr_f[31]), .B(cr2[31]), .Z(n_13194
		));
	notech_ao4 i_76794(.A(n_996), .B(n_13542), .C(n_595), .D(n_1017), .Z(n_55488
		));
	notech_reg wrD_reg_0(.CP(n_61720), .D(n_13200), .CD(n_61023), .Q(wrD[0])
		);
	notech_or2 i_19382(.A(wrD[0]), .B(n_53362), .Z(n_13200));
	notech_nand2 i_99(.A(n_55715), .B(n_13767), .Z(n_55516));
	notech_reg wrD_reg_1(.CP(n_61720), .D(n_13206), .CD(n_61023), .Q(wrD[1])
		);
	notech_mux2 i_19390(.S(n_53362), .A(wrD[1]), .B(data_miss[1]), .Z(n_13206
		));
	notech_nand2 i_100(.A(n_55715), .B(n_13766), .Z(n_55522));
	notech_reg wrD_reg_2(.CP(n_61721), .D(n_13212), .CD(n_61024), .Q(wrD[2])
		);
	notech_mux2 i_19398(.S(n_53362), .A(wrD[2]), .B(data_miss[2]), .Z(n_13212
		));
	notech_nand2 i_101(.A(n_55715), .B(n_13765), .Z(n_55528));
	notech_reg wrD_reg_3(.CP(n_61720), .D(n_13218), .CD(n_61023), .Q(wrD[3])
		);
	notech_mux2 i_19406(.S(n_53362), .A(wrD[3]), .B(data_miss[3]), .Z(n_13218
		));
	notech_nand2 i_102(.A(n_55715), .B(n_13764), .Z(n_55534));
	notech_reg wrD_reg_4(.CP(n_61720), .D(n_13224), .CD(n_61023), .Q(wrD[4])
		);
	notech_mux2 i_19414(.S(n_53362), .A(wrD[4]), .B(data_miss[4]), .Z(n_13224
		));
	notech_nand2 i_103(.A(n_55715), .B(n_13762), .Z(n_55546));
	notech_reg wrD_reg_5(.CP(n_61720), .D(n_13230), .CD(n_61023), .Q(wrD[5])
		);
	notech_mux2 i_19422(.S(n_53362), .A(wrD[5]), .B(n_52185), .Z(n_13230));
	notech_nand2 i_104(.A(n_55715), .B(n_13761), .Z(n_55552));
	notech_reg wrD_reg_6(.CP(n_61720), .D(n_13236), .CD(n_61023), .Q(wrD[6])
		);
	notech_mux2 i_19430(.S(n_53362), .A(wrD[6]), .B(n_52191), .Z(n_13236));
	notech_nand2 i_105(.A(n_55715), .B(n_13760), .Z(n_55558));
	notech_reg wrD_reg_7(.CP(n_61720), .D(n_13242), .CD(n_61023), .Q(wrD[7])
		);
	notech_mux2 i_19438(.S(n_53362), .A(wrD[7]), .B(data_miss[7]), .Z(n_13242
		));
	notech_nand2 i_106(.A(n_55715), .B(n_13759), .Z(n_55564));
	notech_reg wrD_reg_8(.CP(n_61720), .D(n_13248), .CD(n_61023), .Q(wrD[8])
		);
	notech_mux2 i_19446(.S(n_53362), .A(wrD[8]), .B(data_miss[8]), .Z(n_13248
		));
	notech_nand2 i_107(.A(n_55715), .B(n_13758), .Z(n_55570));
	notech_reg wrD_reg_9(.CP(n_61717), .D(n_13254), .CD(n_61020), .Q(wrD[9])
		);
	notech_mux2 i_19454(.S(n_53362), .A(wrD[9]), .B(data_miss[9]), .Z(n_13254
		));
	notech_or2 i_108(.A(data_miss[12]), .B(n_13488), .Z(n_55576));
	notech_reg wrD_reg_10(.CP(n_61717), .D(n_13260), .CD(n_61020), .Q(wrD[10
		]));
	notech_mux2 i_19462(.S(n_53362), .A(wrD[10]), .B(data_miss[10]), .Z(n_13260
		));
	notech_or2 i_109(.A(data_miss[13]), .B(n_13488), .Z(n_55582));
	notech_reg wrD_reg_11(.CP(n_61717), .D(n_13266), .CD(n_61020), .Q(wrD[11
		]));
	notech_mux2 i_19470(.S(n_53362), .A(wrD[11]), .B(data_miss[11]), .Z(n_13266
		));
	notech_or2 i_110(.A(data_miss[14]), .B(n_13488), .Z(n_55588));
	notech_reg wrD_reg_12(.CP(n_61717), .D(n_13272), .CD(n_61020), .Q(wrD[12
		]));
	notech_mux2 i_19478(.S(n_53362), .A(wrD[12]), .B(data_miss[12]), .Z(n_13272
		));
	notech_or2 i_111(.A(data_miss[15]), .B(n_13488), .Z(n_55594));
	notech_reg wrD_reg_13(.CP(n_61717), .D(n_13278), .CD(n_61020), .Q(wrD[13
		]));
	notech_mux2 i_19486(.S(n_53362), .A(wrD[13]), .B(data_miss[13]), .Z(n_13278
		));
	notech_or2 i_112(.A(data_miss[16]), .B(n_13488), .Z(n_55600));
	notech_reg wrD_reg_14(.CP(n_61716), .D(n_13284), .CD(n_61019), .Q(wrD[14
		]));
	notech_mux2 i_19494(.S(n_53362), .A(wrD[14]), .B(data_miss[14]), .Z(n_13284
		));
	notech_or2 i_113(.A(data_miss[17]), .B(n_13488), .Z(n_55606));
	notech_reg wrD_reg_15(.CP(n_61716), .D(n_13290), .CD(n_61019), .Q(wrD[15
		]));
	notech_mux2 i_19502(.S(n_53362), .A(wrD[15]), .B(data_miss[15]), .Z(n_13290
		));
	notech_or2 i_114(.A(data_miss[18]), .B(n_13488), .Z(n_55612));
	notech_reg wrD_reg_16(.CP(n_61717), .D(n_13296), .CD(n_61020), .Q(wrD[16
		]));
	notech_mux2 i_19510(.S(n_53364), .A(wrD[16]), .B(data_miss[16]), .Z(n_13296
		));
	notech_or2 i_115(.A(data_miss[19]), .B(n_13488), .Z(n_55618));
	notech_reg wrD_reg_17(.CP(n_61717), .D(n_13302), .CD(n_61020), .Q(wrD[17
		]));
	notech_mux2 i_19518(.S(n_53364), .A(wrD[17]), .B(data_miss[17]), .Z(n_13302
		));
	notech_or2 i_116(.A(data_miss[20]), .B(n_13488), .Z(n_55624));
	notech_reg wrD_reg_18(.CP(n_61719), .D(n_13308), .CD(n_61022), .Q(wrD[18
		]));
	notech_mux2 i_19526(.S(n_53364), .A(wrD[18]), .B(data_miss[18]), .Z(n_13308
		));
	notech_or2 i_117(.A(data_miss[21]), .B(n_54628), .Z(n_55630));
	notech_reg wrD_reg_19(.CP(n_61719), .D(n_13314), .CD(n_61022), .Q(wrD[19
		]));
	notech_mux2 i_19534(.S(n_53364), .A(wrD[19]), .B(data_miss[19]), .Z(n_13314
		));
	notech_or2 i_118(.A(data_miss[22]), .B(n_54628), .Z(n_55636));
	notech_reg wrD_reg_20(.CP(n_61719), .D(n_13320), .CD(n_61022), .Q(wrD[20
		]));
	notech_mux2 i_19542(.S(n_53364), .A(wrD[20]), .B(data_miss[20]), .Z(n_13320
		));
	notech_or2 i_119(.A(data_miss[23]), .B(n_54628), .Z(n_55642));
	notech_reg wrD_reg_21(.CP(n_61719), .D(n_13326), .CD(n_61022), .Q(wrD[21
		]));
	notech_mux2 i_19550(.S(n_53364), .A(wrD[21]), .B(data_miss[21]), .Z(n_13326
		));
	notech_or2 i_120(.A(data_miss[24]), .B(n_54628), .Z(n_55648));
	notech_reg wrD_reg_22(.CP(n_61719), .D(n_13332), .CD(n_61022), .Q(wrD[22
		]));
	notech_mux2 i_19558(.S(n_53364), .A(wrD[22]), .B(data_miss[22]), .Z(n_13332
		));
	notech_or2 i_121(.A(data_miss[25]), .B(n_54628), .Z(n_55654));
	notech_reg wrD_reg_23(.CP(n_61717), .D(n_13338), .CD(n_61020), .Q(wrD[23
		]));
	notech_mux2 i_19566(.S(n_53364), .A(wrD[23]), .B(data_miss[23]), .Z(n_13338
		));
	notech_or2 i_122(.A(data_miss[26]), .B(n_54628), .Z(n_55660));
	notech_reg wrD_reg_24(.CP(n_61717), .D(n_13344), .CD(n_61020), .Q(wrD[24
		]));
	notech_mux2 i_19574(.S(n_53364), .A(wrD[24]), .B(data_miss[24]), .Z(n_13344
		));
	notech_or2 i_123(.A(data_miss[27]), .B(n_54628), .Z(n_55666));
	notech_reg wrD_reg_25(.CP(n_61717), .D(n_13350), .CD(n_61020), .Q(wrD[25
		]));
	notech_mux2 i_19582(.S(n_53364), .A(wrD[25]), .B(data_miss[25]), .Z(n_13350
		));
	notech_or2 i_124(.A(data_miss[28]), .B(n_13488), .Z(n_55672));
	notech_reg wrD_reg_26(.CP(n_61717), .D(n_13356), .CD(n_61020), .Q(wrD[26
		]));
	notech_mux2 i_19590(.S(n_53364), .A(wrD[26]), .B(data_miss[26]), .Z(n_13356
		));
	notech_or2 i_125(.A(data_miss[29]), .B(n_54628), .Z(n_55678));
	notech_reg wrD_reg_27(.CP(n_61721), .D(n_13362), .CD(n_61024), .Q(wrD[27
		]));
	notech_mux2 i_19598(.S(n_53364), .A(wrD[27]), .B(data_miss[27]), .Z(n_13362
		));
	notech_or2 i_126(.A(data_miss[30]), .B(n_54628), .Z(n_55684));
	notech_reg wrD_reg_28(.CP(n_61726), .D(n_13368), .CD(n_61029), .Q(wrD[28
		]));
	notech_mux2 i_19606(.S(n_53364), .A(wrD[28]), .B(data_miss[28]), .Z(n_13368
		));
	notech_or2 i_127(.A(data_miss[31]), .B(n_54628), .Z(n_55690));
	notech_reg wrD_reg_29(.CP(n_61726), .D(n_13374), .CD(n_61029), .Q(wrD[29
		]));
	notech_mux2 i_19614(.S(n_53364), .A(wrD[29]), .B(data_miss[29]), .Z(n_13374
		));
	notech_ao4 i_3(.A(data_miss[0]), .B(n_989), .C(n_984), .D(n_985), .Z(n_55715
		));
	notech_reg wrD_reg_30(.CP(n_61726), .D(n_13380), .CD(n_61029), .Q(wrD[30
		]));
	notech_mux2 i_19622(.S(n_53364), .A(wrD[30]), .B(data_miss[30]), .Z(n_13380
		));
	notech_reg wrD_reg_31(.CP(n_61726), .D(n_13386), .CD(n_61029), .Q(wrD[31
		]));
	notech_mux2 i_19630(.S(n_53364), .A(wrD[31]), .B(data_miss[31]), .Z(n_13386
		));
	notech_reg owrite_data_reg_0(.CP(n_61726), .D(n_53009), .CD(n_61029), .Q
		(owrite_data[0]));
	notech_reg owrite_data_reg_1(.CP(n_61725), .D(n_53016), .CD(n_61028), .Q
		(owrite_data[1]));
	notech_reg owrite_data_reg_2(.CP(n_61725), .D(n_53023), .CD(n_61028), .Q
		(owrite_data[2]));
	notech_reg owrite_data_reg_3(.CP(n_61726), .D(n_53030), .CD(n_61029), .Q
		(owrite_data[3]));
	notech_reg owrite_data_reg_4(.CP(n_61726), .D(n_53037), .CD(n_61029), .Q
		(owrite_data[4]));
	notech_reg owrite_data_reg_5(.CP(n_61727), .D(n_53044), .CD(n_61030), .Q
		(owrite_data[5]));
	notech_reg owrite_data_reg_6(.CP(n_61727), .D(n_53051), .CD(n_61030), .Q
		(owrite_data[6]));
	notech_reg owrite_data_reg_7(.CP(n_61727), .D(n_53058), .CD(n_61030), .Q
		(owrite_data[7]));
	notech_reg owrite_data_reg_8(.CP(n_61727), .D(n_53065), .CD(n_61030), .Q
		(owrite_data[8]));
	notech_reg owrite_data_reg_9(.CP(n_61727), .D(n_53072), .CD(n_61030), .Q
		(owrite_data[9]));
	notech_reg owrite_data_reg_10(.CP(n_61726), .D(n_53079), .CD(n_61029), .Q
		(owrite_data[10]));
	notech_reg owrite_data_reg_11(.CP(n_61726), .D(n_53086), .CD(n_61029), .Q
		(owrite_data[11]));
	notech_reg owrite_data_reg_12(.CP(n_61726), .D(n_53093), .CD(n_61029), .Q
		(owrite_data[12]));
	notech_reg owrite_data_reg_13(.CP(n_61726), .D(n_53100), .CD(n_61029), .Q
		(owrite_data[13]));
	notech_reg owrite_data_reg_14(.CP(n_61721), .D(n_53107), .CD(n_61024), .Q
		(owrite_data[14]));
	notech_reg owrite_data_reg_15(.CP(n_61721), .D(n_53114), .CD(n_61024), .Q
		(owrite_data[15]));
	notech_reg owrite_data_reg_16(.CP(n_61721), .D(n_53121), .CD(n_61024), .Q
		(owrite_data[16]));
	notech_reg owrite_data_reg_17(.CP(n_61721), .D(n_53128), .CD(n_61024), .Q
		(owrite_data[17]));
	notech_reg owrite_data_reg_18(.CP(n_61721), .D(n_53135), .CD(n_61024), .Q
		(owrite_data[18]));
	notech_reg owrite_data_reg_19(.CP(n_61721), .D(n_53142), .CD(n_61024), .Q
		(owrite_data[19]));
	notech_reg owrite_data_reg_20(.CP(n_61721), .D(n_53149), .CD(n_61024), .Q
		(owrite_data[20]));
	notech_reg owrite_data_reg_21(.CP(n_61721), .D(n_53156), .CD(n_61024), .Q
		(owrite_data[21]));
	notech_reg owrite_data_reg_22(.CP(n_61721), .D(n_53163), .CD(n_61024), .Q
		(owrite_data[22]));
	notech_reg owrite_data_reg_23(.CP(n_61725), .D(n_53170), .CD(n_61028), .Q
		(owrite_data[23]));
	notech_reg owrite_data_reg_24(.CP(n_61725), .D(n_53177), .CD(n_61028), .Q
		(owrite_data[24]));
	notech_reg owrite_data_reg_25(.CP(n_61725), .D(n_53184), .CD(n_61028), .Q
		(owrite_data[25]));
	notech_reg owrite_data_reg_26(.CP(n_61725), .D(n_53191), .CD(n_61028), .Q
		(owrite_data[26]));
	notech_reg owrite_data_reg_27(.CP(n_61725), .D(n_53198), .CD(n_61028), .Q
		(owrite_data[27]));
	notech_reg owrite_data_reg_28(.CP(n_61725), .D(n_53205), .CD(n_61028), .Q
		(owrite_data[28]));
	notech_reg owrite_data_reg_29(.CP(n_61725), .D(n_53212), .CD(n_61028), .Q
		(owrite_data[29]));
	notech_reg owrite_data_reg_30(.CP(n_61725), .D(n_53219), .CD(n_61028), .Q
		(owrite_data[30]));
	notech_reg owrite_data_reg_31(.CP(n_61725), .D(n_53226), .CD(n_61028), .Q
		(owrite_data[31]));
	notech_inv i_21454(.A(n_1050), .Z(n_13457));
	notech_inv i_21455(.A(n_54796), .Z(n_13458));
	notech_inv i_21456(.A(n_1033), .Z(n_13459));
	notech_inv i_21457(.A(n_1016), .Z(n_13460));
	notech_inv i_21458(.A(n_987), .Z(n_13461));
	notech_inv i_21459(.A(n_999), .Z(n_13462));
	notech_inv i_21460(.A(n_53473), .Z(n_13463));
	notech_inv i_21461(.A(n_985), .Z(n_13464));
	notech_inv i_21462(.A(n_983), .Z(n_13465));
	notech_inv i_21463(.A(n_1011), .Z(n_13466));
	notech_inv i_21464(.A(\dir1[10] ), .Z(n_13467));
	notech_inv i_21465(.A(\dir1[11] ), .Z(n_13468));
	notech_inv i_21466(.A(\dir1[12] ), .Z(n_13469));
	notech_inv i_21467(.A(\dir1[13] ), .Z(n_13470));
	notech_inv i_21468(.A(\dir1[14] ), .Z(n_13471));
	notech_inv i_21469(.A(\dir1[15] ), .Z(n_13472));
	notech_inv i_21470(.A(\dir1[16] ), .Z(n_13473));
	notech_inv i_21471(.A(\dir1[17] ), .Z(n_13474));
	notech_inv i_21472(.A(\dir1[18] ), .Z(n_13475));
	notech_inv i_21473(.A(\dir1[19] ), .Z(n_13476));
	notech_inv i_21474(.A(\dir1[20] ), .Z(n_13477));
	notech_inv i_21475(.A(\dir1[21] ), .Z(n_13478));
	notech_inv i_21476(.A(\dir1[22] ), .Z(n_13479));
	notech_inv i_21477(.A(\dir1[23] ), .Z(n_13480));
	notech_inv i_21478(.A(\dir1[24] ), .Z(n_13481));
	notech_inv i_21479(.A(\dir1[25] ), .Z(n_13482));
	notech_inv i_21480(.A(\dir1[26] ), .Z(n_13483));
	notech_inv i_21481(.A(n_494), .Z(n_13484));
	notech_inv i_21482(.A(\dir1[27] ), .Z(n_13485));
	notech_inv i_21483(.A(\dir1[28] ), .Z(n_13486));
	notech_inv i_21484(.A(\dir1[29] ), .Z(n_13487));
	notech_inv i_21485(.A(n_55715), .Z(n_13488));
	notech_inv i_21486(.A(n_536), .Z(n_13489));
	notech_inv i_21487(.A(n_571), .Z(n_13490));
	notech_inv i_21488(.A(\tab12[10] ), .Z(n_13491));
	notech_inv i_21489(.A(\tab12[11] ), .Z(n_13492));
	notech_inv i_21490(.A(\tab12[12] ), .Z(n_13493));
	notech_inv i_21491(.A(\tab12[13] ), .Z(n_13494));
	notech_inv i_21492(.A(\tab12[14] ), .Z(n_13495));
	notech_inv i_21493(.A(\tab12[15] ), .Z(n_13496));
	notech_inv i_21494(.A(\tab12[16] ), .Z(n_13497));
	notech_inv i_21495(.A(\tab12[17] ), .Z(n_13498));
	notech_inv i_21496(.A(n_583), .Z(n_13499));
	notech_inv i_21497(.A(\tab12[18] ), .Z(n_13500));
	notech_inv i_21498(.A(\tab12[19] ), .Z(n_13501));
	notech_inv i_21499(.A(\tab12[20] ), .Z(n_13502));
	notech_inv i_21500(.A(\tab12[21] ), .Z(n_13503));
	notech_inv i_21501(.A(\tab12[22] ), .Z(n_13504));
	notech_inv i_21502(.A(\tab12[23] ), .Z(n_13505));
	notech_inv i_21503(.A(\tab12[24] ), .Z(n_13506));
	notech_inv i_21504(.A(\tab12[25] ), .Z(n_13507));
	notech_inv i_21505(.A(\tab12[26] ), .Z(n_13508));
	notech_inv i_21506(.A(\tab12[27] ), .Z(n_13509));
	notech_inv i_21507(.A(\tab12[28] ), .Z(n_13510));
	notech_inv i_21508(.A(\tab12[29] ), .Z(n_13511));
	notech_inv i_21509(.A(hit_adr12), .Z(n_13512));
	notech_inv i_21510(.A(n_58627), .Z(n_13513));
	notech_inv i_21511(.A(n_606), .Z(n_50997));
	notech_inv i_21512(.A(\tab14[10] ), .Z(n_13515));
	notech_inv i_21513(.A(\tab14[11] ), .Z(n_13516));
	notech_inv i_21514(.A(\tab14[12] ), .Z(n_13517));
	notech_inv i_21515(.A(\tab14[13] ), .Z(n_13518));
	notech_inv i_21516(.A(\tab14[14] ), .Z(n_13519));
	notech_inv i_21517(.A(\tab14[15] ), .Z(n_13520));
	notech_inv i_21518(.A(\tab14[16] ), .Z(n_13521));
	notech_inv i_21519(.A(\tab14[17] ), .Z(n_13522));
	notech_inv i_21520(.A(\tab14[18] ), .Z(n_13523));
	notech_inv i_21521(.A(\tab14[19] ), .Z(n_13524));
	notech_inv i_21522(.A(\tab14[20] ), .Z(n_13525));
	notech_inv i_21523(.A(\tab14[21] ), .Z(n_13526));
	notech_inv i_21524(.A(\tab14[22] ), .Z(n_13527));
	notech_inv i_21525(.A(\tab14[23] ), .Z(n_13528));
	notech_inv i_21526(.A(\tab14[24] ), .Z(n_13529));
	notech_inv i_21527(.A(\tab14[25] ), .Z(n_13530));
	notech_inv i_21528(.A(\tab14[26] ), .Z(n_13531));
	notech_inv i_21529(.A(\tab14[27] ), .Z(n_13532));
	notech_inv i_21530(.A(\tab14[28] ), .Z(n_13533));
	notech_inv i_21531(.A(\tab14[29] ), .Z(n_13534));
	notech_inv i_21532(.A(n_55482), .Z(n_13535));
	notech_inv i_21533(.A(\nx_tab1[0] ), .Z(n_13536));
	notech_inv i_21534(.A(n_55488), .Z(n_13537));
	notech_inv i_21535(.A(\nx_tab1[1] ), .Z(n_13538));
	notech_inv i_21536(.A(n_54104), .Z(n_13539));
	notech_inv i_21537(.A(\nnx_tab1[0] ), .Z(n_13540));
	notech_inv i_21538(.A(n_54110), .Z(n_13541));
	notech_inv i_21539(.A(\nnx_tab1[1] ), .Z(n_13542));
	notech_inv i_21540(.A(\nbus_14031[0] ), .Z(n_13543));
	notech_inv i_21541(.A(\tab22[10] ), .Z(n_13544));
	notech_inv i_21542(.A(\tab22[11] ), .Z(n_13545));
	notech_inv i_21543(.A(\tab22[12] ), .Z(n_13546));
	notech_inv i_21544(.A(\tab22[13] ), .Z(n_13547));
	notech_inv i_21545(.A(\tab22[14] ), .Z(n_13548));
	notech_inv i_21546(.A(\tab22[15] ), .Z(n_13549));
	notech_inv i_21547(.A(\tab22[16] ), .Z(n_13550));
	notech_inv i_21548(.A(\tab22[17] ), .Z(n_13551));
	notech_inv i_21549(.A(\tab22[18] ), .Z(n_13552));
	notech_inv i_21550(.A(\tab22[19] ), .Z(n_13553));
	notech_inv i_21551(.A(\tab22[20] ), .Z(n_13554));
	notech_inv i_21552(.A(\tab22[21] ), .Z(n_13555));
	notech_inv i_21553(.A(\tab22[22] ), .Z(n_13556));
	notech_inv i_21554(.A(\tab22[23] ), .Z(n_13557));
	notech_inv i_21555(.A(\tab22[24] ), .Z(n_13558));
	notech_inv i_21556(.A(\tab22[25] ), .Z(n_13559));
	notech_inv i_21557(.A(\tab22[26] ), .Z(n_13560));
	notech_inv i_21558(.A(\tab22[27] ), .Z(n_13561));
	notech_inv i_21559(.A(\tab22[28] ), .Z(n_13562));
	notech_inv i_21560(.A(\tab22[29] ), .Z(n_13563));
	notech_inv i_21561(.A(hit_adr22), .Z(n_13564));
	notech_inv i_21562(.A(\tab23[10] ), .Z(n_13565));
	notech_inv i_21563(.A(\tab23[11] ), .Z(n_13566));
	notech_inv i_21564(.A(\tab23[12] ), .Z(n_13567));
	notech_inv i_21565(.A(\tab23[13] ), .Z(n_13568));
	notech_inv i_21566(.A(\tab23[14] ), .Z(n_13569));
	notech_inv i_21567(.A(\tab23[15] ), .Z(n_13570));
	notech_inv i_21568(.A(\tab23[16] ), .Z(n_13571));
	notech_inv i_21569(.A(\tab23[17] ), .Z(n_13572));
	notech_inv i_21570(.A(\tab23[18] ), .Z(n_13573));
	notech_inv i_21571(.A(\tab23[19] ), .Z(n_13574));
	notech_inv i_21572(.A(\tab23[20] ), .Z(n_13575));
	notech_inv i_21573(.A(\tab23[21] ), .Z(n_13576));
	notech_inv i_21574(.A(\tab23[22] ), .Z(n_13577));
	notech_inv i_21575(.A(\tab23[23] ), .Z(n_13578));
	notech_inv i_21576(.A(\tab23[24] ), .Z(n_13579));
	notech_inv i_21577(.A(\tab23[25] ), .Z(n_13580));
	notech_inv i_21578(.A(\tab23[26] ), .Z(n_13581));
	notech_inv i_21579(.A(\tab23[27] ), .Z(n_13582));
	notech_inv i_21580(.A(\tab23[28] ), .Z(n_13583));
	notech_inv i_21581(.A(\tab23[29] ), .Z(n_13584));
	notech_inv i_21582(.A(\tab24[10] ), .Z(n_13585));
	notech_inv i_21583(.A(\tab24[11] ), .Z(n_13586));
	notech_inv i_21584(.A(\tab24[12] ), .Z(n_13587));
	notech_inv i_21585(.A(\tab24[13] ), .Z(n_13588));
	notech_inv i_21586(.A(\tab24[14] ), .Z(n_13589));
	notech_inv i_21587(.A(\tab24[15] ), .Z(n_13590));
	notech_inv i_21588(.A(\tab24[16] ), .Z(n_13591));
	notech_inv i_21589(.A(\tab24[17] ), .Z(n_13592));
	notech_inv i_21590(.A(\tab24[18] ), .Z(n_13593));
	notech_inv i_21591(.A(\tab24[19] ), .Z(n_13594));
	notech_inv i_21592(.A(\tab24[20] ), .Z(n_13595));
	notech_inv i_21593(.A(\tab24[21] ), .Z(n_13596));
	notech_inv i_21594(.A(\tab24[22] ), .Z(n_13597));
	notech_inv i_21595(.A(\tab24[23] ), .Z(n_13598));
	notech_inv i_21596(.A(\tab24[24] ), .Z(n_13599));
	notech_inv i_21597(.A(\tab24[25] ), .Z(n_13600));
	notech_inv i_21598(.A(\tab24[26] ), .Z(n_13601));
	notech_inv i_21599(.A(\tab24[27] ), .Z(n_13602));
	notech_inv i_21600(.A(\tab24[28] ), .Z(n_13603));
	notech_inv i_21601(.A(\tab24[29] ), .Z(n_13604));
	notech_inv i_21602(.A(n_54069), .Z(n_13605));
	notech_inv i_21603(.A(\nnx_tab2[0] ), .Z(n_13606));
	notech_inv i_21604(.A(n_54075), .Z(n_13607));
	notech_inv i_21605(.A(\nnx_tab2[1] ), .Z(n_13608));
	notech_inv i_21606(.A(\nbus_14030[0] ), .Z(n_13609));
	notech_inv i_21607(.A(n_55457), .Z(n_13610));
	notech_inv i_21608(.A(\nx_tab2[0] ), .Z(n_13611));
	notech_inv i_21609(.A(n_55463), .Z(n_13612));
	notech_inv i_21610(.A(\nx_tab2[1] ), .Z(n_13613));
	notech_inv i_21611(.A(n_53241), .Z(n_13614));
	notech_inv i_21612(.A(n_54154), .Z(n_13615));
	notech_inv i_21613(.A(fsm[1]), .Z(n_13616));
	notech_inv i_21614(.A(fsm[2]), .Z(n_13617));
	notech_inv i_21615(.A(fsm[3]), .Z(n_13618));
	notech_inv i_21616(.A(n_54189), .Z(n_13619));
	notech_inv i_21617(.A(n_54195), .Z(n_13620));
	notech_inv i_21618(.A(n_54201), .Z(n_13621));
	notech_inv i_21619(.A(n_54207), .Z(n_13622));
	notech_inv i_21620(.A(n_54213), .Z(n_13623));
	notech_inv i_21621(.A(n_54219), .Z(n_13624));
	notech_inv i_21622(.A(n_54225), .Z(n_13625));
	notech_inv i_21623(.A(n_54231), .Z(n_13626));
	notech_inv i_21624(.A(n_54237), .Z(n_13627));
	notech_inv i_21625(.A(n_54243), .Z(n_13628));
	notech_inv i_21626(.A(req_miss), .Z(n_13629));
	notech_inv i_21627(.A(addr_miss[0]), .Z(n_13630));
	notech_inv i_21628(.A(addr_miss[1]), .Z(n_13631));
	notech_inv i_21629(.A(addr_miss[2]), .Z(n_13632));
	notech_inv i_21630(.A(addr_miss[3]), .Z(n_13633));
	notech_inv i_21631(.A(addr_miss[4]), .Z(n_13634));
	notech_inv i_21632(.A(addr_miss[5]), .Z(n_13635));
	notech_inv i_21633(.A(addr_miss[6]), .Z(n_13636));
	notech_inv i_21634(.A(addr_miss[7]), .Z(n_13637));
	notech_inv i_21635(.A(addr_miss[8]), .Z(n_13638));
	notech_inv i_21636(.A(addr_miss[9]), .Z(n_13639));
	notech_inv i_21637(.A(addr_miss[10]), .Z(n_13640));
	notech_inv i_21638(.A(addr_miss[11]), .Z(n_13641));
	notech_inv i_21639(.A(addr_miss[12]), .Z(n_13642));
	notech_inv i_21640(.A(wrA[12]), .Z(n_13643));
	notech_inv i_21641(.A(addr_miss[13]), .Z(n_13644));
	notech_inv i_21642(.A(wrA[13]), .Z(n_13645));
	notech_inv i_21643(.A(addr_miss[14]), .Z(n_13646));
	notech_inv i_21644(.A(wrA[14]), .Z(n_13647));
	notech_inv i_21645(.A(addr_miss[15]), .Z(n_13648));
	notech_inv i_21646(.A(wrA[15]), .Z(n_13649));
	notech_inv i_21647(.A(addr_miss[16]), .Z(n_13650));
	notech_inv i_21648(.A(wrA[16]), .Z(n_13651));
	notech_inv i_21649(.A(addr_miss[17]), .Z(n_13652));
	notech_inv i_21650(.A(wrA[17]), .Z(n_13653));
	notech_inv i_21651(.A(addr_miss[18]), .Z(n_13654));
	notech_inv i_21652(.A(wrA[18]), .Z(n_13655));
	notech_inv i_21653(.A(addr_miss[19]), .Z(n_13656));
	notech_inv i_21654(.A(wrA[19]), .Z(n_13657));
	notech_inv i_21655(.A(addr_miss[20]), .Z(n_13658));
	notech_inv i_21656(.A(wrA[20]), .Z(n_13659));
	notech_inv i_21657(.A(addr_miss[21]), .Z(n_13660));
	notech_inv i_21658(.A(wrA[21]), .Z(n_13661));
	notech_inv i_21659(.A(addr_miss[22]), .Z(n_13662));
	notech_inv i_21660(.A(wrA[22]), .Z(n_13663));
	notech_inv i_21661(.A(addr_miss[23]), .Z(n_13664));
	notech_inv i_21662(.A(wrA[23]), .Z(n_13665));
	notech_inv i_21663(.A(addr_miss[24]), .Z(n_13666));
	notech_inv i_21664(.A(wrA[24]), .Z(n_13667));
	notech_inv i_21665(.A(addr_miss[25]), .Z(n_13668));
	notech_inv i_21666(.A(wrA[25]), .Z(n_13669));
	notech_inv i_21667(.A(addr_miss[26]), .Z(n_13670));
	notech_inv i_21668(.A(wrA[26]), .Z(n_13671));
	notech_inv i_21669(.A(addr_miss[27]), .Z(n_13672));
	notech_inv i_21670(.A(wrA[27]), .Z(n_13673));
	notech_inv i_21671(.A(addr_miss[28]), .Z(n_13674));
	notech_inv i_21672(.A(wrA[28]), .Z(n_13675));
	notech_inv i_21673(.A(addr_miss[29]), .Z(n_13676));
	notech_inv i_21674(.A(wrA[29]), .Z(n_13677));
	notech_inv i_21675(.A(addr_miss[30]), .Z(n_13678));
	notech_inv i_21676(.A(wrA[30]), .Z(n_13679));
	notech_inv i_21677(.A(addr_miss[31]), .Z(n_13680));
	notech_inv i_21678(.A(wrA[31]), .Z(n_13681));
	notech_inv i_21679(.A(n_53845), .Z(n_13682));
	notech_inv i_21680(.A(n_53852), .Z(n_13683));
	notech_inv i_21681(.A(n_53859), .Z(n_13684));
	notech_inv i_21682(.A(n_53866), .Z(n_13685));
	notech_inv i_21683(.A(n_53873), .Z(n_13686));
	notech_inv i_21684(.A(n_53880), .Z(n_13687));
	notech_inv i_21685(.A(n_53887), .Z(n_13688));
	notech_inv i_21686(.A(n_53894), .Z(n_13689));
	notech_inv i_21687(.A(n_53901), .Z(n_13690));
	notech_inv i_21688(.A(n_53908), .Z(n_13691));
	notech_inv i_21689(.A(n_53915), .Z(n_13692));
	notech_inv i_21690(.A(n_53922), .Z(n_13693));
	notech_inv i_21691(.A(n_53929), .Z(n_13694));
	notech_inv i_21692(.A(n_53936), .Z(n_13695));
	notech_inv i_21693(.A(n_53943), .Z(n_13696));
	notech_inv i_21694(.A(n_53950), .Z(n_13697));
	notech_inv i_21695(.A(n_53957), .Z(n_13698));
	notech_inv i_21696(.A(n_53964), .Z(n_13699));
	notech_inv i_21697(.A(n_53971), .Z(n_13700));
	notech_inv i_21698(.A(n_53978), .Z(n_13701));
	notech_inv i_21700(.A(cr3[31]), .Z(n_13703));
	notech_inv i_21701(.A(cr3[30]), .Z(n_13704));
	notech_inv i_21702(.A(cr3[29]), .Z(n_13705));
	notech_inv i_21703(.A(cr3[28]), .Z(n_13706));
	notech_inv i_21704(.A(cr3[27]), .Z(n_13707));
	notech_inv i_21705(.A(cr3[26]), .Z(n_13708));
	notech_inv i_21706(.A(cr3[25]), .Z(n_13709));
	notech_inv i_21707(.A(cr3[24]), .Z(n_13710));
	notech_inv i_21708(.A(cr3[23]), .Z(n_13711));
	notech_inv i_21709(.A(cr3[22]), .Z(n_13712));
	notech_inv i_21710(.A(cr3[21]), .Z(n_13713));
	notech_inv i_21711(.A(cr3[20]), .Z(n_13714));
	notech_inv i_21712(.A(cr3[19]), .Z(n_13715));
	notech_inv i_21713(.A(cr3[18]), .Z(n_13716));
	notech_inv i_21714(.A(cr3[17]), .Z(n_13717));
	notech_inv i_21715(.A(cr3[16]), .Z(n_13718));
	notech_inv i_21716(.A(cr3[15]), .Z(n_13719));
	notech_inv i_21717(.A(cr3[14]), .Z(n_13720));
	notech_inv i_21718(.A(cr3[13]), .Z(n_13721));
	notech_inv i_21719(.A(cr3[12]), .Z(n_13722));
	notech_inv i_21720(.A(iDaddr[0]), .Z(n_13723));
	notech_inv i_21721(.A(iDaddr[1]), .Z(n_13724));
	notech_inv i_21722(.A(iDaddr[2]), .Z(n_13725));
	notech_inv i_21723(.A(iDaddr[3]), .Z(n_13726));
	notech_inv i_21724(.A(iDaddr[4]), .Z(n_13727));
	notech_inv i_21725(.A(iDaddr[5]), .Z(n_13728));
	notech_inv i_21726(.A(iDaddr[6]), .Z(n_13729));
	notech_inv i_21727(.A(iDaddr[7]), .Z(n_13730));
	notech_inv i_21728(.A(iDaddr[8]), .Z(n_13731));
	notech_inv i_21729(.A(iDaddr[9]), .Z(n_13732));
	notech_inv i_21730(.A(iDaddr[10]), .Z(n_13733));
	notech_inv i_21731(.A(iDaddr[11]), .Z(n_13734));
	notech_inv i_21732(.A(iDaddr[12]), .Z(n_13735));
	notech_inv i_21733(.A(iDaddr[13]), .Z(n_13736));
	notech_inv i_21734(.A(iDaddr[14]), .Z(n_13737));
	notech_inv i_21735(.A(iDaddr[15]), .Z(n_13738));
	notech_inv i_21736(.A(iDaddr[16]), .Z(n_13739));
	notech_inv i_21737(.A(iDaddr[17]), .Z(n_13740));
	notech_inv i_21738(.A(iDaddr[18]), .Z(n_13741));
	notech_inv i_21739(.A(iDaddr[19]), .Z(n_13742));
	notech_inv i_21740(.A(iDaddr[20]), .Z(n_13743));
	notech_inv i_21741(.A(iDaddr[21]), .Z(n_13744));
	notech_inv i_21742(.A(iDaddr[22]), .Z(n_13745));
	notech_inv i_21743(.A(iDaddr[23]), .Z(n_13746));
	notech_inv i_21744(.A(iDaddr[24]), .Z(n_13747));
	notech_inv i_21745(.A(iDaddr[25]), .Z(n_13748));
	notech_inv i_21746(.A(iDaddr[26]), .Z(n_13749));
	notech_inv i_21747(.A(iDaddr[27]), .Z(n_13750));
	notech_inv i_21748(.A(iDaddr[28]), .Z(n_13751));
	notech_inv i_21749(.A(iDaddr[29]), .Z(n_13752));
	notech_inv i_21750(.A(iDaddr[30]), .Z(n_13753));
	notech_inv i_21751(.A(iDaddr[31]), .Z(n_13754));
	notech_inv i_21752(.A(cs[1]), .Z(n_13755));
	notech_inv i_21753(.A(cr0[16]), .Z(n_13756));
	notech_inv i_21754(.A(n_977), .Z(n_13757));
	notech_inv i_21755(.A(\dir1_0[9] ), .Z(n_13758));
	notech_inv i_21756(.A(\dir1_0[8] ), .Z(n_13759));
	notech_inv i_21757(.A(\dir1_0[7] ), .Z(n_13760));
	notech_inv i_21758(.A(\dir1_0[6] ), .Z(n_13761));
	notech_inv i_21759(.A(\dir1_0[5] ), .Z(n_13762));
	notech_inv i_21760(.A(\dir1_0[4] ), .Z(n_13763));
	notech_inv i_21761(.A(\dir1_0[3] ), .Z(n_13764));
	notech_inv i_21762(.A(\dir1_0[2] ), .Z(n_13765));
	notech_inv i_21763(.A(\dir1_0[1] ), .Z(n_13766));
	notech_inv i_21764(.A(\dir1_0[0] ), .Z(n_13767));
	notech_inv i_21765(.A(\tab11_0[9] ), .Z(n_13768));
	notech_inv i_21766(.A(\tab11_0[8] ), .Z(n_13769));
	notech_inv i_21767(.A(\tab11_0[7] ), .Z(n_13770));
	notech_inv i_21768(.A(\tab11_0[6] ), .Z(n_13771));
	notech_inv i_21769(.A(\tab11_0[5] ), .Z(n_13772));
	notech_inv i_21770(.A(\tab11_0[4] ), .Z(n_13773));
	notech_inv i_21771(.A(\tab11_0[3] ), .Z(n_13774));
	notech_inv i_21772(.A(\tab11_0[2] ), .Z(n_13775));
	notech_inv i_21773(.A(\tab11_0[1] ), .Z(n_13776));
	notech_inv i_21774(.A(\tab11_0[0] ), .Z(n_13777));
	notech_inv i_21775(.A(oread_ack97032), .Z(oread_ack));
	notech_inv i_21776(.A(hit_tab12), .Z(n_13779));
	notech_inv i_21777(.A(hit_tab23), .Z(n_13780));
	notech_inv i_21778(.A(n_58609), .Z(n_13781));
	notech_inv i_21779(.A(n_58618), .Z(n_13782));
	notech_inv i_21780(.A(n_61604), .Z(n_13783));
	notech_inv i_21781(.A(iread_ack), .Z(n_13784));
	notech_inv i_21782(.A(flush_tlb), .Z(n_13785));
	cmp14_9 t11(.ina({\tab11[33] , \tab11[32] , UNCONNECTED_000, \tab11[30] 
		, \tab11[9] , \tab11[8] , \tab11[7] , \tab11[6] , \tab11[5] , \tab11[4] 
		, \tab11[3] , \tab11[2] , \tab11[1] , \tab11[0] }), .inb({
		UNCONNECTED_001, n_50997, UNCONNECTED_002, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab11), .out2(hit_add11));
	cmp14_8 t24(.ina({\tab24[33] , \tab24[32] , UNCONNECTED_003, \tab24[30] 
		, \tab24[9] , \tab24[8] , \tab24[7] , \tab24[6] , \tab24[5] , \tab24[4] 
		, \tab24[3] , \tab24[2] , \tab24[1] , \tab24[0] }), .inb({
		UNCONNECTED_004, n_50997, UNCONNECTED_005, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab24), .out2(hit_add24));
	cmp14_7 t23(.ina({\tab23[33] , \tab23[32] , UNCONNECTED_006, \tab23[30] 
		, \tab23[9] , \tab23[8] , \tab23[7] , \tab23[6] , \tab23[5] , \tab23[4] 
		, \tab23[3] , \tab23[2] , \tab23[1] , \tab23[0] }), .inb({
		UNCONNECTED_007, n_50997, UNCONNECTED_008, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab23), .out2(hit_add23));
	cmp14_6 t22(.ina({\tab22[33] , \tab22[32] , UNCONNECTED_009, \tab22[30] 
		, \tab22[9] , \tab22[8] , \tab22[7] , \tab22[6] , \tab22[5] , \tab22[4] 
		, \tab22[3] , \tab22[2] , \tab22[1] , \tab22[0] }), .inb({
		UNCONNECTED_010, n_50997, UNCONNECTED_011, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab22), .out2(hit_add22));
	cmp14_5 t21(.ina({\tab21[33] , \tab21[32] , UNCONNECTED_012, \tab21[30] 
		, \tab21[9] , \tab21[8] , \tab21[7] , \tab21[6] , \tab21[5] , \tab21[4] 
		, \tab21[3] , \tab21[2] , \tab21[1] , \tab21[0] }), .inb({
		UNCONNECTED_013, n_50997, UNCONNECTED_014, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab21), .out2(hit_add21));
	cmp14_4 t14(.ina({\tab14[33] , \tab14[32] , UNCONNECTED_015, \tab14[30] 
		, \tab14[9] , \tab14[8] , \tab14[7] , \tab14[6] , \tab14[5] , \tab14[4] 
		, \tab14[3] , \tab14[2] , \tab14[1] , \tab14[0] }), .inb({
		UNCONNECTED_016, n_50997, UNCONNECTED_017, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab14), .out2(hit_add14));
	cmp14_3 t13(.ina({\tab13[33] , \tab13[32] , UNCONNECTED_018, \tab13[30] 
		, \tab13[9] , \tab13[8] , \tab13[7] , \tab13[6] , \tab13[5] , \tab13[4] 
		, \tab13[3] , \tab13[2] , \tab13[1] , \tab13[0] }), .inb({
		UNCONNECTED_019, n_50997, UNCONNECTED_020, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab13), .out2(hit_add13));
	cmp14_2 t12(.ina({\tab12[33] , \tab12[32] , UNCONNECTED_021, \tab12[30] 
		, \tab12[9] , \tab12[8] , \tab12[7] , \tab12[6] , \tab12[5] , \tab12[4] 
		, \tab12[3] , \tab12[2] , \tab12[1] , \tab12[0] }), .inb({
		UNCONNECTED_022, n_50997, UNCONNECTED_023, iwrite_req, \tab11_0[9] 
		, \tab11_0[8] , \tab11_0[7] , \tab11_0[6] , \tab11_0[5] , \tab11_0[4] 
		, \tab11_0[3] , \tab11_0[2] , \tab11_0[1] , \tab11_0[0] }), .out
		(hit_tab12), .out2(hit_add12));
	cmp14_1 d2(.ina({\dir2[33] , UNCONNECTED_024, UNCONNECTED_025, 
		UNCONNECTED_026, \dir2[9] , \dir2[8] , \dir2[7] , \dir2[6] , \dir2[5] 
		, \dir2[4] , \dir2[3] , \dir2[2] , \dir2[1] , \dir2[0] }), .inb(
		{UNCONNECTED_027, UNCONNECTED_028, UNCONNECTED_029, 
		UNCONNECTED_030, \dir1_0[9] , \dir1_0[8] , \dir1_0[7] , \dir1_0[6] 
		, \dir1_0[5] , \dir1_0[4] , \dir1_0[3] , \dir1_0[2] , \dir1_0[1] 
		, \dir1_0[0] }), .out(hit_dir2));
	cmp14_0 d1(.ina({\dir1[33] , UNCONNECTED_031, UNCONNECTED_032, 
		UNCONNECTED_033, \dir1[9] , \dir1[8] , \dir1[7] , \dir1[6] , \dir1[5] 
		, \dir1[4] , \dir1[3] , \dir1[2] , \dir1[1] , \dir1[0] }), .inb(
		{UNCONNECTED_034, UNCONNECTED_035, UNCONNECTED_036, 
		UNCONNECTED_037, \dir1_0[9] , \dir1_0[8] , \dir1_0[7] , \dir1_0[6] 
		, \dir1_0[5] , \dir1_0[4] , \dir1_0[3] , \dir1_0[2] , \dir1_0[1] 
		, \dir1_0[0] }), .out(\hit_dir1[7] ));
	AWDP_INC_34 i_75623(.O0(fsm5_cnt_0), .fsm5_cnt(fsm5_cnt));
endmodule
module AWDP_INC_27(O0, fsm5_cnt);

	output [8:0] O0;
	input [8:0] fsm5_cnt;




	notech_ha2 i_8(.A(fsm5_cnt[8]), .B(n_86), .Z(O0[8]));
	notech_ha2 i_7(.A(fsm5_cnt[7]), .B(n_84), .Z(O0[7]), .CO(n_86));
	notech_ha2 i_6(.A(fsm5_cnt[6]), .B(n_82), .Z(O0[6]), .CO(n_84));
	notech_ha2 i_5(.A(fsm5_cnt[5]), .B(n_80), .Z(O0[5]), .CO(n_82));
	notech_ha2 i_4(.A(fsm5_cnt[4]), .B(n_78), .Z(O0[4]), .CO(n_80));
	notech_ha2 i_3(.A(fsm5_cnt[3]), .B(n_76), .Z(O0[3]), .CO(n_78));
	notech_ha2 i_2(.A(fsm5_cnt[2]), .B(n_74), .Z(O0[2]), .CO(n_76));
	notech_ha2 i_1(.A(fsm5_cnt[1]), .B(fsm5_cnt[0]), .Z(O0[1]), .CO(n_74));
	notech_inv i_0(.A(fsm5_cnt[0]), .Z(O0[0]));
endmodule
module cmp14_10(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_10(.A(inb[2]), .B(ina[2]), .Z(n_34));
	notech_xor2 i_9(.A(inb[4]), .B(ina[4]), .Z(n_33));
	notech_xor2 i_8(.A(inb[6]), .B(ina[6]), .Z(n_32));
	notech_xor2 i_6(.A(inb[3]), .B(ina[3]), .Z(n_31));
	notech_xor2 i_5(.A(inb[5]), .B(ina[5]), .Z(n_30));
	notech_xor2 i_4(.A(inb[7]), .B(ina[7]), .Z(n_29));
	notech_xor2 i_0(.A(inb[9]), .B(ina[9]), .Z(n_55));
	notech_xor2 i_1(.A(inb[8]), .B(ina[8]), .Z(n_56));
	notech_xor2 i_3(.A(inb[1]), .B(ina[1]), .Z(n_57));
	notech_xor2 i_7(.A(inb[0]), .B(ina[0]), .Z(n_58));
	notech_or4 i_38(.A(n_57), .B(n_56), .C(n_55), .D(ina[13]), .Z(n_61));
	notech_or4 i_37(.A(n_34), .B(n_31), .C(n_33), .D(n_30), .Z(n_66));
	notech_or4 i_39(.A(n_32), .B(n_29), .C(n_58), .D(n_66), .Z(n_67));
	notech_nor2 i_2(.A(n_67), .B(n_61), .Z(out));
endmodule
module cmp14_11(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_10(.A(inb[2]), .B(ina[2]), .Z(n_34));
	notech_xor2 i_9(.A(inb[4]), .B(ina[4]), .Z(n_33));
	notech_xor2 i_8(.A(inb[6]), .B(ina[6]), .Z(n_32));
	notech_xor2 i_6(.A(inb[3]), .B(ina[3]), .Z(n_31));
	notech_xor2 i_5(.A(inb[5]), .B(ina[5]), .Z(n_30));
	notech_xor2 i_4(.A(inb[7]), .B(ina[7]), .Z(n_29));
	notech_xor2 i_0(.A(inb[9]), .B(ina[9]), .Z(n_55));
	notech_xor2 i_1(.A(inb[8]), .B(ina[8]), .Z(n_56));
	notech_xor2 i_3(.A(inb[1]), .B(ina[1]), .Z(n_57));
	notech_xor2 i_7(.A(inb[0]), .B(ina[0]), .Z(n_58));
	notech_or4 i_38(.A(n_57), .B(n_56), .C(n_55), .D(ina[13]), .Z(n_61));
	notech_or4 i_37(.A(n_34), .B(n_31), .C(n_33), .D(n_30), .Z(n_66));
	notech_or4 i_39(.A(n_32), .B(n_29), .C(n_58), .D(n_66), .Z(n_67));
	notech_nor2 i_2(.A(n_67), .B(n_61), .Z(out));
endmodule
module cmp14_12(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out297002), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out297002));
	notech_inv i_9514(.A(out297002), .Z(out2));
endmodule
module cmp14_13(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out297001), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out297001));
	notech_inv i_9498(.A(out297001), .Z(out2));
endmodule
module cmp14_14(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out297000), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out297000));
	notech_inv i_9482(.A(out297000), .Z(out2));
endmodule
module cmp14_15(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out296999), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out296999));
	notech_inv i_9466(.A(out296999), .Z(out2));
endmodule
module cmp14_16(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out296998), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out296998));
	notech_inv i_9450(.A(out296998), .Z(out2));
endmodule
module cmp14_17(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out296997), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out296997));
	notech_inv i_9434(.A(out296997), .Z(out2));
endmodule
module cmp14_18(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out296996), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out296996));
	notech_inv i_9418(.A(out296996), .Z(out2));
endmodule
module cmp14_19(ina, inb, out, out2);

	input [13:0] ina;
	input [13:0] inb;
	output out;
	output out2;




	notech_xor2 i_25(.A(inb[5]), .B(ina[5]), .Z(n_59));
	notech_xor2 i_26(.A(inb[4]), .B(ina[4]), .Z(n_60));
	notech_xor2 i_27(.A(inb[3]), .B(ina[3]), .Z(n_62));
	notech_xor2 i_28(.A(inb[2]), .B(ina[2]), .Z(n_63));
	notech_or4 i_38(.A(n_63), .B(n_62), .C(n_60), .D(n_59), .Z(n_65));
	notech_xor2 i_29(.A(inb[1]), .B(ina[1]), .Z(n_66));
	notech_xor2 i_30(.A(inb[0]), .B(ina[0]), .Z(n_67));
	notech_xor2 i_21(.A(inb[9]), .B(ina[9]), .Z(n_69));
	notech_xor2 i_22(.A(inb[8]), .B(ina[8]), .Z(n_70));
	notech_xor2 i_23(.A(inb[7]), .B(ina[7]), .Z(n_72));
	notech_xor2 i_24(.A(inb[6]), .B(ina[6]), .Z(n_73));
	notech_or4 i_37(.A(n_73), .B(n_72), .C(n_70), .D(n_69), .Z(n_75));
	notech_nor2 i_2(.A(ina[13]), .B(out296995), .Z(out));
	notech_or4 i_32(.A(n_67), .B(n_66), .C(n_75), .D(n_65), .Z(out296995));
	notech_inv i_9402(.A(out296995), .Z(out2));
endmodule
module Itlb(clk, rstn, addr_phys, cr3, cr0, data_miss, iDaddr, pg_en, iwrite_data
		, owrite_data, iread_req, iread_ack, iwrite_req, iwrite_ack, iread_sz
		, oread_sz, oread_req, oread_ack, owrite_req, owrite_ack, pg_fault
		, wr_fault, cr2, flush_tlb, cs, pt_fault, busy_ram);

	input clk;
	input rstn;
	output [31:0] addr_phys;
	input [31:0] cr3;
	input [31:0] cr0;
	input [31:0] data_miss;
	input [31:0] iDaddr;
	input pg_en;
	input [31:0] iwrite_data;
	output [31:0] owrite_data;
	input iread_req;
	input iread_ack;
	input iwrite_req;
	input iwrite_ack;
	input [1:0] iread_sz;
	output [1:0] oread_sz;
	output oread_req;
	output oread_ack;
	output owrite_req;
	output owrite_ack;
	output pg_fault;
	output wr_fault;
	output [31:0] cr2;
	input flush_tlb;
	input [31:0] cs;
	output pt_fault;
	input busy_ram;

	wire [3:0] fsm;
	wire [31:0] iDaddr_f;
	wire [1:0] nx_dir;
	wire [8:0] fsm5_cnt_0;
	wire [8:0] fsm5_cnt;



	notech_inv i_15348(.A(n_61637), .Z(n_61691));
	notech_inv i_15347(.A(n_61637), .Z(n_61690));
	notech_inv i_15343(.A(n_61637), .Z(n_61686));
	notech_inv i_15339(.A(n_61637), .Z(n_61682));
	notech_inv i_15338(.A(n_61637), .Z(n_61681));
	notech_inv i_15334(.A(n_61637), .Z(n_61677));
	notech_inv i_15330(.A(n_61637), .Z(n_61673));
	notech_inv i_15329(.A(n_61637), .Z(n_61672));
	notech_inv i_15325(.A(n_61637), .Z(n_61668));
	notech_inv i_15320(.A(n_61637), .Z(n_61663));
	notech_inv i_15319(.A(n_61637), .Z(n_61662));
	notech_inv i_15315(.A(n_61637), .Z(n_61658));
	notech_inv i_15311(.A(n_61637), .Z(n_61654));
	notech_inv i_15310(.A(n_61637), .Z(n_61653));
	notech_inv i_15306(.A(n_61637), .Z(n_61649));
	notech_inv i_15302(.A(n_61637), .Z(n_61645));
	notech_inv i_15301(.A(n_61637), .Z(n_61644));
	notech_inv i_15297(.A(n_61637), .Z(n_61640));
	notech_inv i_15294(.A(clk), .Z(n_61637));
	notech_inv i_15292(.A(n_61609), .Z(n_61635));
	notech_inv i_15291(.A(n_61609), .Z(n_61634));
	notech_inv i_15287(.A(n_61609), .Z(n_61630));
	notech_inv i_15283(.A(n_61609), .Z(n_61626));
	notech_inv i_15282(.A(n_61609), .Z(n_61625));
	notech_inv i_15278(.A(n_61609), .Z(n_61621));
	notech_inv i_15274(.A(n_61609), .Z(n_61617));
	notech_inv i_15273(.A(n_61609), .Z(n_61616));
	notech_inv i_15269(.A(n_61609), .Z(n_61612));
	notech_inv i_15266(.A(clk), .Z(n_61609));
	notech_inv i_15254(.A(n_61589), .Z(n_61595));
	notech_inv i_15253(.A(n_61589), .Z(n_61594));
	notech_inv i_15249(.A(n_61589), .Z(n_61590));
	notech_inv i_15248(.A(pg_en), .Z(n_61589));
	notech_inv i_15244(.A(n_61578), .Z(n_61584));
	notech_inv i_15239(.A(n_61578), .Z(n_61579));
	notech_inv i_15238(.A(fsm[0]), .Z(n_61578));
	notech_inv i_15236(.A(n_61562), .Z(n_61575));
	notech_inv i_15234(.A(n_61562), .Z(n_61573));
	notech_inv i_15231(.A(n_61562), .Z(n_61570));
	notech_inv i_15229(.A(n_61562), .Z(n_61568));
	notech_inv i_15226(.A(n_61562), .Z(n_61565));
	notech_inv i_15224(.A(n_61562), .Z(n_61563));
	notech_inv i_15223(.A(n_551), .Z(n_61562));
	notech_inv i_15198(.A(n_61533), .Z(n_61534));
	notech_inv i_15197(.A(n_878), .Z(n_61533));
	notech_inv i_14821(.A(n_61465), .Z(n_61471));
	notech_inv i_14820(.A(n_61465), .Z(n_61470));
	notech_inv i_14816(.A(n_61465), .Z(n_61466));
	notech_inv i_14815(.A(n_886), .Z(n_61465));
	notech_inv i_14808(.A(n_61456), .Z(n_61457));
	notech_inv i_14807(.A(n_993), .Z(n_61456));
	notech_inv i_14800(.A(n_61447), .Z(n_61448));
	notech_inv i_14799(.A(n_9866), .Z(n_61447));
	notech_inv i_14322(.A(n_60909), .Z(n_60963));
	notech_inv i_14321(.A(n_60909), .Z(n_60962));
	notech_inv i_14317(.A(n_60909), .Z(n_60958));
	notech_inv i_14313(.A(n_60909), .Z(n_60954));
	notech_inv i_14312(.A(n_60909), .Z(n_60953));
	notech_inv i_14308(.A(n_60909), .Z(n_60949));
	notech_inv i_14304(.A(n_60909), .Z(n_60945));
	notech_inv i_14303(.A(n_60909), .Z(n_60944));
	notech_inv i_14299(.A(n_60909), .Z(n_60940));
	notech_inv i_14294(.A(n_60909), .Z(n_60935));
	notech_inv i_14293(.A(n_60909), .Z(n_60934));
	notech_inv i_14289(.A(n_60909), .Z(n_60930));
	notech_inv i_14285(.A(n_60909), .Z(n_60926));
	notech_inv i_14284(.A(n_60909), .Z(n_60925));
	notech_inv i_14280(.A(n_60909), .Z(n_60921));
	notech_inv i_14276(.A(n_60909), .Z(n_60917));
	notech_inv i_14275(.A(n_60909), .Z(n_60916));
	notech_inv i_14271(.A(n_60909), .Z(n_60912));
	notech_inv i_14268(.A(rstn), .Z(n_60909));
	notech_inv i_14266(.A(n_60881), .Z(n_60907));
	notech_inv i_14265(.A(n_60881), .Z(n_60906));
	notech_inv i_14261(.A(n_60881), .Z(n_60902));
	notech_inv i_14257(.A(n_60881), .Z(n_60898));
	notech_inv i_14256(.A(n_60881), .Z(n_60897));
	notech_inv i_14252(.A(n_60881), .Z(n_60893));
	notech_inv i_14248(.A(n_60881), .Z(n_60889));
	notech_inv i_14247(.A(n_60881), .Z(n_60888));
	notech_inv i_14243(.A(n_60881), .Z(n_60884));
	notech_inv i_14240(.A(rstn), .Z(n_60881));
	notech_inv i_14163(.A(n_60794), .Z(n_60795));
	notech_inv i_14162(.A(n_885), .Z(n_60794));
	notech_inv i_14155(.A(n_60785), .Z(n_60786));
	notech_inv i_14154(.A(n_890), .Z(n_60785));
	notech_inv i_13832(.A(n_60440), .Z(n_60441));
	notech_inv i_13831(.A(n_853), .Z(n_60440));
	notech_inv i_13828(.A(n_60431), .Z(n_60436));
	notech_inv i_13824(.A(n_60431), .Z(n_60432));
	notech_inv i_13823(.A(data_miss[0]), .Z(n_60431));
	notech_inv i_13609(.A(n_60112), .Z(n_60113));
	notech_inv i_13608(.A(\nbus_14493[0] ), .Z(n_60112));
	notech_inv i_13599(.A(n_60101), .Z(n_60102));
	notech_inv i_13598(.A(\nbus_14505[0] ), .Z(n_60101));
	notech_inv i_13589(.A(n_60090), .Z(n_60091));
	notech_inv i_13588(.A(\nbus_14494[0] ), .Z(n_60090));
	notech_inv i_13579(.A(n_60079), .Z(n_60080));
	notech_inv i_13578(.A(\nbus_14514[0] ), .Z(n_60079));
	notech_inv i_13569(.A(n_60068), .Z(n_60069));
	notech_inv i_13568(.A(\nbus_14501[0] ), .Z(n_60068));
	notech_inv i_13559(.A(n_60057), .Z(n_60058));
	notech_inv i_13558(.A(\nbus_14492[0] ), .Z(n_60057));
	notech_inv i_13549(.A(n_60046), .Z(n_60047));
	notech_inv i_13548(.A(\nbus_14517[0] ), .Z(n_60046));
	notech_inv i_13539(.A(n_60035), .Z(n_60036));
	notech_inv i_13538(.A(\nbus_14495[0] ), .Z(n_60035));
	notech_inv i_13529(.A(n_60024), .Z(n_60025));
	notech_inv i_13528(.A(\nbus_14502[0] ), .Z(n_60024));
	notech_inv i_13519(.A(n_60013), .Z(n_60014));
	notech_inv i_13518(.A(\nbus_14489[0] ), .Z(n_60013));
	notech_inv i_13490(.A(\nbus_14497[0] ), .Z(n_59983));
	notech_inv i_13485(.A(\nbus_14497[0] ), .Z(n_59977));
	notech_inv i_7757(.A(n_53567), .Z(n_53568));
	notech_inv i_7756(.A(n_808), .Z(n_53567));
	notech_ao3 i_68(.A(n_9985), .B(n_9956), .C(hit_adr24), .Z(n_492));
	notech_nor2 i_66(.A(hit_adr24), .B(\nx_tab2[0] ), .Z(n_490));
	notech_nor2 i_468(.A(hit_adr23), .B(n_490), .Z(n_489));
	notech_nor2 i_78(.A(hit_adr22), .B(n_489), .Z(n_487));
	notech_nand3 i_465(.A(n_60436), .B(n_875), .C(n_891), .Z(n_485));
	notech_or4 i_464(.A(n_899), .B(n_919), .C(n_10033), .D(\nx_tab1[1] ), .Z
		(n_484));
	notech_or4 i_463(.A(n_899), .B(n_919), .C(n_10035), .D(\nx_tab1[0] ), .Z
		(n_483));
	notech_or4 i_462(.A(n_899), .B(n_919), .C(n_10035), .D(n_10033), .Z(n_482
		));
	notech_xor2 i_79(.A(\nnx_tab1[1] ), .B(n_10028), .Z(n_478));
	notech_or4 i_73(.A(hit_adr13), .B(hit_adr14), .C(hit_adr12), .D(hit_adr11
		), .Z(n_476));
	notech_ao3 i_69(.A(n_10035), .B(n_10006), .C(hit_adr14), .Z(n_471));
	notech_nor2 i_67(.A(hit_adr14), .B(\nx_tab1[0] ), .Z(n_469));
	notech_nor2 i_452(.A(hit_adr13), .B(n_469), .Z(n_468));
	notech_nor2 i_80(.A(hit_adr12), .B(n_468), .Z(n_466));
	notech_or4 i_449(.A(n_899), .B(n_919), .C(\nx_tab1[1] ), .D(\nx_tab1[0] 
		), .Z(n_464));
	notech_and2 i_61(.A(fsm5_cnt[7]), .B(n_387), .Z(n_463));
	notech_or4 i_448(.A(fsm5_cnt[8]), .B(n_10181), .C(n_930), .D(n_463), .Z(n_462
		));
	notech_nor2 i_74(.A(n_463), .B(fsm5_cnt[8]), .Z(n_461));
	notech_nand2 i_445(.A(fsm[2]), .B(fsm[1]), .Z(n_459));
	notech_and3 i_51(.A(data_miss[5]), .B(iread_req), .C(n_60436), .Z(n_458)
		);
	notech_and2 i_82(.A(data_miss[5]), .B(n_60436), .Z(n_457));
	notech_ao3 i_85(.A(n_905), .B(iread_req), .C(busy_ram), .Z(n_454));
	notech_mux2 i_84(.S(fsm[3]), .A(n_459), .B(n_61584), .Z(n_453));
	notech_ao4 i_83(.A(n_61584), .B(n_889), .C(n_934), .D(n_896), .Z(n_452)
		);
	notech_or2 i_433(.A(iwrite_ack), .B(n_10058), .Z(n_450));
	notech_nor2 i_58(.A(data_miss[5]), .B(n_10124), .Z(n_449));
	notech_nand2 i_87(.A(n_948), .B(n_450), .Z(n_447));
	notech_mux2 i_86(.S(fsm[3]), .A(n_9867), .B(iwrite_ack), .Z(n_445));
	notech_nand3 i_427(.A(n_61584), .B(cr3[31]), .C(n_885), .Z(n_443));
	notech_nand3 i_424(.A(n_61584), .B(n_885), .C(cr3[30]), .Z(n_442));
	notech_nand3 i_421(.A(n_61584), .B(n_885), .C(cr3[29]), .Z(n_441));
	notech_nand3 i_418(.A(n_61584), .B(n_885), .C(cr3[28]), .Z(n_440));
	notech_nand3 i_415(.A(n_61584), .B(n_885), .C(cr3[27]), .Z(n_439));
	notech_nand3 i_412(.A(n_61584), .B(n_885), .C(cr3[26]), .Z(n_438));
	notech_nand3 i_409(.A(n_61584), .B(n_885), .C(cr3[25]), .Z(n_437));
	notech_nand3 i_406(.A(n_61584), .B(n_885), .C(cr3[24]), .Z(n_436));
	notech_nand3 i_403(.A(n_61584), .B(n_885), .C(cr3[23]), .Z(n_435));
	notech_nand3 i_400(.A(n_61584), .B(n_885), .C(cr3[22]), .Z(n_434));
	notech_nand3 i_397(.A(n_61584), .B(n_885), .C(cr3[21]), .Z(n_433));
	notech_nand3 i_394(.A(n_61584), .B(n_60795), .C(cr3[20]), .Z(n_432));
	notech_nand3 i_391(.A(n_61584), .B(n_60795), .C(cr3[19]), .Z(n_431));
	notech_nand3 i_388(.A(n_61584), .B(n_60795), .C(cr3[18]), .Z(n_430));
	notech_nand3 i_385(.A(n_61584), .B(n_60795), .C(cr3[17]), .Z(n_429));
	notech_nand3 i_382(.A(n_61584), .B(n_60795), .C(cr3[16]), .Z(n_428));
	notech_nand3 i_379(.A(n_61584), .B(n_60795), .C(cr3[15]), .Z(n_427));
	notech_nand3 i_376(.A(n_61579), .B(n_885), .C(cr3[14]), .Z(n_426));
	notech_nand3 i_373(.A(n_61579), .B(n_60795), .C(cr3[13]), .Z(n_425));
	notech_nand3 i_370(.A(n_61579), .B(n_60795), .C(cr3[12]), .Z(n_424));
	notech_nand3 i_344(.A(n_61594), .B(\wrA[2] ), .C(n_61471), .Z(n_400));
	notech_nor2 i_27(.A(n_972), .B(n_10181), .Z(n_399));
	notech_nand3 i_341(.A(n_61594), .B(n_61470), .C(\wrA[3] ), .Z(n_398));
	notech_nand3 i_338(.A(n_61595), .B(n_61471), .C(\wrA[4] ), .Z(n_397));
	notech_nand3 i_335(.A(n_61595), .B(n_61471), .C(\wrA[5] ), .Z(n_396));
	notech_nand3 i_332(.A(n_61595), .B(n_61471), .C(\wrA[6] ), .Z(n_395));
	notech_nand3 i_329(.A(n_61594), .B(n_61470), .C(\wrA[7] ), .Z(n_394));
	notech_nand3 i_326(.A(n_61594), .B(n_61470), .C(\wrA[8] ), .Z(n_393));
	notech_nand3 i_323(.A(n_61594), .B(n_61470), .C(\wrA[9] ), .Z(n_392));
	notech_nand3 i_320(.A(n_61594), .B(n_61470), .C(\wrA[10] ), .Z(n_391));
	notech_nand3 i_317(.A(n_61594), .B(n_61470), .C(\wrA[11] ), .Z(n_390));
	notech_nand2 i_81(.A(n_459), .B(n_10058), .Z(n_389));
	notech_nao3 i_21(.A(flush_tlb), .B(n_61595), .C(n_61573), .Z(n_388));
	notech_or2 i_60(.A(fsm5_cnt[6]), .B(n_386), .Z(n_387));
	notech_and3 i_52(.A(fsm5_cnt[4]), .B(fsm5_cnt[5]), .C(n_385), .Z(n_386)
		);
	notech_or2 i_48(.A(fsm5_cnt[2]), .B(fsm5_cnt[3]), .Z(n_385));
	notech_or4 i_72(.A(hit_adr23), .B(hit_adr24), .C(hit_adr22), .D(hit_adr21
		), .Z(n_497));
	notech_xor2 i_77(.A(\nnx_tab2[1] ), .B(n_9978), .Z(n_499));
	notech_nand3 i_478(.A(n_9868), .B(\nx_tab2[1] ), .C(\nx_tab2[0] ), .Z(n_503
		));
	notech_nand3 i_479(.A(n_9868), .B(\nx_tab2[1] ), .C(n_9983), .Z(n_504)
		);
	notech_nand3 i_480(.A(\nx_tab2[0] ), .B(n_9985), .C(n_9868), .Z(n_505)
		);
	notech_nand3 i_483(.A(n_9868), .B(n_9985), .C(n_9983), .Z(n_508));
	notech_or2 i_484(.A(n_876), .B(n_875), .Z(n_509));
	notech_or4 i_503(.A(n_61579), .B(n_875), .C(n_889), .D(n_887), .Z(n_528)
		);
	notech_or4 i_506(.A(nx_dir[0]), .B(nx_dir[1]), .C(n_887), .D(n_890), .Z(n_531
		));
	notech_or4 i_507(.A(n_61579), .B(n_889), .C(n_887), .D(n_60436), .Z(n_532
		));
	notech_or4 i_830012(.A(fsm[1]), .B(fsm[3]), .C(fsm[2]), .D(n_61579), .Z(n_551
		));
	notech_nand2 i_47(.A(n_61595), .B(n_555), .Z(n_553));
	notech_or4 i_528(.A(fsm[2]), .B(n_884), .C(n_61579), .D(n_883), .Z(n_555
		));
	notech_or4 i_75(.A(hit_tab12), .B(hit_tab11), .C(hit_tab13), .D(hit_tab14
		), .Z(n_557));
	notech_or4 i_76(.A(hit_tab22), .B(hit_tab21), .C(hit_tab24), .D(hit_tab23
		), .Z(n_559));
	notech_nao3 i_96(.A(n_973), .B(\addr_miss[31] ), .C(n_61471), .Z(n_564)
		);
	notech_nao3 i_93(.A(n_994), .B(\tab22[29] ), .C(n_993), .Z(n_567));
	notech_nand3 i_90(.A(n_9866), .B(n_986), .C(\tab13[29] ), .Z(n_570));
	notech_nao3 i_107(.A(n_973), .B(\addr_miss[30] ), .C(n_61471), .Z(n_575)
		);
	notech_nao3 i_104(.A(n_994), .B(\tab22[28] ), .C(n_993), .Z(n_578));
	notech_nand3 i_101(.A(n_9866), .B(n_986), .C(\tab13[28] ), .Z(n_581));
	notech_nao3 i_118(.A(n_973), .B(\addr_miss[29] ), .C(n_61471), .Z(n_586)
		);
	notech_nao3 i_115(.A(n_994), .B(\tab22[27] ), .C(n_993), .Z(n_589));
	notech_nand3 i_112(.A(n_9866), .B(n_986), .C(\tab13[27] ), .Z(n_592));
	notech_nao3 i_129(.A(n_973), .B(\addr_miss[28] ), .C(n_61471), .Z(n_597)
		);
	notech_nao3 i_126(.A(n_994), .B(\tab22[26] ), .C(n_993), .Z(n_600));
	notech_nand3 i_123(.A(n_9866), .B(n_986), .C(\tab13[26] ), .Z(n_603));
	notech_nao3 i_140(.A(n_973), .B(\addr_miss[27] ), .C(n_61471), .Z(n_608)
		);
	notech_nao3 i_137(.A(n_994), .B(\tab22[25] ), .C(n_993), .Z(n_611));
	notech_nand3 i_134(.A(n_9866), .B(n_986), .C(\tab13[25] ), .Z(n_614));
	notech_nao3 i_151(.A(n_973), .B(\addr_miss[26] ), .C(n_61471), .Z(n_619)
		);
	notech_nao3 i_148(.A(n_994), .B(\tab22[24] ), .C(n_993), .Z(n_622));
	notech_nand3 i_145(.A(n_9866), .B(n_986), .C(\tab13[24] ), .Z(n_625));
	notech_nao3 i_162(.A(n_973), .B(\addr_miss[25] ), .C(n_61471), .Z(n_630)
		);
	notech_nao3 i_159(.A(n_994), .B(\tab22[23] ), .C(n_993), .Z(n_633));
	notech_nand3 i_156(.A(n_9866), .B(n_986), .C(\tab13[23] ), .Z(n_636));
	notech_nao3 i_173(.A(n_973), .B(\addr_miss[24] ), .C(n_61471), .Z(n_641)
		);
	notech_nao3 i_170(.A(n_994), .B(\tab22[22] ), .C(n_993), .Z(n_644));
	notech_nand3 i_167(.A(n_9866), .B(n_986), .C(\tab13[22] ), .Z(n_647));
	notech_nao3 i_184(.A(n_973), .B(\addr_miss[23] ), .C(n_61471), .Z(n_652)
		);
	notech_nao3 i_181(.A(n_994), .B(\tab22[21] ), .C(n_993), .Z(n_655));
	notech_nand3 i_178(.A(n_9866), .B(n_986), .C(\tab13[21] ), .Z(n_658));
	notech_nao3 i_195(.A(n_973), .B(\addr_miss[22] ), .C(n_61471), .Z(n_663)
		);
	notech_nao3 i_192(.A(n_994), .B(\tab22[20] ), .C(n_993), .Z(n_666));
	notech_nand3 i_189(.A(n_9866), .B(n_986), .C(\tab13[20] ), .Z(n_669));
	notech_nao3 i_206(.A(n_973), .B(\addr_miss[21] ), .C(n_61470), .Z(n_674)
		);
	notech_nao3 i_203(.A(n_994), .B(\tab22[19] ), .C(n_993), .Z(n_677));
	notech_nand3 i_200(.A(n_9866), .B(n_986), .C(\tab13[19] ), .Z(n_680));
	notech_nao3 i_218(.A(n_973), .B(\addr_miss[20] ), .C(n_61466), .Z(n_685)
		);
	notech_nao3 i_214(.A(n_994), .B(\tab22[18] ), .C(n_61457), .Z(n_688));
	notech_nand3 i_211(.A(n_61448), .B(n_986), .C(\tab13[18] ), .Z(n_691));
	notech_nao3 i_235(.A(n_973), .B(\addr_miss[19] ), .C(n_61466), .Z(n_696)
		);
	notech_nao3 i_232(.A(n_994), .B(\tab22[17] ), .C(n_61457), .Z(n_699));
	notech_nand3 i_229(.A(n_61448), .B(n_986), .C(\tab13[17] ), .Z(n_702));
	notech_nao3 i_246(.A(n_973), .B(\addr_miss[18] ), .C(n_61466), .Z(n_707)
		);
	notech_nao3 i_243(.A(n_994), .B(\tab22[16] ), .C(n_61457), .Z(n_710));
	notech_nand3 i_240(.A(n_61448), .B(n_986), .C(\tab13[16] ), .Z(n_713));
	notech_nao3 i_257(.A(n_973), .B(\addr_miss[17] ), .C(n_61466), .Z(n_718)
		);
	notech_nao3 i_254(.A(n_994), .B(\tab22[15] ), .C(n_61457), .Z(n_721));
	notech_nand3 i_251(.A(n_61448), .B(n_986), .C(\tab13[15] ), .Z(n_724));
	notech_nao3 i_268(.A(n_973), .B(\addr_miss[16] ), .C(n_61466), .Z(n_729)
		);
	notech_nao3 i_265(.A(n_994), .B(\tab22[14] ), .C(n_61457), .Z(n_732));
	notech_nand3 i_262(.A(n_61448), .B(n_986), .C(\tab13[14] ), .Z(n_735));
	notech_nao3 i_279(.A(n_973), .B(\addr_miss[15] ), .C(n_61466), .Z(n_740)
		);
	notech_nao3 i_276(.A(n_994), .B(\tab22[13] ), .C(n_61457), .Z(n_743));
	notech_nand3 i_273(.A(n_61448), .B(n_986), .C(\tab13[13] ), .Z(n_746));
	notech_nao3 i_290(.A(n_973), .B(\addr_miss[14] ), .C(n_61466), .Z(n_751)
		);
	notech_nao3 i_287(.A(n_994), .B(\tab22[12] ), .C(n_61457), .Z(n_754));
	notech_nand3 i_284(.A(n_61448), .B(n_986), .C(\tab13[12] ), .Z(n_757));
	notech_nao3 i_301(.A(n_973), .B(\addr_miss[13] ), .C(n_61466), .Z(n_762)
		);
	notech_nao3 i_298(.A(n_994), .B(\tab22[11] ), .C(n_993), .Z(n_765));
	notech_nand3 i_295(.A(n_9866), .B(n_986), .C(\tab13[11] ), .Z(n_768));
	notech_nao3 i_312(.A(\addr_miss[12] ), .B(n_973), .C(n_61466), .Z(n_773)
		);
	notech_nao3 i_309(.A(\tab22[10] ), .B(n_994), .C(n_61457), .Z(n_776));
	notech_nand3 i_306(.A(n_61448), .B(\tab13[10] ), .C(n_986), .Z(n_779));
	notech_and2 i_8(.A(\wrD[7] ), .B(n_61466), .Z(owrite_data[7]));
	notech_and2 i_7(.A(\wrD[6] ), .B(n_61470), .Z(owrite_data[6]));
	notech_and2 i_6(.A(\wrD[5] ), .B(n_61470), .Z(owrite_data[5]));
	notech_and2 i_522313(.A(\wrD[4] ), .B(n_61470), .Z(owrite_data[4]));
	notech_and2 i_4(.A(\wrD[3] ), .B(n_61470), .Z(owrite_data[3]));
	notech_and2 i_3(.A(\wrD[2] ), .B(n_61470), .Z(owrite_data[2]));
	notech_and2 i_222312(.A(\wrD[1] ), .B(n_61466), .Z(owrite_data[1]));
	notech_and2 i_1(.A(\wrD[0] ), .B(n_61466), .Z(owrite_data[0]));
	notech_nao3 i_80343(.A(n_58573), .B(n_10124), .C(n_887), .Z(n_808));
	notech_or4 i_434(.A(n_854), .B(flush_tlb), .C(n_893), .D(n_906), .Z(n_851
		));
	notech_or4 i_435(.A(fsm[2]), .B(fsm[1]), .C(n_10181), .D(n_10058), .Z(n_852
		));
	notech_nand2 i_81549(.A(n_61595), .B(n_58550), .Z(n_853));
	notech_ao4 i_49(.A(hit_dir2), .B(\hit_dir1[7] ), .C(pg_fault), .D(n_9870
		), .Z(n_854));
	notech_or4 i_439(.A(fsm[1]), .B(fsm[3]), .C(fsm[2]), .D(n_454), .Z(n_855
		));
	notech_nao3 i_444(.A(n_10058), .B(n_9867), .C(iwrite_ack), .Z(n_858));
	notech_and2 i_44(.A(iwrite_ack), .B(n_389), .Z(n_861));
	notech_and2 i_79453(.A(n_58573), .B(n_10124), .Z(n_862));
	notech_ao3 i_79441(.A(fsm5_cnt_0[0]), .B(n_929), .C(n_884), .Z(n_863));
	notech_ao3 i_79442(.A(n_929), .B(fsm5_cnt_0[1]), .C(n_884), .Z(n_864));
	notech_ao3 i_79443(.A(n_929), .B(fsm5_cnt_0[2]), .C(n_884), .Z(n_865));
	notech_ao3 i_79444(.A(n_929), .B(fsm5_cnt_0[3]), .C(n_884), .Z(n_866));
	notech_ao3 i_79445(.A(n_929), .B(fsm5_cnt_0[4]), .C(n_884), .Z(n_867));
	notech_ao3 i_79446(.A(n_929), .B(fsm5_cnt_0[5]), .C(n_884), .Z(n_868));
	notech_ao3 i_79447(.A(n_929), .B(fsm5_cnt_0[6]), .C(n_884), .Z(n_869));
	notech_ao3 i_79448(.A(n_929), .B(fsm5_cnt_0[7]), .C(n_884), .Z(n_870));
	notech_ao3 i_79449(.A(n_929), .B(fsm5_cnt_0[8]), .C(n_884), .Z(n_871));
	notech_or4 i_81050(.A(n_906), .B(n_893), .C(n_904), .D(n_905), .Z(n_872)
		);
	notech_nor2 i_80097(.A(n_896), .B(n_10171), .Z(n_873));
	notech_ao3 i_79280(.A(n_60436), .B(\dir1_0[4] ), .C(n_890), .Z(n_874));
	notech_nor2 i_330010(.A(nx_dir[0]), .B(nx_dir[1]), .Z(n_875));
	notech_or4 i_81648(.A(n_61579), .B(n_889), .C(n_887), .D(n_10124), .Z(n_876
		));
	notech_and2 i_79197(.A(iread_ack), .B(n_553), .Z(oread_ack));
	notech_reg nx_dir_reg_0(.CP(n_61668), .D(n_7016), .CD(n_60940), .Q(nx_dir
		[0]));
	notech_mux2 i_9548(.S(n_876), .A(n_875), .B(nx_dir[0]), .Z(n_7016));
	notech_nand3 i_79169(.A(n_10058), .B(n_9867), .C(n_61595), .Z(n_878));
	notech_reg nx_dir_reg_1(.CP(n_61668), .D(n_7025), .CD(n_60940), .Q(nx_dir
		[1]));
	notech_and2 i_9558(.A(n_876), .B(nx_dir[1]), .Z(n_7025));
	notech_reg iDaddr_f_reg_0(.CP(n_61668), .D(n_7028), .CD(n_60940), .Q(iDaddr_f
		[0]));
	notech_mux2 i_9564(.S(n_61573), .A(iDaddr[0]), .B(iDaddr_f[0]), .Z(n_7028
		));
	notech_reg iDaddr_f_reg_1(.CP(n_61668), .D(n_7034), .CD(n_60940), .Q(iDaddr_f
		[1]));
	notech_mux2 i_9572(.S(n_61573), .A(iDaddr[1]), .B(iDaddr_f[1]), .Z(n_7034
		));
	notech_reg iDaddr_f_reg_2(.CP(n_61663), .D(n_7040), .CD(n_60935), .Q(iDaddr_f
		[2]));
	notech_mux2 i_9580(.S(n_61570), .A(iDaddr[2]), .B(iDaddr_f[2]), .Z(n_7040
		));
	notech_reg iDaddr_f_reg_3(.CP(n_61668), .D(n_7046), .CD(n_60940), .Q(iDaddr_f
		[3]));
	notech_mux2 i_9588(.S(n_61570), .A(iDaddr[3]), .B(iDaddr_f[3]), .Z(n_7046
		));
	notech_ao4 i_79026(.A(n_10183), .B(n_9948), .C(n_10180), .D(n_9945), .Z(n_883
		));
	notech_reg iDaddr_f_reg_4(.CP(n_61668), .D(n_7052), .CD(n_60940), .Q(iDaddr_f
		[4]));
	notech_mux2 i_9596(.S(n_61573), .A(iDaddr[4]), .B(iDaddr_f[4]), .Z(n_7052
		));
	notech_or2 i_30(.A(fsm[1]), .B(fsm[3]), .Z(n_884));
	notech_reg iDaddr_f_reg_5(.CP(n_61668), .D(n_7058), .CD(n_60940), .Q(iDaddr_f
		[5]));
	notech_mux2 i_9604(.S(n_61573), .A(iDaddr[5]), .B(iDaddr_f[5]), .Z(n_7058
		));
	notech_nor2 i_59(.A(fsm[2]), .B(n_884), .Z(n_885));
	notech_reg iDaddr_f_reg_6(.CP(n_61668), .D(n_7064), .CD(n_60940), .Q(iDaddr_f
		[6]));
	notech_mux2 i_9612(.S(n_61573), .A(iDaddr[6]), .B(iDaddr_f[6]), .Z(n_7064
		));
	notech_and3 i_20(.A(fsm[2]), .B(fsm[1]), .C(n_10058), .Z(n_886));
	notech_reg iDaddr_f_reg_7(.CP(n_61668), .D(n_7070), .CD(n_60940), .Q(iDaddr_f
		[7]));
	notech_mux2 i_9620(.S(n_61573), .A(iDaddr[7]), .B(iDaddr_f[7]), .Z(n_7070
		));
	notech_nand2 i_31(.A(iread_ack), .B(n_61595), .Z(n_887));
	notech_reg iDaddr_f_reg_8(.CP(n_61668), .D(n_7076), .CD(n_60940), .Q(iDaddr_f
		[8]));
	notech_mux2 i_9628(.S(n_61573), .A(iDaddr[8]), .B(iDaddr_f[8]), .Z(n_7076
		));
	notech_reg iDaddr_f_reg_9(.CP(n_61668), .D(n_7082), .CD(n_60940), .Q(iDaddr_f
		[9]));
	notech_mux2 i_9636(.S(n_61573), .A(iDaddr[9]), .B(iDaddr_f[9]), .Z(n_7082
		));
	notech_nao3 i_18(.A(fsm[1]), .B(n_10058), .C(fsm[2]), .Z(n_889));
	notech_reg iDaddr_f_reg_10(.CP(n_61668), .D(n_7088), .CD(n_60940), .Q(iDaddr_f
		[10]));
	notech_mux2 i_9644(.S(n_61570), .A(iDaddr[10]), .B(iDaddr_f[10]), .Z(n_7088
		));
	notech_nand2 i_32(.A(n_10057), .B(n_9869), .Z(n_890));
	notech_reg iDaddr_f_reg_11(.CP(n_61668), .D(n_7094), .CD(n_60940), .Q(iDaddr_f
		[11]));
	notech_mux2 i_9652(.S(n_61570), .A(iDaddr[11]), .B(iDaddr_f[11]), .Z(n_7094
		));
	notech_ao3 i_55(.A(iread_ack), .B(n_61595), .C(n_890), .Z(n_891));
	notech_reg iDaddr_f_reg_12(.CP(n_61663), .D(\tab11_0[0] ), .CD(n_60935),
		 .Q(iDaddr_f[12]));
	notech_reg iDaddr_f_reg_13(.CP(n_61663), .D(\tab11_0[1] ), .CD(n_60935),
		 .Q(iDaddr_f[13]));
	notech_or4 i_64(.A(fsm[2]), .B(n_884), .C(n_61579), .D(n_10181), .Z(n_893
		));
	notech_reg iDaddr_f_reg_14(.CP(n_61663), .D(\tab11_0[2] ), .CD(n_60935),
		 .Q(iDaddr_f[14]));
	notech_reg iDaddr_f_reg_15(.CP(n_61663), .D(\tab11_0[3] ), .CD(n_60935),
		 .Q(iDaddr_f[15]));
	notech_nand2 i_802(.A(fsm[2]), .B(n_10057), .Z(n_895));
	notech_reg iDaddr_f_reg_16(.CP(n_61663), .D(\tab11_0[4] ), .CD(n_60935),
		 .Q(iDaddr_f[16]));
	notech_or2 i_79145(.A(n_884), .B(n_895), .Z(n_896));
	notech_reg iDaddr_f_reg_17(.CP(n_61663), .D(\tab11_0[5] ), .CD(n_60935),
		 .Q(iDaddr_f[17]));
	notech_reg iDaddr_f_reg_18(.CP(n_61663), .D(\tab11_0[6] ), .CD(n_60935),
		 .Q(iDaddr_f[18]));
	notech_reg iDaddr_f_reg_19(.CP(n_61663), .D(\tab11_0[7] ), .CD(n_60935),
		 .Q(iDaddr_f[19]));
	notech_or4 i_10(.A(n_887), .B(n_884), .C(n_895), .D(n_10124), .Z(n_899)
		);
	notech_reg iDaddr_f_reg_20(.CP(n_61663), .D(\tab11_0[8] ), .CD(n_60935),
		 .Q(iDaddr_f[20]));
	notech_nand2 i_19(.A(hit_dir2), .B(n_10180), .Z(n_900));
	notech_reg iDaddr_f_reg_21(.CP(n_61663), .D(\tab11_0[9] ), .CD(n_60935),
		 .Q(iDaddr_f[21]));
	notech_or4 i_33(.A(n_896), .B(n_887), .C(n_900), .D(n_10124), .Z(n_901)
		);
	notech_reg iDaddr_f_reg_22(.CP(n_61663), .D(\dir1_0[0] ), .CD(n_60935), 
		.Q(iDaddr_f[22]));
	notech_reg iDaddr_f_reg_23(.CP(n_61663), .D(\dir1_0[1] ), .CD(n_60935), 
		.Q(iDaddr_f[23]));
	notech_reg iDaddr_f_reg_24(.CP(n_61663), .D(\dir1_0[2] ), .CD(n_60935), 
		.Q(iDaddr_f[24]));
	notech_nao3 i_798(.A(n_883), .B(n_10184), .C(flush_tlb), .Z(n_904));
	notech_reg iDaddr_f_reg_25(.CP(n_61663), .D(\dir1_0[3] ), .CD(n_60935), 
		.Q(iDaddr_f[25]));
	notech_and2 i_26(.A(n_10183), .B(n_10180), .Z(n_905));
	notech_reg iDaddr_f_reg_26(.CP(n_61663), .D(\dir1_0[4] ), .CD(n_60935), 
		.Q(iDaddr_f[26]));
	notech_or2 i_45(.A(busy_ram), .B(n_10182), .Z(n_906));
	notech_reg iDaddr_f_reg_27(.CP(n_61668), .D(\dir1_0[5] ), .CD(n_60940), 
		.Q(iDaddr_f[27]));
	notech_reg iDaddr_f_reg_28(.CP(n_61672), .D(\dir1_0[6] ), .CD(n_60944), 
		.Q(iDaddr_f[28]));
	notech_reg iDaddr_f_reg_29(.CP(n_61672), .D(\dir1_0[7] ), .CD(n_60944), 
		.Q(iDaddr_f[29]));
	notech_reg iDaddr_f_reg_30(.CP(n_61672), .D(\dir1_0[8] ), .CD(n_60944), 
		.Q(iDaddr_f[30]));
	notech_reg iDaddr_f_reg_31(.CP(n_61672), .D(\dir1_0[9] ), .CD(n_60944), 
		.Q(iDaddr_f[31]));
	notech_reg_set dir1_reg_0(.CP(n_61672), .D(n_7220), .SD(n_60944), .Q(\dir1[0] 
		));
	notech_mux2 i_9820(.S(\nbus_14492[0] ), .A(\dir1[0] ), .B(n_57419), .Z(n_7220
		));
	notech_nand2 i_79141(.A(n_61579), .B(n_9869), .Z(n_912));
	notech_reg_set dir1_reg_1(.CP(n_61672), .D(n_7226), .SD(n_60944), .Q(\dir1[1] 
		));
	notech_mux2 i_9828(.S(\nbus_14492[0] ), .A(\dir1[1] ), .B(n_57425), .Z(n_7226
		));
	notech_nao3 i_29(.A(n_61579), .B(n_61595), .C(n_889), .Z(n_913));
	notech_reg_set dir1_reg_2(.CP(n_61672), .D(n_7232), .SD(n_60944), .Q(\dir1[2] 
		));
	notech_mux2 i_9836(.S(\nbus_14492[0] ), .A(\dir1[2] ), .B(n_57431), .Z(n_7232
		));
	notech_reg_set dir1_reg_3(.CP(n_61673), .D(n_7238), .SD(n_60945), .Q(\dir1[3] 
		));
	notech_mux2 i_9844(.S(\nbus_14492[0] ), .A(\dir1[3] ), .B(n_57437), .Z(n_7238
		));
	notech_reg dir1_reg_4(.CP(n_61673), .D(n_7244), .CD(n_60945), .Q(\dir1[4] 
		));
	notech_mux2 i_9852(.S(\nbus_14492[0] ), .A(\dir1[4] ), .B(n_874), .Z(n_7244
		));
	notech_or2 i_53(.A(n_912), .B(hit_adr21), .Z(n_916));
	notech_reg_set dir1_reg_5(.CP(n_61673), .D(n_7250), .SD(n_60945), .Q(\dir1[5] 
		));
	notech_mux2 i_9860(.S(\nbus_14492[0] ), .A(\dir1[5] ), .B(n_57449), .Z(n_7250
		));
	notech_or2 i_789(.A(hit_adr22), .B(n_916), .Z(n_917));
	notech_reg_set dir1_reg_6(.CP(n_61673), .D(n_7256), .SD(n_60945), .Q(\dir1[6] 
		));
	notech_mux2 i_9868(.S(\nbus_14492[0] ), .A(\dir1[6] ), .B(n_57455), .Z(n_7256
		));
	notech_reg_set dir1_reg_7(.CP(n_61673), .D(n_7262), .SD(n_60945), .Q(\dir1[7] 
		));
	notech_mux2 i_9876(.S(\nbus_14492[0] ), .A(\dir1[7] ), .B(n_57461), .Z(n_7262
		));
	notech_nand2 i_17(.A(\hit_dir1[7] ), .B(n_10183), .Z(n_919));
	notech_reg_set dir1_reg_8(.CP(n_61673), .D(n_7268), .SD(n_60945), .Q(\dir1[8] 
		));
	notech_mux2 i_9884(.S(\nbus_14492[0] ), .A(\dir1[8] ), .B(n_57467), .Z(n_7268
		));
	notech_or4 i_34(.A(n_896), .B(n_887), .C(n_919), .D(n_10124), .Z(n_920)
		);
	notech_reg_set dir1_reg_9(.CP(n_61673), .D(n_7274), .SD(n_60945), .Q(\dir1[9] 
		));
	notech_mux2 i_9892(.S(\nbus_14492[0] ), .A(\dir1[9] ), .B(n_57473), .Z(n_7274
		));
	notech_reg_set dir1_reg_10(.CP(n_61672), .D(n_7280), .SD(n_60944), .Q(\dir1[10] 
		));
	notech_mux2 i_9900(.S(\nbus_14492[0] ), .A(\dir1[10] ), .B(n_57479), .Z(n_7280
		));
	notech_reg_set dir1_reg_11(.CP(n_61672), .D(n_7286), .SD(n_60944), .Q(\dir1[11] 
		));
	notech_mux2 i_9908(.S(\nbus_14492[0] ), .A(\dir1[11] ), .B(n_57485), .Z(n_7286
		));
	notech_reg_set dir1_reg_12(.CP(n_61672), .D(n_7292), .SD(n_60944), .Q(\dir1[12] 
		));
	notech_mux2 i_9916(.S(\nbus_14492[0] ), .A(\dir1[12] ), .B(n_57491), .Z(n_7292
		));
	notech_reg_set dir1_reg_13(.CP(n_61672), .D(n_7298), .SD(n_60944), .Q(\dir1[13] 
		));
	notech_mux2 i_9924(.S(\nbus_14492[0] ), .A(\dir1[13] ), .B(n_57497), .Z(n_7298
		));
	notech_reg_set dir1_reg_14(.CP(n_61668), .D(n_7304), .SD(n_60940), .Q(\dir1[14] 
		));
	notech_mux2 i_9932(.S(\nbus_14492[0] ), .A(\dir1[14] ), .B(n_57503), .Z(n_7304
		));
	notech_or2 i_54(.A(n_912), .B(hit_adr11), .Z(n_926));
	notech_reg_set dir1_reg_15(.CP(n_61668), .D(n_7310), .SD(n_60940), .Q(\dir1[15] 
		));
	notech_mux2 i_9940(.S(\nbus_14492[0] ), .A(\dir1[15] ), .B(n_57509), .Z(n_7310
		));
	notech_or2 i_784(.A(hit_adr12), .B(n_926), .Z(n_927));
	notech_reg_set dir1_reg_16(.CP(n_61668), .D(n_7316), .SD(n_60940), .Q(\dir1[16] 
		));
	notech_mux2 i_9948(.S(n_60058), .A(\dir1[16] ), .B(n_57515), .Z(n_7316)
		);
	notech_reg_set dir1_reg_17(.CP(n_61668), .D(n_7322), .SD(n_60940), .Q(\dir1[17] 
		));
	notech_mux2 i_9956(.S(n_60058), .A(\dir1[17] ), .B(n_57521), .Z(n_7322)
		);
	notech_and2 i_782(.A(fsm[2]), .B(n_61584), .Z(n_929));
	notech_reg_set dir1_reg_18(.CP(n_61672), .D(n_7328), .SD(n_60944), .Q(\dir1[18] 
		));
	notech_mux2 i_9964(.S(n_60058), .A(\dir1[18] ), .B(n_57527), .Z(n_7328)
		);
	notech_nao3 i_79148(.A(fsm[2]), .B(n_61579), .C(n_884), .Z(n_930));
	notech_reg_set dir1_reg_19(.CP(n_61672), .D(n_7334), .SD(n_60944), .Q(\dir1[19] 
		));
	notech_mux2 i_9972(.S(n_60058), .A(\dir1[19] ), .B(n_57533), .Z(n_7334)
		);
	notech_reg_set dir1_reg_20(.CP(n_61672), .D(n_7340), .SD(n_60944), .Q(\dir1[20] 
		));
	notech_mux2 i_9980(.S(n_60058), .A(\dir1[20] ), .B(n_57539), .Z(n_7340)
		);
	notech_nao3 i_35(.A(n_929), .B(n_61595), .C(n_884), .Z(n_932));
	notech_reg_set dir1_reg_21(.CP(n_61672), .D(n_7346), .SD(n_60944), .Q(\dir1[21] 
		));
	notech_mux2 i_9988(.S(n_60058), .A(\dir1[21] ), .B(n_57545), .Z(n_7346)
		);
	notech_reg_set dir1_reg_22(.CP(n_61672), .D(n_7352), .SD(n_60944), .Q(\dir1[22] 
		));
	notech_mux2 i_9996(.S(n_60058), .A(\dir1[22] ), .B(n_57551), .Z(n_7352)
		);
	notech_and2 i_28(.A(data_miss[5]), .B(iread_req), .Z(n_934));
	notech_reg_set dir1_reg_23(.CP(n_61672), .D(n_7358), .SD(n_60944), .Q(\dir1[23] 
		));
	notech_mux2 i_10004(.S(n_60058), .A(\dir1[23] ), .B(n_57557), .Z(n_7358)
		);
	notech_ao4 i_769(.A(n_896), .B(n_458), .C(n_889), .D(n_457), .Z(n_935)
		);
	notech_reg_set dir1_reg_24(.CP(n_61672), .D(n_7364), .SD(n_60944), .Q(\dir1[24] 
		));
	notech_mux2 i_10012(.S(n_60058), .A(\dir1[24] ), .B(n_57563), .Z(n_7364)
		);
	notech_reg_set dir1_reg_25(.CP(n_61654), .D(n_7370), .SD(n_60926), .Q(\dir1[25] 
		));
	notech_mux2 i_10020(.S(n_60058), .A(\dir1[25] ), .B(n_57569), .Z(n_7370)
		);
	notech_ao4 i_767(.A(n_453), .B(iwrite_ack), .C(n_452), .D(n_10124), .Z(n_937
		));
	notech_reg_set dir1_reg_26(.CP(n_61654), .D(n_7376), .SD(n_60926), .Q(\dir1[26] 
		));
	notech_mux2 i_10028(.S(n_60058), .A(\dir1[26] ), .B(n_57575), .Z(n_7376)
		);
	notech_nand2 i_79134(.A(n_61579), .B(n_60795), .Z(n_938));
	notech_reg_set dir1_reg_27(.CP(n_61658), .D(n_7382), .SD(n_60930), .Q(\dir1[27] 
		));
	notech_mux2 i_10036(.S(n_60058), .A(\dir1[27] ), .B(n_57581), .Z(n_7382)
		);
	notech_reg_set dir1_reg_28(.CP(n_61654), .D(n_7388), .SD(n_60926), .Q(\dir1[28] 
		));
	notech_mux2 i_10044(.S(n_60058), .A(\dir1[28] ), .B(n_57587), .Z(n_7388)
		);
	notech_reg_set dir1_reg_29(.CP(n_61654), .D(n_7394), .SD(n_60926), .Q(\dir1[29] 
		));
	notech_mux2 i_10052(.S(n_60058), .A(\dir1[29] ), .B(n_57593), .Z(n_7394)
		);
	notech_reg_set dir1_reg_33(.CP(n_61654), .D(n_7400), .SD(n_60926), .Q(\dir1[33] 
		));
	notech_mux2 i_10060(.S(n_60058), .A(\dir1[33] ), .B(n_57618), .Z(n_7400)
		);
	notech_reg_set dir2_reg_0(.CP(n_61654), .D(n_7406), .SD(n_60926), .Q(\dir2[0] 
		));
	notech_mux2 i_10068(.S(\nbus_14493[0] ), .A(\dir2[0] ), .B(n_57419), .Z(n_7406
		));
	notech_reg_set dir2_reg_1(.CP(n_61658), .D(n_7412), .SD(n_60930), .Q(\dir2[1] 
		));
	notech_mux2 i_10076(.S(\nbus_14493[0] ), .A(\dir2[1] ), .B(n_57425), .Z(n_7412
		));
	notech_reg_set dir2_reg_2(.CP(n_61658), .D(n_7418), .SD(n_60930), .Q(\dir2[2] 
		));
	notech_mux2 i_10084(.S(\nbus_14493[0] ), .A(\dir2[2] ), .B(n_57431), .Z(n_7418
		));
	notech_and3 i_760(.A(n_852), .B(n_851), .C(n_853), .Z(n_945));
	notech_reg_set dir2_reg_3(.CP(n_61658), .D(n_7424), .SD(n_60930), .Q(\dir2[3] 
		));
	notech_mux2 i_10092(.S(\nbus_14493[0] ), .A(\dir2[3] ), .B(n_57437), .Z(n_7424
		));
	notech_reg dir2_reg_4(.CP(n_61658), .D(n_7430), .CD(n_60930), .Q(\dir2[4] 
		));
	notech_mux2 i_10100(.S(\nbus_14493[0] ), .A(\dir2[4] ), .B(n_874), .Z(n_7430
		));
	notech_or2 i_757(.A(fsm[2]), .B(fsm[3]), .Z(n_947));
	notech_reg_set dir2_reg_5(.CP(n_61658), .D(n_7436), .SD(n_60930), .Q(\dir2[5] 
		));
	notech_mux2 i_10108(.S(\nbus_14493[0] ), .A(\dir2[5] ), .B(n_57449), .Z(n_7436
		));
	notech_ao4 i_756(.A(n_458), .B(n_884), .C(n_449), .D(n_947), .Z(n_948)
		);
	notech_reg_set dir2_reg_6(.CP(n_61658), .D(n_7442), .SD(n_60930), .Q(\dir2[6] 
		));
	notech_mux2 i_10116(.S(\nbus_14493[0] ), .A(\dir2[6] ), .B(n_57455), .Z(n_7442
		));
	notech_or2 i_15(.A(\hit_dir1[7] ), .B(n_912), .Z(n_949));
	notech_reg_set dir2_reg_7(.CP(n_61658), .D(n_7448), .SD(n_60930), .Q(\dir2[7] 
		));
	notech_mux2 i_10124(.S(\nbus_14493[0] ), .A(\dir2[7] ), .B(n_57461), .Z(n_7448
		));
	notech_nao3 i_11(.A(n_61579), .B(\hit_dir1[7] ), .C(n_889), .Z(n_950));
	notech_reg_set dir2_reg_8(.CP(n_61654), .D(n_7454), .SD(n_60926), .Q(\dir2[8] 
		));
	notech_mux2 i_10132(.S(\nbus_14493[0] ), .A(\dir2[8] ), .B(n_57467), .Z(n_7454
		));
	notech_ao4 i_755(.A(n_950), .B(n_9890), .C(n_949), .D(n_9910), .Z(n_951)
		);
	notech_reg_set dir2_reg_9(.CP(n_61654), .D(n_7460), .SD(n_60926), .Q(\dir2[9] 
		));
	notech_mux2 i_10140(.S(\nbus_14493[0] ), .A(\dir2[9] ), .B(n_57473), .Z(n_7460
		));
	notech_ao4 i_754(.A(n_950), .B(n_9889), .C(n_949), .D(n_9909), .Z(n_952)
		);
	notech_reg_set dir2_reg_10(.CP(n_61654), .D(n_7466), .SD(n_60926), .Q(\dir2[10] 
		));
	notech_mux2 i_10148(.S(\nbus_14493[0] ), .A(\dir2[10] ), .B(n_57479), .Z
		(n_7466));
	notech_ao4 i_753(.A(n_950), .B(n_9888), .C(n_949), .D(n_9908), .Z(n_953)
		);
	notech_reg_set dir2_reg_11(.CP(n_61654), .D(n_7472), .SD(n_60926), .Q(\dir2[11] 
		));
	notech_mux2 i_10156(.S(\nbus_14493[0] ), .A(\dir2[11] ), .B(n_57485), .Z
		(n_7472));
	notech_ao4 i_752(.A(n_950), .B(n_9887), .C(n_949), .D(n_9907), .Z(n_954)
		);
	notech_reg_set dir2_reg_12(.CP(n_61654), .D(n_7478), .SD(n_60926), .Q(\dir2[12] 
		));
	notech_mux2 i_10164(.S(\nbus_14493[0] ), .A(\dir2[12] ), .B(n_57491), .Z
		(n_7478));
	notech_ao4 i_751(.A(n_950), .B(n_9886), .C(n_949), .D(n_9906), .Z(n_955)
		);
	notech_reg_set dir2_reg_13(.CP(n_61653), .D(n_7484), .SD(n_60925), .Q(\dir2[13] 
		));
	notech_mux2 i_10172(.S(\nbus_14493[0] ), .A(\dir2[13] ), .B(n_57497), .Z
		(n_7484));
	notech_ao4 i_750(.A(n_950), .B(n_9885), .C(n_949), .D(n_9905), .Z(n_956)
		);
	notech_reg_set dir2_reg_14(.CP(n_61653), .D(n_7490), .SD(n_60925), .Q(\dir2[14] 
		));
	notech_mux2 i_10180(.S(\nbus_14493[0] ), .A(\dir2[14] ), .B(n_57503), .Z
		(n_7490));
	notech_ao4 i_749(.A(n_950), .B(n_9884), .C(n_949), .D(n_9904), .Z(n_957)
		);
	notech_reg_set dir2_reg_15(.CP(n_61653), .D(n_7496), .SD(n_60925), .Q(\dir2[15] 
		));
	notech_mux2 i_10188(.S(\nbus_14493[0] ), .A(\dir2[15] ), .B(n_57509), .Z
		(n_7496));
	notech_ao4 i_748(.A(n_950), .B(n_9883), .C(n_949), .D(n_9903), .Z(n_958)
		);
	notech_reg_set dir2_reg_16(.CP(n_61654), .D(n_7502), .SD(n_60926), .Q(\dir2[16] 
		));
	notech_mux2 i_10196(.S(n_60113), .A(\dir2[16] ), .B(n_57515), .Z(n_7502)
		);
	notech_ao4 i_747(.A(n_950), .B(n_9882), .C(n_949), .D(n_9902), .Z(n_959)
		);
	notech_reg_set dir2_reg_17(.CP(n_61654), .D(n_7508), .SD(n_60926), .Q(\dir2[17] 
		));
	notech_mux2 i_10204(.S(n_60113), .A(\dir2[17] ), .B(n_57521), .Z(n_7508)
		);
	notech_ao4 i_746(.A(n_950), .B(n_9881), .C(n_949), .D(n_9901), .Z(n_960)
		);
	notech_reg_set dir2_reg_18(.CP(n_61654), .D(n_7514), .SD(n_60926), .Q(\dir2[18] 
		));
	notech_mux2 i_10212(.S(n_60113), .A(\dir2[18] ), .B(n_57527), .Z(n_7514)
		);
	notech_ao4 i_745(.A(n_950), .B(n_9880), .C(n_949), .D(n_9900), .Z(n_961)
		);
	notech_reg_set dir2_reg_19(.CP(n_61654), .D(n_7520), .SD(n_60926), .Q(\dir2[19] 
		));
	notech_mux2 i_10220(.S(n_60113), .A(\dir2[19] ), .B(n_57533), .Z(n_7520)
		);
	notech_ao4 i_744(.A(n_950), .B(n_9879), .C(n_949), .D(n_9899), .Z(n_962)
		);
	notech_reg_set dir2_reg_20(.CP(n_61654), .D(n_7526), .SD(n_60926), .Q(\dir2[20] 
		));
	notech_mux2 i_10228(.S(n_60113), .A(\dir2[20] ), .B(n_57539), .Z(n_7526)
		);
	notech_ao4 i_743(.A(n_950), .B(n_9878), .C(n_949), .D(n_9898), .Z(n_963)
		);
	notech_reg_set dir2_reg_21(.CP(n_61654), .D(n_7532), .SD(n_60926), .Q(\dir2[21] 
		));
	notech_mux2 i_10236(.S(n_60113), .A(\dir2[21] ), .B(n_57545), .Z(n_7532)
		);
	notech_ao4 i_742(.A(n_950), .B(n_9877), .C(n_949), .D(n_9897), .Z(n_964)
		);
	notech_reg_set dir2_reg_22(.CP(n_61654), .D(n_7538), .SD(n_60926), .Q(\dir2[22] 
		));
	notech_mux2 i_10244(.S(n_60113), .A(\dir2[22] ), .B(n_57551), .Z(n_7538)
		);
	notech_ao4 i_741(.A(n_950), .B(n_9876), .C(n_949), .D(n_9896), .Z(n_965)
		);
	notech_reg_set dir2_reg_23(.CP(n_61658), .D(n_7544), .SD(n_60930), .Q(\dir2[23] 
		));
	notech_mux2 i_10252(.S(n_60113), .A(\dir2[23] ), .B(n_57557), .Z(n_7544)
		);
	notech_ao4 i_740(.A(n_950), .B(n_9875), .C(n_949), .D(n_9895), .Z(n_966)
		);
	notech_reg_set dir2_reg_24(.CP(n_61662), .D(n_7550), .SD(n_60934), .Q(\dir2[24] 
		));
	notech_mux2 i_10260(.S(n_60113), .A(\dir2[24] ), .B(n_57563), .Z(n_7550)
		);
	notech_ao4 i_739(.A(n_950), .B(n_9874), .C(n_949), .D(n_9894), .Z(n_967)
		);
	notech_reg_set dir2_reg_25(.CP(n_61662), .D(n_7556), .SD(n_60934), .Q(\dir2[25] 
		));
	notech_mux2 i_10268(.S(n_60113), .A(\dir2[25] ), .B(n_57569), .Z(n_7556)
		);
	notech_ao4 i_738(.A(n_950), .B(n_9873), .C(n_949), .D(n_9893), .Z(n_968)
		);
	notech_reg_set dir2_reg_26(.CP(n_61662), .D(n_7562), .SD(n_60934), .Q(\dir2[26] 
		));
	notech_mux2 i_10276(.S(n_60113), .A(\dir2[26] ), .B(n_57575), .Z(n_7562)
		);
	notech_ao4 i_737(.A(n_950), .B(n_9872), .C(n_949), .D(n_9892), .Z(n_969)
		);
	notech_reg_set dir2_reg_27(.CP(n_61662), .D(n_7568), .SD(n_60934), .Q(\dir2[27] 
		));
	notech_mux2 i_10284(.S(n_60113), .A(\dir2[27] ), .B(n_57581), .Z(n_7568)
		);
	notech_ao4 i_736(.A(n_950), .B(n_9871), .C(n_949), .D(n_9891), .Z(n_970)
		);
	notech_reg_set dir2_reg_28(.CP(n_61662), .D(n_7574), .SD(n_60934), .Q(\dir2[28] 
		));
	notech_mux2 i_10292(.S(n_60113), .A(\dir2[28] ), .B(n_57587), .Z(n_7574)
		);
	notech_reg_set dir2_reg_29(.CP(n_61662), .D(n_7580), .SD(n_60934), .Q(\dir2[29] 
		));
	notech_mux2 i_10300(.S(n_60113), .A(\dir2[29] ), .B(n_57593), .Z(n_7580)
		);
	notech_ao3 i_031203(.A(n_61595), .B(n_9870), .C(n_61466), .Z(n_972));
	notech_reg_set dir2_reg_33(.CP(n_61662), .D(n_7586), .SD(n_60934), .Q(\dir2[33] 
		));
	notech_mux2 i_10308(.S(n_60113), .A(\dir2[33] ), .B(n_57618), .Z(n_7586)
		);
	notech_and2 i_725(.A(n_61595), .B(n_883), .Z(n_973));
	notech_reg_set tab21_reg_0(.CP(n_61662), .D(n_7592), .SD(n_60934), .Q(\tab21[0] 
		));
	notech_mux2 i_10316(.S(\nbus_14494[0] ), .A(\tab21[0] ), .B(n_56940), .Z
		(n_7592));
	notech_nao3 i_9(.A(n_61595), .B(n_883), .C(n_61470), .Z(n_974));
	notech_reg_set tab21_reg_1(.CP(n_61663), .D(n_7598), .SD(n_60935), .Q(\tab21[1] 
		));
	notech_mux2 i_10324(.S(\nbus_14494[0] ), .A(\tab21[1] ), .B(n_56946), .Z
		(n_7598));
	notech_ao4 i_724(.A(n_974), .B(n_10069), .C(n_399), .D(n_10125), .Z(n_975
		));
	notech_reg_set tab21_reg_2(.CP(n_61663), .D(n_7604), .SD(n_60935), .Q(\tab21[2] 
		));
	notech_mux2 i_10332(.S(\nbus_14494[0] ), .A(\tab21[2] ), .B(n_56952), .Z
		(n_7604));
	notech_ao4 i_723(.A(n_974), .B(n_10070), .C(n_399), .D(n_10126), .Z(n_976
		));
	notech_reg_set tab21_reg_3(.CP(n_61662), .D(n_7610), .SD(n_60934), .Q(\tab21[3] 
		));
	notech_mux2 i_10340(.S(\nbus_14494[0] ), .A(\tab21[3] ), .B(n_56958), .Z
		(n_7610));
	notech_ao4 i_722(.A(n_974), .B(n_10071), .C(n_399), .D(n_10127), .Z(n_977
		));
	notech_reg tab21_reg_4(.CP(n_61662), .D(n_7616), .CD(n_60934), .Q(\tab21[4] 
		));
	notech_mux2 i_10348(.S(\nbus_14494[0] ), .A(\tab21[4] ), .B(n_873), .Z(n_7616
		));
	notech_ao4 i_721(.A(n_974), .B(n_10072), .C(n_399), .D(n_10128), .Z(n_978
		));
	notech_reg_set tab21_reg_5(.CP(n_61662), .D(n_7622), .SD(n_60934), .Q(\tab21[5] 
		));
	notech_mux2 i_10356(.S(\nbus_14494[0] ), .A(\tab21[5] ), .B(n_56970), .Z
		(n_7622));
	notech_ao4 i_720(.A(n_974), .B(n_10073), .C(n_399), .D(n_10129), .Z(n_979
		));
	notech_reg_set tab21_reg_6(.CP(n_61662), .D(n_7628), .SD(n_60934), .Q(\tab21[6] 
		));
	notech_mux2 i_10364(.S(\nbus_14494[0] ), .A(\tab21[6] ), .B(n_56976), .Z
		(n_7628));
	notech_ao4 i_719(.A(n_974), .B(n_10074), .C(n_399), .D(n_10130), .Z(n_980
		));
	notech_reg_set tab21_reg_7(.CP(n_61662), .D(n_7634), .SD(n_60934), .Q(\tab21[7] 
		));
	notech_mux2 i_10372(.S(\nbus_14494[0] ), .A(\tab21[7] ), .B(n_56982), .Z
		(n_7634));
	notech_ao4 i_718(.A(n_974), .B(n_10075), .C(n_399), .D(n_10131), .Z(n_981
		));
	notech_reg_set tab21_reg_8(.CP(n_61658), .D(n_7640), .SD(n_60930), .Q(\tab21[8] 
		));
	notech_mux2 i_10380(.S(\nbus_14494[0] ), .A(\tab21[8] ), .B(n_56988), .Z
		(n_7640));
	notech_ao4 i_717(.A(n_974), .B(n_10076), .C(n_399), .D(n_10132), .Z(n_982
		));
	notech_reg_set tab21_reg_9(.CP(n_61658), .D(n_7646), .SD(n_60930), .Q(\tab21[9] 
		));
	notech_mux2 i_10388(.S(\nbus_14494[0] ), .A(\tab21[9] ), .B(n_56994), .Z
		(n_7646));
	notech_ao4 i_716(.A(n_974), .B(n_10077), .C(n_399), .D(n_10133), .Z(n_983
		));
	notech_reg_set tab21_reg_10(.CP(n_61658), .D(n_7652), .SD(n_60930), .Q(\tab21[10] 
		));
	notech_mux2 i_10396(.S(\nbus_14494[0] ), .A(\tab21[10] ), .B(n_57000), .Z
		(n_7652));
	notech_ao4 i_715(.A(n_974), .B(n_10078), .C(n_399), .D(n_10134), .Z(n_984
		));
	notech_reg_set tab21_reg_11(.CP(n_61658), .D(n_7658), .SD(n_60930), .Q(\tab21[11] 
		));
	notech_mux2 i_10404(.S(\nbus_14494[0] ), .A(\tab21[11] ), .B(n_57006), .Z
		(n_7658));
	notech_nand2 i_63(.A(\hit_dir1[7] ), .B(n_972), .Z(n_985));
	notech_reg_set tab21_reg_12(.CP(n_61658), .D(n_7664), .SD(n_60930), .Q(\tab21[12] 
		));
	notech_mux2 i_10412(.S(\nbus_14494[0] ), .A(\tab21[12] ), .B(n_57012), .Z
		(n_7664));
	notech_ao3 i_713(.A(hit_tab13), .B(n_10179), .C(hit_tab11), .Z(n_986));
	notech_reg_set tab21_reg_13(.CP(n_61658), .D(n_7670), .SD(n_60930), .Q(\tab21[13] 
		));
	notech_mux2 i_10420(.S(\nbus_14494[0] ), .A(\tab21[13] ), .B(n_57018), .Z
		(n_7670));
	notech_reg_set tab21_reg_14(.CP(n_61658), .D(n_7676), .SD(n_60930), .Q(\tab21[14] 
		));
	notech_mux2 i_10428(.S(\nbus_14494[0] ), .A(\tab21[14] ), .B(n_57024), .Z
		(n_7676));
	notech_or4 i_25(.A(hit_tab12), .B(hit_tab11), .C(hit_tab13), .D(n_985), 
		.Z(n_988));
	notech_reg_set tab21_reg_15(.CP(n_61662), .D(n_7682), .SD(n_60934), .Q(\tab21[15] 
		));
	notech_mux2 i_10436(.S(\nbus_14494[0] ), .A(\tab21[15] ), .B(n_57030), .Z
		(n_7682));
	notech_reg_set tab21_reg_16(.CP(n_61662), .D(n_7688), .SD(n_60934), .Q(\tab21[16] 
		));
	notech_mux2 i_10444(.S(n_60091), .A(\tab21[16] ), .B(n_57036), .Z(n_7688
		));
	notech_nao3 i_24(.A(hit_tab12), .B(n_61448), .C(hit_tab11), .Z(n_990));
	notech_reg_set tab21_reg_17(.CP(n_61662), .D(n_7694), .SD(n_60934), .Q(\tab21[17] 
		));
	notech_mux2 i_10452(.S(n_60091), .A(\tab21[17] ), .B(n_57042), .Z(n_7694
		));
	notech_ao4 i_708(.A(n_9986), .B(n_990), .C(n_988), .D(n_10007), .Z(n_991
		));
	notech_reg_set tab21_reg_18(.CP(n_61662), .D(n_7700), .SD(n_60934), .Q(\tab21[18] 
		));
	notech_mux2 i_10460(.S(n_60091), .A(\tab21[18] ), .B(n_57048), .Z(n_7700
		));
	notech_reg_set tab21_reg_19(.CP(n_61658), .D(n_7706), .SD(n_60930), .Q(\tab21[19] 
		));
	notech_mux2 i_10468(.S(n_60091), .A(\tab21[19] ), .B(n_57054), .Z(n_7706
		));
	notech_or4 i_62(.A(n_61470), .B(\hit_dir1[7] ), .C(n_10181), .D(n_883), 
		.Z(n_993));
	notech_reg_set tab21_reg_20(.CP(n_61658), .D(n_7712), .SD(n_60930), .Q(\tab21[20] 
		));
	notech_mux2 i_10476(.S(n_60091), .A(\tab21[20] ), .B(n_57060), .Z(n_7712
		));
	notech_and2 i_711(.A(hit_tab22), .B(n_10177), .Z(n_994));
	notech_reg_set tab21_reg_21(.CP(n_61662), .D(n_7718), .SD(n_60934), .Q(\tab21[21] 
		));
	notech_mux2 i_10484(.S(n_60091), .A(\tab21[21] ), .B(n_57066), .Z(n_7718
		));
	notech_reg_set tab21_reg_22(.CP(n_61673), .D(n_7724), .SD(n_60945), .Q(\tab21[22] 
		));
	notech_mux2 i_10492(.S(n_60091), .A(\tab21[22] ), .B(n_57072), .Z(n_7724
		));
	notech_nand2 i_22(.A(hit_tab11), .B(n_61448), .Z(n_996));
	notech_reg_set tab21_reg_23(.CP(n_61686), .D(n_7730), .SD(n_60958), .Q(\tab21[23] 
		));
	notech_mux2 i_10500(.S(n_60091), .A(\tab21[23] ), .B(n_57078), .Z(n_7730
		));
	notech_reg_set tab21_reg_24(.CP(n_61686), .D(n_7736), .SD(n_60958), .Q(\tab21[24] 
		));
	notech_mux2 i_10508(.S(n_60091), .A(\tab21[24] ), .B(n_57084), .Z(n_7736
		));
	notech_or4 i_16(.A(hit_tab22), .B(hit_tab21), .C(n_61457), .D(n_10178), 
		.Z(n_998));
	notech_reg_set tab21_reg_25(.CP(n_61686), .D(n_7742), .SD(n_60958), .Q(\tab21[25] 
		));
	notech_mux2 i_10516(.S(n_60091), .A(\tab21[25] ), .B(n_57090), .Z(n_7742
		));
	notech_ao4 i_706(.A(n_998), .B(n_9933), .C(n_996), .D(n_10036), .Z(n_999
		));
	notech_reg_set tab21_reg_26(.CP(n_61686), .D(n_7748), .SD(n_60958), .Q(\tab21[26] 
		));
	notech_mux2 i_10524(.S(n_60091), .A(\tab21[26] ), .B(n_57096), .Z(n_7748
		));
	notech_reg_set tab21_reg_27(.CP(n_61686), .D(n_7754), .SD(n_60958), .Q(\tab21[27] 
		));
	notech_mux2 i_10532(.S(n_60091), .A(\tab21[27] ), .B(n_57102), .Z(n_7754
		));
	notech_and4 i_710(.A(n_999), .B(n_991), .C(n_776), .D(n_779), .Z(n_1001)
		);
	notech_reg_set tab21_reg_28(.CP(n_61686), .D(n_7760), .SD(n_60958), .Q(\tab21[28] 
		));
	notech_mux2 i_10540(.S(n_60091), .A(\tab21[28] ), .B(n_57108), .Z(n_7760
		));
	notech_nao3 i_13(.A(hit_tab21), .B(n_972), .C(\hit_dir1[7] ), .Z(n_1002)
		);
	notech_reg_set tab21_reg_29(.CP(n_61686), .D(n_7766), .SD(n_60958), .Q(\tab21[29] 
		));
	notech_mux2 i_10548(.S(n_60091), .A(\tab21[29] ), .B(n_57114), .Z(n_7766
		));
	notech_or4 i_12(.A(hit_tab22), .B(hit_tab21), .C(hit_tab23), .D(n_61457)
		, .Z(n_1003));
	notech_reg_set tab21_reg_33(.CP(n_61690), .D(n_7772), .SD(n_60962), .Q(\tab21[33] 
		));
	notech_mux2 i_10556(.S(n_60091), .A(\tab21[33] ), .B(n_57138), .Z(n_7772
		));
	notech_ao4 i_703(.A(n_1003), .B(n_9957), .C(n_1002), .D(n_9912), .Z(n_1004
		));
	notech_reg hit_adr21_reg(.CP(n_61690), .D(n_7778), .CD(n_60962), .Q(hit_adr21
		));
	notech_mux2 i_10564(.S(n_872), .A(hit_add21), .B(hit_adr21), .Z(n_7778)
		);
	notech_reg_set tab22_reg_0(.CP(n_61690), .D(n_7784), .SD(n_60962), .Q(\tab22[0] 
		));
	notech_mux2 i_10572(.S(\nbus_14505[0] ), .A(\tab22[0] ), .B(n_56940), .Z
		(n_7784));
	notech_ao4 i_702(.A(n_61590), .B(n_10135), .C(n_878), .D(n_10079), .Z(n_1006
		));
	notech_reg_set tab22_reg_1(.CP(n_61690), .D(n_7790), .SD(n_60962), .Q(\tab22[1] 
		));
	notech_mux2 i_10580(.S(\nbus_14505[0] ), .A(\tab22[1] ), .B(n_56946), .Z
		(n_7790));
	notech_reg_set tab22_reg_2(.CP(n_61686), .D(n_7796), .SD(n_60958), .Q(\tab22[2] 
		));
	notech_mux2 i_10588(.S(\nbus_14505[0] ), .A(\tab22[2] ), .B(n_56952), .Z
		(n_7796));
	notech_ao4 i_699(.A(n_990), .B(n_9987), .C(n_988), .D(n_10008), .Z(n_1008
		));
	notech_reg_set tab22_reg_3(.CP(n_61690), .D(n_7802), .SD(n_60962), .Q(\tab22[3] 
		));
	notech_mux2 i_10596(.S(\nbus_14505[0] ), .A(\tab22[3] ), .B(n_56958), .Z
		(n_7802));
	notech_reg tab22_reg_4(.CP(n_61690), .D(n_7808), .CD(n_60962), .Q(\tab22[4] 
		));
	notech_mux2 i_10604(.S(\nbus_14505[0] ), .A(\tab22[4] ), .B(n_873), .Z(n_7808
		));
	notech_ao4 i_697(.A(n_998), .B(n_9934), .C(n_996), .D(n_10037), .Z(n_1010
		));
	notech_reg_set tab22_reg_5(.CP(n_61686), .D(n_7814), .SD(n_60958), .Q(\tab22[5] 
		));
	notech_mux2 i_10612(.S(\nbus_14505[0] ), .A(\tab22[5] ), .B(n_56970), .Z
		(n_7814));
	notech_reg_set tab22_reg_6(.CP(n_61682), .D(n_7820), .SD(n_60954), .Q(\tab22[6] 
		));
	notech_mux2 i_10620(.S(\nbus_14505[0] ), .A(\tab22[6] ), .B(n_56976), .Z
		(n_7820));
	notech_and4 i_701(.A(n_1010), .B(n_1008), .C(n_765), .D(n_768), .Z(n_1012
		));
	notech_reg_set tab22_reg_7(.CP(n_61686), .D(n_7826), .SD(n_60958), .Q(\tab22[7] 
		));
	notech_mux2 i_10628(.S(\nbus_14505[0] ), .A(\tab22[7] ), .B(n_56982), .Z
		(n_7826));
	notech_ao4 i_694(.A(n_1003), .B(n_9958), .C(n_1002), .D(n_9913), .Z(n_1013
		));
	notech_reg_set tab22_reg_8(.CP(n_61686), .D(n_7832), .SD(n_60958), .Q(\tab22[8] 
		));
	notech_mux2 i_10636(.S(\nbus_14505[0] ), .A(\tab22[8] ), .B(n_56988), .Z
		(n_7832));
	notech_reg_set tab22_reg_9(.CP(n_61682), .D(n_7838), .SD(n_60954), .Q(\tab22[9] 
		));
	notech_mux2 i_10644(.S(\nbus_14505[0] ), .A(\tab22[9] ), .B(n_56994), .Z
		(n_7838));
	notech_ao4 i_693(.A(n_61590), .B(n_10136), .C(n_878), .D(n_10080), .Z(n_1015
		));
	notech_reg_set tab22_reg_10(.CP(n_61682), .D(n_7844), .SD(n_60954), .Q(\tab22[10] 
		));
	notech_mux2 i_10652(.S(\nbus_14505[0] ), .A(\tab22[10] ), .B(n_57000), .Z
		(n_7844));
	notech_reg_set tab22_reg_11(.CP(n_61682), .D(n_7850), .SD(n_60954), .Q(\tab22[11] 
		));
	notech_mux2 i_10660(.S(\nbus_14505[0] ), .A(\tab22[11] ), .B(n_57006), .Z
		(n_7850));
	notech_ao4 i_690(.A(n_990), .B(n_9988), .C(n_988), .D(n_10009), .Z(n_1017
		));
	notech_reg_set tab22_reg_12(.CP(n_61682), .D(n_7856), .SD(n_60954), .Q(\tab22[12] 
		));
	notech_mux2 i_10668(.S(\nbus_14505[0] ), .A(\tab22[12] ), .B(n_57012), .Z
		(n_7856));
	notech_reg_set tab22_reg_13(.CP(n_61686), .D(n_7862), .SD(n_60958), .Q(\tab22[13] 
		));
	notech_mux2 i_10676(.S(\nbus_14505[0] ), .A(\tab22[13] ), .B(n_57018), .Z
		(n_7862));
	notech_ao4 i_688(.A(n_998), .B(n_9935), .C(n_996), .D(n_10038), .Z(n_1019
		));
	notech_reg_set tab22_reg_14(.CP(n_61686), .D(n_7868), .SD(n_60958), .Q(\tab22[14] 
		));
	notech_mux2 i_10684(.S(\nbus_14505[0] ), .A(\tab22[14] ), .B(n_57024), .Z
		(n_7868));
	notech_reg_set tab22_reg_15(.CP(n_61686), .D(n_7874), .SD(n_60958), .Q(\tab22[15] 
		));
	notech_mux2 i_10692(.S(\nbus_14505[0] ), .A(\tab22[15] ), .B(n_57030), .Z
		(n_7874));
	notech_and4 i_692(.A(n_1019), .B(n_1017), .C(n_754), .D(n_757), .Z(n_1021
		));
	notech_reg_set tab22_reg_16(.CP(n_61686), .D(n_7880), .SD(n_60958), .Q(\tab22[16] 
		));
	notech_mux2 i_10700(.S(n_60102), .A(\tab22[16] ), .B(n_57036), .Z(n_7880
		));
	notech_ao4 i_685(.A(n_1003), .B(n_9959), .C(n_1002), .D(n_9914), .Z(n_1022
		));
	notech_reg_set tab22_reg_17(.CP(n_61686), .D(n_7886), .SD(n_60958), .Q(\tab22[17] 
		));
	notech_mux2 i_10708(.S(n_60102), .A(\tab22[17] ), .B(n_57042), .Z(n_7886
		));
	notech_reg_set tab22_reg_18(.CP(n_61686), .D(n_7892), .SD(n_60958), .Q(\tab22[18] 
		));
	notech_mux2 i_10716(.S(n_60102), .A(\tab22[18] ), .B(n_57048), .Z(n_7892
		));
	notech_ao4 i_684(.A(n_61590), .B(n_10137), .C(n_878), .D(n_10081), .Z(n_1024
		));
	notech_reg_set tab22_reg_19(.CP(n_61686), .D(n_7898), .SD(n_60958), .Q(\tab22[19] 
		));
	notech_mux2 i_10724(.S(n_60102), .A(\tab22[19] ), .B(n_57054), .Z(n_7898
		));
	notech_reg_set tab22_reg_20(.CP(n_61690), .D(n_7904), .SD(n_60962), .Q(\tab22[20] 
		));
	notech_mux2 i_10732(.S(n_60102), .A(\tab22[20] ), .B(n_57060), .Z(n_7904
		));
	notech_ao4 i_681(.A(n_990), .B(n_9989), .C(n_988), .D(n_10010), .Z(n_1026
		));
	notech_reg_set tab22_reg_21(.CP(n_61691), .D(n_7910), .SD(n_60963), .Q(\tab22[21] 
		));
	notech_mux2 i_10740(.S(n_60102), .A(\tab22[21] ), .B(n_57066), .Z(n_7910
		));
	notech_reg_set tab22_reg_22(.CP(n_61691), .D(n_7916), .SD(n_60963), .Q(\tab22[22] 
		));
	notech_mux2 i_10748(.S(n_60102), .A(\tab22[22] ), .B(n_57072), .Z(n_7916
		));
	notech_ao4 i_679(.A(n_998), .B(n_9936), .C(n_996), .D(n_10039), .Z(n_1028
		));
	notech_reg_set tab22_reg_23(.CP(n_61691), .D(n_7922), .SD(n_60963), .Q(\tab22[23] 
		));
	notech_mux2 i_10756(.S(n_60102), .A(\tab22[23] ), .B(n_57078), .Z(n_7922
		));
	notech_reg_set tab22_reg_24(.CP(n_61691), .D(n_7928), .SD(n_60963), .Q(\tab22[24] 
		));
	notech_mux2 i_10764(.S(n_60102), .A(\tab22[24] ), .B(n_57084), .Z(n_7928
		));
	notech_and4 i_683(.A(n_1028), .B(n_1026), .C(n_743), .D(n_746), .Z(n_1030
		));
	notech_reg_set tab22_reg_25(.CP(n_61691), .D(n_7934), .SD(n_60963), .Q(\tab22[25] 
		));
	notech_mux2 i_10772(.S(n_60102), .A(\tab22[25] ), .B(n_57090), .Z(n_7934
		));
	notech_ao4 i_676(.A(n_1003), .B(n_9960), .C(n_1002), .D(n_9915), .Z(n_1031
		));
	notech_reg_set tab22_reg_26(.CP(n_61691), .D(n_7940), .SD(n_60963), .Q(\tab22[26] 
		));
	notech_mux2 i_10780(.S(n_60102), .A(\tab22[26] ), .B(n_57096), .Z(n_7940
		));
	notech_reg_set tab22_reg_27(.CP(n_61691), .D(n_7946), .SD(n_60963), .Q(\tab22[27] 
		));
	notech_mux2 i_10788(.S(n_60102), .A(\tab22[27] ), .B(n_57102), .Z(n_7946
		));
	notech_ao4 i_675(.A(n_61590), .B(n_10138), .C(n_878), .D(n_10082), .Z(n_1033
		));
	notech_reg_set tab22_reg_28(.CP(n_61691), .D(n_7952), .SD(n_60963), .Q(\tab22[28] 
		));
	notech_mux2 i_10796(.S(n_60102), .A(\tab22[28] ), .B(n_57108), .Z(n_7952
		));
	notech_reg_set tab22_reg_29(.CP(n_61691), .D(n_7958), .SD(n_60963), .Q(\tab22[29] 
		));
	notech_mux2 i_10804(.S(n_60102), .A(\tab22[29] ), .B(n_57114), .Z(n_7958
		));
	notech_ao4 i_672(.A(n_990), .B(n_9990), .C(n_988), .D(n_10011), .Z(n_1035
		));
	notech_reg_set tab22_reg_33(.CP(n_61691), .D(n_7964), .SD(n_60963), .Q(\tab22[33] 
		));
	notech_mux2 i_10812(.S(n_60102), .A(\tab22[33] ), .B(n_57138), .Z(n_7964
		));
	notech_reg hit_adr22_reg(.CP(n_61691), .D(n_7970), .CD(n_60963), .Q(hit_adr22
		));
	notech_mux2 i_10820(.S(n_872), .A(hit_add22), .B(hit_adr22), .Z(n_7970)
		);
	notech_ao4 i_670(.A(n_998), .B(n_9937), .C(n_996), .D(n_10040), .Z(n_1037
		));
	notech_reg_set tab23_reg_0(.CP(n_61691), .D(n_7976), .SD(n_60963), .Q(\tab23[0] 
		));
	notech_mux2 i_10828(.S(\nbus_14501[0] ), .A(\tab23[0] ), .B(n_56940), .Z
		(n_7976));
	notech_reg_set tab23_reg_1(.CP(n_61691), .D(n_7982), .SD(n_60963), .Q(\tab23[1] 
		));
	notech_mux2 i_10836(.S(\nbus_14501[0] ), .A(\tab23[1] ), .B(n_56946), .Z
		(n_7982));
	notech_and4 i_674(.A(n_1037), .B(n_1035), .C(n_732), .D(n_735), .Z(n_1039
		));
	notech_reg_set tab23_reg_2(.CP(n_61691), .D(n_7988), .SD(n_60963), .Q(\tab23[2] 
		));
	notech_mux2 i_10844(.S(\nbus_14501[0] ), .A(\tab23[2] ), .B(n_56952), .Z
		(n_7988));
	notech_ao4 i_667(.A(n_1003), .B(n_9961), .C(n_1002), .D(n_9916), .Z(n_1040
		));
	notech_reg_set tab23_reg_3(.CP(n_61691), .D(n_7994), .SD(n_60963), .Q(\tab23[3] 
		));
	notech_mux2 i_10852(.S(\nbus_14501[0] ), .A(\tab23[3] ), .B(n_56958), .Z
		(n_7994));
	notech_reg tab23_reg_4(.CP(n_61690), .D(n_8000), .CD(n_60962), .Q(\tab23[4] 
		));
	notech_mux2 i_10860(.S(\nbus_14501[0] ), .A(\tab23[4] ), .B(n_873), .Z(n_8000
		));
	notech_ao4 i_666(.A(n_61590), .B(n_10139), .C(n_878), .D(n_10083), .Z(n_1042
		));
	notech_reg_set tab23_reg_5(.CP(n_61690), .D(n_8006), .SD(n_60962), .Q(\tab23[5] 
		));
	notech_mux2 i_10868(.S(\nbus_14501[0] ), .A(\tab23[5] ), .B(n_56970), .Z
		(n_8006));
	notech_reg_set tab23_reg_6(.CP(n_61690), .D(n_8012), .SD(n_60962), .Q(\tab23[6] 
		));
	notech_mux2 i_10876(.S(\nbus_14501[0] ), .A(\tab23[6] ), .B(n_56976), .Z
		(n_8012));
	notech_ao4 i_663(.A(n_990), .B(n_9991), .C(n_988), .D(n_10012), .Z(n_1044
		));
	notech_reg_set tab23_reg_7(.CP(n_61690), .D(n_8018), .SD(n_60962), .Q(\tab23[7] 
		));
	notech_mux2 i_10884(.S(\nbus_14501[0] ), .A(\tab23[7] ), .B(n_56982), .Z
		(n_8018));
	notech_reg_set tab23_reg_8(.CP(n_61690), .D(n_8024), .SD(n_60962), .Q(\tab23[8] 
		));
	notech_mux2 i_10892(.S(\nbus_14501[0] ), .A(\tab23[8] ), .B(n_56988), .Z
		(n_8024));
	notech_ao4 i_661(.A(n_998), .B(n_9938), .C(n_996), .D(n_10041), .Z(n_1046
		));
	notech_reg_set tab23_reg_9(.CP(n_61690), .D(n_8030), .SD(n_60962), .Q(\tab23[9] 
		));
	notech_mux2 i_10900(.S(\nbus_14501[0] ), .A(\tab23[9] ), .B(n_56994), .Z
		(n_8030));
	notech_reg_set tab23_reg_10(.CP(n_61690), .D(n_8036), .SD(n_60962), .Q(\tab23[10] 
		));
	notech_mux2 i_10908(.S(\nbus_14501[0] ), .A(\tab23[10] ), .B(n_57000), .Z
		(n_8036));
	notech_and4 i_665(.A(n_1046), .B(n_1044), .C(n_721), .D(n_724), .Z(n_1048
		));
	notech_reg_set tab23_reg_11(.CP(n_61691), .D(n_8042), .SD(n_60963), .Q(\tab23[11] 
		));
	notech_mux2 i_10916(.S(\nbus_14501[0] ), .A(\tab23[11] ), .B(n_57006), .Z
		(n_8042));
	notech_ao4 i_658(.A(n_1003), .B(n_9962), .C(n_1002), .D(n_9917), .Z(n_1049
		));
	notech_reg_set tab23_reg_12(.CP(n_61691), .D(n_8048), .SD(n_60963), .Q(\tab23[12] 
		));
	notech_mux2 i_10924(.S(\nbus_14501[0] ), .A(\tab23[12] ), .B(n_57012), .Z
		(n_8048));
	notech_reg_set tab23_reg_13(.CP(n_61691), .D(n_8054), .SD(n_60963), .Q(\tab23[13] 
		));
	notech_mux2 i_10932(.S(\nbus_14501[0] ), .A(\tab23[13] ), .B(n_57018), .Z
		(n_8054));
	notech_ao4 i_657(.A(n_61590), .B(n_10140), .C(n_878), .D(n_10084), .Z(n_1051
		));
	notech_reg_set tab23_reg_14(.CP(n_61690), .D(n_8060), .SD(n_60962), .Q(\tab23[14] 
		));
	notech_mux2 i_10940(.S(\nbus_14501[0] ), .A(\tab23[14] ), .B(n_57024), .Z
		(n_8060));
	notech_reg_set tab23_reg_15(.CP(n_61690), .D(n_8066), .SD(n_60962), .Q(\tab23[15] 
		));
	notech_mux2 i_10948(.S(\nbus_14501[0] ), .A(\tab23[15] ), .B(n_57030), .Z
		(n_8066));
	notech_ao4 i_654(.A(n_990), .B(n_9992), .C(n_988), .D(n_10013), .Z(n_1053
		));
	notech_reg_set tab23_reg_16(.CP(n_61690), .D(n_8072), .SD(n_60962), .Q(\tab23[16] 
		));
	notech_mux2 i_10956(.S(n_60069), .A(\tab23[16] ), .B(n_57036), .Z(n_8072
		));
	notech_reg_set tab23_reg_17(.CP(n_61690), .D(n_8078), .SD(n_60962), .Q(\tab23[17] 
		));
	notech_mux2 i_10964(.S(n_60069), .A(\tab23[17] ), .B(n_57042), .Z(n_8078
		));
	notech_ao4 i_652(.A(n_998), .B(n_9939), .C(n_996), .D(n_10042), .Z(n_1055
		));
	notech_reg_set tab23_reg_18(.CP(n_61677), .D(n_8084), .SD(n_60949), .Q(\tab23[18] 
		));
	notech_mux2 i_10972(.S(n_60069), .A(\tab23[18] ), .B(n_57048), .Z(n_8084
		));
	notech_reg_set tab23_reg_19(.CP(n_61677), .D(n_8090), .SD(n_60949), .Q(\tab23[19] 
		));
	notech_mux2 i_10980(.S(n_60069), .A(\tab23[19] ), .B(n_57054), .Z(n_8090
		));
	notech_and4 i_656(.A(n_1055), .B(n_1053), .C(n_710), .D(n_713), .Z(n_1057
		));
	notech_reg_set tab23_reg_20(.CP(n_61677), .D(n_8096), .SD(n_60949), .Q(\tab23[20] 
		));
	notech_mux2 i_10988(.S(n_60069), .A(\tab23[20] ), .B(n_57060), .Z(n_8096
		));
	notech_ao4 i_649(.A(n_1003), .B(n_9963), .C(n_1002), .D(n_9918), .Z(n_1058
		));
	notech_reg_set tab23_reg_21(.CP(n_61677), .D(n_8102), .SD(n_60949), .Q(\tab23[21] 
		));
	notech_mux2 i_10996(.S(n_60069), .A(\tab23[21] ), .B(n_57066), .Z(n_8102
		));
	notech_reg_set tab23_reg_22(.CP(n_61677), .D(n_8108), .SD(n_60949), .Q(\tab23[22] 
		));
	notech_mux2 i_11004(.S(n_60069), .A(\tab23[22] ), .B(n_57072), .Z(n_8108
		));
	notech_ao4 i_648(.A(n_61590), .B(n_10141), .C(n_878), .D(n_10085), .Z(n_1060
		));
	notech_reg_set tab23_reg_23(.CP(n_61677), .D(n_8114), .SD(n_60949), .Q(\tab23[23] 
		));
	notech_mux2 i_11012(.S(n_60069), .A(\tab23[23] ), .B(n_57078), .Z(n_8114
		));
	notech_reg_set tab23_reg_24(.CP(n_61677), .D(n_8120), .SD(n_60949), .Q(\tab23[24] 
		));
	notech_mux2 i_11020(.S(n_60069), .A(\tab23[24] ), .B(n_57084), .Z(n_8120
		));
	notech_ao4 i_645(.A(n_990), .B(n_9993), .C(n_988), .D(n_10014), .Z(n_1062
		));
	notech_reg_set tab23_reg_25(.CP(n_61677), .D(n_8126), .SD(n_60949), .Q(\tab23[25] 
		));
	notech_mux2 i_11028(.S(n_60069), .A(\tab23[25] ), .B(n_57090), .Z(n_8126
		));
	notech_reg_set tab23_reg_26(.CP(n_61677), .D(n_8132), .SD(n_60949), .Q(\tab23[26] 
		));
	notech_mux2 i_11036(.S(n_60069), .A(\tab23[26] ), .B(n_57096), .Z(n_8132
		));
	notech_ao4 i_643(.A(n_998), .B(n_9941), .C(n_996), .D(n_10043), .Z(n_1064
		));
	notech_reg_set tab23_reg_27(.CP(n_61681), .D(n_8138), .SD(n_60953), .Q(\tab23[27] 
		));
	notech_mux2 i_11044(.S(n_60069), .A(\tab23[27] ), .B(n_57102), .Z(n_8138
		));
	notech_reg_set tab23_reg_28(.CP(n_61677), .D(n_8144), .SD(n_60949), .Q(\tab23[28] 
		));
	notech_mux2 i_11052(.S(n_60069), .A(\tab23[28] ), .B(n_57108), .Z(n_8144
		));
	notech_and4 i_647(.A(n_1064), .B(n_1062), .C(n_699), .D(n_702), .Z(n_1066
		));
	notech_reg_set tab23_reg_29(.CP(n_61677), .D(n_8150), .SD(n_60949), .Q(\tab23[29] 
		));
	notech_mux2 i_11060(.S(n_60069), .A(\tab23[29] ), .B(n_57114), .Z(n_8150
		));
	notech_ao4 i_640(.A(n_1003), .B(n_9964), .C(n_1002), .D(n_9919), .Z(n_1067
		));
	notech_reg_set tab23_reg_33(.CP(n_61677), .D(n_8156), .SD(n_60949), .Q(\tab23[33] 
		));
	notech_mux2 i_11068(.S(n_60069), .A(\tab23[33] ), .B(n_57138), .Z(n_8156
		));
	notech_reg hit_adr23_reg(.CP(n_61677), .D(n_8162), .CD(n_60949), .Q(hit_adr23
		));
	notech_mux2 i_11076(.S(n_872), .A(hit_add23), .B(hit_adr23), .Z(n_8162)
		);
	notech_ao4 i_639(.A(n_61590), .B(n_10142), .C(n_878), .D(n_10086), .Z(n_1069
		));
	notech_reg_set tab24_reg_0(.CP(n_61677), .D(n_8168), .SD(n_60949), .Q(\tab24[0] 
		));
	notech_mux2 i_11084(.S(\nbus_14514[0] ), .A(\tab24[0] ), .B(n_56940), .Z
		(n_8168));
	notech_reg_set tab24_reg_1(.CP(n_61673), .D(n_8174), .SD(n_60945), .Q(\tab24[1] 
		));
	notech_mux2 i_11092(.S(\nbus_14514[0] ), .A(\tab24[1] ), .B(n_56946), .Z
		(n_8174));
	notech_ao4 i_636(.A(n_990), .B(n_9994), .C(n_988), .D(n_10015), .Z(n_1071
		));
	notech_reg_set tab24_reg_2(.CP(n_61673), .D(n_8180), .SD(n_60945), .Q(\tab24[2] 
		));
	notech_mux2 i_11100(.S(\nbus_14514[0] ), .A(\tab24[2] ), .B(n_56952), .Z
		(n_8180));
	notech_reg_set tab24_reg_3(.CP(n_61673), .D(n_8186), .SD(n_60945), .Q(\tab24[3] 
		));
	notech_mux2 i_11108(.S(\nbus_14514[0] ), .A(\tab24[3] ), .B(n_56958), .Z
		(n_8186));
	notech_ao4 i_634(.A(n_998), .B(n_9942), .C(n_996), .D(n_10044), .Z(n_1073
		));
	notech_reg tab24_reg_4(.CP(n_61673), .D(n_8192), .CD(n_60945), .Q(\tab24[4] 
		));
	notech_mux2 i_11116(.S(\nbus_14514[0] ), .A(\tab24[4] ), .B(n_873), .Z(n_8192
		));
	notech_reg_set tab24_reg_5(.CP(n_61673), .D(n_8198), .SD(n_60945), .Q(\tab24[5] 
		));
	notech_mux2 i_11124(.S(\nbus_14514[0] ), .A(\tab24[5] ), .B(n_56970), .Z
		(n_8198));
	notech_and4 i_638(.A(n_1073), .B(n_1071), .C(n_688), .D(n_691), .Z(n_1075
		));
	notech_reg_set tab24_reg_6(.CP(n_61673), .D(n_8204), .SD(n_60945), .Q(\tab24[6] 
		));
	notech_mux2 i_11132(.S(\nbus_14514[0] ), .A(\tab24[6] ), .B(n_56976), .Z
		(n_8204));
	notech_ao4 i_631(.A(n_1003), .B(n_9965), .C(n_1002), .D(n_9920), .Z(n_1076
		));
	notech_reg_set tab24_reg_7(.CP(n_61673), .D(n_8210), .SD(n_60945), .Q(\tab24[7] 
		));
	notech_mux2 i_11140(.S(\nbus_14514[0] ), .A(\tab24[7] ), .B(n_56982), .Z
		(n_8210));
	notech_reg_set tab24_reg_8(.CP(n_61677), .D(n_8216), .SD(n_60949), .Q(\tab24[8] 
		));
	notech_mux2 i_11148(.S(\nbus_14514[0] ), .A(\tab24[8] ), .B(n_56988), .Z
		(n_8216));
	notech_ao4 i_630(.A(n_61590), .B(n_10143), .C(n_878), .D(n_10087), .Z(n_1078
		));
	notech_reg_set tab24_reg_9(.CP(n_61677), .D(n_8222), .SD(n_60949), .Q(\tab24[9] 
		));
	notech_mux2 i_11156(.S(\nbus_14514[0] ), .A(\tab24[9] ), .B(n_56994), .Z
		(n_8222));
	notech_reg_set tab24_reg_10(.CP(n_61677), .D(n_8228), .SD(n_60949), .Q(\tab24[10] 
		));
	notech_mux2 i_11164(.S(\nbus_14514[0] ), .A(\tab24[10] ), .B(n_57000), .Z
		(n_8228));
	notech_ao4 i_627(.A(n_990), .B(n_9995), .C(n_988), .D(n_10016), .Z(n_1080
		));
	notech_reg_set tab24_reg_11(.CP(n_61677), .D(n_8234), .SD(n_60949), .Q(\tab24[11] 
		));
	notech_mux2 i_11172(.S(\nbus_14514[0] ), .A(\tab24[11] ), .B(n_57006), .Z
		(n_8234));
	notech_reg_set tab24_reg_12(.CP(n_61673), .D(n_8240), .SD(n_60945), .Q(\tab24[12] 
		));
	notech_mux2 i_11180(.S(\nbus_14514[0] ), .A(\tab24[12] ), .B(n_57012), .Z
		(n_8240));
	notech_ao4 i_625(.A(n_998), .B(n_9943), .C(n_996), .D(n_10045), .Z(n_1082
		));
	notech_reg_set tab24_reg_13(.CP(n_61673), .D(n_8246), .SD(n_60945), .Q(\tab24[13] 
		));
	notech_mux2 i_11188(.S(\nbus_14514[0] ), .A(\tab24[13] ), .B(n_57018), .Z
		(n_8246));
	notech_reg_set tab24_reg_14(.CP(n_61673), .D(n_8252), .SD(n_60945), .Q(\tab24[14] 
		));
	notech_mux2 i_11196(.S(\nbus_14514[0] ), .A(\tab24[14] ), .B(n_57024), .Z
		(n_8252));
	notech_and4 i_629(.A(n_1082), .B(n_1080), .C(n_677), .D(n_680), .Z(n_1084
		));
	notech_reg_set tab24_reg_15(.CP(n_61681), .D(n_8258), .SD(n_60953), .Q(\tab24[15] 
		));
	notech_mux2 i_11204(.S(\nbus_14514[0] ), .A(\tab24[15] ), .B(n_57030), .Z
		(n_8258));
	notech_ao4 i_622(.A(n_1003), .B(n_9966), .C(n_1002), .D(n_9921), .Z(n_1085
		));
	notech_reg_set tab24_reg_16(.CP(n_61682), .D(n_8264), .SD(n_60954), .Q(\tab24[16] 
		));
	notech_mux2 i_11212(.S(n_60080), .A(\tab24[16] ), .B(n_57036), .Z(n_8264
		));
	notech_reg_set tab24_reg_17(.CP(n_61682), .D(n_8270), .SD(n_60954), .Q(\tab24[17] 
		));
	notech_mux2 i_11220(.S(n_60080), .A(\tab24[17] ), .B(n_57042), .Z(n_8270
		));
	notech_ao4 i_621(.A(n_61590), .B(n_10144), .C(n_878), .D(n_10088), .Z(n_1087
		));
	notech_reg_set tab24_reg_18(.CP(n_61682), .D(n_8276), .SD(n_60954), .Q(\tab24[18] 
		));
	notech_mux2 i_11228(.S(n_60080), .A(\tab24[18] ), .B(n_57048), .Z(n_8276
		));
	notech_reg_set tab24_reg_19(.CP(n_61682), .D(n_8282), .SD(n_60954), .Q(\tab24[19] 
		));
	notech_mux2 i_11236(.S(n_60080), .A(\tab24[19] ), .B(n_57054), .Z(n_8282
		));
	notech_ao4 i_618(.A(n_990), .B(n_9996), .C(n_988), .D(n_10017), .Z(n_1089
		));
	notech_reg_set tab24_reg_20(.CP(n_61681), .D(n_8288), .SD(n_60953), .Q(\tab24[20] 
		));
	notech_mux2 i_11244(.S(n_60080), .A(\tab24[20] ), .B(n_57060), .Z(n_8288
		));
	notech_reg_set tab24_reg_21(.CP(n_61682), .D(n_8294), .SD(n_60954), .Q(\tab24[21] 
		));
	notech_mux2 i_11252(.S(n_60080), .A(\tab24[21] ), .B(n_57066), .Z(n_8294
		));
	notech_ao4 i_616(.A(n_998), .B(n_9944), .C(n_996), .D(n_10046), .Z(n_1091
		));
	notech_reg_set tab24_reg_22(.CP(n_61682), .D(n_8300), .SD(n_60954), .Q(\tab24[22] 
		));
	notech_mux2 i_11260(.S(n_60080), .A(\tab24[22] ), .B(n_57072), .Z(n_8300
		));
	notech_reg_set tab24_reg_23(.CP(n_61682), .D(n_8306), .SD(n_60954), .Q(\tab24[23] 
		));
	notech_mux2 i_11268(.S(n_60080), .A(\tab24[23] ), .B(n_57078), .Z(n_8306
		));
	notech_and4 i_620(.A(n_1091), .B(n_1089), .C(n_666), .D(n_669), .Z(n_1093
		));
	notech_reg_set tab24_reg_24(.CP(n_61682), .D(n_8312), .SD(n_60954), .Q(\tab24[24] 
		));
	notech_mux2 i_11276(.S(n_60080), .A(\tab24[24] ), .B(n_57084), .Z(n_8312
		));
	notech_ao4 i_613(.A(n_1003), .B(n_9967), .C(n_1002), .D(n_9922), .Z(n_1094
		));
	notech_reg_set tab24_reg_25(.CP(n_61682), .D(n_8318), .SD(n_60954), .Q(\tab24[25] 
		));
	notech_mux2 i_11284(.S(n_60080), .A(\tab24[25] ), .B(n_57090), .Z(n_8318
		));
	notech_reg_set tab24_reg_26(.CP(n_61682), .D(n_8324), .SD(n_60954), .Q(\tab24[26] 
		));
	notech_mux2 i_11292(.S(n_60080), .A(\tab24[26] ), .B(n_57096), .Z(n_8324
		));
	notech_ao4 i_612(.A(n_61590), .B(n_10145), .C(n_878), .D(n_10089), .Z(n_1096
		));
	notech_reg_set tab24_reg_27(.CP(n_61682), .D(n_8330), .SD(n_60954), .Q(\tab24[27] 
		));
	notech_mux2 i_11300(.S(n_60080), .A(\tab24[27] ), .B(n_57102), .Z(n_8330
		));
	notech_reg_set tab24_reg_28(.CP(n_61682), .D(n_8336), .SD(n_60954), .Q(\tab24[28] 
		));
	notech_mux2 i_11308(.S(n_60080), .A(\tab24[28] ), .B(n_57108), .Z(n_8336
		));
	notech_ao4 i_609(.A(n_990), .B(n_9997), .C(n_988), .D(n_10018), .Z(n_1098
		));
	notech_reg_set tab24_reg_29(.CP(n_61682), .D(n_8342), .SD(n_60954), .Q(\tab24[29] 
		));
	notech_mux2 i_11316(.S(n_60080), .A(\tab24[29] ), .B(n_57114), .Z(n_8342
		));
	notech_reg_set tab24_reg_33(.CP(n_61681), .D(n_8348), .SD(n_60953), .Q(\tab24[33] 
		));
	notech_mux2 i_11324(.S(n_60080), .A(\tab24[33] ), .B(n_57138), .Z(n_8348
		));
	notech_ao4 i_607(.A(n_998), .B(n_9946), .C(n_996), .D(n_10047), .Z(n_1100
		));
	notech_reg_set nnx_tab2_reg_0(.CP(n_61681), .D(n_8354), .SD(n_60953), .Q
		(\nnx_tab2[0] ));
	notech_mux2 i_11332(.S(n_9981), .A(\nnx_tab2[0] ), .B(n_9977), .Z(n_8354
		));
	notech_reg nnx_tab2_reg_1(.CP(n_61681), .D(n_8360), .CD(n_60953), .Q(\nnx_tab2[1] 
		));
	notech_mux2 i_11340(.S(n_9981), .A(\nnx_tab2[1] ), .B(n_9979), .Z(n_8360
		));
	notech_and4 i_611(.A(n_1100), .B(n_1098), .C(n_655), .D(n_658), .Z(n_1102
		));
	notech_reg hit_adr24_reg(.CP(n_61681), .D(n_8366), .CD(n_60953), .Q(hit_adr24
		));
	notech_mux2 i_11348(.S(n_872), .A(hit_add24), .B(hit_adr24), .Z(n_8366)
		);
	notech_ao4 i_604(.A(n_1003), .B(n_9968), .C(n_1002), .D(n_9923), .Z(n_1103
		));
	notech_reg nx_tab2_reg_0(.CP(n_61681), .D(n_8372), .CD(n_60953), .Q(\nx_tab2[0] 
		));
	notech_mux2 i_11356(.S(\nbus_14516[0] ), .A(\nx_tab2[0] ), .B(n_9982), .Z
		(n_8372));
	notech_reg nx_tab2_reg_1(.CP(n_61681), .D(n_8378), .CD(n_60953), .Q(\nx_tab2[1] 
		));
	notech_mux2 i_11364(.S(\nbus_14516[0] ), .A(\nx_tab2[1] ), .B(n_9984), .Z
		(n_8378));
	notech_ao4 i_603(.A(n_61594), .B(n_10146), .C(n_61534), .D(n_10090), .Z(n_1105
		));
	notech_reg hit_adr11_reg(.CP(n_61681), .D(n_8384), .CD(n_60953), .Q(hit_adr11
		));
	notech_mux2 i_11372(.S(n_872), .A(hit_add11), .B(hit_adr11), .Z(n_8384)
		);
	notech_reg_set tab12_reg_0(.CP(n_61681), .D(n_8390), .SD(n_60953), .Q(\tab12[0] 
		));
	notech_mux2 i_11380(.S(\nbus_14517[0] ), .A(\tab12[0] ), .B(n_56940), .Z
		(n_8390));
	notech_ao4 i_600(.A(n_990), .B(n_9998), .C(n_988), .D(n_10019), .Z(n_1107
		));
	notech_reg_set tab12_reg_1(.CP(n_61681), .D(n_8396), .SD(n_60953), .Q(\tab12[1] 
		));
	notech_mux2 i_11388(.S(\nbus_14517[0] ), .A(\tab12[1] ), .B(n_56946), .Z
		(n_8396));
	notech_reg_set tab12_reg_2(.CP(n_61681), .D(n_8402), .SD(n_60953), .Q(\tab12[2] 
		));
	notech_mux2 i_11396(.S(\nbus_14517[0] ), .A(\tab12[2] ), .B(n_56952), .Z
		(n_8402));
	notech_ao4 i_598(.A(n_998), .B(n_9947), .C(n_996), .D(n_10048), .Z(n_1109
		));
	notech_reg_set tab12_reg_3(.CP(n_61681), .D(n_8408), .SD(n_60953), .Q(\tab12[3] 
		));
	notech_mux2 i_11404(.S(\nbus_14517[0] ), .A(\tab12[3] ), .B(n_56958), .Z
		(n_8408));
	notech_reg tab12_reg_4(.CP(n_61681), .D(n_8414), .CD(n_60953), .Q(\tab12[4] 
		));
	notech_mux2 i_11412(.S(\nbus_14517[0] ), .A(\tab12[4] ), .B(n_873), .Z(n_8414
		));
	notech_and4 i_602(.A(n_1109), .B(n_1107), .C(n_644), .D(n_647), .Z(n_1111
		));
	notech_reg_set tab12_reg_5(.CP(n_61681), .D(n_8420), .SD(n_60953), .Q(\tab12[5] 
		));
	notech_mux2 i_11420(.S(\nbus_14517[0] ), .A(\tab12[5] ), .B(n_56970), .Z
		(n_8420));
	notech_ao4 i_595(.A(n_1003), .B(n_9969), .C(n_1002), .D(n_9924), .Z(n_1112
		));
	notech_reg_set tab12_reg_6(.CP(n_61681), .D(n_8426), .SD(n_60953), .Q(\tab12[6] 
		));
	notech_mux2 i_11428(.S(\nbus_14517[0] ), .A(\tab12[6] ), .B(n_56976), .Z
		(n_8426));
	notech_reg_set tab12_reg_7(.CP(n_61681), .D(n_8432), .SD(n_60953), .Q(\tab12[7] 
		));
	notech_mux2 i_11436(.S(\nbus_14517[0] ), .A(\tab12[7] ), .B(n_56982), .Z
		(n_8432));
	notech_ao4 i_594(.A(n_61594), .B(n_10147), .C(n_61534), .D(n_10091), .Z(n_1114
		));
	notech_reg_set tab12_reg_8(.CP(n_61653), .D(n_8438), .SD(n_60925), .Q(\tab12[8] 
		));
	notech_mux2 i_11444(.S(\nbus_14517[0] ), .A(\tab12[8] ), .B(n_56988), .Z
		(n_8438));
	notech_reg_set tab12_reg_9(.CP(n_61625), .D(n_8444), .SD(n_60897), .Q(\tab12[9] 
		));
	notech_mux2 i_11452(.S(\nbus_14517[0] ), .A(\tab12[9] ), .B(n_56994), .Z
		(n_8444));
	notech_ao4 i_591(.A(n_990), .B(n_9999), .C(n_988), .D(n_10020), .Z(n_1116
		));
	notech_reg_set tab12_reg_10(.CP(n_61625), .D(n_8450), .SD(n_60897), .Q(\tab12[10] 
		));
	notech_mux2 i_11460(.S(\nbus_14517[0] ), .A(\tab12[10] ), .B(n_57000), .Z
		(n_8450));
	notech_reg_set tab12_reg_11(.CP(n_61626), .D(n_8456), .SD(n_60898), .Q(\tab12[11] 
		));
	notech_mux2 i_11468(.S(\nbus_14517[0] ), .A(\tab12[11] ), .B(n_57006), .Z
		(n_8456));
	notech_ao4 i_589(.A(n_998), .B(n_9949), .C(n_996), .D(n_10049), .Z(n_1118
		));
	notech_reg_set tab12_reg_12(.CP(n_61625), .D(n_8462), .SD(n_60897), .Q(\tab12[12] 
		));
	notech_mux2 i_11476(.S(\nbus_14517[0] ), .A(\tab12[12] ), .B(n_57012), .Z
		(n_8462));
	notech_reg_set tab12_reg_13(.CP(n_61625), .D(n_8468), .SD(n_60897), .Q(\tab12[13] 
		));
	notech_mux2 i_11484(.S(\nbus_14517[0] ), .A(\tab12[13] ), .B(n_57018), .Z
		(n_8468));
	notech_and4 i_593(.A(n_1118), .B(n_1116), .C(n_633), .D(n_636), .Z(n_1120
		));
	notech_reg_set tab12_reg_14(.CP(n_61625), .D(n_8474), .SD(n_60897), .Q(\tab12[14] 
		));
	notech_mux2 i_11492(.S(\nbus_14517[0] ), .A(\tab12[14] ), .B(n_57024), .Z
		(n_8474));
	notech_ao4 i_586(.A(n_1003), .B(n_9970), .C(n_1002), .D(n_9925), .Z(n_1121
		));
	notech_reg_set tab12_reg_15(.CP(n_61625), .D(n_8480), .SD(n_60897), .Q(\tab12[15] 
		));
	notech_mux2 i_11500(.S(\nbus_14517[0] ), .A(\tab12[15] ), .B(n_57030), .Z
		(n_8480));
	notech_reg_set tab12_reg_16(.CP(n_61626), .D(n_8486), .SD(n_60898), .Q(\tab12[16] 
		));
	notech_mux2 i_11508(.S(n_60047), .A(\tab12[16] ), .B(n_57036), .Z(n_8486
		));
	notech_ao4 i_585(.A(n_61594), .B(n_10148), .C(n_61534), .D(n_10092), .Z(n_1123
		));
	notech_reg_set tab12_reg_17(.CP(n_61626), .D(n_8492), .SD(n_60898), .Q(\tab12[17] 
		));
	notech_mux2 i_11516(.S(n_60047), .A(\tab12[17] ), .B(n_57042), .Z(n_8492
		));
	notech_reg_set tab12_reg_18(.CP(n_61626), .D(n_8498), .SD(n_60898), .Q(\tab12[18] 
		));
	notech_mux2 i_11524(.S(n_60047), .A(\tab12[18] ), .B(n_57048), .Z(n_8498
		));
	notech_ao4 i_582(.A(n_990), .B(n_10000), .C(n_988), .D(n_10021), .Z(n_1125
		));
	notech_reg_set tab12_reg_19(.CP(n_61626), .D(n_8504), .SD(n_60898), .Q(\tab12[19] 
		));
	notech_mux2 i_11532(.S(n_60047), .A(\tab12[19] ), .B(n_57054), .Z(n_8504
		));
	notech_reg_set tab12_reg_20(.CP(n_61626), .D(n_8510), .SD(n_60898), .Q(\tab12[20] 
		));
	notech_mux2 i_11540(.S(n_60047), .A(\tab12[20] ), .B(n_57060), .Z(n_8510
		));
	notech_ao4 i_580(.A(n_998), .B(n_9950), .C(n_996), .D(n_10050), .Z(n_1127
		));
	notech_reg_set tab12_reg_21(.CP(n_61626), .D(n_8516), .SD(n_60898), .Q(\tab12[21] 
		));
	notech_mux2 i_11548(.S(n_60047), .A(\tab12[21] ), .B(n_57066), .Z(n_8516
		));
	notech_reg_set tab12_reg_22(.CP(n_61626), .D(n_8522), .SD(n_60898), .Q(\tab12[22] 
		));
	notech_mux2 i_11556(.S(n_60047), .A(\tab12[22] ), .B(n_57072), .Z(n_8522
		));
	notech_and4 i_584(.A(n_1127), .B(n_1125), .C(n_622), .D(n_625), .Z(n_1129
		));
	notech_reg_set tab12_reg_23(.CP(n_61625), .D(n_8528), .SD(n_60897), .Q(\tab12[23] 
		));
	notech_mux2 i_11564(.S(n_60047), .A(\tab12[23] ), .B(n_57078), .Z(n_8528
		));
	notech_ao4 i_577(.A(n_1003), .B(n_9971), .C(n_1002), .D(n_9927), .Z(n_1130
		));
	notech_reg_set tab12_reg_24(.CP(n_61621), .D(n_8534), .SD(n_60893), .Q(\tab12[24] 
		));
	notech_mux2 i_11572(.S(n_60047), .A(\tab12[24] ), .B(n_57084), .Z(n_8534
		));
	notech_reg_set tab12_reg_25(.CP(n_61625), .D(n_8540), .SD(n_60897), .Q(\tab12[25] 
		));
	notech_mux2 i_11580(.S(n_60047), .A(\tab12[25] ), .B(n_57090), .Z(n_8540
		));
	notech_ao4 i_576(.A(n_61594), .B(n_10149), .C(n_61534), .D(n_10093), .Z(n_1132
		));
	notech_reg_set tab12_reg_26(.CP(n_61625), .D(n_8546), .SD(n_60897), .Q(\tab12[26] 
		));
	notech_mux2 i_11588(.S(n_60047), .A(\tab12[26] ), .B(n_57096), .Z(n_8546
		));
	notech_reg_set tab12_reg_27(.CP(n_61621), .D(n_8552), .SD(n_60893), .Q(\tab12[27] 
		));
	notech_mux2 i_11596(.S(n_60047), .A(\tab12[27] ), .B(n_57102), .Z(n_8552
		));
	notech_ao4 i_573(.A(n_990), .B(n_10001), .C(n_988), .D(n_10022), .Z(n_1134
		));
	notech_reg_set tab12_reg_28(.CP(n_61621), .D(n_8558), .SD(n_60893), .Q(\tab12[28] 
		));
	notech_mux2 i_11604(.S(n_60047), .A(\tab12[28] ), .B(n_57108), .Z(n_8558
		));
	notech_reg_set tab12_reg_29(.CP(n_61621), .D(n_8564), .SD(n_60893), .Q(\tab12[29] 
		));
	notech_mux2 i_11612(.S(n_60047), .A(\tab12[29] ), .B(n_57114), .Z(n_8564
		));
	notech_ao4 i_571(.A(n_998), .B(n_9951), .C(n_996), .D(n_10051), .Z(n_1136
		));
	notech_reg_set tab12_reg_33(.CP(n_61621), .D(n_8570), .SD(n_60893), .Q(\tab12[33] 
		));
	notech_mux2 i_11620(.S(n_60047), .A(\tab12[33] ), .B(n_57138), .Z(n_8570
		));
	notech_reg hit_adr12_reg(.CP(n_61625), .D(n_8576), .CD(n_60897), .Q(hit_adr12
		));
	notech_mux2 i_11628(.S(n_872), .A(hit_add12), .B(hit_adr12), .Z(n_8576)
		);
	notech_and4 i_575(.A(n_1136), .B(n_1134), .C(n_611), .D(n_614), .Z(n_1138
		));
	notech_reg_set tab13_reg_0(.CP(n_61625), .D(n_8582), .SD(n_60897), .Q(\tab13[0] 
		));
	notech_mux2 i_11636(.S(\nbus_14502[0] ), .A(\tab13[0] ), .B(n_56940), .Z
		(n_8582));
	notech_ao4 i_568(.A(n_1003), .B(n_9972), .C(n_1002), .D(n_9928), .Z(n_1139
		));
	notech_reg_set tab13_reg_1(.CP(n_61625), .D(n_8588), .SD(n_60897), .Q(\tab13[1] 
		));
	notech_mux2 i_11644(.S(\nbus_14502[0] ), .A(\tab13[1] ), .B(n_56946), .Z
		(n_8588));
	notech_reg_set tab13_reg_2(.CP(n_61625), .D(n_8594), .SD(n_60897), .Q(\tab13[2] 
		));
	notech_mux2 i_11652(.S(\nbus_14502[0] ), .A(\tab13[2] ), .B(n_56952), .Z
		(n_8594));
	notech_ao4 i_567(.A(n_61594), .B(n_10150), .C(n_61534), .D(n_10094), .Z(n_1141
		));
	notech_reg_set tab13_reg_3(.CP(n_61625), .D(n_8600), .SD(n_60897), .Q(\tab13[3] 
		));
	notech_mux2 i_11660(.S(\nbus_14502[0] ), .A(\tab13[3] ), .B(n_56958), .Z
		(n_8600));
	notech_reg tab13_reg_4(.CP(n_61625), .D(n_8606), .CD(n_60897), .Q(\tab13[4] 
		));
	notech_mux2 i_11668(.S(\nbus_14502[0] ), .A(\tab13[4] ), .B(n_873), .Z(n_8606
		));
	notech_ao4 i_564(.A(n_990), .B(n_10002), .C(n_988), .D(n_10023), .Z(n_1143
		));
	notech_reg_set tab13_reg_5(.CP(n_61625), .D(n_8612), .SD(n_60897), .Q(\tab13[5] 
		));
	notech_mux2 i_11676(.S(\nbus_14502[0] ), .A(\tab13[5] ), .B(n_56970), .Z
		(n_8612));
	notech_reg_set tab13_reg_6(.CP(n_61626), .D(n_8618), .SD(n_60898), .Q(\tab13[6] 
		));
	notech_mux2 i_11684(.S(\nbus_14502[0] ), .A(\tab13[6] ), .B(n_56976), .Z
		(n_8618));
	notech_ao4 i_562(.A(n_998), .B(n_9952), .C(n_996), .D(n_10052), .Z(n_1145
		));
	notech_reg_set tab13_reg_7(.CP(n_61630), .D(n_8624), .SD(n_60902), .Q(\tab13[7] 
		));
	notech_mux2 i_11692(.S(\nbus_14502[0] ), .A(\tab13[7] ), .B(n_56982), .Z
		(n_8624));
	notech_reg_set tab13_reg_8(.CP(n_61630), .D(n_8630), .SD(n_60902), .Q(\tab13[8] 
		));
	notech_mux2 i_11700(.S(\nbus_14502[0] ), .A(\tab13[8] ), .B(n_56988), .Z
		(n_8630));
	notech_and4 i_566(.A(n_1145), .B(n_1143), .C(n_600), .D(n_603), .Z(n_1147
		));
	notech_reg_set tab13_reg_9(.CP(n_61630), .D(n_8636), .SD(n_60902), .Q(\tab13[9] 
		));
	notech_mux2 i_11708(.S(\nbus_14502[0] ), .A(\tab13[9] ), .B(n_56994), .Z
		(n_8636));
	notech_ao4 i_559(.A(n_1003), .B(n_9973), .C(n_1002), .D(n_9929), .Z(n_1148
		));
	notech_reg_set tab13_reg_10(.CP(n_61630), .D(n_8642), .SD(n_60902), .Q(\tab13[10] 
		));
	notech_mux2 i_11716(.S(\nbus_14502[0] ), .A(\tab13[10] ), .B(n_57000), .Z
		(n_8642));
	notech_reg_set tab13_reg_11(.CP(n_61630), .D(n_8648), .SD(n_60902), .Q(\tab13[11] 
		));
	notech_mux2 i_11724(.S(\nbus_14502[0] ), .A(\tab13[11] ), .B(n_57006), .Z
		(n_8648));
	notech_ao4 i_558(.A(n_61590), .B(n_10151), .C(n_61534), .D(n_10095), .Z(n_1150
		));
	notech_reg_set tab13_reg_12(.CP(n_61630), .D(n_8654), .SD(n_60902), .Q(\tab13[12] 
		));
	notech_mux2 i_11732(.S(\nbus_14502[0] ), .A(\tab13[12] ), .B(n_57012), .Z
		(n_8654));
	notech_reg_set tab13_reg_13(.CP(n_61630), .D(n_8660), .SD(n_60902), .Q(\tab13[13] 
		));
	notech_mux2 i_11740(.S(\nbus_14502[0] ), .A(\tab13[13] ), .B(n_57018), .Z
		(n_8660));
	notech_ao4 i_555(.A(n_990), .B(n_10003), .C(n_988), .D(n_10024), .Z(n_1152
		));
	notech_reg_set tab13_reg_14(.CP(n_61634), .D(n_8666), .SD(n_60906), .Q(\tab13[14] 
		));
	notech_mux2 i_11748(.S(\nbus_14502[0] ), .A(\tab13[14] ), .B(n_57024), .Z
		(n_8666));
	notech_reg_set tab13_reg_15(.CP(n_61634), .D(n_8672), .SD(n_60906), .Q(\tab13[15] 
		));
	notech_mux2 i_11756(.S(\nbus_14502[0] ), .A(\tab13[15] ), .B(n_57030), .Z
		(n_8672));
	notech_ao4 i_553(.A(n_998), .B(n_9953), .C(n_996), .D(n_10053), .Z(n_1154
		));
	notech_reg_set tab13_reg_16(.CP(n_61634), .D(n_8678), .SD(n_60906), .Q(\tab13[16] 
		));
	notech_mux2 i_11764(.S(n_60025), .A(\tab13[16] ), .B(n_57036), .Z(n_8678
		));
	notech_reg_set tab13_reg_17(.CP(n_61630), .D(n_8684), .SD(n_60902), .Q(\tab13[17] 
		));
	notech_mux2 i_11772(.S(n_60025), .A(\tab13[17] ), .B(n_57042), .Z(n_8684
		));
	notech_and4 i_557(.A(n_1154), .B(n_1152), .C(n_589), .D(n_592), .Z(n_1156
		));
	notech_reg_set tab13_reg_18(.CP(n_61630), .D(n_8690), .SD(n_60902), .Q(\tab13[18] 
		));
	notech_mux2 i_11780(.S(n_60025), .A(\tab13[18] ), .B(n_57048), .Z(n_8690
		));
	notech_ao4 i_550(.A(n_1003), .B(n_9974), .C(n_1002), .D(n_9930), .Z(n_1157
		));
	notech_reg_set tab13_reg_19(.CP(n_61630), .D(n_8696), .SD(n_60902), .Q(\tab13[19] 
		));
	notech_mux2 i_11788(.S(n_60025), .A(\tab13[19] ), .B(n_57054), .Z(n_8696
		));
	notech_reg_set tab13_reg_20(.CP(n_61630), .D(n_8702), .SD(n_60902), .Q(\tab13[20] 
		));
	notech_mux2 i_11796(.S(n_60025), .A(\tab13[20] ), .B(n_57060), .Z(n_8702
		));
	notech_ao4 i_549(.A(n_61590), .B(n_10152), .C(n_61534), .D(n_10096), .Z(n_1159
		));
	notech_reg_set tab13_reg_21(.CP(n_61630), .D(n_8708), .SD(n_60902), .Q(\tab13[21] 
		));
	notech_mux2 i_11804(.S(n_60025), .A(\tab13[21] ), .B(n_57066), .Z(n_8708
		));
	notech_reg_set tab13_reg_22(.CP(n_61626), .D(n_8714), .SD(n_60898), .Q(\tab13[22] 
		));
	notech_mux2 i_11812(.S(n_60025), .A(\tab13[22] ), .B(n_57072), .Z(n_8714
		));
	notech_ao4 i_546(.A(n_990), .B(n_10004), .C(n_988), .D(n_10025), .Z(n_1161
		));
	notech_reg_set tab13_reg_23(.CP(n_61626), .D(n_8720), .SD(n_60898), .Q(\tab13[23] 
		));
	notech_mux2 i_11820(.S(n_60025), .A(\tab13[23] ), .B(n_57078), .Z(n_8720
		));
	notech_reg_set tab13_reg_24(.CP(n_61626), .D(n_8726), .SD(n_60898), .Q(\tab13[24] 
		));
	notech_mux2 i_11828(.S(n_60025), .A(\tab13[24] ), .B(n_57084), .Z(n_8726
		));
	notech_ao4 i_544(.A(n_998), .B(n_9954), .C(n_996), .D(n_10054), .Z(n_1163
		));
	notech_reg_set tab13_reg_25(.CP(n_61626), .D(n_8732), .SD(n_60898), .Q(\tab13[25] 
		));
	notech_mux2 i_11836(.S(n_60025), .A(\tab13[25] ), .B(n_57090), .Z(n_8732
		));
	notech_reg_set tab13_reg_26(.CP(n_61626), .D(n_8738), .SD(n_60898), .Q(\tab13[26] 
		));
	notech_mux2 i_11844(.S(n_60025), .A(\tab13[26] ), .B(n_57096), .Z(n_8738
		));
	notech_and4 i_548(.A(n_1163), .B(n_1161), .C(n_578), .D(n_581), .Z(n_1165
		));
	notech_reg_set tab13_reg_27(.CP(n_61626), .D(n_8744), .SD(n_60898), .Q(\tab13[27] 
		));
	notech_mux2 i_11852(.S(n_60025), .A(\tab13[27] ), .B(n_57102), .Z(n_8744
		));
	notech_ao4 i_541(.A(n_1003), .B(n_9975), .C(n_1002), .D(n_9931), .Z(n_1166
		));
	notech_reg_set tab13_reg_28(.CP(n_61626), .D(n_8750), .SD(n_60898), .Q(\tab13[28] 
		));
	notech_mux2 i_11860(.S(n_60025), .A(\tab13[28] ), .B(n_57108), .Z(n_8750
		));
	notech_reg_set tab13_reg_29(.CP(n_61630), .D(n_8756), .SD(n_60902), .Q(\tab13[29] 
		));
	notech_mux2 i_11868(.S(n_60025), .A(\tab13[29] ), .B(n_57114), .Z(n_8756
		));
	notech_ao4 i_540(.A(n_61590), .B(n_10153), .C(n_878), .D(n_10097), .Z(n_1168
		));
	notech_reg_set tab13_reg_33(.CP(n_61630), .D(n_8762), .SD(n_60902), .Q(\tab13[33] 
		));
	notech_mux2 i_11876(.S(n_60025), .A(\tab13[33] ), .B(n_57138), .Z(n_8762
		));
	notech_reg hit_adr13_reg(.CP(n_61630), .D(n_8768), .CD(n_60902), .Q(hit_adr13
		));
	notech_mux2 i_11884(.S(n_872), .A(hit_add13), .B(hit_adr13), .Z(n_8768)
		);
	notech_ao4 i_537(.A(n_990), .B(n_10005), .C(n_988), .D(n_10026), .Z(n_1170
		));
	notech_reg_set tab14_reg_0(.CP(n_61630), .D(n_8774), .SD(n_60902), .Q(\tab14[0] 
		));
	notech_mux2 i_11892(.S(\nbus_14489[0] ), .A(\tab14[0] ), .B(n_56940), .Z
		(n_8774));
	notech_reg_set tab14_reg_1(.CP(n_61626), .D(n_8780), .SD(n_60898), .Q(\tab14[1] 
		));
	notech_mux2 i_11900(.S(\nbus_14489[0] ), .A(\tab14[1] ), .B(n_56946), .Z
		(n_8780));
	notech_ao4 i_535(.A(n_998), .B(n_9955), .C(n_996), .D(n_10055), .Z(n_1172
		));
	notech_reg_set tab14_reg_2(.CP(n_61630), .D(n_8786), .SD(n_60902), .Q(\tab14[2] 
		));
	notech_mux2 i_11908(.S(\nbus_14489[0] ), .A(\tab14[2] ), .B(n_56952), .Z
		(n_8786));
	notech_reg_set tab14_reg_3(.CP(n_61630), .D(n_8792), .SD(n_60902), .Q(\tab14[3] 
		));
	notech_mux2 i_11916(.S(\nbus_14489[0] ), .A(\tab14[3] ), .B(n_56958), .Z
		(n_8792));
	notech_and4 i_539(.A(n_1172), .B(n_1170), .C(n_567), .D(n_570), .Z(n_1174
		));
	notech_reg tab14_reg_4(.CP(n_61616), .D(n_8798), .CD(n_60888), .Q(\tab14[4] 
		));
	notech_mux2 i_11924(.S(\nbus_14489[0] ), .A(\tab14[4] ), .B(n_873), .Z(n_8798
		));
	notech_ao4 i_532(.A(n_1003), .B(n_9976), .C(n_1002), .D(n_9932), .Z(n_1175
		));
	notech_reg_set tab14_reg_5(.CP(n_61616), .D(n_8804), .SD(n_60888), .Q(\tab14[5] 
		));
	notech_mux2 i_11932(.S(\nbus_14489[0] ), .A(\tab14[5] ), .B(n_56970), .Z
		(n_8804));
	notech_reg_set tab14_reg_6(.CP(n_61616), .D(n_8810), .SD(n_60888), .Q(\tab14[6] 
		));
	notech_mux2 i_11940(.S(\nbus_14489[0] ), .A(\tab14[6] ), .B(n_56976), .Z
		(n_8810));
	notech_ao4 i_531(.A(n_61594), .B(n_10154), .C(n_61534), .D(n_10098), .Z(n_1177
		));
	notech_reg_set tab14_reg_7(.CP(n_61616), .D(n_8816), .SD(n_60888), .Q(\tab14[7] 
		));
	notech_mux2 i_11948(.S(\nbus_14489[0] ), .A(\tab14[7] ), .B(n_56982), .Z
		(n_8816));
	notech_reg_set tab14_reg_8(.CP(n_61612), .D(n_8822), .SD(n_60884), .Q(\tab14[8] 
		));
	notech_mux2 i_11956(.S(\nbus_14489[0] ), .A(\tab14[8] ), .B(n_56988), .Z
		(n_8822));
	notech_ao4 i_79167(.A(n_10102), .B(n_10181), .C(n_9940), .D(n_10182), .Z
		(oread_req97003));
	notech_reg_set tab14_reg_9(.CP(n_61616), .D(n_8828), .SD(n_60888), .Q(\tab14[9] 
		));
	notech_mux2 i_11964(.S(\nbus_14489[0] ), .A(\tab14[9] ), .B(n_56994), .Z
		(n_8828));
	notech_nand3 i_80446(.A(n_532), .B(n_388), .C(n_531), .Z(\nbus_14492[0] 
		));
	notech_reg_set tab14_reg_10(.CP(n_61616), .D(n_8834), .SD(n_60888), .Q(\tab14[10] 
		));
	notech_mux2 i_11972(.S(\nbus_14489[0] ), .A(\tab14[10] ), .B(n_57000), .Z
		(n_8834));
	notech_nand3 i_80682(.A(n_532), .B(n_388), .C(n_528), .Z(\nbus_14493[0] 
		));
	notech_reg_set tab14_reg_11(.CP(n_61616), .D(n_8840), .SD(n_60888), .Q(\tab14[11] 
		));
	notech_mux2 i_11980(.S(\nbus_14489[0] ), .A(\tab14[11] ), .B(n_57006), .Z
		(n_8840));
	notech_nand3 i_80794(.A(n_509), .B(n_388), .C(n_508), .Z(\nbus_14494[0] 
		));
	notech_reg_set tab14_reg_12(.CP(n_61616), .D(n_8846), .SD(n_60888), .Q(\tab14[12] 
		));
	notech_mux2 i_11988(.S(\nbus_14489[0] ), .A(\tab14[12] ), .B(n_57012), .Z
		(n_8846));
	notech_nand3 i_81438(.A(n_509), .B(n_388), .C(n_505), .Z(\nbus_14505[0] 
		));
	notech_reg_set tab14_reg_13(.CP(n_61616), .D(n_8852), .SD(n_60888), .Q(\tab14[13] 
		));
	notech_mux2 i_11996(.S(\nbus_14489[0] ), .A(\tab14[13] ), .B(n_57018), .Z
		(n_8852));
	notech_nand3 i_81214(.A(n_509), .B(n_388), .C(n_504), .Z(\nbus_14501[0] 
		));
	notech_reg_set tab14_reg_14(.CP(n_61616), .D(n_8858), .SD(n_60888), .Q(\tab14[14] 
		));
	notech_mux2 i_12004(.S(\nbus_14489[0] ), .A(\tab14[14] ), .B(n_57024), .Z
		(n_8858));
	notech_nand3 i_81672(.A(n_509), .B(n_388), .C(n_503), .Z(\nbus_14514[0] 
		));
	notech_reg_set tab14_reg_15(.CP(n_61616), .D(n_8864), .SD(n_60888), .Q(\tab14[15] 
		));
	notech_mux2 i_12012(.S(\nbus_14489[0] ), .A(\tab14[15] ), .B(n_57030), .Z
		(n_8864));
	notech_ao4 i_81830(.A(n_899), .B(n_900), .C(n_913), .D(n_9926), .Z(\nbus_14515[0] 
		));
	notech_reg_set tab14_reg_16(.CP(n_61616), .D(n_8870), .SD(n_60888), .Q(\tab14[16] 
		));
	notech_mux2 i_12020(.S(n_60014), .A(\tab14[16] ), .B(n_57036), .Z(n_8870
		));
	notech_nand2 i_81847(.A(n_913), .B(n_901), .Z(\nbus_14516[0] ));
	notech_reg_set tab14_reg_17(.CP(n_61616), .D(n_8876), .SD(n_60888), .Q(\tab14[17] 
		));
	notech_mux2 i_12028(.S(n_60014), .A(\tab14[17] ), .B(n_57042), .Z(n_8876
		));
	notech_nand3 i_81866(.A(n_485), .B(n_388), .C(n_484), .Z(\nbus_14517[0] 
		));
	notech_reg_set tab14_reg_18(.CP(n_61612), .D(n_8882), .SD(n_60884), .Q(\tab14[18] 
		));
	notech_mux2 i_12036(.S(n_60014), .A(\tab14[18] ), .B(n_57048), .Z(n_8882
		));
	notech_nand3 i_81326(.A(n_485), .B(n_388), .C(n_483), .Z(\nbus_14502[0] 
		));
	notech_reg_set tab14_reg_19(.CP(n_61612), .D(n_8888), .SD(n_60884), .Q(\tab14[19] 
		));
	notech_mux2 i_12044(.S(n_60014), .A(\tab14[19] ), .B(n_57054), .Z(n_8888
		));
	notech_nand3 i_80190(.A(n_485), .B(n_388), .C(n_482), .Z(\nbus_14489[0] 
		));
	notech_reg_set tab14_reg_20(.CP(n_61612), .D(n_8894), .SD(n_60884), .Q(\tab14[20] 
		));
	notech_mux2 i_12052(.S(n_60014), .A(\tab14[20] ), .B(n_57060), .Z(n_8894
		));
	notech_ao4 i_80328(.A(n_899), .B(n_919), .C(n_913), .D(n_9911), .Z(\nbus_14490[0] 
		));
	notech_reg_set tab14_reg_21(.CP(n_61612), .D(n_8900), .SD(n_60884), .Q(\tab14[21] 
		));
	notech_mux2 i_12060(.S(n_60014), .A(\tab14[21] ), .B(n_57066), .Z(n_8900
		));
	notech_nand2 i_81165(.A(n_913), .B(n_920), .Z(\nbus_14499[0] ));
	notech_reg_set tab14_reg_22(.CP(n_61612), .D(n_8906), .SD(n_60884), .Q(\tab14[22] 
		));
	notech_mux2 i_12068(.S(n_60014), .A(\tab14[22] ), .B(n_57072), .Z(n_8906
		));
	notech_nand3 i_80906(.A(n_485), .B(n_388), .C(n_464), .Z(\nbus_14495[0] 
		));
	notech_reg_set tab14_reg_23(.CP(n_61612), .D(n_8912), .SD(n_60884), .Q(\tab14[23] 
		));
	notech_mux2 i_12076(.S(n_60014), .A(\tab14[23] ), .B(n_57078), .Z(n_8912
		));
	notech_nand2 i_81177(.A(n_893), .B(n_462), .Z(\nbus_14500[0] ));
	notech_reg_set tab14_reg_24(.CP(n_61612), .D(n_8918), .SD(n_60884), .Q(\tab14[24] 
		));
	notech_mux2 i_12084(.S(n_60014), .A(\tab14[24] ), .B(n_57084), .Z(n_8918
		));
	notech_ao4 i_81812(.A(n_461), .B(n_932), .C(n_887), .D(n_10099), .Z(n_59950
		));
	notech_reg_set tab14_reg_25(.CP(n_61612), .D(n_8924), .SD(n_60884), .Q(\tab14[25] 
		));
	notech_mux2 i_12092(.S(n_60014), .A(\tab14[25] ), .B(n_57090), .Z(n_8924
		));
	notech_nand3 i_81025(.A(n_61534), .B(n_59950), .C(n_945), .Z(\nbus_14496[0] 
		));
	notech_reg_set tab14_reg_26(.CP(n_61612), .D(n_8930), .SD(n_60884), .Q(\tab14[26] 
		));
	notech_mux2 i_12100(.S(n_60014), .A(\tab14[26] ), .B(n_57096), .Z(n_8930
		));
	notech_nand2 i_79654(.A(n_938), .B(n_912), .Z(n_58550));
	notech_reg_set tab14_reg_27(.CP(n_61612), .D(n_8936), .SD(n_60884), .Q(\tab14[27] 
		));
	notech_mux2 i_12108(.S(n_60014), .A(\tab14[27] ), .B(n_57102), .Z(n_8936
		));
	notech_ao4 i_81061(.A(n_876), .B(data_miss[5]), .C(n_899), .D(n_934), .Z
		(\nbus_14497[0] ));
	notech_reg_set tab14_reg_28(.CP(n_61612), .D(n_8942), .SD(n_60884), .Q(\tab14[28] 
		));
	notech_mux2 i_12116(.S(n_60014), .A(\tab14[28] ), .B(n_57108), .Z(n_8942
		));
	notech_ao4 i_81043(.A(n_10181), .B(n_10101), .C(n_887), .D(n_10099), .Z(n_58547
		));
	notech_reg_set tab14_reg_29(.CP(n_61612), .D(n_8948), .SD(n_60884), .Q(\tab14[29] 
		));
	notech_mux2 i_12124(.S(n_60014), .A(\tab14[29] ), .B(n_57114), .Z(n_8948
		));
	notech_nand2 i_322380(.A(n_975), .B(n_400), .Z(addr_phys[2]));
	notech_reg_set tab14_reg_33(.CP(n_61612), .D(n_8954), .SD(n_60884), .Q(\tab14[33] 
		));
	notech_mux2 i_12132(.S(n_60014), .A(\tab14[33] ), .B(n_57138), .Z(n_8954
		));
	notech_nand2 i_422381(.A(n_976), .B(n_398), .Z(addr_phys[3]));
	notech_reg hit_adr14_reg(.CP(n_61612), .D(n_8960), .CD(n_60884), .Q(hit_adr14
		));
	notech_mux2 i_12140(.S(n_872), .A(hit_add14), .B(hit_adr14), .Z(n_8960)
		);
	notech_nand2 i_522382(.A(n_977), .B(n_397), .Z(addr_phys[4]));
	notech_reg_set nnx_tab1_reg_0(.CP(n_61612), .D(n_8966), .SD(n_60884), .Q
		(\nnx_tab1[0] ));
	notech_mux2 i_12148(.S(n_10031), .A(\nnx_tab1[0] ), .B(n_10027), .Z(n_8966
		));
	notech_nand2 i_622383(.A(n_978), .B(n_396), .Z(addr_phys[5]));
	notech_reg nnx_tab1_reg_1(.CP(n_61616), .D(n_8972), .CD(n_60888), .Q(\nnx_tab1[1] 
		));
	notech_mux2 i_12156(.S(n_10031), .A(\nnx_tab1[1] ), .B(n_10029), .Z(n_8972
		));
	notech_nand2 i_722384(.A(n_979), .B(n_395), .Z(addr_phys[6]));
	notech_reg nx_tab1_reg_0(.CP(n_61621), .D(n_8978), .CD(n_60893), .Q(\nx_tab1[0] 
		));
	notech_mux2 i_12164(.S(\nbus_14499[0] ), .A(\nx_tab1[0] ), .B(n_10032), 
		.Z(n_8978));
	notech_nand2 i_822385(.A(n_980), .B(n_394), .Z(addr_phys[7]));
	notech_reg nx_tab1_reg_1(.CP(n_61621), .D(n_8984), .CD(n_60893), .Q(\nx_tab1[1] 
		));
	notech_mux2 i_12172(.S(\nbus_14499[0] ), .A(\nx_tab1[1] ), .B(n_10034), 
		.Z(n_8984));
	notech_nand2 i_922386(.A(n_981), .B(n_393), .Z(addr_phys[8]));
	notech_reg_set tab11_reg_0(.CP(n_61621), .D(n_8990), .SD(n_60893), .Q(\tab11[0] 
		));
	notech_mux2 i_12180(.S(\nbus_14495[0] ), .A(\tab11[0] ), .B(n_56940), .Z
		(n_8990));
	notech_nand2 i_1022387(.A(n_982), .B(n_392), .Z(addr_phys[9]));
	notech_reg_set tab11_reg_1(.CP(n_61621), .D(n_8996), .SD(n_60893), .Q(\tab11[1] 
		));
	notech_mux2 i_12188(.S(\nbus_14495[0] ), .A(\tab11[1] ), .B(n_56946), .Z
		(n_8996));
	notech_nand2 i_1122388(.A(n_983), .B(n_391), .Z(addr_phys[10]));
	notech_reg_set tab11_reg_2(.CP(n_61617), .D(n_9002), .SD(n_60889), .Q(\tab11[2] 
		));
	notech_mux2 i_12196(.S(\nbus_14495[0] ), .A(\tab11[2] ), .B(n_56952), .Z
		(n_9002));
	notech_nand2 i_1222389(.A(n_984), .B(n_390), .Z(addr_phys[11]));
	notech_reg_set tab11_reg_3(.CP(n_61617), .D(n_9008), .SD(n_60889), .Q(\tab11[3] 
		));
	notech_mux2 i_12204(.S(\nbus_14495[0] ), .A(\tab11[3] ), .B(n_56958), .Z
		(n_9008));
	notech_and4 i_1322390(.A(n_1004), .B(n_1006), .C(n_1001), .D(n_773), .Z(addr_phys_1297004
		));
	notech_reg tab11_reg_4(.CP(n_61617), .D(n_9014), .CD(n_60889), .Q(\tab11[4] 
		));
	notech_mux2 i_12212(.S(\nbus_14495[0] ), .A(\tab11[4] ), .B(n_873), .Z(n_9014
		));
	notech_and4 i_1422391(.A(n_1013), .B(n_1015), .C(n_1012), .D(n_762), .Z(addr_phys_1397005
		));
	notech_reg_set tab11_reg_5(.CP(n_61621), .D(n_9020), .SD(n_60893), .Q(\tab11[5] 
		));
	notech_mux2 i_12220(.S(\nbus_14495[0] ), .A(\tab11[5] ), .B(n_56970), .Z
		(n_9020));
	notech_and4 i_1522392(.A(n_1022), .B(n_1024), .C(n_1021), .D(n_751), .Z(addr_phys_1497006
		));
	notech_reg_set tab11_reg_6(.CP(n_61621), .D(n_9026), .SD(n_60893), .Q(\tab11[6] 
		));
	notech_mux2 i_12228(.S(\nbus_14495[0] ), .A(\tab11[6] ), .B(n_56976), .Z
		(n_9026));
	notech_and4 i_1622393(.A(n_1031), .B(n_1033), .C(n_1030), .D(n_740), .Z(addr_phys_1597007
		));
	notech_reg_set tab11_reg_7(.CP(n_61621), .D(n_9032), .SD(n_60893), .Q(\tab11[7] 
		));
	notech_mux2 i_12236(.S(\nbus_14495[0] ), .A(\tab11[7] ), .B(n_56982), .Z
		(n_9032));
	notech_and4 i_1722394(.A(n_1040), .B(n_1042), .C(n_1039), .D(n_729), .Z(addr_phys_1697008
		));
	notech_reg_set tab11_reg_8(.CP(n_61621), .D(n_9038), .SD(n_60893), .Q(\tab11[8] 
		));
	notech_mux2 i_12244(.S(\nbus_14495[0] ), .A(\tab11[8] ), .B(n_56988), .Z
		(n_9038));
	notech_and4 i_1822395(.A(n_1049), .B(n_1051), .C(n_1048), .D(n_718), .Z(addr_phys_1797009
		));
	notech_reg_set tab11_reg_9(.CP(n_61621), .D(n_9044), .SD(n_60893), .Q(\tab11[9] 
		));
	notech_mux2 i_12252(.S(\nbus_14495[0] ), .A(\tab11[9] ), .B(n_56994), .Z
		(n_9044));
	notech_and4 i_1922396(.A(n_1058), .B(n_1060), .C(n_1057), .D(n_707), .Z(addr_phys_1897010
		));
	notech_reg_set tab11_reg_10(.CP(n_61621), .D(n_9050), .SD(n_60893), .Q(\tab11[10] 
		));
	notech_mux2 i_12260(.S(\nbus_14495[0] ), .A(\tab11[10] ), .B(n_57000), .Z
		(n_9050));
	notech_and4 i_2022397(.A(n_1067), .B(n_1069), .C(n_1066), .D(n_696), .Z(addr_phys_1997011
		));
	notech_reg_set tab11_reg_11(.CP(n_61621), .D(n_9056), .SD(n_60893), .Q(\tab11[11] 
		));
	notech_mux2 i_12268(.S(\nbus_14495[0] ), .A(\tab11[11] ), .B(n_57006), .Z
		(n_9056));
	notech_and4 i_2122398(.A(n_1076), .B(n_1078), .C(n_1075), .D(n_685), .Z(addr_phys_2097012
		));
	notech_reg_set tab11_reg_12(.CP(n_61617), .D(n_9062), .SD(n_60889), .Q(\tab11[12] 
		));
	notech_mux2 i_12276(.S(\nbus_14495[0] ), .A(\tab11[12] ), .B(n_57012), .Z
		(n_9062));
	notech_and4 i_2222399(.A(n_1085), .B(n_1087), .C(n_1084), .D(n_674), .Z(addr_phys_2197013
		));
	notech_reg_set tab11_reg_13(.CP(n_61617), .D(n_9068), .SD(n_60889), .Q(\tab11[13] 
		));
	notech_mux2 i_12284(.S(\nbus_14495[0] ), .A(\tab11[13] ), .B(n_57018), .Z
		(n_9068));
	notech_and4 i_2322400(.A(n_1094), .B(n_1096), .C(n_1093), .D(n_663), .Z(addr_phys_2297014
		));
	notech_reg_set tab11_reg_14(.CP(n_61617), .D(n_9074), .SD(n_60889), .Q(\tab11[14] 
		));
	notech_mux2 i_12292(.S(\nbus_14495[0] ), .A(\tab11[14] ), .B(n_57024), .Z
		(n_9074));
	notech_and4 i_2422401(.A(n_1103), .B(n_1105), .C(n_1102), .D(n_652), .Z(addr_phys_2397015
		));
	notech_reg_set tab11_reg_15(.CP(n_61617), .D(n_9080), .SD(n_60889), .Q(\tab11[15] 
		));
	notech_mux2 i_12300(.S(\nbus_14495[0] ), .A(\tab11[15] ), .B(n_57030), .Z
		(n_9080));
	notech_and4 i_2522402(.A(n_1112), .B(n_1114), .C(n_1111), .D(n_641), .Z(addr_phys_2497016
		));
	notech_reg_set tab11_reg_16(.CP(n_61617), .D(n_9086), .SD(n_60889), .Q(\tab11[16] 
		));
	notech_mux2 i_12308(.S(n_60036), .A(\tab11[16] ), .B(n_57036), .Z(n_9086
		));
	notech_and4 i_2622403(.A(n_1121), .B(n_1123), .C(n_1120), .D(n_630), .Z(addr_phys_2597017
		));
	notech_reg_set tab11_reg_17(.CP(n_61616), .D(n_9092), .SD(n_60888), .Q(\tab11[17] 
		));
	notech_mux2 i_12316(.S(n_60036), .A(\tab11[17] ), .B(n_57042), .Z(n_9092
		));
	notech_and4 i_2722404(.A(n_1130), .B(n_1132), .C(n_1129), .D(n_619), .Z(addr_phys_2697018
		));
	notech_reg_set tab11_reg_18(.CP(n_61616), .D(n_9098), .SD(n_60888), .Q(\tab11[18] 
		));
	notech_mux2 i_12324(.S(n_60036), .A(\tab11[18] ), .B(n_57048), .Z(n_9098
		));
	notech_and4 i_2822405(.A(n_1139), .B(n_1141), .C(n_1138), .D(n_608), .Z(addr_phys_2797019
		));
	notech_reg_set tab11_reg_19(.CP(n_61617), .D(n_9104), .SD(n_60889), .Q(\tab11[19] 
		));
	notech_mux2 i_12332(.S(n_60036), .A(\tab11[19] ), .B(n_57054), .Z(n_9104
		));
	notech_and4 i_2922406(.A(n_1148), .B(n_1150), .C(n_1147), .D(n_597), .Z(addr_phys_2897020
		));
	notech_reg_set tab11_reg_20(.CP(n_61617), .D(n_9110), .SD(n_60889), .Q(\tab11[20] 
		));
	notech_mux2 i_12340(.S(n_60036), .A(\tab11[20] ), .B(n_57060), .Z(n_9110
		));
	notech_and4 i_3022407(.A(n_1157), .B(n_1159), .C(n_1156), .D(n_586), .Z(addr_phys_2997021
		));
	notech_reg_set tab11_reg_21(.CP(n_61617), .D(n_9116), .SD(n_60889), .Q(\tab11[21] 
		));
	notech_mux2 i_12348(.S(n_60036), .A(\tab11[21] ), .B(n_57066), .Z(n_9116
		));
	notech_and4 i_3122408(.A(n_1166), .B(n_1168), .C(n_1165), .D(n_575), .Z(addr_phys_3097022
		));
	notech_reg_set tab11_reg_22(.CP(n_61617), .D(n_9122), .SD(n_60889), .Q(\tab11[22] 
		));
	notech_mux2 i_12356(.S(n_60036), .A(\tab11[22] ), .B(n_57072), .Z(n_9122
		));
	notech_and4 i_3222409(.A(n_1175), .B(n_1177), .C(n_1174), .D(n_564), .Z(addr_phys_3197023
		));
	notech_reg_set tab11_reg_23(.CP(n_61617), .D(n_9128), .SD(n_60889), .Q(\tab11[23] 
		));
	notech_mux2 i_12364(.S(n_60036), .A(\tab11[23] ), .B(n_57078), .Z(n_9128
		));
	notech_mux2 i_122921(.S(n_61570), .A(iDaddr[12]), .B(iDaddr_f[12]), .Z(\tab11_0[0] 
		));
	notech_reg_set tab11_reg_24(.CP(n_61617), .D(n_9134), .SD(n_60889), .Q(\tab11[24] 
		));
	notech_mux2 i_12372(.S(n_60036), .A(\tab11[24] ), .B(n_57084), .Z(n_9134
		));
	notech_mux2 i_222922(.S(n_61570), .A(iDaddr[13]), .B(iDaddr_f[13]), .Z(\tab11_0[1] 
		));
	notech_reg_set tab11_reg_25(.CP(n_61617), .D(n_9140), .SD(n_60889), .Q(\tab11[25] 
		));
	notech_mux2 i_12380(.S(n_60036), .A(\tab11[25] ), .B(n_57090), .Z(n_9140
		));
	notech_mux2 i_322923(.S(n_61570), .A(iDaddr[14]), .B(iDaddr_f[14]), .Z(\tab11_0[2] 
		));
	notech_reg_set tab11_reg_26(.CP(n_61617), .D(n_9146), .SD(n_60889), .Q(\tab11[26] 
		));
	notech_mux2 i_12388(.S(n_60036), .A(\tab11[26] ), .B(n_57096), .Z(n_9146
		));
	notech_mux2 i_422924(.S(n_61570), .A(iDaddr[15]), .B(iDaddr_f[15]), .Z(\tab11_0[3] 
		));
	notech_reg_set tab11_reg_27(.CP(n_61634), .D(n_9152), .SD(n_60906), .Q(\tab11[27] 
		));
	notech_mux2 i_12396(.S(n_60036), .A(\tab11[27] ), .B(n_57102), .Z(n_9152
		));
	notech_mux2 i_522925(.S(n_61570), .A(iDaddr[16]), .B(iDaddr_f[16]), .Z(\tab11_0[4] 
		));
	notech_reg_set tab11_reg_28(.CP(n_61645), .D(n_9158), .SD(n_60917), .Q(\tab11[28] 
		));
	notech_mux2 i_12404(.S(n_60036), .A(\tab11[28] ), .B(n_57108), .Z(n_9158
		));
	notech_mux2 i_622926(.S(n_61570), .A(iDaddr[17]), .B(iDaddr_f[17]), .Z(\tab11_0[5] 
		));
	notech_reg_set tab11_reg_29(.CP(n_61645), .D(n_9164), .SD(n_60917), .Q(\tab11[29] 
		));
	notech_mux2 i_12412(.S(n_60036), .A(\tab11[29] ), .B(n_57114), .Z(n_9164
		));
	notech_mux2 i_722927(.S(n_61570), .A(iDaddr[18]), .B(iDaddr_f[18]), .Z(\tab11_0[6] 
		));
	notech_reg_set tab11_reg_33(.CP(n_61645), .D(n_9170), .SD(n_60917), .Q(\tab11[33] 
		));
	notech_mux2 i_12420(.S(n_60036), .A(\tab11[33] ), .B(n_57138), .Z(n_9170
		));
	notech_mux2 i_822928(.S(n_61570), .A(iDaddr[19]), .B(iDaddr_f[19]), .Z(\tab11_0[7] 
		));
	notech_reg fsm5_cnt_reg_0(.CP(n_61645), .D(n_9176), .CD(n_60917), .Q(fsm5_cnt
		[0]));
	notech_mux2 i_12428(.S(\nbus_14500[0] ), .A(fsm5_cnt[0]), .B(n_863), .Z(n_9176
		));
	notech_mux2 i_922929(.S(n_61570), .A(iDaddr[20]), .B(iDaddr_f[20]), .Z(\tab11_0[8] 
		));
	notech_reg fsm5_cnt_reg_1(.CP(n_61645), .D(n_9182), .CD(n_60917), .Q(fsm5_cnt
		[1]));
	notech_mux2 i_12436(.S(\nbus_14500[0] ), .A(fsm5_cnt[1]), .B(n_864), .Z(n_9182
		));
	notech_mux2 i_1022930(.S(n_61570), .A(iDaddr[21]), .B(iDaddr_f[21]), .Z(\tab11_0[9] 
		));
	notech_reg fsm5_cnt_reg_2(.CP(n_61645), .D(n_9188), .CD(n_60917), .Q(fsm5_cnt
		[2]));
	notech_mux2 i_12444(.S(\nbus_14500[0] ), .A(fsm5_cnt[2]), .B(n_865), .Z(n_9188
		));
	notech_mux2 i_1122931(.S(n_61575), .A(iDaddr[22]), .B(iDaddr_f[22]), .Z(\dir1_0[0] 
		));
	notech_reg fsm5_cnt_reg_3(.CP(n_61645), .D(n_9194), .CD(n_60917), .Q(fsm5_cnt
		[3]));
	notech_mux2 i_12452(.S(\nbus_14500[0] ), .A(fsm5_cnt[3]), .B(n_866), .Z(n_9194
		));
	notech_mux2 i_1222932(.S(n_61575), .A(iDaddr[23]), .B(iDaddr_f[23]), .Z(\dir1_0[1] 
		));
	notech_reg fsm5_cnt_reg_4(.CP(n_61645), .D(n_9200), .CD(n_60917), .Q(fsm5_cnt
		[4]));
	notech_mux2 i_12460(.S(\nbus_14500[0] ), .A(fsm5_cnt[4]), .B(n_867), .Z(n_9200
		));
	notech_mux2 i_1322933(.S(n_61575), .A(iDaddr[24]), .B(iDaddr_f[24]), .Z(\dir1_0[2] 
		));
	notech_reg fsm5_cnt_reg_5(.CP(n_61649), .D(n_9206), .CD(n_60921), .Q(fsm5_cnt
		[5]));
	notech_mux2 i_12468(.S(\nbus_14500[0] ), .A(fsm5_cnt[5]), .B(n_868), .Z(n_9206
		));
	notech_mux2 i_1422934(.S(n_61575), .A(iDaddr[25]), .B(iDaddr_f[25]), .Z(\dir1_0[3] 
		));
	notech_reg fsm5_cnt_reg_6(.CP(n_61649), .D(n_9212), .CD(n_60921), .Q(fsm5_cnt
		[6]));
	notech_mux2 i_12476(.S(\nbus_14500[0] ), .A(fsm5_cnt[6]), .B(n_869), .Z(n_9212
		));
	notech_mux2 i_1522935(.S(n_61575), .A(iDaddr[26]), .B(iDaddr_f[26]), .Z(\dir1_0[4] 
		));
	notech_reg fsm5_cnt_reg_7(.CP(n_61645), .D(n_9218), .CD(n_60917), .Q(fsm5_cnt
		[7]));
	notech_mux2 i_12484(.S(\nbus_14500[0] ), .A(fsm5_cnt[7]), .B(n_870), .Z(n_9218
		));
	notech_mux2 i_1622936(.S(n_61575), .A(iDaddr[27]), .B(iDaddr_f[27]), .Z(\dir1_0[5] 
		));
	notech_reg fsm5_cnt_reg_8(.CP(n_61645), .D(n_9224), .CD(n_60917), .Q(fsm5_cnt
		[8]));
	notech_mux2 i_12492(.S(\nbus_14500[0] ), .A(fsm5_cnt[8]), .B(n_871), .Z(n_9224
		));
	notech_mux2 i_1722937(.S(n_61575), .A(iDaddr[28]), .B(iDaddr_f[28]), .Z(\dir1_0[6] 
		));
	notech_reg pg_fault_reg(.CP(n_61645), .D(n_9230), .CD(n_60917), .Q(pg_fault
		));
	notech_mux2 i_12500(.S(n_10056), .A(pg_fault), .B(n_862), .Z(n_9230));
	notech_mux2 i_1822938(.S(n_61575), .A(iDaddr[29]), .B(iDaddr_f[29]), .Z(\dir1_0[7] 
		));
	notech_reg fsm_reg_0(.CP(n_61645), .D(n_9236), .CD(n_60917), .Q(fsm[0])
		);
	notech_mux2 i_12508(.S(\nbus_14496[0] ), .A(n_61579), .B(n_58520), .Z(n_9236
		));
	notech_mux2 i_1922939(.S(n_61575), .A(iDaddr[30]), .B(iDaddr_f[30]), .Z(\dir1_0[8] 
		));
	notech_reg fsm_reg_1(.CP(n_61645), .D(n_9242), .CD(n_60917), .Q(fsm[1])
		);
	notech_mux2 i_12516(.S(\nbus_14496[0] ), .A(fsm[1]), .B(n_58526), .Z(n_9242
		));
	notech_mux2 i_2022940(.S(n_61575), .A(iDaddr[31]), .B(iDaddr_f[31]), .Z(\dir1_0[9] 
		));
	notech_reg fsm_reg_2(.CP(n_61644), .D(n_9248), .CD(n_60916), .Q(fsm[2])
		);
	notech_mux2 i_12524(.S(\nbus_14496[0] ), .A(fsm[2]), .B(n_58532), .Z(n_9248
		));
	notech_nand3 i_79273(.A(n_60436), .B(n_61575), .C(n_10165), .Z(n_57419)
		);
	notech_reg fsm_reg_3(.CP(n_61644), .D(n_9254), .CD(n_60916), .Q(fsm[3])
		);
	notech_mux2 i_12532(.S(\nbus_14496[0] ), .A(fsm[3]), .B(n_861), .Z(n_9254
		));
	notech_nand3 i_79275(.A(n_60436), .B(n_61575), .C(n_10164), .Z(n_57425)
		);
	notech_reg addr_miss_reg_2(.CP(n_61644), .D(n_9260), .CD(n_60916), .Q(\addr_miss[2] 
		));
	notech_mux2 i_12540(.S(n_853), .A(n_10059), .B(\addr_miss[2] ), .Z(n_9260
		));
	notech_nand3 i_79277(.A(n_60436), .B(n_61573), .C(n_10163), .Z(n_57431)
		);
	notech_reg addr_miss_reg_3(.CP(n_61644), .D(n_9266), .CD(n_60916), .Q(\addr_miss[3] 
		));
	notech_mux2 i_12548(.S(n_853), .A(n_10060), .B(\addr_miss[3] ), .Z(n_9266
		));
	notech_nand3 i_79279(.A(n_60436), .B(n_61573), .C(n_10162), .Z(n_57437)
		);
	notech_reg addr_miss_reg_4(.CP(n_61644), .D(n_9272), .CD(n_60916), .Q(\addr_miss[4] 
		));
	notech_mux2 i_12556(.S(n_853), .A(n_10061), .B(\addr_miss[4] ), .Z(n_9272
		));
	notech_nand3 i_79283(.A(n_60436), .B(n_61573), .C(n_10160), .Z(n_57449)
		);
	notech_reg addr_miss_reg_5(.CP(n_61644), .D(n_9278), .CD(n_60916), .Q(\addr_miss[5] 
		));
	notech_mux2 i_12564(.S(n_853), .A(n_10062), .B(\addr_miss[5] ), .Z(n_9278
		));
	notech_nand3 i_79285(.A(n_60436), .B(n_61573), .C(n_10159), .Z(n_57455)
		);
	notech_reg addr_miss_reg_6(.CP(n_61644), .D(n_9284), .CD(n_60916), .Q(\addr_miss[6] 
		));
	notech_mux2 i_12572(.S(n_853), .A(n_10063), .B(\addr_miss[6] ), .Z(n_9284
		));
	notech_nand3 i_79287(.A(n_60436), .B(n_61573), .C(n_10158), .Z(n_57461)
		);
	notech_reg addr_miss_reg_7(.CP(n_61645), .D(n_9290), .CD(n_60917), .Q(\addr_miss[7] 
		));
	notech_mux2 i_12580(.S(n_853), .A(n_10064), .B(\addr_miss[7] ), .Z(n_9290
		));
	notech_nand3 i_79289(.A(n_60436), .B(n_61573), .C(n_10157), .Z(n_57467)
		);
	notech_reg addr_miss_reg_8(.CP(n_61645), .D(n_9296), .CD(n_60917), .Q(\addr_miss[8] 
		));
	notech_mux2 i_12588(.S(n_853), .A(n_10065), .B(\addr_miss[8] ), .Z(n_9296
		));
	notech_nand3 i_79291(.A(n_60436), .B(n_61575), .C(n_10156), .Z(n_57473)
		);
	notech_reg addr_miss_reg_9(.CP(n_61645), .D(n_9302), .CD(n_60917), .Q(\addr_miss[9] 
		));
	notech_mux2 i_12596(.S(n_853), .A(n_10066), .B(\addr_miss[9] ), .Z(n_9302
		));
	notech_nao3 i_79293(.A(n_61575), .B(n_60436), .C(data_miss[12]), .Z(n_57479
		));
	notech_reg addr_miss_reg_10(.CP(n_61645), .D(n_9308), .CD(n_60917), .Q(\addr_miss[10] 
		));
	notech_mux2 i_12604(.S(n_853), .A(n_10067), .B(\addr_miss[10] ), .Z(n_9308
		));
	notech_nao3 i_79295(.A(n_61575), .B(n_60436), .C(data_miss[13]), .Z(n_57485
		));
	notech_reg addr_miss_reg_11(.CP(n_61644), .D(n_9314), .CD(n_60916), .Q(\addr_miss[11] 
		));
	notech_mux2 i_12612(.S(n_853), .A(n_10068), .B(\addr_miss[11] ), .Z(n_9314
		));
	notech_nao3 i_79297(.A(n_61573), .B(n_60436), .C(data_miss[14]), .Z(n_57491
		));
	notech_reg addr_miss_reg_12(.CP(n_61644), .D(n_9320), .CD(n_60916), .Q(\addr_miss[12] 
		));
	notech_mux2 i_12620(.S(n_853), .A(n_59588), .B(\addr_miss[12] ), .Z(n_9320
		));
	notech_nao3 i_79299(.A(n_61575), .B(n_60436), .C(data_miss[15]), .Z(n_57497
		));
	notech_reg addr_miss_reg_13(.CP(n_61645), .D(n_9326), .CD(n_60917), .Q(\addr_miss[13] 
		));
	notech_mux2 i_12628(.S(n_853), .A(n_59594), .B(\addr_miss[13] ), .Z(n_9326
		));
	notech_nao3 i_79301(.A(n_61570), .B(n_60432), .C(data_miss[16]), .Z(n_57503
		));
	notech_reg addr_miss_reg_14(.CP(n_61649), .D(n_9332), .CD(n_60921), .Q(\addr_miss[14] 
		));
	notech_mux2 i_12636(.S(n_853), .A(n_59600), .B(\addr_miss[14] ), .Z(n_9332
		));
	notech_nao3 i_79303(.A(n_61565), .B(n_60432), .C(data_miss[17]), .Z(n_57509
		));
	notech_reg addr_miss_reg_15(.CP(n_61653), .D(n_9338), .CD(n_60925), .Q(\addr_miss[15] 
		));
	notech_mux2 i_12644(.S(n_853), .A(n_59606), .B(\addr_miss[15] ), .Z(n_9338
		));
	notech_nao3 i_79305(.A(n_61565), .B(n_60432), .C(data_miss[18]), .Z(n_57515
		));
	notech_reg addr_miss_reg_16(.CP(n_61653), .D(n_9344), .CD(n_60925), .Q(\addr_miss[16] 
		));
	notech_mux2 i_12652(.S(n_853), .A(n_59612), .B(\addr_miss[16] ), .Z(n_9344
		));
	notech_nao3 i_79307(.A(n_61565), .B(n_60432), .C(data_miss[19]), .Z(n_57521
		));
	notech_reg addr_miss_reg_17(.CP(n_61653), .D(n_9350), .CD(n_60925), .Q(\addr_miss[17] 
		));
	notech_mux2 i_12660(.S(n_60441), .A(n_59618), .B(\addr_miss[17] ), .Z(n_9350
		));
	notech_nao3 i_79309(.A(n_61563), .B(n_60432), .C(data_miss[20]), .Z(n_57527
		));
	notech_reg addr_miss_reg_18(.CP(n_61653), .D(n_9356), .CD(n_60925), .Q(\addr_miss[18] 
		));
	notech_mux2 i_12668(.S(n_60441), .A(n_59624), .B(\addr_miss[18] ), .Z(n_9356
		));
	notech_nao3 i_79311(.A(n_61563), .B(n_60432), .C(data_miss[21]), .Z(n_57533
		));
	notech_reg addr_miss_reg_19(.CP(n_61653), .D(n_9362), .CD(n_60925), .Q(\addr_miss[19] 
		));
	notech_mux2 i_12676(.S(n_60441), .A(n_59630), .B(\addr_miss[19] ), .Z(n_9362
		));
	notech_nao3 i_79313(.A(n_61565), .B(n_60432), .C(data_miss[22]), .Z(n_57539
		));
	notech_reg addr_miss_reg_20(.CP(n_61653), .D(n_9368), .CD(n_60925), .Q(\addr_miss[20] 
		));
	notech_mux2 i_12684(.S(n_60441), .A(n_59636), .B(\addr_miss[20] ), .Z(n_9368
		));
	notech_nao3 i_79315(.A(n_61565), .B(n_60432), .C(data_miss[23]), .Z(n_57545
		));
	notech_reg addr_miss_reg_21(.CP(n_61653), .D(n_9374), .CD(n_60925), .Q(\addr_miss[21] 
		));
	notech_mux2 i_12692(.S(n_60441), .A(n_59642), .B(\addr_miss[21] ), .Z(n_9374
		));
	notech_nao3 i_79317(.A(n_61565), .B(n_60432), .C(data_miss[24]), .Z(n_57551
		));
	notech_reg addr_miss_reg_22(.CP(n_61653), .D(n_9380), .CD(n_60925), .Q(\addr_miss[22] 
		));
	notech_mux2 i_12700(.S(n_60441), .A(n_59648), .B(\addr_miss[22] ), .Z(n_9380
		));
	notech_nao3 i_79319(.A(n_61565), .B(n_60432), .C(data_miss[25]), .Z(n_57557
		));
	notech_reg addr_miss_reg_23(.CP(n_61653), .D(n_9386), .CD(n_60925), .Q(\addr_miss[23] 
		));
	notech_mux2 i_12708(.S(n_60441), .A(n_59654), .B(\addr_miss[23] ), .Z(n_9386
		));
	notech_nao3 i_79321(.A(n_61565), .B(n_60432), .C(data_miss[26]), .Z(n_57563
		));
	notech_reg addr_miss_reg_24(.CP(n_61653), .D(n_9392), .CD(n_60925), .Q(\addr_miss[24] 
		));
	notech_mux2 i_12716(.S(n_60441), .A(n_59660), .B(\addr_miss[24] ), .Z(n_9392
		));
	notech_nao3 i_79323(.A(n_61565), .B(n_60432), .C(data_miss[27]), .Z(n_57569
		));
	notech_reg addr_miss_reg_25(.CP(n_61653), .D(n_9398), .CD(n_60925), .Q(\addr_miss[25] 
		));
	notech_mux2 i_12724(.S(n_60441), .A(n_59666), .B(\addr_miss[25] ), .Z(n_9398
		));
	notech_nao3 i_79325(.A(n_61563), .B(n_60432), .C(data_miss[28]), .Z(n_57575
		));
	notech_reg addr_miss_reg_26(.CP(n_61653), .D(n_9404), .CD(n_60925), .Q(\addr_miss[26] 
		));
	notech_mux2 i_12732(.S(n_60441), .A(n_59672), .B(\addr_miss[26] ), .Z(n_9404
		));
	notech_nao3 i_79327(.A(n_61563), .B(n_60432), .C(data_miss[29]), .Z(n_57581
		));
	notech_reg addr_miss_reg_27(.CP(n_61653), .D(n_9410), .CD(n_60925), .Q(\addr_miss[27] 
		));
	notech_mux2 i_12740(.S(n_60441), .A(n_59678), .B(\addr_miss[27] ), .Z(n_9410
		));
	notech_nao3 i_79329(.A(n_61563), .B(n_60432), .C(data_miss[30]), .Z(n_57587
		));
	notech_reg addr_miss_reg_28(.CP(n_61653), .D(n_9416), .CD(n_60925), .Q(\addr_miss[28] 
		));
	notech_mux2 i_12748(.S(n_60441), .A(n_59684), .B(\addr_miss[28] ), .Z(n_9416
		));
	notech_nao3 i_79331(.A(n_61563), .B(n_60432), .C(data_miss[31]), .Z(n_57593
		));
	notech_reg addr_miss_reg_29(.CP(n_61649), .D(n_9422), .CD(n_60921), .Q(\addr_miss[29] 
		));
	notech_mux2 i_12756(.S(n_60441), .A(n_59690), .B(\addr_miss[29] ), .Z(n_9422
		));
	notech_nand2 i_79337(.A(n_61563), .B(n_60432), .Z(n_57618));
	notech_reg addr_miss_reg_30(.CP(n_61649), .D(n_9428), .CD(n_60921), .Q(\addr_miss[30] 
		));
	notech_mux2 i_12764(.S(n_60441), .A(n_59696), .B(\addr_miss[30] ), .Z(n_9428
		));
	notech_nand2 i_79574(.A(n_896), .B(n_890), .Z(n_58573));
	notech_reg addr_miss_reg_31(.CP(n_61649), .D(n_9434), .CD(n_60921), .Q(\addr_miss[31] 
		));
	notech_mux2 i_12772(.S(n_60441), .A(n_59702), .B(\addr_miss[31] ), .Z(n_9434
		));
	notech_ao4 i_79467(.A(n_938), .B(n_10165), .C(n_912), .D(n_10175), .Z(n_59528
		));
	notech_reg wrA_reg_2(.CP(n_61649), .D(n_9440), .CD(n_60921), .Q(\wrA[2] 
		));
	notech_mux2 i_12780(.S(n_59983), .A(\wrA[2] ), .B(\addr_miss[2] ), .Z(n_9440
		));
	notech_ao4 i_79470(.A(n_938), .B(n_10164), .C(n_912), .D(n_10174), .Z(n_59534
		));
	notech_reg wrA_reg_3(.CP(n_61649), .D(n_9446), .CD(n_60921), .Q(\wrA[3] 
		));
	notech_mux2 i_12788(.S(n_59983), .A(\wrA[3] ), .B(\addr_miss[3] ), .Z(n_9446
		));
	notech_ao4 i_79473(.A(n_938), .B(n_10163), .C(n_912), .D(n_10173), .Z(n_59540
		));
	notech_reg wrA_reg_4(.CP(n_61649), .D(n_9452), .CD(n_60921), .Q(\wrA[4] 
		));
	notech_mux2 i_12796(.S(n_59983), .A(\wrA[4] ), .B(\addr_miss[4] ), .Z(n_9452
		));
	notech_ao4 i_79476(.A(n_938), .B(n_10162), .C(n_912), .D(n_10172), .Z(n_59546
		));
	notech_reg wrA_reg_5(.CP(n_61649), .D(n_9458), .CD(n_60921), .Q(\wrA[5] 
		));
	notech_mux2 i_12804(.S(n_59983), .A(\wrA[5] ), .B(\addr_miss[5] ), .Z(n_9458
		));
	notech_ao4 i_79479(.A(n_938), .B(n_10161), .C(n_912), .D(n_10171), .Z(n_59552
		));
	notech_reg wrA_reg_6(.CP(n_61649), .D(n_9464), .CD(n_60921), .Q(\wrA[6] 
		));
	notech_mux2 i_12812(.S(n_59983), .A(\wrA[6] ), .B(\addr_miss[6] ), .Z(n_9464
		));
	notech_ao4 i_79482(.A(n_938), .B(n_10160), .C(n_912), .D(n_10170), .Z(n_59558
		));
	notech_reg wrA_reg_7(.CP(n_61649), .D(n_9470), .CD(n_60921), .Q(\wrA[7] 
		));
	notech_mux2 i_12820(.S(n_59983), .A(\wrA[7] ), .B(\addr_miss[7] ), .Z(n_9470
		));
	notech_ao4 i_79485(.A(n_938), .B(n_10159), .C(n_912), .D(n_10169), .Z(n_59564
		));
	notech_reg wrA_reg_8(.CP(n_61649), .D(n_9476), .CD(n_60921), .Q(\wrA[8] 
		));
	notech_mux2 i_12828(.S(n_59983), .A(\wrA[8] ), .B(\addr_miss[8] ), .Z(n_9476
		));
	notech_ao4 i_79488(.A(n_938), .B(n_10158), .C(n_912), .D(n_10168), .Z(n_59570
		));
	notech_reg wrA_reg_9(.CP(n_61649), .D(n_9482), .CD(n_60921), .Q(\wrA[9] 
		));
	notech_mux2 i_12836(.S(n_59983), .A(\wrA[9] ), .B(\addr_miss[9] ), .Z(n_9482
		));
	notech_ao4 i_79491(.A(n_938), .B(n_10157), .C(n_912), .D(n_10167), .Z(n_59576
		));
	notech_reg wrA_reg_10(.CP(n_61649), .D(n_9488), .CD(n_60921), .Q(\wrA[10] 
		));
	notech_mux2 i_12844(.S(n_59983), .A(\wrA[10] ), .B(\addr_miss[10] ), .Z(n_9488
		));
	notech_ao4 i_79494(.A(n_938), .B(n_10156), .C(n_912), .D(n_10166), .Z(n_59582
		));
	notech_reg wrA_reg_11(.CP(n_61649), .D(n_9494), .CD(n_60921), .Q(\wrA[11] 
		));
	notech_mux2 i_12852(.S(n_59983), .A(\wrA[11] ), .B(\addr_miss[11] ), .Z(n_9494
		));
	notech_nand2 i_79497(.A(n_970), .B(n_424), .Z(n_59588));
	notech_reg wrA_reg_12(.CP(n_61649), .D(n_9500), .CD(n_60921), .Q(\wrA[12] 
		));
	notech_mux2 i_12860(.S(n_59983), .A(\wrA[12] ), .B(\addr_miss[12] ), .Z(n_9500
		));
	notech_nand2 i_79500(.A(n_969), .B(n_425), .Z(n_59594));
	notech_reg wrA_reg_13(.CP(n_61649), .D(n_9506), .CD(n_60921), .Q(\wrA[13] 
		));
	notech_mux2 i_12868(.S(n_59983), .A(\wrA[13] ), .B(\addr_miss[13] ), .Z(n_9506
		));
	notech_nand2 i_79503(.A(n_968), .B(n_426), .Z(n_59600));
	notech_reg wrA_reg_14(.CP(n_61635), .D(n_9512), .CD(n_60907), .Q(\wrA[14] 
		));
	notech_mux2 i_12876(.S(n_59983), .A(\wrA[14] ), .B(\addr_miss[14] ), .Z(n_9512
		));
	notech_nand2 i_79506(.A(n_967), .B(n_427), .Z(n_59606));
	notech_reg wrA_reg_15(.CP(n_61635), .D(n_9518), .CD(n_60907), .Q(\wrA[15] 
		));
	notech_mux2 i_12884(.S(n_59983), .A(\wrA[15] ), .B(\addr_miss[15] ), .Z(n_9518
		));
	notech_nand2 i_79509(.A(n_966), .B(n_428), .Z(n_59612));
	notech_reg wrA_reg_16(.CP(n_61635), .D(n_9524), .CD(n_60907), .Q(\wrA[16] 
		));
	notech_mux2 i_12892(.S(n_59983), .A(\wrA[16] ), .B(\addr_miss[16] ), .Z(n_9524
		));
	notech_nand2 i_79512(.A(n_965), .B(n_429), .Z(n_59618));
	notech_reg wrA_reg_17(.CP(n_61635), .D(n_9530), .CD(n_60907), .Q(\wrA[17] 
		));
	notech_mux2 i_12900(.S(n_59983), .A(\wrA[17] ), .B(\addr_miss[17] ), .Z(n_9530
		));
	notech_nand2 i_79515(.A(n_964), .B(n_430), .Z(n_59624));
	notech_reg wrA_reg_18(.CP(n_61635), .D(n_9536), .CD(n_60907), .Q(\wrA[18] 
		));
	notech_mux2 i_12908(.S(n_59983), .A(\wrA[18] ), .B(\addr_miss[18] ), .Z(n_9536
		));
	notech_nand2 i_79518(.A(n_963), .B(n_431), .Z(n_59630));
	notech_reg wrA_reg_19(.CP(n_61635), .D(n_9542), .CD(n_60907), .Q(\wrA[19] 
		));
	notech_mux2 i_12916(.S(n_59983), .A(\wrA[19] ), .B(\addr_miss[19] ), .Z(n_9542
		));
	notech_nand2 i_79521(.A(n_962), .B(n_432), .Z(n_59636));
	notech_reg wrA_reg_20(.CP(n_61635), .D(n_9548), .CD(n_60907), .Q(\wrA[20] 
		));
	notech_mux2 i_12924(.S(n_59983), .A(\wrA[20] ), .B(\addr_miss[20] ), .Z(n_9548
		));
	notech_nand2 i_79524(.A(n_961), .B(n_433), .Z(n_59642));
	notech_reg wrA_reg_21(.CP(n_61635), .D(n_9554), .CD(n_60907), .Q(\wrA[21] 
		));
	notech_mux2 i_12932(.S(n_59977), .A(\wrA[21] ), .B(\addr_miss[21] ), .Z(n_9554
		));
	notech_nand2 i_79527(.A(n_960), .B(n_434), .Z(n_59648));
	notech_reg wrA_reg_22(.CP(n_61635), .D(n_9560), .CD(n_60907), .Q(\wrA[22] 
		));
	notech_mux2 i_12940(.S(n_59977), .A(\wrA[22] ), .B(\addr_miss[22] ), .Z(n_9560
		));
	notech_nand2 i_79530(.A(n_959), .B(n_435), .Z(n_59654));
	notech_reg wrA_reg_23(.CP(n_61635), .D(n_9566), .CD(n_60907), .Q(\wrA[23] 
		));
	notech_mux2 i_12948(.S(n_59977), .A(\wrA[23] ), .B(\addr_miss[23] ), .Z(n_9566
		));
	notech_nand2 i_79533(.A(n_958), .B(n_436), .Z(n_59660));
	notech_reg wrA_reg_24(.CP(n_61635), .D(n_9572), .CD(n_60907), .Q(\wrA[24] 
		));
	notech_mux2 i_12956(.S(n_59977), .A(\wrA[24] ), .B(\addr_miss[24] ), .Z(n_9572
		));
	notech_nand2 i_79536(.A(n_957), .B(n_437), .Z(n_59666));
	notech_reg wrA_reg_25(.CP(n_61635), .D(n_9578), .CD(n_60907), .Q(\wrA[25] 
		));
	notech_mux2 i_12964(.S(n_59977), .A(\wrA[25] ), .B(\addr_miss[25] ), .Z(n_9578
		));
	notech_nand2 i_79539(.A(n_956), .B(n_438), .Z(n_59672));
	notech_reg wrA_reg_26(.CP(n_61635), .D(n_9584), .CD(n_60907), .Q(\wrA[26] 
		));
	notech_mux2 i_12972(.S(n_59977), .A(\wrA[26] ), .B(\addr_miss[26] ), .Z(n_9584
		));
	notech_nand2 i_79542(.A(n_955), .B(n_439), .Z(n_59678));
	notech_reg wrA_reg_27(.CP(n_61635), .D(n_9590), .CD(n_60907), .Q(\wrA[27] 
		));
	notech_mux2 i_12980(.S(n_59977), .A(\wrA[27] ), .B(\addr_miss[27] ), .Z(n_9590
		));
	notech_nand2 i_79545(.A(n_954), .B(n_440), .Z(n_59684));
	notech_reg wrA_reg_28(.CP(n_61635), .D(n_9596), .CD(n_60907), .Q(\wrA[28] 
		));
	notech_mux2 i_12988(.S(n_59977), .A(\wrA[28] ), .B(\addr_miss[28] ), .Z(n_9596
		));
	notech_nand2 i_79548(.A(n_953), .B(n_441), .Z(n_59690));
	notech_reg wrA_reg_29(.CP(n_61634), .D(n_9602), .CD(n_60906), .Q(\wrA[29] 
		));
	notech_mux2 i_12996(.S(n_59977), .A(\wrA[29] ), .B(\addr_miss[29] ), .Z(n_9602
		));
	notech_nand2 i_79551(.A(n_952), .B(n_442), .Z(n_59696));
	notech_reg wrA_reg_30(.CP(n_61634), .D(n_9608), .CD(n_60906), .Q(\wrA[30] 
		));
	notech_mux2 i_13004(.S(n_59977), .A(\wrA[30] ), .B(\addr_miss[30] ), .Z(n_9608
		));
	notech_nand2 i_79554(.A(n_951), .B(n_443), .Z(n_59702));
	notech_reg wrA_reg_31(.CP(n_61634), .D(n_9614), .CD(n_60906), .Q(\wrA[31] 
		));
	notech_mux2 i_13012(.S(n_59977), .A(\wrA[31] ), .B(\addr_miss[31] ), .Z(n_9614
		));
	notech_ao4 i_79933(.A(n_912), .B(n_9983), .C(n_896), .D(\nnx_tab2[0] ), 
		.Z(n_59976));
	notech_reg wrD_reg_0(.CP(n_61634), .D(n_9620), .CD(n_60906), .Q(\wrD[0] 
		));
	notech_mux2 i_13020(.S(n_59977), .A(\wrD[0] ), .B(n_58573), .Z(n_9620)
		);
	notech_ao4 i_79936(.A(n_912), .B(n_9985), .C(n_896), .D(n_499), .Z(n_59982
		));
	notech_reg wrD_reg_1(.CP(n_61634), .D(n_9626), .CD(n_60906), .Q(\wrD[1] 
		));
	notech_mux2 i_13028(.S(n_59983), .A(\wrD[1] ), .B(data_miss[1]), .Z(n_9626
		));
	notech_ao4 i_79947(.A(n_896), .B(n_9978), .C(n_487), .D(n_916), .Z(n_60001
		));
	notech_reg wrD_reg_2(.CP(n_61634), .D(n_9632), .CD(n_60906), .Q(\wrD[2] 
		));
	notech_mux2 i_13036(.S(n_59977), .A(\wrD[2] ), .B(data_miss[2]), .Z(n_9632
		));
	notech_ao4 i_79950(.A(n_896), .B(n_9980), .C(n_492), .D(n_917), .Z(n_60007
		));
	notech_reg wrD_reg_3(.CP(n_61634), .D(n_9638), .CD(n_60906), .Q(\wrD[3] 
		));
	notech_mux2 i_13044(.S(n_59977), .A(\wrD[3] ), .B(data_miss[3]), .Z(n_9638
		));
	notech_nand3 i_80090(.A(n_890), .B(n_61563), .C(n_10175), .Z(n_56940));
	notech_reg wrD_reg_4(.CP(n_61634), .D(n_9644), .CD(n_60906), .Q(\wrD[4] 
		));
	notech_mux2 i_13052(.S(n_59977), .A(\wrD[4] ), .B(data_miss[4]), .Z(n_9644
		));
	notech_nand3 i_80092(.A(n_890), .B(n_61563), .C(n_10174), .Z(n_56946));
	notech_reg wrD_reg_5(.CP(n_61634), .D(n_9650), .CD(n_60906), .Q(\wrD[5] 
		));
	notech_mux2 i_13060(.S(n_59977), .A(\wrD[5] ), .B(n_58573), .Z(n_9650)
		);
	notech_nand3 i_80094(.A(n_890), .B(n_61563), .C(n_10173), .Z(n_56952));
	notech_reg wrD_reg_6(.CP(n_61634), .D(n_9656), .CD(n_60906), .Q(\wrD[6] 
		));
	notech_mux2 i_13068(.S(n_59977), .A(\wrD[6] ), .B(data_miss[6]), .Z(n_9656
		));
	notech_nand3 i_80096(.A(n_890), .B(n_61563), .C(n_10172), .Z(n_56958));
	notech_reg wrD_reg_7(.CP(n_61634), .D(n_9662), .CD(n_60906), .Q(\wrD[7] 
		));
	notech_mux2 i_13076(.S(n_59977), .A(\wrD[7] ), .B(data_miss[7]), .Z(n_9662
		));
	notech_nand3 i_80100(.A(n_890), .B(n_61563), .C(n_10170), .Z(n_56970));
	notech_reg req_miss_reg(.CP(n_61634), .D(n_9668), .CD(n_60906), .Q(req_miss
		));
	notech_mux2 i_13084(.S(n_10103), .A(req_miss), .B(n_58550), .Z(n_9668)
		);
	notech_nand3 i_80102(.A(n_890), .B(n_61563), .C(n_10169), .Z(n_56976));
	notech_reg cr2_reg_0(.CP(n_61634), .D(n_9674), .CD(n_60906), .Q(cr2[0])
		);
	notech_mux2 i_13092(.S(n_808), .A(iDaddr_f[0]), .B(cr2[0]), .Z(n_9674)
		);
	notech_nand3 i_80104(.A(n_890), .B(n_61563), .C(n_10168), .Z(n_56982));
	notech_reg cr2_reg_1(.CP(n_61634), .D(n_9680), .CD(n_60906), .Q(cr2[1])
		);
	notech_mux2 i_13100(.S(n_808), .A(iDaddr_f[1]), .B(cr2[1]), .Z(n_9680)
		);
	notech_nand3 i_80106(.A(n_890), .B(n_61568), .C(n_10167), .Z(n_56988));
	notech_reg cr2_reg_2(.CP(n_61635), .D(n_9686), .CD(n_60907), .Q(cr2[2])
		);
	notech_mux2 i_13108(.S(n_808), .A(iDaddr_f[2]), .B(cr2[2]), .Z(n_9686)
		);
	notech_nand3 i_80108(.A(n_890), .B(n_61568), .C(n_10166), .Z(n_56994));
	notech_reg cr2_reg_3(.CP(n_61640), .D(n_9692), .CD(n_60912), .Q(cr2[3])
		);
	notech_mux2 i_13116(.S(n_808), .A(iDaddr_f[3]), .B(cr2[3]), .Z(n_9692)
		);
	notech_nao3 i_80110(.A(n_890), .B(n_61568), .C(data_miss[12]), .Z(n_57000
		));
	notech_reg cr2_reg_4(.CP(n_61644), .D(n_9698), .CD(n_60916), .Q(cr2[4])
		);
	notech_mux2 i_13124(.S(n_808), .A(iDaddr_f[4]), .B(cr2[4]), .Z(n_9698)
		);
	notech_nao3 i_80112(.A(n_890), .B(n_61568), .C(data_miss[13]), .Z(n_57006
		));
	notech_reg cr2_reg_5(.CP(n_61644), .D(n_9704), .CD(n_60916), .Q(cr2[5])
		);
	notech_mux2 i_13132(.S(n_808), .A(iDaddr_f[5]), .B(cr2[5]), .Z(n_9704)
		);
	notech_nao3 i_80114(.A(n_890), .B(n_61568), .C(data_miss[14]), .Z(n_57012
		));
	notech_reg cr2_reg_6(.CP(n_61640), .D(n_9710), .CD(n_60912), .Q(cr2[6])
		);
	notech_mux2 i_13140(.S(n_808), .A(iDaddr_f[6]), .B(cr2[6]), .Z(n_9710)
		);
	notech_nao3 i_80116(.A(n_890), .B(n_61568), .C(data_miss[15]), .Z(n_57018
		));
	notech_reg cr2_reg_7(.CP(n_61640), .D(n_9716), .CD(n_60912), .Q(cr2[7])
		);
	notech_mux2 i_13148(.S(n_808), .A(iDaddr_f[7]), .B(cr2[7]), .Z(n_9716)
		);
	notech_nao3 i_80118(.A(n_60786), .B(n_61568), .C(data_miss[16]), .Z(n_57024
		));
	notech_reg cr2_reg_8(.CP(n_61640), .D(n_9722), .CD(n_60912), .Q(cr2[8])
		);
	notech_mux2 i_13156(.S(n_808), .A(iDaddr_f[8]), .B(cr2[8]), .Z(n_9722)
		);
	notech_nao3 i_80120(.A(n_60786), .B(n_61570), .C(data_miss[17]), .Z(n_57030
		));
	notech_reg cr2_reg_9(.CP(n_61640), .D(n_9728), .CD(n_60912), .Q(cr2[9])
		);
	notech_mux2 i_13164(.S(n_808), .A(iDaddr_f[9]), .B(cr2[9]), .Z(n_9728)
		);
	notech_nao3 i_80122(.A(n_60786), .B(n_61568), .C(data_miss[18]), .Z(n_57036
		));
	notech_reg cr2_reg_10(.CP(n_61644), .D(n_9734), .CD(n_60916), .Q(cr2[10]
		));
	notech_mux2 i_13172(.S(n_808), .A(iDaddr_f[10]), .B(cr2[10]), .Z(n_9734)
		);
	notech_nao3 i_80124(.A(n_60786), .B(n_61568), .C(data_miss[19]), .Z(n_57042
		));
	notech_reg cr2_reg_11(.CP(n_61644), .D(n_9740), .CD(n_60916), .Q(cr2[11]
		));
	notech_mux2 i_13180(.S(n_808), .A(iDaddr_f[11]), .B(cr2[11]), .Z(n_9740)
		);
	notech_nao3 i_80126(.A(n_60786), .B(n_61568), .C(data_miss[20]), .Z(n_57048
		));
	notech_reg cr2_reg_12(.CP(n_61644), .D(n_9746), .CD(n_60916), .Q(cr2[12]
		));
	notech_mux2 i_13188(.S(n_808), .A(iDaddr_f[12]), .B(cr2[12]), .Z(n_9746)
		);
	notech_nao3 i_80128(.A(n_60786), .B(n_61568), .C(data_miss[21]), .Z(n_57054
		));
	notech_reg cr2_reg_13(.CP(n_61644), .D(n_9752), .CD(n_60916), .Q(cr2[13]
		));
	notech_mux2 i_13196(.S(n_808), .A(iDaddr_f[13]), .B(cr2[13]), .Z(n_9752)
		);
	notech_nao3 i_80130(.A(n_60786), .B(n_61565), .C(data_miss[22]), .Z(n_57060
		));
	notech_reg cr2_reg_14(.CP(n_61644), .D(n_9758), .CD(n_60916), .Q(cr2[14]
		));
	notech_mux2 i_13204(.S(n_808), .A(iDaddr_f[14]), .B(cr2[14]), .Z(n_9758)
		);
	notech_nao3 i_80132(.A(n_60786), .B(n_61565), .C(data_miss[23]), .Z(n_57066
		));
	notech_reg cr2_reg_15(.CP(n_61644), .D(n_9764), .CD(n_60916), .Q(cr2[15]
		));
	notech_mux2 i_13212(.S(n_808), .A(iDaddr_f[15]), .B(cr2[15]), .Z(n_9764)
		);
	notech_nao3 i_80134(.A(n_60786), .B(n_61565), .C(data_miss[24]), .Z(n_57072
		));
	notech_reg cr2_reg_16(.CP(n_61644), .D(n_9770), .CD(n_60916), .Q(cr2[16]
		));
	notech_mux2 i_13220(.S(n_53568), .A(iDaddr_f[16]), .B(cr2[16]), .Z(n_9770
		));
	notech_nao3 i_80136(.A(n_60786), .B(n_61565), .C(data_miss[25]), .Z(n_57078
		));
	notech_reg cr2_reg_17(.CP(n_61640), .D(n_9776), .CD(n_60912), .Q(cr2[17]
		));
	notech_mux2 i_13228(.S(n_53568), .A(iDaddr_f[17]), .B(cr2[17]), .Z(n_9776
		));
	notech_nao3 i_80138(.A(n_60786), .B(n_61565), .C(data_miss[26]), .Z(n_57084
		));
	notech_reg cr2_reg_18(.CP(n_61640), .D(n_9782), .CD(n_60912), .Q(cr2[18]
		));
	notech_mux2 i_13236(.S(n_53568), .A(iDaddr_f[18]), .B(cr2[18]), .Z(n_9782
		));
	notech_nao3 i_80140(.A(n_890), .B(n_61565), .C(data_miss[27]), .Z(n_57090
		));
	notech_reg cr2_reg_19(.CP(n_61640), .D(n_9788), .CD(n_60912), .Q(cr2[19]
		));
	notech_mux2 i_13244(.S(n_53568), .A(iDaddr_f[19]), .B(cr2[19]), .Z(n_9788
		));
	notech_nao3 i_80142(.A(n_60786), .B(n_61568), .C(data_miss[28]), .Z(n_57096
		));
	notech_reg cr2_reg_20(.CP(n_61640), .D(n_9794), .CD(n_60912), .Q(cr2[20]
		));
	notech_mux2 i_13252(.S(n_53568), .A(iDaddr_f[20]), .B(cr2[20]), .Z(n_9794
		));
	notech_nao3 i_80144(.A(n_60786), .B(n_61568), .C(data_miss[29]), .Z(n_57102
		));
	notech_reg cr2_reg_21(.CP(n_61640), .D(n_9800), .CD(n_60912), .Q(cr2[21]
		));
	notech_mux2 i_13260(.S(n_53568), .A(iDaddr_f[21]), .B(cr2[21]), .Z(n_9800
		));
	notech_nao3 i_80146(.A(n_60786), .B(n_61568), .C(data_miss[30]), .Z(n_57108
		));
	notech_reg cr2_reg_22(.CP(n_61635), .D(n_9806), .CD(n_60907), .Q(cr2[22]
		));
	notech_mux2 i_13268(.S(n_53568), .A(iDaddr_f[22]), .B(cr2[22]), .Z(n_9806
		));
	notech_nao3 i_80148(.A(n_60786), .B(n_61568), .C(data_miss[31]), .Z(n_57114
		));
	notech_reg cr2_reg_23(.CP(n_61635), .D(n_9812), .CD(n_60907), .Q(cr2[23]
		));
	notech_mux2 i_13276(.S(n_53568), .A(iDaddr_f[23]), .B(cr2[23]), .Z(n_9812
		));
	notech_nand2 i_80154(.A(n_60786), .B(n_61568), .Z(n_57138));
	notech_reg cr2_reg_24(.CP(n_61640), .D(n_9818), .CD(n_60912), .Q(cr2[24]
		));
	notech_mux2 i_13284(.S(n_53568), .A(iDaddr_f[24]), .B(cr2[24]), .Z(n_9818
		));
	notech_ao4 i_80162(.A(n_912), .B(n_10033), .C(n_896), .D(\nnx_tab1[0] ),
		 .Z(n_57194));
	notech_reg cr2_reg_25(.CP(n_61640), .D(n_9824), .CD(n_60912), .Q(cr2[25]
		));
	notech_mux2 i_13292(.S(n_53568), .A(iDaddr_f[25]), .B(cr2[25]), .Z(n_9824
		));
	notech_ao4 i_80165(.A(n_912), .B(n_10035), .C(n_896), .D(n_478), .Z(n_57200
		));
	notech_reg cr2_reg_26(.CP(n_61640), .D(n_9830), .CD(n_60912), .Q(cr2[26]
		));
	notech_mux2 i_13300(.S(n_53568), .A(iDaddr_f[26]), .B(cr2[26]), .Z(n_9830
		));
	notech_ao4 i_80172(.A(n_896), .B(n_10028), .C(n_466), .D(n_926), .Z(n_58780
		));
	notech_reg cr2_reg_27(.CP(n_61640), .D(n_9836), .CD(n_60912), .Q(cr2[27]
		));
	notech_mux2 i_13308(.S(n_53568), .A(iDaddr_f[27]), .B(cr2[27]), .Z(n_9836
		));
	notech_ao4 i_80175(.A(n_896), .B(n_10030), .C(n_471), .D(n_927), .Z(n_58786
		));
	notech_reg cr2_reg_28(.CP(n_61640), .D(n_9842), .CD(n_60912), .Q(cr2[28]
		));
	notech_mux2 i_13316(.S(n_53568), .A(iDaddr_f[28]), .B(cr2[28]), .Z(n_9842
		));
	notech_nand3 i_43(.A(n_912), .B(n_935), .C(n_858), .Z(n_58532));
	notech_reg cr2_reg_29(.CP(n_61640), .D(n_9848), .CD(n_60912), .Q(cr2[29]
		));
	notech_mux2 i_13324(.S(n_53568), .A(iDaddr_f[29]), .B(cr2[29]), .Z(n_9848
		));
	notech_nand3 i_42(.A(n_938), .B(n_855), .C(n_937), .Z(n_58526));
	notech_reg cr2_reg_30(.CP(n_61640), .D(n_9854), .CD(n_60912), .Q(cr2[30]
		));
	notech_mux2 i_13332(.S(n_53568), .A(iDaddr_f[30]), .B(cr2[30]), .Z(n_9854
		));
	notech_mux2 i_41(.S(n_61579), .A(n_447), .B(n_445), .Z(n_58520));
	notech_reg cr2_reg_31(.CP(n_61640), .D(n_9860), .CD(n_60912), .Q(cr2[31]
		));
	notech_mux2 i_13340(.S(n_53568), .A(iDaddr_f[31]), .B(cr2[31]), .Z(n_9860
		));
	notech_inv i_14822(.A(n_985), .Z(n_9866));
	notech_inv i_14823(.A(n_459), .Z(n_9867));
	notech_inv i_14824(.A(n_901), .Z(n_9868));
	notech_inv i_14825(.A(n_889), .Z(n_9869));
	notech_inv i_14826(.A(n_883), .Z(n_9870));
	notech_inv i_14827(.A(\dir1[10] ), .Z(n_9871));
	notech_inv i_14828(.A(\dir1[11] ), .Z(n_9872));
	notech_inv i_14829(.A(\dir1[12] ), .Z(n_9873));
	notech_inv i_14830(.A(\dir1[13] ), .Z(n_9874));
	notech_inv i_14831(.A(\dir1[14] ), .Z(n_9875));
	notech_inv i_14832(.A(\dir1[15] ), .Z(n_9876));
	notech_inv i_14833(.A(\dir1[16] ), .Z(n_9877));
	notech_inv i_14834(.A(\dir1[17] ), .Z(n_9878));
	notech_inv i_14835(.A(\dir1[18] ), .Z(n_9879));
	notech_inv i_14836(.A(\dir1[19] ), .Z(n_9880));
	notech_inv i_14837(.A(\dir1[20] ), .Z(n_9881));
	notech_inv i_14838(.A(\dir1[21] ), .Z(n_9882));
	notech_inv i_14839(.A(\dir1[22] ), .Z(n_9883));
	notech_inv i_14840(.A(\dir1[23] ), .Z(n_9884));
	notech_inv i_14841(.A(\dir1[24] ), .Z(n_9885));
	notech_inv i_14842(.A(\dir1[25] ), .Z(n_9886));
	notech_inv i_14843(.A(\dir1[26] ), .Z(n_9887));
	notech_inv i_14844(.A(\dir1[27] ), .Z(n_9888));
	notech_inv i_14845(.A(\dir1[28] ), .Z(n_9889));
	notech_inv i_14846(.A(\dir1[29] ), .Z(n_9890));
	notech_inv i_14847(.A(\dir2[10] ), .Z(n_9891));
	notech_inv i_14848(.A(\dir2[11] ), .Z(n_9892));
	notech_inv i_14849(.A(\dir2[12] ), .Z(n_9893));
	notech_inv i_14850(.A(\dir2[13] ), .Z(n_9894));
	notech_inv i_14851(.A(\dir2[14] ), .Z(n_9895));
	notech_inv i_14852(.A(\dir2[15] ), .Z(n_9896));
	notech_inv i_14853(.A(\dir2[16] ), .Z(n_9897));
	notech_inv i_14854(.A(\dir2[17] ), .Z(n_9898));
	notech_inv i_14855(.A(\dir2[18] ), .Z(n_9899));
	notech_inv i_14856(.A(\dir2[19] ), .Z(n_9900));
	notech_inv i_14857(.A(\dir2[20] ), .Z(n_9901));
	notech_inv i_14858(.A(\dir2[21] ), .Z(n_9902));
	notech_inv i_14859(.A(\dir2[22] ), .Z(n_9903));
	notech_inv i_14860(.A(\dir2[23] ), .Z(n_9904));
	notech_inv i_14861(.A(\dir2[24] ), .Z(n_9905));
	notech_inv i_14862(.A(\dir2[25] ), .Z(n_9906));
	notech_inv i_14863(.A(\dir2[26] ), .Z(n_9907));
	notech_inv i_14864(.A(\dir2[27] ), .Z(n_9908));
	notech_inv i_14865(.A(\dir2[28] ), .Z(n_9909));
	notech_inv i_14866(.A(\dir2[29] ), .Z(n_9910));
	notech_inv i_14867(.A(n_476), .Z(n_9911));
	notech_inv i_14868(.A(\tab21[10] ), .Z(n_9912));
	notech_inv i_14869(.A(\tab21[11] ), .Z(n_9913));
	notech_inv i_14870(.A(\tab21[12] ), .Z(n_9914));
	notech_inv i_14871(.A(\tab21[13] ), .Z(n_9915));
	notech_inv i_14872(.A(\tab21[14] ), .Z(n_9916));
	notech_inv i_14873(.A(\tab21[15] ), .Z(n_9917));
	notech_inv i_14874(.A(\tab21[16] ), .Z(n_9918));
	notech_inv i_14875(.A(\tab21[17] ), .Z(n_9919));
	notech_inv i_14876(.A(\tab21[18] ), .Z(n_9920));
	notech_inv i_14877(.A(\tab21[19] ), .Z(n_9921));
	notech_inv i_14878(.A(\tab21[20] ), .Z(n_9922));
	notech_inv i_14879(.A(\tab21[21] ), .Z(n_9923));
	notech_inv i_14880(.A(\tab21[22] ), .Z(n_9924));
	notech_inv i_14881(.A(\tab21[23] ), .Z(n_9925));
	notech_inv i_14882(.A(n_497), .Z(n_9926));
	notech_inv i_14883(.A(\tab21[24] ), .Z(n_9927));
	notech_inv i_14884(.A(\tab21[25] ), .Z(n_9928));
	notech_inv i_14885(.A(\tab21[26] ), .Z(n_9929));
	notech_inv i_14886(.A(\tab21[27] ), .Z(n_9930));
	notech_inv i_14887(.A(\tab21[28] ), .Z(n_9931));
	notech_inv i_14888(.A(\tab21[29] ), .Z(n_9932));
	notech_inv i_14889(.A(\tab23[10] ), .Z(n_9933));
	notech_inv i_14890(.A(\tab23[11] ), .Z(n_9934));
	notech_inv i_14891(.A(\tab23[12] ), .Z(n_9935));
	notech_inv i_14892(.A(\tab23[13] ), .Z(n_9936));
	notech_inv i_14893(.A(\tab23[14] ), .Z(n_9937));
	notech_inv i_14894(.A(\tab23[15] ), .Z(n_9938));
	notech_inv i_14895(.A(\tab23[16] ), .Z(n_9939));
	notech_inv i_14896(.A(n_553), .Z(n_9940));
	notech_inv i_14897(.A(\tab23[17] ), .Z(n_9941));
	notech_inv i_14898(.A(\tab23[18] ), .Z(n_9942));
	notech_inv i_14899(.A(\tab23[19] ), .Z(n_9943));
	notech_inv i_14900(.A(\tab23[20] ), .Z(n_9944));
	notech_inv i_14901(.A(n_557), .Z(n_9945));
	notech_inv i_14902(.A(\tab23[21] ), .Z(n_9946));
	notech_inv i_14903(.A(\tab23[22] ), .Z(n_9947));
	notech_inv i_14904(.A(n_559), .Z(n_9948));
	notech_inv i_14905(.A(\tab23[23] ), .Z(n_9949));
	notech_inv i_14906(.A(\tab23[24] ), .Z(n_9950));
	notech_inv i_14907(.A(\tab23[25] ), .Z(n_9951));
	notech_inv i_14908(.A(\tab23[26] ), .Z(n_9952));
	notech_inv i_14909(.A(\tab23[27] ), .Z(n_9953));
	notech_inv i_14910(.A(\tab23[28] ), .Z(n_9954));
	notech_inv i_14911(.A(\tab23[29] ), .Z(n_9955));
	notech_inv i_14912(.A(hit_adr23), .Z(n_9956));
	notech_inv i_14913(.A(\tab24[10] ), .Z(n_9957));
	notech_inv i_14914(.A(\tab24[11] ), .Z(n_9958));
	notech_inv i_14915(.A(\tab24[12] ), .Z(n_9959));
	notech_inv i_14916(.A(\tab24[13] ), .Z(n_9960));
	notech_inv i_14917(.A(\tab24[14] ), .Z(n_9961));
	notech_inv i_14918(.A(\tab24[15] ), .Z(n_9962));
	notech_inv i_14919(.A(\tab24[16] ), .Z(n_9963));
	notech_inv i_14920(.A(\tab24[17] ), .Z(n_9964));
	notech_inv i_14921(.A(\tab24[18] ), .Z(n_9965));
	notech_inv i_14922(.A(\tab24[19] ), .Z(n_9966));
	notech_inv i_14923(.A(\tab24[20] ), .Z(n_9967));
	notech_inv i_14924(.A(\tab24[21] ), .Z(n_9968));
	notech_inv i_14925(.A(\tab24[22] ), .Z(n_9969));
	notech_inv i_14926(.A(\tab24[23] ), .Z(n_9970));
	notech_inv i_14927(.A(\tab24[24] ), .Z(n_9971));
	notech_inv i_14928(.A(\tab24[25] ), .Z(n_9972));
	notech_inv i_14929(.A(\tab24[26] ), .Z(n_9973));
	notech_inv i_14930(.A(\tab24[27] ), .Z(n_9974));
	notech_inv i_14931(.A(\tab24[28] ), .Z(n_9975));
	notech_inv i_14932(.A(\tab24[29] ), .Z(n_9976));
	notech_inv i_14933(.A(n_59976), .Z(n_9977));
	notech_inv i_14934(.A(\nnx_tab2[0] ), .Z(n_9978));
	notech_inv i_14935(.A(n_59982), .Z(n_9979));
	notech_inv i_14936(.A(\nnx_tab2[1] ), .Z(n_9980));
	notech_inv i_14937(.A(\nbus_14515[0] ), .Z(n_9981));
	notech_inv i_14938(.A(n_60001), .Z(n_9982));
	notech_inv i_14939(.A(\nx_tab2[0] ), .Z(n_9983));
	notech_inv i_14940(.A(n_60007), .Z(n_9984));
	notech_inv i_14941(.A(\nx_tab2[1] ), .Z(n_9985));
	notech_inv i_14942(.A(\tab12[10] ), .Z(n_9986));
	notech_inv i_14943(.A(\tab12[11] ), .Z(n_9987));
	notech_inv i_14944(.A(\tab12[12] ), .Z(n_9988));
	notech_inv i_14945(.A(\tab12[13] ), .Z(n_9989));
	notech_inv i_14946(.A(\tab12[14] ), .Z(n_9990));
	notech_inv i_14947(.A(\tab12[15] ), .Z(n_9991));
	notech_inv i_14948(.A(\tab12[16] ), .Z(n_9992));
	notech_inv i_14949(.A(\tab12[17] ), .Z(n_9993));
	notech_inv i_14950(.A(\tab12[18] ), .Z(n_9994));
	notech_inv i_14951(.A(\tab12[19] ), .Z(n_9995));
	notech_inv i_14952(.A(\tab12[20] ), .Z(n_9996));
	notech_inv i_14953(.A(\tab12[21] ), .Z(n_9997));
	notech_inv i_14954(.A(\tab12[22] ), .Z(n_9998));
	notech_inv i_14955(.A(\tab12[23] ), .Z(n_9999));
	notech_inv i_14956(.A(\tab12[24] ), .Z(n_10000));
	notech_inv i_14957(.A(\tab12[25] ), .Z(n_10001));
	notech_inv i_14958(.A(\tab12[26] ), .Z(n_10002));
	notech_inv i_14959(.A(\tab12[27] ), .Z(n_10003));
	notech_inv i_14960(.A(\tab12[28] ), .Z(n_10004));
	notech_inv i_14961(.A(\tab12[29] ), .Z(n_10005));
	notech_inv i_14962(.A(hit_adr13), .Z(n_10006));
	notech_inv i_14963(.A(\tab14[10] ), .Z(n_10007));
	notech_inv i_14964(.A(\tab14[11] ), .Z(n_10008));
	notech_inv i_14965(.A(\tab14[12] ), .Z(n_10009));
	notech_inv i_14966(.A(\tab14[13] ), .Z(n_10010));
	notech_inv i_14967(.A(\tab14[14] ), .Z(n_10011));
	notech_inv i_14968(.A(\tab14[15] ), .Z(n_10012));
	notech_inv i_14969(.A(\tab14[16] ), .Z(n_10013));
	notech_inv i_14970(.A(\tab14[17] ), .Z(n_10014));
	notech_inv i_14971(.A(\tab14[18] ), .Z(n_10015));
	notech_inv i_14972(.A(\tab14[19] ), .Z(n_10016));
	notech_inv i_14973(.A(\tab14[20] ), .Z(n_10017));
	notech_inv i_14974(.A(\tab14[21] ), .Z(n_10018));
	notech_inv i_14975(.A(\tab14[22] ), .Z(n_10019));
	notech_inv i_14976(.A(\tab14[23] ), .Z(n_10020));
	notech_inv i_14977(.A(\tab14[24] ), .Z(n_10021));
	notech_inv i_14978(.A(\tab14[25] ), .Z(n_10022));
	notech_inv i_14979(.A(\tab14[26] ), .Z(n_10023));
	notech_inv i_14980(.A(\tab14[27] ), .Z(n_10024));
	notech_inv i_14981(.A(\tab14[28] ), .Z(n_10025));
	notech_inv i_14982(.A(\tab14[29] ), .Z(n_10026));
	notech_inv i_14983(.A(n_57194), .Z(n_10027));
	notech_inv i_14984(.A(\nnx_tab1[0] ), .Z(n_10028));
	notech_inv i_14985(.A(n_57200), .Z(n_10029));
	notech_inv i_14986(.A(\nnx_tab1[1] ), .Z(n_10030));
	notech_inv i_14987(.A(\nbus_14490[0] ), .Z(n_10031));
	notech_inv i_14988(.A(n_58780), .Z(n_10032));
	notech_inv i_14989(.A(\nx_tab1[0] ), .Z(n_10033));
	notech_inv i_14990(.A(n_58786), .Z(n_10034));
	notech_inv i_14991(.A(\nx_tab1[1] ), .Z(n_10035));
	notech_inv i_14992(.A(\tab11[10] ), .Z(n_10036));
	notech_inv i_14993(.A(\tab11[11] ), .Z(n_10037));
	notech_inv i_14994(.A(\tab11[12] ), .Z(n_10038));
	notech_inv i_14995(.A(\tab11[13] ), .Z(n_10039));
	notech_inv i_14996(.A(\tab11[14] ), .Z(n_10040));
	notech_inv i_14997(.A(\tab11[15] ), .Z(n_10041));
	notech_inv i_14998(.A(\tab11[16] ), .Z(n_10042));
	notech_inv i_14999(.A(\tab11[17] ), .Z(n_10043));
	notech_inv i_15000(.A(\tab11[18] ), .Z(n_10044));
	notech_inv i_15001(.A(\tab11[19] ), .Z(n_10045));
	notech_inv i_15002(.A(\tab11[20] ), .Z(n_10046));
	notech_inv i_15003(.A(\tab11[21] ), .Z(n_10047));
	notech_inv i_15004(.A(\tab11[22] ), .Z(n_10048));
	notech_inv i_15005(.A(\tab11[23] ), .Z(n_10049));
	notech_inv i_15006(.A(\tab11[24] ), .Z(n_10050));
	notech_inv i_15007(.A(\tab11[25] ), .Z(n_10051));
	notech_inv i_15008(.A(\tab11[26] ), .Z(n_10052));
	notech_inv i_15009(.A(\tab11[27] ), .Z(n_10053));
	notech_inv i_15010(.A(\tab11[28] ), .Z(n_10054));
	notech_inv i_15011(.A(\tab11[29] ), .Z(n_10055));
	notech_inv i_15012(.A(n_59950), .Z(n_10056));
	notech_inv i_15013(.A(n_61579), .Z(n_10057));
	notech_inv i_15014(.A(fsm[3]), .Z(n_10058));
	notech_inv i_15015(.A(n_59528), .Z(n_10059));
	notech_inv i_15016(.A(n_59534), .Z(n_10060));
	notech_inv i_15017(.A(n_59540), .Z(n_10061));
	notech_inv i_15018(.A(n_59546), .Z(n_10062));
	notech_inv i_15019(.A(n_59552), .Z(n_10063));
	notech_inv i_15020(.A(n_59558), .Z(n_10064));
	notech_inv i_15021(.A(n_59564), .Z(n_10065));
	notech_inv i_15022(.A(n_59570), .Z(n_10066));
	notech_inv i_15023(.A(n_59576), .Z(n_10067));
	notech_inv i_15024(.A(n_59582), .Z(n_10068));
	notech_inv i_15025(.A(\addr_miss[2] ), .Z(n_10069));
	notech_inv i_15026(.A(\addr_miss[3] ), .Z(n_10070));
	notech_inv i_15027(.A(\addr_miss[4] ), .Z(n_10071));
	notech_inv i_15028(.A(\addr_miss[5] ), .Z(n_10072));
	notech_inv i_15029(.A(\addr_miss[6] ), .Z(n_10073));
	notech_inv i_15030(.A(\addr_miss[7] ), .Z(n_10074));
	notech_inv i_15031(.A(\addr_miss[8] ), .Z(n_10075));
	notech_inv i_15032(.A(\addr_miss[9] ), .Z(n_10076));
	notech_inv i_15033(.A(\addr_miss[10] ), .Z(n_10077));
	notech_inv i_15034(.A(\addr_miss[11] ), .Z(n_10078));
	notech_inv i_15035(.A(\wrA[12] ), .Z(n_10079));
	notech_inv i_15036(.A(\wrA[13] ), .Z(n_10080));
	notech_inv i_15037(.A(\wrA[14] ), .Z(n_10081));
	notech_inv i_15038(.A(\wrA[15] ), .Z(n_10082));
	notech_inv i_15039(.A(\wrA[16] ), .Z(n_10083));
	notech_inv i_15040(.A(\wrA[17] ), .Z(n_10084));
	notech_inv i_15041(.A(\wrA[18] ), .Z(n_10085));
	notech_inv i_15042(.A(\wrA[19] ), .Z(n_10086));
	notech_inv i_15043(.A(\wrA[20] ), .Z(n_10087));
	notech_inv i_15044(.A(\wrA[21] ), .Z(n_10088));
	notech_inv i_15045(.A(\wrA[22] ), .Z(n_10089));
	notech_inv i_15046(.A(\wrA[23] ), .Z(n_10090));
	notech_inv i_15047(.A(\wrA[24] ), .Z(n_10091));
	notech_inv i_15048(.A(\wrA[25] ), .Z(n_10092));
	notech_inv i_15049(.A(\wrA[26] ), .Z(n_10093));
	notech_inv i_15050(.A(\wrA[27] ), .Z(n_10094));
	notech_inv i_15051(.A(\wrA[28] ), .Z(n_10095));
	notech_inv i_15052(.A(\wrA[29] ), .Z(n_10096));
	notech_inv i_15053(.A(\wrA[30] ), .Z(n_10097));
	notech_inv i_15054(.A(\wrA[31] ), .Z(n_10098));
	notech_inv i_15055(.A(n_58573), .Z(n_10099));
	notech_inv i_15057(.A(n_58550), .Z(n_10101));
	notech_inv i_15058(.A(req_miss), .Z(n_10102));
	notech_inv i_15059(.A(n_58547), .Z(n_10103));
	notech_inv i_15060(.A(addr_phys_3197023), .Z(addr_phys[31]));
	notech_inv i_15061(.A(addr_phys_3097022), .Z(addr_phys[30]));
	notech_inv i_15062(.A(addr_phys_2997021), .Z(addr_phys[29]));
	notech_inv i_15063(.A(addr_phys_2897020), .Z(addr_phys[28]));
	notech_inv i_15064(.A(addr_phys_2797019), .Z(addr_phys[27]));
	notech_inv i_15065(.A(addr_phys_2697018), .Z(addr_phys[26]));
	notech_inv i_15066(.A(addr_phys_2597017), .Z(addr_phys[25]));
	notech_inv i_15067(.A(addr_phys_2497016), .Z(addr_phys[24]));
	notech_inv i_15068(.A(addr_phys_2397015), .Z(addr_phys[23]));
	notech_inv i_15069(.A(addr_phys_2297014), .Z(addr_phys[22]));
	notech_inv i_15070(.A(addr_phys_2197013), .Z(addr_phys[21]));
	notech_inv i_15071(.A(addr_phys_2097012), .Z(addr_phys[20]));
	notech_inv i_15072(.A(addr_phys_1997011), .Z(addr_phys[19]));
	notech_inv i_15073(.A(addr_phys_1897010), .Z(addr_phys[18]));
	notech_inv i_15074(.A(addr_phys_1797009), .Z(addr_phys[17]));
	notech_inv i_15075(.A(addr_phys_1697008), .Z(addr_phys[16]));
	notech_inv i_15076(.A(addr_phys_1597007), .Z(addr_phys[15]));
	notech_inv i_15077(.A(addr_phys_1497006), .Z(addr_phys[14]));
	notech_inv i_15078(.A(addr_phys_1397005), .Z(addr_phys[13]));
	notech_inv i_15079(.A(addr_phys_1297004), .Z(addr_phys[12]));
	notech_inv i_15080(.A(n_60432), .Z(n_10124));
	notech_inv i_15081(.A(iDaddr[2]), .Z(n_10125));
	notech_inv i_15082(.A(iDaddr[3]), .Z(n_10126));
	notech_inv i_15083(.A(iDaddr[4]), .Z(n_10127));
	notech_inv i_15084(.A(iDaddr[5]), .Z(n_10128));
	notech_inv i_15085(.A(iDaddr[6]), .Z(n_10129));
	notech_inv i_15086(.A(iDaddr[7]), .Z(n_10130));
	notech_inv i_15087(.A(iDaddr[8]), .Z(n_10131));
	notech_inv i_15088(.A(iDaddr[9]), .Z(n_10132));
	notech_inv i_15089(.A(iDaddr[10]), .Z(n_10133));
	notech_inv i_15090(.A(iDaddr[11]), .Z(n_10134));
	notech_inv i_15091(.A(iDaddr[12]), .Z(n_10135));
	notech_inv i_15092(.A(iDaddr[13]), .Z(n_10136));
	notech_inv i_15093(.A(iDaddr[14]), .Z(n_10137));
	notech_inv i_15094(.A(iDaddr[15]), .Z(n_10138));
	notech_inv i_15095(.A(iDaddr[16]), .Z(n_10139));
	notech_inv i_15096(.A(iDaddr[17]), .Z(n_10140));
	notech_inv i_15097(.A(iDaddr[18]), .Z(n_10141));
	notech_inv i_15098(.A(iDaddr[19]), .Z(n_10142));
	notech_inv i_15099(.A(iDaddr[20]), .Z(n_10143));
	notech_inv i_15100(.A(iDaddr[21]), .Z(n_10144));
	notech_inv i_15101(.A(iDaddr[22]), .Z(n_10145));
	notech_inv i_15102(.A(iDaddr[23]), .Z(n_10146));
	notech_inv i_15103(.A(iDaddr[24]), .Z(n_10147));
	notech_inv i_15104(.A(iDaddr[25]), .Z(n_10148));
	notech_inv i_15105(.A(iDaddr[26]), .Z(n_10149));
	notech_inv i_15106(.A(iDaddr[27]), .Z(n_10150));
	notech_inv i_15107(.A(iDaddr[28]), .Z(n_10151));
	notech_inv i_15108(.A(iDaddr[29]), .Z(n_10152));
	notech_inv i_15109(.A(iDaddr[30]), .Z(n_10153));
	notech_inv i_15110(.A(iDaddr[31]), .Z(n_10154));
	notech_inv i_15111(.A(n_61534), .Z(owrite_req));
	notech_inv i_15112(.A(\dir1_0[9] ), .Z(n_10156));
	notech_inv i_15113(.A(\dir1_0[8] ), .Z(n_10157));
	notech_inv i_15114(.A(\dir1_0[7] ), .Z(n_10158));
	notech_inv i_15115(.A(\dir1_0[6] ), .Z(n_10159));
	notech_inv i_15116(.A(\dir1_0[5] ), .Z(n_10160));
	notech_inv i_15117(.A(\dir1_0[4] ), .Z(n_10161));
	notech_inv i_15118(.A(\dir1_0[3] ), .Z(n_10162));
	notech_inv i_15119(.A(\dir1_0[2] ), .Z(n_10163));
	notech_inv i_15120(.A(\dir1_0[1] ), .Z(n_10164));
	notech_inv i_15121(.A(\dir1_0[0] ), .Z(n_10165));
	notech_inv i_15122(.A(\tab11_0[9] ), .Z(n_10166));
	notech_inv i_15123(.A(\tab11_0[8] ), .Z(n_10167));
	notech_inv i_15124(.A(\tab11_0[7] ), .Z(n_10168));
	notech_inv i_15125(.A(\tab11_0[6] ), .Z(n_10169));
	notech_inv i_15126(.A(\tab11_0[5] ), .Z(n_10170));
	notech_inv i_15127(.A(\tab11_0[4] ), .Z(n_10171));
	notech_inv i_15128(.A(\tab11_0[3] ), .Z(n_10172));
	notech_inv i_15129(.A(\tab11_0[2] ), .Z(n_10173));
	notech_inv i_15130(.A(\tab11_0[1] ), .Z(n_10174));
	notech_inv i_15131(.A(\tab11_0[0] ), .Z(n_10175));
	notech_inv i_15132(.A(oread_req97003), .Z(oread_req));
	notech_inv i_15133(.A(hit_tab21), .Z(n_10177));
	notech_inv i_15134(.A(hit_tab23), .Z(n_10178));
	notech_inv i_15135(.A(hit_tab12), .Z(n_10179));
	notech_inv i_15136(.A(\hit_dir1[7] ), .Z(n_10180));
	notech_inv i_15137(.A(n_61594), .Z(n_10181));
	notech_inv i_15138(.A(iread_req), .Z(n_10182));
	notech_inv i_15139(.A(hit_dir2), .Z(n_10183));
	notech_inv i_15140(.A(pg_fault), .Z(n_10184));
	cmp14_19 t11(.ina({\tab11[33] , UNCONNECTED_000, UNCONNECTED_001, 
		UNCONNECTED_002, \tab11[9] , \tab11[8] , \tab11[7] , \tab11[6] ,
		 \tab11[5] , \tab11[4] , \tab11[3] , \tab11[2] , \tab11[1] , \tab11[0] 
		}), .inb({UNCONNECTED_003, UNCONNECTED_004, UNCONNECTED_005, 
		UNCONNECTED_006, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab11), .out2(hit_add11));
	cmp14_18 t14(.ina({\tab14[33] , UNCONNECTED_007, UNCONNECTED_008, 
		UNCONNECTED_009, \tab14[9] , \tab14[8] , \tab14[7] , \tab14[6] ,
		 \tab14[5] , \tab14[4] , \tab14[3] , \tab14[2] , \tab14[1] , \tab14[0] 
		}), .inb({UNCONNECTED_010, UNCONNECTED_011, UNCONNECTED_012, 
		UNCONNECTED_013, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab14), .out2(hit_add14));
	cmp14_17 t13(.ina({\tab13[33] , UNCONNECTED_014, UNCONNECTED_015, 
		UNCONNECTED_016, \tab13[9] , \tab13[8] , \tab13[7] , \tab13[6] ,
		 \tab13[5] , \tab13[4] , \tab13[3] , \tab13[2] , \tab13[1] , \tab13[0] 
		}), .inb({UNCONNECTED_017, UNCONNECTED_018, UNCONNECTED_019, 
		UNCONNECTED_020, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab13), .out2(hit_add13));
	cmp14_16 t12(.ina({\tab12[33] , UNCONNECTED_021, UNCONNECTED_022, 
		UNCONNECTED_023, \tab12[9] , \tab12[8] , \tab12[7] , \tab12[6] ,
		 \tab12[5] , \tab12[4] , \tab12[3] , \tab12[2] , \tab12[1] , \tab12[0] 
		}), .inb({UNCONNECTED_024, UNCONNECTED_025, UNCONNECTED_026, 
		UNCONNECTED_027, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab12), .out2(hit_add12));
	cmp14_15 t24(.ina({\tab24[33] , UNCONNECTED_028, UNCONNECTED_029, 
		UNCONNECTED_030, \tab24[9] , \tab24[8] , \tab24[7] , \tab24[6] ,
		 \tab24[5] , \tab24[4] , \tab24[3] , \tab24[2] , \tab24[1] , \tab24[0] 
		}), .inb({UNCONNECTED_031, UNCONNECTED_032, UNCONNECTED_033, 
		UNCONNECTED_034, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab24), .out2(hit_add24));
	cmp14_14 t23(.ina({\tab23[33] , UNCONNECTED_035, UNCONNECTED_036, 
		UNCONNECTED_037, \tab23[9] , \tab23[8] , \tab23[7] , \tab23[6] ,
		 \tab23[5] , \tab23[4] , \tab23[3] , \tab23[2] , \tab23[1] , \tab23[0] 
		}), .inb({UNCONNECTED_038, UNCONNECTED_039, UNCONNECTED_040, 
		UNCONNECTED_041, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab23), .out2(hit_add23));
	cmp14_13 t22(.ina({\tab22[33] , UNCONNECTED_042, UNCONNECTED_043, 
		UNCONNECTED_044, \tab22[9] , \tab22[8] , \tab22[7] , \tab22[6] ,
		 \tab22[5] , \tab22[4] , \tab22[3] , \tab22[2] , \tab22[1] , \tab22[0] 
		}), .inb({UNCONNECTED_045, UNCONNECTED_046, UNCONNECTED_047, 
		UNCONNECTED_048, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab22), .out2(hit_add22));
	cmp14_12 t21(.ina({\tab21[33] , UNCONNECTED_049, UNCONNECTED_050, 
		UNCONNECTED_051, \tab21[9] , \tab21[8] , \tab21[7] , \tab21[6] ,
		 \tab21[5] , \tab21[4] , \tab21[3] , \tab21[2] , \tab21[1] , \tab21[0] 
		}), .inb({UNCONNECTED_052, UNCONNECTED_053, UNCONNECTED_054, 
		UNCONNECTED_055, \tab11_0[9] , \tab11_0[8] , \tab11_0[7] , \tab11_0[6] 
		, \tab11_0[5] , \tab11_0[4] , \tab11_0[3] , \tab11_0[2] , \tab11_0[1] 
		, \tab11_0[0] }), .out(hit_tab21), .out2(hit_add21));
	cmp14_11 d2(.ina({\dir2[33] , UNCONNECTED_056, UNCONNECTED_057, 
		UNCONNECTED_058, \dir2[9] , \dir2[8] , \dir2[7] , \dir2[6] , \dir2[5] 
		, \dir2[4] , \dir2[3] , \dir2[2] , \dir2[1] , \dir2[0] }), .inb(
		{UNCONNECTED_059, UNCONNECTED_060, UNCONNECTED_061, 
		UNCONNECTED_062, \dir1_0[9] , \dir1_0[8] , \dir1_0[7] , \dir1_0[6] 
		, \dir1_0[5] , \dir1_0[4] , \dir1_0[3] , \dir1_0[2] , \dir1_0[1] 
		, \dir1_0[0] }), .out(hit_dir2));
	cmp14_10 d1(.ina({\dir1[33] , UNCONNECTED_063, UNCONNECTED_064, 
		UNCONNECTED_065, \dir1[9] , \dir1[8] , \dir1[7] , \dir1[6] , \dir1[5] 
		, \dir1[4] , \dir1[3] , \dir1[2] , \dir1[1] , \dir1[0] }), .inb(
		{UNCONNECTED_066, UNCONNECTED_067, UNCONNECTED_068, 
		UNCONNECTED_069, \dir1_0[9] , \dir1_0[8] , \dir1_0[7] , \dir1_0[6] 
		, \dir1_0[5] , \dir1_0[4] , \dir1_0[3] , \dir1_0[2] , \dir1_0[1] 
		, \dir1_0[0] }), .out(\hit_dir1[7] ));
	AWDP_INC_27 i_79020(.O0(fsm5_cnt_0), .fsm5_cnt(fsm5_cnt));
endmodule
module AWDP_partition_1(O0, mod_dec, sib_dec, displc, imm_sz, pfx_sz, twobyte, fpu);
    output [5:0] O0;
    input  mod_dec;
    input  sib_dec;
    input [2:0] displc;
    input [2:0] imm_sz;
    input [4:0] pfx_sz;
    input  twobyte;
    input  fpu;
    // Line 404
    wire [6:0] N18;
    // Line 404
    wire [5:0] N26;
    // Line 211
    wire [5:0] O0;
    // Line 404
    wire [7:0] N21;
    // Line 405
    wire [5:0] N16;

    // Line 404
    assign N18 = N16 + 7'h1 + mod_dec;
    // Line 404
    assign N26 = N21 + imm_sz;
    // Line 211
    assign O0 = N26;
    // Line 404
    assign N21 = N18 + displc + sib_dec;
    // Line 405
    assign N16 = pfx_sz + twobyte + fpu;
endmodule

module deco8(in8, indic);

	input [7:0] in8;
	output [72:0] indic;

	wire \indic[10] ;
	wire \indic[14] ;
	wire \indic[15] ;
	wire \indic[22] ;
	wire \indic[0] ;
	wire \indic[1] ;
	wire \indic[2] ;
	wire \indic[3] ;
	wire \indic[4] ;
	wire \indic[5] ;
	wire \indic[6] ;
	wire \indic[7] ;
	wire \indic[8] ;
	wire \indic[9] ;
	wire \indic[11] ;
	wire \indic[12] ;
	wire \indic[13] ;
	wire \indic[16] ;
	wire \indic[17] ;
	wire \indic[18] ;
	wire \indic[19] ;
	wire \indic[20] ;
	wire \indic[21] ;
	wire \indic[23] ;
	wire \indic[24] ;
	wire \indic[25] ;
	wire \indic[26] ;
	wire \indic[27] ;
	wire \indic[28] ;
	wire \indic[29] ;
	wire \indic[30] ;
	wire \indic[32] ;
	wire \indic[33] ;
	wire \indic[34] ;
	wire \indic[35] ;
	wire \indic[36] ;
	wire \indic[37] ;
	wire \indic[38] ;
	wire \indic[39] ;
	wire \indic[40] ;
	wire \indic[41] ;
	wire \indic[42] ;
	wire \indic[43] ;
	wire \indic[44] ;
	wire \indic[45] ;
	wire \indic[46] ;
	wire \indic[47] ;
	wire \indic[48] ;
	wire \indic[49] ;
	wire \indic[50] ;
	wire \indic[51] ;
	wire \indic[53] ;
	wire \indic[54] ;
	wire \indic[55] ;
	wire \indic[56] ;
	wire \indic[57] ;
	wire \indic[58] ;
	wire \indic[59] ;
	wire \indic[60] ;
	wire \indic[61] ;
	wire \indic[62] ;
	wire \indic[63] ;
	wire \indic[64] ;
	wire \indic[67] ;
	wire \indic[68] ;
	wire \indic[69] ;
	wire \indic[70] ;
	wire \indic[71] ;
	wire \indic[72] ;


	assign indic[10] = \indic[10] ;
	assign indic[14] = \indic[14] ;
	assign indic[15] = \indic[15] ;
	assign indic[22] = \indic[22] ;
	assign indic[0] = \indic[0] ;
	assign indic[1] = \indic[1] ;
	assign indic[2] = \indic[2] ;
	assign indic[3] = \indic[3] ;
	assign indic[4] = \indic[4] ;
	assign indic[5] = \indic[5] ;
	assign indic[6] = \indic[6] ;
	assign indic[7] = \indic[7] ;
	assign indic[8] = \indic[8] ;
	assign indic[9] = \indic[9] ;
	assign indic[11] = \indic[11] ;
	assign indic[12] = \indic[12] ;
	assign indic[13] = \indic[13] ;
	assign indic[16] = \indic[16] ;
	assign indic[17] = \indic[17] ;
	assign indic[18] = \indic[18] ;
	assign indic[19] = \indic[19] ;
	assign indic[20] = \indic[20] ;
	assign indic[21] = \indic[21] ;
	assign indic[23] = \indic[23] ;
	assign indic[24] = \indic[24] ;
	assign indic[25] = \indic[25] ;
	assign indic[26] = \indic[26] ;
	assign indic[27] = \indic[27] ;
	assign indic[28] = \indic[28] ;
	assign indic[29] = \indic[29] ;
	assign indic[30] = \indic[30] ;
	assign indic[32] = \indic[32] ;
	assign indic[33] = \indic[33] ;
	assign indic[34] = \indic[34] ;
	assign indic[66] = \indic[35] ;
	assign indic[35] = \indic[35] ;
	assign indic[36] = \indic[36] ;
	assign indic[37] = \indic[37] ;
	assign indic[38] = \indic[38] ;
	assign indic[39] = \indic[39] ;
	assign indic[40] = \indic[40] ;
	assign indic[52] = \indic[41] ;
	assign indic[41] = \indic[41] ;
	assign indic[42] = \indic[42] ;
	assign indic[43] = \indic[43] ;
	assign indic[44] = \indic[44] ;
	assign indic[45] = \indic[45] ;
	assign indic[46] = \indic[46] ;
	assign indic[47] = \indic[47] ;
	assign indic[48] = \indic[48] ;
	assign indic[49] = \indic[49] ;
	assign indic[65] = \indic[50] ;
	assign indic[50] = \indic[50] ;
	assign indic[51] = \indic[51] ;
	assign indic[53] = \indic[53] ;
	assign indic[54] = \indic[54] ;
	assign indic[55] = \indic[55] ;
	assign indic[56] = \indic[56] ;
	assign indic[57] = \indic[57] ;
	assign indic[58] = \indic[58] ;
	assign indic[59] = \indic[59] ;
	assign indic[60] = \indic[60] ;
	assign indic[61] = \indic[61] ;
	assign indic[62] = \indic[62] ;
	assign indic[63] = \indic[63] ;
	assign indic[64] = \indic[64] ;
	assign indic[67] = \indic[67] ;
	assign indic[68] = \indic[68] ;
	assign indic[69] = \indic[69] ;
	assign indic[70] = \indic[70] ;
	assign indic[71] = \indic[71] ;
	assign indic[72] = \indic[72] ;

	notech_and3 i_79(.A(in8[6]), .B(in8[7]), .C(n_75), .Z(n_102));
	notech_and3 i_77(.A(n_29904), .B(n_29905), .C(in8[3]), .Z(n_96));
	notech_and2 i_80(.A(n_29904), .B(n_29903), .Z(n_93));
	notech_and2 i_97(.A(n_29905), .B(n_29903), .Z(n_92));
	notech_and2 i_96(.A(in8[0]), .B(in8[2]), .Z(n_90));
	notech_and4 i_72(.A(in8[6]), .B(in8[7]), .C(in8[4]), .D(n_29907), .Z(n_88
		));
	notech_and3 i_69(.A(in8[6]), .B(in8[7]), .C(n_85), .Z(n_86));
	notech_nor2 i_78(.A(in8[4]), .B(in8[5]), .Z(n_85));
	notech_and2 i_86(.A(n_29903), .B(in8[2]), .Z(n_80));
	notech_and2 i_88(.A(n_78), .B(in8[1]), .Z(n_79));
	notech_nor2 i_71(.A(in8[7]), .B(in8[6]), .Z(n_78));
	notech_nor2 i_70(.A(in8[4]), .B(n_29907), .Z(n_75));
	notech_and3 i_15(.A(in8[0]), .B(in8[3]), .C(in8[2]), .Z(n_73));
	notech_and3 i_10(.A(n_29906), .B(in8[1]), .C(n_29905), .Z(n_72));
	notech_and2 i_23(.A(in8[6]), .B(in8[7]), .Z(n_71));
	notech_and2 i_14(.A(n_29906), .B(n_29905), .Z(n_70));
	notech_and4 i_116(.A(n_92), .B(in8[1]), .C(n_29907), .D(in8[3]), .Z(n_113
		));
	notech_nand3 i_119(.A(\indic[4] ), .B(n_29906), .C(in8[0]), .Z(n_116));
	notech_and4 i_070324(.A(n_71), .B(\indic[41] ), .C(n_29906), .D(n_29905)
		, .Z(\indic[0] ));
	notech_and4 i_1(.A(n_75), .B(\indic[24] ), .C(n_29906), .D(in8[2]), .Z(\indic[1] 
		));
	notech_and4 i_2(.A(n_80), .B(in8[3]), .C(in8[5]), .D(n_79), .Z(\indic[2] 
		));
	notech_and4 i_3(.A(\indic[6] ), .B(n_80), .C(n_78), .D(in8[5]), .Z(\indic[3] 
		));
	notech_and2 i_4(.A(n_78), .B(n_29905), .Z(\indic[4] ));
	notech_and3 i_5(.A(n_75), .B(\indic[24] ), .C(n_29905), .Z(\indic[5] )
		);
	notech_and2 i_6(.A(n_29906), .B(in8[1]), .Z(\indic[6] ));
	notech_and2 i_7(.A(in8[0]), .B(in8[3]), .Z(\indic[7] ));
	notech_ao3 i_8(.A(in8[7]), .B(n_85), .C(in8[6]), .Z(\indic[8] ));
	notech_and4 i_9(.A(in8[6]), .B(in8[7]), .C(n_85), .D(n_29906), .Z(\indic[9] 
		));
	notech_and4 i_11(.A(in8[4]), .B(n_71), .C(n_70), .D(n_29907), .Z(\indic[11] 
		));
	notech_and4 i_12(.A(n_71), .B(\indic[41] ), .C(in8[2]), .D(in8[1]), .Z(\indic[12] 
		));
	notech_ao3 i_13(.A(n_78), .B(n_29907), .C(in8[4]), .Z(\indic[13] ));
	notech_and3 i_16(.A(in8[4]), .B(n_78), .C(in8[5]), .Z(\indic[16] ));
	notech_and4 i_17(.A(n_90), .B(\indic[28] ), .C(n_29906), .D(in8[1]), .Z(\indic[17] 
		));
	notech_ao3 i_18(.A(in8[7]), .B(n_75), .C(in8[6]), .Z(\indic[18] ));
	notech_and2 i_19(.A(n_29904), .B(n_29905), .Z(\indic[19] ));
	notech_and3 i_20(.A(n_29905), .B(n_29903), .C(in8[1]), .Z(\indic[60] )
		);
	notech_and4 i_21(.A(in8[6]), .B(in8[7]), .C(n_85), .D(in8[3]), .Z(\indic[20] 
		));
	notech_and3 i_22(.A(n_29904), .B(n_29903), .C(in8[2]), .Z(\indic[21] )
		);
	notech_and3 i_24(.A(n_78), .B(in8[0]), .C(in8[2]), .Z(\indic[23] ));
	notech_and2 i_25(.A(in8[6]), .B(n_29908), .Z(\indic[24] ));
	notech_nor2 i_26(.A(in8[6]), .B(n_29908), .Z(\indic[25] ));
	notech_and4 i_27(.A(n_78), .B(n_29904), .C(n_29903), .D(in8[2]), .Z(\indic[26] 
		));
	notech_and3 i_28(.A(in8[3]), .B(\indic[5] ), .C(in8[1]), .Z(\indic[27] )
		);
	notech_and3 i_29(.A(in8[4]), .B(\indic[24] ), .C(in8[5]), .Z(\indic[28] 
		));
	notech_ao3 i_30(.A(\indic[43] ), .B(n_29904), .C(in8[0]), .Z(\indic[29] 
		));
	notech_and4 i_31(.A(n_85), .B(in8[0]), .C(\indic[25] ), .D(n_72), .Z(\indic[30] 
		));
	notech_ao3 i_32(.A(\indic[18] ), .B(n_96), .C(in8[0]), .Z(\indic[32] )
		);
	notech_and4 i_33(.A(in8[4]), .B(\indic[25] ), .C(in8[5]), .D(n_29906), .Z
		(\indic[33] ));
	notech_and4 i_34(.A(n_71), .B(n_85), .C(n_70), .D(n_29904), .Z(\indic[34] 
		));
	notech_and3 i_35(.A(n_73), .B(n_86), .C(n_29904), .Z(\indic[36] ));
	notech_and4 i_36(.A(in8[2]), .B(n_29904), .C(n_88), .D(n_29906), .Z(\indic[37] 
		));
	notech_ao3 i_37(.A(n_71), .B(n_75), .C(in8[3]), .Z(\indic[38] ));
	notech_and4 i_38(.A(n_102), .B(in8[1]), .C(\indic[7] ), .D(n_29905), .Z(\indic[39] 
		));
	notech_and4 i_39(.A(\indic[6] ), .B(n_71), .C(\indic[41] ), .D(n_80), .Z
		(\indic[40] ));
	notech_and4 i_40(.A(n_86), .B(n_29905), .C(n_29903), .D(in8[1]), .Z(\indic[42] 
		));
	notech_and4 i_41(.A(\indic[25] ), .B(n_85), .C(n_29906), .D(n_29905), .Z
		(\indic[43] ));
	notech_and4 i_42(.A(n_78), .B(in8[0]), .C(in8[2]), .D(n_29904), .Z(\indic[44] 
		));
	notech_and4 i_43(.A(in8[4]), .B(\indic[25] ), .C(in8[5]), .D(in8[3]), .Z
		(\indic[45] ));
	notech_and4 i_44(.A(in8[6]), .B(in8[7]), .C(n_75), .D(n_96), .Z(\indic[46] 
		));
	notech_and3 i_45(.A(n_75), .B(\indic[24] ), .C(n_96), .Z(\indic[47] ));
	notech_and4 i_46(.A(\indic[25] ), .B(n_75), .C(n_29906), .D(n_29905), .Z
		(\indic[48] ));
	notech_and3 i_47(.A(\indic[25] ), .B(n_96), .C(in8[5]), .Z(\indic[49] )
		);
	notech_and4 i_48(.A(\indic[6] ), .B(n_71), .C(\indic[41] ), .D(n_90), .Z
		(\indic[51] ));
	notech_and2 i_49(.A(in8[4]), .B(in8[5]), .Z(\indic[41] ));
	notech_and3 i_50(.A(\indic[45] ), .B(in8[1]), .C(n_92), .Z(\indic[53] )
		);
	notech_and4 i_51(.A(n_85), .B(n_78), .C(in8[1]), .D(n_73), .Z(\indic[54] 
		));
	notech_and4 i_52(.A(n_93), .B(\indic[41] ), .C(\indic[24] ), .D(n_70), .Z
		(\indic[55] ));
	notech_ao3 i_53(.A(\indic[18] ), .B(\indic[21] ), .C(in8[3]), .Z(\indic[56] 
		));
	notech_ao3 i_54(.A(n_72), .B(n_86), .C(in8[0]), .Z(\indic[57] ));
	notech_and3 i_55(.A(in8[2]), .B(\indic[9] ), .C(n_93), .Z(\indic[58] )
		);
	notech_and4 i_56(.A(in8[0]), .B(in8[2]), .C(\indic[9] ), .D(n_29904), .Z
		(\indic[59] ));
	notech_and4 i_57(.A(in8[4]), .B(n_71), .C(in8[3]), .D(n_29907), .Z(\indic[61] 
		));
	notech_and4 i_58(.A(n_75), .B(\indic[24] ), .C(\indic[6] ), .D(n_80), .Z
		(\indic[62] ));
	notech_and4 i_59(.A(\indic[6] ), .B(n_71), .C(\indic[41] ), .D(n_29905),
		 .Z(\indic[63] ));
	notech_and4 i_60(.A(n_92), .B(in8[3]), .C(n_102), .D(in8[1]), .Z(\indic[64] 
		));
	notech_and4 i_61(.A(\indic[6] ), .B(n_86), .C(in8[0]), .D(in8[2]), .Z(\indic[50] 
		));
	notech_and4 i_62(.A(n_86), .B(n_29903), .C(in8[2]), .D(\indic[6] ), .Z(\indic[35] 
		));
	notech_and4 i_63(.A(\indic[6] ), .B(n_90), .C(n_75), .D(\indic[24] ), .Z
		(\indic[67] ));
	notech_and3 i_64(.A(in8[4]), .B(\indic[25] ), .C(n_113), .Z(\indic[68] )
		);
	notech_ao3 i_65(.A(n_85), .B(n_29904), .C(n_116), .Z(\indic[69] ));
	notech_and4 i_66(.A(\indic[18] ), .B(n_29904), .C(n_29903), .D(in8[2]), 
		.Z(\indic[70] ));
	notech_and4 i_67(.A(n_72), .B(\indic[25] ), .C(n_85), .D(n_29903), .Z(\indic[71] 
		));
	notech_and4 i_68(.A(n_72), .B(\indic[41] ), .C(\indic[25] ), .D(n_29903)
		, .Z(\indic[72] ));
	notech_inv i_33206(.A(in8[0]), .Z(n_29903));
	notech_inv i_33207(.A(in8[1]), .Z(n_29904));
	notech_inv i_33208(.A(in8[2]), .Z(n_29905));
	notech_inv i_33209(.A(in8[3]), .Z(n_29906));
	notech_inv i_33210(.A(in8[5]), .Z(n_29907));
	notech_inv i_33211(.A(in8[7]), .Z(n_29908));
	notech_inv i_33212(.A(n_70), .Z(\indic[14] ));
	notech_inv i_33213(.A(n_71), .Z(\indic[22] ));
	notech_inv i_33214(.A(n_72), .Z(\indic[10] ));
	notech_inv i_33215(.A(n_73), .Z(\indic[15] ));
endmodule
module deco_rm(in8, indic);

	input [7:0] in8;
	output [7:0] indic;




	notech_nand2 i_1(.A(in8[7]), .B(in8[6]), .Z(indic[1]));
	notech_and3 i_070325(.A(in8[2]), .B(n_29915), .C(n_29914), .Z(indic[0])
		);
	notech_and4 i_2(.A(in8[2]), .B(in8[0]), .C(indic[7]), .D(n_29914), .Z(indic
		[2]));
	notech_and2 i_3(.A(in8[7]), .B(n_29913), .Z(indic[3]));
	notech_nor2 i_4(.A(in8[7]), .B(n_29913), .Z(indic[4]));
	notech_nor2 i_5(.A(in8[5]), .B(in8[4]), .Z(indic[5]));
	notech_and4 i_6(.A(indic[7]), .B(in8[2]), .C(in8[1]), .D(n_29915), .Z(indic
		[6]));
	notech_nor2 i_7(.A(in8[7]), .B(in8[6]), .Z(indic[7]));
	notech_inv i_33225(.A(in8[6]), .Z(n_29913));
	notech_inv i_33226(.A(in8[1]), .Z(n_29914));
	notech_inv i_33227(.A(in8[0]), .Z(n_29915));
endmodule
module udecox(op, modrm, twobyte, cpl, adz, opz, jsz, udeco, fpu, emul, ipg_fault
		);

	input [7:0] op;
	input [7:0] modrm;
	input twobyte;
	input [1:0] cpl;
	input adz;
	input [2:0] opz;
	input [3:0] jsz;
	output [127:0] udeco;
	input fpu;
	input emul;
	input ipg_fault;

	wire n_4024;
	wire \udeco[0] ;
	wire \udeco[1] ;
	wire \udeco[2] ;
	wire \udeco[3] ;
	wire \udeco[4] ;
	wire \udeco[5] ;
	wire \udeco[6] ;
	wire \udeco[8] ;
	wire \udeco[9] ;
	wire \udeco[10] ;
	wire \udeco[11] ;
	wire \udeco[12] ;
	wire \udeco[13] ;
	wire \udeco[14] ;
	wire \udeco[15] ;
	wire \udeco[16] ;
	wire \udeco[17] ;
	wire \udeco[18] ;
	wire \udeco[19] ;
	wire \udeco[20] ;
	wire \udeco[21] ;
	wire \udeco[22] ;
	wire \udeco[23] ;
	wire \udeco[24] ;
	wire \udeco[25] ;
	wire \udeco[26] ;
	wire \udeco[27] ;
	wire \udeco[28] ;
	wire \udeco[29] ;
	wire \udeco[30] ;
	wire \udeco[31] ;
	wire \udeco[32] ;
	wire \udeco[33] ;
	wire \udeco[34] ;
	wire \udeco[35] ;
	wire \udeco[36] ;
	wire \udeco[37] ;
	wire \udeco[38] ;
	wire \udeco[39] ;
	wire \udeco[40] ;
	wire \udeco[41] ;
	wire \udeco[42] ;
	wire \udeco[43] ;
	wire \udeco[44] ;
	wire \udeco[45] ;
	wire \udeco[46] ;
	wire \udeco[47] ;
	wire \udeco[48] ;
	wire \udeco[49] ;
	wire \udeco[50] ;
	wire \udeco[51] ;
	wire \udeco[52] ;
	wire \udeco[53] ;
	wire \udeco[54] ;
	wire \udeco[55] ;
	wire \udeco[56] ;
	wire \udeco[57] ;
	wire \udeco[58] ;
	wire \udeco[59] ;
	wire \udeco[60] ;
	wire \udeco[61] ;
	wire \udeco[62] ;
	wire \udeco[63] ;
	wire \udeco[64] ;
	wire \udeco[65] ;
	wire \udeco[66] ;
	wire \udeco[67] ;
	wire \udeco[68] ;
	wire \udeco[69] ;
	wire \udeco[70] ;
	wire \udeco[71] ;
	wire \udeco[72] ;
	wire \udeco[73] ;
	wire \udeco[74] ;
	wire \udeco[75] ;
	wire \udeco[77] ;
	wire \udeco[78] ;
	wire \udeco[80] ;
	wire \udeco[81] ;
	wire \udeco[82] ;
	wire \udeco[83] ;
	wire \udeco[84] ;
	wire \udeco[85] ;
	wire \udeco[86] ;
	wire \udeco[87] ;
	wire \udeco[88] ;
	wire \udeco[89] ;
	wire \udeco[90] ;
	wire \udeco[91] ;
	wire \udeco[92] ;
	wire \udeco[93] ;
	wire \udeco[95] ;
	wire \udeco[96] ;
	wire \udeco[98] ;
	wire \udeco[99] ;
	wire \udeco[100] ;
	wire \udeco[101] ;
	wire \udeco[102] ;
	wire \udeco[103] ;
	wire \udeco[104] ;
	wire \udeco[105] ;
	wire \udeco[106] ;
	wire \udeco[107] ;
	wire \udeco[108] ;
	wire \udeco[109] ;
	wire \udeco[110] ;
	wire \udeco[112] ;
	wire \udeco[113] ;
	wire \udeco[114] ;
	wire \udeco[115] ;
	wire \udeco[116] ;
	wire \udeco[117] ;
	wire \udeco[118] ;
	wire \udeco[119] ;
	wire \udeco[120] ;
	wire \udeco[121] ;
	wire \udeco[122] ;
	wire \udeco[123] ;
	wire \udeco[124] ;
	wire \udeco[125] ;
	wire \udeco[126] ;
	wire \udeco[127] ;


	assign udeco[111] = n_4024;
	assign udeco[0] = \udeco[0] ;
	assign udeco[1] = \udeco[1] ;
	assign udeco[2] = \udeco[2] ;
	assign udeco[3] = \udeco[3] ;
	assign udeco[4] = \udeco[4] ;
	assign udeco[5] = \udeco[5] ;
	assign udeco[7] = \udeco[6] ;
	assign udeco[6] = \udeco[6] ;
	assign udeco[8] = \udeco[8] ;
	assign udeco[9] = \udeco[9] ;
	assign udeco[10] = \udeco[10] ;
	assign udeco[11] = \udeco[11] ;
	assign udeco[12] = \udeco[12] ;
	assign udeco[13] = \udeco[13] ;
	assign udeco[14] = \udeco[14] ;
	assign udeco[15] = \udeco[15] ;
	assign udeco[16] = \udeco[16] ;
	assign udeco[17] = \udeco[17] ;
	assign udeco[18] = \udeco[18] ;
	assign udeco[19] = \udeco[19] ;
	assign udeco[20] = \udeco[20] ;
	assign udeco[21] = \udeco[21] ;
	assign udeco[22] = \udeco[22] ;
	assign udeco[23] = \udeco[23] ;
	assign udeco[24] = \udeco[24] ;
	assign udeco[25] = \udeco[25] ;
	assign udeco[26] = \udeco[26] ;
	assign udeco[27] = \udeco[27] ;
	assign udeco[28] = \udeco[28] ;
	assign udeco[29] = \udeco[29] ;
	assign udeco[30] = \udeco[30] ;
	assign udeco[31] = \udeco[31] ;
	assign udeco[32] = \udeco[32] ;
	assign udeco[33] = \udeco[33] ;
	assign udeco[34] = \udeco[34] ;
	assign udeco[35] = \udeco[35] ;
	assign udeco[36] = \udeco[36] ;
	assign udeco[37] = \udeco[37] ;
	assign udeco[38] = \udeco[38] ;
	assign udeco[39] = \udeco[39] ;
	assign udeco[40] = \udeco[40] ;
	assign udeco[41] = \udeco[41] ;
	assign udeco[42] = \udeco[42] ;
	assign udeco[43] = \udeco[43] ;
	assign udeco[44] = \udeco[44] ;
	assign udeco[45] = \udeco[45] ;
	assign udeco[46] = \udeco[46] ;
	assign udeco[47] = \udeco[47] ;
	assign udeco[48] = \udeco[48] ;
	assign udeco[49] = \udeco[49] ;
	assign udeco[50] = \udeco[50] ;
	assign udeco[51] = \udeco[51] ;
	assign udeco[52] = \udeco[52] ;
	assign udeco[53] = \udeco[53] ;
	assign udeco[54] = \udeco[54] ;
	assign udeco[55] = \udeco[55] ;
	assign udeco[56] = \udeco[56] ;
	assign udeco[57] = \udeco[57] ;
	assign udeco[58] = \udeco[58] ;
	assign udeco[59] = \udeco[59] ;
	assign udeco[60] = \udeco[60] ;
	assign udeco[61] = \udeco[61] ;
	assign udeco[62] = \udeco[62] ;
	assign udeco[63] = \udeco[63] ;
	assign udeco[64] = \udeco[64] ;
	assign udeco[65] = \udeco[65] ;
	assign udeco[66] = \udeco[66] ;
	assign udeco[67] = \udeco[67] ;
	assign udeco[68] = \udeco[68] ;
	assign udeco[69] = \udeco[69] ;
	assign udeco[70] = \udeco[70] ;
	assign udeco[71] = \udeco[71] ;
	assign udeco[72] = \udeco[72] ;
	assign udeco[73] = \udeco[73] ;
	assign udeco[76] = \udeco[74] ;
	assign udeco[74] = \udeco[74] ;
	assign udeco[75] = \udeco[75] ;
	assign udeco[77] = \udeco[77] ;
	assign udeco[79] = \udeco[78] ;
	assign udeco[78] = \udeco[78] ;
	assign udeco[80] = \udeco[80] ;
	assign udeco[81] = \udeco[81] ;
	assign udeco[82] = \udeco[82] ;
	assign udeco[83] = \udeco[83] ;
	assign udeco[84] = \udeco[84] ;
	assign udeco[85] = \udeco[85] ;
	assign udeco[86] = \udeco[86] ;
	assign udeco[87] = \udeco[87] ;
	assign udeco[88] = \udeco[88] ;
	assign udeco[89] = \udeco[89] ;
	assign udeco[90] = \udeco[90] ;
	assign udeco[91] = \udeco[91] ;
	assign udeco[92] = \udeco[92] ;
	assign udeco[94] = \udeco[93] ;
	assign udeco[93] = \udeco[93] ;
	assign udeco[95] = \udeco[95] ;
	assign udeco[96] = \udeco[96] ;
	assign udeco[98] = \udeco[98] ;
	assign udeco[99] = \udeco[99] ;
	assign udeco[97] = \udeco[100] ;
	assign udeco[100] = \udeco[100] ;
	assign udeco[101] = \udeco[101] ;
	assign udeco[102] = \udeco[102] ;
	assign udeco[103] = \udeco[103] ;
	assign udeco[104] = \udeco[104] ;
	assign udeco[105] = \udeco[105] ;
	assign udeco[106] = \udeco[106] ;
	assign udeco[107] = \udeco[107] ;
	assign udeco[108] = \udeco[108] ;
	assign udeco[109] = \udeco[109] ;
	assign udeco[110] = \udeco[110] ;
	assign udeco[112] = \udeco[112] ;
	assign udeco[113] = \udeco[113] ;
	assign udeco[114] = \udeco[114] ;
	assign udeco[115] = \udeco[115] ;
	assign udeco[116] = \udeco[116] ;
	assign udeco[117] = \udeco[117] ;
	assign udeco[118] = \udeco[118] ;
	assign udeco[119] = \udeco[119] ;
	assign udeco[120] = \udeco[120] ;
	assign udeco[121] = \udeco[121] ;
	assign udeco[122] = \udeco[122] ;
	assign udeco[123] = \udeco[123] ;
	assign udeco[124] = \udeco[124] ;
	assign udeco[125] = \udeco[125] ;
	assign udeco[126] = \udeco[126] ;
	assign udeco[127] = \udeco[127] ;

	notech_inv i_11453(.A(n_57920), .Z(n_57925));
	notech_inv i_11449(.A(n_57920), .Z(n_57921));
	notech_inv i_11448(.A(op[0]), .Z(n_57920));
	notech_inv i_11445(.A(n_57921), .Z(n_57916));
	notech_inv i_11444(.A(n_57921), .Z(n_57915));
	notech_inv i_11439(.A(n_57921), .Z(n_57910));
	notech_inv i_11435(.A(n_57898), .Z(n_57905));
	notech_inv i_11434(.A(n_57898), .Z(n_57904));
	notech_inv i_11429(.A(n_57898), .Z(n_57899));
	notech_inv i_11428(.A(op[3]), .Z(n_57898));
	notech_inv i_11421(.A(n_57889), .Z(n_57890));
	notech_inv i_11420(.A(n_2286), .Z(n_57889));
	notech_inv i_11417(.A(n_57876), .Z(n_57885));
	notech_inv i_11413(.A(n_57876), .Z(n_57881));
	notech_inv i_11409(.A(n_57876), .Z(n_57877));
	notech_inv i_11408(.A(op[6]), .Z(n_57876));
	notech_inv i_11405(.A(n_57867), .Z(n_57872));
	notech_inv i_11401(.A(n_57867), .Z(n_57868));
	notech_inv i_11400(.A(op[4]), .Z(n_57867));
	notech_inv i_11393(.A(n_57858), .Z(n_57859));
	notech_inv i_11392(.A(n_30110), .Z(n_57858));
	notech_inv i_11389(.A(n_57849), .Z(n_57854));
	notech_inv i_11385(.A(n_57849), .Z(n_57850));
	notech_inv i_11384(.A(op[5]), .Z(n_57849));
	notech_inv i_11381(.A(n_57840), .Z(n_57845));
	notech_inv i_11377(.A(n_57840), .Z(n_57841));
	notech_inv i_11376(.A(op[2]), .Z(n_57840));
	notech_inv i_11363(.A(n_57824), .Z(n_57825));
	notech_inv i_11362(.A(n_30108), .Z(n_57824));
	notech_inv i_11359(.A(n_57815), .Z(n_57820));
	notech_inv i_11355(.A(n_57815), .Z(n_57816));
	notech_inv i_11354(.A(op[1]), .Z(n_57815));
	notech_inv i_11351(.A(n_57799), .Z(n_57811));
	notech_inv i_11350(.A(n_57799), .Z(n_57810));
	notech_inv i_11345(.A(n_57799), .Z(n_57805));
	notech_inv i_11340(.A(n_57799), .Z(n_57800));
	notech_inv i_11339(.A(n_2328), .Z(n_57799));
	notech_inv i_11335(.A(n_57904), .Z(n_57794));
	notech_inv i_11330(.A(n_57904), .Z(n_57789));
	notech_inv i_11322(.A(n_57779), .Z(n_57780));
	notech_inv i_11321(.A(n_30111), .Z(n_57779));
	notech_inv i_11314(.A(n_57770), .Z(n_57771));
	notech_inv i_11313(.A(n_2325), .Z(n_57770));
	notech_inv i_11306(.A(n_57761), .Z(n_57762));
	notech_inv i_11305(.A(n_2271), .Z(n_57761));
	notech_inv i_11298(.A(n_57752), .Z(n_57753));
	notech_inv i_11297(.A(n_30107), .Z(n_57752));
	notech_inv i_11290(.A(n_57743), .Z(n_57744));
	notech_inv i_11289(.A(n_29925), .Z(n_57743));
	notech_inv i_11282(.A(n_57734), .Z(n_57735));
	notech_inv i_11281(.A(n_2282), .Z(n_57734));
	notech_inv i_11274(.A(n_57725), .Z(n_57726));
	notech_inv i_11273(.A(modrm[5]), .Z(n_57725));
	notech_inv i_11266(.A(n_57716), .Z(n_57717));
	notech_inv i_11265(.A(n_30117), .Z(n_57716));
	notech_inv i_11254(.A(n_57702), .Z(n_57703));
	notech_inv i_11253(.A(n_2360), .Z(n_57702));
	notech_inv i_11246(.A(n_57693), .Z(n_57694));
	notech_inv i_11245(.A(n_2410), .Z(n_57693));
	notech_and4 i_1531(.A(n_2839), .B(n_1543), .C(n_2931), .D(n_2924), .Z(n_2934
		));
	notech_ao3 i_1534(.A(n_2934), .B(n_2904), .C(n_30025), .Z(n_2936));
	notech_and2 i_793(.A(n_2179), .B(n_1603), .Z(n_2937));
	notech_and4 i_1535(.A(n_2663), .B(n_2352), .C(n_2937), .D(n_2567), .Z(n_2939
		));
	notech_and4 i_1546(.A(n_3993), .B(n_4040), .C(n_3733), .D(n_1907), .Z(n_2942
		));
	notech_and4 i_306(.A(n_2137), .B(n_2942), .C(n_2026), .D(n_3984), .Z(n_2945
		));
	notech_and3 i_770(.A(n_2638), .B(n_2014), .C(n_1896), .Z(n_2946));
	notech_and4 i_1552(.A(n_4019), .B(n_2080), .C(n_2945), .D(n_2946), .Z(n_2949
		));
	notech_and4 i_1557(.A(n_2189), .B(n_2206), .C(n_2028), .D(n_2457), .Z(n_2953
		));
	notech_and4 i_245(.A(n_2611), .B(n_2949), .C(n_2953), .D(n_2484), .Z(n_2955
		));
	notech_and4 i_1561(.A(n_2435), .B(n_2631), .C(n_1953), .D(n_2030), .Z(n_2958
		));
	notech_and4 i_303(.A(n_2141), .B(n_4013), .C(n_2058), .D(n_2958), .Z(n_2959
		));
	notech_and3 i_1569(.A(n_2033), .B(n_2032), .C(n_4020), .Z(n_2961));
	notech_and4 i_1572(.A(n_2176), .B(n_1837), .C(n_2034), .D(n_2961), .Z(n_2964
		));
	notech_and4 i_724(.A(n_2332), .B(n_2964), .C(n_2091), .D(n_3972), .Z(n_2967
		));
	notech_and4 i_521(.A(n_29992), .B(n_29957), .C(n_29991), .D(n_2031), .Z(n_2969
		));
	notech_ao4 i_1576(.A(n_3963), .B(n_2574), .C(n_2362), .D(n_2331), .Z(n_2970
		));
	notech_and4 i_1578(.A(n_3992), .B(n_1895), .C(n_2970), .D(n_3672), .Z(n_2972
		));
	notech_and4 i_1581(.A(n_2972), .B(n_2406), .C(n_2969), .D(n_2967), .Z(n_2975
		));
	notech_ao3 i_653(.A(n_2668), .B(n_3777), .C(n_29929), .Z(n_2978));
	notech_and4 i_1607(.A(n_843), .B(n_1332), .C(n_2494), .D(n_2046), .Z(n_2983
		));
	notech_and3 i_1611(.A(n_3994), .B(n_2983), .C(n_1340), .Z(n_2985));
	notech_and4 i_1615(.A(n_1329), .B(n_2021), .C(n_2562), .D(n_2985), .Z(n_2987
		));
	notech_ao4 i_510(.A(n_2098), .B(n_2101), .C(n_4065), .D(n_2027), .Z(n_2988
		));
	notech_ao4 i_1598(.A(n_29995), .B(n_30042), .C(adz), .D(n_2305), .Z(n_2989
		));
	notech_and4 i_1596(.A(n_2040), .B(n_2219), .C(n_29979), .D(n_2041), .Z(n_2992
		));
	notech_and4 i_1600(.A(n_2042), .B(n_2045), .C(n_2989), .D(n_2992), .Z(n_2995
		));
	notech_and4 i_1603(.A(n_2195), .B(n_4022), .C(n_2995), .D(n_1346), .Z(n_2999
		));
	notech_and4 i_1610(.A(n_2050), .B(n_2999), .C(n_2051), .D(n_2053), .Z(n_3002
		));
	notech_and4 i_1616(.A(n_3002), .B(n_1728), .C(n_2665), .D(n_2246), .Z(n_3005
		));
	notech_ao4 i_1633(.A(n_29995), .B(n_2574), .C(n_30053), .D(n_2355), .Z(n_3008
		));
	notech_ao3 i_1635(.A(n_2829), .B(n_3008), .C(n_3820), .Z(n_3010));
	notech_and4 i_244(.A(n_2392), .B(n_2967), .C(n_3955), .D(n_3010), .Z(n_3013
		));
	notech_and4 i_1640(.A(n_2435), .B(n_2631), .C(n_1526), .D(n_4025), .Z(n_3015
		));
	notech_and4 i_1643(.A(n_3015), .B(n_2379), .C(n_2852), .D(n_1905), .Z(n_3018
		));
	notech_and2 i_726(.A(n_3890), .B(n_2238), .Z(n_3021));
	notech_and4 i_1656(.A(n_1855), .B(n_1854), .C(n_4028), .D(n_2071), .Z(n_3023
		));
	notech_and4 i_1662(.A(n_2073), .B(n_3023), .C(n_1656), .D(n_2076), .Z(n_3026
		));
	notech_ao3 i_1669(.A(n_3026), .B(n_3021), .C(n_2077), .Z(n_3028));
	notech_and3 i_176(.A(n_4026), .B(n_1284), .C(n_4027), .Z(n_3030));
	notech_and4 i_1672(.A(n_3977), .B(n_1306), .C(n_3030), .D(n_3028), .Z(n_3033
		));
	notech_and4 i_1653(.A(n_2252), .B(n_222291111), .C(n_2188), .D(n_2070), 
		.Z(n_3039));
	notech_and4 i_1659(.A(n_2190), .B(n_3039), .C(n_2709), .D(n_2072), .Z(n_3042
		));
	notech_and4 i_1668(.A(n_3042), .B(n_4029), .C(n_2074), .D(n_1290), .Z(n_3045
		));
	notech_and4 i_1671(.A(n_3045), .B(n_2075), .C(n_2598), .D(n_4005), .Z(n_3046
		));
	notech_and4 i_1675(.A(n_4055), .B(n_1857), .C(n_3046), .D(n_3033), .Z(n_3048
		));
	notech_and2 i_549(.A(n_2264), .B(n_1911), .Z(n_3049));
	notech_and4 i_1677(.A(n_3049), .B(n_3048), .C(n_2789), .D(n_29930), .Z(n_3052
		));
	notech_and4 i_1679(.A(n_1329), .B(n_2021), .C(n_2826), .D(n_3052), .Z(n_3054
		));
	notech_and3 i_210(.A(n_4027), .B(n_4036), .C(n_4076), .Z(n_3056));
	notech_and4 i_1720(.A(n_2151), .B(n_3992), .C(n_3977), .D(n_29965), .Z(n_3059
		));
	notech_and2 i_624(.A(n_4017), .B(n_4019), .Z(n_3061));
	notech_and3 i_556(.A(n_2192), .B(n_4017), .C(n_3981), .Z(n_3062));
	notech_and4 i_1527(.A(n_1434), .B(n_2928), .C(n_29959), .D(n_4016), .Z(n_2931
		));
	notech_and3 i_206(.A(n_29978), .B(n_1958), .C(n_2377), .Z(n_3064));
	notech_ao4 i_1780(.A(n_30058), .B(n_57916), .C(n_30100), .D(n_30115), .Z
		(n_3067));
	notech_and3 i_1782(.A(n_3067), .B(n_2086), .C(n_3980), .Z(n_3069));
	notech_and4 i_1787(.A(n_4047), .B(n_223489126), .C(n_3069), .D(n_2305), 
		.Z(n_3072));
	notech_ao4 i_1788(.A(n_2124), .B(n_57794), .C(n_2333), .D(n_2359), .Z(n_3073
		));
	notech_and4 i_1792(.A(n_4017), .B(n_3073), .C(n_3072), .D(n_4019), .Z(n_3075
		));
	notech_and4 i_1799(.A(n_3075), .B(n_3967), .C(n_2090), .D(n_3064), .Z(n_3078
		));
	notech_and2 i_4702(.A(n_29961), .B(n_4082), .Z(n_3079));
	notech_and4 i_1789(.A(n_3079), .B(n_2087), .C(n_2089), .D(n_1624), .Z(n_3083
		));
	notech_and4 i_1795(.A(n_3083), .B(n_2579), .C(n_2609), .D(n_3981), .Z(n_3086
		));
	notech_and4 i_1800(.A(n_2663), .B(n_3086), .C(n_2978), .D(n_2091), .Z(n_3089
		));
	notech_and4 i_1803(.A(n_3089), .B(n_3078), .C(n_5254), .D(n_29986), .Z(n_3091
		));
	notech_and2 i_1808(.A(n_4040), .B(n_733), .Z(n_3095));
	notech_and4 i_258(.A(n_4002), .B(n_1332), .C(n_1329), .D(n_3095), .Z(n_3098
		));
	notech_ao3 i_809(.A(n_4055), .B(n_2097), .C(n_2100), .Z(n_3102));
	notech_ao4 i_560(.A(n_2499), .B(n_2485), .C(n_2596), .D(n_2302), .Z(n_3103
		));
	notech_and4 i_1821(.A(n_1984), .B(n_1801), .C(n_2159), .D(n_2104), .Z(n_3105
		));
	notech_and3 i_20372292(.A(n_2206), .B(n_4028), .C(n_2790), .Z(n_3107));
	notech_and3 i_296(.A(n_3965), .B(n_2579), .C(n_29989), .Z(n_2928));
	notech_and3 i_64772262(.A(n_2238), .B(n_4053), .C(n_2159), .Z(n_3109));
	notech_and4 i_1864(.A(n_3109), .B(n_222191110), .C(n_3107), .D(n_29994),
		 .Z(n_3111));
	notech_and4 i_1869(.A(n_3111), .B(n_2327), .C(n_2103), .D(n_29961), .Z(n_3114
		));
	notech_and4 i_1874(.A(n_29978), .B(n_4044), .C(n_3114), .D(n_4027), .Z(n_3117
		));
	notech_and4 i_1877(.A(n_2057), .B(n_1794), .C(n_2105), .D(n_3117), .Z(n_3119
		));
	notech_and4 i_1884(.A(n_3119), .B(n_2480), .C(n_2108), .D(n_2572), .Z(n_3122
		));
	notech_and2 i_719(.A(n_2218), .B(n_3970), .Z(n_3124));
	notech_and4 i_1887(.A(n_3970), .B(n_3122), .C(n_2218), .D(n_2116), .Z(n_3126
		));
	notech_ao3 i_317(.A(n_2609), .B(n_1792), .C(n_1795), .Z(n_3128));
	notech_and4 i_1871(.A(n_1932), .B(n_2123), .C(n_4041), .D(n_4043), .Z(n_3131
		));
	notech_and4 i_1879(.A(n_3131), .B(n_2107), .C(n_2104), .D(n_2106), .Z(n_3134
		));
	notech_and4 i_1883(.A(n_2176), .B(n_2195), .C(n_1970), .D(n_3134), .Z(n_3136
		));
	notech_and4 i_1888(.A(n_30063), .B(n_3128), .C(n_3136), .D(n_29959), .Z(n_3138
		));
	notech_and4 i_1891(.A(n_3098), .B(n_3126), .C(n_2109), .D(n_3138), .Z(n_3141
		));
	notech_and2 i_4754(.A(n_2688), .B(n_3739), .Z(n_3143));
	notech_and4 i_1924(.A(n_2579), .B(n_1970), .C(n_222891117), .D(n_2125), 
		.Z(n_3145));
	notech_and4 i_1917(.A(n_3061), .B(n_4032), .C(n_3981), .D(n_2122), .Z(n_3150
		));
	notech_and4 i_1919(.A(n_574), .B(n_4046), .C(n_2121), .D(n_3150), .Z(n_3151
		));
	notech_ao4 i_746(.A(n_2297), .B(n_2118), .C(n_2382), .D(n_2325), .Z(n_3152
		));
	notech_and4 i_444(.A(n_1855), .B(n_1854), .C(n_2111), .D(n_2255), .Z(n_3154
		));
	notech_and3 i_1904(.A(n_2119), .B(n_223489126), .C(n_30100), .Z(n_3157)
		);
	notech_and4 i_1908(.A(n_2627), .B(n_29961), .C(n_2364), .D(n_3157), .Z(n_3160
		));
	notech_and4 i_1910(.A(n_3154), .B(n_3160), .C(n_3992), .D(n_2120), .Z(n_3162
		));
	notech_and4 i_1918(.A(n_3152), .B(n_709), .C(n_3162), .D(n_2465), .Z(n_3165
		));
	notech_and4 i_1923(.A(n_673), .B(n_3165), .C(n_3151), .D(n_960), .Z(n_3168
		));
	notech_and4 i_1927(.A(n_3168), .B(n_703), .C(n_2126), .D(n_3145), .Z(n_3171
		));
	notech_nand2 i_441(.A(n_2625), .B(n_3779), .Z(n_3174));
	notech_and4 i_817(.A(n_2631), .B(n_1780), .C(n_2137), .D(n_29931), .Z(n_3177
		));
	notech_and3 i_811(.A(n_4058), .B(n_2049), .C(n_2129), .Z(n_3178));
	notech_and2 i_234(.A(n_3178), .B(n_2130), .Z(n_3179));
	notech_and3 i_1937(.A(n_2141), .B(n_2131), .C(n_29972), .Z(n_3181));
	notech_and4 i_1940(.A(n_2258), .B(n_3975), .C(n_3181), .D(n_29946), .Z(n_3184
		));
	notech_and3 i_1988(.A(n_3982), .B(n_29958), .C(n_455), .Z(n_3187));
	notech_and4 i_1981(.A(n_3977), .B(n_2377), .C(n_2134), .D(n_2978), .Z(n_3193
		));
	notech_and4 i_1986(.A(n_2218), .B(n_3970), .C(n_3193), .D(n_444), .Z(n_3195
		));
	notech_and3 i_37472278(.A(n_2104), .B(n_3154), .C(n_4046), .Z(n_3197));
	notech_ao4 i_1972(.A(n_2400), .B(n_2497), .C(n_2278), .D(n_2339), .Z(n_3200
		));
	notech_and4 i_1974(.A(n_3197), .B(n_2216), .C(n_4051), .D(n_3200), .Z(n_3201
		));
	notech_and4 i_1976(.A(n_29978), .B(n_4019), .C(n_3201), .D(n_1923), .Z(n_3204
		));
	notech_and4 i_1983(.A(n_3204), .B(n_2579), .C(n_2395), .D(n_3021), .Z(n_3207
		));
	notech_and4 i_1985(.A(n_4002), .B(n_1526), .C(n_3207), .D(n_2166), .Z(n_3208
		));
	notech_and4 i_1991(.A(n_2522), .B(n_3208), .C(n_3195), .D(n_2352), .Z(n_3211
		));
	notech_and4 i_1993(.A(n_3177), .B(n_3187), .C(n_3211), .D(n_2893), .Z(n_3213
		));
	notech_and4 i_2032(.A(n_2555), .B(n_1873), .C(n_3102), .D(n_3178), .Z(n_3217
		));
	notech_and4 i_2039(.A(n_3217), .B(n_2352), .C(n_2308), .D(n_2294), .Z(n_3219
		));
	notech_and4 i_2030(.A(n_3021), .B(n_2513), .C(n_3972), .D(n_2144), .Z(n_3223
		));
	notech_ao3 i_2013(.A(n_4028), .B(n_1829), .C(n_2142), .Z(n_3225));
	notech_and4 i_2007(.A(n_2433), .B(n_4048), .C(n_1263), .D(n_696), .Z(n_3227
		));
	notech_and4 i_2010(.A(n_2140), .B(n_4014), .C(n_2141), .D(n_3227), .Z(n_3230
		));
	notech_and4 i_2015(.A(n_3230), .B(n_4051), .C(n_3225), .D(n_29972), .Z(n_3233
		));
	notech_and4 i_2019(.A(n_1656), .B(n_4007), .C(n_3233), .D(n_29955), .Z(n_3236
		));
	notech_and3 i_2020(.A(n_1958), .B(n_4022), .C(n_29946), .Z(n_3240));
	notech_and4 i_2026(.A(n_3103), .B(n_3240), .C(n_2143), .D(n_29962), .Z(n_3243
		));
	notech_and4 i_2028(.A(n_3236), .B(n_3243), .C(n_3697), .D(n_2614), .Z(n_3244
		));
	notech_and4 i_2037(.A(n_3244), .B(n_466), .C(n_2854), .D(n_3223), .Z(n_3247
		));
	notech_and4 i_259(.A(n_3970), .B(n_2136), .C(n_2137), .D(n_1332), .Z(n_3250
		));
	notech_ao4 i_571(.A(n_2139), .B(n_30057), .C(n_2458), .D(n_2275), .Z(n_3252
		));
	notech_and4 i_2038(.A(n_3252), .B(n_3250), .C(n_2145), .D(n_455), .Z(n_3254
		));
	notech_and4 i_2042(.A(n_3254), .B(n_3247), .C(n_3219), .D(n_2834), .Z(n_3257
		));
	notech_ao4 i_171(.A(n_2278), .B(n_2154), .C(n_2318), .D(n_2161), .Z(n_3261
		));
	notech_and3 i_2073(.A(n_3970), .B(n_2166), .C(n_2168), .Z(n_3263));
	notech_and4 i_2082(.A(n_2065), .B(n_3261), .C(n_3263), .D(n_1623), .Z(n_3266
		));
	notech_and4 i_2091(.A(n_2538), .B(n_2663), .C(n_2173), .D(n_3266), .Z(n_3269
		));
	notech_and4 i_2097(.A(n_3979), .B(n_3269), .C(n_4032), .D(n_3984), .Z(n_3271
		));
	notech_and4 i_2105(.A(n_3271), .B(n_2526), .C(n_3179), .D(n_2175), .Z(n_3273
		));
	notech_and4 i_764(.A(n_2234), .B(n_4005), .C(n_2159), .D(n_4004), .Z(n_3275
		));
	notech_ao4 i_627(.A(n_30051), .B(n_2517), .C(n_3963), .D(n_2407), .Z(n_3276
		));
	notech_or4 i_98(.A(n_2403), .B(n_2311), .C(n_57845), .D(n_30107), .Z(n_3277
		));
	notech_and2 i_360472311(.A(n_1797), .B(n_2106), .Z(n_3279));
	notech_ao4 i_1502(.A(n_2140), .B(n_57925), .C(n_2433), .D(n_57905), .Z(n_2925
		));
	notech_and3 i_38272277(.A(n_1993), .B(n_2665), .C(n_3143), .Z(n_3280));
	notech_ao3 i_2067(.A(n_3280), .B(n_3279), .C(n_30091), .Z(n_3282));
	notech_and3 i_2068(.A(n_1925), .B(n_3107), .C(n_3282), .Z(n_3283));
	notech_and4 i_2072(.A(n_2516), .B(n_3283), .C(n_2163), .D(n_1828), .Z(n_3286
		));
	notech_and4 i_2079(.A(n_3286), .B(n_2170), .C(n_3276), .D(n_2169), .Z(n_3289
		));
	notech_ao4 i_777(.A(n_2495), .B(n_2376), .C(n_2337), .D(n_29968), .Z(n_3290
		));
	notech_and4 i_2083(.A(n_3290), .B(n_2076), .C(n_3289), .D(n_3890), .Z(n_3293
		));
	notech_and4 i_2087(.A(n_3975), .B(n_4037), .C(n_2172), .D(n_2174), .Z(n_3297
		));
	notech_and4 i_2092(.A(n_3293), .B(n_1526), .C(n_2639), .D(n_3297), .Z(n_3299
		));
	notech_and4 i_2103(.A(n_673), .B(n_3299), .C(n_3275), .D(n_3177), .Z(n_3302
		));
	notech_and4 i_2096(.A(n_3987), .B(n_2029), .C(n_3128), .D(n_1712), .Z(n_3307
		));
	notech_and4 i_2104(.A(n_3252), .B(n_3307), .C(n_2563), .D(n_497), .Z(n_3309
		));
	notech_ao4 i_2112(.A(n_2329), .B(n_2448), .C(n_2407), .D(n_2408), .Z(n_3312
		));
	notech_and2 i_2127(.A(n_2188), .B(n_4013), .Z(n_3316));
	notech_and4 i_2130(.A(n_2189), .B(n_2234), .C(n_2190), .D(n_3316), .Z(n_3319
		));
	notech_and4 i_2139(.A(n_2192), .B(n_3319), .C(n_4051), .D(n_3290), .Z(n_3322
		));
	notech_ao4 i_2131(.A(n_2278), .B(n_30066), .C(n_30043), .D(n_2531), .Z(n_3323
		));
	notech_and4 i_2140(.A(n_3323), .B(n_2631), .C(n_3276), .D(n_29952), .Z(n_3326
		));
	notech_and4 i_2150(.A(n_3326), .B(n_3322), .C(n_2196), .D(n_29989), .Z(n_3329
		));
	notech_and4 i_2138(.A(n_2193), .B(n_223489126), .C(n_2327), .D(n_29954),
		 .Z(n_3333));
	notech_and4 i_2147(.A(n_3333), .B(n_1892), .C(n_3672), .D(n_1806), .Z(n_3336
		));
	notech_and4 i_2154(.A(n_3329), .B(n_2380), .C(n_2377), .D(n_3336), .Z(n_3338
		));
	notech_and4 i_2162(.A(n_2198), .B(n_3056), .C(n_1970), .D(n_3338), .Z(n_3340
		));
	notech_and4 i_2172(.A(n_3340), .B(n_3728), .C(n_493), .D(n_2200), .Z(n_3343
		));
	notech_ao4 i_2144(.A(n_2186), .B(n_57794), .C(n_1819), .D(n_2285), .Z(n_3347
		));
	notech_and4 i_2152(.A(n_3347), .B(n_2195), .C(n_2639), .D(n_2565), .Z(n_3349
		));
	notech_and4 i_2160(.A(n_2723), .B(n_3349), .C(n_2533), .D(n_2197), .Z(n_3351
		));
	notech_and4 i_2167(.A(n_2663), .B(n_3351), .C(n_2945), .D(n_2183), .Z(n_3353
		));
	notech_and3 i_453(.A(n_4032), .B(n_2365), .C(n_2181), .Z(n_3355));
	notech_and4 i_2161(.A(n_4034), .B(n_2465), .C(n_4053), .D(n_1924), .Z(n_3358
		));
	notech_and4 i_1529(.A(n_2921), .B(n_2534), .C(n_2620), .D(n_2656), .Z(n_2924
		));
	notech_and3 i_3668(.A(n_4031), .B(n_4056), .C(n_29986), .Z(n_3360));
	notech_and4 i_2168(.A(n_497), .B(n_3358), .C(n_3360), .D(n_2199), .Z(n_3362
		));
	notech_and4 i_2173(.A(n_3362), .B(n_533), .C(n_3353), .D(n_3355), .Z(n_3364
		));
	notech_and3 i_2177(.A(n_2258), .B(n_3739), .C(n_2202), .Z(n_3367));
	notech_and4 i_375(.A(n_3049), .B(n_2790), .C(n_3367), .D(n_1905), .Z(n_3370
		));
	notech_and4 i_2203(.A(n_4005), .B(n_2532), .C(n_2218), .D(n_3779), .Z(n_3373
		));
	notech_ao4 i_488(.A(n_2412), .B(n_30067), .C(n_2455), .D(n_2297), .Z(n_3374
		));
	notech_and4 i_2195(.A(n_2637), .B(n_3374), .C(n_3965), .D(n_2207), .Z(n_3377
		));
	notech_and4 i_2186(.A(n_4048), .B(n_3109), .C(n_2516), .D(n_2206), .Z(n_3381
		));
	notech_and4 i_2189(.A(n_1855), .B(n_3381), .C(n_1854), .D(n_29954), .Z(n_3383
		));
	notech_and4 i_2192(.A(n_2668), .B(n_3383), .C(n_3973), .D(n_29951), .Z(n_3385
		));
	notech_and4 i_2199(.A(n_3385), .B(n_3377), .C(n_2305), .D(n_4056), .Z(n_3388
		));
	notech_ao4 i_815(.A(n_2205), .B(n_2285), .C(n_2331), .D(n_2586), .Z(n_3389
		));
	notech_and4 i_2202(.A(n_3777), .B(n_4055), .C(n_3389), .D(n_3388), .Z(n_3392
		));
	notech_and4 i_2205(.A(n_1796), .B(n_3392), .C(n_3373), .D(n_4029), .Z(n_3394
		));
	notech_and4 i_2208(.A(n_3250), .B(n_3394), .C(n_960), .D(n_3370), .Z(n_3397
		));
	notech_and2 i_408972310(.A(n_4079), .B(n_1984), .Z(n_3402));
	notech_and4 i_59972269(.A(n_2192), .B(n_2305), .C(n_29972), .D(n_29951),
		 .Z(n_3403));
	notech_and4 i_2219(.A(n_3403), .B(n_3402), .C(n_4048), .D(n_2668), .Z(n_3406
		));
	notech_and4 i_2222(.A(n_4058), .B(n_3406), .C(n_3838), .D(n_2216), .Z(n_3408
		));
	notech_and4 i_2225(.A(n_3408), .B(n_4029), .C(n_2217), .D(n_730), .Z(n_3411
		));
	notech_and4 i_2228(.A(n_2218), .B(n_3411), .C(n_3030), .D(n_3981), .Z(n_3413
		));
	notech_and4 i_2232(.A(n_3413), .B(n_2538), .C(n_2111), .D(n_29959), .Z(n_3415
		));
	notech_and4 i_2233(.A(n_2395), .B(n_218), .C(n_4049), .D(n_2411), .Z(n_3419
		));
	notech_and4 i_2236(.A(n_2534), .B(n_3415), .C(n_3250), .D(n_3419), .Z(n_3421
		));
	notech_ao4 i_2214(.A(n_30051), .B(n_2594), .C(n_2391), .D(n_29968), .Z(n_3422
		));
	notech_and4 i_2239(.A(n_204), .B(n_3421), .C(n_3370), .D(n_2379), .Z(n_3425
		));
	notech_and4 i_2281(.A(n_3994), .B(n_204), .C(n_3370), .D(n_4085), .Z(n_3429
		));
	notech_ao4 i_2258(.A(n_2678), .B(n_30111), .C(n_2485), .D(n_2689), .Z(n_3430
		));
	notech_and4 i_2261(.A(n_2631), .B(n_3374), .C(n_3430), .D(n_2222), .Z(n_3433
		));
	notech_and4 i_2253(.A(n_3998), .B(n_2220), .C(n_3402), .D(n_29990), .Z(n_3437
		));
	notech_and4 i_2257(.A(n_2221), .B(n_2130), .C(n_2223), .D(n_3437), .Z(n_3440
		));
	notech_and4 i_2264(.A(n_3975), .B(n_3103), .C(n_3389), .D(n_3440), .Z(n_3443
		));
	notech_and4 i_2268(.A(n_3433), .B(n_3443), .C(n_2116), .D(n_29965), .Z(n_3445
		));
	notech_and4 i_2269(.A(n_3030), .B(n_1130), .C(n_2695), .D(n_2854), .Z(n_3449
		));
	notech_and4 i_2274(.A(n_2675), .B(n_3449), .C(n_3445), .D(n_29960), .Z(n_3451
		));
	notech_and4 i_2272(.A(n_2076), .B(n_2080), .C(n_3275), .D(n_29946), .Z(n_3452
		));
	notech_and4 i_2278(.A(n_444), .B(n_960), .C(n_2722), .D(n_2226), .Z(n_3457
		));
	notech_and4 i_2280(.A(n_2534), .B(n_3452), .C(n_3451), .D(n_3457), .Z(n_3458
		));
	notech_and4 i_2326(.A(n_2294), .B(n_2587), .C(n_1340), .D(n_2228), .Z(n_3463
		));
	notech_and4 i_2330(.A(n_3994), .B(n_3463), .C(n_29960), .D(n_2850), .Z(n_3465
		));
	notech_ao4 i_2300(.A(n_2363), .B(n_2412), .C(n_2065), .D(n_30107), .Z(n_3466
		));
	notech_and4 i_2308(.A(n_3466), .B(n_3154), .C(n_2598), .D(n_4037), .Z(n_3469
		));
	notech_and4 i_2318(.A(n_3469), .B(n_2614), .C(n_1332), .D(n_29944), .Z(n_3472
		));
	notech_and4 i_2312(.A(n_2238), .B(n_4031), .C(n_2239), .D(n_2099), .Z(n_3475
		));
	notech_and4 i_2321(.A(n_4034), .B(n_3475), .C(n_3062), .D(n_3472), .Z(n_3478
		));
	notech_and2 i_631(.A(n_2229), .B(n_3965), .Z(n_3481));
	notech_and4 i_2297(.A(n_2231), .B(n_3279), .C(n_2232), .D(n_2233), .Z(n_3485
		));
	notech_and4 i_2301(.A(n_4028), .B(n_3485), .C(n_223489126), .D(n_4044), 
		.Z(n_3488));
	notech_and4 i_2307(.A(n_3488), .B(n_2394), .C(n_2237), .D(n_4084), .Z(n_3490
		));
	notech_and4 i_2310(.A(n_4007), .B(n_29951), .C(n_1936), .D(n_3490), .Z(n_3491
		));
	notech_and4 i_2317(.A(n_2572), .B(n_29958), .C(n_3481), .D(n_3491), .Z(n_3494
		));
	notech_and4 i_2322(.A(n_4076), .B(n_3494), .C(n_2615), .D(n_3128), .Z(n_3496
		));
	notech_and4 i_2327(.A(n_3496), .B(n_3252), .C(n_2240), .D(n_3478), .Z(n_3498
		));
	notech_and4 i_2331(.A(n_1329), .B(n_2021), .C(n_3498), .D(n_2898), .Z(n_3500
		));
	notech_and2 i_2381(.A(n_2723), .B(n_2946), .Z(n_3507));
	notech_ao4 i_2368(.A(n_57916), .B(n_2250), .C(n_2285), .D(n_2245), .Z(n_3508
		));
	notech_and2 i_21972291(.A(n_4007), .B(n_4047), .Z(n_3510));
	notech_and4 i_2356(.A(n_1193), .B(n_1833), .C(n_3510), .D(n_29947), .Z(n_3513
		));
	notech_and4 i_2359(.A(n_2252), .B(n_3513), .C(n_2253), .D(n_2254), .Z(n_3516
		));
	notech_ao3 i_2361(.A(n_3516), .B(n_2255), .C(n_1807), .Z(n_3518));
	notech_and4 i_2364(.A(n_4058), .B(n_2256), .C(n_2257), .D(n_3518), .Z(n_3521
		));
	notech_and4 i_2367(.A(n_2233), .B(n_1938), .C(n_3521), .D(n_2571), .Z(n_3523
		));
	notech_and4 i_2374(.A(n_2263), .B(n_3523), .C(n_3508), .D(n_2262), .Z(n_3525
		));
	notech_and4 i_2375(.A(n_4017), .B(n_4019), .C(n_4022), .D(n_2264), .Z(n_3528
		));
	notech_and4 i_2379(.A(n_2206), .B(n_733), .C(n_2265), .D(n_3528), .Z(n_3530
		));
	notech_and4 i_2384(.A(n_3525), .B(n_3530), .C(n_3507), .D(n_2266), .Z(n_3532
		));
	notech_ao4 i_2366(.A(n_30051), .B(n_30042), .C(n_2285), .D(n_2288), .Z(n_3534
		));
	notech_and4 i_2377(.A(n_3534), .B(n_3261), .C(n_2532), .D(n_3481), .Z(n_3537
		));
	notech_and4 i_2385(.A(n_4046), .B(n_3537), .C(n_3967), .D(n_29986), .Z(n_3540
		));
	notech_and4 i_2390(.A(n_3540), .B(n_3532), .C(n_466), .D(n_2790), .Z(n_3542
		));
	notech_and4 i_2391(.A(n_2304), .B(n_960), .C(n_3542), .D(n_2267), .Z(n_3543
		));
	notech_and3 i_3610(.A(n_223489126), .B(n_1792), .C(n_3355), .Z(n_3545)
		);
	notech_and4 i_2394(.A(n_68), .B(n_901), .C(n_3543), .D(n_3545), .Z(n_3548
		));
	notech_ao3 i_2425(.A(n_894), .B(n_2620), .C(n_30020), .Z(n_3552));
	notech_and4 i_2431(.A(n_2826), .B(n_3452), .C(n_2157), .D(n_3552), .Z(n_3553
		));
	notech_and4 i_2432(.A(n_2884), .B(n_1728), .C(n_2379), .D(n_2850), .Z(n_3556
		));
	notech_and3 i_2433(.A(n_4016), .B(n_2498), .C(n_3972), .Z(n_3558));
	notech_and4 i_2440(.A(n_3556), .B(n_3553), .C(n_3558), .D(n_2937), .Z(n_3560
		));
	notech_and4 i_2416(.A(n_3062), .B(n_2560), .C(n_2610), .D(n_2829), .Z(n_3564
		));
	notech_and4 i_2400(.A(n_3107), .B(n_2614), .C(n_2269), .D(n_29990), .Z(n_3567
		));
	notech_and4 i_2404(.A(n_2516), .B(n_2638), .C(n_3567), .D(n_1985), .Z(n_3570
		));
	notech_and4 i_2407(.A(n_3570), .B(n_2709), .C(n_2631), .D(n_3834), .Z(n_3572
		));
	notech_and4 i_2411(.A(n_4058), .B(n_2049), .C(n_2457), .D(n_3572), .Z(n_3574
		));
	notech_and4 i_2408(.A(n_2678), .B(n_2791), .C(n_730), .D(n_1958), .Z(n_3576
		));
	notech_and4 i_2415(.A(n_3576), .B(n_3779), .C(n_3574), .D(n_2099), .Z(n_3579
		));
	notech_and4 i_2420(.A(n_2555), .B(n_3579), .C(n_3564), .D(n_2557), .Z(n_3581
		));
	notech_and4 i_2423(.A(n_2686), .B(n_2675), .C(n_2526), .D(n_3581), .Z(n_3584
		));
	notech_and4 i_2434(.A(n_2903), .B(n_3584), .C(n_2654), .D(n_2702), .Z(n_3586
		));
	notech_and4 i_2435(.A(n_2572), .B(n_2415), .C(n_2309), .D(n_1969), .Z(n_3588
		));
	notech_and4 i_2441(.A(n_2904), .B(n_3588), .C(n_3586), .D(n_2664), .Z(n_3591
		));
	notech_and4 i_1522(.A(n_2572), .B(n_2906), .C(n_2513), .D(n_2918), .Z(n_2921
		));
	notech_or2 i_104572318(.A(n_3957), .B(n_2401), .Z(n_208149053));
	notech_and2 i_186(.A(n_2689), .B(n_2501), .Z(n_3957));
	notech_ao3 i_117072317(.A(n_29924), .B(n_29921), .C(n_3277), .Z(n_207949052
		));
	notech_nao3 i_23111409(.A(n_57905), .B(n_2397), .C(n_2282), .Z(n_1984)
		);
	notech_or4 i_860(.A(n_2282), .B(n_2407), .C(n_57845), .D(n_30107), .Z(n_4079
		));
	notech_and2 i_5672305(.A(n_29962), .B(n_30122), .Z(n_1960));
	notech_and4 i_62525(.A(n_2688), .B(n_2684), .C(n_2662), .D(n_1996), .Z(n_4024
		));
	notech_nor2 i_14(.A(n_2182), .B(n_2185), .Z(n_3971));
	notech_nao3 i_448(.A(modrm[5]), .B(n_29922), .C(n_2325), .Z(n_4027));
	notech_or4 i_23110638(.A(n_2311), .B(n_57905), .C(n_57916), .D(n_30051),
		 .Z(n_4047));
	notech_or2 i_462(.A(n_3957), .B(n_2355), .Z(n_4007));
	notech_or4 i_23111094(.A(n_2383), .B(n_2486), .C(n_2290), .D(n_2292), .Z
		(n_4055));
	notech_and2 i_28472286(.A(n_4022), .B(n_29987), .Z(n_1114));
	notech_or4 i_409(.A(n_2292), .B(n_57925), .C(n_57905), .D(n_30066), .Z(n_4022
		));
	notech_nor2 i_23111397(.A(n_2299), .B(n_2339), .Z(n_4088));
	notech_nor2 i_67172284(.A(n_2101), .B(n_2485), .Z(n_204849027));
	notech_or4 i_359(.A(n_57810), .B(n_2313), .C(n_2389), .D(n_2303), .Z(n_4046
		));
	notech_ao4 i_45772275(.A(n_2118), .B(n_2363), .C(n_2278), .D(n_2339), .Z
		(n_1193));
	notech_or4 i_23111394(.A(n_2339), .B(n_57905), .C(n_57916), .D(n_2271), 
		.Z(n_4044));
	notech_or4 i_8(.A(n_2360), .B(n_2280), .C(n_2282), .D(n_2363), .Z(n_4056
		));
	notech_and4 i_1518(.A(n_4017), .B(n_2915), .C(n_2628), .D(n_3996), .Z(n_2918
		));
	notech_and3 i_55872271(.A(n_4031), .B(n_4036), .C(n_1637), .Z(n_696));
	notech_ao3 i_188(.A(n_29924), .B(n_29956), .C(n_2297), .Z(n_4050));
	notech_nand2 i_63972264(.A(n_3107), .B(n_2614), .Z(n_1086));
	notech_and2 i_68872259(.A(n_4048), .B(n_2195), .Z(n_1925));
	notech_or4 i_23110875(.A(n_57810), .B(n_30110), .C(n_30072), .D(n_57905)
		, .Z(n_4048));
	notech_or4 i_853(.A(n_2311), .B(n_57925), .C(n_57794), .D(n_29995), .Z(n_2305
		));
	notech_or4 i_23110863(.A(n_2286), .B(n_2383), .C(n_30110), .D(n_30072), 
		.Z(n_3993));
	notech_ao3 i_23110755(.A(n_57916), .B(n_57794), .C(n_2464), .Z(n_3969)
		);
	notech_and3 i_79572248(.A(n_4064), .B(n_2377), .C(n_4040), .Z(n_1263));
	notech_or4 i_23110869(.A(n_57810), .B(n_2428), .C(n_57845), .D(n_57820),
		 .Z(n_4040));
	notech_and3 i_816(.A(n_2707), .B(n_2598), .C(n_2704), .Z(n_4071));
	notech_and2 i_541(.A(n_2516), .B(n_3733), .Z(n_4070));
	notech_or4 i_38(.A(n_2410), .B(n_2372), .C(n_4090), .D(n_30117), .Z(n_3984
		));
	notech_and4 i_1515(.A(n_2912), .B(n_2709), .C(n_3980), .D(n_3931), .Z(n_2915
		));
	notech_and4 i_337(.A(n_2310), .B(n_29926), .C(n_57854), .D(n_29919), .Z(n_3974
		));
	notech_or2 i_685(.A(n_2400), .B(n_4072), .Z(n_4030));
	notech_or4 i_23110608(.A(n_2286), .B(n_2311), .C(n_30051), .D(n_30121), 
		.Z(n_4093));
	notech_and4 i_1511(.A(n_2285), .B(n_4014), .C(n_3838), .D(n_2909), .Z(n_2912
		));
	notech_nand3 i_1279(.A(n_57916), .B(n_57904), .C(n_29956), .Z(n_4064));
	notech_or4 i_1053(.A(n_57885), .B(n_57854), .C(n_57872), .D(n_2355), .Z(n_4076
		));
	notech_or4 i_23110878(.A(n_57885), .B(n_2382), .C(n_57854), .D(n_57872),
		 .Z(n_4002));
	notech_or4 i_670(.A(n_2214), .B(n_2497), .C(n_30115), .D(n_30116), .Z(n_4086
		));
	notech_nor2 i_10(.A(n_3935), .B(n_2577), .Z(n_3978));
	notech_or4 i_23111091(.A(n_2360), .B(n_57810), .C(n_2333), .D(n_29968), 
		.Z(n_4026));
	notech_or4 i_11(.A(n_2360), .B(n_2280), .C(n_2282), .D(n_1818), .Z(n_4031
		));
	notech_nor2 i_19(.A(n_4090), .B(n_30057), .Z(n_3986));
	notech_ao3 i_255(.A(n_29924), .B(n_30059), .C(n_2101), .Z(n_4060));
	notech_and4 i_1508(.A(n_4013), .B(n_2255), .C(n_29973), .D(n_29948), .Z(n_2909
		));
	notech_and4 i_1519(.A(n_2162), .B(n_2623), .C(n_4082), .D(n_2019), .Z(n_2906
		));
	notech_or4 i_447(.A(n_57811), .B(n_2519), .C(n_57845), .D(n_30107), .Z(n_4014
		));
	notech_and2 i_412(.A(n_2206), .B(n_4028), .Z(n_2124));
	notech_and2 i_330(.A(n_2359), .B(n_2355), .Z(n_4072));
	notech_and4 i_155(.A(n_3967), .B(n_2171), .C(n_2479), .D(n_2014), .Z(n_2904
		));
	notech_and2 i_613(.A(n_3965), .B(n_3994), .Z(n_2903));
	notech_nao3 i_466(.A(n_30117), .B(n_29922), .C(n_2325), .Z(n_4036));
	notech_ao3 i_93(.A(n_3895), .B(adz), .C(n_2348), .Z(n_4001));
	notech_nor2 i_843(.A(n_2382), .B(n_30057), .Z(n_4080));
	notech_or4 i_139(.A(n_2360), .B(n_57811), .C(n_30004), .D(n_1802), .Z(n_4017
		));
	notech_and3 i_1429(.A(n_2516), .B(n_1890), .C(n_2264), .Z(n_2900));
	notech_or4 i_660(.A(n_2410), .B(n_2037), .C(n_3954), .D(modrm[5]), .Z(n_4053
		));
	notech_and2 i_272(.A(n_2400), .B(n_30053), .Z(n_3958));
	notech_nao3 i_526(.A(n_2397), .B(n_29925), .C(n_2276), .Z(n_4013));
	notech_and2 i_17(.A(n_4067), .B(n_29979), .Z(n_2151));
	notech_or2 i_248(.A(n_3836), .B(n_3957), .Z(n_3994));
	notech_and2 i_772(.A(n_2557), .B(n_2555), .Z(n_2899));
	notech_and4 i_177(.A(n_4008), .B(n_2894), .C(n_29946), .D(n_2895), .Z(n_2898
		));
	notech_ao4 i_239(.A(n_2410), .B(n_2403), .C(n_2325), .D(n_2282), .Z(n_2398
		));
	notech_ao3 i_243(.A(n_2380), .B(n_1951), .C(n_30047), .Z(n_1942));
	notech_and3 i_654(.A(n_2709), .B(n_2071), .C(n_2587), .Z(n_1856));
	notech_and4 i_304(.A(n_2379), .B(n_2699), .C(n_2483), .D(n_1870), .Z(n_1865
		));
	notech_and3 i_260(.A(n_29990), .B(n_1921), .C(n_29962), .Z(n_1834));
	notech_nor2 i_481(.A(n_4057), .B(n_30023), .Z(n_1950));
	notech_and2 i_4450(.A(n_3803), .B(n_3982), .Z(n_1014));
	notech_and2 i_4611(.A(n_4031), .B(n_4036), .Z(n_853));
	notech_and4 i_166(.A(n_4055), .B(n_2538), .C(n_2663), .D(n_3059), .Z(n_872
		));
	notech_and3 i_268(.A(n_2216), .B(n_4037), .C(n_4038), .Z(n_738));
	notech_ao4 i_744(.A(n_3957), .B(n_2485), .C(n_30051), .D(n_2519), .Z(n_811
		));
	notech_and2 i_1433(.A(n_2014), .B(n_2305), .Z(n_2895));
	notech_and4 i_3961(.A(n_3838), .B(n_3973), .C(n_3987), .D(n_4029), .Z(n_2894
		));
	notech_and4 i_162(.A(n_3665), .B(n_1915), .C(n_2212), .D(n_1728), .Z(n_2893
		));
	notech_ao3 i_23111286(.A(n_30115), .B(n_30116), .C(n_2113), .Z(n_4091)
		);
	notech_and4 i_384(.A(n_2654), .B(n_2887), .C(n_1951), .D(n_2619), .Z(n_2890
		));
	notech_and2 i_420(.A(n_2384), .B(n_2382), .Z(n_4090));
	notech_ao3 i_136(.A(n_57925), .B(n_57904), .C(n_2464), .Z(n_4089));
	notech_or4 i_15(.A(n_2315), .B(n_2330), .C(n_2214), .D(n_1900), .Z(n_4087
		));
	notech_or4 i_23111403(.A(n_2289), .B(n_2280), .C(n_2338), .D(n_29925), .Z
		(n_4085));
	notech_nand3 i_274(.A(n_2037), .B(n_2287), .C(n_2375), .Z(n_4084));
	notech_or4 i_33(.A(n_2360), .B(n_57810), .C(n_3935), .D(n_30121), .Z(n_4082
		));
	notech_and2 i_238(.A(n_2517), .B(n_2407), .Z(n_3935));
	notech_and4 i_1439(.A(n_2049), .B(n_2500), .C(n_2510), .D(n_29986), .Z(n_2887
		));
	notech_nao3 i_2969(.A(n_57885), .B(n_2272), .C(n_2403), .Z(n_3733));
	notech_or4 i_1256(.A(n_2282), .B(n_2300), .C(n_30110), .D(n_30072), .Z(n_4067
		));
	notech_or4 i_1265(.A(n_2346), .B(n_2302), .C(n_30117), .D(n_2374), .Z(n_4066
		));
	notech_and2 i_331(.A(n_3277), .B(n_2318), .Z(n_4065));
	notech_or4 i_1294(.A(n_2286), .B(n_2311), .C(n_30051), .D(adz), .Z(n_4062
		));
	notech_or2 i_1295(.A(n_2410), .B(n_2403), .Z(n_4061));
	notech_nor2 i_586(.A(n_3836), .B(n_2101), .Z(n_4059));
	notech_and2 i_207(.A(n_2497), .B(n_2359), .Z(n_3836));
	notech_or4 i_62(.A(n_2276), .B(n_1902), .C(n_2316), .D(n_2289), .Z(n_4058
		));
	notech_ao3 i_23110701(.A(n_57885), .B(n_2272), .C(n_2330), .Z(n_4057));
	notech_ao3 i_201(.A(n_29924), .B(n_29956), .C(n_2275), .Z(n_4054));
	notech_and3 i_355(.A(n_3777), .B(n_4046), .C(n_4034), .Z(n_2884));
	notech_and2 i_332(.A(n_2485), .B(n_2401), .Z(n_3954));
	notech_ao3 i_848(.A(n_29925), .B(n_2296), .C(n_2393), .Z(n_4052));
	notech_or4 i_235(.A(n_2289), .B(n_2338), .C(n_2271), .D(n_2280), .Z(n_4051
		));
	notech_and2 i_487(.A(n_3777), .B(n_4046), .Z(n_2883));
	notech_or2 i_368(.A(n_2285), .B(n_2128), .Z(n_4049));
	notech_ao3 i_23110866(.A(n_57872), .B(n_2324), .C(n_2368), .Z(n_4045));
	notech_or2 i_859(.A(n_2278), .B(n_2337), .Z(n_4043));
	notech_or4 i_669(.A(n_2360), .B(n_57810), .C(n_2486), .D(n_29968), .Z(n_4041
		));
	notech_or2 i_1025(.A(n_2285), .B(n_2095), .Z(n_4038));
	notech_or2 i_35(.A(n_1819), .B(n_2285), .Z(n_4037));
	notech_nor2 i_216(.A(n_2485), .B(n_2215), .Z(n_4035));
	notech_or4 i_25(.A(n_57810), .B(n_2313), .C(n_2389), .D(n_2291), .Z(n_4034
		));
	notech_ao3 i_31(.A(n_29924), .B(n_2349), .C(n_2297), .Z(n_4033));
	notech_or4 i_36(.A(n_2348), .B(n_2360), .C(n_2282), .D(n_1812), .Z(n_4032
		));
	notech_or4 i_23110662(.A(n_2292), .B(n_57925), .C(n_57904), .D(n_29969),
		 .Z(n_4029));
	notech_nand3 i_212(.A(n_29925), .B(n_2530), .C(n_30107), .Z(n_4028));
	notech_or4 i_123(.A(n_2469), .B(n_30060), .C(n_30121), .D(n_30045), .Z(n_4025
		));
	notech_ao3 i_680(.A(modrm[2]), .B(n_2271), .C(n_2564), .Z(n_4023));
	notech_or4 i_1109(.A(n_2347), .B(n_2289), .C(n_3963), .D(n_30111), .Z(n_4020
		));
	notech_and2 i_343(.A(n_30051), .B(n_29995), .Z(n_3963));
	notech_or4 i_23111421(.A(n_2289), .B(n_30004), .C(n_2284), .D(n_2271), .Z
		(n_4019));
	notech_and4 i_23011453(.A(emul), .B(fpu), .C(n_30119), .D(n_2469), .Z(n_4018
		));
	notech_nao3 i_318(.A(n_29924), .B(n_29928), .C(n_2101), .Z(n_4016));
	notech_nor2 i_388(.A(n_3958), .B(n_4072), .Z(n_4015));
	notech_and4 i_1404(.A(n_2834), .B(n_2880), .C(n_2009), .D(n_2010), .Z(n_2881
		));
	notech_and4 i_1403(.A(n_1920), .B(n_2847), .C(n_1870), .D(n_30013), .Z(n_2880
		));
	notech_and4 i_27(.A(emul), .B(fpu), .C(n_30119), .D(n_29923), .Z(n_4011)
		);
	notech_and3 i_23011465(.A(cpl[1]), .B(cpl[0]), .C(ipg_fault), .Z(n_4010)
		);
	notech_and2 i_20(.A(n_29923), .B(ipg_fault), .Z(n_4009));
	notech_or4 i_1117(.A(n_2410), .B(n_2037), .C(n_30117), .D(n_2401), .Z(n_4008
		));
	notech_ao3 i_249(.A(n_57885), .B(n_2272), .C(n_2381), .Z(n_4006));
	notech_nand3 i_133(.A(n_3895), .B(n_57872), .C(n_2324), .Z(n_4005));
	notech_nand2 i_407(.A(n_2330), .B(n_2381), .Z(n_3895));
	notech_or4 i_464(.A(n_57810), .B(n_2519), .C(n_57845), .D(n_57820), .Z(n_4004
		));
	notech_nor2 i_141(.A(n_2244), .B(n_2523), .Z(n_4003));
	notech_and2 i_411(.A(n_2485), .B(n_2497), .Z(n_3845));
	notech_or4 i_217(.A(n_2403), .B(n_2316), .C(n_2311), .D(n_2290), .Z(n_3998
		));
	notech_nao3 i_668(.A(n_29926), .B(adz), .C(n_2519), .Z(n_3996));
	notech_or4 i_1399(.A(n_30075), .B(n_30025), .C(n_2875), .D(n_30029), .Z(n_2878
		));
	notech_or4 i_23111106(.A(n_2289), .B(n_2325), .C(n_2271), .D(n_30051), .Z
		(n_3992));
	notech_or4 i_229(.A(n_2348), .B(n_2360), .C(n_2282), .D(n_2331), .Z(n_3991
		));
	notech_nor2 i_538(.A(n_2278), .B(n_2393), .Z(n_3990));
	notech_or4 i_231(.A(n_57810), .B(n_2316), .C(n_2389), .D(n_2291), .Z(n_3987
		));
	notech_ao3 i_23111160(.A(n_57794), .B(n_57925), .C(n_2318), .Z(n_3985)
		);
	notech_nao3 i_285(.A(n_29924), .B(n_30056), .C(n_2101), .Z(n_3982));
	notech_or4 i_42(.A(n_2311), .B(n_3963), .C(n_57915), .D(n_57794), .Z(n_3981
		));
	notech_or4 i_16(.A(n_57810), .B(n_3935), .C(n_2283), .D(n_30121), .Z(n_3980
		));
	notech_or4 i_125(.A(n_2360), .B(n_57810), .C(n_3935), .D(adz), .Z(n_3979
		));
	notech_or4 i_370(.A(n_2290), .B(n_2292), .C(n_2383), .D(n_2333), .Z(n_3977
		));
	notech_or4 i_498(.A(n_2360), .B(n_57810), .C(n_2325), .D(n_2299), .Z(n_3975
		));
	notech_nao3 i_2992(.A(modrm[2]), .B(n_2530), .C(n_29925), .Z(n_3973));
	notech_or4 i_51(.A(n_2410), .B(n_2373), .C(n_4090), .D(n_30117), .Z(n_3972
		));
	notech_or4 i_23110590(.A(n_2360), .B(n_57810), .C(n_2289), .D(n_2410), .Z
		(n_3970));
	notech_ao3 i_23110725(.A(n_57885), .B(n_2272), .C(n_2368), .Z(n_3968));
	notech_or4 i_338(.A(n_57810), .B(n_2316), .C(n_30004), .D(n_2303), .Z(n_3967
		));
	notech_or4 i_128(.A(n_30004), .B(n_57915), .C(n_57794), .D(n_29995), .Z(n_3965
		));
	notech_or4 i_23110593(.A(n_57811), .B(n_2621), .C(n_57820), .D(n_30108),
		 .Z(n_3964));
	notech_and2 i_147(.A(n_3867), .B(n_1875), .Z(n_2380));
	notech_or4 i_1297(.A(n_57915), .B(n_57794), .C(adz), .D(n_30060), .Z(n_3867
		));
	notech_and2 i_3098(.A(n_4062), .B(n_4093), .Z(n_2366));
	notech_ao3 i_30(.A(n_30108), .B(n_30107), .C(n_57811), .Z(n_2354));
	notech_ao3 i_37(.A(n_30108), .B(n_57820), .C(n_57811), .Z(n_2369));
	notech_nand2 i_3157(.A(n_2327), .B(n_29958), .Z(n_2307));
	notech_or4 i_1392(.A(n_30041), .B(n_30071), .C(n_2873), .D(n_30015), .Z(n_2875
		));
	notech_and2 i_415(.A(n_2286), .B(n_2290), .Z(n_3961));
	notech_ao3 i_256(.A(n_2385), .B(n_30117), .C(n_2410), .Z(n_3959));
	notech_ao3 i_89(.A(n_30115), .B(modrm[4]), .C(n_2214), .Z(n_2210));
	notech_or4 i_3282(.A(n_2386), .B(n_57925), .C(n_57794), .D(n_30110), .Z(n_2182
		));
	notech_or4 i_3297(.A(n_2386), .B(n_57915), .C(n_57794), .D(n_30110), .Z(n_2167
		));
	notech_nand2 i_3299(.A(n_29992), .B(n_29957), .Z(n_2165));
	notech_nand3 i_1388(.A(n_2538), .B(n_2111), .C(n_2872), .Z(n_2873));
	notech_or4 i_110(.A(n_2280), .B(n_2282), .C(n_57820), .D(n_30108), .Z(n_2118
		));
	notech_or4 i_3446(.A(n_57915), .B(n_57794), .C(n_2271), .D(n_30073), .Z(n_2018
		));
	notech_and4 i_1384(.A(n_1815), .B(n_4005), .C(n_2870), .D(n_2789), .Z(n_2872
		));
	notech_nor2 i_23111376(.A(n_2564), .B(n_2271), .Z(n_1987));
	notech_and2 i_12(.A(n_4025), .B(n_29989), .Z(n_1953));
	notech_and4 i_23110713(.A(adz), .B(n_2296), .C(n_2469), .D(n_2466), .Z(n_3950
		));
	notech_and4 i_1381(.A(n_2171), .B(n_2867), .C(n_2857), .D(n_2022), .Z(n_2870
		));
	notech_and3 i_3727(.A(n_3996), .B(n_2579), .C(n_4082), .Z(n_1737));
	notech_and4 i_1377(.A(n_1656), .B(n_2627), .C(n_2863), .D(n_1623), .Z(n_2867
		));
	notech_nand3 i_699(.A(n_4031), .B(n_4056), .C(n_2611), .Z(n_3956));
	notech_and2 i_3849(.A(n_3838), .B(n_4028), .Z(n_1615));
	notech_nand3 i_198(.A(n_29925), .B(n_30107), .C(n_2536), .Z(n_3838));
	notech_and4 i_3919(.A(n_2579), .B(n_1970), .C(n_3998), .D(n_29990), .Z(n_1545
		));
	notech_and2 i_72(.A(n_2063), .B(n_2969), .Z(n_3955));
	notech_or4 i_861(.A(n_57811), .B(n_2865), .C(n_57820), .D(n_30108), .Z(n_3803
		));
	notech_and2 i_4744(.A(n_3739), .B(n_2195), .Z(n_720));
	notech_or4 i_467(.A(n_57881), .B(n_57854), .C(n_57872), .D(n_2401), .Z(n_3739
		));
	notech_or2 i_273(.A(n_1858), .B(n_3963), .Z(n_3880));
	notech_and3 i_5210(.A(n_1829), .B(n_1828), .C(n_4084), .Z(n_254));
	notech_nand3 i_4(.A(n_57881), .B(n_57854), .C(n_57872), .Z(n_2410));
	notech_or4 i_1350(.A(n_2347), .B(n_2244), .C(n_30111), .D(adz), .Z(n_2865
		));
	notech_nand3 i_60(.A(n_57916), .B(n_57904), .C(n_29925), .Z(n_2302));
	notech_nand3 i_65(.A(n_57925), .B(n_57904), .C(n_29925), .Z(n_2275));
	notech_nao3 i_23(.A(n_30107), .B(n_57845), .C(n_57811), .Z(n_2383));
	notech_or4 i_18(.A(n_2372), .B(n_2214), .C(n_2330), .D(n_2504), .Z(n_3931
		));
	notech_and2 i_21(.A(n_30122), .B(n_1919), .Z(n_1951));
	notech_and2 i_22(.A(n_223489126), .B(n_1792), .Z(n_2017));
	notech_and3 i_24(.A(n_57885), .B(n_30111), .C(n_30110), .Z(n_2397));
	notech_nand3 i_61(.A(n_57794), .B(n_57925), .C(n_29925), .Z(n_2278));
	notech_and3 i_76(.A(n_57916), .B(n_57794), .C(n_29925), .Z(n_3908));
	notech_ao4 i_26(.A(n_2278), .B(n_2458), .C(n_2455), .D(n_29968), .Z(n_2123
		));
	notech_and2 i_29(.A(n_2141), .B(n_4013), .Z(n_2065));
	notech_nand2 i_74(.A(opz[1]), .B(n_2322), .Z(n_2320));
	notech_and2 i_34(.A(n_4031), .B(n_4056), .Z(n_2116));
	notech_and4 i_1374(.A(n_3964), .B(n_4004), .C(n_2860), .D(n_2676), .Z(n_2863
		));
	notech_and2 i_53(.A(n_2192), .B(n_4017), .Z(n_2176));
	notech_and2 i_57(.A(n_2071), .B(n_1835), .Z(n_2171));
	notech_and3 i_58(.A(n_2233), .B(n_1938), .C(n_4079), .Z(n_2049));
	notech_and3 i_80(.A(n_2629), .B(n_29975), .C(n_29973), .Z(n_2357));
	notech_and4 i_1371(.A(n_2435), .B(n_3998), .C(n_2008), .D(n_2630), .Z(n_2860
		));
	notech_nand3 i_97(.A(n_2062), .B(adz), .C(n_29926), .Z(n_3890));
	notech_nand3 i_122(.A(n_29992), .B(n_29957), .C(n_29991), .Z(n_2164));
	notech_or4 i_167(.A(n_57811), .B(n_2316), .C(n_30004), .D(n_2291), .Z(n_3876
		));
	notech_ao4 i_130(.A(n_2278), .B(n_2346), .C(n_2275), .D(n_2393), .Z(n_1958
		));
	notech_or4 i_131(.A(fpu), .B(twobyte), .C(ipg_fault), .D(op[7]), .Z(n_2403
		));
	notech_and4 i_135(.A(n_2623), .B(n_3964), .C(n_3965), .D(n_2380), .Z(n_2332
		));
	notech_and3 i_146(.A(n_2327), .B(n_29958), .C(n_2305), .Z(n_2304));
	notech_and2 i_160(.A(n_1918), .B(n_1794), .Z(n_1978));
	notech_ao3 i_704(.A(n_4014), .B(n_1921), .C(n_29927), .Z(n_2857));
	notech_and4 i_170(.A(n_3876), .B(n_2609), .C(n_2663), .D(n_2500), .Z(n_901
		));
	notech_and4 i_175(.A(n_1874), .B(n_2702), .C(n_2900), .D(n_29931), .Z(n_1504
		));
	notech_nand2 i_182(.A(n_30116), .B(modrm[3]), .Z(n_2315));
	notech_and4 i_191(.A(n_57885), .B(n_30111), .C(n_57872), .D(n_2369), .Z(n_3846
		));
	notech_and2 i_204(.A(n_3994), .B(n_29960), .Z(n_1999));
	notech_ao4 i_208(.A(n_2290), .B(n_2447), .C(n_29995), .D(n_2448), .Z(n_2327
		));
	notech_and2 i_211(.A(n_2308), .B(n_2294), .Z(n_2058));
	notech_or4 i_469(.A(n_2410), .B(n_2315), .C(n_2382), .D(n_30117), .Z(n_3834
		));
	notech_and2 i_214(.A(n_3996), .B(n_4082), .Z(n_1972));
	notech_and3 i_220(.A(n_4002), .B(n_1797), .C(n_4017), .Z(n_1777));
	notech_and4 i_309(.A(n_2638), .B(n_2014), .C(n_2192), .D(n_29944), .Z(n_2854
		));
	notech_ao4 i_225(.A(n_1879), .B(n_2488), .C(n_2037), .D(n_2489), .Z(n_2024
		));
	notech_and2 i_240(.A(n_4014), .B(n_2005), .Z(n_1624));
	notech_and2 i_241(.A(n_2057), .B(n_1794), .Z(n_1290));
	notech_nor2 i_862(.A(n_2400), .B(n_2098), .Z(n_3820));
	notech_and2 i_252(.A(n_1985), .B(n_29977), .Z(n_1678));
	notech_and4 i_364(.A(n_2394), .B(n_1958), .C(n_2065), .D(n_2285), .Z(n_2852
		));
	notech_and4 i_261(.A(n_2094), .B(n_4026), .C(n_2155), .D(n_1825), .Z(n_497
		));
	notech_and4 i_263(.A(n_2394), .B(n_1958), .C(n_2026), .D(n_2925), .Z(n_1434
		));
	notech_and4 i_265(.A(n_2179), .B(n_3312), .C(n_3179), .D(n_2180), .Z(n_493
		));
	notech_and4 i_267(.A(n_2398), .B(n_1545), .C(n_29972), .D(n_29951), .Z(n_68
		));
	notech_and4 i_270(.A(n_2639), .B(n_3184), .C(n_3179), .D(n_2937), .Z(n_537
		));
	notech_and2 i_271(.A(n_29955), .B(n_29954), .Z(n_2099));
	notech_ao4 i_278(.A(n_2244), .B(n_2523), .C(n_30053), .D(n_2485), .Z(n_2212
		));
	notech_and2 i_279(.A(n_4041), .B(n_1896), .Z(n_2094));
	notech_and3 i_280(.A(n_1993), .B(n_2665), .C(n_2688), .Z(n_1718));
	notech_and3 i_289(.A(n_2046), .B(n_1912), .C(n_1914), .Z(n_1993));
	notech_and2 i_295(.A(n_2136), .B(n_2978), .Z(n_1329));
	notech_and2 i_299(.A(n_3803), .B(n_29988), .Z(n_1623));
	notech_and4 i_477(.A(n_2151), .B(n_2166), .C(n_2588), .D(n_1890), .Z(n_2850
		));
	notech_and4 i_305(.A(n_2678), .B(n_2791), .C(n_1857), .D(n_533), .Z(n_530
		));
	notech_and4 i_1396(.A(n_2707), .B(n_2352), .C(n_2839), .D(n_2844), .Z(n_2847
		));
	notech_and2 i_314(.A(n_3977), .B(n_4086), .Z(n_1332));
	notech_and4 i_323(.A(n_208149053), .B(n_4049), .C(n_29955), .D(n_3981), 
		.Z(n_444));
	notech_and3 i_324(.A(n_2663), .B(n_2183), .C(n_3422), .Z(n_204));
	notech_and2 i_333(.A(n_4032), .B(n_2365), .Z(n_1905));
	notech_ao4 i_341(.A(n_2400), .B(n_3845), .C(n_3958), .D(n_2401), .Z(n_2157
		));
	notech_and4 i_357(.A(n_3996), .B(n_4014), .C(n_4082), .D(n_3980), .Z(n_1970
		));
	notech_or4 i_360(.A(n_57811), .B(n_2316), .C(n_2389), .D(n_2303), .Z(n_3779
		));
	notech_or4 i_406(.A(n_2389), .B(n_2290), .C(n_2292), .D(n_29995), .Z(n_3777
		));
	notech_and4 i_1391(.A(n_2465), .B(n_2198), .C(n_2842), .D(n_2831), .Z(n_2844
		));
	notech_or4 i_367(.A(n_3956), .B(n_30044), .C(n_30012), .D(n_30038), .Z(n_3773
		));
	notech_and3 i_371(.A(n_2157), .B(n_1930), .C(n_2625), .Z(n_1870));
	notech_and4 i_1386(.A(n_4084), .B(n_2377), .C(n_2827), .D(n_1712), .Z(n_2842
		));
	notech_and3 i_379(.A(n_2231), .B(n_1833), .C(n_1936), .Z(n_1780));
	notech_and4 i_381(.A(n_3739), .B(n_2195), .C(n_2264), .D(n_719), .Z(n_717
		));
	notech_mux2 i_391(.S(n_57820), .A(modrm[0]), .B(modrm[3]), .Z(n_3763));
	notech_nor2 i_395(.A(n_2301), .B(n_3908), .Z(n_3761));
	notech_mux2 i_397(.S(n_57820), .A(n_30115), .B(n_30113), .Z(n_3760));
	notech_nao3 i_401(.A(n_57872), .B(n_30117), .C(n_2386), .Z(n_2214));
	notech_and3 i_402(.A(n_223489126), .B(n_1792), .C(n_29965), .Z(n_2015)
		);
	notech_and2 i_413(.A(n_3838), .B(n_3973), .Z(n_2076));
	notech_and3 i_421(.A(n_4062), .B(n_4093), .C(n_29961), .Z(n_2022));
	notech_nao3 i_852(.A(n_2385), .B(n_30056), .C(n_2214), .Z(n_3751));
	notech_and2 i_425(.A(n_3751), .B(n_29989), .Z(n_1526));
	notech_and2 i_428(.A(n_4055), .B(n_1857), .Z(n_2029));
	notech_and2 i_437(.A(n_29980), .B(n_29960), .Z(n_1728));
	notech_ao4 i_440(.A(n_2501), .B(n_2382), .C(n_57811), .D(n_2646), .Z(n_733
		));
	notech_and4 i_310(.A(n_4002), .B(n_2195), .C(n_2414), .D(n_2597), .Z(n_2839
		));
	notech_and2 i_454(.A(n_2073), .B(n_2202), .Z(n_2162));
	notech_and4 i_455(.A(n_3979), .B(n_1970), .C(n_29988), .D(n_1978), .Z(n_1969
		));
	notech_and2 i_474(.A(n_3979), .B(n_3980), .Z(n_1816));
	notech_or4 i_835(.A(n_2214), .B(n_2384), .C(modrm[3]), .D(n_30116), .Z(n_3736
		));
	notech_and2 i_476(.A(n_2587), .B(n_1851), .Z(n_1603));
	notech_nand2 i_479(.A(n_3998), .B(n_29990), .Z(n_1967));
	notech_and4 i_492(.A(n_3967), .B(n_3987), .C(n_1796), .D(n_4029), .Z(n_3728
		));
	notech_or4 i_493(.A(n_57811), .B(n_2286), .C(n_57845), .D(n_30107), .Z(n_2368
		));
	notech_and3 i_501(.A(n_29972), .B(n_29951), .C(n_2305), .Z(n_1924));
	notech_and2 i_508(.A(n_2327), .B(n_4047), .Z(n_1923));
	notech_and4 i_515(.A(n_29978), .B(n_1958), .C(n_2377), .D(n_29959), .Z(n_960
		));
	notech_nao3 i_532(.A(n_29925), .B(n_2375), .C(n_2286), .Z(n_2113));
	notech_and2 i_792(.A(n_2411), .B(n_1603), .Z(n_2834));
	notech_or4 i_536(.A(n_57885), .B(n_2338), .C(n_57872), .D(n_30111), .Z(n_2234
		));
	notech_and2 i_545(.A(n_2216), .B(n_30058), .Z(n_1656));
	notech_and2 i_550(.A(n_2132), .B(n_2789), .Z(n_455));
	notech_and4 i_555(.A(n_4027), .B(n_4036), .C(n_4076), .D(n_2091), .Z(n_894
		));
	notech_and4 i_562(.A(n_2233), .B(n_1938), .C(n_4079), .D(n_4058), .Z(n_2047
		));
	notech_and3 i_567(.A(n_3838), .B(n_3973), .C(n_1798), .Z(n_3697));
	notech_and3 i_692(.A(n_4025), .B(n_29989), .C(n_2357), .Z(n_2831));
	notech_and2 i_606(.A(n_2380), .B(n_30122), .Z(n_1593));
	notech_and3 i_94(.A(n_3992), .B(n_1895), .C(n_1831), .Z(n_2829));
	notech_ao4 i_604(.A(n_2387), .B(n_30055), .C(n_2382), .D(n_30057), .Z(n_2827
		));
	notech_ao4 i_618(.A(n_30051), .B(n_2407), .C(n_2485), .D(n_30053), .Z(n_1306
		));
	notech_and2 i_625(.A(n_3982), .B(n_29958), .Z(n_1537));
	notech_and3 i_634(.A(n_3993), .B(n_4040), .C(n_2103), .Z(n_730));
	notech_and3 i_637(.A(n_3992), .B(n_2123), .C(n_29946), .Z(n_1712));
	notech_and4 i_780(.A(n_1949), .B(n_1796), .C(n_3880), .D(n_29931), .Z(n_2826
		));
	notech_or2 i_658(.A(n_3958), .B(n_2355), .Z(n_3672));
	notech_or4 i_659(.A(n_2316), .B(n_2276), .C(n_2373), .D(n_2333), .Z(n_2052
		));
	notech_or2 i_684(.A(n_2400), .B(n_2359), .Z(n_3665));
	notech_ao4 i_708(.A(n_2400), .B(n_3845), .C(n_30060), .D(n_2286), .Z(n_1543
		));
	notech_or4 i_729(.A(n_4010), .B(n_4018), .C(n_3950), .D(n_4015), .Z(n_1262
		));
	notech_and2 i_736(.A(n_3979), .B(n_4032), .Z(n_861));
	notech_and2 i_748(.A(n_2246), .B(n_1984), .Z(n_520));
	notech_and2 i_750(.A(n_2665), .B(n_2394), .Z(n_719));
	notech_and3 i_751(.A(n_2790), .B(n_1993), .C(n_3105), .Z(n_703));
	notech_ao4 i_753(.A(n_2291), .B(n_30066), .C(n_2118), .D(n_2363), .Z(n_673
		));
	notech_and2 i_755(.A(n_4002), .B(n_4048), .Z(n_2080));
	notech_ao4 i_757(.A(n_2422), .B(n_2384), .C(n_2499), .D(n_2382), .Z(n_574
		));
	notech_and2 i_768(.A(n_1936), .B(n_29951), .Z(n_215));
	notech_and3 i_769(.A(n_4041), .B(n_4036), .C(n_2056), .Z(n_1284));
	notech_and3 i_779(.A(n_3880), .B(n_3374), .C(n_2213), .Z(n_218));
	notech_and2 i_781(.A(n_2206), .B(n_733), .Z(n_709));
	notech_and3 i_782(.A(n_2625), .B(n_3779), .C(n_2073), .Z(n_533));
	notech_and3 i_791(.A(n_3979), .B(n_3980), .C(n_4082), .Z(n_1815));
	notech_or4 i_1318(.A(n_30079), .B(n_2817), .C(n_1998), .D(n_2000), .Z(n_2820
		));
	notech_and3 i_804(.A(n_4055), .B(n_2538), .C(n_3834), .Z(n_1340));
	notech_and3 i_810(.A(n_2166), .B(n_2108), .C(n_2380), .Z(n_466));
	notech_and3 i_812(.A(n_1886), .B(n_2686), .C(n_1887), .Z(n_2246));
	notech_and4 i_813(.A(n_3834), .B(n_2036), .C(n_1924), .D(n_3984), .Z(n_1920
		));
	notech_and3 i_818(.A(n_2025), .B(n_2103), .C(n_4027), .Z(n_1346));
	notech_and4 i_2932(.A(n_4047), .B(n_2091), .C(n_1999), .D(n_29980), .Z(n_1996
		));
	notech_or4 i_1315(.A(n_30020), .B(n_30037), .C(n_30074), .D(n_2814), .Z(n_2817
		));
	notech_nao3 i_1313(.A(n_1678), .B(n_2588), .C(n_2812), .Z(n_2814));
	notech_or4 i_1311(.A(n_1997), .B(n_30049), .C(n_2809), .D(n_2078), .Z(n_2812
		));
	notech_nao3 i_1308(.A(n_3777), .B(n_2808), .C(n_222391112), .Z(n_2809)
		);
	notech_and4 i_1307(.A(n_3665), .B(n_1923), .C(n_2804), .D(n_29985), .Z(n_2808
		));
	notech_and4 i_1304(.A(n_2627), .B(n_1995), .C(n_3965), .D(n_2801), .Z(n_2804
		));
	notech_ao3 i_1300(.A(n_2799), .B(n_2216), .C(n_1933), .Z(n_2801));
	notech_and4 i_1298(.A(n_2516), .B(n_2797), .C(n_3998), .D(n_2794), .Z(n_2799
		));
	notech_and4 i_1292(.A(n_29975), .B(n_29973), .C(n_1990), .D(n_1994), .Z(n_2797
		));
	notech_ao4 i_1290(.A(n_57916), .B(n_2734), .C(n_2140), .D(n_57794), .Z(n_2794
		));
	notech_and2 i_237(.A(n_2791), .B(n_2790), .Z(n_2792));
	notech_ao4 i_486(.A(n_2384), .B(n_30053), .C(n_2403), .D(n_30004), .Z(n_2791
		));
	notech_and2 i_43(.A(n_2789), .B(n_1982), .Z(n_2790));
	notech_and3 i_349(.A(n_1901), .B(n_4087), .C(n_3931), .Z(n_2789));
	notech_or4 i_1262(.A(n_222991118), .B(n_1975), .C(n_1976), .D(n_2782), .Z
		(n_2785));
	notech_nand3 i_1259(.A(n_2780), .B(n_2729), .C(n_222791116), .Z(n_2782)
		);
	notech_and4 i_1257(.A(n_2778), .B(n_2212), .C(n_29946), .D(n_2532), .Z(n_2780
		));
	notech_and4 i_1254(.A(n_2765), .B(n_1978), .C(n_2136), .D(n_2777), .Z(n_2778
		));
	notech_and4 i_1253(.A(n_2192), .B(n_2775), .C(n_2744), .D(n_2305), .Z(n_2777
		));
	notech_and4 i_1248(.A(n_1877), .B(n_2772), .C(n_3996), .D(n_29957), .Z(n_2775
		));
	notech_and4 i_1245(.A(n_2768), .B(n_3993), .C(n_2771), .D(n_29990), .Z(n_2772
		));
	notech_ao4 i_1244(.A(n_2458), .B(n_2299), .C(n_2383), .D(n_2621), .Z(n_2771
		));
	notech_ao4 i_1240(.A(n_2734), .B(n_30107), .C(n_2140), .D(n_30110), .Z(n_2768
		));
	notech_and3 i_173(.A(n_2216), .B(n_2733), .C(n_2730), .Z(n_2765));
	notech_and4 i_3740(.A(n_223489126), .B(n_1792), .C(n_2151), .D(n_29965),
		 .Z(n_2760));
	notech_and4 i_226(.A(n_29980), .B(n_29960), .C(n_2091), .D(n_3994), .Z(n_2759
		));
	notech_and2 i_478(.A(n_1993), .B(n_2665), .Z(n_2757));
	notech_and4 i_1213(.A(n_2751), .B(n_222791116), .C(n_2729), .D(n_1955), 
		.Z(n_2754));
	notech_and4 i_1210(.A(n_30063), .B(n_2749), .C(n_29990), .D(n_1954), .Z(n_2751
		));
	notech_and4 i_1208(.A(n_1930), .B(n_2741), .C(n_2747), .D(n_1737), .Z(n_2749
		));
	notech_and4 i_1206(.A(n_1949), .B(n_2744), .C(n_1952), .D(n_2743), .Z(n_2747
		));
	notech_and2 i_251(.A(n_1932), .B(n_30021), .Z(n_2744));
	notech_and2 i_138(.A(n_2192), .B(n_2305), .Z(n_2743));
	notech_and4 i_1203(.A(n_2730), .B(n_2731), .C(n_3965), .D(n_2739), .Z(n_2741
		));
	notech_and4 i_1200(.A(n_3993), .B(n_3992), .C(n_2736), .D(n_3980), .Z(n_2739
		));
	notech_and3 i_1194(.A(n_2733), .B(n_2234), .C(n_1947), .Z(n_2736));
	notech_ao4 i_218(.A(n_2403), .B(n_2389), .C(n_57811), .D(n_2646), .Z(n_2734
		));
	notech_ao4 i_543(.A(n_29995), .B(n_2446), .C(n_2325), .D(n_2282), .Z(n_2733
		));
	notech_ao4 i_1196(.A(n_2166), .B(n_30090), .C(n_2290), .D(n_2464), .Z(n_2731
		));
	notech_ao4 i_696(.A(n_2318), .B(n_2286), .C(n_29995), .D(n_2519), .Z(n_2730
		));
	notech_and4 i_157(.A(n_4084), .B(n_2377), .C(n_3751), .D(n_2727), .Z(n_2729
		));
	notech_ao4 i_1154(.A(n_2118), .B(n_2027), .C(n_2362), .D(n_2331), .Z(n_2727
		));
	notech_and4 i_1173(.A(n_29978), .B(n_1780), .C(n_2395), .D(n_2414), .Z(n_2726
		));
	notech_and2 i_485(.A(n_4002), .B(n_1797), .Z(n_2723));
	notech_and3 i_300(.A(n_3967), .B(n_2171), .C(n_2479), .Z(n_2722));
	notech_and4 i_1182(.A(n_2141), .B(n_4013), .C(n_2015), .D(n_1941), .Z(n_2719
		));
	notech_and4 i_348(.A(n_2195), .B(n_2714), .C(n_2611), .D(n_2713), .Z(n_2717
		));
	notech_ao4 i_1177(.A(n_2384), .B(n_1937), .C(n_2052), .D(n_2331), .Z(n_2714
		));
	notech_and2 i_701(.A(n_4016), .B(n_3972), .Z(n_2713));
	notech_and2 i_452(.A(n_1798), .B(n_2111), .Z(n_2709));
	notech_and4 i_387(.A(n_2190), .B(n_3973), .C(n_2463), .D(n_2675), .Z(n_2707
		));
	notech_and2 i_646(.A(n_2703), .B(n_2543), .Z(n_2704));
	notech_and4 i_473(.A(n_1873), .B(n_2555), .C(n_1874), .D(n_2702), .Z(n_2703
		));
	notech_and2 i_233(.A(n_1800), .B(n_2563), .Z(n_2702));
	notech_and4 i_1127(.A(n_2417), .B(n_2695), .C(n_2198), .D(n_2696), .Z(n_2699
		));
	notech_and4 i_1124(.A(n_2073), .B(n_4067), .C(n_2202), .D(n_29979), .Z(n_2696
		));
	notech_and2 i_399(.A(n_1796), .B(n_4029), .Z(n_2695));
	notech_and2 i_566(.A(n_2157), .B(n_1930), .Z(n_2694));
	notech_and3 i_3466(.A(n_3994), .B(n_29960), .C(n_29980), .Z(n_2690));
	notech_or4 i_101(.A(n_2386), .B(n_2037), .C(n_30110), .D(n_30117), .Z(n_2689
		));
	notech_and2 i_288(.A(n_2246), .B(n_2264), .Z(n_2688));
	notech_ao4 i_376(.A(n_2553), .B(n_2685), .C(n_2557), .D(n_2037), .Z(n_2686
		));
	notech_nand2 i_936(.A(n_1885), .B(modrm[1]), .Z(n_2685));
	notech_and4 i_711(.A(n_2681), .B(n_2675), .C(n_2665), .D(n_2664), .Z(n_2684
		));
	notech_and4 i_1021(.A(n_2179), .B(n_2678), .C(n_2457), .D(n_2022), .Z(n_2681
		));
	notech_and3 i_193(.A(n_2676), .B(n_2189), .C(n_2190), .Z(n_2678));
	notech_and2 i_54(.A(n_2188), .B(n_1907), .Z(n_2676));
	notech_and4 i_358(.A(n_4055), .B(n_1857), .C(n_3977), .D(n_2673), .Z(n_2675
		));
	notech_and4 i_877(.A(n_1855), .B(n_1854), .C(n_2668), .D(n_2238), .Z(n_2673
		));
	notech_ao4 i_137(.A(n_2667), .B(n_2300), .C(n_2666), .D(n_2292), .Z(n_2668
		));
	notech_nand2 i_868(.A(n_2530), .B(n_57820), .Z(n_2667));
	notech_nand2 i_867(.A(n_30107), .B(n_2536), .Z(n_2666));
	notech_and2 i_758(.A(n_2024), .B(n_1911), .Z(n_2665));
	notech_and2 i_614(.A(n_2663), .B(n_2352), .Z(n_2664));
	notech_ao4 i_52(.A(n_2291), .B(n_2052), .C(n_2278), .D(n_2337), .Z(n_2663
		));
	notech_and4 i_1111(.A(n_2484), .B(n_2549), .C(n_2483), .D(n_2661), .Z(n_2662
		));
	notech_and4 i_1108(.A(n_2658), .B(n_2619), .C(n_2607), .D(n_2567), .Z(n_2661
		));
	notech_and4 i_1100(.A(n_2654), .B(n_2157), .C(n_2650), .D(n_2656), .Z(n_2658
		));
	notech_and2 i_602(.A(n_2655), .B(n_4025), .Z(n_2656));
	notech_ao4 i_356(.A(n_2391), .B(n_2303), .C(n_2291), .D(n_29969), .Z(n_2655
		));
	notech_and2 i_293(.A(n_2030), .B(n_3991), .Z(n_2654));
	notech_and4 i_1093(.A(n_2648), .B(n_2643), .C(n_2304), .D(n_2620), .Z(n_2650
		));
	notech_and4 i_383(.A(n_4002), .B(n_4048), .C(n_2076), .D(n_29946), .Z(n_2648
		));
	notech_or4 i_997(.A(n_57885), .B(n_57854), .C(n_30110), .D(n_57904), .Z(n_2646
		));
	notech_and4 i_1087(.A(n_2625), .B(n_2634), .C(n_2332), .D(n_2641), .Z(n_2643
		));
	notech_and4 i_1084(.A(n_4058), .B(n_2049), .C(n_2639), .D(n_3981), .Z(n_2641
		));
	notech_and2 i_242(.A(n_2638), .B(n_2014), .Z(n_2639));
	notech_ao4 i_215(.A(n_2325), .B(n_2384), .C(n_2383), .D(n_2428), .Z(n_2638
		));
	notech_and2 i_616(.A(n_2233), .B(n_1938), .Z(n_2637));
	notech_and4 i_1081(.A(n_2631), .B(n_2628), .C(n_2357), .D(n_29989), .Z(n_2634
		));
	notech_and3 i_302(.A(n_2433), .B(n_2140), .C(n_4064), .Z(n_2631));
	notech_and2 i_569(.A(n_2433), .B(n_2140), .Z(n_2630));
	notech_nor2 i_426(.A(n_4010), .B(n_4018), .Z(n_2629));
	notech_and3 i_774(.A(n_3993), .B(n_4040), .C(n_3733), .Z(n_2628));
	notech_and2 i_410(.A(n_3993), .B(n_4040), .Z(n_2627));
	notech_and2 i_134(.A(n_1877), .B(n_1831), .Z(n_2625));
	notech_and2 i_45(.A(n_29972), .B(n_29951), .Z(n_2623));
	notech_or4 i_923(.A(n_2386), .B(n_30110), .C(n_57925), .D(n_57905), .Z(n_2621
		));
	notech_and2 i_509(.A(n_3987), .B(n_4029), .Z(n_2620));
	notech_and4 i_36690983(.A(n_2611), .B(n_2379), .C(n_2614), .D(n_2616), .Z
		(n_2619));
	notech_and4 i_978(.A(n_4027), .B(n_4036), .C(n_29955), .D(n_29954), .Z(n_2616
		));
	notech_and2 i_783(.A(n_4027), .B(n_4036), .Z(n_2615));
	notech_and3 i_430(.A(n_4041), .B(n_1896), .C(n_4026), .Z(n_2614));
	notech_and4 i_196(.A(n_4044), .B(n_2609), .C(n_2108), .D(n_29987), .Z(n_2611
		));
	notech_and4 i_802(.A(n_4044), .B(n_4051), .C(n_29987), .D(n_4085), .Z(n_2610
		));
	notech_and2 i_458(.A(n_4051), .B(n_4085), .Z(n_2609));
	notech_and4 i_1102(.A(n_2572), .B(n_1969), .C(n_2605), .D(n_2309), .Z(n_2607
		));
	notech_and4 i_63(.A(n_2591), .B(n_2602), .C(n_2588), .D(n_2587), .Z(n_2605
		));
	notech_and4 i_1076(.A(n_3931), .B(n_2598), .C(n_2171), .D(n_2601), .Z(n_2602
		));
	notech_and3 i_1075(.A(n_2192), .B(n_4017), .C(n_2195), .Z(n_2601));
	notech_and3 i_199(.A(n_2103), .B(n_2159), .C(n_1851), .Z(n_2598));
	notech_and2 i_830(.A(n_2103), .B(n_2159), .Z(n_2597));
	notech_or4 i_823(.A(n_57811), .B(n_2486), .C(n_57845), .D(n_30107), .Z(n_2596
		));
	notech_or4 i_863(.A(n_2302), .B(n_57872), .C(n_30072), .D(modrm[5]), .Z(n_2594
		));
	notech_and4 i_787(.A(n_2162), .B(n_29992), .C(n_29957), .D(n_29991), .Z(n_2591
		));
	notech_and3 i_598(.A(n_3970), .B(n_1806), .C(n_29962), .Z(n_2588));
	notech_and2 i_152(.A(n_1825), .B(n_2070), .Z(n_2587));
	notech_or4 i_1069(.A(n_57811), .B(n_2283), .C(n_30004), .D(n_30117), .Z(n_2586
		));
	notech_and3 i_223(.A(n_3979), .B(n_29988), .C(n_1978), .Z(n_2579));
	notech_or4 i_910(.A(n_57811), .B(n_30108), .C(n_30107), .D(adz), .Z(n_2577
		));
	notech_or4 i_663(.A(n_57885), .B(n_57872), .C(n_30111), .D(n_30045), .Z(n_2574
		));
	notech_and4 i_378(.A(n_1984), .B(n_1801), .C(n_4019), .D(n_30058), .Z(n_2572
		));
	notech_and2 i_517(.A(n_1984), .B(n_1801), .Z(n_2571));
	notech_and2 i_3478(.A(n_4019), .B(n_30058), .Z(n_2569));
	notech_and3 i_377(.A(n_2565), .B(n_2563), .C(n_2562), .Z(n_2567));
	notech_and3 i_759(.A(n_4067), .B(n_2166), .C(n_29979), .Z(n_2565));
	notech_or4 i_499(.A(n_57885), .B(n_2282), .C(n_57854), .D(n_30110), .Z(n_2564
		));
	notech_ao4 i_442(.A(n_2494), .B(n_2315), .C(n_2489), .D(n_2373), .Z(n_2563
		));
	notech_and4 i_723(.A(n_1873), .B(n_2555), .C(n_1874), .D(n_1800), .Z(n_2562
		));
	notech_or4 i_108(.A(n_2497), .B(n_2333), .C(modrm[1]), .D(modrm[0]), .Z(n_2560
		));
	notech_or4 i_109(.A(n_2497), .B(n_2333), .C(modrm[1]), .D(n_30113), .Z(n_2557
		));
	notech_and2 i_291(.A(n_1869), .B(n_1871), .Z(n_2555));
	notech_or2 i_496(.A(n_2497), .B(n_2333), .Z(n_2553));
	notech_and4 i_1101(.A(n_2510), .B(n_2500), .C(n_2547), .D(n_2498), .Z(n_2549
		));
	notech_and4 i_1095(.A(n_2534), .B(n_2522), .C(n_2526), .D(n_2545), .Z(n_2547
		));
	notech_and4 i_1088(.A(n_2538), .B(n_2111), .C(n_3982), .D(n_2543), .Z(n_2545
		));
	notech_and2 i_433(.A(n_3880), .B(n_29931), .Z(n_2543));
	notech_nor2 i_832(.A(n_2486), .B(n_2288), .Z(n_2542));
	notech_ao3 i_829(.A(modrm[2]), .B(n_2287), .C(n_2333), .Z(n_2541));
	notech_and3 i_608(.A(n_1798), .B(n_1796), .C(n_2111), .Z(n_2539));
	notech_and2 i_190(.A(n_1798), .B(n_1796), .Z(n_2538));
	notech_and4 i_84(.A(n_57916), .B(n_2431), .C(n_30108), .D(n_30117), .Z(n_2536
		));
	notech_and4 i_362(.A(n_2206), .B(n_4028), .C(n_2532), .D(n_3777), .Z(n_2534
		));
	notech_and4 i_638(.A(n_2206), .B(n_4028), .C(n_3992), .D(n_2123), .Z(n_2533
		));
	notech_and2 i_423(.A(n_3992), .B(n_2123), .Z(n_2532));
	notech_nand2 i_963(.A(n_30107), .B(n_29925), .Z(n_2531));
	notech_and4 i_83(.A(n_2431), .B(n_57916), .C(n_30108), .D(modrm[5]), .Z(n_2530
		));
	notech_and4 i_315(.A(n_3665), .B(n_2216), .C(n_3672), .D(n_2212), .Z(n_2526
		));
	notech_nand3 i_833(.A(n_2310), .B(n_29926), .C(n_57854), .Z(n_2523));
	notech_and4 i_298(.A(n_4004), .B(n_2398), .C(n_2513), .D(n_2518), .Z(n_2522
		));
	notech_or4 i_187(.A(n_57885), .B(n_2244), .C(n_57872), .D(n_30111), .Z(n_2519
		));
	notech_and2 i_713(.A(n_2516), .B(n_1890), .Z(n_2518));
	notech_or4 i_495(.A(n_57885), .B(n_2289), .C(n_57872), .D(n_30111), .Z(n_2517
		));
	notech_and2 i_903(.A(n_2515), .B(n_2032), .Z(n_2516));
	notech_or4 i_580(.A(n_2279), .B(n_57811), .C(n_30110), .D(n_57905), .Z(n_2515
		));
	notech_and2 i_703(.A(n_2234), .B(n_4005), .Z(n_2513));
	notech_and2 i_392(.A(n_2289), .B(n_30045), .Z(n_2512));
	notech_and4 i_380(.A(n_1901), .B(n_4087), .C(n_2198), .D(n_3972), .Z(n_2510
		));
	notech_or4 i_991(.A(n_2410), .B(modrm[3]), .C(modrm[4]), .D(modrm[5]), .Z
		(n_2505));
	notech_xor2 i_432(.A(n_30118), .B(modrm[7]), .Z(n_2504));
	notech_or4 i_90(.A(n_2410), .B(modrm[3]), .C(n_30116), .D(n_30117), .Z(n_2501
		));
	notech_and2 i_213(.A(n_3834), .B(n_3984), .Z(n_2500));
	notech_or4 i_87(.A(n_2386), .B(n_2315), .C(n_30110), .D(n_30117), .Z(n_2499
		));
	notech_and2 i_771(.A(n_1993), .B(n_1915), .Z(n_2498));
	notech_or4 i_48(.A(n_2329), .B(n_2292), .C(n_57925), .D(n_57905), .Z(n_2497
		));
	notech_and2 i_418(.A(n_2373), .B(n_2372), .Z(n_2495));
	notech_or4 i_578(.A(n_2486), .B(n_2485), .C(modrm[1]), .D(n_30113), .Z(n_2494
		));
	notech_and2 i_403(.A(n_30115), .B(n_30116), .Z(n_2492));
	notech_or4 i_885(.A(n_57872), .B(n_30072), .C(n_30117), .D(modrm[1]), .Z
		(n_2490));
	notech_or2 i_106(.A(n_2488), .B(modrm[0]), .Z(n_2489));
	notech_or4 i_836(.A(n_2325), .B(n_2485), .C(n_30117), .D(n_30114), .Z(n_2488
		));
	notech_or4 i_40(.A(n_57885), .B(n_57854), .C(n_57872), .D(n_30117), .Z(n_2486
		));
	notech_or4 i_49(.A(n_2329), .B(n_2300), .C(n_57925), .D(n_57905), .Z(n_2485
		));
	notech_and4 i_799(.A(n_1919), .B(n_3998), .C(n_29986), .D(n_29990), .Z(n_2484
		));
	notech_and4 i_319(.A(n_3967), .B(n_2480), .C(n_2479), .D(n_2415), .Z(n_2483
		));
	notech_ao4 i_129(.A(n_2027), .B(n_2393), .C(n_2346), .D(n_2387), .Z(n_2480
		));
	notech_and2 i_611(.A(n_3876), .B(n_4022), .Z(n_2479));
	notech_nand3 i_803(.A(n_2450), .B(n_2036), .C(n_2474), .Z(n_2475));
	notech_and3 i_795(.A(n_247289127), .B(n_2465), .C(n_1848), .Z(n_2474));
	notech_and3 i_800(.A(n_4025), .B(n_29975), .C(n_29973), .Z(n_247289127)
		);
	notech_and2 i_831(.A(cpl[1]), .B(cpl[0]), .Z(n_2469));
	notech_ao3 i_408(.A(n_57885), .B(n_2272), .C(n_2383), .Z(n_2466));
	notech_and4 i_504(.A(n_3965), .B(n_29992), .C(n_29957), .D(n_29991), .Z(n_2465
		));
	notech_or4 i_530(.A(n_57811), .B(n_30004), .C(n_57845), .D(n_30107), .Z(n_2464
		));
	notech_and4 i_119(.A(n_2189), .B(n_2206), .C(n_2179), .D(n_2457), .Z(n_2463
		));
	notech_or4 i_528(.A(n_57885), .B(n_57854), .C(n_57872), .D(n_29995), .Z(n_2458
		));
	notech_and3 i_316(.A(n_2255), .B(n_1805), .C(n_3975), .Z(n_2457));
	notech_or4 i_99(.A(n_57811), .B(n_57872), .C(n_30072), .D(n_57845), .Z(n_2455
		));
	notech_ao3 i_470(.A(n_3970), .B(n_1806), .C(n_1807), .Z(n_2450));
	notech_nand3 i_150(.A(n_2310), .B(n_57854), .C(n_29919), .Z(n_2448));
	notech_or4 i_849(.A(n_57810), .B(n_2311), .C(n_57845), .D(n_57753), .Z(n_2447
		));
	notech_nao3 i_457(.A(n_57925), .B(n_57905), .C(n_2311), .Z(n_2446));
	notech_or4 i_801(.A(n_29966), .B(n_30049), .C(n_2442), .D(n_3986), .Z(n_2445
		));
	notech_nao3 i_784(.A(n_2440), .B(n_2430), .C(n_1846), .Z(n_2442));
	notech_and4 i_775(.A(n_1843), .B(n_2437), .C(n_2140), .D(n_29990), .Z(n_2440
		));
	notech_and4 i_761(.A(n_2435), .B(n_1960), .C(n_3993), .D(n_2305), .Z(n_2437
		));
	notech_and2 i_44972276(.A(n_2234), .B(n_2398), .Z(n_2435));
	notech_and2 i_69072258(.A(n_3993), .B(n_2305), .Z(n_2434));
	notech_or2 i_250(.A(n_2403), .B(n_2389), .Z(n_2433));
	notech_nor2 i_579(.A(n_57885), .B(n_2403), .Z(n_2431));
	notech_ao4 i_773(.A(n_30108), .B(n_1842), .C(n_2383), .D(n_2428), .Z(n_2430
		));
	notech_or4 i_527(.A(n_57916), .B(n_57794), .C(n_30110), .D(n_30072), .Z(n_2428
		));
	notech_and3 i_674(.A(n_30110), .B(n_2324), .C(n_2369), .Z(n_2427));
	notech_and4 i_636(.A(n_4062), .B(n_4093), .C(n_29961), .D(n_29972), .Z(n_2426
		));
	notech_or4 i_352(.A(n_2386), .B(n_2372), .C(n_57859), .D(n_30117), .Z(n_2422
		));
	notech_and4 i_127(.A(n_57885), .B(n_30111), .C(n_57859), .D(n_2354), .Z(n_2418
		));
	notech_and2 i_594(.A(n_1938), .B(n_1835), .Z(n_2417));
	notech_and3 i_450(.A(n_2137), .B(n_2045), .C(n_2411), .Z(n_2415));
	notech_and2 i_307(.A(n_2137), .B(n_2045), .Z(n_2414));
	notech_and2 i_398(.A(n_2302), .B(n_30067), .Z(n_2413));
	notech_or4 i_194(.A(n_57805), .B(n_2325), .C(n_57820), .D(n_30108), .Z(n_2412
		));
	notech_and3 i_142(.A(n_2231), .B(n_1833), .C(n_2026), .Z(n_2411));
	notech_nao3 i_730(.A(n_30108), .B(n_57820), .C(n_2276), .Z(n_2408));
	notech_or4 i_77(.A(n_57885), .B(n_2290), .C(n_57872), .D(n_30111), .Z(n_2407
		));
	notech_and4 i_246(.A(n_2395), .B(n_2402), .C(n_2392), .D(n_2379), .Z(n_2406
		));
	notech_ao4 i_725(.A(n_2401), .B(n_3958), .C(n_3963), .D(n_2396), .Z(n_2402
		));
	notech_or4 i_67(.A(n_2329), .B(n_57905), .C(n_57916), .D(n_29925), .Z(n_2401
		));
	notech_and2 i_390(.A(n_30057), .B(n_2399), .Z(n_2400));
	notech_or4 i_96(.A(n_2410), .B(n_30115), .C(n_30116), .D(modrm[5]), .Z(n_2399
		));
	notech_or4 i_691(.A(n_57881), .B(n_2299), .C(n_57854), .D(n_57868), .Z(n_2396
		));
	notech_and3 i_434(.A(n_1829), .B(n_1828), .C(n_1958), .Z(n_2395));
	notech_ao4 i_132(.A(n_2297), .B(n_2393), .C(n_2346), .D(n_2299), .Z(n_2394
		));
	notech_or4 i_107(.A(n_2347), .B(n_2313), .C(n_2282), .D(n_30111), .Z(n_2393
		));
	notech_ao4 i_778(.A(n_2391), .B(n_2387), .C(n_30053), .D(n_4090), .Z(n_2392
		));
	notech_and2 i_429(.A(n_29969), .B(n_30055), .Z(n_2391));
	notech_and4 i_100(.A(n_57881), .B(n_30111), .C(n_57868), .D(n_2354), .Z(n_2390
		));
	notech_nand3 i_664(.A(n_57881), .B(n_30111), .C(n_57868), .Z(n_2389));
	notech_and2 i_185(.A(n_2278), .B(n_2299), .Z(n_2387));
	notech_nand2 i_369(.A(n_57881), .B(n_57854), .Z(n_2386));
	notech_nand2 i_419(.A(n_2372), .B(n_2315), .Z(n_2385));
	notech_nao3 i_95(.A(modrm[6]), .B(modrm[7]), .C(n_2381), .Z(n_2384));
	notech_or4 i_85(.A(n_2329), .B(n_57916), .C(n_57794), .D(n_2271), .Z(n_2382
		));
	notech_or4 i_661(.A(n_57805), .B(n_2283), .C(n_57916), .D(n_57794), .Z(n_2381
		));
	notech_and4 i_325(.A(n_4031), .B(n_4056), .C(n_4084), .D(n_2377), .Z(n_2379
		));
	notech_and2 i_339(.A(n_4066), .B(n_29953), .Z(n_2377));
	notech_or4 i_344(.A(n_2286), .B(n_29925), .C(n_2346), .D(n_30117), .Z(n_2376
		));
	notech_nor2 i_705(.A(n_2346), .B(n_57717), .Z(n_2375));
	notech_xor2 i_389(.A(n_30116), .B(modrm[3]), .Z(n_2374));
	notech_nand2 i_46(.A(n_30115), .B(modrm[4]), .Z(n_2373));
	notech_nand2 i_183(.A(n_30115), .B(n_30116), .Z(n_2372));
	notech_or4 i_693(.A(n_2279), .B(n_57820), .C(n_30108), .D(n_57859), .Z(n_2371
		));
	notech_and2 i_168(.A(n_1817), .B(n_2364), .Z(n_2365));
	notech_and2 i_756(.A(n_3991), .B(n_1813), .Z(n_2364));
	notech_and2 i_459(.A(n_2275), .B(n_2302), .Z(n_2363));
	notech_or4 i_86(.A(n_2347), .B(n_2360), .C(n_2282), .D(n_30111), .Z(n_2362
		));
	notech_nand2 i_535(.A(n_57753), .B(n_57845), .Z(n_2360));
	notech_or4 i_71(.A(n_2329), .B(n_57925), .C(n_57905), .D(n_2271), .Z(n_2359
		));
	notech_or4 i_66(.A(n_2329), .B(n_57905), .C(n_57916), .D(n_2271), .Z(n_2355
		));
	notech_and4 i_64(.A(n_223489126), .B(n_1792), .C(n_29965), .D(n_1797), .Z
		(n_2352));
	notech_or4 i_577(.A(n_2348), .B(n_2284), .C(n_30045), .D(n_29925), .Z(n_2350
		));
	notech_nor2 i_111(.A(n_2348), .B(n_2284), .Z(n_2349));
	notech_nao3 i_13(.A(n_57859), .B(n_57850), .C(n_57881), .Z(n_2348));
	notech_or2 i_600(.A(n_57881), .B(n_57868), .Z(n_2347));
	notech_or4 i_79(.A(n_2282), .B(n_2280), .C(n_57845), .D(n_57753), .Z(n_2346
		));
	notech_and4 i_351(.A(n_2141), .B(n_4013), .C(n_2058), .D(n_2343), .Z(n_2344
		));
	notech_and4 i_683(.A(n_2340), .B(n_2233), .C(n_2195), .D(n_2099), .Z(n_2343
		));
	notech_and2 i_513(.A(n_4044), .B(n_29987), .Z(n_2340));
	notech_nao3 i_671(.A(n_57877), .B(n_2272), .C(n_2338), .Z(n_2339));
	notech_nao3 i_151(.A(n_30108), .B(n_57753), .C(n_2282), .Z(n_2338));
	notech_or4 i_585(.A(n_2316), .B(n_2276), .C(n_2037), .D(n_2333), .Z(n_2337
		));
	notech_or4 i_32(.A(n_57877), .B(n_57850), .C(n_57868), .D(modrm[5]), .Z(n_2333
		));
	notech_nao3 i_574(.A(modrm[7]), .B(modrm[6]), .C(n_2290), .Z(n_2331));
	notech_or4 i_121(.A(n_57800), .B(n_2283), .C(n_57925), .D(n_57794), .Z(n_2330
		));
	notech_nao3 i_1(.A(n_57845), .B(n_57820), .C(n_57800), .Z(n_2329));
	notech_or4 i_0(.A(twobyte), .B(fpu), .C(ipg_fault), .D(n_30112), .Z(n_2328
		));
	notech_nao3 i_3(.A(n_57780), .B(n_57859), .C(n_57877), .Z(n_2325));
	notech_nor2 i_449(.A(n_57881), .B(n_57850), .Z(n_2324));
	notech_nor2 i_599(.A(opz[0]), .B(opz[2]), .Z(n_2322));
	notech_and2 i_73(.A(opz[2]), .B(n_2319), .Z(n_2321));
	notech_nor2 i_597(.A(opz[0]), .B(opz[1]), .Z(n_2319));
	notech_or4 i_92(.A(n_2403), .B(n_2311), .C(n_57845), .D(n_57820), .Z(n_2318
		));
	notech_nand2 i_584(.A(n_30108), .B(n_57753), .Z(n_2316));
	notech_nand2 i_446(.A(n_57825), .B(n_57820), .Z(n_2313));
	notech_nand3 i_41(.A(n_57877), .B(n_57859), .C(n_57850), .Z(n_2311));
	notech_and2 i_382(.A(n_57881), .B(n_57859), .Z(n_2310));
	notech_and4 i_436(.A(n_2141), .B(n_4013), .C(n_2308), .D(n_2294), .Z(n_2309
		));
	notech_and3 i_657(.A(n_4037), .B(n_1820), .C(n_1824), .Z(n_2308));
	notech_ao4 i_405(.A(n_2290), .B(n_2300), .C(n_2289), .D(n_29925), .Z(n_2303
		));
	notech_ao3 i_91(.A(n_57916), .B(n_57794), .C(n_2300), .Z(n_2301));
	notech_nao3 i_282(.A(modrm[7]), .B(modrm[6]), .C(modrm[2]), .Z(n_2300)
		);
	notech_nand3 i_68(.A(n_57789), .B(n_57925), .C(n_2271), .Z(n_2299));
	notech_nand3 i_59(.A(n_57925), .B(n_57905), .C(n_2271), .Z(n_2297));
	notech_and2 i_5(.A(n_57921), .B(n_57905), .Z(n_2296));
	notech_nao3 i_468(.A(modrm[2]), .B(n_2271), .C(n_2286), .Z(n_2295));
	notech_and2 i_790(.A(n_2258), .B(n_1821), .Z(n_2294));
	notech_nao3 i_88(.A(n_57916), .B(n_57789), .C(n_2292), .Z(n_2293));
	notech_nand3 i_276(.A(modrm[7]), .B(modrm[2]), .C(modrm[6]), .Z(n_2292)
		);
	notech_and2 i_393(.A(n_2278), .B(n_29968), .Z(n_2291));
	notech_nand2 i_2(.A(n_57915), .B(n_57789), .Z(n_2290));
	notech_nand2 i_6(.A(n_57789), .B(n_57921), .Z(n_2289));
	notech_or4 i_590(.A(modrm[2]), .B(n_57921), .C(n_57789), .D(n_29925), .Z
		(n_2288));
	notech_and4 i_120(.A(modrm[7]), .B(n_57910), .C(n_57905), .D(modrm[6]), 
		.Z(n_2287));
	notech_nand2 i_772375(.A(n_57910), .B(n_57905), .Z(n_2286));
	notech_or4 i_75(.A(n_57735), .B(n_2280), .C(n_57825), .D(n_57753), .Z(n_2285
		));
	notech_nao3 i_856(.A(n_57841), .B(n_57820), .C(n_57735), .Z(n_2284));
	notech_nand2 i_589(.A(n_57841), .B(n_57820), .Z(n_2283));
	notech_or4 i_9(.A(fpu), .B(ipg_fault), .C(n_30112), .D(n_30120), .Z(n_2282
		));
	notech_nao3 i_44(.A(n_57850), .B(n_57868), .C(n_57881), .Z(n_2280));
	notech_or2 i_593(.A(n_57881), .B(n_57780), .Z(n_2279));
	notech_or4 i_857(.A(fpu), .B(ipg_fault), .C(op[7]), .D(n_30120), .Z(n_2276
		));
	notech_and2 i_537(.A(n_57780), .B(n_57859), .Z(n_2272));
	notech_and2 i_230(.A(modrm[7]), .B(modrm[6]), .Z(n_2271));
	notech_and4 i_281(.A(n_3591), .B(n_3560), .C(n_717), .D(n_1593), .Z(n_2270
		));
	notech_or2 i_2397(.A(n_2398), .B(n_57910), .Z(n_2269));
	notech_nand3 i_308(.A(n_2757), .B(n_3548), .C(n_1951), .Z(\udeco[8] ));
	notech_nand2 i_2345(.A(modrm[3]), .B(n_3174), .Z(n_2267));
	notech_nao3 i_2349(.A(opz[1]), .B(n_2322), .C(n_2247), .Z(n_2266));
	notech_or4 i_2341(.A(n_2410), .B(n_2373), .C(n_3954), .D(n_57717), .Z(n_2265
		));
	notech_or2 i_335(.A(n_2485), .B(n_2333), .Z(n_2264));
	notech_or4 i_2350(.A(n_57805), .B(n_2248), .C(n_57841), .D(n_57820), .Z(n_2263
		));
	notech_nand2 i_2353(.A(n_57899), .B(n_2251), .Z(n_2262));
	notech_or4 i_144(.A(n_2286), .B(modrm[2]), .C(n_2285), .D(n_57744), .Z(n_2258
		));
	notech_or4 i_2344(.A(n_2412), .B(n_57910), .C(n_57789), .D(n_2271), .Z(n_2257
		));
	notech_or4 i_2342(.A(n_57805), .B(n_2316), .C(n_2389), .D(n_2278), .Z(n_2256
		));
	notech_or4 i_23111193(.A(n_2313), .B(n_57910), .C(n_2271), .D(n_30065), 
		.Z(n_2255));
	notech_or4 i_2351(.A(n_57805), .B(n_57816), .C(n_57825), .D(n_2249), .Z(n_2254
		));
	notech_or4 i_2346(.A(n_2347), .B(n_2338), .C(n_2512), .D(n_57780), .Z(n_2253
		));
	notech_or4 i_822(.A(n_2280), .B(n_57805), .C(n_57899), .D(n_57841), .Z(n_2252
		));
	notech_nand2 i_202(.A(n_2433), .B(n_2678), .Z(n_2251));
	notech_and3 i_203(.A(n_2141), .B(n_4013), .C(n_2140), .Z(n_2250));
	notech_and2 i_205(.A(n_2448), .B(n_2243), .Z(n_2249));
	notech_ao4 i_209(.A(n_2486), .B(n_2288), .C(n_2348), .D(n_2289), .Z(n_2248
		));
	notech_ao4 i_219(.A(n_2318), .B(n_2297), .C(n_2401), .D(n_2101), .Z(n_2247
		));
	notech_ao3 i_222(.A(n_2275), .B(n_2302), .C(n_2301), .Z(n_2245));
	notech_and2 i_404(.A(n_57890), .B(n_30045), .Z(n_2244));
	notech_nao3 i_2339(.A(n_2310), .B(n_57850), .C(n_2244), .Z(n_2243));
	notech_and4 i_320(.A(n_2484), .B(n_2703), .C(n_3500), .D(n_3465), .Z(n_2241
		));
	notech_nand2 i_2293(.A(n_3174), .B(modrm[4]), .Z(n_2240));
	notech_or4 i_2294(.A(n_2410), .B(n_2373), .C(n_2230), .D(n_57717), .Z(n_2239
		));
	notech_or4 i_287(.A(n_2383), .B(n_2486), .C(n_2290), .D(n_2300), .Z(n_2238
		));
	notech_nand2 i_2291(.A(n_57868), .B(n_30032), .Z(n_2237));
	notech_or4 i_23111322(.A(n_2348), .B(n_2320), .C(n_2275), .D(n_2284), .Z
		(n_223489126));
	notech_or4 i_23111436(.A(n_57744), .B(n_2337), .C(n_57921), .D(n_57899),
		 .Z(n_2233));
	notech_or4 i_2290(.A(n_2285), .B(n_57910), .C(n_57789), .D(n_2271), .Z(n_2232
		));
	notech_or4 i_23111388(.A(n_2347), .B(n_2290), .C(n_2408), .D(n_57780), .Z
		(n_2231));
	notech_and2 i_200(.A(n_2382), .B(n_2485), .Z(n_2230));
	notech_or4 i_2286(.A(n_57890), .B(n_2329), .C(n_2325), .D(n_57762), .Z(n_2229
		));
	notech_or4 i_2285(.A(n_2285), .B(n_57899), .C(n_57910), .D(n_57744), .Z(n_2228
		));
	notech_and4 i_334(.A(n_2694), .B(n_3458), .C(n_3429), .D(n_2704), .Z(n_2227
		));
	notech_nand2 i_2248(.A(n_3174), .B(modrm[5]), .Z(n_2226));
	notech_nao3 i_2249(.A(n_29924), .B(n_30056), .C(n_2499), .Z(n_2223));
	notech_or2 i_2243(.A(n_2065), .B(n_57825), .Z(n_2222));
	notech_or4 i_2247(.A(n_2360), .B(n_57800), .C(n_57771), .D(n_2297), .Z(n_2221
		));
	notech_or4 i_2250(.A(n_2316), .B(n_2276), .C(n_2289), .D(n_2280), .Z(n_2220
		));
	notech_and4 i_345(.A(n_2904), .B(n_2703), .C(n_2484), .D(n_3425), .Z(n_221989125
		));
	notech_or4 i_149(.A(n_2244), .B(n_2185), .C(n_57859), .D(n_2386), .Z(n_2218
		));
	notech_or2 i_2216(.A(n_2065), .B(n_57789), .Z(n_2217));
	notech_or4 i_23110650(.A(n_2329), .B(n_57899), .C(n_57910), .D(n_2389), 
		.Z(n_2216));
	notech_and4 i_431(.A(n_2689), .B(n_2501), .C(n_2499), .D(n_2422), .Z(n_2215
		));
	notech_or2 i_2215(.A(n_2215), .B(n_2359), .Z(n_2213));
	notech_and4 i_363(.A(n_2484), .B(n_3397), .C(n_2904), .D(n_2704), .Z(n_2208
		));
	notech_or2 i_2183(.A(n_2215), .B(n_2497), .Z(n_2207));
	notech_or4 i_23111190(.A(n_2316), .B(n_57910), .C(n_30065), .D(n_57762),
		 .Z(n_2206));
	notech_and2 i_353(.A(n_2295), .B(n_2293), .Z(n_2205));
	notech_or4 i_361(.A(n_57890), .B(n_2292), .C(n_2329), .D(n_30053), .Z(n_2202
		));
	notech_nand3 i_385(.A(n_3364), .B(n_3343), .C(n_1951), .Z(\udeco[16] )
		);
	notech_nao3 i_2126(.A(opz[1]), .B(n_2322), .C(n_2187), .Z(n_2200));
	notech_or2 i_2123(.A(n_2883), .B(n_30115), .Z(n_2199));
	notech_or2 i_297(.A(n_4090), .B(n_30053), .Z(n_2198));
	notech_or4 i_2125(.A(n_2373), .B(n_57717), .C(n_2410), .D(n_2115), .Z(n_2197
		));
	notech_or4 i_2120(.A(n_57694), .B(n_2037), .C(n_3954), .D(n_57717), .Z(n_2196
		));
	notech_or4 i_153(.A(n_57881), .B(n_2330), .C(n_57854), .D(n_57868), .Z(n_2195
		));
	notech_or4 i_2119(.A(n_2292), .B(n_2285), .C(n_57921), .D(n_57899), .Z(n_2193
		));
	notech_or4 i_677(.A(n_30004), .B(n_57899), .C(n_57910), .D(n_30051), .Z(n_2192
		));
	notech_or2 i_2982(.A(n_2300), .B(n_30043), .Z(n_2190));
	notech_or4 i_1241(.A(n_57910), .B(n_30065), .C(n_57841), .D(n_57744), .Z
		(n_2189));
	notech_or4 i_179(.A(n_57881), .B(n_2403), .C(n_2360), .D(n_57921), .Z(n_2188
		));
	notech_ao4 i_181(.A(n_4065), .B(n_2297), .C(n_2098), .D(n_2101), .Z(n_2187
		));
	notech_and2 i_524(.A(n_2668), .B(n_3154), .Z(n_2186));
	notech_and3 i_394(.A(n_2383), .B(n_30051), .C(n_29995), .Z(n_2185));
	notech_or4 i_2116(.A(n_2285), .B(n_57921), .C(n_57899), .D(n_57762), .Z(n_2183
		));
	notech_nao3 i_2115(.A(opz[1]), .B(n_2322), .C(n_2350), .Z(n_2181));
	notech_nand3 i_2110(.A(n_3895), .B(n_57854), .C(n_2310), .Z(n_2180));
	notech_or4 i_39(.A(n_2458), .B(n_57915), .C(n_57789), .D(n_57762), .Z(n_2179
		));
	notech_and4 i_400(.A(n_3309), .B(n_3302), .C(n_3273), .D(n_2562), .Z(n_2177
		));
	notech_or2 i_2061(.A(n_2883), .B(n_30116), .Z(n_2175));
	notech_or4 i_2060(.A(n_57694), .B(n_2373), .C(n_3836), .D(n_57717), .Z(n_2174
		));
	notech_nand2 i_2064(.A(n_57868), .B(n_30078), .Z(n_2173));
	notech_nao3 i_2062(.A(n_2321), .B(n_30059), .C(n_2101), .Z(n_2172));
	notech_or4 i_2063(.A(n_2403), .B(n_2161), .C(n_2313), .D(n_2311), .Z(n_2170
		));
	notech_or4 i_2058(.A(n_57694), .B(n_2037), .C(n_57717), .D(n_2355), .Z(n_2169
		));
	notech_nao3 i_2056(.A(n_2385), .B(n_29922), .C(n_2214), .Z(n_2168));
	notech_or4 i_227(.A(n_57771), .B(n_57762), .C(n_30045), .D(n_30051), .Z(n_2166
		));
	notech_or4 i_2059(.A(n_57921), .B(n_57899), .C(n_57762), .D(n_29969), .Z
		(n_2163));
	notech_ao4 i_518(.A(n_2297), .B(n_30073), .C(n_2275), .D(n_2149), .Z(n_2161
		));
	notech_or4 i_224(.A(n_57890), .B(n_2486), .C(n_57762), .D(n_29995), .Z(n_2159
		));
	notech_or4 i_2050(.A(n_57800), .B(n_2594), .C(n_57841), .D(n_57816), .Z(n_2155
		));
	notech_and2 i_290(.A(n_2285), .B(n_29969), .Z(n_2154));
	notech_and2 i_328(.A(n_2320), .B(n_30073), .Z(n_2149));
	notech_and4 i_414(.A(n_2757), .B(n_3257), .C(n_1504), .D(n_520), .Z(n_2146
		));
	notech_or2 i_2004(.A(n_2883), .B(n_57717), .Z(n_2145));
	notech_or4 i_2002(.A(n_57694), .B(n_2037), .C(n_3836), .D(n_57717), .Z(n_2144
		));
	notech_nand2 i_2005(.A(n_57854), .B(n_30078), .Z(n_2143));
	notech_and3 i_2003(.A(n_2287), .B(n_2375), .C(n_2385), .Z(n_2142));
	notech_nao3 i_1250(.A(n_2397), .B(n_57762), .C(n_2276), .Z(n_2141));
	notech_or4 i_180(.A(n_57881), .B(n_2403), .C(n_2283), .D(n_57850), .Z(n_2140
		));
	notech_and3 i_326(.A(n_2485), .B(n_2401), .C(n_2497), .Z(n_2139));
	notech_or4 i_675(.A(n_57703), .B(n_57800), .C(n_57771), .D(n_2027), .Z(n_2137
		));
	notech_or2 i_591(.A(n_2497), .B(n_30053), .Z(n_2136));
	notech_and4 i_438(.A(n_530), .B(n_2703), .C(n_3213), .D(n_537), .Z(n_2135
		));
	notech_or4 i_1968(.A(n_57694), .B(n_2373), .C(n_3954), .D(modrm[5]), .Z(n_2134
		));
	notech_or4 i_1967(.A(n_57921), .B(n_57899), .C(n_57762), .D(n_30066), .Z
		(n_2132));
	notech_nao3 i_1935(.A(n_30115), .B(n_30116), .C(n_2376), .Z(n_2131));
	notech_or4 i_1934(.A(n_57694), .B(n_2373), .C(n_2384), .D(n_57717), .Z(n_2130
		));
	notech_or4 i_1933(.A(n_57703), .B(n_57800), .C(n_57771), .D(n_2302), .Z(n_2129
		));
	notech_ao3 i_1931(.A(n_2299), .B(n_2297), .C(n_2301), .Z(n_2128));
	notech_and4 i_48310341(.A(n_719), .B(n_3171), .C(n_3143), .D(n_1950), .Z
		(n_2127));
	notech_nand3 i_1902(.A(opz[1]), .B(n_2322), .C(n_2117), .Z(n_2126));
	notech_or2 i_1898(.A(n_3728), .B(n_30115), .Z(n_2125));
	notech_or4 i_1901(.A(n_57694), .B(n_2037), .C(n_2115), .D(n_57717), .Z(n_2122
		));
	notech_or2 i_1899(.A(n_3697), .B(n_57789), .Z(n_2121));
	notech_or2 i_1897(.A(n_2151), .B(n_57915), .Z(n_2120));
	notech_or2 i_1900(.A(n_2052), .B(n_29968), .Z(n_2119));
	notech_nand2 i_169(.A(n_2988), .B(n_2350), .Z(n_2117));
	notech_and3 i_174(.A(n_2497), .B(n_2359), .C(n_2355), .Z(n_2115));
	notech_nand3 i_124(.A(n_57744), .B(n_57816), .C(n_2536), .Z(n_2111));
	notech_nao3 i_472(.A(n_1718), .B(n_3141), .C(n_4024), .Z(\udeco[25] ));
	notech_nand2 i_1860(.A(modrm[4]), .B(n_29981), .Z(n_2109));
	notech_or4 i_838(.A(n_57881), .B(n_57850), .C(n_57868), .D(n_2098), .Z(n_2108
		));
	notech_nand2 i_1861(.A(n_57868), .B(n_29982), .Z(n_2107));
	notech_nao3 i_1197(.A(opz[2]), .B(n_2319), .C(n_2350), .Z(n_2106));
	notech_or2 i_1858(.A(n_2151), .B(n_57753), .Z(n_2105));
	notech_nao3 i_827(.A(n_2287), .B(n_2375), .C(n_2374), .Z(n_2104));
	notech_or4 i_47(.A(n_2596), .B(n_57921), .C(n_57789), .D(n_57762), .Z(n_2103
		));
	notech_ao3 i_16372320(.A(opz[2]), .B(n_2319), .C(n_2083), .Z(n_2102));
	notech_and2 i_633(.A(n_2499), .B(n_2422), .Z(n_2101));
	notech_ao3 i_1824(.A(n_29924), .B(n_29928), .C(n_2499), .Z(n_2100));
	notech_and2 i_329(.A(n_2401), .B(n_2355), .Z(n_2098));
	notech_or4 i_1823(.A(n_57694), .B(n_2315), .C(n_3836), .D(n_57717), .Z(n_2097
		));
	notech_and4 i_1811(.A(n_2278), .B(n_2275), .C(n_29968), .D(n_2293), .Z(n_2095
		));
	notech_and4 i_546(.A(n_3091), .B(n_2903), .C(n_30104), .D(n_30064), .Z(n_2092
		));
	notech_or2 i_416(.A(n_3957), .B(n_2098), .Z(n_2091));
	notech_nao3 i_1775(.A(opz[1]), .B(n_2322), .C(n_2083), .Z(n_2090));
	notech_or4 i_1776(.A(n_2348), .B(n_57703), .C(n_57735), .D(n_2291), .Z(n_2089
		));
	notech_or4 i_1778(.A(n_2311), .B(n_3963), .C(n_57921), .D(n_57899), .Z(n_2087
		));
	notech_or4 i_1777(.A(n_57703), .B(n_2280), .C(n_57735), .D(n_30067), .Z(n_2086
		));
	notech_ao4 i_516(.A(n_2101), .B(n_2355), .C(n_4065), .D(n_2027), .Z(n_2083
		));
	notech_nand3 i_745(.A(n_3054), .B(n_2079), .C(n_30122), .Z(\udeco[108] )
		);
	notech_nand2 i_1646(.A(opz[0]), .B(n_2067), .Z(n_2079));
	notech_nor2 i_192(.A(n_2400), .B(n_3845), .Z(n_2078));
	notech_ao4 i_1647(.A(n_2418), .B(n_30069), .C(n_2301), .D(n_3908), .Z(n_2077
		));
	notech_or2 i_1648(.A(n_2359), .B(n_2069), .Z(n_2075));
	notech_or2 i_1645(.A(n_2523), .B(n_3961), .Z(n_2074));
	notech_or4 i_55(.A(modrm[2]), .B(n_2330), .C(n_57744), .D(n_30053), .Z(n_2073
		));
	notech_or4 i_1649(.A(n_2347), .B(n_57890), .C(n_3963), .D(n_57780), .Z(n_2072
		));
	notech_or4 i_23110740(.A(n_30004), .B(n_2329), .C(n_2331), .D(modrm[5]),
		 .Z(n_2071));
	notech_or4 i_23110743(.A(n_2586), .B(n_57925), .C(n_57899), .D(n_57744),
		 .Z(n_2070));
	notech_and3 i_163(.A(n_2400), .B(n_30004), .C(n_30053), .Z(n_2069));
	notech_nand3 i_165(.A(n_3018), .B(n_3013), .C(n_2955), .Z(n_2067));
	notech_or4 i_1629(.A(n_57800), .B(n_2574), .C(n_57841), .D(n_57753), .Z(n_2063
		));
	notech_nand2 i_1627(.A(n_2407), .B(n_2061), .Z(n_2062));
	notech_or4 i_254(.A(n_57881), .B(n_57890), .C(n_57868), .D(n_57780), .Z(n_2061
		));
	notech_and2 i_294(.A(n_2383), .B(n_2329), .Z(n_2059));
	notech_nao3 i_1622(.A(n_29926), .B(n_30121), .C(n_2407), .Z(n_2057));
	notech_or4 i_1620(.A(n_57800), .B(n_2407), .C(n_57841), .D(n_57816), .Z(n_2056
		));
	notech_and4 i_762(.A(n_3005), .B(n_2987), .C(n_2054), .D(n_30122), .Z(n_2055
		));
	notech_nand2 i_1590(.A(opz[1]), .B(n_30083), .Z(n_2054));
	notech_nao3 i_1586(.A(opz[1]), .B(n_2322), .C(n_2988), .Z(n_2053));
	notech_or2 i_1584(.A(adz), .B(n_2036), .Z(n_2051));
	notech_nao3 i_1585(.A(n_30113), .B(n_2037), .C(n_2488), .Z(n_2050));
	notech_or4 i_1228(.A(n_2485), .B(n_2490), .C(n_2492), .D(modrm[0]), .Z(n_2046
		));
	notech_or4 i_854(.A(n_57703), .B(n_57800), .C(n_57771), .D(n_2413), .Z(n_2045
		));
	notech_or4 i_1589(.A(n_57800), .B(n_2313), .C(n_2486), .D(n_2288), .Z(n_2042
		));
	notech_or4 i_1592(.A(n_57771), .B(n_3963), .C(n_57717), .D(n_2295), .Z(n_2041
		));
	notech_or4 i_1587(.A(n_57805), .B(n_2428), .C(n_57825), .D(n_57753), .Z(n_2040
		));
	notech_and4 i_158(.A(n_2309), .B(n_2958), .C(n_2975), .D(n_2955), .Z(n_2038
		));
	notech_nand2 i_564(.A(modrm[3]), .B(modrm[4]), .Z(n_2037));
	notech_and3 i_197(.A(n_2327), .B(n_4047), .C(n_3981), .Z(n_2036));
	notech_nand3 i_1566(.A(n_57881), .B(n_2272), .C(n_29928), .Z(n_2034));
	notech_or2 i_1567(.A(n_2523), .B(n_2512), .Z(n_2033));
	notech_or4 i_826(.A(n_2279), .B(n_57805), .C(n_57859), .D(n_57789), .Z(n_2032
		));
	notech_or4 i_1562(.A(n_2347), .B(n_2512), .C(n_57780), .D(n_2059), .Z(n_2031
		));
	notech_or4 i_1282(.A(n_2348), .B(n_57735), .C(n_1888), .D(n_57703), .Z(n_2030
		));
	notech_or4 i_1553(.A(n_3963), .B(n_2027), .C(n_57868), .D(n_30072), .Z(n_2028
		));
	notech_and2 i_301(.A(n_2275), .B(n_2297), .Z(n_2027));
	notech_or4 i_845(.A(n_2313), .B(n_57735), .C(n_2348), .D(n_2387), .Z(n_2026
		));
	notech_or4 i_1543(.A(n_2214), .B(n_2497), .C(modrm[3]), .D(n_30116), .Z(n_2025
		));
	notech_or4 i_1541(.A(n_2280), .B(n_57805), .C(n_57904), .D(n_57825), .Z(n_2021
		));
	notech_and4 i_796(.A(n_2939), .B(n_2936), .C(n_1718), .D(n_2890), .Z(n_2020
		));
	notech_or2 i_1174(.A(n_2400), .B(n_2401), .Z(n_2019));
	notech_or4 i_834(.A(n_57890), .B(n_57859), .C(n_30072), .D(n_29995), .Z(n_2014
		));
	notech_ao4 i_178(.A(n_2542), .B(n_2541), .C(n_2369), .D(n_2354), .Z(n_2013
		));
	notech_nand3 i_873(.A(n_2881), .B(n_1593), .C(n_2011), .Z(\udeco[117] )
		);
	notech_nand2 i_1366(.A(n_30034), .B(n_30085), .Z(n_2011));
	notech_nand2 i_1367(.A(modrm[4]), .B(n_3773), .Z(n_2010));
	notech_nand2 i_1368(.A(modrm[1]), .B(n_2007), .Z(n_2009));
	notech_or4 i_1365(.A(n_57735), .B(n_30004), .C(n_57794), .D(n_57753), .Z
		(n_2008));
	notech_nand3 i_140(.A(n_2099), .B(n_3736), .C(n_2654), .Z(n_2007));
	notech_mux2 i_396(.S(n_57816), .A(n_30116), .B(n_30114), .Z(n_2006));
	notech_or4 i_1361(.A(n_57703), .B(n_57805), .C(n_2519), .D(n_30121), .Z(n_2005
		));
	notech_or4 i_90810263(.A(n_2002), .B(n_2001), .C(n_2820), .D(n_1180), .Z
		(\udeco[120] ));
	notech_and2 i_1287(.A(n_3763), .B(n_1968), .Z(n_2002));
	notech_and2 i_1281(.A(n_29971), .B(n_29970), .Z(n_2001));
	notech_and2 i_1285(.A(modrm[0]), .B(n_30086), .Z(n_2000));
	notech_and2 i_1286(.A(modrm[3]), .B(n_1988), .Z(n_1998));
	notech_nor2 i_1288(.A(n_2362), .B(n_1989), .Z(n_1997));
	notech_or4 i_1141(.A(n_57703), .B(n_2280), .C(n_57735), .D(n_2413), .Z(n_1995
		));
	notech_or4 i_1280(.A(n_57810), .B(n_2517), .C(n_57845), .D(n_57816), .Z(n_1994
		));
	notech_or4 i_1284(.A(n_2347), .B(n_2338), .C(n_2244), .D(n_57780), .Z(n_1990
		));
	notech_and4 i_116(.A(n_2275), .B(n_2297), .C(n_2278), .D(n_2299), .Z(n_1989
		));
	notech_nand3 i_118(.A(n_2480), .B(n_1777), .C(n_2415), .Z(n_1988));
	notech_and4 i_655(.A(n_2309), .B(n_2760), .C(n_2717), .D(n_2759), .Z(n_1986
		));
	notech_or4 i_1275(.A(n_2315), .B(n_2214), .C(n_2330), .D(n_57744), .Z(n_1985
		));
	notech_or2 i_1273(.A(n_2382), .B(n_30053), .Z(n_1982));
	notech_or4 i_1272(.A(n_2372), .B(n_2214), .C(n_2330), .D(n_57744), .Z(n_1981
		));
	notech_or4 i_908(.A(n_1979), .B(n_1321), .C(n_1977), .D(n_2785), .Z(\udeco[121] 
		));
	notech_and2 i_1239(.A(n_1968), .B(n_30087), .Z(n_1979));
	notech_and2 i_1231(.A(n_29970), .B(n_30085), .Z(n_1977));
	notech_and2 i_1237(.A(modrm[1]), .B(n_30086), .Z(n_1976));
	notech_and2 i_1238(.A(modrm[4]), .B(n_1964), .Z(n_1975));
	notech_nand3 i_114(.A(n_2688), .B(n_2757), .C(n_2166), .Z(n_1968));
	notech_mux2 i_422(.S(n_57816), .A(n_30114), .B(n_30116), .Z(n_1965));
	notech_nand3 i_115(.A(n_2395), .B(n_1777), .C(n_2415), .Z(n_1964));
	notech_or4 i_483(.A(n_1326), .B(n_222991118), .C(n_1956), .D(n_30026), .Z
		(\udeco[122] ));
	notech_and2 i_1192(.A(modrm[2]), .B(n_1946), .Z(n_1956));
	notech_nand2 i_1191(.A(modrm[5]), .B(n_1945), .Z(n_1955));
	notech_nand2 i_1189(.A(n_1944), .B(n_30061), .Z(n_1954));
	notech_or4 i_1190(.A(n_2387), .B(n_57868), .C(n_30072), .D(n_29995), .Z(n_1952
		));
	notech_or4 i_1187(.A(n_57810), .B(n_57771), .C(n_57845), .D(n_3761), .Z(n_1949
		));
	notech_or2 i_1186(.A(n_2734), .B(n_57825), .Z(n_1947));
	notech_nand3 i_104(.A(n_2719), .B(n_2717), .C(n_2091), .Z(n_1946));
	notech_nand3 i_112(.A(n_2723), .B(n_4017), .C(n_2726), .Z(n_1945));
	notech_mux2 i_506(.S(n_57816), .A(n_57726), .B(modrm[2]), .Z(n_1944));
	notech_mux2 i_505(.S(n_57816), .A(modrm[2]), .B(n_57726), .Z(n_1943));
	notech_or2 i_1180(.A(n_1940), .B(n_2285), .Z(n_1941));
	notech_and4 i_113(.A(n_2027), .B(n_2387), .C(n_2302), .D(n_29968), .Z(n_1940
		));
	notech_or4 i_23111442(.A(n_57744), .B(n_2052), .C(n_57921), .D(n_57904),
		 .Z(n_1938));
	notech_and2 i_313(.A(n_2422), .B(n_2325), .Z(n_1937));
	notech_or4 i_1170(.A(n_2393), .B(n_57904), .C(n_57915), .D(n_29925), .Z(n_1936
		));
	notech_and4 i_1157(.A(n_57868), .B(n_2324), .C(n_2296), .D(n_29926), .Z(n_1933
		));
	notech_or2 i_1156(.A(n_2101), .B(n_2382), .Z(n_1932));
	notech_or2 i_1123(.A(n_3845), .B(n_30053), .Z(n_1930));
	notech_or4 i_1116(.A(n_57703), .B(n_57805), .C(n_30004), .D(n_2289), .Z(n_1921
		));
	notech_or4 i_1057(.A(n_2214), .B(n_2382), .C(n_30115), .D(n_30116), .Z(n_1919
		));
	notech_or4 i_1044(.A(n_2348), .B(n_30045), .C(adz), .D(n_2059), .Z(n_1918
		));
	notech_or4 i_284(.A(n_57805), .B(n_2286), .C(n_57816), .D(n_57825), .Z(n_1917
		));
	notech_and2 i_1042(.A(n_2330), .B(n_1917), .Z(n_1916));
	notech_or2 i_1030(.A(n_3836), .B(n_30053), .Z(n_1915));
	notech_or2 i_1028(.A(n_2494), .B(n_1913), .Z(n_1914));
	notech_and3 i_311(.A(n_2373), .B(n_2372), .C(n_2037), .Z(n_1913));
	notech_nao3 i_1027(.A(n_30113), .B(n_2385), .C(n_2488), .Z(n_1912));
	notech_or2 i_1018(.A(n_2497), .B(n_2486), .Z(n_1911));
	notech_or4 i_1011(.A(n_57816), .B(n_57825), .C(n_57915), .D(n_30065), .Z
		(n_1907));
	notech_ao4 i_1003(.A(n_2037), .B(n_2486), .C(n_57859), .D(n_2279), .Z(n_1902
		));
	notech_or4 i_992(.A(n_2330), .B(modrm[6]), .C(modrm[7]), .D(n_2505), .Z(n_1901
		));
	notech_and2 i_989(.A(modrm[6]), .B(modrm[7]), .Z(n_1900));
	notech_or4 i_975(.A(n_2412), .B(n_57904), .C(n_57915), .D(n_57762), .Z(n_1896
		));
	notech_or4 i_968(.A(n_2458), .B(n_57904), .C(n_57915), .D(n_57762), .Z(n_1895
		));
	notech_or4 i_956(.A(n_2313), .B(n_57735), .C(n_2280), .D(n_2387), .Z(n_1892
		));
	notech_or2 i_946(.A(n_3935), .B(n_3963), .Z(n_1890));
	notech_and4 i_940(.A(n_2027), .B(n_2387), .C(n_29968), .D(n_2413), .Z(n_1888
		));
	notech_or4 i_938(.A(modrm[1]), .B(n_2553), .C(n_30113), .D(n_2495), .Z(n_1887
		));
	notech_or4 i_937(.A(modrm[1]), .B(n_2553), .C(modrm[0]), .D(n_2492), .Z(n_1886
		));
	notech_mux2 i_321(.S(modrm[0]), .A(n_1882), .B(n_2037), .Z(n_1885));
	notech_nand3 i_322(.A(n_2372), .B(n_2315), .C(n_2037), .Z(n_1882));
	notech_nand2 i_932(.A(n_2037), .B(modrm[0]), .Z(n_1879));
	notech_or4 i_922(.A(n_2300), .B(n_2455), .C(n_57921), .D(n_57904), .Z(n_1877
		));
	notech_or4 i_913(.A(n_2360), .B(n_57805), .C(n_30004), .D(n_57890), .Z(n_1875
		));
	notech_or4 i_898(.A(modrm[1]), .B(n_2553), .C(modrm[0]), .D(n_2372), .Z(n_1874
		));
	notech_or4 i_897(.A(modrm[1]), .B(n_2553), .C(n_2315), .D(n_30113), .Z(n_1873
		));
	notech_mux2 i_312(.S(modrm[0]), .A(n_2373), .B(n_2037), .Z(n_1872));
	notech_or4 i_894(.A(n_2497), .B(n_2333), .C(n_1872), .D(n_30114), .Z(n_1871
		));
	notech_or4 i_893(.A(n_2485), .B(n_2372), .C(n_2490), .D(modrm[0]), .Z(n_1869
		));
	notech_ao4 i_881(.A(n_2333), .B(n_2288), .C(n_2486), .D(n_2295), .Z(n_1858
		));
	notech_or4 i_875(.A(n_2383), .B(n_2333), .C(n_2290), .D(n_2300), .Z(n_1857
		));
	notech_nao3 i_870(.A(n_57753), .B(n_2530), .C(n_2300), .Z(n_1855));
	notech_nao3 i_869(.A(n_57816), .B(n_2536), .C(n_2292), .Z(n_1854));
	notech_or4 i_825(.A(n_57771), .B(n_2302), .C(n_3963), .D(n_57726), .Z(n_1851
		));
	notech_or4 i_954(.A(n_2475), .B(n_2445), .C(n_1849), .D(n_1838), .Z(\udeco[126] 
		));
	notech_and2 i_752(.A(modrm[2]), .B(n_30092), .Z(n_1849));
	notech_nand2 i_741(.A(n_1943), .B(n_30061), .Z(n_1848));
	notech_and4 i_743(.A(n_57744), .B(n_1944), .C(n_2296), .D(n_2427), .Z(n_1846
		));
	notech_or2 i_740(.A(n_2433), .B(n_57904), .Z(n_1843));
	notech_and2 i_69(.A(n_2032), .B(n_3733), .Z(n_1842));
	notech_and4 i_81(.A(n_1837), .B(n_2417), .C(n_2415), .D(n_2406), .Z(n_1841
		));
	notech_and4 i_82(.A(n_2352), .B(n_2344), .C(n_1905), .D(n_1825), .Z(n_1840
		));
	notech_and2 i_749(.A(n_57726), .B(n_30093), .Z(n_1838));
	notech_or4 i_735(.A(n_57805), .B(n_2316), .C(n_30004), .D(n_2387), .Z(n_1837
		));
	notech_nand3 i_734(.A(n_57881), .B(n_2272), .C(n_30056), .Z(n_1835));
	notech_or4 i_731(.A(n_2276), .B(n_2407), .C(n_57845), .D(n_57816), .Z(n_1833
		));
	notech_or4 i_673(.A(n_2299), .B(n_3963), .C(n_57868), .D(n_30072), .Z(n_1831
		));
	notech_or4 i_718(.A(n_2393), .B(n_57915), .C(n_57789), .D(n_57744), .Z(n_1829
		));
	notech_or4 i_717(.A(n_2313), .B(n_57735), .C(n_2280), .D(n_2299), .Z(n_1828
		));
	notech_nao3 i_851(.A(n_57881), .B(n_2272), .C(n_4072), .Z(n_1825));
	notech_or2 i_656(.A(n_2303), .B(n_2285), .Z(n_1824));
	notech_and3 i_340(.A(n_2278), .B(n_2293), .C(n_29968), .Z(n_1822));
	notech_or2 i_652(.A(n_2285), .B(n_1822), .Z(n_1821));
	notech_or2 i_651(.A(n_2285), .B(n_2027), .Z(n_1820));
	notech_and2 i_647(.A(n_2295), .B(n_2302), .Z(n_1819));
	notech_and2 i_286(.A(n_2297), .B(n_30067), .Z(n_1818));
	notech_or4 i_621(.A(n_2348), .B(n_57703), .C(n_57735), .D(n_1818), .Z(n_1817
		));
	notech_or4 i_620(.A(n_2348), .B(n_57703), .C(n_57735), .D(n_2299), .Z(n_1813
		));
	notech_and4 i_615(.A(n_2278), .B(n_2275), .C(n_2302), .D(n_29968), .Z(n_1812
		));
	notech_ao3 i_531(.A(n_57868), .B(n_2324), .C(n_2330), .Z(n_1807));
	notech_or4 i_529(.A(n_57694), .B(n_2185), .C(n_57915), .D(n_57789), .Z(n_1806
		));
	notech_or4 i_502(.A(n_57805), .B(n_57771), .C(n_2297), .D(n_57845), .Z(n_1805
		));
	notech_and2 i_463(.A(n_2289), .B(n_2290), .Z(n_1802));
	notech_or2 i_23111433(.A(n_2337), .B(n_29968), .Z(n_1801));
	notech_or4 i_184(.A(n_2488), .B(n_30115), .C(n_30116), .D(n_30113), .Z(n_1800
		));
	notech_nand3 i_145(.A(n_57744), .B(n_2530), .C(n_57816), .Z(n_1798));
	notech_or4 i_839(.A(n_2313), .B(n_57735), .C(n_2280), .D(n_2290), .Z(n_1797
		));
	notech_or4 i_855(.A(n_2292), .B(n_2455), .C(n_57921), .D(n_57904), .Z(n_1796
		));
	notech_ao3 i_1104(.A(n_30056), .B(n_2321), .C(n_2101), .Z(n_1795));
	notech_or4 i_1225(.A(adz), .B(n_57780), .C(n_2347), .D(n_1916), .Z(n_1794
		));
	notech_or4 i_1291(.A(n_57805), .B(n_2448), .C(n_57841), .D(n_57816), .Z(n_1793
		));
	notech_or4 i_1233(.A(n_2347), .B(n_2284), .C(n_2018), .D(n_57780), .Z(n_1792
		));
	notech_nand3 i_520(.A(n_2278), .B(n_2299), .C(n_3761), .Z(n_1791));
	notech_and4 i_78571572(.A(n_1778), .B(n_3280), .C(n_3109), .D(n_1785), .Z
		(n_1789));
	notech_and4 i_78171576(.A(n_1950), .B(n_1638), .C(n_738), .D(n_3994), .Z
		(n_1785));
	notech_and4 i_78071577(.A(n_811), .B(n_3098), .C(n_2579), .D(n_3079), .Z
		(n_1778));
	notech_and4 i_11572301(.A(n_2571), .B(n_4013), .C(n_2394), .D(n_2365), .Z
		(n_1770));
	notech_and4 i_67371658(.A(n_1741), .B(n_1738), .C(n_176189124), .D(n_29994
		), .Z(n_1762));
	notech_and4 i_67071659(.A(n_1745), .B(n_1744), .C(n_1759), .D(n_1702), .Z
		(n_176189124));
	notech_and4 i_66871661(.A(n_3993), .B(n_1757), .C(n_2305), .D(n_1751), .Z
		(n_1759));
	notech_and4 i_66071668(.A(n_1793), .B(n_2894), .C(n_2136), .D(n_3152), .Z
		(n_1757));
	notech_and4 i_65971669(.A(n_2609), .B(n_2928), .C(n_1792), .D(n_2629), .Z
		(n_1751));
	notech_ao4 i_65871670(.A(n_30058), .B(n_57753), .C(n_30057), .D(n_4072),
		 .Z(n_1745));
	notech_ao4 i_65671671(.A(n_30060), .B(n_1802), .C(n_2124), .D(n_57859), 
		.Z(n_1744));
	notech_and4 i_66271666(.A(n_30102), .B(n_69847849), .C(n_29945), .D(n_2365
		), .Z(n_1741));
	notech_and4 i_66171667(.A(n_4056), .B(n_4036), .C(n_872), .D(n_29985), .Z
		(n_1738));
	notech_and3 i_31372283(.A(n_4014), .B(n_208149053), .C(n_29964), .Z(n_1734
		));
	notech_and4 i_46571827(.A(n_2894), .B(n_4055), .C(n_1725), .D(n_1699), .Z
		(n_1730));
	notech_and4 i_46071831(.A(n_4030), .B(n_2569), .C(n_1950), .D(n_29958), 
		.Z(n_1725));
	notech_nand3 i_25472288(.A(n_2076), .B(n_4055), .C(n_2620), .Z(n_1722)
		);
	notech_ao3 i_46471828(.A(n_1719), .B(n_1714), .C(n_1640), .Z(n_1721));
	notech_and4 i_45971832(.A(n_4031), .B(n_1014), .C(n_3993), .D(n_29986), 
		.Z(n_1719));
	notech_and4 i_45871833(.A(n_4026), .B(n_2760), .C(n_2479), .D(n_2690), .Z
		(n_1714));
	notech_and4 i_31272285(.A(n_4007), .B(n_4047), .C(n_2340), .D(n_2609), .Z
		(n_1709));
	notech_and4 i_11672300(.A(n_4086), .B(n_2538), .C(n_29988), .D(n_1704), 
		.Z(n_1708));
	notech_and3 i_8172303(.A(n_4002), .B(n_4076), .C(n_4027), .Z(n_1704));
	notech_and4 i_73572253(.A(n_29978), .B(n_1958), .C(n_2377), .D(n_29957),
		 .Z(n_1702));
	notech_and2 i_62272265(.A(n_2365), .B(n_29955), .Z(n_1699));
	notech_and4 i_13972115(.A(n_1801), .B(n_3402), .C(n_1694), .D(n_4093), .Z
		(n_1695));
	notech_and4 i_13772117(.A(n_2664), .B(n_2637), .C(n_2357), .D(n_3124), .Z
		(n_1694));
	notech_or4 i_13872116(.A(n_1795), .B(n_4024), .C(n_1626), .D(n_1625), .Z
		(n_1689));
	notech_and4 i_12572129(.A(n_2611), .B(n_2949), .C(n_2166), .D(n_2463), .Z
		(n_1684));
	notech_and4 i_12672128(.A(n_3013), .B(n_2480), .C(n_2729), .D(n_2959), .Z
		(n_1681));
	notech_ao3 i_8772160(.A(n_2743), .B(n_2623), .C(n_1675), .Z(n_1676));
	notech_nand3 i_32672281(.A(n_2019), .B(n_1616), .C(n_1618), .Z(n_1675)
		);
	notech_and4 i_8572162(.A(n_1671), .B(n_1668), .C(n_1664), .D(n_1661), .Z
		(n_1673));
	notech_and4 i_8072165(.A(n_247289127), .B(n_2045), .C(n_2591), .D(n_4030
		), .Z(n_1671));
	notech_and4 i_7972166(.A(n_2588), .B(n_3360), .C(n_2627), .D(n_29946), .Z
		(n_1668));
	notech_and4 i_7872167(.A(n_2744), .B(n_2140), .C(n_2516), .D(n_1942), .Z
		(n_1664));
	notech_ao3 i_7772168(.A(n_29930), .B(n_1619), .C(n_30079), .Z(n_1661));
	notech_and4 i_5972184(.A(n_4048), .B(n_164989123), .C(n_2036), .D(n_1653
		), .Z(n_1654));
	notech_and4 i_5772186(.A(n_30102), .B(n_2831), .C(n_2450), .D(n_2426), .Z
		(n_1653));
	notech_and2 i_5072192(.A(n_2398), .B(n_1834), .Z(n_164989123));
	notech_and4 i_5872185(.A(n_1644), .B(n_2305), .C(n_1612), .D(n_3984), .Z
		(n_1647));
	notech_ao4 i_5372189(.A(n_2166), .B(n_2006), .C(n_4071), .D(n_1965), .Z(n_1644
		));
	notech_nand3 i_52372274(.A(n_4025), .B(n_2629), .C(n_29989), .Z(n_1640)
		);
	notech_and4 i_50272327(.A(n_1770), .B(n_1789), .C(n_1709), .D(n_3197), .Z
		(n_1639));
	notech_or2 i_77371582(.A(n_2151), .B(n_57789), .Z(n_1638));
	notech_or2 i_71171633(.A(n_3958), .B(n_2359), .Z(n_1637));
	notech_nand3 i_55372332(.A(n_1762), .B(n_1734), .C(n_1629), .Z(\udeco[33] 
		));
	notech_nand2 i_64471679(.A(modrm[4]), .B(n_221891108), .Z(n_1629));
	notech_and4 i_60372340(.A(n_1730), .B(n_1709), .C(n_1708), .D(n_1721), .Z
		(n_1628));
	notech_or4 i_77672369(.A(n_1689), .B(n_1621), .C(n_30098), .D(n_2102), .Z
		(\udeco[110] ));
	notech_and2 i_12972125(.A(adz), .B(n_30089), .Z(n_1626));
	notech_and2 i_12872126(.A(adz), .B(n_29984), .Z(n_1625));
	notech_and4 i_372239(.A(n_2484), .B(n_1684), .C(n_1681), .D(n_1995), .Z(n_1622
		));
	notech_and2 i_13072124(.A(opz[2]), .B(n_30123), .Z(n_1621));
	notech_and4 i_91572372(.A(n_1676), .B(n_1673), .C(n_29947), .D(n_2435), 
		.Z(n_1620));
	notech_or4 i_6872176(.A(n_2289), .B(n_57771), .C(n_57744), .D(n_30051), 
		.Z(n_1619));
	notech_or4 i_6572179(.A(n_2311), .B(n_57915), .C(n_57789), .D(n_30051), 
		.Z(n_1618));
	notech_nao3 i_6672178(.A(n_57915), .B(n_57904), .C(n_3277), .Z(n_1616)
		);
	notech_and4 i_94372373(.A(n_1654), .B(n_1647), .C(n_1613), .D(n_1606), .Z
		(n_1614));
	notech_nand2 i_4772195(.A(modrm[1]), .B(n_30124), .Z(n_1613));
	notech_or2 i_4572197(.A(n_4070), .B(n_57753), .Z(n_1612));
	notech_and4 i_072242(.A(n_4034), .B(n_1865), .C(n_1604), .D(n_2883), .Z(n_1608
		));
	notech_nand3 i_62542(.A(n_2398), .B(n_2380), .C(n_29951), .Z(\udeco[4] )
		);
	notech_and4 i_62775(.A(n_2366), .B(n_1960), .C(n_29988), .D(n_122990279)
		, .Z(udeco_7397047));
	notech_and2 i_1072232(.A(modrm[4]), .B(n_30008), .Z(n_118490236));
	notech_or4 i_62806(.A(n_4024), .B(n_214991049), .C(n_3971), .D(n_118490236
		), .Z(\udeco[84] ));
	notech_and2 i_1372229(.A(n_57726), .B(n_30008), .Z(n_118590237));
	notech_or4 i_62811(.A(n_3971), .B(n_4045), .C(n_118590237), .D(n_123490283
		), .Z(\udeco[85] ));
	notech_nao3 i_10372314(.A(n_1960), .B(n_3998), .C(n_4057), .Z(\udeco[88] 
		));
	notech_or2 i_62823(.A(\udeco[88] ), .B(\udeco[5] ), .Z(\udeco[89] ));
	notech_or4 i_6972313(.A(n_30047), .B(\udeco[5] ), .C(n_30023), .D(n_3971
		), .Z(\udeco[91] ));
	notech_nao3 i_62826(.A(n_29962), .B(n_29990), .C(n_30054), .Z(\udeco[92] 
		));
	notech_nao3 i_11372312(.A(n_3998), .B(n_29962), .C(n_30054), .Z(\udeco[90] 
		));
	notech_or2 i_62828(.A(n_4057), .B(\udeco[90] ), .Z(\udeco[93] ));
	notech_or2 i_62829(.A(n_4057), .B(\udeco[91] ), .Z(\udeco[95] ));
	notech_nao3 i_62830(.A(n_3998), .B(n_1960), .C(n_4010), .Z(\udeco[96] )
		);
	notech_or2 i_62832(.A(n_4010), .B(\udeco[88] ), .Z(\udeco[98] ));
	notech_or4 i_62834(.A(n_4024), .B(n_4057), .C(n_3971), .D(n_3985), .Z(\udeco[100] 
		));
	notech_and4 i_62835(.A(n_30063), .B(n_2623), .C(n_1960), .D(n_29990), .Z
		(udeco_10197046));
	notech_or4 i_62836(.A(n_4018), .B(n_3950), .C(\udeco[88] ), .D(n_4010), 
		.Z(\udeco[102] ));
	notech_nao3 i_28672374(.A(n_30125), .B(n_124590294), .C(n_124090289), .Z
		(\udeco[127] ));
	notech_nand3 i_272240(.A(n_2099), .B(n_3736), .C(n_1905), .Z(n_118690238
		));
	notech_nor2 i_9072157(.A(n_1984), .B(n_30108), .Z(n_118790239));
	notech_nand2 i_9172156(.A(n_57726), .B(n_3956), .Z(n_118890240));
	notech_and2 i_9272155(.A(modrm[2]), .B(n_118690238), .Z(n_118990241));
	notech_or4 i_88072371(.A(n_124090289), .B(n_126190307), .C(n_125490301),
		 .D(n_125190298), .Z(\udeco[118] ));
	notech_or4 i_69872370(.A(n_4024), .B(n_4057), .C(n_1675), .D(n_30000), .Z
		(\udeco[115] ));
	notech_or4 i_56172368(.A(n_128790328), .B(n_30003), .C(n_127390316), .D(n_207949052
		), .Z(\udeco[107] ));
	notech_nao3 i_16272095(.A(n_57904), .B(n_2397), .C(n_2403), .Z(n_119090242
		));
	notech_or4 i_16472094(.A(n_57694), .B(n_4090), .C(n_2315), .D(modrm[5]),
		 .Z(n_119190243));
	notech_nand2 i_16872091(.A(opz[2]), .B(n_29974), .Z(n_119290244));
	notech_nand3 i_20272367(.A(n_119190243), .B(n_119090242), .C(n_129790337
		), .Z(\udeco[106] ));
	notech_or2 i_17872083(.A(n_2278), .B(n_2052), .Z(n_119490245));
	notech_nand2 i_17972082(.A(opz[1]), .B(n_29974), .Z(n_119590246));
	notech_nand3 i_72572366(.A(n_119190243), .B(n_130990344), .C(n_119090242
		), .Z(\udeco[105] ));
	notech_and4 i_20572365(.A(n_1969), .B(n_2623), .C(n_1960), .D(n_30063), 
		.Z(udeco_10397045));
	notech_and2 i_19272069(.A(modrm[7]), .B(n_30008), .Z(n_119690247));
	notech_or4 i_72172364(.A(n_30054), .B(n_214991049), .C(n_3971), .D(n_119690247
		), .Z(\udeco[87] ));
	notech_and2 i_19572066(.A(modrm[6]), .B(n_30008), .Z(n_119790248));
	notech_or4 i_72110266(.A(n_30054), .B(n_214991049), .C(n_3971), .D(n_119790248
		), .Z(\udeco[86] ));
	notech_or4 i_62833(.A(n_4024), .B(n_4057), .C(n_4010), .D(n_3971), .Z(\udeco[99] 
		));
	notech_nand2 i_19972062(.A(modrm[3]), .B(n_30008), .Z(n_119890249));
	notech_or4 i_71872363(.A(n_214991049), .B(n_4009), .C(\udeco[99] ), .D(n_131590350
		), .Z(\udeco[83] ));
	notech_nand2 i_21172055(.A(modrm[2]), .B(n_30008), .Z(n_120190252));
	notech_nand3 i_71572362(.A(n_131890353), .B(n_131790352), .C(n_132290355
		), .Z(\udeco[82] ));
	notech_or4 i_21772049(.A(n_2386), .B(n_57890), .C(n_57859), .D(n_29995),
		 .Z(n_120290253));
	notech_or4 i_22072047(.A(n_57805), .B(n_2182), .C(n_57816), .D(n_57825),
		 .Z(n_120490255));
	notech_and2 i_22172046(.A(modrm[1]), .B(n_30008), .Z(n_120590256));
	notech_or4 i_71272361(.A(n_30101), .B(n_120590256), .C(n_30054), .D(n_133190361
		), .Z(\udeco[81] ));
	notech_or4 i_22272360(.A(n_4011), .B(n_4018), .C(\udeco[91] ), .D(n_30005
		), .Z(\udeco[80] ));
	notech_nao3 i_10472307(.A(n_122990279), .B(n_1960), .C(n_133790365), .Z(\udeco[74] 
		));
	notech_or4 i_21610269(.A(n_29950), .B(n_29949), .C(\udeco[74] ), .D(n_3968
		), .Z(\udeco[78] ));
	notech_nao3 i_20510272(.A(n_29992), .B(n_30125), .C(n_133890366), .Z(\udeco[77] 
		));
	notech_or4 i_22872359(.A(n_133890366), .B(n_1326), .C(n_3971), .D(n_3978
		), .Z(\udeco[75] ));
	notech_nand3 i_22210281(.A(n_131790352), .B(n_135390376), .C(n_122990279
		), .Z(\udeco[72] ));
	notech_or4 i_70972358(.A(n_124090289), .B(n_136290384), .C(n_29949), .D(n_3969
		), .Z(\udeco[70] ));
	notech_nao3 i_11472306(.A(n_29975), .B(n_29957), .C(n_136290384), .Z(\udeco[71] 
		));
	notech_or4 i_70572357(.A(n_4009), .B(n_3969), .C(n_136290384), .D(n_3968
		), .Z(\udeco[68] ));
	notech_or4 i_20972356(.A(n_29949), .B(\udeco[71] ), .C(\udeco[5] ), .D(n_214991049
		), .Z(\udeco[67] ));
	notech_or4 i_20210288(.A(n_4045), .B(n_136290384), .C(n_136390385), .D(n_29950
		), .Z(\udeco[69] ));
	notech_or2 i_70272355(.A(n_4057), .B(\udeco[69] ), .Z(\udeco[66] ));
	notech_or4 i_69810292(.A(n_135690378), .B(n_30028), .C(n_136090382), .D(n_137390394
		), .Z(\udeco[65] ));
	notech_or4 i_69810296(.A(n_135690378), .B(n_30028), .C(n_136090382), .D(n_137790398
		), .Z(\udeco[64] ));
	notech_or4 i_69472354(.A(n_4054), .B(n_139390411), .C(n_4015), .D(n_138990407
		), .Z(\udeco[63] ));
	notech_or4 i_68372353(.A(n_121190261), .B(n_139390411), .C(n_124090289),
		 .D(n_138990407), .Z(\udeco[62] ));
	notech_nao3 i_68972352(.A(n_140090418), .B(n_30007), .C(n_124090289), .Z
		(\udeco[61] ));
	notech_or4 i_59272351(.A(n_140590422), .B(n_140290420), .C(n_4015), .D(n_4054
		), .Z(\udeco[60] ));
	notech_nand3 i_68310301(.A(n_138490402), .B(n_141290429), .C(n_30006), .Z
		(\udeco[59] ));
	notech_nand3 i_67872350(.A(n_2579), .B(n_138490402), .C(n_142390438), .Z
		(\udeco[58] ));
	notech_or4 i_67272349(.A(n_135890380), .B(n_135790379), .C(n_140290420),
		 .D(n_142690440), .Z(\udeco[57] ));
	notech_ao4 i_105872245(.A(n_2210), .B(n_3959), .C(n_30059), .D(n_29922),
		 .Z(n_121190261));
	notech_or4 i_66772348(.A(n_142990443), .B(n_121190261), .C(n_143290446),
		 .D(n_140290420), .Z(\udeco[56] ));
	notech_or4 i_66210306(.A(n_144190454), .B(n_4011), .C(n_1640), .D(n_30091
		), .Z(\udeco[55] ));
	notech_nao3 i_65772347(.A(n_143890451), .B(n_144890461), .C(n_124090289)
		, .Z(\udeco[54] ));
	notech_or4 i_65272346(.A(n_30012), .B(n_146190473), .C(n_221891108), .D(n_30028
		), .Z(\udeco[53] ));
	notech_or4 i_64572345(.A(n_146490476), .B(n_30091), .C(n_30011), .D(n_122890278
		), .Z(\udeco[52] ));
	notech_or4 i_64172344(.A(n_135890380), .B(n_135790379), .C(n_30091), .D(n_148390489
		), .Z(\udeco[51] ));
	notech_ao3 i_39471893(.A(n_30116), .B(modrm[3]), .C(n_2113), .Z(n_121290262
		));
	notech_or4 i_63572343(.A(n_30028), .B(n_30012), .C(n_124090289), .D(n_149990503
		), .Z(\udeco[50] ));
	notech_or4 i_41171876(.A(n_2118), .B(n_57921), .C(n_57789), .D(n_57762),
		 .Z(n_121390263));
	notech_nao3 i_61972342(.A(n_150990512), .B(n_143890451), .C(n_30091), .Z
		(\udeco[48] ));
	notech_or4 i_62372341(.A(n_152490527), .B(n_151290515), .C(n_139190409),
		 .D(n_29996), .Z(\udeco[47] ));
	notech_or4 i_61910310(.A(n_1640), .B(n_30017), .C(n_152790529), .D(n_153690537
		), .Z(\udeco[46] ));
	notech_or4 i_61572339(.A(n_155190547), .B(n_151790520), .C(n_154990545),
		 .D(n_29996), .Z(\udeco[44] ));
	notech_or4 i_35372338(.A(n_221891108), .B(n_29993), .C(n_30022), .D(n_157290565
		), .Z(\udeco[43] ));
	notech_or2 i_49871794(.A(n_5254), .B(n_57717), .Z(n_121490264));
	notech_or4 i_60972337(.A(n_30022), .B(n_157490567), .C(n_159190581), .D(n_29997
		), .Z(\udeco[42] ));
	notech_or4 i_60310317(.A(n_30091), .B(n_151790520), .C(n_161090596), .D(n_135990381
		), .Z(\udeco[41] ));
	notech_ao4 i_472238(.A(n_4065), .B(n_2320), .C(n_57735), .D(n_2371), .Z(n_121890268
		));
	notech_nor2 i_54371756(.A(n_5254), .B(n_30115), .Z(n_121990269));
	notech_nor2 i_54471755(.A(n_2275), .B(n_121890268), .Z(n_122090270));
	notech_or4 i_59672336(.A(n_161690601), .B(n_162590607), .C(n_152790529),
		 .D(n_151290515), .Z(\udeco[40] ));
	notech_nand3 i_59210322(.A(n_163990618), .B(n_163690615), .C(n_163290612
		), .Z(\udeco[39] ));
	notech_or4 i_58772335(.A(n_164890627), .B(n_164590624), .C(n_155190547),
		 .D(n_30027), .Z(\udeco[38] ));
	notech_nao3 i_57572334(.A(n_1734), .B(n_166590641), .C(n_221891108), .Z(\udeco[36] 
		));
	notech_nao3 i_61071702(.A(n_57744), .B(n_57904), .C(n_2564), .Z(n_122190271
		));
	notech_and4 i_56872333(.A(n_1193), .B(n_168390658), .C(n_167590651), .D(n_1734
		), .Z(udeco_3597044));
	notech_nand3 i_53972331(.A(n_170790679), .B(n_169190666), .C(n_1960), .Z
		(\udeco[31] ));
	notech_or4 i_53172330(.A(n_221891108), .B(n_30040), .C(n_204849027), .D(n_172790695
		), .Z(\udeco[30] ));
	notech_and4 i_52272329(.A(n_169090665), .B(n_1770), .C(n_174390708), .D(n_3109
		), .Z(udeco_2997043));
	notech_and4 i_51272328(.A(n_175090714), .B(n_176290724), .C(n_3510), .D(n_169190666
		), .Z(udeco_2897042));
	notech_or4 i_78871569(.A(n_2347), .B(n_2338), .C(n_3961), .D(n_57780), .Z
		(n_122290272));
	notech_nao3 i_46172326(.A(n_179190743), .B(n_1699), .C(n_30036), .Z(\udeco[22] 
		));
	notech_and4 i_45172325(.A(n_179490746), .B(n_182090769), .C(n_1925), .D(n_222291111
		), .Z(udeco_2197041));
	notech_or4 i_42472324(.A(n_30040), .B(n_30091), .C(n_30039), .D(n_184390787
		), .Z(\udeco[19] ));
	notech_and4 i_37272323(.A(n_185990802), .B(n_185590799), .C(n_185390797)
		, .D(n_3403), .Z(udeco_1597040));
	notech_and4 i_36972322(.A(n_187290812), .B(n_186790809), .C(n_151890521)
		, .D(n_3403), .Z(udeco_1497039));
	notech_nor2 i_88671476(.A(n_3954), .B(n_3958), .Z(n_122390273));
	notech_and4 i_35310360(.A(n_188090820), .B(n_187790817), .C(n_189290832)
		, .D(n_29964), .Z(udeco_1297038));
	notech_nand2 i_29510365(.A(n_68), .B(n_30048), .Z(\udeco[6] ));
	notech_or2 i_91271450(.A(n_2398), .B(n_57789), .Z(n_122490274));
	notech_nand3 i_29072321(.A(n_122490274), .B(n_29972), .C(n_30048), .Z(\udeco[3] 
		));
	notech_nor2 i_91671447(.A(n_2398), .B(n_57825), .Z(n_122590275));
	notech_or4 i_29010369(.A(n_1967), .B(n_30049), .C(n_122590275), .D(n_189790837
		), .Z(\udeco[2] ));
	notech_nor2 i_92071443(.A(n_2398), .B(n_57753), .Z(n_122690276));
	notech_or4 i_28610374(.A(n_190090839), .B(n_4006), .C(n_122690276), .D(n_30050
		), .Z(\udeco[1] ));
	notech_nand2 i_35472280(.A(n_1958), .B(n_4066), .Z(n_122890278));
	notech_and3 i_68672260(.A(n_3992), .B(n_3876), .C(n_29998), .Z(n_122990279
		));
	notech_nao3 i_1572227(.A(n_1950), .B(n_2380), .C(n_214991049), .Z(n_123490283
		));
	notech_nao3 i_6372304(.A(n_29975), .B(n_29973), .C(n_1640), .Z(n_124090289
		));
	notech_and4 i_3472208(.A(n_4017), .B(n_1920), .C(n_2450), .D(n_29991), .Z
		(n_124390292));
	notech_and4 i_3672206(.A(n_4048), .B(n_2195), .C(n_124390292), .D(n_2435
		), .Z(n_124590294));
	notech_or4 i_10072147(.A(n_30016), .B(n_4003), .C(n_1180), .D(n_3985), .Z
		(n_125190298));
	notech_or4 i_10172146(.A(n_222591114), .B(n_30084), .C(n_30088), .D(n_4080
		), .Z(n_125490301));
	notech_and4 i_9972148(.A(n_2516), .B(n_3733), .C(n_2332), .D(n_118890240
		), .Z(n_125890305));
	notech_or4 i_10672143(.A(n_118790239), .B(n_118990241), .C(n_3974), .D(n_29999
		), .Z(n_126190307));
	notech_and4 i_11272137(.A(n_1543), .B(n_1923), .C(n_4061), .D(n_1545), .Z
		(n_126990312));
	notech_or4 i_15272103(.A(n_222991118), .B(n_30001), .C(n_1262), .D(n_30002
		), .Z(n_127390316));
	notech_and4 i_15372102(.A(n_4084), .B(n_3991), .C(n_2162), .D(n_4004), .Z
		(n_127690319));
	notech_nand2 i_14472110(.A(n_4061), .B(n_2792), .Z(n_128190324));
	notech_or4 i_15472101(.A(n_4024), .B(n_29976), .C(n_29963), .D(n_128190324
		), .Z(n_128390326));
	notech_or4 i_16072097(.A(n_30094), .B(n_4009), .C(n_128390326), .D(n_30036
		), .Z(n_128790328));
	notech_and4 i_17572086(.A(n_1678), .B(n_208390990), .C(n_2623), .D(n_29990
		), .Z(n_129690336));
	notech_and4 i_17672085(.A(n_129690336), .B(n_29975), .C(n_4087), .D(n_119290244
		), .Z(n_129790337));
	notech_and4 i_18572076(.A(n_4043), .B(n_4087), .C(n_1678), .D(n_208390990
		), .Z(n_130190339));
	notech_and3 i_18472077(.A(n_2049), .B(n_3998), .C(n_119590246), .Z(n_130790342
		));
	notech_and4 i_18772074(.A(n_119490245), .B(n_130790342), .C(n_130190339)
		, .D(n_2380), .Z(n_130990344));
	notech_nao3 i_20472060(.A(n_4093), .B(n_119890249), .C(n_29950), .Z(n_131590350
		));
	notech_and2 i_69172257(.A(n_2366), .B(n_30122), .Z(n_131790352));
	notech_ao4 i_21372053(.A(n_2383), .B(n_2167), .C(n_3963), .D(n_2182), .Z
		(n_131890353));
	notech_and4 i_21472052(.A(n_29992), .B(n_29988), .C(n_2357), .D(n_120190252
		), .Z(n_132290355));
	notech_ao4 i_22572043(.A(n_2383), .B(n_2182), .C(n_2167), .D(n_30051), .Z
		(n_133090360));
	notech_nand3 i_22772041(.A(n_120290253), .B(n_133090360), .C(n_29988), .Z
		(n_133190361));
	notech_ao4 i_23372037(.A(n_1953), .B(n_30113), .C(n_2577), .D(n_3935), .Z
		(n_133490363));
	notech_nao3 i_80372247(.A(n_2629), .B(n_1953), .C(n_4011), .Z(n_133790365
		));
	notech_nao3 i_16972294(.A(n_5254), .B(n_29998), .C(n_133790365), .Z(n_133890366
		));
	notech_and3 i_25072020(.A(n_3970), .B(n_120490255), .C(n_30058), .Z(n_134990372
		));
	notech_ao4 i_24972021(.A(n_29995), .B(n_2167), .C(n_57694), .D(n_2368), 
		.Z(n_135190374));
	notech_and4 i_25272018(.A(n_135190374), .B(n_2151), .C(n_30095), .D(n_134990372
		), .Z(n_135390376));
	notech_nand2 i_55172272(.A(n_2123), .B(n_4034), .Z(n_135690378));
	notech_or2 i_80572246(.A(n_135690378), .B(n_30028), .Z(n_135790379));
	notech_or2 i_25772015(.A(n_29983), .B(n_4024), .Z(n_135890380));
	notech_or4 i_15672297(.A(n_4024), .B(n_29983), .C(n_135690378), .D(n_30028
		), .Z(n_135990381));
	notech_nand3 i_64272263(.A(n_4056), .B(n_4044), .C(n_3964), .Z(n_136090382
		));
	notech_or4 i_235572243(.A(n_4091), .B(n_136090382), .C(n_135890380), .D(n_135790379
		), .Z(n_136290384));
	notech_or4 i_25972013(.A(n_4011), .B(n_1640), .C(n_4009), .D(n_3969), .Z
		(n_136390385));
	notech_nand3 i_65172261(.A(n_5254), .B(n_2377), .C(n_1958), .Z(n_136890390
		));
	notech_or2 i_73072255(.A(n_29983), .B(n_30023), .Z(n_136990391));
	notech_or4 i_27272001(.A(n_30047), .B(n_3978), .C(n_136990391), .D(n_136890390
		), .Z(n_137390394));
	notech_or4 i_27771996(.A(n_30047), .B(n_4091), .C(n_136990391), .D(n_133790365
		), .Z(n_137790398));
	notech_and4 i_8272302(.A(n_2094), .B(n_210391008), .C(n_2569), .D(n_1905
		), .Z(n_138490402));
	notech_and4 i_28571989(.A(n_3979), .B(n_29991), .C(n_29957), .D(n_1978),
		 .Z(n_138790405));
	notech_nand3 i_11772299(.A(n_138490402), .B(n_138790405), .C(n_1193), .Z
		(n_138990407));
	notech_and2 i_62072267(.A(n_29959), .B(n_29954), .Z(n_139090408));
	notech_or2 i_59772270(.A(n_4006), .B(n_4024), .Z(n_139190409));
	notech_or4 i_28871987(.A(n_4024), .B(n_4006), .C(n_4091), .D(n_30018), .Z
		(n_139390411));
	notech_and4 i_29771979(.A(n_2327), .B(n_2623), .C(n_29958), .D(n_2305), 
		.Z(n_139790415));
	notech_and4 i_30071976(.A(n_139790415), .B(n_131790352), .C(n_139090408)
		, .D(n_30006), .Z(n_140090418));
	notech_nand2 i_62172266(.A(n_2579), .B(n_138490402), .Z(n_140290420));
	notech_or4 i_30471972(.A(n_4006), .B(n_4091), .C(n_222491113), .D(n_30018
		), .Z(n_140590422));
	notech_and4 i_31171965(.A(n_1978), .B(n_30102), .C(n_2304), .D(n_1816), 
		.Z(n_141190428));
	notech_and4 i_31471964(.A(n_141190428), .B(n_1953), .C(n_2623), .D(n_29959
		), .Z(n_141290429));
	notech_and3 i_81472244(.A(n_29961), .B(n_29954), .C(n_2380), .Z(n_141590432
		));
	notech_and4 i_32171957(.A(n_139790415), .B(n_30102), .C(n_2357), .D(n_30009
		), .Z(n_142190436));
	notech_and4 i_32571954(.A(n_30006), .B(n_1193), .C(n_141590432), .D(n_142190436
		), .Z(n_142390438));
	notech_nao3 i_32971951(.A(n_29958), .B(n_139090408), .C(n_4091), .Z(n_142690440
		));
	notech_nao3 i_33571945(.A(n_1953), .B(n_1950), .C(n_4009), .Z(n_142990443
		));
	notech_or4 i_33671944(.A(n_4091), .B(n_2307), .C(n_29983), .D(n_2165), .Z
		(n_143290446));
	notech_and4 i_32272282(.A(n_4031), .B(n_69847849), .C(n_2304), .D(n_29972
		), .Z(n_143890451));
	notech_or4 i_34471936(.A(n_3986), .B(n_210191006), .C(n_30035), .D(n_30010
		), .Z(n_144190454));
	notech_and4 i_35071930(.A(n_29978), .B(n_29987), .C(n_2365), .D(n_1972),
		 .Z(n_144690459));
	notech_and4 i_35271928(.A(n_30064), .B(n_144690459), .C(n_29998), .D(n_29986
		), .Z(n_144890461));
	notech_nand2 i_35871924(.A(n_222791116), .B(n_4016), .Z(n_145190463));
	notech_and4 i_36471918(.A(n_2365), .B(n_2099), .C(n_2327), .D(n_29987), 
		.Z(n_145590467));
	notech_nao3 i_36771916(.A(n_145590467), .B(n_2380), .C(n_145190463), .Z(n_145690468
		));
	notech_or4 i_36671917(.A(n_4045), .B(n_210191006), .C(n_4091), .D(n_29984
		), .Z(n_145990471));
	notech_or4 i_37071914(.A(n_145990471), .B(n_30094), .C(n_4009), .D(n_145690468
		), .Z(n_146190473));
	notech_or4 i_37871908(.A(n_30096), .B(n_30080), .C(n_30082), .D(n_4024),
		 .Z(n_146490476));
	notech_and4 i_37971907(.A(n_3360), .B(n_2099), .C(n_69847849), .D(n_29957
		), .Z(n_146990479));
	notech_and4 i_38871899(.A(n_222791116), .B(n_1737), .C(n_5254), .D(n_4031
		), .Z(n_147990486));
	notech_and4 i_38971898(.A(n_3982), .B(n_147990486), .C(n_2614), .D(n_29972
		), .Z(n_148190487));
	notech_nand3 i_39171896(.A(n_148190487), .B(n_141590432), .C(n_1702), .Z
		(n_148390489));
	notech_or4 i_39571892(.A(n_4023), .B(n_30081), .C(n_30094), .D(n_3990), 
		.Z(n_148690492));
	notech_or4 i_40471883(.A(n_121290262), .B(n_148690492), .C(n_1326), .D(n_4045
		), .Z(n_148890494));
	notech_or4 i_40371884(.A(n_4091), .B(n_3968), .C(n_4088), .D(n_30014), .Z
		(n_149590500));
	notech_or4 i_40571882(.A(n_209691002), .B(n_4052), .C(n_145190463), .D(n_149590500
		), .Z(n_149790501));
	notech_or4 i_40871879(.A(n_148890494), .B(n_30035), .C(n_149790501), .D(n_135690378
		), .Z(n_149990503));
	notech_and4 i_41771870(.A(n_3979), .B(n_2366), .C(n_30102), .D(n_210091005
		), .Z(n_150390507));
	notech_ao3 i_41671871(.A(n_210491009), .B(n_121390263), .C(n_222391112),
		 .Z(n_150790510));
	notech_and4 i_41971868(.A(n_150390507), .B(n_150790510), .C(n_2380), .D(n_29988
		), .Z(n_150990512));
	notech_nand3 i_25372289(.A(n_843), .B(n_4047), .C(n_4067), .Z(n_151290515
		));
	notech_and4 i_42871860(.A(n_4051), .B(n_4007), .C(n_4025), .D(n_4085), .Z
		(n_151690519));
	notech_nand3 i_17472293(.A(n_3993), .B(n_4055), .C(n_151690519), .Z(n_151790520
		));
	notech_and2 i_73772252(.A(n_29980), .B(n_29965), .Z(n_151890521));
	notech_and4 i_43271856(.A(n_4019), .B(n_1014), .C(n_2116), .D(n_29986), 
		.Z(n_152190524));
	notech_nao3 i_43371855(.A(n_29975), .B(n_152190524), .C(n_4088), .Z(n_152290525
		));
	notech_or4 i_43671852(.A(n_4035), .B(n_151790520), .C(n_4033), .D(n_152290525
		), .Z(n_152490527));
	notech_nand2 i_73872251(.A(n_4085), .B(n_1704), .Z(n_152790529));
	notech_and4 i_44371845(.A(n_3982), .B(n_1623), .C(n_29975), .D(n_29987),
		 .Z(n_153390534));
	notech_and4 i_44471844(.A(n_3064), .B(n_3360), .C(n_153390534), .D(n_29954
		), .Z(n_153490535));
	notech_or2 i_44671842(.A(n_139190409), .B(n_30033), .Z(n_153690537));
	notech_and4 i_47371819(.A(n_2017), .B(n_29965), .C(n_29980), .D(n_3980),
		 .Z(n_154290540));
	notech_and4 i_47471818(.A(n_5254), .B(n_4019), .C(n_3064), .D(n_2304), .Z
		(n_154790543));
	notech_nao3 i_47671816(.A(n_154790543), .B(n_154290540), .C(n_151290515)
		, .Z(n_154990545));
	notech_or4 i_36572279(.A(n_4050), .B(n_4054), .C(n_4059), .D(n_4024), .Z
		(n_155190547));
	notech_or4 i_48771805(.A(n_4023), .B(n_4059), .C(n_30097), .D(n_223091119
		), .Z(n_155890553));
	notech_or4 i_49271800(.A(n_1987), .B(n_30068), .C(n_1722), .D(n_155890553
		), .Z(n_156090555));
	notech_nand3 i_48371809(.A(n_1798), .B(n_1796), .C(n_4025), .Z(n_156390557
		));
	notech_or4 i_48971803(.A(n_2307), .B(n_222391112), .C(n_30081), .D(n_30105
		), .Z(n_156790561));
	notech_or4 i_49171801(.A(n_30096), .B(n_4050), .C(n_156390557), .D(n_156790561
		), .Z(n_156890562));
	notech_or4 i_49571797(.A(n_156090555), .B(n_156890562), .C(n_1086), .D(n_30033
		), .Z(n_157290565));
	notech_or4 i_51071783(.A(n_4035), .B(n_4033), .C(n_29983), .D(n_30023), 
		.Z(n_157490567));
	notech_and4 i_50671787(.A(n_210391008), .B(n_69847849), .C(n_2365), .D(n_3993
		), .Z(n_158390573));
	notech_and4 i_50871785(.A(n_3994), .B(n_3996), .C(n_158390573), .D(n_121490264
		), .Z(n_158490574));
	notech_and4 i_50771786(.A(n_2623), .B(n_29991), .C(n_29992), .D(n_4030),
		 .Z(n_158890578));
	notech_and4 i_51371781(.A(n_158890578), .B(n_141590432), .C(n_2116), .D(n_29975
		), .Z(n_159090580));
	notech_nand3 i_51571779(.A(n_222291111), .B(n_158490574), .C(n_159090580
		), .Z(n_159190581));
	notech_ao4 i_52871768(.A(n_5254), .B(n_30116), .C(n_4065), .D(n_2018), .Z
		(n_159490583));
	notech_and4 i_52971767(.A(n_1728), .B(n_4032), .C(n_4056), .D(n_4082), .Z
		(n_159790586));
	notech_and4 i_53071766(.A(n_2760), .B(n_3064), .C(n_214591046), .D(n_29955
		), .Z(n_160190590));
	notech_and4 i_53271765(.A(n_2569), .B(n_29958), .C(n_222791116), .D(n_4086
		), .Z(n_160690593));
	notech_and4 i_53571762(.A(n_160690593), .B(n_160190590), .C(n_159790586)
		, .D(n_159490583), .Z(n_160890595));
	notech_nand2 i_53671761(.A(n_160890595), .B(n_1704), .Z(n_161090596));
	notech_or4 i_55671745(.A(n_156390557), .B(n_4006), .C(n_30099), .D(n_122090270
		), .Z(n_161690601));
	notech_and4 i_55271748(.A(n_1014), .B(n_1951), .C(n_4007), .D(n_1815), .Z
		(n_162290606));
	notech_or4 i_55571746(.A(n_4001), .B(n_2164), .C(n_121990269), .D(n_30024
		), .Z(n_162590607));
	notech_and4 i_57171733(.A(n_2036), .B(n_2569), .C(n_29957), .D(n_30122),
		 .Z(n_163290612));
	notech_and4 i_56971735(.A(n_1332), .B(n_3967), .C(n_212091022), .D(n_211791020
		), .Z(n_163690615));
	notech_and4 i_57071734(.A(n_2176), .B(n_3979), .C(n_901), .D(n_3965), .Z
		(n_163990618));
	notech_and4 i_58071725(.A(n_2176), .B(n_901), .C(n_894), .D(n_212491025)
		, .Z(n_164490623));
	notech_nand3 i_58271723(.A(n_2036), .B(n_164490623), .C(n_29988), .Z(n_164590624
		));
	notech_or4 i_58171724(.A(n_30088), .B(n_1987), .C(n_30096), .D(n_4060), 
		.Z(n_164890627));
	notech_and4 i_60171709(.A(n_2569), .B(n_2015), .C(n_214591046), .D(n_29959
		), .Z(n_165390631));
	notech_and4 i_59871711(.A(n_1329), .B(n_3977), .C(n_861), .D(n_1537), .Z
		(n_165890634));
	notech_and4 i_59171715(.A(n_2663), .B(n_2327), .C(n_214091041), .D(n_853
		), .Z(n_165990635));
	notech_and4 i_60271708(.A(n_3967), .B(n_3965), .C(n_165990635), .D(n_165890634
		), .Z(n_166290638));
	notech_and4 i_60671705(.A(n_166290638), .B(n_165390631), .C(n_30019), .D
		(n_3107), .Z(n_166590641));
	notech_and4 i_63071689(.A(n_69847849), .B(n_1816), .C(n_29992), .D(n_29987
		), .Z(n_166990645));
	notech_and4 i_62771692(.A(n_222691115), .B(n_4051), .C(n_4029), .D(n_872
		), .Z(n_167390649));
	notech_and4 i_63371686(.A(n_167390649), .B(n_166990645), .C(n_2305), .D(n_122190271
		), .Z(n_167590651));
	notech_and4 i_61471698(.A(n_3062), .B(n_2500), .C(n_3736), .D(n_1905), .Z
		(n_167790653));
	notech_and4 i_62971690(.A(n_3994), .B(n_1593), .C(n_1329), .D(n_29985), 
		.Z(n_168290657));
	notech_and4 i_63271687(.A(n_2076), .B(n_4036), .C(n_167790653), .D(n_168290657
		), .Z(n_168390658));
	notech_and4 i_68171651(.A(n_3970), .B(n_1806), .C(n_730), .D(n_3079), .Z
		(n_168890663));
	notech_and4 i_68471649(.A(n_733), .B(n_738), .C(n_168890663), .D(n_3197)
		, .Z(n_169090665));
	notech_and2 i_26972287(.A(n_3109), .B(n_169090665), .Z(n_169190666));
	notech_and4 i_70171640(.A(n_2327), .B(n_4032), .C(n_853), .D(n_214091041
		), .Z(n_169490669));
	notech_and4 i_69971642(.A(n_717), .B(n_2246), .C(n_4014), .D(n_4013), .Z
		(n_169790672));
	notech_and3 i_69271646(.A(n_1984), .B(n_1801), .C(n_1993), .Z(n_169890673
		));
	notech_and4 i_70371639(.A(n_4034), .B(n_169790672), .C(n_4085), .D(n_169890673
		), .Z(n_170390676));
	notech_and4 i_70771636(.A(n_222291111), .B(n_169490669), .C(n_208149053)
		, .D(n_170390676), .Z(n_170790679));
	notech_and4 i_72371625(.A(n_214391044), .B(n_3992), .C(n_202790942), .D(n_692
		), .Z(n_171690685));
	notech_nand3 i_72771622(.A(n_171690685), .B(n_2627), .C(n_29961), .Z(n_171790686
		));
	notech_and4 i_72471624(.A(n_709), .B(n_719), .C(n_703), .D(n_4008), .Z(n_172190689
		));
	notech_and4 i_72671623(.A(n_2760), .B(n_4032), .C(n_3143), .D(n_3980), .Z
		(n_172490692));
	notech_or4 i_73371618(.A(n_30031), .B(n_171790686), .C(n_155190547), .D(n_30030
		), .Z(n_172790695));
	notech_and4 i_74771607(.A(n_4041), .B(n_4036), .C(n_720), .D(n_673), .Z(n_173390699
		));
	notech_and4 i_74871606(.A(n_214391044), .B(n_4028), .C(n_1718), .D(n_222891117
		), .Z(n_173890703));
	notech_and2 i_74571609(.A(n_1332), .B(n_212091022), .Z(n_174090705));
	notech_and4 i_75171603(.A(n_222691115), .B(n_4029), .C(n_174090705), .D(n_173890703
		), .Z(n_174290707));
	notech_and4 i_75271602(.A(n_173390699), .B(n_174290707), .C(n_1950), .D(n_29962
		), .Z(n_174390708));
	notech_and4 i_76371591(.A(n_2099), .B(n_4016), .C(n_4026), .D(n_2538), .Z
		(n_174790712));
	notech_and4 i_76871587(.A(n_4055), .B(n_2894), .C(n_174790712), .D(n_1770
		), .Z(n_175090714));
	notech_and4 i_76171593(.A(n_1290), .B(n_4014), .C(n_720), .D(n_1999), .Z
		(n_175690718));
	notech_and4 i_76271592(.A(n_1718), .B(n_3967), .C(n_29985), .D(n_2760), 
		.Z(n_175990721));
	notech_and4 i_77071585(.A(n_175990721), .B(n_175690718), .C(n_1960), .D(n_29964
		), .Z(n_176290724));
	notech_and2 i_77572249(.A(n_1434), .B(n_122290272), .Z(n_176690727));
	notech_and4 i_79871560(.A(n_4053), .B(n_200290921), .C(n_4027), .D(n_1615
		), .Z(n_177590733));
	notech_and4 i_80171557(.A(n_493), .B(n_4084), .C(n_177590733), .D(n_497)
		, .Z(n_177690734));
	notech_and2 i_79371564(.A(n_4038), .B(n_191190849), .Z(n_178190736));
	notech_and4 i_80071558(.A(n_1537), .B(n_2760), .C(n_2928), .D(n_2571), .Z
		(n_178790740));
	notech_and4 i_80271556(.A(n_178190736), .B(n_178790740), .C(n_2080), .D(n_1996
		), .Z(n_178990741));
	notech_and4 i_80871552(.A(n_177690734), .B(n_176690727), .C(n_3280), .D(n_178990741
		), .Z(n_179190743));
	notech_and4 i_82871533(.A(n_2928), .B(n_853), .C(n_730), .D(n_4047), .Z(n_179490746
		));
	notech_and4 i_82371538(.A(n_2678), .B(n_2791), .C(n_533), .D(n_2884), .Z
		(n_180090751));
	notech_and4 i_81271548(.A(n_2631), .B(n_1780), .C(n_2137), .D(n_2757), .Z
		(n_180390754));
	notech_and4 i_82571536(.A(n_2157), .B(n_2212), .C(n_4049), .D(n_2029), .Z
		(n_180790758));
	notech_and4 i_83071531(.A(n_574), .B(n_466), .C(n_180390754), .D(n_180790758
		), .Z(n_180890759));
	notech_and4 i_83371528(.A(n_4004), .B(n_2538), .C(n_180090751), .D(n_180890759
		), .Z(n_180990760));
	notech_and4 i_82671535(.A(n_3987), .B(n_537), .C(n_202090937), .D(n_1777
		), .Z(n_181290763));
	notech_and4 i_82771534(.A(n_3973), .B(n_4037), .C(n_1504), .D(n_4005), .Z
		(n_181790766));
	notech_and4 i_83671525(.A(n_181790766), .B(n_181290763), .C(n_2435), .D(n_180990760
		), .Z(n_182090769));
	notech_and4 i_85671505(.A(n_2398), .B(n_4004), .C(n_4084), .D(n_1923), .Z
		(n_182490772));
	notech_and4 i_85171510(.A(n_4002), .B(n_4076), .C(n_2377), .D(n_4064), .Z
		(n_183090777));
	notech_and4 i_85271509(.A(n_1970), .B(n_1526), .C(n_530), .D(n_2058), .Z
		(n_183590781));
	notech_ao3 i_84371518(.A(n_2216), .B(n_455), .C(n_1987), .Z(n_183890783)
		);
	notech_and4 i_85871503(.A(n_183590781), .B(n_1603), .C(n_3975), .D(n_183890783
		), .Z(n_184190785));
	notech_and4 i_86171500(.A(n_4017), .B(n_183090777), .C(n_184190785), .D(n_2380
		), .Z(n_184290786));
	notech_nand3 i_86371498(.A(n_182490772), .B(n_176690727), .C(n_184290786
		), .Z(n_184390787));
	notech_ao4 i_84571516(.A(n_3957), .B(n_3954), .C(n_3963), .D(n_2517), .Z
		(n_184590789));
	notech_and4 i_85571506(.A(n_3993), .B(n_493), .C(n_3973), .D(n_4085), .Z
		(n_184990793));
	notech_and4 i_85971502(.A(n_1306), .B(n_184590789), .C(n_184990793), .D(n_1340
		), .Z(n_185090794));
	notech_and3 i_76672250(.A(n_2141), .B(n_4013), .C(n_2484), .Z(n_185390797
		));
	notech_and4 i_86971492(.A(n_3374), .B(n_3880), .C(n_4079), .D(n_3981), .Z
		(n_185590799));
	notech_and4 i_87071491(.A(n_4046), .B(n_4053), .C(n_2171), .D(n_4058), .Z
		(n_185990802));
	notech_and4 i_87871483(.A(n_4084), .B(n_2394), .C(n_520), .D(n_3982), .Z
		(n_186490807));
	notech_and4 i_88371479(.A(n_444), .B(n_4046), .C(n_186490807), .D(n_185390797
		), .Z(n_186790809));
	notech_and4 i_87971482(.A(n_2024), .B(n_2047), .C(n_1780), .D(n_201490933
		), .Z(n_187290812));
	notech_and4 i_89671466(.A(n_1346), .B(n_204), .C(n_1284), .D(n_215), .Z(n_187790817
		));
	notech_and4 i_89771465(.A(n_2171), .B(n_530), .C(n_218), .D(n_254), .Z(n_188090820
		));
	notech_and4 i_89871464(.A(n_3975), .B(n_4085), .C(n_29987), .D(n_1615), 
		.Z(n_188590825));
	notech_ao3 i_89571467(.A(n_1130), .B(n_29965), .C(n_122390273), .Z(n_188990829
		));
	notech_and3 i_89971463(.A(n_69847849), .B(n_4004), .C(n_188990829), .Z(n_189090830
		));
	notech_and4 i_90471458(.A(n_189090830), .B(n_185390797), .C(n_2434), .D(n_188590825
		), .Z(n_189290832));
	notech_nao3 i_90671456(.A(n_1919), .B(n_29986), .C(n_2164), .Z(n_189490834
		));
	notech_or4 i_90971453(.A(n_29966), .B(n_189490834), .C(n_29984), .D(n_30046
		), .Z(n_189690836));
	notech_or4 i_14872298(.A(n_4011), .B(n_1640), .C(n_4009), .D(n_189690836
		), .Z(n_189790837));
	notech_or4 i_15872296(.A(n_124090289), .B(n_30047), .C(\udeco[5] ), .D(n_189690836
		), .Z(n_190090839));
	notech_nand3 i_10392112(.A(n_3779), .B(n_1865), .C(n_194990882), .Z(n_190890846
		));
	notech_and4 i_10292113(.A(n_2352), .B(n_2654), .C(n_1856), .D(n_2344), .Z
		(n_190990847));
	notech_or4 i_118392115(.A(n_57805), .B(n_3935), .C(n_57841), .D(n_57753)
		, .Z(n_191190849));
	notech_nand2 i_114092117(.A(modrm[3]), .B(n_30052), .Z(n_191390851));
	notech_and2 i_113792118(.A(n_3763), .B(n_29970), .Z(n_191490852));
	notech_and2 i_113992119(.A(modrm[0]), .B(n_190890846), .Z(n_191590853)
		);
	notech_or4 i_92992120(.A(n_1321), .B(n_191490852), .C(n_191590853), .D(n_30062
		), .Z(\udeco[124] ));
	notech_and3 i_33692122(.A(n_2302), .B(n_30067), .C(n_29968), .Z(n_191790855
		));
	notech_or4 i_116492123(.A(n_2348), .B(n_57703), .C(n_57735), .D(n_191790855
		), .Z(n_191890856));
	notech_nao3 i_116392124(.A(n_29924), .B(n_29921), .C(n_2318), .Z(n_191990857
		));
	notech_and4 i_89292125(.A(n_199890917), .B(n_199490914), .C(n_2694), .D(n_1942
		), .Z(udeco_11997037));
	notech_nand3 i_14892126(.A(n_3736), .B(n_2099), .C(n_1905), .Z(n_192190858
		));
	notech_or4 i_141092128(.A(n_57805), .B(n_2316), .C(n_2389), .D(n_3761), 
		.Z(n_192690860));
	notech_nand2 i_141292129(.A(modrm[0]), .B(n_192190858), .Z(n_192790861)
		);
	notech_and2 i_140992130(.A(modrm[3]), .B(n_3773), .Z(n_192990862));
	notech_and2 i_141192131(.A(n_29971), .B(n_30034), .Z(n_193090863));
	notech_or4 i_85092132(.A(n_1321), .B(n_192990862), .C(n_30070), .D(n_193090863
		), .Z(\udeco[116] ));
	notech_or4 i_144392133(.A(n_57694), .B(n_2373), .C(n_57717), .D(n_2401),
		 .Z(n_193190864));
	notech_and4 i_84292134(.A(n_204590959), .B(n_201790935), .C(n_2684), .D(n_2890
		), .Z(udeco_11497036));
	notech_and4 i_82092135(.A(n_2704), .B(n_2684), .C(n_207790985), .D(n_2890
		), .Z(udeco_11397035));
	notech_or4 i_168292136(.A(n_57694), .B(n_2373), .C(n_3845), .D(n_57726),
		 .Z(n_193290865));
	notech_or4 i_168692137(.A(n_57805), .B(n_2313), .C(n_57890), .D(n_2348),
		 .Z(n_193390866));
	notech_and2 i_168592138(.A(opz[0]), .B(n_29974), .Z(n_193490867));
	notech_or4 i_66292139(.A(n_193490867), .B(n_209290999), .C(n_30079), .D(n_30076
		), .Z(\udeco[104] ));
	notech_and2 i_12692140(.A(n_3992), .B(n_3876), .Z(n_5254));
	notech_nao3 i_62892144(.A(n_211491018), .B(n_5254), .C(n_210191006), .Z(\udeco[49] 
		));
	notech_or4 i_172392145(.A(n_57694), .B(n_2037), .C(n_4072), .D(n_57726),
		 .Z(n_193890871));
	notech_and4 i_58292146(.A(n_193890871), .B(n_213891039), .C(n_1593), .D(n_894
		), .Z(udeco_3797034));
	notech_nao3 i_175092149(.A(n_29924), .B(n_30059), .C(n_2499), .Z(n_194190874
		));
	notech_or2 i_174792150(.A(n_2124), .B(n_57780), .Z(n_194290875));
	notech_or4 i_174992151(.A(n_57694), .B(n_2315), .C(n_57717), .D(n_3836),
		 .Z(n_194390876));
	notech_nao3 i_56110330(.A(n_216891063), .B(n_214391044), .C(n_1326), .Z(\udeco[34] 
		));
	notech_or2 i_182692152(.A(n_2151), .B(n_57825), .Z(n_194490877));
	notech_or2 i_182892153(.A(n_3697), .B(n_57780), .Z(n_194590878));
	notech_or2 i_182792154(.A(n_3728), .B(n_57717), .Z(n_194690879));
	notech_nao3 i_49492155(.A(n_717), .B(n_219691088), .C(n_1326), .Z(\udeco[26] 
		));
	notech_and4 i_47210352(.A(n_520), .B(n_537), .C(n_2567), .D(n_221591105)
		, .Z(udeco_2397033));
	notech_nao3 i_34692156(.A(n_1951), .B(n_2380), .C(n_4057), .Z(n_1326));
	notech_or4 i_17292158(.A(n_1326), .B(n_30084), .C(n_29967), .D(n_3978), 
		.Z(n_1321));
	notech_ao3 i_113192160(.A(n_3777), .B(n_3987), .C(n_3846), .Z(n_194990882
		));
	notech_ao4 i_114292164(.A(n_57915), .B(n_4070), .C(n_2348), .D(n_2338), 
		.Z(n_195690886));
	notech_ao4 i_114392165(.A(n_2166), .B(n_3760), .C(n_30051), .D(n_3935), 
		.Z(n_195790887));
	notech_and4 i_114692168(.A(n_195790887), .B(n_195690886), .C(n_3834), .D
		(n_247289127), .Z(n_196290890));
	notech_and4 i_114992171(.A(n_2450), .B(n_196290890), .C(n_1834), .D(n_191390851
		), .Z(n_196590893));
	notech_and3 i_116692175(.A(n_2676), .B(n_191990857), .C(n_191890856), .Z
		(n_197390897));
	notech_nand2 i_14392177(.A(n_2629), .B(n_29989), .Z(n_1249));
	notech_nand2 i_22192179(.A(n_30102), .B(n_29992), .Z(n_1180));
	notech_and4 i_26692182(.A(n_2216), .B(n_2709), .C(n_2151), .D(n_30058), 
		.Z(n_1130));
	notech_and4 i_133192183(.A(n_2231), .B(n_1833), .C(n_2188), .D(n_1907), 
		.Z(n_197790901));
	notech_and4 i_133392186(.A(n_2630), .B(n_3733), .C(n_3993), .D(n_197790901
		), .Z(n_198190904));
	notech_and4 i_133692189(.A(n_198190904), .B(n_2638), .C(n_1130), .D(n_2065
		), .Z(n_198590907));
	notech_and3 i_133892191(.A(n_4002), .B(n_2166), .C(n_2829), .Z(n_198890909
		));
	notech_and4 i_134092193(.A(n_2827), .B(n_198590907), .C(n_198890909), .D
		(n_2414), .Z(n_199090911));
	notech_and4 i_134692196(.A(n_2826), .B(n_199090911), .C(n_2707), .D(n_1920
		), .Z(n_199490914));
	notech_and4 i_134592199(.A(n_2522), .B(n_2831), .C(n_2510), .D(n_2605), 
		.Z(n_199890917));
	notech_and2 i_61092202(.A(n_4029), .B(n_3967), .Z(n_200290921));
	notech_ao4 i_141392203(.A(n_1984), .B(n_57915), .C(n_2383), .D(n_2865), 
		.Z(n_200390922));
	notech_and4 i_141692206(.A(n_200390922), .B(n_2857), .C(n_192690860), .D
		(n_29972), .Z(n_200690925));
	notech_and4 i_141892208(.A(n_2479), .B(n_200690925), .C(n_29990), .D(n_30063
		), .Z(n_200890927));
	notech_and4 i_142192211(.A(n_200290921), .B(n_200890927), .C(n_2884), .D
		(n_192790861), .Z(n_201190930));
	notech_and2 i_61292214(.A(n_1993), .B(n_4040), .Z(n_201490933));
	notech_and4 i_146692216(.A(n_1993), .B(n_4040), .C(n_2309), .D(n_2483), 
		.Z(n_201790935));
	notech_and4 i_25792218(.A(n_1886), .B(n_2686), .C(n_2572), .D(n_2899), .Z
		(n_202090937));
	notech_and4 i_71092223(.A(n_4007), .B(n_3672), .C(n_1537), .D(n_193190864
		), .Z(n_202790942));
	notech_and4 i_144892226(.A(n_2629), .B(n_3964), .C(n_2709), .D(n_29975),
		 .Z(n_203190945));
	notech_and4 i_145192229(.A(n_2765), .B(n_3867), .C(n_203190945), .D(n_2124
		), .Z(n_203490948));
	notech_and3 i_145392231(.A(n_1949), .B(n_1796), .C(n_3880), .Z(n_203690950
		));
	notech_and4 i_145692233(.A(n_3777), .B(n_203490948), .C(n_1526), .D(n_203690950
		), .Z(n_203890952));
	notech_and4 i_145992236(.A(n_203890952), .B(n_198890909), .C(n_2655), .D
		(n_202790942), .Z(n_204190955));
	notech_and4 i_146592239(.A(n_2903), .B(n_2605), .C(n_204190955), .D(n_1504
		), .Z(n_204490958));
	notech_and4 i_146792240(.A(n_2898), .B(n_202090937), .C(n_2893), .D(n_204490958
		), .Z(n_204590959));
	notech_and4 i_148692246(.A(n_3994), .B(n_2839), .C(n_202790942), .D(n_2852
		), .Z(n_205490965));
	notech_ao3 i_147292249(.A(n_2516), .B(n_29973), .C(n_4010), .Z(n_205790968
		));
	notech_and4 i_147592252(.A(n_2765), .B(n_3931), .C(n_3751), .D(n_205790968
		), .Z(n_206190971));
	notech_and4 i_147892255(.A(n_2625), .B(n_2176), .C(n_206190971), .D(n_2591
		), .Z(n_206490974));
	notech_and4 i_148292258(.A(n_2332), .B(n_206490974), .C(n_2534), .D(n_2539
		), .Z(n_206890977));
	notech_and4 i_148792260(.A(n_2572), .B(n_1969), .C(n_206890977), .D(n_2656
		), .Z(n_207090979));
	notech_and4 i_149092263(.A(n_2722), .B(n_2898), .C(n_207090979), .D(n_2850
		), .Z(n_207390982));
	notech_and4 i_149292264(.A(n_4040), .B(n_205490965), .C(n_207390982), .D
		(n_1993), .Z(n_207490983));
	notech_and4 i_149492266(.A(n_2834), .B(n_2893), .C(n_207490983), .D(n_2688
		), .Z(n_207790985));
	notech_and2 i_72092269(.A(n_3973), .B(n_4029), .Z(n_843));
	notech_and4 i_26492272(.A(n_2327), .B(n_193290865), .C(n_3665), .D(n_30122
		), .Z(n_208390990));
	notech_and4 i_168992275(.A(n_3998), .B(n_193390866), .C(n_3890), .D(n_29975
		), .Z(n_208690993));
	notech_and4 i_169292278(.A(n_208690993), .B(n_1290), .C(n_2162), .D(n_2380
		), .Z(n_208990996));
	notech_or4 i_169592281(.A(n_3820), .B(n_29976), .C(n_1249), .D(n_30077),
		 .Z(n_209290999));
	notech_nand3 i_4353(.A(n_223489126), .B(n_1792), .C(n_1999), .Z(n_209691002
		));
	notech_and4 i_4356(.A(n_29978), .B(n_4019), .C(n_29979), .D(n_1972), .Z(n_210091005
		));
	notech_or4 i_37392286(.A(n_30096), .B(n_30080), .C(n_30082), .D(n_1180),
		 .Z(n_210191006));
	notech_and2 i_4347(.A(n_4026), .B(n_3982), .Z(n_69847849));
	notech_and2 i_4298(.A(n_3838), .B(n_3987), .Z(n_210391008));
	notech_ao4 i_65092288(.A(n_2113), .B(n_2373), .C(n_2278), .D(n_2346), .Z
		(n_210491009));
	notech_ao4 i_170692289(.A(n_2275), .B(n_2118), .C(n_2564), .D(n_57762), 
		.Z(n_210591010));
	notech_and4 i_170992292(.A(n_210591010), .B(n_210491009), .C(n_4031), .D
		(n_1816), .Z(n_210891013));
	notech_and4 i_171392295(.A(n_2340), .B(n_210891013), .C(n_2099), .D(n_210391008
		), .Z(n_211191016));
	notech_and4 i_171592297(.A(n_4032), .B(n_4030), .C(n_211191016), .D(n_69847849
		), .Z(n_211491018));
	notech_and4 i_80792299(.A(n_4076), .B(n_193890871), .C(n_2615), .D(n_2091
		), .Z(n_211791020));
	notech_ao3 i_4572(.A(n_4014), .B(n_1329), .C(n_29927), .Z(n_212091022)
		);
	notech_and4 i_173892302(.A(n_872), .B(n_2500), .C(n_212091022), .D(n_200290921
		), .Z(n_212291024));
	notech_and2 i_74292303(.A(n_3994), .B(n_4085), .Z(n_692));
	notech_and3 i_4510(.A(n_2629), .B(n_4086), .C(n_29989), .Z(n_212491025)
		);
	notech_and4 i_172692307(.A(n_3973), .B(n_3736), .C(n_4031), .D(n_1114), 
		.Z(n_212891029));
	notech_and4 i_172992310(.A(n_212891029), .B(n_2743), .C(n_3061), .D(n_29980
		), .Z(n_213191032));
	notech_and4 i_173392313(.A(n_4034), .B(n_213191032), .C(n_2465), .D(n_861
		), .Z(n_213491035));
	notech_and4 i_173792315(.A(n_2036), .B(n_1014), .C(n_213491035), .D(n_30104
		), .Z(n_213691037));
	notech_and4 i_174092317(.A(n_3994), .B(n_213691037), .C(n_212291024), .D
		(n_4085), .Z(n_213891039));
	notech_and4 i_4614(.A(n_2192), .B(n_4017), .C(n_2500), .D(n_3981), .Z(n_214091041
		));
	notech_and4 i_4656(.A(n_2663), .B(n_2327), .C(n_214091041), .D(n_30063),
		 .Z(n_214391044));
	notech_ao3 i_4531(.A(n_4041), .B(n_1896), .C(n_222391112), .Z(n_214591046
		));
	notech_nand2 i_351092324(.A(n_29992), .B(n_29988), .Z(n_214991049));
	notech_ao4 i_175192325(.A(n_57825), .B(n_30058), .C(n_57717), .D(n_30100
		), .Z(n_215091050));
	notech_and4 i_175492328(.A(n_215091050), .B(n_3992), .C(n_194190874), .D
		(n_30095), .Z(n_215491053));
	notech_and4 i_175992331(.A(n_215491053), .B(n_194290875), .C(n_2017), .D
		(n_194390876), .Z(n_215891056));
	notech_and4 i_176092332(.A(n_811), .B(n_2340), .C(n_214591046), .D(n_215891056
		), .Z(n_215991057));
	notech_and4 i_176392334(.A(n_4055), .B(n_2538), .C(n_843), .D(n_215991057
		), .Z(n_216191059));
	notech_and4 i_176492335(.A(n_2099), .B(n_216191059), .C(n_3736), .D(n_2116
		), .Z(n_216291060));
	notech_and4 i_176792338(.A(n_960), .B(n_894), .C(n_2903), .D(n_216291060
		), .Z(n_216891063));
	notech_and3 i_184492341(.A(n_3102), .B(n_738), .C(n_2588), .Z(n_217291066
		));
	notech_and4 i_184892343(.A(n_30063), .B(n_217291066), .C(n_3098), .D(n_29959
		), .Z(n_217491068));
	notech_and4 i_183192347(.A(n_4026), .B(n_4041), .C(n_4013), .D(n_3980), 
		.Z(n_217991072));
	notech_and3 i_183492349(.A(n_217991072), .B(n_2305), .C(n_29985), .Z(n_218191074
		));
	notech_and4 i_183892351(.A(n_1290), .B(n_194490877), .C(n_218191074), .D
		(n_194590878), .Z(n_218491076));
	notech_and4 i_183992355(.A(n_3103), .B(n_853), .C(n_2099), .D(n_2533), .Z
		(n_218891080));
	notech_and4 i_184392357(.A(n_218891080), .B(n_2465), .C(n_218491076), .D
		(n_2015), .Z(n_219091082));
	notech_and4 i_184992360(.A(n_219091082), .B(n_222891117), .C(n_29986), .D
		(n_194690879), .Z(n_219391085));
	notech_and4 i_185292363(.A(n_703), .B(n_2246), .C(n_219391085), .D(n_217491068
		), .Z(n_219691088));
	notech_and4 i_195592367(.A(n_3049), .B(n_2723), .C(n_2928), .D(n_2024), 
		.Z(n_220091092));
	notech_and3 i_194792370(.A(n_4048), .B(n_4047), .C(n_4019), .Z(n_220391095
		));
	notech_and4 i_195092373(.A(n_2365), .B(n_3739), .C(n_4049), .D(n_220391095
		), .Z(n_220691098));
	notech_and4 i_195692376(.A(n_2212), .B(n_2522), .C(n_200290921), .D(n_220691098
		), .Z(n_220991101));
	notech_and4 i_195992378(.A(n_2157), .B(n_220991101), .C(n_3177), .D(n_220091092
		), .Z(n_221191103));
	notech_and4 i_196192380(.A(n_1993), .B(n_4040), .C(n_221191103), .D(n_530
		), .Z(n_221591105));
	notech_nand3 i_20072319(.A(n_2123), .B(n_4034), .C(n_4022), .Z(n_221891108
		));
	notech_and2 i_413972309(.A(n_29961), .B(n_4062), .Z(n_2219));
	notech_and3 i_4288(.A(n_3992), .B(n_3876), .C(n_2377), .Z(n_222191110)
		);
	notech_and3 i_61772268(.A(n_4067), .B(n_4022), .C(n_29979), .Z(n_222291111
		));
	notech_and4 i_172241(.A(n_2344), .B(n_3279), .C(n_3545), .D(n_1856), .Z(n_1607
		));
	notech_ao3 i_16192383(.A(n_30121), .B(n_3895), .C(n_2348), .Z(n_222391112
		));
	notech_or2 i_3625(.A(n_4089), .B(n_4024), .Z(n_222491113));
	notech_nand3 i_3834(.A(n_2073), .B(n_2202), .C(n_4082), .Z(n_222591114)
		);
	notech_ao4 i_4638(.A(n_2303), .B(n_30066), .C(n_30055), .D(n_2291), .Z(n_222691115
		));
	notech_nand2 i_4672196(.A(modrm[4]), .B(n_30141), .Z(n_1606));
	notech_ao4 i_41792384(.A(n_4072), .B(n_30053), .C(n_30057), .D(n_4090), 
		.Z(n_222791116));
	notech_ao4 i_55992385(.A(n_3954), .B(n_3957), .C(n_2339), .D(n_2299), .Z
		(n_222891117));
	notech_nand3 i_69592386(.A(n_2587), .B(n_197390897), .C(n_2722), .Z(n_222991118
		));
	notech_nand3 i_79792387(.A(n_4086), .B(n_4044), .C(n_30063), .Z(n_223091119
		));
	notech_nand2 i_4172201(.A(n_2390), .B(n_1791), .Z(n_1604));
	notech_inv i_34962(.A(n_1614), .Z(\udeco[125] ));
	notech_inv i_34963(.A(n_1620), .Z(\udeco[123] ));
	notech_inv i_34964(.A(n_1628), .Z(\udeco[45] ));
	notech_inv i_34965(.A(n_1802), .Z(n_29919));
	notech_inv i_34966(.A(n_1639), .Z(\udeco[27] ));
	notech_inv i_34967(.A(n_2027), .Z(n_29921));
	notech_inv i_34968(.A(n_2359), .Z(n_29922));
	notech_inv i_34969(.A(n_2469), .Z(n_29923));
	notech_inv i_34970(.A(n_2149), .Z(n_29924));
	notech_inv i_34971(.A(n_57762), .Z(n_29925));
	notech_inv i_34972(.A(n_2059), .Z(n_29926));
	notech_inv i_34973(.A(n_2005), .Z(n_29927));
	notech_inv i_34974(.A(n_2098), .Z(n_29928));
	notech_inv i_34975(.A(n_2202), .Z(n_29929));
	notech_inv i_34976(.A(n_2078), .Z(n_29930));
	notech_inv i_34977(.A(n_2013), .Z(n_29931));
	notech_inv i_34978(.A(n_2020), .Z(\udeco[112] ));
	notech_inv i_34979(.A(n_2055), .Z(\udeco[109] ));
	notech_inv i_34980(.A(n_2092), .Z(\udeco[32] ));
	notech_inv i_34981(.A(n_2127), .Z(\udeco[24] ));
	notech_inv i_34982(.A(n_2135), .Z(\udeco[20] ));
	notech_inv i_34983(.A(n_2146), .Z(\udeco[18] ));
	notech_inv i_34984(.A(n_2177), .Z(\udeco[17] ));
	notech_inv i_34985(.A(n_2208), .Z(\udeco[13] ));
	notech_inv i_34986(.A(n_221989125), .Z(\udeco[11] ));
	notech_inv i_34987(.A(n_2227), .Z(\udeco[10] ));
	notech_inv i_34988(.A(n_2241), .Z(\udeco[9] ));
	notech_inv i_34989(.A(n_2270), .Z(\udeco[0] ));
	notech_inv i_34990(.A(n_4003), .Z(n_29944));
	notech_inv i_34991(.A(n_4080), .Z(n_29945));
	notech_inv i_34992(.A(n_3974), .Z(n_29946));
	notech_inv i_34993(.A(n_207949052), .Z(n_29947));
	notech_inv i_34994(.A(n_4018), .Z(n_29948));
	notech_inv i_34995(.A(n_4093), .Z(n_29949));
	notech_inv i_34996(.A(n_4062), .Z(n_29950));
	notech_inv i_34997(.A(n_4057), .Z(n_29951));
	notech_inv i_34998(.A(n_4052), .Z(n_29952));
	notech_inv i_34999(.A(n_4091), .Z(n_29953));
	notech_inv i_35000(.A(n_4054), .Z(n_29954));
	notech_inv i_35001(.A(n_4050), .Z(n_29955));
	notech_inv i_35002(.A(n_4065), .Z(n_29956));
	notech_inv i_35003(.A(n_3969), .Z(n_29957));
	notech_inv i_35004(.A(n_4060), .Z(n_29958));
	notech_inv i_35005(.A(n_4015), .Z(n_29959));
	notech_inv i_35006(.A(n_4059), .Z(n_29960));
	notech_inv i_35007(.A(n_4045), .Z(n_29961));
	notech_inv i_35008(.A(n_3971), .Z(n_29962));
	notech_inv i_35009(.A(n_3981), .Z(n_29963));
	notech_inv i_35010(.A(n_204849027), .Z(n_29964));
	notech_inv i_35011(.A(n_4033), .Z(n_29965));
	notech_inv i_35012(.A(n_3984), .Z(n_29966));
	notech_inv i_35013(.A(n_4082), .Z(n_29967));
	notech_inv i_35014(.A(n_3908), .Z(n_29968));
	notech_inv i_35015(.A(n_3846), .Z(n_29969));
	notech_inv i_35016(.A(n_4071), .Z(n_29970));
	notech_inv i_35017(.A(n_3760), .Z(n_29971));
	notech_inv i_35018(.A(n_4006), .Z(n_29972));
	notech_inv i_35019(.A(n_4011), .Z(n_29973));
	notech_inv i_35020(.A(n_3955), .Z(n_29974));
	notech_inv i_35021(.A(n_4009), .Z(n_29975));
	notech_inv i_35022(.A(n_3972), .Z(n_29976));
	notech_inv i_35023(.A(n_3820), .Z(n_29977));
	notech_inv i_35024(.A(n_3990), .Z(n_29978));
	notech_inv i_35025(.A(n_4023), .Z(n_29979));
	notech_inv i_35026(.A(n_4035), .Z(n_29980));
	notech_inv i_35027(.A(n_3728), .Z(n_29981));
	notech_inv i_35028(.A(n_3697), .Z(n_29982));
	notech_inv i_35029(.A(n_3980), .Z(n_29983));
	notech_inv i_35030(.A(n_2305), .Z(n_29984));
	notech_inv i_35031(.A(n_4001), .Z(n_29985));
	notech_inv i_35032(.A(n_3986), .Z(n_29986));
	notech_inv i_35033(.A(n_4088), .Z(n_29987));
	notech_inv i_35034(.A(n_3978), .Z(n_29988));
	notech_inv i_35035(.A(n_3950), .Z(n_29989));
	notech_inv i_35036(.A(n_3985), .Z(n_29990));
	notech_inv i_35037(.A(n_4089), .Z(n_29991));
	notech_inv i_35038(.A(n_3968), .Z(n_29992));
	notech_inv i_35039(.A(n_4085), .Z(n_29993));
	notech_inv i_35040(.A(n_2102), .Z(n_29994));
	notech_inv i_35041(.A(n_2354), .Z(n_29995));
	notech_inv i_35042(.A(n_1708), .Z(n_29996));
	notech_inv i_35043(.A(n_1709), .Z(n_29997));
	notech_inv i_35044(.A(n_122890278), .Z(n_29998));
	notech_inv i_35045(.A(n_125890305), .Z(n_29999));
	notech_inv i_35046(.A(n_126990312), .Z(n_30000));
	notech_inv i_35047(.A(n_1712), .Z(n_30001));
	notech_inv i_35048(.A(n_1870), .Z(n_30002));
	notech_inv i_35049(.A(n_127690319), .Z(n_30003));
	notech_inv i_35050(.A(n_2397), .Z(n_30004));
	notech_inv i_35051(.A(n_133490363), .Z(n_30005));
	notech_inv i_35052(.A(n_136890390), .Z(n_30006));
	notech_inv i_35053(.A(n_138990407), .Z(n_30007));
	notech_inv i_35054(.A(n_1953), .Z(n_30008));
	notech_inv i_35055(.A(n_121190261), .Z(n_30009));
	notech_inv i_35056(.A(n_143890451), .Z(n_30010));
	notech_inv i_35057(.A(n_146990479), .Z(n_30011));
	notech_inv i_35058(.A(n_2614), .Z(n_30012));
	notech_inv i_35059(.A(n_2878), .Z(n_30013));
	notech_inv i_35060(.A(n_1978), .Z(n_30014));
	notech_inv i_35061(.A(n_2854), .Z(n_30015));
	notech_inv i_35062(.A(n_1623), .Z(n_30016));
	notech_inv i_35063(.A(n_153490535), .Z(n_30017));
	notech_inv i_35064(.A(n_2304), .Z(n_30018));
	notech_inv i_35065(.A(n_155190547), .Z(n_30019));
	notech_inv i_35066(.A(n_1981), .Z(n_30020));
	notech_inv i_35067(.A(n_1933), .Z(n_30021));
	notech_inv i_35068(.A(n_1704), .Z(n_30022));
	notech_inv i_35069(.A(n_1951), .Z(n_30023));
	notech_inv i_35070(.A(n_162290606), .Z(n_30024));
	notech_inv i_35071(.A(n_2759), .Z(n_30025));
	notech_inv i_35072(.A(n_2754), .Z(n_30026));
	notech_inv i_35073(.A(n_1702), .Z(n_30027));
	notech_inv i_35074(.A(n_3107), .Z(n_30028));
	notech_inv i_35075(.A(n_2713), .Z(n_30029));
	notech_inv i_35076(.A(n_172190689), .Z(n_30030));
	notech_inv i_35077(.A(n_172490692), .Z(n_30031));
	notech_inv i_35078(.A(n_2678), .Z(n_30032));
	notech_inv i_35079(.A(n_3510), .Z(n_30033));
	notech_inv i_35080(.A(n_1718), .Z(n_30034));
	notech_inv i_35081(.A(n_1699), .Z(n_30035));
	notech_inv i_35082(.A(n_1263), .Z(n_30036));
	notech_inv i_35083(.A(n_2620), .Z(n_30037));
	notech_inv i_35084(.A(n_2615), .Z(n_30038));
	notech_inv i_35085(.A(n_185090794), .Z(n_30039));
	notech_inv i_35086(.A(n_696), .Z(n_30040));
	notech_inv i_35087(.A(n_2543), .Z(n_30041));
	notech_inv i_35088(.A(n_2541), .Z(n_30042));
	notech_inv i_35089(.A(n_2536), .Z(n_30043));
	notech_inv i_35090(.A(n_1615), .Z(n_30044));
	notech_inv i_35091(.A(n_2296), .Z(n_30045));
	notech_inv i_35092(.A(n_1923), .Z(n_30046));
	notech_inv i_35093(.A(n_2022), .Z(n_30047));
	notech_inv i_35094(.A(n_190090839), .Z(n_30048));
	notech_inv i_35095(.A(n_2426), .Z(n_30049));
	notech_inv i_35096(.A(n_1969), .Z(n_30050));
	notech_inv i_35097(.A(n_2369), .Z(n_30051));
	notech_inv i_35098(.A(n_190990847), .Z(n_30052));
	notech_inv i_35099(.A(n_3959), .Z(n_30053));
	notech_inv i_35100(.A(n_1942), .Z(n_30054));
	notech_inv i_35101(.A(n_2390), .Z(n_30055));
	notech_inv i_35102(.A(n_2401), .Z(n_30056));
	notech_inv i_35103(.A(n_2210), .Z(n_30057));
	notech_inv i_35104(.A(n_1987), .Z(n_30058));
	notech_inv i_35105(.A(n_2355), .Z(n_30059));
	notech_inv i_35106(.A(n_2466), .Z(n_30060));
	notech_inv i_35107(.A(n_2463), .Z(n_30061));
	notech_inv i_35108(.A(n_196590893), .Z(n_30062));
	notech_inv i_35109(.A(n_1249), .Z(n_30063));
	notech_inv i_35110(.A(n_1180), .Z(n_30064));
	notech_inv i_35111(.A(n_2431), .Z(n_30065));
	notech_inv i_35112(.A(n_2418), .Z(n_30066));
	notech_inv i_35113(.A(n_2287), .Z(n_30067));
	notech_inv i_35114(.A(n_1905), .Z(n_30068));
	notech_inv i_35115(.A(n_2391), .Z(n_30069));
	notech_inv i_35116(.A(n_201190930), .Z(n_30070));
	notech_inv i_35117(.A(n_2852), .Z(n_30071));
	notech_inv i_35118(.A(n_2324), .Z(n_30072));
	notech_inv i_35119(.A(n_2321), .Z(n_30073));
	notech_inv i_35120(.A(n_2656), .Z(n_30074));
	notech_inv i_35121(.A(n_2850), .Z(n_30075));
	notech_inv i_35122(.A(n_208390990), .Z(n_30076));
	notech_inv i_35123(.A(n_208990996), .Z(n_30077));
	notech_inv i_35124(.A(n_2186), .Z(n_30078));
	notech_inv i_35125(.A(n_2792), .Z(n_30079));
	notech_inv i_35126(.A(n_1999), .Z(n_30080));
	notech_inv i_35127(.A(n_1972), .Z(n_30081));
	notech_inv i_35128(.A(n_210091005), .Z(n_30082));
	notech_inv i_35129(.A(n_2038), .Z(n_30083));
	notech_inv i_35130(.A(n_1816), .Z(n_30084));
	notech_inv i_35131(.A(n_2006), .Z(n_30085));
	notech_inv i_35132(.A(n_1986), .Z(n_30086));
	notech_inv i_35133(.A(n_1965), .Z(n_30087));
	notech_inv i_35134(.A(n_1624), .Z(n_30088));
	notech_inv i_35135(.A(n_2036), .Z(n_30089));
	notech_inv i_35136(.A(n_1943), .Z(n_30090));
	notech_inv i_35137(.A(n_1114), .Z(n_30091));
	notech_inv i_35138(.A(n_1841), .Z(n_30092));
	notech_inv i_35139(.A(n_1840), .Z(n_30093));
	notech_inv i_35140(.A(n_2116), .Z(n_30094));
	notech_inv i_35141(.A(n_214991049), .Z(n_30095));
	notech_inv i_35142(.A(n_2017), .Z(n_30096));
	notech_inv i_35143(.A(n_960), .Z(n_30097));
	notech_inv i_35144(.A(n_1695), .Z(n_30098));
	notech_inv i_35145(.A(n_2365), .Z(n_30099));
	notech_inv i_35146(.A(n_221891108), .Z(n_30100));
	notech_inv i_35147(.A(n_2357), .Z(n_30101));
	notech_inv i_35148(.A(n_222491113), .Z(n_30102));
	notech_inv i_35149(.A(n_2380), .Z(\udeco[5] ));
	notech_inv i_35150(.A(n_223091119), .Z(n_30104));
	notech_inv i_35151(.A(n_1950), .Z(n_30105));
	notech_inv i_35153(.A(n_57816), .Z(n_30107));
	notech_inv i_35154(.A(n_57845), .Z(n_30108));
	notech_inv i_35156(.A(n_57868), .Z(n_30110));
	notech_inv i_35157(.A(n_57854), .Z(n_30111));
	notech_inv i_35158(.A(op[7]), .Z(n_30112));
	notech_inv i_35159(.A(modrm[0]), .Z(n_30113));
	notech_inv i_35160(.A(modrm[1]), .Z(n_30114));
	notech_inv i_35161(.A(modrm[3]), .Z(n_30115));
	notech_inv i_35162(.A(modrm[4]), .Z(n_30116));
	notech_inv i_35163(.A(n_57726), .Z(n_30117));
	notech_inv i_35164(.A(modrm[6]), .Z(n_30118));
	notech_inv i_35165(.A(ipg_fault), .Z(n_30119));
	notech_inv i_35166(.A(twobyte), .Z(n_30120));
	notech_inv i_35167(.A(adz), .Z(n_30121));
	notech_inv i_35168(.A(n_4024), .Z(n_30122));
	notech_inv i_35169(.A(n_1622), .Z(n_30123));
	notech_inv i_35170(.A(n_1608), .Z(n_30124));
	notech_inv i_35171(.A(\udeco[91] ), .Z(n_30125));
	notech_inv i_35172(.A(udeco_7397047), .Z(\udeco[73] ));
	notech_inv i_35173(.A(udeco_10197046), .Z(\udeco[101] ));
	notech_inv i_35174(.A(udeco_10397045), .Z(\udeco[103] ));
	notech_inv i_35175(.A(udeco_3597044), .Z(\udeco[35] ));
	notech_inv i_35176(.A(udeco_2997043), .Z(\udeco[29] ));
	notech_inv i_35177(.A(udeco_2897042), .Z(\udeco[28] ));
	notech_inv i_35178(.A(udeco_2197041), .Z(\udeco[21] ));
	notech_inv i_35179(.A(udeco_1597040), .Z(\udeco[15] ));
	notech_inv i_35180(.A(udeco_1497039), .Z(\udeco[14] ));
	notech_inv i_35181(.A(udeco_1297038), .Z(\udeco[12] ));
	notech_inv i_35182(.A(udeco_11997037), .Z(\udeco[119] ));
	notech_inv i_35183(.A(udeco_11497036), .Z(\udeco[114] ));
	notech_inv i_35184(.A(udeco_11397035), .Z(\udeco[113] ));
	notech_inv i_35185(.A(udeco_3797034), .Z(\udeco[37] ));
	notech_inv i_35186(.A(udeco_2397033), .Z(\udeco[23] ));
	notech_inv i_35187(.A(n_1607), .Z(n_30141));
endmodule
module deco(clk, rstn, useq_ptr, in128, adz, pc_req, ivect, int_main, iack, ie, pg_fault
		, ipg_fault, cpl, cr0, valid_len, to_vliw, lenpc_out, immediate,
		 to_acu, operand_size, reps, over_seg, valid_op, term, start, ready_vliw
		);

	input clk;
	input rstn;
	output [3:0] useq_ptr;
	input [127:0] in128;
	input adz;
	input pc_req;
	input [7:0] ivect;
	input int_main;
	output iack;
	input ie;
	input pg_fault;
	input ipg_fault;
	input [1:0] cpl;
	input [31:0] cr0;
	input [5:0] valid_len;
	output [127:0] to_vliw;
	output [31:0] lenpc_out;
	output [63:0] immediate;
	output [210:0] to_acu;
	output [2:0] operand_size;
	output [2:0] reps;
	output [5:0] over_seg;
	output valid_op;
	input term;
	output start;
	input ready_vliw;

	wire [210:0] to_acu2;
	wire [2:0] opz2;
	wire [31:0] lenpc2;
	wire [210:0] to_acu1;
	wire [127:0] inst_deco1;
	wire [127:0] inst_deco2;
	wire [2:0] reps1;
	wire [3:0] i_ptr;
	wire [5:0] int_excl;
	wire [1:0] idx_deco;
	wire [2:0] reps2;
	wire [7:0] ififo_rvect1;
	wire [4:0] fsm;
	wire [31:0] lenpc1;
	wire [2:0] opz1;
	wire [210:0] to_acu0;
	wire [127:0] inst_deco;
	wire [2:0] opz0;
	wire [2:0] reps0;
	wire [31:0] lenpc;
	wire [7:0] ififo_rvect2;
	wire [7:0] ififo_rvect3;
	wire [7:0] ififo_rvect4;
	wire [127:0] udeco;
	wire [2:0] displc;
	wire [2:0] opz;
	wire [2:0] imm_sz;
	wire [4:0] pfx_sz;



	notech_inv i_15638(.A(n_61909), .Z(n_61972));
	notech_inv i_15636(.A(n_61909), .Z(n_61970));
	notech_inv i_15633(.A(n_61909), .Z(n_61967));
	notech_inv i_15631(.A(n_61909), .Z(n_61965));
	notech_inv i_15628(.A(n_61909), .Z(n_61962));
	notech_inv i_15626(.A(n_61909), .Z(n_61960));
	notech_inv i_15622(.A(n_61909), .Z(n_61956));
	notech_inv i_15620(.A(n_61909), .Z(n_61954));
	notech_inv i_15617(.A(n_61909), .Z(n_61951));
	notech_inv i_15615(.A(n_61909), .Z(n_61949));
	notech_inv i_15612(.A(n_61909), .Z(n_61946));
	notech_inv i_15610(.A(n_61909), .Z(n_61944));
	notech_inv i_15606(.A(n_61909), .Z(n_61940));
	notech_inv i_15604(.A(n_61909), .Z(n_61938));
	notech_inv i_15601(.A(n_61909), .Z(n_61935));
	notech_inv i_15599(.A(n_61909), .Z(n_61933));
	notech_inv i_15596(.A(n_61909), .Z(n_61930));
	notech_inv i_15594(.A(n_61909), .Z(n_61928));
	notech_inv i_15590(.A(n_61911), .Z(n_61924));
	notech_inv i_15588(.A(n_61911), .Z(n_61922));
	notech_inv i_15585(.A(n_61911), .Z(n_61919));
	notech_inv i_15583(.A(n_61911), .Z(n_61917));
	notech_inv i_15580(.A(n_61911), .Z(n_61914));
	notech_inv i_15578(.A(n_61911), .Z(n_61912));
	notech_inv i_15577(.A(n_61910), .Z(n_61911));
	notech_inv i_15576(.A(n_61909), .Z(n_61910));
	notech_inv i_15575(.A(clk), .Z(n_61909));
	notech_inv i_15573(.A(n_61844), .Z(n_61907));
	notech_inv i_15571(.A(n_61844), .Z(n_61905));
	notech_inv i_15568(.A(n_61844), .Z(n_61902));
	notech_inv i_15566(.A(n_61844), .Z(n_61900));
	notech_inv i_15563(.A(n_61844), .Z(n_61897));
	notech_inv i_15561(.A(n_61844), .Z(n_61895));
	notech_inv i_15557(.A(n_61844), .Z(n_61891));
	notech_inv i_15555(.A(n_61844), .Z(n_61889));
	notech_inv i_15552(.A(n_61844), .Z(n_61886));
	notech_inv i_15550(.A(n_61844), .Z(n_61884));
	notech_inv i_15547(.A(n_61844), .Z(n_61881));
	notech_inv i_15545(.A(n_61844), .Z(n_61879));
	notech_inv i_15541(.A(n_61844), .Z(n_61875));
	notech_inv i_15539(.A(n_61844), .Z(n_61873));
	notech_inv i_15536(.A(n_61844), .Z(n_61870));
	notech_inv i_15534(.A(n_61844), .Z(n_61868));
	notech_inv i_15531(.A(n_61844), .Z(n_61865));
	notech_inv i_15529(.A(n_61844), .Z(n_61863));
	notech_inv i_15525(.A(n_61846), .Z(n_61859));
	notech_inv i_15523(.A(n_61846), .Z(n_61857));
	notech_inv i_15520(.A(n_61846), .Z(n_61854));
	notech_inv i_15518(.A(n_61846), .Z(n_61852));
	notech_inv i_15515(.A(n_61846), .Z(n_61849));
	notech_inv i_15513(.A(n_61846), .Z(n_61847));
	notech_inv i_15512(.A(n_61868), .Z(n_61846));
	notech_inv i_15510(.A(clk), .Z(n_61844));
	notech_inv i_15508(.A(n_61779), .Z(n_61842));
	notech_inv i_15506(.A(n_61779), .Z(n_61840));
	notech_inv i_15503(.A(n_61779), .Z(n_61837));
	notech_inv i_15501(.A(n_61779), .Z(n_61835));
	notech_inv i_15498(.A(n_61779), .Z(n_61832));
	notech_inv i_15496(.A(n_61779), .Z(n_61830));
	notech_inv i_15492(.A(n_61779), .Z(n_61826));
	notech_inv i_15490(.A(n_61779), .Z(n_61824));
	notech_inv i_15487(.A(n_61779), .Z(n_61821));
	notech_inv i_15485(.A(n_61779), .Z(n_61819));
	notech_inv i_15482(.A(n_61779), .Z(n_61816));
	notech_inv i_15480(.A(n_61779), .Z(n_61814));
	notech_inv i_15476(.A(n_61779), .Z(n_61810));
	notech_inv i_15474(.A(n_61779), .Z(n_61808));
	notech_inv i_15471(.A(n_61779), .Z(n_61805));
	notech_inv i_15469(.A(n_61779), .Z(n_61803));
	notech_inv i_15466(.A(n_61779), .Z(n_61800));
	notech_inv i_15464(.A(n_61779), .Z(n_61798));
	notech_inv i_15460(.A(n_61781), .Z(n_61794));
	notech_inv i_15458(.A(n_61781), .Z(n_61792));
	notech_inv i_15455(.A(n_61781), .Z(n_61789));
	notech_inv i_15453(.A(n_61781), .Z(n_61787));
	notech_inv i_15450(.A(n_61781), .Z(n_61784));
	notech_inv i_15448(.A(n_61781), .Z(n_61782));
	notech_inv i_15447(.A(n_61803), .Z(n_61781));
	notech_inv i_15445(.A(clk), .Z(n_61779));
	notech_inv i_14767(.A(n_61348), .Z(n_61412));
	notech_inv i_14765(.A(n_61348), .Z(n_61410));
	notech_inv i_14764(.A(n_61348), .Z(n_61409));
	notech_inv i_14760(.A(n_61348), .Z(n_61405));
	notech_inv i_14759(.A(n_61348), .Z(n_61404));
	notech_inv i_14755(.A(n_61348), .Z(n_61400));
	notech_inv i_14754(.A(n_61348), .Z(n_61399));
	notech_inv i_14750(.A(n_61348), .Z(n_61395));
	notech_inv i_14748(.A(n_61348), .Z(n_61393));
	notech_inv i_14745(.A(n_61348), .Z(n_61390));
	notech_inv i_14743(.A(n_61348), .Z(n_61388));
	notech_inv i_14740(.A(n_61348), .Z(n_61385));
	notech_inv i_14738(.A(n_61348), .Z(n_61383));
	notech_inv i_14734(.A(n_61348), .Z(n_61379));
	notech_inv i_14732(.A(n_61348), .Z(n_61377));
	notech_inv i_14729(.A(n_61348), .Z(n_61374));
	notech_inv i_14727(.A(n_61348), .Z(n_61372));
	notech_inv i_14724(.A(n_61348), .Z(n_61369));
	notech_inv i_14722(.A(n_61348), .Z(n_61367));
	notech_inv i_14718(.A(n_61350), .Z(n_61363));
	notech_inv i_14716(.A(n_61350), .Z(n_61361));
	notech_inv i_14713(.A(n_61350), .Z(n_61358));
	notech_inv i_14711(.A(n_61350), .Z(n_61356));
	notech_inv i_14708(.A(n_61350), .Z(n_61353));
	notech_inv i_14706(.A(n_61350), .Z(n_61351));
	notech_inv i_14705(.A(n_61367), .Z(n_61350));
	notech_inv i_14703(.A(rstn), .Z(n_61348));
	notech_inv i_14701(.A(n_61283), .Z(n_61346));
	notech_inv i_14699(.A(n_61283), .Z(n_61344));
	notech_inv i_14696(.A(n_61283), .Z(n_61341));
	notech_inv i_14694(.A(n_61283), .Z(n_61339));
	notech_inv i_14691(.A(n_61283), .Z(n_61336));
	notech_inv i_14689(.A(n_61283), .Z(n_61334));
	notech_inv i_14685(.A(n_61283), .Z(n_61330));
	notech_inv i_14683(.A(n_61283), .Z(n_61328));
	notech_inv i_14680(.A(n_61283), .Z(n_61325));
	notech_inv i_14678(.A(n_61283), .Z(n_61323));
	notech_inv i_14675(.A(n_61283), .Z(n_61320));
	notech_inv i_14673(.A(n_61283), .Z(n_61318));
	notech_inv i_14669(.A(n_61283), .Z(n_61314));
	notech_inv i_14667(.A(n_61283), .Z(n_61312));
	notech_inv i_14664(.A(n_61283), .Z(n_61309));
	notech_inv i_14662(.A(n_61283), .Z(n_61307));
	notech_inv i_14659(.A(n_61283), .Z(n_61304));
	notech_inv i_14657(.A(n_61283), .Z(n_61302));
	notech_inv i_14653(.A(n_61285), .Z(n_61298));
	notech_inv i_14651(.A(n_61285), .Z(n_61296));
	notech_inv i_14648(.A(n_61285), .Z(n_61293));
	notech_inv i_14646(.A(n_61285), .Z(n_61291));
	notech_inv i_14643(.A(n_61285), .Z(n_61288));
	notech_inv i_14641(.A(n_61285), .Z(n_61286));
	notech_inv i_14640(.A(n_61307), .Z(n_61285));
	notech_inv i_14638(.A(rstn), .Z(n_61283));
	notech_inv i_14636(.A(n_61218), .Z(n_61281));
	notech_inv i_14634(.A(n_61218), .Z(n_61279));
	notech_inv i_14631(.A(n_61218), .Z(n_61276));
	notech_inv i_14629(.A(n_61218), .Z(n_61274));
	notech_inv i_14626(.A(n_61218), .Z(n_61271));
	notech_inv i_14624(.A(n_61218), .Z(n_61269));
	notech_inv i_14620(.A(n_61218), .Z(n_61265));
	notech_inv i_14618(.A(n_61218), .Z(n_61263));
	notech_inv i_14615(.A(n_61218), .Z(n_61260));
	notech_inv i_14613(.A(n_61218), .Z(n_61258));
	notech_inv i_14610(.A(n_61218), .Z(n_61255));
	notech_inv i_14608(.A(n_61218), .Z(n_61253));
	notech_inv i_14604(.A(n_61218), .Z(n_61249));
	notech_inv i_14602(.A(n_61218), .Z(n_61247));
	notech_inv i_14599(.A(n_61218), .Z(n_61244));
	notech_inv i_14597(.A(n_61218), .Z(n_61242));
	notech_inv i_14594(.A(n_61218), .Z(n_61239));
	notech_inv i_14592(.A(n_61218), .Z(n_61237));
	notech_inv i_14588(.A(n_61220), .Z(n_61233));
	notech_inv i_14586(.A(n_61220), .Z(n_61231));
	notech_inv i_14583(.A(n_61220), .Z(n_61228));
	notech_inv i_14581(.A(n_61220), .Z(n_61226));
	notech_inv i_14578(.A(n_61220), .Z(n_61223));
	notech_inv i_14576(.A(n_61220), .Z(n_61221));
	notech_inv i_14575(.A(n_61242), .Z(n_61220));
	notech_inv i_14573(.A(rstn), .Z(n_61218));
	notech_inv i_14088(.A(n_60649), .Z(n_60714));
	notech_inv i_14087(.A(n_60649), .Z(n_60713));
	notech_inv i_14082(.A(n_60649), .Z(n_60708));
	notech_inv i_14077(.A(n_60649), .Z(n_60703));
	notech_inv i_14076(.A(n_60649), .Z(n_60702));
	notech_inv i_14071(.A(n_60649), .Z(n_60697));
	notech_inv i_14066(.A(n_60649), .Z(n_60692));
	notech_inv i_14065(.A(n_60649), .Z(n_60691));
	notech_inv i_14060(.A(n_60649), .Z(n_60686));
	notech_inv i_14054(.A(n_60649), .Z(n_60680));
	notech_inv i_14053(.A(n_60649), .Z(n_60679));
	notech_inv i_14048(.A(n_60649), .Z(n_60674));
	notech_inv i_14043(.A(n_60649), .Z(n_60669));
	notech_inv i_14042(.A(n_60649), .Z(n_60668));
	notech_inv i_14037(.A(n_60649), .Z(n_60663));
	notech_inv i_14032(.A(n_60649), .Z(n_60658));
	notech_inv i_14031(.A(n_60649), .Z(n_60657));
	notech_inv i_14026(.A(n_60649), .Z(n_60652));
	notech_inv i_14023(.A(term), .Z(n_60649));
	notech_inv i_14020(.A(n_60615), .Z(n_60646));
	notech_inv i_14019(.A(n_60615), .Z(n_60645));
	notech_inv i_14014(.A(n_60615), .Z(n_60640));
	notech_inv i_14009(.A(n_60615), .Z(n_60635));
	notech_inv i_14008(.A(n_60615), .Z(n_60634));
	notech_inv i_14003(.A(n_60615), .Z(n_60629));
	notech_inv i_13998(.A(n_60615), .Z(n_60624));
	notech_inv i_13997(.A(n_60615), .Z(n_60623));
	notech_inv i_13992(.A(n_60615), .Z(n_60618));
	notech_inv i_13989(.A(term), .Z(n_60615));
	notech_inv i_13182(.A(n_59679), .Z(n_59695));
	notech_inv i_13180(.A(n_59679), .Z(n_59693));
	notech_inv i_13179(.A(n_59679), .Z(n_59692));
	notech_inv i_13175(.A(n_59679), .Z(n_59688));
	notech_inv i_13173(.A(n_59679), .Z(n_59686));
	notech_inv i_13170(.A(n_59679), .Z(n_59683));
	notech_inv i_13168(.A(n_59679), .Z(n_59681));
	notech_inv i_13167(.A(n_59679), .Z(n_59680));
	notech_inv i_13166(.A(n_2055), .Z(n_59679));
	notech_inv i_13157(.A(n_59668), .Z(n_59669));
	notech_inv i_13156(.A(n_2124), .Z(n_59668));
	notech_inv i_13153(.A(n_59599), .Z(n_59664));
	notech_inv i_13152(.A(n_59599), .Z(n_59663));
	notech_inv i_13147(.A(n_59599), .Z(n_59658));
	notech_inv i_13142(.A(n_59599), .Z(n_59653));
	notech_inv i_13141(.A(n_59599), .Z(n_59652));
	notech_inv i_13136(.A(n_59599), .Z(n_59647));
	notech_inv i_13131(.A(n_59599), .Z(n_59642));
	notech_inv i_13130(.A(n_59599), .Z(n_59641));
	notech_inv i_13125(.A(n_59599), .Z(n_59636));
	notech_inv i_13119(.A(n_59599), .Z(n_59630));
	notech_inv i_13118(.A(n_59599), .Z(n_59629));
	notech_inv i_13113(.A(n_59599), .Z(n_59624));
	notech_inv i_13108(.A(n_59599), .Z(n_59619));
	notech_inv i_13107(.A(n_59599), .Z(n_59618));
	notech_inv i_13102(.A(n_59599), .Z(n_59613));
	notech_inv i_13097(.A(n_59599), .Z(n_59608));
	notech_inv i_13096(.A(n_59599), .Z(n_59607));
	notech_inv i_13091(.A(n_59599), .Z(n_59602));
	notech_inv i_13088(.A(n_40195), .Z(n_59599));
	notech_inv i_13085(.A(n_59565), .Z(n_59596));
	notech_inv i_13084(.A(n_59565), .Z(n_59595));
	notech_inv i_13079(.A(n_59565), .Z(n_59590));
	notech_inv i_13073(.A(n_59565), .Z(n_59584));
	notech_inv i_13068(.A(n_59565), .Z(n_59579));
	notech_inv i_13062(.A(n_59565), .Z(n_59573));
	notech_inv i_13057(.A(n_59565), .Z(n_59568));
	notech_inv i_13054(.A(n_40195), .Z(n_59565));
	notech_inv i_12369(.A(n_58828), .Z(n_58882));
	notech_inv i_12368(.A(n_58828), .Z(n_58881));
	notech_inv i_12364(.A(n_58828), .Z(n_58877));
	notech_inv i_12360(.A(n_58828), .Z(n_58873));
	notech_inv i_12359(.A(n_58828), .Z(n_58872));
	notech_inv i_12355(.A(n_58828), .Z(n_58868));
	notech_inv i_12351(.A(n_58828), .Z(n_58864));
	notech_inv i_12350(.A(n_58828), .Z(n_58863));
	notech_inv i_12346(.A(n_58828), .Z(n_58859));
	notech_inv i_12341(.A(n_58828), .Z(n_58854));
	notech_inv i_12340(.A(n_58828), .Z(n_58853));
	notech_inv i_12336(.A(n_58828), .Z(n_58849));
	notech_inv i_12332(.A(n_58828), .Z(n_58845));
	notech_inv i_12331(.A(n_58828), .Z(n_58844));
	notech_inv i_12327(.A(n_58828), .Z(n_58840));
	notech_inv i_12323(.A(n_58828), .Z(n_58836));
	notech_inv i_12322(.A(n_58828), .Z(n_58835));
	notech_inv i_12318(.A(n_58828), .Z(n_58831));
	notech_inv i_12315(.A(n_2828), .Z(n_58828));
	notech_inv i_12313(.A(n_58800), .Z(n_58826));
	notech_inv i_12312(.A(n_58800), .Z(n_58825));
	notech_inv i_12308(.A(n_58800), .Z(n_58821));
	notech_inv i_12299(.A(n_58811), .Z(n_58812));
	notech_inv i_12298(.A(n_58810), .Z(n_58811));
	notech_inv i_12297(.A(n_58800), .Z(n_58810));
	notech_inv i_12290(.A(n_58802), .Z(n_58803));
	notech_inv i_12289(.A(n_58801), .Z(n_58802));
	notech_inv i_12288(.A(n_58800), .Z(n_58801));
	notech_inv i_12287(.A(n_2828), .Z(n_58800));
	notech_inv i_12285(.A(n_58709), .Z(n_58797));
	notech_inv i_12283(.A(n_58709), .Z(n_58795));
	notech_inv i_12280(.A(n_58709), .Z(n_58792));
	notech_inv i_12278(.A(n_58709), .Z(n_58790));
	notech_inv i_12274(.A(n_58709), .Z(n_58786));
	notech_inv i_12272(.A(n_58709), .Z(n_58784));
	notech_inv i_12269(.A(n_58709), .Z(n_58781));
	notech_inv i_12267(.A(n_58709), .Z(n_58779));
	notech_inv i_12263(.A(n_58709), .Z(n_58775));
	notech_inv i_12261(.A(n_58709), .Z(n_58773));
	notech_inv i_12258(.A(n_58709), .Z(n_58770));
	notech_inv i_12256(.A(n_58709), .Z(n_58768));
	notech_inv i_12252(.A(n_58709), .Z(n_58764));
	notech_inv i_12250(.A(n_58709), .Z(n_58762));
	notech_inv i_12247(.A(n_58709), .Z(n_58759));
	notech_inv i_12245(.A(n_58709), .Z(n_58757));
	notech_inv i_12240(.A(n_58744), .Z(n_58752));
	notech_inv i_12238(.A(n_58744), .Z(n_58750));
	notech_inv i_12235(.A(n_58744), .Z(n_58747));
	notech_inv i_12233(.A(n_58744), .Z(n_58745));
	notech_inv i_12232(.A(n_58790), .Z(n_58744));
	notech_inv i_12229(.A(n_58744), .Z(n_58741));
	notech_inv i_12227(.A(n_58744), .Z(n_58739));
	notech_inv i_12224(.A(n_58744), .Z(n_58736));
	notech_inv i_12222(.A(n_58744), .Z(n_58734));
	notech_inv i_12218(.A(n_58744), .Z(n_58730));
	notech_inv i_12216(.A(n_58744), .Z(n_58728));
	notech_inv i_12213(.A(n_58744), .Z(n_58725));
	notech_inv i_12211(.A(n_58744), .Z(n_58723));
	notech_inv i_12207(.A(n_58709), .Z(n_58719));
	notech_inv i_12205(.A(n_58709), .Z(n_58717));
	notech_inv i_12202(.A(n_58709), .Z(n_58714));
	notech_inv i_12200(.A(n_58709), .Z(n_58712));
	notech_inv i_12197(.A(n_2829), .Z(n_58709));
	notech_inv i_12195(.A(n_58664), .Z(n_58707));
	notech_inv i_12193(.A(n_58664), .Z(n_58705));
	notech_inv i_12190(.A(n_58664), .Z(n_58702));
	notech_inv i_12188(.A(n_58664), .Z(n_58700));
	notech_inv i_12184(.A(n_58664), .Z(n_58696));
	notech_inv i_12182(.A(n_58664), .Z(n_58694));
	notech_inv i_12179(.A(n_58664), .Z(n_58691));
	notech_inv i_12177(.A(n_58664), .Z(n_58689));
	notech_inv i_12173(.A(n_58664), .Z(n_58685));
	notech_inv i_12171(.A(n_58664), .Z(n_58683));
	notech_inv i_12168(.A(n_58664), .Z(n_58680));
	notech_inv i_12166(.A(n_58664), .Z(n_58678));
	notech_inv i_12161(.A(n_58664), .Z(n_58673));
	notech_inv i_12160(.A(n_58664), .Z(n_58672));
	notech_inv i_12155(.A(n_58664), .Z(n_58667));
	notech_inv i_12152(.A(n_2829), .Z(n_58664));
	notech_inv i_11970(.A(n_58463), .Z(n_58479));
	notech_inv i_11968(.A(n_58463), .Z(n_58477));
	notech_inv i_11967(.A(n_58463), .Z(n_58476));
	notech_inv i_11963(.A(n_58463), .Z(n_58472));
	notech_inv i_11961(.A(n_58463), .Z(n_58470));
	notech_inv i_11958(.A(n_58463), .Z(n_58467));
	notech_inv i_11956(.A(n_58463), .Z(n_58465));
	notech_inv i_11955(.A(n_58463), .Z(n_58464));
	notech_inv i_11954(.A(n_5768), .Z(n_58463));
	notech_inv i_11947(.A(n_58454), .Z(n_58455));
	notech_inv i_11946(.A(n_3146), .Z(n_58454));
	notech_inv i_11944(.A(n_58433), .Z(n_58451));
	notech_inv i_11942(.A(n_58433), .Z(n_58449));
	notech_inv i_11939(.A(n_58433), .Z(n_58446));
	notech_inv i_11937(.A(n_58433), .Z(n_58444));
	notech_inv i_11934(.A(n_58433), .Z(n_58441));
	notech_inv i_11932(.A(n_58433), .Z(n_58439));
	notech_inv i_11929(.A(n_58433), .Z(n_58436));
	notech_inv i_11927(.A(n_58433), .Z(n_58434));
	notech_inv i_11926(.A(n_3145), .Z(n_58433));
	notech_inv i_11919(.A(n_58424), .Z(n_58425));
	notech_inv i_11918(.A(n_3246), .Z(n_58424));
	notech_inv i_11911(.A(n_58415), .Z(n_58416));
	notech_inv i_11910(.A(n_21291841), .Z(n_58415));
	notech_inv i_11903(.A(n_58406), .Z(n_58407));
	notech_inv i_11902(.A(n_38330), .Z(n_58406));
	notech_inv i_11900(.A(n_58387), .Z(n_58403));
	notech_inv i_11898(.A(n_58387), .Z(n_58401));
	notech_inv i_11897(.A(n_58387), .Z(n_58400));
	notech_inv i_11893(.A(n_58387), .Z(n_58396));
	notech_inv i_11891(.A(n_58387), .Z(n_58394));
	notech_inv i_11888(.A(n_58387), .Z(n_58391));
	notech_inv i_11886(.A(n_58387), .Z(n_58389));
	notech_inv i_11885(.A(n_58387), .Z(n_58388));
	notech_inv i_11884(.A(n_5276), .Z(n_58387));
	notech_inv i_11263(.A(n_57711), .Z(n_57713));
	notech_inv i_11262(.A(n_57711), .Z(n_57712));
	notech_inv i_11261(.A(in128[10]), .Z(n_57711));
	notech_inv i_11242(.A(n_57624), .Z(n_57689));
	notech_inv i_11241(.A(n_57624), .Z(n_57688));
	notech_inv i_11236(.A(n_57624), .Z(n_57683));
	notech_inv i_11231(.A(n_57624), .Z(n_57678));
	notech_inv i_11230(.A(n_57624), .Z(n_57677));
	notech_inv i_11225(.A(n_57624), .Z(n_57672));
	notech_inv i_11220(.A(n_57624), .Z(n_57667));
	notech_inv i_11219(.A(n_57624), .Z(n_57666));
	notech_inv i_11214(.A(n_57624), .Z(n_57661));
	notech_inv i_11208(.A(n_57624), .Z(n_57655));
	notech_inv i_11207(.A(n_57624), .Z(n_57654));
	notech_inv i_11202(.A(n_57624), .Z(n_57649));
	notech_inv i_11197(.A(n_57624), .Z(n_57644));
	notech_inv i_11196(.A(n_57624), .Z(n_57643));
	notech_inv i_11191(.A(n_57624), .Z(n_57638));
	notech_inv i_11186(.A(n_57624), .Z(n_57633));
	notech_inv i_11185(.A(n_57624), .Z(n_57632));
	notech_inv i_11180(.A(n_57624), .Z(n_57627));
	notech_inv i_11177(.A(\nbus_13549[0] ), .Z(n_57624));
	notech_inv i_11174(.A(n_57590), .Z(n_57621));
	notech_inv i_11173(.A(n_57590), .Z(n_57620));
	notech_inv i_11163(.A(n_57590), .Z(n_57610));
	notech_inv i_11162(.A(n_57590), .Z(n_57609));
	notech_inv i_11157(.A(n_57590), .Z(n_57604));
	notech_inv i_11152(.A(n_57590), .Z(n_57599));
	notech_inv i_11151(.A(n_57590), .Z(n_57598));
	notech_inv i_11146(.A(n_57590), .Z(n_57593));
	notech_inv i_11143(.A(\nbus_13549[0] ), .Z(n_57590));
	notech_inv i_11141(.A(n_57499), .Z(n_57587));
	notech_inv i_11139(.A(n_57499), .Z(n_57585));
	notech_inv i_11136(.A(n_57499), .Z(n_57582));
	notech_inv i_11134(.A(n_57499), .Z(n_57580));
	notech_inv i_11130(.A(n_57499), .Z(n_57576));
	notech_inv i_11128(.A(n_57499), .Z(n_57574));
	notech_inv i_11125(.A(n_57499), .Z(n_57571));
	notech_inv i_11123(.A(n_57499), .Z(n_57569));
	notech_inv i_11119(.A(n_57499), .Z(n_57565));
	notech_inv i_11117(.A(n_57499), .Z(n_57563));
	notech_inv i_11114(.A(n_57499), .Z(n_57560));
	notech_inv i_11112(.A(n_57499), .Z(n_57558));
	notech_inv i_11108(.A(n_57499), .Z(n_57554));
	notech_inv i_11106(.A(n_57499), .Z(n_57552));
	notech_inv i_11103(.A(n_57499), .Z(n_57549));
	notech_inv i_11101(.A(n_57499), .Z(n_57547));
	notech_inv i_11096(.A(n_57534), .Z(n_57542));
	notech_inv i_11094(.A(n_57534), .Z(n_57540));
	notech_inv i_11091(.A(n_57534), .Z(n_57537));
	notech_inv i_11089(.A(n_57534), .Z(n_57535));
	notech_inv i_11088(.A(n_57580), .Z(n_57534));
	notech_inv i_11085(.A(n_57534), .Z(n_57531));
	notech_inv i_11083(.A(n_57534), .Z(n_57529));
	notech_inv i_11080(.A(n_57534), .Z(n_57526));
	notech_inv i_11078(.A(n_57534), .Z(n_57524));
	notech_inv i_11074(.A(n_57534), .Z(n_57520));
	notech_inv i_11072(.A(n_57534), .Z(n_57518));
	notech_inv i_11069(.A(n_57534), .Z(n_57515));
	notech_inv i_11067(.A(n_57534), .Z(n_57513));
	notech_inv i_11063(.A(n_57499), .Z(n_57509));
	notech_inv i_11061(.A(n_57499), .Z(n_57507));
	notech_inv i_11058(.A(n_57499), .Z(n_57504));
	notech_inv i_11056(.A(n_57499), .Z(n_57502));
	notech_inv i_11053(.A(n_5409), .Z(n_57499));
	notech_inv i_11051(.A(n_57454), .Z(n_57497));
	notech_inv i_11049(.A(n_57454), .Z(n_57495));
	notech_inv i_11046(.A(n_57454), .Z(n_57492));
	notech_inv i_11044(.A(n_57454), .Z(n_57490));
	notech_inv i_11040(.A(n_57454), .Z(n_57486));
	notech_inv i_11038(.A(n_57454), .Z(n_57484));
	notech_inv i_11035(.A(n_57454), .Z(n_57481));
	notech_inv i_11033(.A(n_57454), .Z(n_57479));
	notech_inv i_11029(.A(n_57454), .Z(n_57475));
	notech_inv i_11027(.A(n_57454), .Z(n_57473));
	notech_inv i_11023(.A(n_57454), .Z(n_57469));
	notech_inv i_11017(.A(n_57454), .Z(n_57463));
	notech_inv i_11016(.A(n_57454), .Z(n_57462));
	notech_inv i_11011(.A(n_57454), .Z(n_57457));
	notech_inv i_11008(.A(n_5409), .Z(n_57454));
	notech_inv i_10332(.A(n_56588), .Z(n_56589));
	notech_inv i_10331(.A(n_2849), .Z(n_56588));
	notech_inv i_9038(.A(n_55059), .Z(n_55060));
	notech_inv i_9037(.A(n_162893249), .Z(n_55059));
	notech_inv i_9028(.A(n_55048), .Z(n_55049));
	notech_inv i_9027(.A(\nbus_13535[0] ), .Z(n_55048));
	notech_inv i_9011(.A(n_55030), .Z(n_55031));
	notech_inv i_9010(.A(\nbus_13539[0] ), .Z(n_55030));
	notech_inv i_9006(.A(n_55030), .Z(n_55026));
	notech_inv i_9002(.A(n_55030), .Z(n_55022));
	notech_inv i_8997(.A(n_55030), .Z(n_55017));
	notech_inv i_8993(.A(n_55030), .Z(n_55013));
	notech_inv i_8983(.A(n_55002), .Z(n_55003));
	notech_inv i_8982(.A(n_54983), .Z(n_55002));
	notech_inv i_8978(.A(n_55002), .Z(n_54998));
	notech_inv i_8974(.A(n_55002), .Z(n_54994));
	notech_inv i_8969(.A(n_55002), .Z(n_54989));
	notech_inv i_8965(.A(n_55002), .Z(n_54985));
	notech_inv i_8963(.A(n_55030), .Z(n_54983));
	notech_inv i_8955(.A(n_54974), .Z(n_54975));
	notech_inv i_8954(.A(n_54955), .Z(n_54974));
	notech_inv i_8950(.A(n_54974), .Z(n_54970));
	notech_inv i_8946(.A(n_54974), .Z(n_54966));
	notech_inv i_8941(.A(n_54974), .Z(n_54961));
	notech_inv i_8937(.A(n_54974), .Z(n_54957));
	notech_inv i_8935(.A(n_55030), .Z(n_54955));
	notech_inv i_8361(.A(n_54202), .Z(n_54267));
	notech_inv i_8360(.A(n_54202), .Z(n_54266));
	notech_inv i_8355(.A(n_54202), .Z(n_54261));
	notech_inv i_8350(.A(n_54202), .Z(n_54256));
	notech_inv i_8349(.A(n_54202), .Z(n_54255));
	notech_inv i_8344(.A(n_54202), .Z(n_54250));
	notech_inv i_8339(.A(n_54202), .Z(n_54245));
	notech_inv i_8338(.A(n_54202), .Z(n_54244));
	notech_inv i_8333(.A(n_54202), .Z(n_54239));
	notech_inv i_8327(.A(n_54202), .Z(n_54233));
	notech_inv i_8326(.A(n_54202), .Z(n_54232));
	notech_inv i_8321(.A(n_54202), .Z(n_54227));
	notech_inv i_8316(.A(n_54202), .Z(n_54222));
	notech_inv i_8315(.A(n_54202), .Z(n_54221));
	notech_inv i_8310(.A(n_54202), .Z(n_54216));
	notech_inv i_8305(.A(n_54202), .Z(n_54211));
	notech_inv i_8304(.A(n_54202), .Z(n_54210));
	notech_inv i_8299(.A(n_54202), .Z(n_54205));
	notech_inv i_8296(.A(\nbus_13538[0] ), .Z(n_54202));
	notech_inv i_8293(.A(n_54168), .Z(n_54199));
	notech_inv i_8292(.A(n_54168), .Z(n_54198));
	notech_inv i_8282(.A(n_54168), .Z(n_54188));
	notech_inv i_8281(.A(n_54168), .Z(n_54187));
	notech_inv i_8276(.A(n_54168), .Z(n_54182));
	notech_inv i_8271(.A(n_54168), .Z(n_54177));
	notech_inv i_8270(.A(n_54168), .Z(n_54176));
	notech_inv i_8265(.A(n_54168), .Z(n_54171));
	notech_inv i_8262(.A(\nbus_13538[0] ), .Z(n_54168));
	notech_inv i_7911(.A(n_53823), .Z(n_53824));
	notech_inv i_7910(.A(n_2887), .Z(n_53823));
	notech_inv i_7903(.A(n_53814), .Z(n_53815));
	notech_inv i_7902(.A(n_2898), .Z(n_53814));
	notech_inv i_7895(.A(n_53805), .Z(n_53806));
	notech_inv i_7894(.A(n_39845), .Z(n_53805));
	notech_inv i_7887(.A(n_53796), .Z(n_53797));
	notech_inv i_7886(.A(n_2885), .Z(n_53796));
	notech_inv i_7879(.A(n_53787), .Z(n_53788));
	notech_inv i_7878(.A(n_3108), .Z(n_53787));
	notech_inv i_7871(.A(n_53726), .Z(n_53727));
	notech_inv i_7870(.A(n_3097), .Z(n_53726));
	notech_ao4 i_322120(.A(n_58757), .B(n_40191), .C(n_57547), .D(n_39830), 
		.Z(n_3240));
	notech_ao4 i_222119(.A(n_58757), .B(n_40192), .C(n_57547), .D(n_39829), 
		.Z(n_3241));
	notech_ao3 i_2942(.A(n_59636), .B(\nbus_12535[1] ), .C(n_58859), .Z(n_3242
		));
	notech_ao4 i_122118(.A(n_58757), .B(n_40194), .C(n_57547), .D(n_39828), 
		.Z(n_3243));
	notech_ao3 i_2941(.A(n_59636), .B(\nbus_12535[0] ), .C(n_58859), .Z(n_3244
		));
	notech_ao4 i_21126540(.A(n_58757), .B(n_40102), .C(n_57547), .D(n_39820)
		, .Z(n_3245));
	notech_ao3 i_2945(.A(n_59636), .B(\nbus_12535[4] ), .C(n_58859), .Z(n_3239
		));
	notech_and2 i_775002(.A(n_2056), .B(n_40193), .Z(n_3246));
	notech_ao4 i_522122(.A(n_58757), .B(n_40189), .C(n_57547), .D(n_39832), 
		.Z(n_3238));
	notech_nao3 i_21275000(.A(n_59636), .B(n_40193), .C(n_1481), .Z(n_3247)
		);
	notech_nao3 i_8(.A(n_59636), .B(n_40193), .C(n_58859), .Z(n_5768));
	notech_nand2 i_3(.A(n_2124), .B(n_59636), .Z(n_5409));
	notech_and2 i_203(.A(n_5415), .B(n_5396), .Z(n_1994));
	notech_ao3 i_2946(.A(n_59636), .B(\nbus_12535[5] ), .C(n_58859), .Z(n_3237
		));
	notech_nand3 i_11(.A(n_40193), .B(n_59641), .C(n_38330), .Z(n_5276));
	notech_or4 i_152(.A(n_2833), .B(pg_fault), .C(pc_req), .D(n_2217), .Z(n_2056
		));
	notech_or2 i_6369(.A(idx_deco[1]), .B(idx_deco[0]), .Z(n_5396));
	notech_nor2 i_66845(.A(idx_deco[1]), .B(n_38656), .Z(n_5408));
	notech_ao4 i_622123(.A(n_58752), .B(n_40188), .C(n_57542), .D(n_39833), 
		.Z(n_3236));
	notech_nand2 i_625657(.A(n_59692), .B(n_1621), .Z(n_3235));
	notech_nor2 i_32173380(.A(n_1977), .B(n_58752), .Z(n_3248));
	notech_ao3 i_38973379(.A(n_59641), .B(in128[54]), .C(n_58859), .Z(n_3249
		));
	notech_ao3 i_46273377(.A(n_59636), .B(in128[86]), .C(n_58859), .Z(n_3250
		));
	notech_and4 i_223228(.A(n_1979), .B(n_1982), .C(n_2067), .D(n_1980), .Z(n_3251
		));
	notech_ao4 i_12725522(.A(n_58752), .B(n_39988), .C(n_57542), .D(n_38870)
		, .Z(n_3252));
	notech_ao4 i_12625521(.A(n_58757), .B(n_39987), .C(n_57542), .D(n_38868)
		, .Z(n_3253));
	notech_ao4 i_12525520(.A(n_58752), .B(n_39986), .C(n_57547), .D(n_38867)
		, .Z(n_3254));
	notech_ao4 i_12425519(.A(n_58757), .B(n_39985), .C(n_57547), .D(n_38865)
		, .Z(n_3255));
	notech_ao4 i_12325518(.A(n_58757), .B(n_39984), .C(n_57547), .D(n_38864)
		, .Z(n_3256));
	notech_ao4 i_12225517(.A(n_58757), .B(n_39983), .C(n_57547), .D(n_38862)
		, .Z(n_3257));
	notech_ao4 i_12125516(.A(n_58759), .B(n_39982), .C(n_57549), .D(n_38861)
		, .Z(n_3258));
	notech_ao4 i_12025515(.A(n_58759), .B(n_39981), .C(n_57549), .D(n_38859)
		, .Z(n_3259));
	notech_ao4 i_11925514(.A(n_58757), .B(n_39980), .C(n_57549), .D(n_38858)
		, .Z(n_3260));
	notech_ao4 i_11825513(.A(n_58757), .B(n_39979), .C(n_57547), .D(n_38856)
		, .Z(n_3261));
	notech_ao4 i_11725512(.A(n_58757), .B(n_39978), .C(n_57547), .D(n_38855)
		, .Z(n_3262));
	notech_ao4 i_11625511(.A(n_58757), .B(n_39977), .C(n_57547), .D(n_38853)
		, .Z(n_3263));
	notech_ao4 i_11525510(.A(n_58757), .B(n_39976), .C(n_57547), .D(n_38852)
		, .Z(n_3264));
	notech_ao4 i_11425509(.A(n_58752), .B(n_39975), .C(n_57547), .D(n_38850)
		, .Z(n_3265));
	notech_ao4 i_11325508(.A(n_58750), .B(n_39974), .C(n_57542), .D(n_38849)
		, .Z(n_3266));
	notech_ao4 i_11225507(.A(n_58750), .B(n_39973), .C(n_57540), .D(n_38847)
		, .Z(n_3267));
	notech_ao4 i_11125506(.A(n_58750), .B(n_39972), .C(n_57540), .D(n_38846)
		, .Z(n_3268));
	notech_ao4 i_11025505(.A(n_58750), .B(n_39971), .C(n_57540), .D(n_38844)
		, .Z(n_3269));
	notech_ao4 i_10925504(.A(n_58750), .B(n_39970), .C(n_57540), .D(n_38843)
		, .Z(n_3270));
	notech_ao4 i_10825503(.A(n_58750), .B(n_39969), .C(n_57540), .D(n_38841)
		, .Z(n_3271));
	notech_ao4 i_10725502(.A(n_58750), .B(n_39968), .C(n_57540), .D(n_38840)
		, .Z(n_3272));
	notech_ao4 i_10625501(.A(n_58750), .B(n_39967), .C(n_57540), .D(n_38838)
		, .Z(n_3273));
	notech_ao4 i_10525500(.A(n_58750), .B(n_39966), .C(n_57540), .D(n_38837)
		, .Z(n_3274));
	notech_ao4 i_10325498(.A(n_58750), .B(n_39964), .C(n_57540), .D(n_38833)
		, .Z(n_3275));
	notech_ao4 i_10225497(.A(n_58752), .B(n_39963), .C(n_57540), .D(n_38831)
		, .Z(n_3276));
	notech_ao4 i_10125496(.A(n_58752), .B(n_39962), .C(n_57542), .D(n_38830)
		, .Z(n_3277));
	notech_ao4 i_10025495(.A(n_58752), .B(n_39961), .C(n_57542), .D(n_38828)
		, .Z(n_3278));
	notech_ao4 i_9925494(.A(n_58752), .B(n_39960), .C(n_57542), .D(n_38827),
		 .Z(n_3279));
	notech_ao4 i_9825493(.A(n_58752), .B(n_39959), .C(n_57542), .D(n_38825),
		 .Z(n_3280));
	notech_ao4 i_9725492(.A(n_58752), .B(n_39958), .C(n_57542), .D(n_38824),
		 .Z(n_3281));
	notech_ao4 i_9625491(.A(n_58750), .B(n_39957), .C(n_57542), .D(n_38822),
		 .Z(n_3282));
	notech_ao4 i_9525490(.A(n_58752), .B(n_39956), .C(n_57542), .D(n_38821),
		 .Z(n_3283));
	notech_ao4 i_9425489(.A(n_58752), .B(n_39955), .C(n_57542), .D(n_38819),
		 .Z(n_3284));
	notech_ao4 i_9325488(.A(n_58752), .B(n_39954), .C(n_57542), .D(n_38818),
		 .Z(n_3285));
	notech_ao4 i_9225487(.A(n_58759), .B(n_39953), .C(n_57542), .D(n_38816),
		 .Z(n_3286));
	notech_ao4 i_9125486(.A(n_58764), .B(n_39952), .C(n_57554), .D(n_38815),
		 .Z(n_3287));
	notech_ao4 i_9025485(.A(n_58764), .B(n_39951), .C(n_57554), .D(n_38813),
		 .Z(n_3288));
	notech_ao4 i_8925484(.A(n_58764), .B(n_39950), .C(n_57554), .D(n_38812),
		 .Z(n_3289));
	notech_ao4 i_8825483(.A(n_58764), .B(n_39949), .C(n_57554), .D(n_38810),
		 .Z(n_3290));
	notech_ao4 i_8725482(.A(n_58764), .B(n_39948), .C(n_57554), .D(n_38809),
		 .Z(n_3291));
	notech_ao4 i_8625481(.A(n_58762), .B(n_39947), .C(n_57552), .D(n_38807),
		 .Z(n_3292));
	notech_ao4 i_8525480(.A(n_58762), .B(n_39946), .C(n_57552), .D(n_38806),
		 .Z(n_3293));
	notech_ao4 i_8425479(.A(n_58762), .B(n_39945), .C(n_57552), .D(n_38804),
		 .Z(n_3294));
	notech_ao4 i_8325478(.A(n_58764), .B(n_39944), .C(n_57554), .D(n_38803),
		 .Z(n_3295));
	notech_ao4 i_8225477(.A(n_58762), .B(n_39943), .C(n_57552), .D(n_38801),
		 .Z(n_3296));
	notech_ao4 i_8125476(.A(n_58764), .B(n_39942), .C(n_57554), .D(n_38800),
		 .Z(n_3297));
	notech_ao4 i_8025475(.A(n_58764), .B(n_39941), .C(n_57554), .D(n_38798),
		 .Z(n_3298));
	notech_ao4 i_7925474(.A(n_58764), .B(n_39940), .C(n_57554), .D(n_38797),
		 .Z(n_3299));
	notech_ao4 i_7825473(.A(n_58768), .B(n_39939), .C(n_57558), .D(n_38795),
		 .Z(n_3300));
	notech_ao4 i_7725472(.A(n_58768), .B(n_39938), .C(n_57558), .D(n_38794),
		 .Z(n_3301));
	notech_ao4 i_7625471(.A(n_58764), .B(n_39937), .C(n_57554), .D(n_38792),
		 .Z(n_3302));
	notech_ao4 i_7525470(.A(n_58764), .B(n_39936), .C(n_57554), .D(n_38791),
		 .Z(n_3303));
	notech_ao3 i_3382(.A(n_59636), .B(udeco[74]), .C(n_58859), .Z(n_3304));
	notech_ao4 i_7425469(.A(n_58764), .B(n_39935), .C(n_57554), .D(n_38789),
		 .Z(n_3305));
	notech_ao4 i_7325468(.A(n_58764), .B(n_39934), .C(n_57554), .D(n_38788),
		 .Z(n_3306));
	notech_ao3 i_3380(.A(n_59636), .B(udeco[72]), .C(n_58859), .Z(n_3307));
	notech_ao4 i_7225467(.A(n_58764), .B(n_39933), .C(n_57554), .D(n_38786),
		 .Z(n_3308));
	notech_ao4 i_7125466(.A(n_58762), .B(n_39932), .C(n_57552), .D(n_38785),
		 .Z(n_3309));
	notech_ao4 i_7025465(.A(n_58759), .B(n_39931), .C(n_57549), .D(n_38783),
		 .Z(n_3310));
	notech_ao4 i_6925464(.A(n_58759), .B(n_39930), .C(n_57549), .D(n_38782),
		 .Z(n_3311));
	notech_ao4 i_6825463(.A(n_58759), .B(n_39929), .C(n_57549), .D(n_38780),
		 .Z(n_3312));
	notech_ao3 i_3375(.A(n_59636), .B(udeco[67]), .C(n_58859), .Z(n_3313));
	notech_ao4 i_6725462(.A(n_58759), .B(n_39928), .C(n_57549), .D(n_38779),
		 .Z(n_3314));
	notech_ao4 i_6625461(.A(n_58759), .B(n_39927), .C(n_57549), .D(n_38777),
		 .Z(n_3315));
	notech_ao4 i_6525460(.A(n_58759), .B(n_39926), .C(n_57549), .D(n_38776),
		 .Z(n_3316));
	notech_ao3 i_3372(.A(n_59630), .B(udeco[64]), .C(n_58859), .Z(n_3317));
	notech_ao4 i_6425459(.A(n_58759), .B(n_39925), .C(n_57549), .D(n_38774),
		 .Z(n_3318));
	notech_ao4 i_6325458(.A(n_58759), .B(n_39924), .C(n_57549), .D(n_38773),
		 .Z(n_3319));
	notech_ao4 i_6225457(.A(n_58759), .B(n_39923), .C(n_57549), .D(n_38771),
		 .Z(n_3320));
	notech_ao3 i_3369(.A(n_59630), .B(udeco[61]), .C(n_58854), .Z(n_3321));
	notech_ao4 i_6125456(.A(n_58759), .B(n_39922), .C(n_57549), .D(n_38770),
		 .Z(n_3322));
	notech_ao3 i_3368(.A(n_59630), .B(udeco[60]), .C(n_58854), .Z(n_3323));
	notech_ao4 i_6025455(.A(n_58762), .B(n_39921), .C(n_57552), .D(n_38768),
		 .Z(n_3324));
	notech_ao3 i_3367(.A(n_59630), .B(udeco[59]), .C(n_58854), .Z(n_3325));
	notech_ao4 i_5925454(.A(n_58762), .B(n_39920), .C(n_57552), .D(n_38767),
		 .Z(n_3326));
	notech_ao3 i_3366(.A(n_59630), .B(udeco[58]), .C(n_58854), .Z(n_3327));
	notech_ao4 i_5825453(.A(n_58762), .B(n_39919), .C(n_57552), .D(n_38765),
		 .Z(n_3328));
	notech_ao3 i_3365(.A(n_59630), .B(udeco[57]), .C(n_58854), .Z(n_3329));
	notech_ao4 i_5725452(.A(n_58762), .B(n_39918), .C(n_57552), .D(n_38764),
		 .Z(n_3330));
	notech_ao3 i_3364(.A(n_59630), .B(udeco[56]), .C(n_58854), .Z(n_3331));
	notech_ao4 i_5625451(.A(n_58762), .B(n_39917), .C(n_57552), .D(n_38762),
		 .Z(n_3332));
	notech_ao3 i_3363(.A(n_59630), .B(udeco[55]), .C(n_58854), .Z(n_3333));
	notech_ao4 i_5525450(.A(n_58762), .B(n_39916), .C(n_57552), .D(n_38761),
		 .Z(n_3334));
	notech_ao3 i_3362(.A(n_59636), .B(udeco[54]), .C(n_58859), .Z(n_3335));
	notech_ao4 i_5425449(.A(n_58759), .B(n_39915), .C(n_57549), .D(n_38759),
		 .Z(n_3336));
	notech_ao3 i_3361(.A(n_59630), .B(udeco[53]), .C(n_58854), .Z(n_3337));
	notech_ao4 i_5325448(.A(n_58762), .B(n_39914), .C(n_57552), .D(n_38758),
		 .Z(n_3338));
	notech_ao3 i_3360(.A(n_59630), .B(udeco[52]), .C(n_58854), .Z(n_3339));
	notech_ao4 i_5225447(.A(n_58762), .B(n_39913), .C(n_57552), .D(n_38756),
		 .Z(n_3340));
	notech_ao3 i_3359(.A(n_59630), .B(udeco[51]), .C(n_58854), .Z(n_3341));
	notech_ao4 i_5125446(.A(n_58762), .B(n_39912), .C(n_57552), .D(n_38755),
		 .Z(n_3342));
	notech_ao3 i_3358(.A(n_59641), .B(udeco[50]), .C(n_58859), .Z(n_3343));
	notech_ao4 i_5025445(.A(n_58739), .B(n_39911), .C(n_57540), .D(n_38753),
		 .Z(n_3344));
	notech_ao3 i_3357(.A(n_59642), .B(udeco[49]), .C(n_58863), .Z(n_3345));
	notech_ao4 i_4925444(.A(n_58739), .B(n_39910), .C(n_57529), .D(n_38752),
		 .Z(n_3346));
	notech_ao3 i_3356(.A(n_59642), .B(udeco[48]), .C(n_58864), .Z(n_3347));
	notech_ao4 i_4825443(.A(n_58739), .B(n_39909), .C(n_57529), .D(n_38750),
		 .Z(n_3348));
	notech_ao3 i_3355(.A(n_59642), .B(udeco[47]), .C(n_58863), .Z(n_3349));
	notech_ao4 i_4725442(.A(n_58739), .B(n_39908), .C(n_57529), .D(n_38749),
		 .Z(n_3350));
	notech_ao3 i_3354(.A(n_59641), .B(udeco[46]), .C(n_58863), .Z(n_3351));
	notech_ao4 i_4625441(.A(n_58739), .B(n_39907), .C(n_57529), .D(n_38747),
		 .Z(n_3352));
	notech_ao3 i_3353(.A(n_59641), .B(udeco[45]), .C(n_58863), .Z(n_3353));
	notech_ao4 i_4525440(.A(n_58736), .B(n_39906), .C(n_57529), .D(n_38746),
		 .Z(n_3354));
	notech_ao3 i_3352(.A(n_59642), .B(udeco[44]), .C(n_58864), .Z(n_3355));
	notech_ao4 i_4425439(.A(n_58736), .B(n_39905), .C(n_57526), .D(n_38744),
		 .Z(n_3356));
	notech_ao3 i_3351(.A(n_59642), .B(udeco[43]), .C(n_58864), .Z(n_3357));
	notech_ao4 i_4325438(.A(n_58736), .B(n_39904), .C(n_57526), .D(n_38743),
		 .Z(n_3358));
	notech_ao3 i_3350(.A(n_59642), .B(udeco[42]), .C(n_58864), .Z(n_3359));
	notech_ao4 i_4225437(.A(n_58739), .B(n_39903), .C(n_57529), .D(n_38741),
		 .Z(n_3360));
	notech_ao3 i_3349(.A(n_59642), .B(udeco[41]), .C(n_58864), .Z(n_3361));
	notech_ao4 i_4125436(.A(n_58739), .B(n_39902), .C(n_57529), .D(n_38740),
		 .Z(n_3362));
	notech_ao3 i_3348(.A(n_59642), .B(udeco[40]), .C(n_58864), .Z(n_3363));
	notech_ao4 i_4025435(.A(n_58739), .B(n_39901), .C(n_57529), .D(n_38738),
		 .Z(n_3364));
	notech_ao3 i_3347(.A(n_59642), .B(udeco[39]), .C(n_58864), .Z(n_3365));
	notech_ao4 i_3925434(.A(n_58739), .B(n_39900), .C(n_57531), .D(n_38737),
		 .Z(n_3366));
	notech_ao3 i_3346(.A(n_59642), .B(udeco[38]), .C(n_58863), .Z(n_3367));
	notech_ao4 i_3825433(.A(n_58741), .B(n_39899), .C(n_57529), .D(n_38735),
		 .Z(n_3368));
	notech_ao3 i_3345(.A(n_59641), .B(udeco[37]), .C(n_58863), .Z(n_3369));
	notech_ao4 i_3725432(.A(n_58741), .B(n_39898), .C(n_57531), .D(n_38734),
		 .Z(n_3370));
	notech_ao3 i_3344(.A(n_59641), .B(udeco[36]), .C(n_58863), .Z(n_3371));
	notech_ao4 i_3625431(.A(n_58741), .B(n_39897), .C(n_57531), .D(n_38732),
		 .Z(n_3372));
	notech_ao3 i_3343(.A(n_59641), .B(udeco[35]), .C(n_58859), .Z(n_3373));
	notech_ao4 i_3525430(.A(n_58739), .B(n_39896), .C(n_57531), .D(n_38731),
		 .Z(n_3374));
	notech_ao3 i_3342(.A(n_59641), .B(udeco[34]), .C(n_58863), .Z(n_3375));
	notech_ao4 i_3425429(.A(n_58739), .B(n_39895), .C(n_57529), .D(n_38729),
		 .Z(n_3376));
	notech_ao3 i_3341(.A(n_59641), .B(udeco[33]), .C(n_58863), .Z(n_3377));
	notech_ao4 i_3325428(.A(n_58739), .B(n_39894), .C(n_57529), .D(n_38728),
		 .Z(n_3378));
	notech_ao3 i_3340(.A(n_59641), .B(udeco[32]), .C(n_58863), .Z(n_3379));
	notech_ao4 i_3225427(.A(n_58739), .B(n_39893), .C(n_57529), .D(n_38726),
		 .Z(n_3380));
	notech_ao3 i_3339(.A(n_59641), .B(udeco[31]), .C(n_58863), .Z(n_3381));
	notech_ao4 i_3125426(.A(n_58739), .B(n_39892), .C(n_57529), .D(n_38725),
		 .Z(n_3382));
	notech_ao3 i_3338(.A(n_59641), .B(udeco[30]), .C(n_58863), .Z(n_3383));
	notech_ao4 i_3025425(.A(n_58736), .B(n_39891), .C(n_57529), .D(n_38723),
		 .Z(n_3384));
	notech_ao3 i_3337(.A(n_59641), .B(udeco[29]), .C(n_58863), .Z(n_3385));
	notech_ao4 i_2925424(.A(n_58734), .B(n_39890), .C(n_57526), .D(n_38722),
		 .Z(n_3386));
	notech_ao3 i_3336(.A(n_59641), .B(udeco[28]), .C(n_58863), .Z(n_3387));
	notech_ao4 i_2825423(.A(n_58734), .B(n_39889), .C(n_57524), .D(n_38720),
		 .Z(n_3388));
	notech_ao3 i_3335(.A(n_59641), .B(udeco[27]), .C(n_58854), .Z(n_3389));
	notech_ao4 i_2725422(.A(n_58734), .B(n_39888), .C(n_57524), .D(n_38719),
		 .Z(n_3390));
	notech_ao3 i_3334(.A(n_59641), .B(udeco[26]), .C(n_58849), .Z(n_3391));
	notech_ao4 i_2625421(.A(n_58734), .B(n_39887), .C(n_57524), .D(n_38717),
		 .Z(n_3392));
	notech_ao3 i_3333(.A(n_59641), .B(udeco[25]), .C(n_58849), .Z(n_3393));
	notech_ao4 i_2525420(.A(n_58734), .B(n_39886), .C(n_57526), .D(n_38716),
		 .Z(n_3394));
	notech_ao3 i_3332(.A(n_59630), .B(udeco[24]), .C(n_58845), .Z(n_3395));
	notech_ao4 i_2425419(.A(n_58734), .B(n_39885), .C(n_57524), .D(n_38714),
		 .Z(n_3396));
	notech_ao3 i_3331(.A(n_59624), .B(udeco[23]), .C(n_58845), .Z(n_3397));
	notech_ao4 i_2325418(.A(n_58734), .B(n_39884), .C(n_57524), .D(n_38713),
		 .Z(n_3398));
	notech_ao3 i_3330(.A(n_59624), .B(udeco[22]), .C(n_58845), .Z(n_3399));
	notech_ao4 i_2225417(.A(n_58734), .B(n_39883), .C(n_57524), .D(n_38711),
		 .Z(n_3400));
	notech_ao3 i_3329(.A(n_59624), .B(udeco[21]), .C(n_58849), .Z(n_3401));
	notech_ao4 i_2125416(.A(n_58734), .B(n_39882), .C(n_57524), .D(n_38710),
		 .Z(n_3402));
	notech_ao3 i_3328(.A(n_59619), .B(udeco[20]), .C(n_58849), .Z(n_3403));
	notech_ao4 i_2025415(.A(n_58734), .B(n_39881), .C(n_57524), .D(n_38708),
		 .Z(n_3404));
	notech_ao3 i_3327(.A(n_59619), .B(udeco[19]), .C(n_58849), .Z(n_3405));
	notech_ao4 i_1925414(.A(n_58736), .B(n_39880), .C(n_57524), .D(n_38707),
		 .Z(n_3406));
	notech_ao3 i_3326(.A(n_59624), .B(udeco[18]), .C(n_58849), .Z(n_3407));
	notech_ao4 i_1825413(.A(n_58736), .B(n_39879), .C(n_57526), .D(n_38705),
		 .Z(n_3408));
	notech_ao3 i_3325(.A(n_59624), .B(udeco[17]), .C(n_58849), .Z(n_3409));
	notech_ao4 i_1725412(.A(n_58736), .B(n_39878), .C(n_57526), .D(n_38704),
		 .Z(n_3410));
	notech_ao3 i_3324(.A(n_59624), .B(udeco[16]), .C(n_58849), .Z(n_3411));
	notech_ao4 i_1625411(.A(n_58736), .B(n_39877), .C(n_57526), .D(n_38702),
		 .Z(n_3412));
	notech_ao3 i_3323(.A(n_59624), .B(udeco[15]), .C(n_58845), .Z(n_3413));
	notech_ao4 i_1525410(.A(n_58736), .B(n_39876), .C(n_57526), .D(n_38701),
		 .Z(n_3414));
	notech_ao3 i_3322(.A(n_59624), .B(udeco[14]), .C(n_58845), .Z(n_3415));
	notech_ao4 i_1425409(.A(n_58736), .B(n_39875), .C(n_57526), .D(n_38699),
		 .Z(n_3416));
	notech_ao3 i_3321(.A(n_59624), .B(udeco[13]), .C(n_58845), .Z(n_3417));
	notech_ao4 i_1325408(.A(n_58736), .B(n_39874), .C(n_57526), .D(n_38698),
		 .Z(n_3418));
	notech_ao3 i_3320(.A(n_59624), .B(udeco[12]), .C(n_58845), .Z(n_3419));
	notech_ao4 i_1225407(.A(n_58736), .B(n_39873), .C(n_57526), .D(n_38696),
		 .Z(n_3420));
	notech_ao3 i_3319(.A(n_59619), .B(udeco[11]), .C(n_58845), .Z(n_3421));
	notech_ao4 i_1125406(.A(n_58736), .B(n_39872), .C(n_57526), .D(n_38695),
		 .Z(n_3422));
	notech_ao3 i_3318(.A(n_59619), .B(udeco[10]), .C(n_58845), .Z(n_3423));
	notech_ao4 i_1025405(.A(n_58736), .B(n_39871), .C(n_57526), .D(n_38693),
		 .Z(n_3424));
	notech_ao3 i_3317(.A(n_59619), .B(udeco[9]), .C(n_58845), .Z(n_3425));
	notech_ao4 i_925404(.A(n_58741), .B(n_39870), .C(n_57526), .D(n_38692), 
		.Z(n_3426));
	notech_ao3 i_3316(.A(n_59619), .B(udeco[8]), .C(n_58845), .Z(n_3427));
	notech_ao4 i_825403(.A(n_58747), .B(n_39869), .C(n_57537), .D(n_38690), 
		.Z(n_3428));
	notech_ao3 i_3315(.A(n_59619), .B(udeco[7]), .C(n_58845), .Z(n_3429));
	notech_ao4 i_725402(.A(n_58747), .B(n_39868), .C(n_57537), .D(n_38689), 
		.Z(n_3430));
	notech_ao3 i_3314(.A(n_59619), .B(udeco[6]), .C(n_58845), .Z(n_3431));
	notech_ao4 i_625401(.A(n_58747), .B(n_39867), .C(n_57537), .D(n_38687), 
		.Z(n_3432));
	notech_ao3 i_3313(.A(n_59619), .B(udeco[5]), .C(n_58845), .Z(n_3433));
	notech_ao4 i_525400(.A(n_58747), .B(n_39866), .C(n_57537), .D(n_38686), 
		.Z(n_3434));
	notech_ao3 i_3312(.A(n_59619), .B(udeco[4]), .C(n_58849), .Z(n_3435));
	notech_ao4 i_425399(.A(n_58747), .B(n_39865), .C(n_57537), .D(n_38684), 
		.Z(n_3436));
	notech_ao3 i_3311(.A(n_59619), .B(udeco[3]), .C(n_58853), .Z(n_3437));
	notech_ao4 i_325398(.A(n_58745), .B(n_39864), .C(n_57535), .D(n_38683), 
		.Z(n_3438));
	notech_ao3 i_3310(.A(n_59619), .B(udeco[2]), .C(n_58853), .Z(n_3439));
	notech_ao4 i_225397(.A(n_58745), .B(n_39863), .C(n_57535), .D(n_38681), 
		.Z(n_3440));
	notech_ao3 i_3309(.A(n_59619), .B(udeco[1]), .C(n_58853), .Z(n_3441));
	notech_ao4 i_125396(.A(n_58745), .B(n_39862), .C(n_57535), .D(n_38680), 
		.Z(n_3442));
	notech_ao3 i_3308(.A(n_59619), .B(udeco[0]), .C(n_58853), .Z(n_3443));
	notech_ao4 i_20826326(.A(n_58747), .B(n_40099), .C(n_57537), .D(n_39417)
		, .Z(n_3444));
	notech_ao3 i_11373263(.A(n_59619), .B(in128[124]), .C(n_58853), .Z(n_3445
		));
	notech_ao4 i_20426322(.A(n_58747), .B(n_40095), .C(n_57537), .D(n_39411)
		, .Z(n_3446));
	notech_ao3 i_11773259(.A(n_59624), .B(in128[120]), .C(n_58853), .Z(n_3447
		));
	notech_ao4 i_20326321(.A(n_58747), .B(n_40094), .C(n_57537), .D(n_39409)
		, .Z(n_3448));
	notech_ao3 i_11873258(.A(n_59629), .B(in128[119]), .C(n_58854), .Z(n_3449
		));
	notech_ao4 i_20126319(.A(n_58747), .B(n_40092), .C(n_57537), .D(n_39406)
		, .Z(n_3450));
	notech_ao3 i_12073256(.A(n_59629), .B(in128[117]), .C(n_58854), .Z(n_3451
		));
	notech_ao4 i_20026318(.A(n_58750), .B(n_40091), .C(n_57540), .D(n_39405)
		, .Z(n_3452));
	notech_ao3 i_12173255(.A(n_59629), .B(in128[116]), .C(n_58854), .Z(n_3453
		));
	notech_ao4 i_19926317(.A(n_58750), .B(n_40090), .C(n_57540), .D(n_39403)
		, .Z(n_3454));
	notech_ao3 i_12273254(.A(n_59629), .B(in128[115]), .C(n_58853), .Z(n_3455
		));
	notech_ao4 i_19826316(.A(n_58750), .B(n_40089), .C(n_57540), .D(n_39402)
		, .Z(n_3456));
	notech_ao3 i_12373253(.A(n_59629), .B(in128[114]), .C(n_58853), .Z(n_3457
		));
	notech_ao4 i_17926297(.A(n_58747), .B(n_40070), .C(n_57537), .D(n_39373)
		, .Z(n_3458));
	notech_ao3 i_14273234(.A(n_59629), .B(in128[95]), .C(n_58849), .Z(n_3459
		));
	notech_ao4 i_17626294(.A(n_58747), .B(n_40067), .C(n_57537), .D(n_39369)
		, .Z(n_3460));
	notech_ao3 i_14573231(.A(n_59630), .B(in128[92]), .C(n_58849), .Z(n_3461
		));
	notech_ao4 i_17426292(.A(n_58747), .B(n_40065), .C(n_57537), .D(n_39366)
		, .Z(n_3462));
	notech_ao3 i_14773229(.A(n_59630), .B(in128[90]), .C(n_58849), .Z(n_3463
		));
	notech_ao4 i_17326291(.A(n_58747), .B(n_40064), .C(n_57537), .D(n_39364)
		, .Z(n_3464));
	notech_ao3 i_14873228(.A(n_59630), .B(in128[89]), .C(n_58849), .Z(n_3465
		));
	notech_ao4 i_16926287(.A(n_58747), .B(n_40060), .C(n_57537), .D(n_39359)
		, .Z(n_3466));
	notech_ao3 i_1473362(.A(n_59630), .B(in128[85]), .C(n_58849), .Z(n_3467)
		);
	notech_ao4 i_16826286(.A(n_58745), .B(n_40059), .C(n_57535), .D(n_39357)
		, .Z(n_3468));
	notech_ao3 i_3073346(.A(n_59630), .B(in128[84]), .C(n_58853), .Z(n_3469)
		);
	notech_ao4 i_16726285(.A(n_58741), .B(n_40058), .C(n_57531), .D(n_39356)
		, .Z(n_3470));
	notech_ao3 i_2573351(.A(n_59630), .B(in128[83]), .C(n_58853), .Z(n_3471)
		);
	notech_ao4 i_16626284(.A(n_58741), .B(n_40057), .C(n_57531), .D(n_39355)
		, .Z(n_3472));
	notech_ao3 i_2273354(.A(n_59629), .B(in128[82]), .C(n_58853), .Z(n_3473)
		);
	notech_ao4 i_16526283(.A(n_58741), .B(n_40056), .C(n_57531), .D(n_39354)
		, .Z(n_3474));
	notech_ao3 i_2073356(.A(n_59629), .B(in128[81]), .C(n_58853), .Z(n_3475)
		);
	notech_ao4 i_16426282(.A(n_58741), .B(n_40055), .C(n_57531), .D(n_39353)
		, .Z(n_3476));
	notech_ao3 i_6273314(.A(n_59629), .B(in128[80]), .C(n_58853), .Z(n_3477)
		);
	notech_ao4 i_14726265(.A(n_58741), .B(n_40038), .C(n_57531), .D(n_39336)
		, .Z(n_3478));
	notech_ao3 i_7073306(.A(n_59629), .B(in128[63]), .C(n_58853), .Z(n_3479)
		);
	notech_ao4 i_13926257(.A(n_58741), .B(n_40030), .C(n_57531), .D(n_39328)
		, .Z(n_3480));
	notech_ao3 i_8273294(.A(n_59624), .B(in128[55]), .C(n_58877), .Z(n_3481)
		);
	notech_ao4 i_12826246(.A(n_58741), .B(n_40019), .C(n_57531), .D(n_39312)
		, .Z(n_3482));
	notech_ao3 i_6473312(.A(n_59629), .B(in128[44]), .C(n_58877), .Z(n_3483)
		);
	notech_ao4 i_12726245(.A(n_58741), .B(n_40018), .C(n_57531), .D(n_39311)
		, .Z(n_3484));
	notech_ao3 i_7573301(.A(n_59629), .B(in128[43]), .C(n_58877), .Z(n_3485)
		);
	notech_ao4 i_12626244(.A(n_58741), .B(n_40017), .C(n_57531), .D(n_39309)
		, .Z(n_3486));
	notech_ao4 i_12526243(.A(n_58741), .B(n_40016), .C(n_57531), .D(n_39308)
		, .Z(n_3487));
	notech_ao3 i_4673330(.A(n_59629), .B(in128[41]), .C(n_58877), .Z(n_3488)
		);
	notech_ao4 i_12426242(.A(n_58745), .B(n_40015), .C(n_57535), .D(n_39307)
		, .Z(n_3489));
	notech_ao3 i_7973297(.A(n_59629), .B(in128[40]), .C(n_58877), .Z(n_3490)
		);
	notech_ao4 i_11326231(.A(n_58745), .B(n_40004), .C(n_57535), .D(n_39292)
		, .Z(n_3491));
	notech_ao3 i_5373323(.A(n_59629), .B(in128[29]), .C(n_58877), .Z(n_3492)
		);
	notech_ao4 i_10726225(.A(n_58745), .B(n_39998), .C(n_57535), .D(n_39283)
		, .Z(n_3493));
	notech_ao4 i_10126219(.A(n_58745), .B(n_39992), .C(n_57535), .D(n_39274)
		, .Z(n_3494));
	notech_ao4 i_10026218(.A(n_58745), .B(n_39991), .C(n_57535), .D(n_39272)
		, .Z(n_3495));
	notech_ao4 i_9926217(.A(n_58745), .B(n_40172), .C(n_57535), .D(n_39271),
		 .Z(n_3496));
	notech_ao4 i_9826216(.A(n_58745), .B(n_40173), .C(n_57535), .D(n_39269),
		 .Z(n_3497));
	notech_ao4 i_9726215(.A(n_58745), .B(n_40206), .C(n_57535), .D(n_39268),
		 .Z(n_3498));
	notech_ao4 i_9626214(.A(n_58745), .B(n_40207), .C(n_57535), .D(n_39266),
		 .Z(n_3499));
	notech_ao4 i_9526213(.A(n_58745), .B(n_40208), .C(n_57535), .D(n_39265),
		 .Z(n_3500));
	notech_ao4 i_9426212(.A(n_58790), .B(n_40197), .C(n_57558), .D(n_39263),
		 .Z(n_3501));
	notech_ao4 i_9326211(.A(n_58786), .B(n_40196), .C(n_57580), .D(n_39262),
		 .Z(n_3502));
	notech_ao4 i_9226210(.A(n_58790), .B(n_40174), .C(n_57580), .D(n_39260),
		 .Z(n_3503));
	notech_ao4 i_9126209(.A(n_58790), .B(n_40202), .C(n_57580), .D(n_39259),
		 .Z(n_3504));
	notech_ao4 i_8726205(.A(n_58790), .B(n_40198), .C(n_57580), .D(n_39253),
		 .Z(n_3505));
	notech_ao4 i_8626204(.A(n_58786), .B(n_40175), .C(n_57580), .D(n_39251),
		 .Z(n_3506));
	notech_ao4 i_8526203(.A(n_58786), .B(n_40176), .C(n_57576), .D(n_39250),
		 .Z(n_3507));
	notech_ao4 i_8226200(.A(n_58786), .B(n_40178), .C(n_57576), .D(n_39244),
		 .Z(n_3508));
	notech_ao4 i_8126199(.A(n_58786), .B(n_40179), .C(n_57576), .D(n_39243),
		 .Z(n_3509));
	notech_ao4 i_7026188(.A(n_58786), .B(n_40166), .C(n_57576), .D(n_39226),
		 .Z(n_3510));
	notech_ao3 i_10373273(.A(n_59629), .B(\to_acu2_0[69] ), .C(n_58881), .Z(n_3511
		));
	notech_ao4 i_6826186(.A(n_58790), .B(n_40107), .C(n_57576), .D(n_39223),
		 .Z(n_3512));
	notech_ao3 i_15073226(.A(n_59629), .B(\to_acu2_0[67] ), .C(n_58881), .Z(n_3513
		));
	notech_ao4 i_6726185(.A(n_58790), .B(n_40108), .C(n_57580), .D(n_39222),
		 .Z(n_3514));
	notech_ao3 i_15173225(.A(n_59629), .B(\to_acu2_0[66] ), .C(n_58881), .Z(n_3515
		));
	notech_ao4 i_6626184(.A(n_58790), .B(n_40109), .C(n_57580), .D(n_39220),
		 .Z(n_3516));
	notech_ao3 i_15273224(.A(n_59642), .B(\to_acu2_0[65] ), .C(n_58881), .Z(n_3517
		));
	notech_ao4 i_6526183(.A(n_58790), .B(n_40110), .C(n_57580), .D(n_39219),
		 .Z(n_3518));
	notech_ao3 i_15373223(.A(n_59663), .B(\to_acu2_0[64] ), .C(n_58881), .Z(n_3519
		));
	notech_ao4 i_2926147(.A(n_58790), .B(n_40163), .C(n_57582), .D(n_39166),
		 .Z(n_3520));
	notech_ao3 i_8873288(.A(n_59663), .B(\to_acu2_0[28] ), .C(n_58877), .Z(n_3521
		));
	notech_ao4 i_2826146(.A(n_58790), .B(n_40159), .C(n_57580), .D(n_39164),
		 .Z(n_3522));
	notech_ao3 i_8773289(.A(n_59663), .B(\to_acu2_0[27] ), .C(n_58877), .Z(n_3523
		));
	notech_ao4 i_2726145(.A(n_58790), .B(n_40160), .C(n_57580), .D(n_39163),
		 .Z(n_3524));
	notech_ao3 i_5573321(.A(n_59658), .B(\to_acu2_0[26] ), .C(n_58873), .Z(n_3525
		));
	notech_ao4 i_2626144(.A(n_58790), .B(n_40162), .C(n_57580), .D(n_39161),
		 .Z(n_3526));
	notech_ao3 i_8673290(.A(n_59658), .B(\to_acu2_0[25] ), .C(n_58873), .Z(n_3527
		));
	notech_ao4 i_2526143(.A(n_58790), .B(n_40161), .C(n_57580), .D(n_39160),
		 .Z(n_3528));
	notech_ao3 i_8573291(.A(n_59663), .B(\to_acu2_0[24] ), .C(n_58873), .Z(n_3529
		));
	notech_ao4 i_2426142(.A(n_58790), .B(n_40157), .C(n_57580), .D(n_39158),
		 .Z(n_3530));
	notech_ao3 i_10273274(.A(n_59663), .B(\to_acu2_0[23] ), .C(n_58877), .Z(n_3531
		));
	notech_ao4 i_2326141(.A(n_58786), .B(n_40158), .C(n_57580), .D(n_39157),
		 .Z(n_3532));
	notech_ao3 i_10173275(.A(n_59663), .B(\to_acu2_0[22] ), .C(n_58877), .Z(n_3533
		));
	notech_ao4 i_1526133(.A(n_58784), .B(n_40150), .C(n_57576), .D(n_39145),
		 .Z(n_3534));
	notech_ao3 i_9673280(.A(n_59663), .B(\to_acu2_0[14] ), .C(n_58877), .Z(n_3535
		));
	notech_ao4 i_1426132(.A(n_58784), .B(n_40151), .C(n_57574), .D(n_39143),
		 .Z(n_3536));
	notech_ao3 i_3773339(.A(n_59663), .B(\to_acu2_0[13] ), .C(n_58877), .Z(n_3537
		));
	notech_ao4 i_1326131(.A(n_58784), .B(n_40154), .C(n_57574), .D(n_39142),
		 .Z(n_3538));
	notech_ao3 i_8373293(.A(n_59663), .B(\to_acu2_0[12] ), .C(n_58877), .Z(n_3539
		));
	notech_ao4 i_926127(.A(n_58784), .B(n_40167), .C(n_57574), .D(n_39136), 
		.Z(n_3540));
	notech_ao3 i_9373283(.A(n_59663), .B(\to_acu2_0[8] ), .C(n_58877), .Z(n_3541
		));
	notech_ao4 i_526123(.A(n_58784), .B(n_40209), .C(n_57574), .D(n_39130), 
		.Z(n_3542));
	notech_ao3 i_1373363(.A(n_59658), .B(\to_acu2_0[4] ), .C(n_58881), .Z(n_3543
		));
	notech_ao4 i_326121(.A(n_58784), .B(n_40147), .C(n_57574), .D(n_39127), 
		.Z(n_3544));
	notech_ao3 i_5673320(.A(n_59658), .B(\to_acu2_0[2] ), .C(n_58882), .Z(n_3545
		));
	notech_ao4 i_126119(.A(n_58784), .B(n_40214), .C(n_57574), .D(n_39124), 
		.Z(n_3546));
	notech_ao3 i_3173345(.A(n_59658), .B(\to_acu2_0[0] ), .C(n_58882), .Z(n_3547
		));
	notech_ao4 i_527805(.A(n_58784), .B(n_225793362), .C(n_57574), .D(n_38514
		), .Z(n_3548));
	notech_ao4 i_327803(.A(n_58784), .B(n_224193378), .C(n_57574), .D(n_38512
		), .Z(n_3549));
	notech_ao4 i_227802(.A(n_58784), .B(n_223393386), .C(n_57574), .D(n_38511
		), .Z(n_3550));
	notech_ao4 i_21026539(.A(n_58786), .B(n_40101), .C(n_57574), .D(n_39818)
		, .Z(n_3551));
	notech_ao3 i_11173265(.A(n_59658), .B(in128[126]), .C(n_58882), .Z(n_3552
		));
	notech_ao4 i_20926538(.A(n_58786), .B(n_40100), .C(n_57576), .D(n_39816)
		, .Z(n_3553));
	notech_ao3 i_11273264(.A(n_59653), .B(in128[125]), .C(n_58882), .Z(n_3554
		));
	notech_ao4 i_20826537(.A(n_58786), .B(n_40099), .C(n_57576), .D(n_39814)
		, .Z(n_3555));
	notech_ao4 i_20726536(.A(n_58786), .B(n_40098), .C(n_57576), .D(n_39813)
		, .Z(n_3556));
	notech_ao3 i_11473262(.A(n_59653), .B(in128[123]), .C(n_58882), .Z(n_3557
		));
	notech_ao4 i_20626535(.A(n_58786), .B(n_40097), .C(n_57576), .D(n_39811)
		, .Z(n_3558));
	notech_ao3 i_11573261(.A(n_59653), .B(in128[122]), .C(n_58882), .Z(n_3559
		));
	notech_ao4 i_20526534(.A(n_58784), .B(n_40096), .C(n_57576), .D(n_39809)
		, .Z(n_3560));
	notech_ao3 i_11673260(.A(n_59658), .B(in128[121]), .C(n_58882), .Z(n_3561
		));
	notech_ao4 i_20426533(.A(n_58784), .B(n_40095), .C(n_57574), .D(n_39807)
		, .Z(n_3562));
	notech_ao4 i_20326532(.A(n_58784), .B(n_40094), .C(n_57574), .D(n_39806)
		, .Z(n_3563));
	notech_ao4 i_20226531(.A(n_58786), .B(n_40093), .C(n_57576), .D(n_39805)
		, .Z(n_3564));
	notech_ao3 i_11973257(.A(n_59658), .B(in128[118]), .C(n_58882), .Z(n_3565
		));
	notech_ao4 i_20126530(.A(n_58786), .B(n_40092), .C(n_57576), .D(n_39803)
		, .Z(n_3566));
	notech_ao4 i_20026529(.A(n_58792), .B(n_40091), .C(n_57576), .D(n_39802)
		, .Z(n_3567));
	notech_ao4 i_19926528(.A(n_58797), .B(n_40090), .C(n_57587), .D(n_39801)
		, .Z(n_3568));
	notech_ao4 i_19826527(.A(n_58795), .B(n_40089), .C(n_57585), .D(n_39800)
		, .Z(n_3569));
	notech_ao4 i_19726526(.A(n_58797), .B(n_40088), .C(n_57587), .D(n_39799)
		, .Z(n_3570));
	notech_ao3 i_12473252(.A(n_59658), .B(in128[113]), .C(n_58882), .Z(n_3571
		));
	notech_ao4 i_19626525(.A(n_58797), .B(n_40087), .C(n_57587), .D(n_39797)
		, .Z(n_3572));
	notech_ao3 i_12573251(.A(n_59658), .B(in128[112]), .C(n_58882), .Z(n_3573
		));
	notech_ao4 i_19526524(.A(n_58797), .B(n_40086), .C(n_57587), .D(n_39795)
		, .Z(n_3574));
	notech_ao3 i_12673250(.A(n_59658), .B(in128[111]), .C(n_58882), .Z(n_3575
		));
	notech_ao4 i_19426523(.A(n_58795), .B(n_40085), .C(n_57585), .D(n_39793)
		, .Z(n_3576));
	notech_ao3 i_12773249(.A(n_59658), .B(in128[110]), .C(n_58881), .Z(n_3577
		));
	notech_ao4 i_19326522(.A(n_58795), .B(n_40084), .C(n_57585), .D(n_39791)
		, .Z(n_3578));
	notech_ao3 i_12873248(.A(n_59663), .B(in128[109]), .C(n_58881), .Z(n_3579
		));
	notech_ao4 i_19226521(.A(n_58795), .B(n_40083), .C(n_57585), .D(n_39789)
		, .Z(n_3580));
	notech_ao3 i_12973247(.A(n_59664), .B(in128[108]), .C(n_58881), .Z(n_3581
		));
	notech_ao4 i_19126520(.A(n_58795), .B(n_40082), .C(n_57585), .D(n_39787)
		, .Z(n_3582));
	notech_ao3 i_13073246(.A(n_59664), .B(in128[107]), .C(n_58881), .Z(n_3583
		));
	notech_ao4 i_19026519(.A(n_58795), .B(n_40081), .C(n_57585), .D(n_39785)
		, .Z(n_3584));
	notech_ao3 i_13173245(.A(n_59664), .B(in128[106]), .C(n_58881), .Z(n_3585
		));
	notech_ao4 i_18926518(.A(n_58797), .B(n_40080), .C(n_57587), .D(n_39783)
		, .Z(n_3586));
	notech_ao3 i_13273244(.A(n_59664), .B(in128[105]), .C(n_58881), .Z(n_3587
		));
	notech_ao4 i_18826517(.A(n_58797), .B(n_40079), .C(n_57587), .D(n_39781)
		, .Z(n_3588));
	notech_ao3 i_13373243(.A(n_59664), .B(in128[104]), .C(n_58882), .Z(n_3589
		));
	notech_ao4 i_18726516(.A(n_58797), .B(n_40078), .C(n_57587), .D(n_39779)
		, .Z(n_3590));
	notech_ao3 i_13473242(.A(n_59664), .B(in128[103]), .C(n_58882), .Z(n_3591
		));
	notech_ao4 i_18626515(.A(n_58797), .B(n_40077), .C(n_57587), .D(n_39777)
		, .Z(n_3592));
	notech_ao3 i_13573241(.A(n_59664), .B(in128[102]), .C(n_58882), .Z(n_3593
		));
	notech_ao4 i_18526514(.A(n_58797), .B(n_40076), .C(n_57587), .D(n_39775)
		, .Z(n_3594));
	notech_ao3 i_13673240(.A(n_59664), .B(in128[101]), .C(n_58881), .Z(n_3595
		));
	notech_ao4 i_18426513(.A(n_58797), .B(n_40075), .C(n_57587), .D(n_39773)
		, .Z(n_3596));
	notech_ao3 i_13773239(.A(n_59664), .B(in128[100]), .C(n_58881), .Z(n_3597
		));
	notech_ao4 i_18326512(.A(n_58797), .B(n_40074), .C(n_57587), .D(n_39771)
		, .Z(n_3598));
	notech_ao3 i_13873238(.A(n_59664), .B(in128[99]), .C(n_58873), .Z(n_3599
		));
	notech_ao4 i_18226511(.A(n_58797), .B(n_40073), .C(n_57587), .D(n_39769)
		, .Z(n_3600));
	notech_ao3 i_13973237(.A(n_59664), .B(in128[98]), .C(n_58868), .Z(n_3601
		));
	notech_ao4 i_18126510(.A(n_58797), .B(n_40072), .C(n_57587), .D(n_39767)
		, .Z(n_3602));
	notech_ao3 i_14073236(.A(n_59664), .B(in128[97]), .C(n_58868), .Z(n_3603
		));
	notech_ao4 i_18026509(.A(n_58797), .B(n_40071), .C(n_57587), .D(n_39765)
		, .Z(n_3604));
	notech_ao3 i_14173235(.A(n_59664), .B(in128[96]), .C(n_58868), .Z(n_3605
		));
	notech_ao4 i_17926508(.A(n_58795), .B(n_40070), .C(n_57585), .D(n_39763)
		, .Z(n_3606));
	notech_ao4 i_17826507(.A(n_58792), .B(n_40069), .C(n_57582), .D(n_39762)
		, .Z(n_3607));
	notech_ao3 i_14373233(.A(n_59663), .B(in128[94]), .C(n_58868), .Z(n_3608
		));
	notech_ao4 i_17726506(.A(n_58792), .B(n_40068), .C(n_57582), .D(n_39760)
		, .Z(n_3609));
	notech_ao3 i_14473232(.A(n_59663), .B(in128[93]), .C(n_58868), .Z(n_3610
		));
	notech_ao4 i_17626505(.A(n_58792), .B(n_40067), .C(n_57582), .D(n_39758)
		, .Z(n_3611));
	notech_ao4 i_17526504(.A(n_58792), .B(n_40066), .C(n_57582), .D(n_39757)
		, .Z(n_3612));
	notech_ao3 i_14673230(.A(n_59663), .B(in128[91]), .C(n_58868), .Z(n_3613
		));
	notech_ao4 i_17426503(.A(n_58792), .B(n_40065), .C(n_57582), .D(n_39755)
		, .Z(n_3614));
	notech_ao4 i_17326502(.A(n_58792), .B(n_40064), .C(n_57582), .D(n_39754)
		, .Z(n_3615));
	notech_ao4 i_17226501(.A(n_58792), .B(n_40063), .C(n_57582), .D(n_39753)
		, .Z(n_3616));
	notech_ao3 i_14973227(.A(n_59663), .B(in128[88]), .C(n_58868), .Z(n_3617
		));
	notech_ao4 i_17126500(.A(n_58792), .B(n_40062), .C(n_57582), .D(n_39751)
		, .Z(n_3618));
	notech_ao3 i_5873318(.A(n_59663), .B(in128[87]), .C(n_58872), .Z(n_3619)
		);
	notech_ao4 i_16926498(.A(n_58792), .B(n_40060), .C(n_57582), .D(n_39748)
		, .Z(n_3620));
	notech_ao4 i_16826497(.A(n_58792), .B(n_40059), .C(n_57582), .D(n_39747)
		, .Z(n_3621));
	notech_ao4 i_16726496(.A(n_58795), .B(n_40058), .C(n_57585), .D(n_39746)
		, .Z(n_3622));
	notech_ao4 i_16626495(.A(n_58795), .B(n_40057), .C(n_57585), .D(n_39745)
		, .Z(n_3623));
	notech_ao4 i_16526494(.A(n_58795), .B(n_40056), .C(n_57585), .D(n_39744)
		, .Z(n_3624));
	notech_ao4 i_16426493(.A(n_58795), .B(n_40055), .C(n_57585), .D(n_39743)
		, .Z(n_3625));
	notech_ao4 i_16326492(.A(n_58795), .B(n_40054), .C(n_57585), .D(n_39742)
		, .Z(n_3626));
	notech_ao3 i_6373313(.A(n_59663), .B(in128[79]), .C(n_58868), .Z(n_3627)
		);
	notech_ao4 i_16226491(.A(n_58792), .B(n_40053), .C(n_57582), .D(n_39740)
		, .Z(n_3628));
	notech_ao3 i_4473332(.A(n_59664), .B(in128[78]), .C(n_58868), .Z(n_3629)
		);
	notech_ao4 i_16126490(.A(n_58792), .B(n_40052), .C(n_57582), .D(n_39738)
		, .Z(n_3630));
	notech_ao3 i_1773359(.A(n_59664), .B(in128[77]), .C(n_58868), .Z(n_3631)
		);
	notech_ao4 i_16026489(.A(n_58792), .B(n_40051), .C(n_57582), .D(n_39736)
		, .Z(n_3632));
	notech_ao3 i_6073316(.A(n_59664), .B(in128[76]), .C(n_58864), .Z(n_3633)
		);
	notech_ao4 i_15926488(.A(n_58795), .B(n_40050), .C(n_57585), .D(n_39734)
		, .Z(n_3634));
	notech_ao3 i_4273334(.A(n_59663), .B(in128[75]), .C(n_58864), .Z(n_3635)
		);
	notech_ao4 i_15826487(.A(n_58795), .B(n_40049), .C(n_57585), .D(n_39732)
		, .Z(n_3636));
	notech_ao3 i_7273304(.A(n_59664), .B(in128[74]), .C(n_58864), .Z(n_3637)
		);
	notech_ao4 i_15726486(.A(n_58773), .B(n_40048), .C(n_57574), .D(n_39730)
		, .Z(n_3638));
	notech_ao3 i_3273344(.A(n_59664), .B(in128[73]), .C(n_58864), .Z(n_3639)
		);
	notech_ao4 i_15626485(.A(n_58773), .B(n_40047), .C(n_57563), .D(n_39728)
		, .Z(n_3640));
	notech_ao3 i_7673300(.A(n_59653), .B(in128[72]), .C(n_58864), .Z(n_3641)
		);
	notech_ao4 i_15526484(.A(n_58773), .B(n_40046), .C(n_57563), .D(n_39726)
		, .Z(n_3642));
	notech_ao3 i_5473322(.A(n_59647), .B(in128[71]), .C(n_58864), .Z(n_3643)
		);
	notech_ao4 i_15426483(.A(n_58773), .B(n_40045), .C(n_57563), .D(n_39724)
		, .Z(n_3644));
	notech_ao3 i_3673340(.A(n_59647), .B(in128[70]), .C(n_58868), .Z(n_3645)
		);
	notech_ao4 i_15326482(.A(n_58773), .B(n_40044), .C(n_57563), .D(n_39722)
		, .Z(n_3646));
	notech_ao3 i_1573361(.A(n_59647), .B(in128[69]), .C(n_58868), .Z(n_3647)
		);
	notech_ao4 i_15226481(.A(n_58770), .B(n_40043), .C(n_57563), .D(n_39720)
		, .Z(n_3648));
	notech_ao3 i_3873338(.A(n_59647), .B(in128[68]), .C(n_58868), .Z(n_3649)
		);
	notech_ao4 i_15126480(.A(n_58770), .B(n_40042), .C(n_57560), .D(n_39718)
		, .Z(n_3650));
	notech_ao3 i_8073296(.A(n_59647), .B(in128[67]), .C(n_58864), .Z(n_3651)
		);
	notech_ao4 i_15026479(.A(n_58770), .B(n_40041), .C(n_57560), .D(n_39716)
		, .Z(n_3652));
	notech_ao3 i_4073336(.A(n_59647), .B(in128[66]), .C(n_58868), .Z(n_3653)
		);
	notech_ao4 i_14926478(.A(n_58770), .B(n_40040), .C(n_57560), .D(n_39714)
		, .Z(n_3654));
	notech_ao3 i_3973337(.A(n_59652), .B(in128[65]), .C(n_58872), .Z(n_3655)
		);
	notech_ao4 i_14826477(.A(n_58770), .B(n_40039), .C(n_57563), .D(n_39712)
		, .Z(n_3656));
	notech_ao3 i_2873348(.A(n_59652), .B(in128[64]), .C(n_58873), .Z(n_3657)
		);
	notech_ao4 i_14626475(.A(n_58773), .B(n_40037), .C(n_57560), .D(n_39709)
		, .Z(n_3658));
	notech_ao3 i_6973307(.A(n_59652), .B(in128[62]), .C(n_58873), .Z(n_3659)
		);
	notech_ao4 i_14526474(.A(n_58773), .B(n_40036), .C(n_57563), .D(n_39707)
		, .Z(n_3660));
	notech_ao3 i_1673360(.A(n_59652), .B(in128[61]), .C(n_58873), .Z(n_3661)
		);
	notech_ao4 i_14426473(.A(n_58773), .B(n_40035), .C(n_57563), .D(n_39705)
		, .Z(n_3662));
	notech_ao3 i_6873308(.A(n_59652), .B(in128[60]), .C(n_58872), .Z(n_3663)
		);
	notech_ao4 i_14326472(.A(n_58775), .B(n_40034), .C(n_57563), .D(n_39703)
		, .Z(n_3664));
	notech_ao3 i_6773309(.A(n_59652), .B(in128[59]), .C(n_58873), .Z(n_3665)
		);
	notech_ao4 i_14226471(.A(n_58773), .B(n_40033), .C(n_57565), .D(n_39701)
		, .Z(n_3666));
	notech_ao3 i_4573331(.A(n_59647), .B(in128[58]), .C(n_58873), .Z(n_3667)
		);
	notech_ao4 i_14126470(.A(n_58773), .B(n_40032), .C(n_57565), .D(n_39699)
		, .Z(n_3668));
	notech_ao3 i_6673310(.A(n_59642), .B(in128[57]), .C(n_58873), .Z(n_3669)
		);
	notech_ao4 i_14026469(.A(n_58773), .B(n_40031), .C(n_57563), .D(n_39697)
		, .Z(n_3670));
	notech_ao3 i_6573311(.A(n_59642), .B(in128[56]), .C(n_58873), .Z(n_3671)
		);
	notech_ao4 i_13726466(.A(n_58773), .B(n_40028), .C(n_57563), .D(n_39692)
		, .Z(n_3672));
	notech_ao3 i_1873358(.A(n_59642), .B(in128[53]), .C(n_58873), .Z(n_3673)
		);
	notech_ao4 i_13626465(.A(n_58773), .B(n_40027), .C(n_57563), .D(n_39690)
		, .Z(n_3674));
	notech_ao3 i_4773329(.A(n_59642), .B(in128[52]), .C(n_58873), .Z(n_3675)
		);
	notech_ao4 i_13526464(.A(n_58773), .B(n_40026), .C(n_57563), .D(n_39688)
		, .Z(n_3676));
	notech_ao3 i_7173305(.A(n_59642), .B(in128[51]), .C(n_58873), .Z(n_3677)
		);
	notech_ao4 i_13426463(.A(n_58770), .B(n_40025), .C(n_57563), .D(n_39686)
		, .Z(n_3678));
	notech_ao3 i_7373303(.A(n_59642), .B(in128[50]), .C(n_58872), .Z(n_3679)
		);
	notech_ao4 i_13326462(.A(n_58768), .B(n_40024), .C(n_57560), .D(n_39684)
		, .Z(n_3680));
	notech_ao3 i_8173295(.A(n_59647), .B(in128[49]), .C(n_58872), .Z(n_3681)
		);
	notech_ao4 i_13226461(.A(n_58768), .B(n_40023), .C(n_57558), .D(n_39682)
		, .Z(n_3682));
	notech_ao3 i_7873298(.A(n_59647), .B(in128[48]), .C(n_58872), .Z(n_3683)
		);
	notech_ao4 i_13126460(.A(n_58768), .B(n_40022), .C(n_57558), .D(n_39680)
		, .Z(n_3684));
	notech_ao3 i_5773319(.A(n_59647), .B(in128[47]), .C(n_58872), .Z(n_3685)
		);
	notech_ao4 i_12926458(.A(n_58768), .B(n_40020), .C(n_57558), .D(n_39676)
		, .Z(n_3686));
	notech_ao3 i_1973357(.A(n_59642), .B(in128[45]), .C(n_58872), .Z(n_3687)
		);
	notech_ao4 i_12826457(.A(n_58768), .B(n_40019), .C(n_57558), .D(n_39674)
		, .Z(n_3688));
	notech_ao4 i_12726456(.A(n_58768), .B(n_40018), .C(n_57558), .D(n_39673)
		, .Z(n_3689));
	notech_ao4 i_12526454(.A(n_58768), .B(n_40016), .C(n_57558), .D(n_39671)
		, .Z(n_3690));
	notech_ao4 i_12426453(.A(n_58768), .B(n_40015), .C(n_57558), .D(n_39670)
		, .Z(n_3691));
	notech_ao4 i_12026449(.A(n_58768), .B(n_40011), .C(n_57558), .D(n_39663)
		, .Z(n_3692));
	notech_ao3 i_7473302(.A(n_59647), .B(in128[36]), .C(n_58872), .Z(n_3693)
		);
	notech_ao4 i_11826447(.A(n_58768), .B(n_40009), .C(n_57558), .D(n_39658)
		, .Z(n_3694));
	notech_ao3 i_5973317(.A(n_59647), .B(in128[34]), .C(n_58872), .Z(n_3695)
		);
	notech_ao4 i_11326442(.A(n_58770), .B(n_40004), .C(n_57558), .D(n_39646)
		, .Z(n_3696));
	notech_ao4 i_7026399(.A(n_58770), .B(n_40166), .C(n_57560), .D(n_39575),
		 .Z(n_3697));
	notech_ao4 i_6826397(.A(n_58770), .B(n_40107), .C(n_57560), .D(n_39572),
		 .Z(n_3698));
	notech_ao4 i_6726396(.A(n_58770), .B(n_40108), .C(n_57560), .D(n_39571),
		 .Z(n_3699));
	notech_ao4 i_6626395(.A(n_58770), .B(n_40109), .C(n_57560), .D(n_39569),
		 .Z(n_3700));
	notech_ao4 i_6526394(.A(n_58768), .B(n_40110), .C(n_57560), .D(n_39568),
		 .Z(n_3701));
	notech_ao4 i_6426393(.A(n_58768), .B(n_40111), .C(n_57560), .D(n_39567),
		 .Z(n_3702));
	notech_ao3 i_15473222(.A(n_59652), .B(\to_acu2_0[63] ), .C(n_58872), .Z(n_3703
		));
	notech_ao4 i_6326392(.A(n_58770), .B(n_40165), .C(n_57558), .D(n_39565),
		 .Z(n_3704));
	notech_ao3 i_10473272(.A(n_59653), .B(\to_acu2_0[62] ), .C(n_58872), .Z(n_3705
		));
	notech_ao4 i_6226391(.A(n_58770), .B(n_40145), .C(n_57560), .D(n_39563),
		 .Z(n_3706));
	notech_ao3 i_9173285(.A(n_59653), .B(\to_acu2_0[61] ), .C(n_58872), .Z(n_3707
		));
	notech_ao4 i_6126390(.A(n_58770), .B(n_40112), .C(n_57560), .D(n_39561),
		 .Z(n_3708));
	notech_ao3 i_15573221(.A(n_59653), .B(\to_acu2_0[60] ), .C(n_58872), .Z(n_3709
		));
	notech_ao4 i_6026389(.A(n_58775), .B(n_40129), .C(n_57560), .D(n_39559),
		 .Z(n_3710));
	notech_ao3 i_9073286(.A(n_59653), .B(\to_acu2_0[59] ), .C(n_58844), .Z(n_3711
		));
	notech_ao4 i_5926388(.A(n_58781), .B(n_40122), .C(n_57571), .D(n_39557),
		 .Z(n_3712));
	notech_ao3 i_5073326(.A(n_59653), .B(\to_acu2_0[58] ), .C(n_58810), .Z(n_3713
		));
	notech_ao4 i_5826387(.A(n_58781), .B(n_40123), .C(n_57571), .D(n_39555),
		 .Z(n_3714));
	notech_ao3 i_3473342(.A(n_59653), .B(\to_acu2_0[57] ), .C(n_58810), .Z(n_3715
		));
	notech_ao4 i_5726386(.A(n_58781), .B(n_40120), .C(n_57571), .D(n_39553),
		 .Z(n_3716));
	notech_ao3 i_9273284(.A(n_59653), .B(\to_acu2_0[56] ), .C(n_58810), .Z(n_3717
		));
	notech_ao4 i_5626385(.A(n_58781), .B(n_40127), .C(n_57571), .D(n_39551),
		 .Z(n_3718));
	notech_ao3 i_4373333(.A(n_59653), .B(\to_acu2_0[55] ), .C(n_58810), .Z(n_3719
		));
	notech_ao4 i_5526384(.A(n_58781), .B(n_40128), .C(n_57571), .D(n_39549),
		 .Z(n_3720));
	notech_ao3 i_2373353(.A(n_59653), .B(\to_acu2_0[54] ), .C(n_58810), .Z(n_3721
		));
	notech_ao4 i_5426383(.A(n_58779), .B(n_40126), .C(n_57569), .D(n_39547),
		 .Z(n_3722));
	notech_ao3 i_4973327(.A(n_59653), .B(\to_acu2_0[53] ), .C(n_58810), .Z(n_3723
		));
	notech_ao4 i_5326382(.A(n_58779), .B(n_40124), .C(n_57569), .D(n_39545),
		 .Z(n_3724));
	notech_ao3 i_3373343(.A(n_59653), .B(\to_acu2_0[52] ), .C(n_58810), .Z(n_3725
		));
	notech_ao4 i_5226381(.A(n_58779), .B(n_40125), .C(n_57569), .D(n_39543),
		 .Z(n_3726));
	notech_ao3 i_2673350(.A(n_59653), .B(\to_acu2_0[51] ), .C(n_58810), .Z(n_3727
		));
	notech_ao4 i_5126380(.A(n_58779), .B(n_40121), .C(n_57569), .D(n_39540),
		 .Z(n_3728));
	notech_ao3 i_5173325(.A(n_59653), .B(\to_acu2_0[50] ), .C(n_58810), .Z(n_3729
		));
	notech_ao4 i_5026379(.A(n_58779), .B(n_40113), .C(n_57569), .D(n_39538),
		 .Z(n_3730));
	notech_ao3 i_15673220(.A(n_59652), .B(\to_acu2_0[49] ), .C(n_58810), .Z(n_3731
		));
	notech_ao4 i_4926378(.A(n_58781), .B(n_40131), .C(n_57571), .D(n_39535),
		 .Z(n_3732));
	notech_ao3 i_8973287(.A(n_59652), .B(\to_acu2_0[48] ), .C(n_58810), .Z(n_3733
		));
	notech_ao4 i_4826377(.A(n_58781), .B(n_40144), .C(n_57571), .D(n_39533),
		 .Z(n_3734));
	notech_ao3 i_7773299(.A(n_59652), .B(\to_acu2_0[47] ), .C(n_58812), .Z(n_3735
		));
	notech_ao4 i_4726376(.A(n_58781), .B(n_40142), .C(n_57571), .D(n_39530),
		 .Z(n_3736));
	notech_ao3 i_5273324(.A(n_59652), .B(\to_acu2_0[46] ), .C(n_58812), .Z(n_3737
		));
	notech_ao4 i_4626375(.A(n_58784), .B(n_40143), .C(n_57574), .D(n_39528),
		 .Z(n_3738));
	notech_ao3 i_3573341(.A(n_59652), .B(\to_acu2_0[45] ), .C(n_58812), .Z(n_3739
		));
	notech_ao4 i_4526374(.A(n_58781), .B(n_40141), .C(n_57571), .D(n_39525),
		 .Z(n_3740));
	notech_ao3 i_2773349(.A(n_59652), .B(\to_acu2_0[44] ), .C(n_58812), .Z(n_3741
		));
	notech_ao4 i_4426373(.A(n_58781), .B(n_40139), .C(n_57571), .D(n_39523),
		 .Z(n_3742));
	notech_ao3 i_2473352(.A(n_59652), .B(\to_acu2_0[43] ), .C(n_58812), .Z(n_3743
		));
	notech_ao4 i_4326372(.A(n_58781), .B(n_40140), .C(n_57571), .D(n_39520),
		 .Z(n_3744));
	notech_ao3 i_2173355(.A(n_59652), .B(\to_acu2_0[42] ), .C(n_58812), .Z(n_3745
		));
	notech_ao4 i_4226371(.A(n_58781), .B(n_40138), .C(n_57571), .D(n_39518),
		 .Z(n_3746));
	notech_ao3 i_11073266(.A(n_59653), .B(\to_acu2_0[41] ), .C(n_58810), .Z(n_3747
		));
	notech_ao4 i_4126370(.A(n_58781), .B(n_40136), .C(n_57571), .D(n_39515),
		 .Z(n_3748));
	notech_ao3 i_16373213(.A(n_59652), .B(\to_acu2_0[40] ), .C(n_58810), .Z(n_3749
		));
	notech_ao4 i_3926368(.A(n_58781), .B(n_40137), .C(n_57571), .D(n_39512),
		 .Z(n_3750));
	notech_ao3 i_10973267(.A(n_59652), .B(\to_acu2_0[38] ), .C(n_58810), .Z(n_3751
		));
	notech_ao4 i_3826367(.A(n_58779), .B(n_40134), .C(n_57569), .D(n_39509),
		 .Z(n_3752));
	notech_ao3 i_10873268(.A(n_59652), .B(\to_acu2_0[37] ), .C(n_58812), .Z(n_3753
		));
	notech_ao4 i_3726366(.A(n_58775), .B(n_40135), .C(n_57565), .D(n_39507),
		 .Z(n_3754));
	notech_ao3 i_10773269(.A(n_59619), .B(\to_acu2_0[36] ), .C(n_58812), .Z(n_3755
		));
	notech_ao4 i_3626365(.A(n_58775), .B(n_40132), .C(n_57565), .D(n_39504),
		 .Z(n_3756));
	notech_ao3 i_10673270(.A(n_59584), .B(\to_acu2_0[35] ), .C(n_58810), .Z(n_3757
		));
	notech_ao4 i_3526364(.A(n_58775), .B(n_40133), .C(n_57565), .D(n_39502),
		 .Z(n_3758));
	notech_ao3 i_10573271(.A(n_59584), .B(\to_acu2_0[34] ), .C(n_58821), .Z(n_3759
		));
	notech_ao4 i_3426363(.A(n_58775), .B(n_40114), .C(n_57565), .D(n_39499),
		 .Z(n_3760));
	notech_ao3 i_15773219(.A(n_59584), .B(\to_acu2_0[33] ), .C(n_58821), .Z(n_3761
		));
	notech_ao4 i_3326362(.A(n_58775), .B(n_40115), .C(n_57565), .D(n_39497),
		 .Z(n_3762));
	notech_ao3 i_15873218(.A(n_59584), .B(\to_acu2_0[32] ), .C(n_58821), .Z(n_3763
		));
	notech_ao4 i_3226361(.A(n_58775), .B(n_40116), .C(n_57565), .D(n_39494),
		 .Z(n_3764));
	notech_ao3 i_15973217(.A(n_59584), .B(\to_acu2_0[31] ), .C(n_58821), .Z(n_3765
		));
	notech_ao4 i_3126360(.A(n_58775), .B(n_40117), .C(n_57565), .D(n_39492),
		 .Z(n_3766));
	notech_ao3 i_16073216(.A(n_59584), .B(\to_acu2_0[30] ), .C(n_58821), .Z(n_3767
		));
	notech_ao4 i_3026359(.A(n_58775), .B(n_40118), .C(n_57565), .D(n_39489),
		 .Z(n_3768));
	notech_ao3 i_16173215(.A(n_59584), .B(\to_acu2_0[29] ), .C(n_58825), .Z(n_3769
		));
	notech_ao4 i_2926358(.A(n_58775), .B(n_40163), .C(n_57565), .D(n_39487),
		 .Z(n_3770));
	notech_ao4 i_2826357(.A(n_58775), .B(n_40159), .C(n_57565), .D(n_39485),
		 .Z(n_3771));
	notech_ao4 i_2726356(.A(n_58779), .B(n_40160), .C(n_57569), .D(n_39483),
		 .Z(n_3772));
	notech_ao4 i_2626355(.A(n_58779), .B(n_40162), .C(n_57569), .D(n_39481),
		 .Z(n_3773));
	notech_ao4 i_2526354(.A(n_58779), .B(n_40161), .C(n_57569), .D(n_39479),
		 .Z(n_3774));
	notech_ao4 i_2426353(.A(n_58779), .B(n_40157), .C(n_57569), .D(n_39477),
		 .Z(n_3775));
	notech_ao4 i_2326352(.A(n_58779), .B(n_40158), .C(n_57569), .D(n_39475),
		 .Z(n_3776));
	notech_ao4 i_2226351(.A(n_58775), .B(n_40156), .C(n_57565), .D(n_39473),
		 .Z(n_3777));
	notech_ao3 i_10073276(.A(n_59584), .B(\to_acu2_0[21] ), .C(n_58825), .Z(n_3778
		));
	notech_ao4 i_2126350(.A(n_58775), .B(n_40155), .C(n_57565), .D(n_39470),
		 .Z(n_3779));
	notech_ao3 i_8473292(.A(n_59584), .B(\to_acu2_0[20] ), .C(n_58825), .Z(n_3780
		));
	notech_ao4 i_1926348(.A(n_58779), .B(n_40153), .C(n_57569), .D(n_39465),
		 .Z(n_3781));
	notech_ao3 i_9973277(.A(n_59584), .B(\to_acu2_0[18] ), .C(n_58825), .Z(n_3782
		));
	notech_ao4 i_1826347(.A(n_58779), .B(n_40152), .C(n_57569), .D(n_39463),
		 .Z(n_3783));
	notech_ao3 i_9873278(.A(n_59584), .B(\to_acu2_0[17] ), .C(n_58825), .Z(n_3784
		));
	notech_ao4 i_1726346(.A(n_58779), .B(n_40164), .C(n_57569), .D(n_39460),
		 .Z(n_3785));
	notech_ao3 i_4173335(.A(n_59584), .B(\to_acu2_0[16] ), .C(n_58825), .Z(n_3786
		));
	notech_ao4 i_1626345(.A(n_58689), .B(n_40149), .C(n_57479), .D(n_39458),
		 .Z(n_3787));
	notech_ao3 i_9773279(.A(n_59584), .B(\to_acu2_0[15] ), .C(n_58821), .Z(n_3788
		));
	notech_ao4 i_1526344(.A(n_58689), .B(n_40150), .C(n_57479), .D(n_39455),
		 .Z(n_3789));
	notech_ao4 i_1426343(.A(n_58689), .B(n_40151), .C(n_57479), .D(n_39453),
		 .Z(n_3790));
	notech_ao4 i_1326342(.A(n_58689), .B(n_40154), .C(n_57479), .D(n_39451),
		 .Z(n_3791));
	notech_ao4 i_1226341(.A(n_58689), .B(n_40168), .C(n_57479), .D(n_39449),
		 .Z(n_3792));
	notech_ao3 i_9573281(.A(n_59579), .B(\to_acu2_0[11] ), .C(n_58821), .Z(n_3793
		));
	notech_ao4 i_1126340(.A(n_58689), .B(n_40169), .C(n_57479), .D(n_39447),
		 .Z(n_3794));
	notech_ao3 i_9473282(.A(n_59579), .B(\to_acu2_0[10] ), .C(n_58810), .Z(n_3795
		));
	notech_ao4 i_1026339(.A(n_58689), .B(n_40170), .C(n_57479), .D(n_39444),
		 .Z(n_3796));
	notech_ao3 i_4873328(.A(n_59579), .B(\to_acu2_0[9] ), .C(n_58810), .Z(n_3797
		));
	notech_ao4 i_926338(.A(n_58689), .B(n_40167), .C(n_57479), .D(n_39442), 
		.Z(n_3798));
	notech_ao4 i_826337(.A(n_58689), .B(n_40146), .C(n_57479), .D(n_39440), 
		.Z(n_3799));
	notech_ao3 i_16573211(.A(n_59579), .B(\to_acu2_0[7] ), .C(n_58810), .Z(n_3800
		));
	notech_ao4 i_726336(.A(n_58689), .B(n_40119), .C(n_57479), .D(n_39437), 
		.Z(n_3801));
	notech_ao3 i_16273214(.A(n_59579), .B(\to_acu2_0[6] ), .C(n_58821), .Z(n_3802
		));
	notech_ao4 i_626335(.A(n_58691), .B(n_40130), .C(n_57481), .D(n_39435), 
		.Z(n_3803));
	notech_ao3 i_2973347(.A(n_59579), .B(\to_acu2_0[5] ), .C(n_58821), .Z(n_3804
		));
	notech_ao4 i_526334(.A(n_58691), .B(n_40209), .C(n_57481), .D(n_39432), 
		.Z(n_3805));
	notech_ao4 i_426333(.A(n_58691), .B(n_40212), .C(n_57481), .D(n_39430), 
		.Z(n_3806));
	notech_ao3 i_16673210(.A(n_59584), .B(\to_acu2_0[3] ), .C(n_58821), .Z(n_3807
		));
	notech_ao4 i_326332(.A(n_58691), .B(n_40147), .C(n_57481), .D(n_39428), 
		.Z(n_3808));
	notech_ao4 i_226331(.A(n_58691), .B(n_40148), .C(n_57481), .D(n_39426), 
		.Z(n_3809));
	notech_ao3 i_6173315(.A(n_59584), .B(\to_acu2_0[1] ), .C(n_58821), .Z(n_3810
		));
	notech_ao4 i_126330(.A(n_58689), .B(n_40214), .C(n_57479), .D(n_39423), 
		.Z(n_3811));
	notech_ao4 i_123152(.A(n_40175), .B(n_39249), .C(n_57479), .D(n_38674), 
		.Z(n_3812));
	notech_and3 i_773369(.A(n_250691353), .B(n_38431), .C(n_38428), .Z(n_3813
		));
	notech_nand2 i_925660(.A(n_59692), .B(n_1620), .Z(n_3234));
	notech_nand2 i_1125662(.A(n_59692), .B(n_1619), .Z(n_3233));
	notech_nand2 i_1225663(.A(n_59692), .B(n_1618), .Z(n_3232));
	notech_nand2 i_1325664(.A(n_59692), .B(n_1617), .Z(n_3231));
	notech_or2 i_528(.A(n_5717), .B(n_251191358), .Z(n_9089));
	notech_nao3 i_166(.A(db67), .B(n_41571), .C(n_5674), .Z(n_5304));
	notech_nand2 i_22(.A(n_2864), .B(n_40171), .Z(n_5674));
	notech_nao3 i_27(.A(db67), .B(n_59584), .C(n_2849), .Z(n_5726));
	notech_ao4 i_65995(.A(n_2140), .B(n_2874), .C(n_2872), .D(n_39849), .Z(n_2058
		));
	notech_ao3 i_427204(.A(n_59579), .B(\nbus_12535[3] ), .C(n_58821), .Z(n_2057
		));
	notech_nand2 i_1092391(.A(n_40193), .B(pc_req), .Z(n_2055));
	notech_ao3 i_240(.A(n_59579), .B(\to_acu2_0[77] ), .C(n_58821), .Z(n_2054
		));
	notech_ao3 i_241(.A(n_59584), .B(in128[3]), .C(n_58812), .Z(n_2053));
	notech_ao3 i_242(.A(n_59584), .B(in128[4]), .C(n_58803), .Z(n_2052));
	notech_ao3 i_243(.A(n_59595), .B(in128[5]), .C(n_58803), .Z(n_2051));
	notech_ao3 i_244(.A(n_59595), .B(in128[6]), .C(n_58803), .Z(n_2050));
	notech_ao3 i_245(.A(n_59595), .B(in128[7]), .C(n_58803), .Z(n_2049));
	notech_ao3 i_289(.A(n_59595), .B(sib_dec), .C(n_58803), .Z(n_2048));
	notech_ao3 i_290(.A(n_59595), .B(mod_dec), .C(n_58803), .Z(n_2047));
	notech_nor2 i_307(.A(n_2163), .B(n_58689), .Z(n_2046));
	notech_nor2 i_308(.A(n_2176), .B(n_58689), .Z(n_2045));
	notech_nor2 i_309(.A(n_2186), .B(n_58691), .Z(n_2044));
	notech_nor2 i_310(.A(n_2196), .B(n_58689), .Z(n_2043));
	notech_nor2 i_311(.A(n_2206), .B(n_58685), .Z(n_2042));
	notech_ao3 i_358(.A(n_59595), .B(\to_acu2_0[80] ), .C(n_58801), .Z(n_2041
		));
	notech_ao3 i_360(.A(n_59595), .B(\to_acu2_0[75] ), .C(n_58801), .Z(n_2040
		));
	notech_ao3 i_361(.A(n_59595), .B(\to_acu2_0[70] ), .C(n_58801), .Z(n_2039
		));
	notech_ao3 i_362(.A(n_59595), .B(\to_acu2_0[79] ), .C(n_58803), .Z(n_2038
		));
	notech_ao3 i_363(.A(n_59595), .B(\to_acu2_0[78] ), .C(n_58801), .Z(n_2037
		));
	notech_ao3 i_364(.A(n_59595), .B(\to_acu2_0[76] ), .C(n_58803), .Z(n_2036
		));
	notech_ao3 i_365(.A(n_59595), .B(\to_acu2_0[72] ), .C(n_58803), .Z(n_2035
		));
	notech_ao3 i_366(.A(n_59590), .B(\to_acu2_0[68] ), .C(n_58803), .Z(n_2034
		));
	notech_ao3 i_375(.A(n_59590), .B(\to_acu2_0[19] ), .C(n_58803), .Z(n_2033
		));
	notech_ao3 i_378(.A(n_59590), .B(n_57713), .C(n_58803), .Z(n_2032));
	notech_ao3 i_379(.A(n_59590), .B(in128[23]), .C(n_58803), .Z(n_2031));
	notech_ao3 i_380(.A(n_59584), .B(in128[27]), .C(n_58803), .Z(n_2030));
	notech_ao3 i_382(.A(n_59584), .B(in128[28]), .C(n_58803), .Z(n_2029));
	notech_ao3 i_383(.A(n_59590), .B(in128[16]), .C(n_58803), .Z(n_2028));
	notech_nand2 i_1525666(.A(n_59692), .B(n_1616), .Z(n_3230));
	notech_ao3 i_390(.A(n_59590), .B(in128[2]), .C(n_58803), .Z(n_2027));
	notech_ao3 i_391(.A(n_59590), .B(in128[20]), .C(n_58803), .Z(n_2026));
	notech_ao3 i_393(.A(n_59590), .B(in128[33]), .C(n_58801), .Z(n_2025));
	notech_ao3 i_394(.A(n_59590), .B(in128[32]), .C(n_58812), .Z(n_2024));
	notech_ao3 i_398(.A(n_59590), .B(in128[37]), .C(n_58812), .Z(n_2023));
	notech_ao3 i_401(.A(n_59590), .B(in128[38]), .C(n_58812), .Z(n_2022));
	notech_ao3 i_404(.A(n_59579), .B(in128[42]), .C(n_58801), .Z(n_2021));
	notech_ao3 i_407(.A(n_59568), .B(in128[35]), .C(n_58801), .Z(n_2020));
	notech_ao3 i_414(.A(n_59568), .B(in128[31]), .C(n_58812), .Z(n_2019));
	notech_ao3 i_424(.A(n_59568), .B(in128[22]), .C(n_58812), .Z(n_2018));
	notech_ao3 i_426(.A(n_59568), .B(in128[25]), .C(n_58812), .Z(n_2017));
	notech_ao3 i_427(.A(n_59568), .B(in128[8]), .C(n_58812), .Z(n_2016));
	notech_ao3 i_428(.A(n_59568), .B(in128[14]), .C(n_58812), .Z(n_2015));
	notech_ao3 i_429(.A(n_59573), .B(in128[9]), .C(n_58812), .Z(n_2014));
	notech_ao3 i_431(.A(n_59573), .B(\to_acu2_0[73] ), .C(n_58801), .Z(n_2013
		));
	notech_ao3 i_433(.A(n_59573), .B(in128[39]), .C(n_58801), .Z(n_2012));
	notech_ao3 i_435(.A(n_59568), .B(in128[18]), .C(n_58801), .Z(n_2011));
	notech_nand2 i_1625667(.A(n_59692), .B(n_1615), .Z(n_3229));
	notech_ao3 i_439(.A(n_59573), .B(\to_acu2_0[71] ), .C(n_58801), .Z(n_2010
		));
	notech_ao3 i_441(.A(n_59573), .B(in128[30]), .C(n_58801), .Z(n_2009));
	notech_ao3 i_444(.A(n_59568), .B(in128[46]), .C(n_58801), .Z(n_2008));
	notech_ao3 i_448(.A(n_59568), .B(\to_acu2_0[74] ), .C(n_58801), .Z(n_2007
		));
	notech_ao3 i_453(.A(n_59568), .B(in128[19]), .C(n_58801), .Z(n_2006));
	notech_ao3 i_455(.A(n_59568), .B(in128[17]), .C(n_58801), .Z(n_2005));
	notech_ao3 i_463(.A(n_59568), .B(in128[13]), .C(n_58801), .Z(n_2004));
	notech_ao3 i_465(.A(n_59568), .B(in128[26]), .C(n_58801), .Z(n_2003));
	notech_ao3 i_470(.A(n_59568), .B(in128[0]), .C(n_58836), .Z(n_2002));
	notech_nand2 i_1725668(.A(n_59692), .B(n_1614), .Z(n_3228));
	notech_ao3 i_471(.A(n_59568), .B(in128[21]), .C(n_58836), .Z(n_2001));
	notech_ao3 i_482(.A(n_59568), .B(in128[12]), .C(n_58836), .Z(n_2000));
	notech_ao3 i_483(.A(n_59568), .B(in128[15]), .C(n_58836), .Z(n_1999));
	notech_ao3 i_490(.A(n_59568), .B(in128[11]), .C(n_58836), .Z(n_1998));
	notech_ao3 i_491(.A(n_59568), .B(in128[24]), .C(n_58836), .Z(n_1997));
	notech_and2 i_199(.A(twobyte), .B(n_40171), .Z(n_1996));
	notech_nand2 i_1825669(.A(n_59692), .B(n_1613), .Z(n_3227));
	notech_nand2 i_1925670(.A(n_59692), .B(n_1612), .Z(n_3226));
	notech_ao4 i_1(.A(n_2833), .B(n_38415), .C(n_2834), .D(n_38661), .Z(n_1995
		));
	notech_nand2 i_6350(.A(idx_deco[1]), .B(n_38656), .Z(n_5415));
	notech_and2 i_95610216(.A(\to_acu2_0[0] ), .B(\to_acu2_0[1] ), .Z(n_5717
		));
	notech_nand2 i_2025671(.A(n_59693), .B(n_1611), .Z(n_3225));
	notech_ao3 i_327203(.A(n_59568), .B(\nbus_12535[2] ), .C(n_58840), .Z(n_45035
		));
	notech_ao3 i_285(.A(n_59573), .B(in128[127]), .C(n_58840), .Z(n_48359)
		);
	notech_ao3 i_63(.A(n_59579), .B(udeco[62]), .C(n_58840), .Z(n_42534));
	notech_ao3 i_64(.A(n_59579), .B(udeco[63]), .C(n_58836), .Z(n_42540));
	notech_ao3 i_66(.A(n_59579), .B(udeco[65]), .C(n_58840), .Z(n_42552));
	notech_ao3 i_67(.A(n_59573), .B(udeco[66]), .C(n_58835), .Z(n_42558));
	notech_ao3 i_69(.A(n_59579), .B(udeco[68]), .C(n_58836), .Z(n_42570));
	notech_ao3 i_70(.A(n_59579), .B(udeco[69]), .C(n_58835), .Z(n_42576));
	notech_ao3 i_71(.A(n_59579), .B(udeco[70]), .C(n_58835), .Z(n_42582));
	notech_ao3 i_72(.A(n_59579), .B(udeco[71]), .C(n_58835), .Z(n_42588));
	notech_ao3 i_74(.A(n_59579), .B(udeco[73]), .C(n_58836), .Z(n_42600));
	notech_ao3 i_76(.A(n_59579), .B(udeco[75]), .C(n_58836), .Z(n_42612));
	notech_ao3 i_77(.A(n_59579), .B(udeco[76]), .C(n_58836), .Z(n_42618));
	notech_ao3 i_78(.A(n_59579), .B(udeco[77]), .C(n_58836), .Z(n_42624));
	notech_ao3 i_79(.A(n_59573), .B(udeco[78]), .C(n_58836), .Z(n_42630));
	notech_ao3 i_80(.A(n_59573), .B(udeco[79]), .C(n_58836), .Z(n_42636));
	notech_ao3 i_81(.A(n_59573), .B(udeco[80]), .C(n_58840), .Z(n_42642));
	notech_ao3 i_82(.A(n_59573), .B(udeco[81]), .C(n_58844), .Z(n_42648));
	notech_ao3 i_83(.A(n_59573), .B(udeco[82]), .C(n_58844), .Z(n_42654));
	notech_ao3 i_84(.A(n_59573), .B(udeco[83]), .C(n_58844), .Z(n_42660));
	notech_ao3 i_85(.A(n_59573), .B(udeco[84]), .C(n_58844), .Z(n_42666));
	notech_ao3 i_86(.A(n_59573), .B(udeco[85]), .C(n_58844), .Z(n_42672));
	notech_ao3 i_87(.A(n_59573), .B(udeco[86]), .C(n_58844), .Z(n_42678));
	notech_ao3 i_88(.A(n_59573), .B(udeco[87]), .C(n_58844), .Z(n_42684));
	notech_ao3 i_89(.A(n_59573), .B(udeco[88]), .C(n_58844), .Z(n_42690));
	notech_ao3 i_90(.A(n_59573), .B(udeco[89]), .C(n_58844), .Z(n_42696));
	notech_ao3 i_91(.A(n_59573), .B(udeco[90]), .C(n_58844), .Z(n_42702));
	notech_ao3 i_92(.A(n_59595), .B(udeco[91]), .C(n_58844), .Z(n_42708));
	notech_ao3 i_93(.A(n_59608), .B(udeco[92]), .C(n_58840), .Z(n_42714));
	notech_ao3 i_94(.A(n_59608), .B(udeco[93]), .C(n_58840), .Z(n_42720));
	notech_ao3 i_95(.A(n_59608), .B(udeco[94]), .C(n_58840), .Z(n_42726));
	notech_ao3 i_96(.A(n_59608), .B(udeco[95]), .C(n_58840), .Z(n_42732));
	notech_ao3 i_97(.A(n_59608), .B(udeco[96]), .C(n_58840), .Z(n_42738));
	notech_ao3 i_98(.A(n_59608), .B(udeco[97]), .C(n_58840), .Z(n_42744));
	notech_ao3 i_99(.A(n_59613), .B(udeco[98]), .C(n_58844), .Z(n_42750));
	notech_ao3 i_100(.A(n_59613), .B(udeco[99]), .C(n_58844), .Z(n_42756));
	notech_ao3 i_101(.A(n_59613), .B(udeco[100]), .C(n_58840), .Z(n_42762)
		);
	notech_ao3 i_102(.A(n_59613), .B(udeco[101]), .C(n_58840), .Z(n_42768)
		);
	notech_ao3 i_103(.A(n_59613), .B(udeco[102]), .C(n_58840), .Z(n_42774)
		);
	notech_ao3 i_105(.A(n_59613), .B(udeco[104]), .C(n_58835), .Z(n_42786)
		);
	notech_ao3 i_106(.A(n_59608), .B(udeco[105]), .C(n_58826), .Z(n_42792)
		);
	notech_ao3 i_107(.A(n_59608), .B(udeco[106]), .C(n_58826), .Z(n_42798)
		);
	notech_ao3 i_108(.A(n_59608), .B(udeco[107]), .C(n_58826), .Z(n_42804)
		);
	notech_ao3 i_109(.A(n_59608), .B(udeco[108]), .C(n_58826), .Z(n_42810)
		);
	notech_ao3 i_110(.A(n_59607), .B(udeco[109]), .C(n_58826), .Z(n_42816)
		);
	notech_ao3 i_111(.A(n_59608), .B(udeco[110]), .C(n_58826), .Z(n_42822)
		);
	notech_ao3 i_112(.A(n_59608), .B(udeco[111]), .C(n_58826), .Z(n_42828)
		);
	notech_ao3 i_113(.A(n_59608), .B(udeco[112]), .C(n_58826), .Z(n_42834)
		);
	notech_ao3 i_114(.A(n_59608), .B(udeco[113]), .C(n_58826), .Z(n_42840)
		);
	notech_ao3 i_115(.A(n_59608), .B(udeco[114]), .C(n_58826), .Z(n_42846)
		);
	notech_ao3 i_116(.A(n_59608), .B(udeco[115]), .C(n_58826), .Z(n_42852)
		);
	notech_ao3 i_117(.A(n_59608), .B(udeco[116]), .C(n_58825), .Z(n_42858)
		);
	notech_ao3 i_118(.A(n_59608), .B(udeco[117]), .C(n_58825), .Z(n_42864)
		);
	notech_ao3 i_119(.A(n_59613), .B(udeco[118]), .C(n_58825), .Z(n_42870)
		);
	notech_ao3 i_120(.A(n_59618), .B(udeco[119]), .C(n_58825), .Z(n_42876)
		);
	notech_ao3 i_121(.A(n_59618), .B(udeco[120]), .C(n_58825), .Z(n_42882)
		);
	notech_ao3 i_122(.A(n_59618), .B(udeco[121]), .C(n_58825), .Z(n_42888)
		);
	notech_ao3 i_123(.A(n_59618), .B(udeco[122]), .C(n_58826), .Z(n_42894)
		);
	notech_ao3 i_124(.A(n_59618), .B(udeco[123]), .C(n_58826), .Z(n_42900)
		);
	notech_ao3 i_125(.A(n_59618), .B(udeco[124]), .C(n_58826), .Z(n_42906)
		);
	notech_ao3 i_126(.A(n_59618), .B(udeco[125]), .C(n_58825), .Z(n_42912)
		);
	notech_ao3 i_127(.A(n_59619), .B(udeco[126]), .C(n_58825), .Z(n_42918)
		);
	notech_ao3 i_208(.A(n_59619), .B(udeco[103]), .C(n_58831), .Z(n_42780)
		);
	notech_nand2 i_2125672(.A(n_59693), .B(n_1610), .Z(n_3224));
	notech_nor2 i_292(.A(n_2225), .B(n_58683), .Z(n_44631));
	notech_nor2 i_293(.A(n_223393386), .B(n_58683), .Z(n_44637));
	notech_nor2 i_294(.A(n_224193378), .B(n_58685), .Z(n_44643));
	notech_nor2 i_295(.A(n_224993370), .B(n_58685), .Z(n_44649));
	notech_nor2 i_296(.A(n_225793362), .B(n_58685), .Z(n_44655));
	notech_nor2 i_297(.A(n_226593354), .B(n_58683), .Z(n_44661));
	notech_nor2 i_298(.A(n_227393346), .B(n_58683), .Z(n_44667));
	notech_nor2 i_299(.A(n_228191128), .B(n_58683), .Z(n_44673));
	notech_nor2 i_300(.A(n_228991136), .B(n_58683), .Z(n_44679));
	notech_nor2 i_301(.A(n_229791144), .B(n_58683), .Z(n_44685));
	notech_nor2 i_302(.A(n_230591152), .B(n_58685), .Z(n_44691));
	notech_nor2 i_303(.A(n_231391160), .B(n_58685), .Z(n_44697));
	notech_nor2 i_304(.A(n_232191168), .B(n_58685), .Z(n_44703));
	notech_nor2 i_305(.A(n_232991176), .B(n_58685), .Z(n_44709));
	notech_nor2 i_306(.A(n_233791184), .B(n_58685), .Z(n_44715));
	notech_nor2 i_312(.A(n_234891195), .B(n_58685), .Z(n_44751));
	notech_nor2 i_313(.A(n_235891205), .B(n_58685), .Z(n_44757));
	notech_nor2 i_314(.A(n_236891215), .B(n_58685), .Z(n_44763));
	notech_nor2 i_315(.A(n_237891225), .B(n_58685), .Z(n_44769));
	notech_nor2 i_316(.A(n_238991236), .B(n_58685), .Z(n_44775));
	notech_nor2 i_317(.A(n_239991246), .B(n_58691), .Z(n_44781));
	notech_nor2 i_318(.A(n_240991256), .B(n_58696), .Z(n_44787));
	notech_nor2 i_319(.A(n_241991266), .B(n_58696), .Z(n_44793));
	notech_nor2 i_320(.A(n_242991276), .B(n_58696), .Z(n_44799));
	notech_nor2 i_322(.A(n_243991286), .B(n_58696), .Z(n_44811));
	notech_nor2 i_323(.A(n_245091297), .B(n_58696), .Z(n_44817));
	notech_nor2 i_324(.A(n_3097), .B(n_39661), .Z(n_44823));
	notech_nor2 i_325(.A(n_3097), .B(n_39654), .Z(n_44829));
	notech_nor2 i_326(.A(n_3097), .B(n_39647), .Z(n_44835));
	notech_nor2 i_327(.A(n_3097), .B(n_39643), .Z(n_44841));
	notech_nor2 i_328(.A(n_3097), .B(n_39636), .Z(n_44847));
	notech_nor2 i_329(.A(n_3097), .B(n_39632), .Z(n_44853));
	notech_nor2 i_330(.A(n_3097), .B(n_39625), .Z(n_44859));
	notech_nor2 i_331(.A(n_3097), .B(n_39619), .Z(n_44865));
	notech_nor2 i_332(.A(n_3108), .B(n_39615), .Z(n_44871));
	notech_nor2 i_333(.A(n_3108), .B(n_39612), .Z(n_44877));
	notech_nor2 i_334(.A(n_3108), .B(n_39610), .Z(n_44883));
	notech_nor2 i_335(.A(n_3108), .B(n_39607), .Z(n_44889));
	notech_nor2 i_336(.A(n_3108), .B(n_39605), .Z(n_44895));
	notech_nor2 i_337(.A(n_3108), .B(n_39601), .Z(n_44901));
	notech_nor2 i_338(.A(n_3108), .B(n_39595), .Z(n_44907));
	notech_nor2 i_339(.A(n_3108), .B(n_39593), .Z(n_44913));
	notech_or2 i_515(.A(n_5761), .B(n_1996), .Z(n_1987));
	notech_nor2 i_163(.A(twobyte), .B(fpu), .Z(n_5761));
	notech_nand2 i_2225673(.A(n_59692), .B(n_1609), .Z(n_3223));
	notech_nand2 i_2325674(.A(n_59692), .B(n_1608), .Z(n_3222));
	notech_nor2 i_2462(.A(int_excl[5]), .B(n_260791454), .Z(n_1981));
	notech_nand2 i_2425675(.A(n_59692), .B(n_1607), .Z(n_3221));
	notech_or2 i_210235(.A(n_2058), .B(n_1981), .Z(n_5392));
	notech_or4 i_4329(.A(n_2219), .B(n_2958), .C(\to_acu2_0[3] ), .D(\to_acu2_0[2] 
		), .Z(n_5299));
	notech_nand2 i_2525676(.A(n_59692), .B(n_1606), .Z(n_3220));
	notech_nand2 i_65724(.A(n_2819), .B(n_2816), .Z(n_1973));
	notech_nand2 i_65731(.A(n_40185), .B(n_40183), .Z(n_1972));
	notech_nand3 i_5525706(.A(n_59692), .B(n_3246), .C(n_1605), .Z(n_3219)
		);
	notech_ao3 i_226(.A(udeco[103]), .B(rep), .C(n_58696), .Z(n_49769));
	notech_nand2 i_5825709(.A(n_59688), .B(n_1604), .Z(n_3218));
	notech_ao3 i_287(.A(n_59618), .B(repz), .C(n_58835), .Z(n_49763));
	notech_ao3 i_3434(.A(n_59618), .B(udeco[127]), .C(n_58835), .Z(n_42924)
		);
	notech_nor2 i_286(.A(n_58696), .B(n_39118), .Z(n_46109));
	notech_nand2 i_7325724(.A(n_59688), .B(n_1603), .Z(n_3217));
	notech_nand2 i_3730128(.A(n_1801), .B(n_38638), .Z(n_1821));
	notech_or4 i_3830129(.A(int_excl[1]), .B(int_excl[0]), .C(int_excl[2]), 
		.D(int_excl[3]), .Z(n_1820));
	notech_nor2 i_13(.A(n_2849), .B(pc_req), .Z(n_41571));
	notech_and2 i_32(.A(n_2084), .B(n_40184), .Z(n_1810));
	notech_nor2 i_156(.A(int_excl[1]), .B(int_excl[0]), .Z(n_1801));
	notech_nand2 i_190(.A(n_2081), .B(n_2080), .Z(n_1787));
	notech_nand3 i_224(.A(n_58835), .B(n_2833), .C(n_59618), .Z(n_1781));
	notech_xor2 i_6333(.A(i_ptr[3]), .B(n_2837), .Z(n_9538));
	notech_xor2 i_6334(.A(n_2836), .B(n_2839), .Z(n_9539));
	notech_xor2 i_6336(.A(imm_sz[0]), .B(i_ptr[0]), .Z(n_1741));
	notech_nand3 i_8325734(.A(n_16150155), .B(n_1601), .C(n_1529), .Z(n_3216
		));
	notech_nand3 i_8425735(.A(n_16150155), .B(n_1599), .C(n_1532), .Z(n_3215
		));
	notech_nand3 i_8525736(.A(n_59688), .B(n_1597), .C(n_1535), .Z(n_3214)
		);
	notech_nand3 i_8625737(.A(n_59688), .B(n_1595), .C(n_1538), .Z(n_3213)
		);
	notech_nand3 i_8825739(.A(n_59688), .B(n_1593), .C(n_1541), .Z(n_3212)
		);
	notech_nand2 i_9325744(.A(n_59688), .B(n_1592), .Z(n_3211));
	notech_nand2 i_9425745(.A(n_59688), .B(n_1591), .Z(n_3210));
	notech_nand2 i_9525746(.A(n_59688), .B(n_1590), .Z(n_3209));
	notech_nand2 i_9725748(.A(n_59692), .B(n_1589), .Z(n_3208));
	notech_nand2 i_9825749(.A(n_59688), .B(n_1588), .Z(n_3207));
	notech_nand3 i_10025751(.A(n_59692), .B(n_1418), .C(n_1587), .Z(n_3206)
		);
	notech_and4 i_11425765(.A(n_59692), .B(n_1418), .C(n_1585), .D(n_1556), 
		.Z(n_3205));
	notech_nand3 i_11525766(.A(n_16150155), .B(n_21191840), .C(n_1584), .Z(n_3204
		));
	notech_nand2 i_11625767(.A(n_59688), .B(n_1583), .Z(n_3203));
	notech_ao4 i_123146(.A(n_58696), .B(n_40104), .C(n_57481), .D(n_39822), 
		.Z(n_3202));
	notech_ao3 i_39275003(.A(n_59618), .B(opz[0]), .C(n_58831), .Z(n_3201)
		);
	notech_ao4 i_223147(.A(n_58696), .B(n_40105), .C(n_57481), .D(n_39823), 
		.Z(n_3200));
	notech_ao3 i_48475004(.A(n_59613), .B(opz[1]), .C(n_58831), .Z(n_3199)
		);
	notech_ao4 i_127801(.A(n_58696), .B(n_2225), .C(n_57481), .D(n_38509), .Z
		(n_3198));
	notech_ao4 i_427804(.A(n_58700), .B(n_224993370), .C(n_57479), .D(n_38513
		), .Z(n_3197));
	notech_ao4 i_627806(.A(n_58700), .B(n_226593354), .C(n_57475), .D(n_38515
		), .Z(n_3196));
	notech_ao4 i_727807(.A(n_58700), .B(n_227393346), .C(n_57475), .D(n_38518
		), .Z(n_3195));
	notech_ao4 i_827808(.A(n_58700), .B(n_228191128), .C(n_57475), .D(n_38520
		), .Z(n_3194));
	notech_ao4 i_927809(.A(n_58700), .B(n_228991136), .C(n_57475), .D(n_38522
		), .Z(n_3193));
	notech_ao4 i_1027810(.A(n_58696), .B(n_229791144), .C(n_57475), .D(n_38524
		), .Z(n_3192));
	notech_ao4 i_1127811(.A(n_58696), .B(n_230591152), .C(n_57473), .D(n_38526
		), .Z(n_3191));
	notech_ao4 i_1227812(.A(n_58696), .B(n_231391160), .C(n_57473), .D(n_38528
		), .Z(n_3190));
	notech_ao4 i_1327813(.A(n_58700), .B(n_232191168), .C(n_57473), .D(n_38530
		), .Z(n_3189));
	notech_ao4 i_1427814(.A(n_58696), .B(n_232991176), .C(n_57473), .D(n_38532
		), .Z(n_3188));
	notech_ao4 i_1527815(.A(n_58694), .B(n_233791184), .C(n_57473), .D(n_38534
		), .Z(n_3187));
	notech_ao4 i_1627816(.A(n_58691), .B(n_2163), .C(n_57475), .D(n_38536), 
		.Z(n_3186));
	notech_ao4 i_1727817(.A(n_58691), .B(n_2176), .C(n_57475), .D(n_38538), 
		.Z(n_3185));
	notech_ao4 i_1827818(.A(n_58694), .B(n_2186), .C(n_57475), .D(n_38540), 
		.Z(n_3184));
	notech_ao4 i_1927819(.A(n_58694), .B(n_2196), .C(n_57479), .D(n_38542), 
		.Z(n_3183));
	notech_ao4 i_2127821(.A(n_58694), .B(n_234891195), .C(n_57475), .D(n_38546
		), .Z(n_3182));
	notech_ao4 i_2227822(.A(n_58691), .B(n_235891205), .C(n_57475), .D(n_38548
		), .Z(n_3181));
	notech_ao4 i_2327823(.A(n_58691), .B(n_236891215), .C(n_57475), .D(n_38550
		), .Z(n_3180));
	notech_ao4 i_2427824(.A(n_58691), .B(n_237891225), .C(n_57475), .D(n_38552
		), .Z(n_3179));
	notech_ao4 i_2527825(.A(n_238991236), .B(n_58691), .C(n_57475), .D(n_38554
		), .Z(n_3178));
	notech_ao4 i_2627826(.A(n_239991246), .B(n_58691), .C(n_57475), .D(n_38556
		), .Z(n_3177));
	notech_ao4 i_2827828(.A(n_241991266), .B(n_58694), .C(n_57486), .D(n_38560
		), .Z(n_3176));
	notech_ao4 i_2927829(.A(n_242991276), .B(n_58694), .C(n_57486), .D(n_38562
		), .Z(n_3175));
	notech_ao4 i_3127831(.A(n_243991286), .B(n_58694), .C(n_57486), .D(n_38566
		), .Z(n_3174));
	notech_ao4 i_3227832(.A(n_245091297), .B(n_58694), .C(n_57486), .D(n_38568
		), .Z(n_3173));
	notech_ao4 i_3327833(.A(n_3097), .B(n_39661), .C(n_57486), .D(n_38570), 
		.Z(n_3172));
	notech_ao4 i_3427834(.A(n_3097), .B(n_39654), .C(n_57486), .D(n_38572), 
		.Z(n_3171));
	notech_ao4 i_3527835(.A(n_3097), .B(n_39647), .C(n_57486), .D(n_38574), 
		.Z(n_3170));
	notech_ao4 i_3627836(.A(n_3097), .B(n_39643), .C(n_57486), .D(n_38576), 
		.Z(n_3169));
	notech_ao4 i_3727837(.A(n_53727), .B(n_39636), .C(n_57486), .D(n_38578),
		 .Z(n_3168));
	notech_ao4 i_3827838(.A(n_53727), .B(n_39632), .C(n_57486), .D(n_38580),
		 .Z(n_3167));
	notech_ao4 i_3927839(.A(n_53727), .B(n_39625), .C(n_57490), .D(n_38583),
		 .Z(n_3166));
	notech_ao4 i_4027840(.A(n_53727), .B(n_39619), .C(n_57490), .D(n_38585),
		 .Z(n_3165));
	notech_ao4 i_4127841(.A(n_3108), .B(n_39615), .C(n_57490), .D(n_38588), 
		.Z(n_3164));
	notech_ao4 i_4227842(.A(n_3108), .B(n_39612), .C(n_57490), .D(n_38590), 
		.Z(n_3163));
	notech_ao4 i_4327843(.A(n_3108), .B(n_39610), .C(n_57490), .D(n_38592), 
		.Z(n_3162));
	notech_ao4 i_4427844(.A(n_3108), .B(n_39607), .C(n_57486), .D(n_38594), 
		.Z(n_3161));
	notech_ao4 i_4527845(.A(n_53788), .B(n_39605), .C(n_57486), .D(n_38596),
		 .Z(n_3160));
	notech_ao4 i_4627846(.A(n_53788), .B(n_39601), .C(n_57486), .D(n_38598),
		 .Z(n_3159));
	notech_ao4 i_4727847(.A(n_53788), .B(n_39595), .C(n_57490), .D(n_38600),
		 .Z(n_3158));
	notech_ao4 i_4827848(.A(n_53788), .B(n_39593), .C(n_57490), .D(n_38602),
		 .Z(n_3157));
	notech_ao4 i_7126189(.A(n_58694), .B(n_40204), .C(n_57486), .D(n_39228),
		 .Z(n_3156));
	notech_ao4 i_7226190(.A(n_58694), .B(n_40205), .C(n_57484), .D(n_39229),
		 .Z(n_3155));
	notech_ao4 i_7326191(.A(n_58694), .B(n_40185), .C(n_57481), .D(n_39231),
		 .Z(n_3154));
	notech_ao4 i_7426192(.A(n_58694), .B(n_40184), .C(n_57484), .D(n_39232),
		 .Z(n_3153));
	notech_ao4 i_7526193(.A(n_58694), .B(n_40211), .C(n_57484), .D(n_39234),
		 .Z(n_3152));
	notech_ao4 i_7626194(.A(n_58694), .B(n_40203), .C(n_57484), .D(n_39235),
		 .Z(n_3151));
	notech_ao4 i_7726195(.A(n_58672), .B(n_40183), .C(n_57481), .D(n_39237),
		 .Z(n_3150));
	notech_ao4 i_7826196(.A(n_58672), .B(n_40182), .C(n_57481), .D(n_39238),
		 .Z(n_3149));
	notech_ao4 i_7926197(.A(n_58672), .B(n_40181), .C(n_57481), .D(n_39240),
		 .Z(n_3148));
	notech_ao4 i_8026198(.A(n_58673), .B(n_40180), .C(n_57481), .D(n_39241),
		 .Z(n_3147));
	notech_nao3 i_6337(.A(n_2076), .B(n_40171), .C(twobyte), .Z(n_1740));
	notech_and3 i_20075005(.A(n_2120), .B(n_2076), .C(n_5761), .Z(n_17550169
		));
	notech_and2 i_22375006(.A(n_1574), .B(n_1474), .Z(n_3146));
	notech_and3 i_14375007(.A(n_59688), .B(n_2141), .C(n_18050174), .Z(n_5765
		));
	notech_and3 i_72700(.A(n_3146), .B(n_40193), .C(n_59613), .Z(n_3145));
	notech_ao3 i_74298(.A(n_18050174), .B(n_1568), .C(n_1475), .Z(n_3144));
	notech_ao3 i_75545(.A(n_58476), .B(n_1577), .C(n_2120), .Z(n_3143));
	notech_and3 i_70818(.A(n_16150155), .B(n_1572), .C(n_1565), .Z(n_3142)
		);
	notech_ao3 i_72382(.A(n_18050174), .B(n_1568), .C(n_1483), .Z(n_3141));
	notech_and4 i_70837(.A(n_59688), .B(n_2141), .C(n_18050174), .D(n_1484),
		 .Z(n_3140));
	notech_and2 i_72234(.A(n_59688), .B(n_2129), .Z(n_3139));
	notech_ao3 i_70765(.A(n_1489), .B(n_5765), .C(n_2123), .Z(n_3138));
	notech_and4 i_70743(.A(n_59693), .B(n_18050174), .C(n_2141), .D(n_1485),
		 .Z(n_3137));
	notech_and4 i_71564(.A(n_18050174), .B(n_1568), .C(n_1489), .D(n_2128), 
		.Z(n_3136));
	notech_nand2 i_1359(.A(n_2867), .B(n_1476), .Z(n_3134));
	notech_ao4 i_1336(.A(n_39117), .B(n_261691463), .C(n_261591462), .D(n_5304
		), .Z(n_3130));
	notech_nand3 i_1332(.A(n_38431), .B(n_38428), .C(n_38434), .Z(n_3128));
	notech_nand3 i_3965(.A(db67), .B(n_41571), .C(n_250691353), .Z(n_3120)
		);
	notech_ao3 i_1133(.A(\fpu_modrm[2] ), .B(\fpu_indrm[0] ), .C(\fpu_modrm[1] 
		), .Z(n_3119));
	notech_ao4 i_1129(.A(n_250391350), .B(in128[55]), .C(n_3095), .D(in128[
		63]), .Z(n_3116));
	notech_ao4 i_1125(.A(n_250091347), .B(in128[54]), .C(n_3095), .D(in128[
		62]), .Z(n_3115));
	notech_ao4 i_1121(.A(n_249791344), .B(in128[53]), .C(n_3095), .D(in128[
		61]), .Z(n_3114));
	notech_ao4 i_1117(.A(n_249491341), .B(in128[52]), .C(n_3095), .D(in128[
		60]), .Z(n_3113));
	notech_ao4 i_1113(.A(n_249191338), .B(in128[51]), .C(n_3095), .D(in128[
		59]), .Z(n_3112));
	notech_ao4 i_1109(.A(n_248891335), .B(in128[50]), .C(n_3095), .D(in128[
		58]), .Z(n_3111));
	notech_ao4 i_1105(.A(n_248591332), .B(in128[49]), .C(n_3095), .D(in128[
		57]), .Z(n_3110));
	notech_ao4 i_1101(.A(n_248291329), .B(in128[48]), .C(n_3095), .D(in128[
		56]), .Z(n_3109));
	notech_nao3 i_7(.A(n_59618), .B(n_248191328), .C(n_58835), .Z(n_3108));
	notech_and4 i_183(.A(imm_sz[2]), .B(n_2914), .C(n_245391300), .D(n_2915)
		, .Z(n_3107));
	notech_ao4 i_1095(.A(n_247891325), .B(in128[55]), .C(n_247791324), .D(in128
		[47]), .Z(n_3105));
	notech_ao4 i_1091(.A(n_247491321), .B(in128[54]), .C(n_247791324), .D(in128
		[46]), .Z(n_3104));
	notech_ao4 i_1087(.A(n_247191318), .B(in128[53]), .C(n_247791324), .D(in128
		[45]), .Z(n_3103));
	notech_ao4 i_1083(.A(n_246891315), .B(in128[52]), .C(n_247791324), .D(in128
		[44]), .Z(n_3102));
	notech_ao4 i_1079(.A(n_246591312), .B(in128[51]), .C(n_247791324), .D(in128
		[43]), .Z(n_3101));
	notech_ao4 i_1075(.A(n_246291309), .B(in128[50]), .C(n_247791324), .D(in128
		[42]), .Z(n_3100));
	notech_ao4 i_1071(.A(n_245991306), .B(in128[49]), .C(n_247791324), .D(in128
		[41]), .Z(n_3099));
	notech_ao4 i_1067(.A(n_245691303), .B(in128[48]), .C(n_247791324), .D(in128
		[40]), .Z(n_3098));
	notech_nao3 i_2(.A(n_59613), .B(n_245591302), .C(n_58835), .Z(n_3097));
	notech_ao3 i_154(.A(n_2890), .B(n_2900), .C(n_2897), .Z(n_3095));
	notech_ao4 i_1055(.A(n_3060), .B(n_40022), .C(n_2921), .D(n_40030), .Z(n_3091
		));
	notech_ao4 i_1054(.A(n_2923), .B(n_40054), .C(n_2922), .D(n_40038), .Z(n_3090
		));
	notech_ao4 i_1043(.A(n_3060), .B(n_40021), .C(n_2921), .D(n_40029), .Z(n_3086
		));
	notech_ao4 i_1042(.A(n_2923), .B(n_40053), .C(n_2922), .D(n_40037), .Z(n_3085
		));
	notech_ao4 i_1031(.A(n_3060), .B(n_40019), .C(n_2921), .D(n_40027), .Z(n_3081
		));
	notech_ao4 i_1030(.A(n_2923), .B(n_40051), .C(n_2922), .D(n_40035), .Z(n_3080
		));
	notech_ao4 i_1019(.A(n_3060), .B(n_40018), .C(n_2921), .D(n_40026), .Z(n_3076
		));
	notech_ao4 i_1018(.A(n_2923), .B(n_40050), .C(n_2922), .D(n_40034), .Z(n_3075
		));
	notech_ao4 i_1007(.A(n_3060), .B(n_40017), .C(n_2921), .D(n_40025), .Z(n_3071
		));
	notech_ao4 i_1006(.A(n_2923), .B(n_40049), .C(n_2922), .D(n_40033), .Z(n_3070
		));
	notech_ao4 i_995(.A(n_3060), .B(n_40016), .C(n_2921), .D(n_40024), .Z(n_3066
		));
	notech_ao4 i_994(.A(n_2923), .B(n_40048), .C(n_2922), .D(n_40032), .Z(n_3065
		));
	notech_ao4 i_983(.A(n_3060), .B(n_40015), .C(n_2921), .D(n_40023), .Z(n_3061
		));
	notech_or2 i_184(.A(n_2924), .B(n_238191228), .Z(n_3060));
	notech_ao4 i_982(.A(n_2923), .B(n_40047), .C(n_2922), .D(n_40031), .Z(n_3057
		));
	notech_and2 i_969(.A(n_237491221), .B(n_3052), .Z(n_3053));
	notech_ao4 i_968(.A(n_2924), .B(n_40014), .C(n_2923), .D(n_40046), .Z(n_3052
		));
	notech_and2 i_951(.A(n_236491211), .B(n_3047), .Z(n_3048));
	notech_ao4 i_950(.A(n_2924), .B(n_40013), .C(n_2923), .D(n_40045), .Z(n_3047
		));
	notech_and2 i_939(.A(n_235491201), .B(n_3042), .Z(n_3043));
	notech_ao4 i_938(.A(n_2924), .B(n_40012), .C(n_2923), .D(n_40044), .Z(n_3042
		));
	notech_and2 i_927(.A(n_234491191), .B(n_3037), .Z(n_3038));
	notech_ao4 i_926(.A(n_2924), .B(n_40011), .C(n_2923), .D(n_40043), .Z(n_3037
		));
	notech_ao4 i_919(.A(n_40037), .B(n_2918), .C(n_40005), .D(n_2916), .Z(n_3035
		));
	notech_and2 i_917(.A(n_3032), .B(n_233691183), .Z(n_3033));
	notech_ao4 i_916(.A(n_40029), .B(n_2907), .C(n_2905), .D(n_40045), .Z(n_3032
		));
	notech_ao4 i_909(.A(n_2918), .B(n_40036), .C(n_2916), .D(n_40004), .Z(n_3030
		));
	notech_and2 i_907(.A(n_3027), .B(n_232891175), .Z(n_3028));
	notech_ao4 i_906(.A(n_2907), .B(n_40028), .C(n_2905), .D(n_40044), .Z(n_3027
		));
	notech_ao4 i_899(.A(n_2918), .B(n_40035), .C(n_2916), .D(n_40003), .Z(n_3025
		));
	notech_and2 i_897(.A(n_3022), .B(n_232091167), .Z(n_3023));
	notech_ao4 i_896(.A(n_2907), .B(n_40027), .C(n_2905), .D(n_40043), .Z(n_3022
		));
	notech_ao4 i_889(.A(n_2918), .B(n_40034), .C(n_2916), .D(n_40002), .Z(n_3020
		));
	notech_and2 i_887(.A(n_3017), .B(n_231291159), .Z(n_3018));
	notech_ao4 i_886(.A(n_2907), .B(n_40026), .C(n_2905), .D(n_40042), .Z(n_3017
		));
	notech_ao4 i_879(.A(n_2918), .B(n_40033), .C(n_2916), .D(n_40001), .Z(n_3015
		));
	notech_and2 i_877(.A(n_3012), .B(n_230491151), .Z(n_3013));
	notech_ao4 i_876(.A(n_2907), .B(n_40025), .C(n_2905), .D(n_40041), .Z(n_3012
		));
	notech_ao4 i_869(.A(n_2918), .B(n_40032), .C(n_2916), .D(n_40000), .Z(n_3010
		));
	notech_and2 i_867(.A(n_3007), .B(n_229691143), .Z(n_3008));
	notech_ao4 i_866(.A(n_2907), .B(n_40024), .C(n_2905), .D(n_40040), .Z(n_3007
		));
	notech_ao4 i_859(.A(n_2918), .B(n_40031), .C(n_2916), .D(n_39999), .Z(n_3005
		));
	notech_and2 i_857(.A(n_3002), .B(n_228891135), .Z(n_3003));
	notech_ao4 i_856(.A(n_2907), .B(n_40023), .C(n_2905), .D(n_40039), .Z(n_3002
		));
	notech_ao4 i_849(.A(n_2906), .B(n_40022), .C(n_2898), .D(n_40172), .Z(n_3000
		));
	notech_and2 i_847(.A(n_2997), .B(n_228091127), .Z(n_2998));
	notech_ao4 i_846(.A(n_2904), .B(n_40038), .C(n_39834), .D(n_40030), .Z(n_2997
		));
	notech_ao4 i_839(.A(n_2906), .B(n_40021), .C(n_2898), .D(n_40173), .Z(n_2995
		));
	notech_and2 i_837(.A(n_2992), .B(n_227293347), .Z(n_2993));
	notech_ao4 i_836(.A(n_2904), .B(n_40037), .C(n_40029), .D(n_39834), .Z(n_2992
		));
	notech_ao4 i_829(.A(n_2906), .B(n_40020), .C(n_2898), .D(n_40206), .Z(n_2990
		));
	notech_and2 i_827(.A(n_2987), .B(n_226493355), .Z(n_2988));
	notech_ao4 i_826(.A(n_2904), .B(n_40036), .C(n_39834), .D(n_40028), .Z(n_2987
		));
	notech_ao4 i_819(.A(n_2906), .B(n_40019), .C(n_2898), .D(n_40207), .Z(n_2985
		));
	notech_and2 i_817(.A(n_2982), .B(n_225693363), .Z(n_2983));
	notech_ao4 i_816(.A(n_2904), .B(n_40035), .C(n_39834), .D(n_40027), .Z(n_2982
		));
	notech_ao4 i_809(.A(n_2906), .B(n_40018), .C(n_2898), .D(n_40208), .Z(n_2980
		));
	notech_and2 i_807(.A(n_2977), .B(n_224893371), .Z(n_2978));
	notech_ao4 i_806(.A(n_2904), .B(n_40034), .C(n_39834), .D(n_40026), .Z(n_2977
		));
	notech_ao4 i_799(.A(n_2906), .B(n_40017), .C(n_2898), .D(n_40197), .Z(n_2975
		));
	notech_and2 i_797(.A(n_2972), .B(n_224093379), .Z(n_2973));
	notech_ao4 i_796(.A(n_2904), .B(n_40033), .C(n_39834), .D(n_40025), .Z(n_2972
		));
	notech_ao4 i_789(.A(n_2906), .B(n_40016), .C(n_2898), .D(n_40196), .Z(n_2970
		));
	notech_and2 i_787(.A(n_2967), .B(n_223293387), .Z(n_2968));
	notech_ao4 i_786(.A(n_2904), .B(n_40032), .C(n_39834), .D(n_40024), .Z(n_2967
		));
	notech_ao4 i_779(.A(n_2906), .B(n_40015), .C(n_40174), .D(n_2898), .Z(n_2965
		));
	notech_and2 i_777(.A(n_2962), .B(n_2224), .Z(n_2963));
	notech_ao4 i_776(.A(n_2904), .B(n_40031), .C(n_40023), .D(n_39834), .Z(n_2962
		));
	notech_ao4 i_19273382(.A(db67), .B(n_39117), .C(n_1991), .D(n_38434), .Z
		(n_2961));
	notech_nao3 i_540(.A(\to_acu2_0[0] ), .B(\to_acu2_0[1] ), .C(n_251191358
		), .Z(n_2958));
	notech_nand3 i_65819(.A(n_2212), .B(n_2955), .C(n_2078), .Z(n_2957));
	notech_and4 i_696(.A(n_40164), .B(n_40163), .C(n_40162), .D(n_40161), .Z
		(n_2955));
	notech_and4 i_690(.A(n_40164), .B(n_40155), .C(n_40187), .D(n_40154), .Z
		(n_2950));
	notech_and2 i_633(.A(n_2202), .B(n_2943), .Z(n_2944));
	notech_ao4 i_632(.A(n_2924), .B(n_40010), .C(n_2923), .D(n_40042), .Z(n_2943
		));
	notech_and2 i_621(.A(n_2192), .B(n_2938), .Z(n_2939));
	notech_ao4 i_620(.A(n_2924), .B(n_40009), .C(n_2923), .D(n_40041), .Z(n_2938
		));
	notech_and2 i_609(.A(n_2182), .B(n_2933), .Z(n_2934));
	notech_ao4 i_608(.A(n_2924), .B(n_40008), .C(n_2923), .D(n_40040), .Z(n_2933
		));
	notech_or4 i_148(.A(imm_sz[0]), .B(imm_sz[1]), .C(n_2890), .D(n_2897), .Z
		(n_2929));
	notech_nand2 i_147(.A(n_2884), .B(n_39838), .Z(n_2928));
	notech_and2 i_596(.A(n_2171), .B(n_2925), .Z(n_2926));
	notech_ao4 i_595(.A(n_2924), .B(n_40007), .C(n_2923), .D(n_40039), .Z(n_2925
		));
	notech_nand2 i_187(.A(n_2914), .B(n_2167), .Z(n_2924));
	notech_nand2 i_151(.A(n_2884), .B(n_2917), .Z(n_2923));
	notech_nao3 i_149(.A(n_2887), .B(n_2884), .C(n_39845), .Z(n_2922));
	notech_or4 i_155(.A(imm_sz[0]), .B(imm_sz[1]), .C(n_2887), .D(n_39845), 
		.Z(n_2921));
	notech_ao4 i_587(.A(n_2918), .B(n_40038), .C(n_2916), .D(n_40006), .Z(n_2919
		));
	notech_or2 i_180(.A(n_2885), .B(n_39834), .Z(n_2918));
	notech_and4 i_131(.A(n_2891), .B(n_2887), .C(n_39841), .D(n_39835), .Z(n_2917
		));
	notech_nand2 i_178(.A(n_2914), .B(n_2162), .Z(n_2916));
	notech_and2 i_142(.A(n_2885), .B(n_2161), .Z(n_2915));
	notech_and4 i_18(.A(n_39841), .B(n_2891), .C(n_2887), .D(n_2890), .Z(n_2914
		));
	notech_and2 i_581(.A(n_2908), .B(n_2160), .Z(n_2909));
	notech_ao4 i_580(.A(n_2907), .B(n_40030), .C(n_2905), .D(n_40046), .Z(n_2908
		));
	notech_or2 i_186(.A(n_2885), .B(n_2906), .Z(n_2907));
	notech_or2 i_104(.A(n_2897), .B(n_2890), .Z(n_2906));
	notech_or2 i_181(.A(n_2885), .B(n_2904), .Z(n_2905));
	notech_or4 i_132(.A(n_2887), .B(n_2891), .C(n_2890), .D(n_2155), .Z(n_2904
		));
	notech_ao3 i_830084(.A(imm_sz[1]), .B(imm_sz[2]), .C(imm_sz[0]), .Z(n_2900
		));
	notech_or2 i_21(.A(n_2897), .B(n_39835), .Z(n_2898));
	notech_nao3 i_574(.A(n_2891), .B(n_39841), .C(n_2887), .Z(n_2897));
	notech_and2 i_130(.A(n_2887), .B(n_2893), .Z(n_2894));
	notech_ao3 i_19(.A(n_39841), .B(n_2890), .C(n_2891), .Z(n_2893));
	notech_xor2 i_2230078(.A(displc[1]), .B(n_2888), .Z(n_2891));
	notech_xor2 i_2330079(.A(displc[2]), .B(n_2889), .Z(n_2890));
	notech_nand2 i_352(.A(displc[1]), .B(n_39846), .Z(n_2889));
	notech_ao4 i_2831(.A(n_2146), .B(n_40177), .C(n_40178), .D(n_39861), .Z(n_2888
		));
	notech_or2 i_2130077(.A(n_2154), .B(n_2153), .Z(n_2887));
	notech_xor2 i_217(.A(n_40177), .B(sib_dec), .Z(n_2886));
	notech_nor2 i_4(.A(n_2884), .B(n_2143), .Z(n_2885));
	notech_nor2 i_630081(.A(imm_sz[0]), .B(imm_sz[1]), .Z(n_2884));
	notech_nao3 i_546(.A(ie), .B(n_40193), .C(ipg_fault), .Z(n_2882));
	notech_and2 i_541(.A(n_38628), .B(n_38627), .Z(n_2878));
	notech_and4 i_543(.A(n_38631), .B(n_38630), .C(n_38634), .D(n_38633), .Z
		(n_2877));
	notech_ao3 i_20173381(.A(n_59613), .B(in128[1]), .C(n_58835), .Z(n_47603
		));
	notech_nand2 i_532(.A(n_60686), .B(term_f), .Z(n_2874));
	notech_nao3 i_530(.A(n_38656), .B(n_39847), .C(idx_deco[1]), .Z(n_2873)
		);
	notech_nao3 i_27074739(.A(cpl[0]), .B(cpl[1]), .C(n_2056), .Z(n_21191840
		));
	notech_nao3 i_28774722(.A(cpl[0]), .B(cpl[1]), .C(n_3246), .Z(n_21291841
		));
	notech_or2 i_29674713(.A(n_3246), .B(n_161751607), .Z(n_21391842));
	notech_and2 i_35774652(.A(n_17550169), .B(\to_acu2_0[71] ), .Z(n_21791846
		));
	notech_or4 i_35874651(.A(n_58476), .B(idx_deco[1]), .C(n_2138), .D(idx_deco
		[0]), .Z(n_21891847));
	notech_or4 i_35974650(.A(idx_deco[1]), .B(n_58476), .C(n_38656), .D(n_2138
		), .Z(n_21991848));
	notech_nao3 i_36074649(.A(idx_deco[1]), .B(n_38656), .C(n_18050174), .Z(n_22091849
		));
	notech_and2 i_122673785(.A(n_17550169), .B(\to_acu2_0[70] ), .Z(n_108192702
		));
	notech_and2 i_123473777(.A(n_17550169), .B(\to_acu2_0[75] ), .Z(n_108292703
		));
	notech_and2 i_289092617(.A(lenpc1[8]), .B(n_38330), .Z(n_108392704));
	notech_and2 i_289192618(.A(lenpc1[9]), .B(n_38330), .Z(n_108492705));
	notech_and2 i_289292619(.A(lenpc1[10]), .B(n_38330), .Z(n_108592706));
	notech_and2 i_289392620(.A(lenpc1[11]), .B(n_38330), .Z(n_108692707));
	notech_and2 i_289492621(.A(lenpc1[12]), .B(n_38330), .Z(n_108792708));
	notech_and2 i_289592622(.A(lenpc1[13]), .B(n_38330), .Z(n_108892709));
	notech_and2 i_289692623(.A(lenpc1[14]), .B(n_38330), .Z(n_108992710));
	notech_and2 i_289792624(.A(lenpc1[15]), .B(n_38330), .Z(n_109092711));
	notech_and2 i_289892625(.A(lenpc1[16]), .B(n_38330), .Z(n_109192712));
	notech_and2 i_289992626(.A(lenpc1[17]), .B(n_38330), .Z(n_109292713));
	notech_and2 i_290092627(.A(lenpc1[18]), .B(n_38330), .Z(n_109392714));
	notech_and2 i_290192628(.A(lenpc1[19]), .B(n_38330), .Z(n_109492715));
	notech_and2 i_290292629(.A(lenpc1[20]), .B(n_38330), .Z(n_109592716));
	notech_and2 i_290392630(.A(lenpc1[21]), .B(n_58407), .Z(n_109692717));
	notech_and2 i_290492631(.A(lenpc1[22]), .B(n_58407), .Z(n_109792718));
	notech_and2 i_290592632(.A(lenpc1[23]), .B(n_58407), .Z(n_109892719));
	notech_and2 i_290692633(.A(lenpc1[24]), .B(n_58407), .Z(n_109992720));
	notech_and2 i_290792634(.A(lenpc1[25]), .B(n_58407), .Z(n_110092721));
	notech_and2 i_290892635(.A(lenpc1[26]), .B(n_58407), .Z(n_110192722));
	notech_and2 i_290992636(.A(lenpc1[27]), .B(n_58407), .Z(n_110292723));
	notech_and2 i_291092637(.A(lenpc1[28]), .B(n_58407), .Z(n_110392724));
	notech_and2 i_291192638(.A(lenpc1[29]), .B(n_58407), .Z(n_110492725));
	notech_and2 i_291292639(.A(lenpc1[30]), .B(n_38330), .Z(n_110592726));
	notech_and2 i_291392640(.A(lenpc1[31]), .B(n_58407), .Z(n_110692727));
	notech_and3 i_293092641(.A(n_2124), .B(lenpc2[21]), .C(n_59613), .Z(n_110792728
		));
	notech_and3 i_293192642(.A(n_2124), .B(lenpc2[22]), .C(n_59618), .Z(n_110892729
		));
	notech_and3 i_293292643(.A(n_2124), .B(lenpc2[23]), .C(n_59618), .Z(n_110992730
		));
	notech_and3 i_293392644(.A(n_2124), .B(lenpc2[24]), .C(n_59618), .Z(n_111092731
		));
	notech_and3 i_293492645(.A(n_2124), .B(lenpc2[25]), .C(n_59618), .Z(n_111192732
		));
	notech_and3 i_293592646(.A(n_2124), .B(lenpc2[26]), .C(n_59618), .Z(n_111292733
		));
	notech_nao3 i_18274818(.A(n_2847), .B(inst_deco1[80]), .C(n_1995), .Z(n_123192852
		));
	notech_ao3 i_18574815(.A(n_2847), .B(inst_deco1[81]), .C(n_1995), .Z(n_123492855
		));
	notech_nao3 i_20374800(.A(n_2847), .B(inst_deco1[86]), .C(n_1995), .Z(n_123792858
		));
	notech_nao3 i_25174758(.A(n_2847), .B(inst_deco1[106]), .C(n_1995), .Z(n_126492885
		));
	notech_and3 i_309592647(.A(n_2124), .B(to_acu2[39]), .C(n_59618), .Z(n_130392924
		));
	notech_and3 i_288592648(.A(n_39847), .B(n_1473), .C(n_1741), .Z(useq_ptr
		[0]));
	notech_and3 i_288392649(.A(n_39847), .B(n_1473), .C(n_9539), .Z(useq_ptr
		[2]));
	notech_ao3 i_288292650(.A(n_1473), .B(n_39847), .C(n_9538), .Z(useq_ptr[
		3]));
	notech_ao4 i_142673585(.A(n_58400), .B(n_39116), .C(n_58476), .D(n_39989
		), .Z(n_130892929));
	notech_ao4 i_142573586(.A(n_58400), .B(n_39114), .C(n_58476), .D(n_39988
		), .Z(n_131092931));
	notech_ao4 i_142473587(.A(n_58400), .B(n_39112), .C(n_58476), .D(n_39987
		), .Z(n_131192932));
	notech_ao4 i_142373588(.A(n_58400), .B(n_39110), .C(n_58476), .D(n_39986
		), .Z(n_131292933));
	notech_ao4 i_142273589(.A(n_58400), .B(n_39108), .C(n_58476), .D(n_39985
		), .Z(n_131392934));
	notech_ao4 i_142173590(.A(n_58400), .B(n_39106), .C(n_58477), .D(n_39984
		), .Z(n_131592936));
	notech_ao4 i_142073591(.A(n_58400), .B(n_39104), .C(n_58476), .D(n_39983
		), .Z(n_131692937));
	notech_ao4 i_141973592(.A(n_58400), .B(n_39102), .C(n_58477), .D(n_39982
		), .Z(n_131792938));
	notech_ao4 i_141873593(.A(n_58401), .B(n_39100), .C(n_58477), .D(n_39981
		), .Z(n_131892939));
	notech_ao4 i_141773594(.A(n_58401), .B(n_39098), .C(n_58476), .D(n_39980
		), .Z(n_131992940));
	notech_ao4 i_141673595(.A(n_58400), .B(n_39096), .C(n_58476), .D(n_39979
		), .Z(n_132092941));
	notech_ao4 i_141573596(.A(n_58400), .B(n_39094), .C(n_58476), .D(n_39978
		), .Z(n_132192942));
	notech_ao4 i_141073601(.A(n_58400), .B(n_39087), .C(n_58476), .D(n_39974
		), .Z(n_132392944));
	notech_ao4 i_140873603(.A(n_58400), .B(n_39085), .C(n_58472), .D(n_39973
		), .Z(n_132592946));
	notech_ao4 i_140773604(.A(n_58400), .B(n_39083), .C(n_58472), .D(n_39972
		), .Z(n_132692947));
	notech_ao4 i_140673605(.A(n_58396), .B(n_39081), .C(n_58472), .D(n_39971
		), .Z(n_132792948));
	notech_ao4 i_140573606(.A(n_58396), .B(n_39079), .C(n_58472), .D(n_39970
		), .Z(n_132892949));
	notech_ao4 i_140473607(.A(n_58396), .B(n_39077), .C(n_58472), .D(n_39969
		), .Z(n_132992950));
	notech_ao4 i_140373608(.A(n_58472), .B(n_39968), .C(n_161751607), .D(n_40193
		), .Z(n_133092951));
	notech_ao4 i_140173610(.A(n_58396), .B(n_39074), .C(n_58472), .D(n_39967
		), .Z(n_133292953));
	notech_ao4 i_140073611(.A(n_58396), .B(n_39072), .C(n_58472), .D(n_39966
		), .Z(n_133392954));
	notech_ao4 i_139973612(.A(n_58396), .B(n_39070), .C(n_58476), .D(n_39965
		), .Z(n_133492955));
	notech_ao4 i_139873613(.A(n_58396), .B(n_39067), .C(n_58476), .D(n_39964
		), .Z(n_133592956));
	notech_ao4 i_139773614(.A(n_58400), .B(n_39065), .C(n_58476), .D(n_39963
		), .Z(n_133692957));
	notech_ao4 i_139673615(.A(n_58400), .B(n_39063), .C(n_58476), .D(n_39962
		), .Z(n_133792958));
	notech_ao4 i_139473617(.A(n_58400), .B(n_39059), .C(n_58472), .D(n_39960
		), .Z(n_133892959));
	notech_ao4 i_139173620(.A(n_58396), .B(n_39053), .C(n_58472), .D(n_39957
		), .Z(n_133992960));
	notech_ao4 i_138773624(.A(n_58396), .B(n_39045), .C(n_58476), .D(n_39953
		), .Z(n_134092961));
	notech_ao4 i_138673625(.A(n_58396), .B(n_39043), .C(n_58472), .D(n_39952
		), .Z(n_134192962));
	notech_ao4 i_138573626(.A(n_58396), .B(n_39041), .C(n_58477), .D(n_39951
		), .Z(n_134292963));
	notech_ao4 i_138473627(.A(n_58401), .B(n_39039), .C(n_58479), .D(n_39950
		), .Z(n_134392964));
	notech_ao4 i_138173630(.A(n_58479), .B(n_39948), .C(n_2056), .D(n_38633)
		, .Z(n_134492965));
	notech_ao4 i_137173640(.A(n_58479), .B(n_39943), .C(n_2056), .D(n_38625)
		, .Z(n_134692967));
	notech_ao4 i_136973642(.A(n_58479), .B(n_39942), .C(n_2056), .D(n_38624)
		, .Z(n_134892969));
	notech_ao4 i_136773644(.A(n_58403), .B(n_39029), .C(n_58479), .D(n_39941
		), .Z(n_135092971));
	notech_ao4 i_136673645(.A(n_58403), .B(n_39027), .C(n_58479), .D(n_39940
		), .Z(n_135192972));
	notech_ao4 i_136573646(.A(n_58403), .B(n_39025), .C(n_58479), .D(n_39939
		), .Z(n_135292973));
	notech_ao4 i_136473647(.A(n_58403), .B(n_39023), .C(n_58479), .D(n_39938
		), .Z(n_135392974));
	notech_ao4 i_136373648(.A(n_58403), .B(n_39021), .C(n_58479), .D(n_39937
		), .Z(n_135492975));
	notech_ao4 i_136273649(.A(n_58403), .B(n_39019), .C(n_58479), .D(n_39936
		), .Z(n_135592976));
	notech_ao4 i_136173650(.A(n_58403), .B(n_39017), .C(n_58479), .D(n_39935
		), .Z(n_135692977));
	notech_ao4 i_135973652(.A(n_58403), .B(n_39013), .C(n_58479), .D(n_39933
		), .Z(n_135792978));
	notech_ao4 i_135873653(.A(n_58403), .B(n_39011), .C(n_58479), .D(n_39932
		), .Z(n_135892979));
	notech_ao4 i_135773654(.A(n_58403), .B(n_39009), .C(n_58479), .D(n_39931
		), .Z(n_135992980));
	notech_ao4 i_135673655(.A(n_58403), .B(n_39007), .C(n_58479), .D(n_39930
		), .Z(n_136092981));
	notech_ao4 i_135573656(.A(n_58403), .B(n_39005), .C(n_58479), .D(n_39929
		), .Z(n_136192982));
	notech_ao4 i_135473657(.A(n_58403), .B(n_39003), .C(n_58477), .D(n_39928
		), .Z(n_136292983));
	notech_ao4 i_135373658(.A(n_58403), .B(n_39001), .C(n_58477), .D(n_39927
		), .Z(n_136392984));
	notech_ao4 i_135273659(.A(n_58403), .B(n_38999), .C(n_58477), .D(n_39926
		), .Z(n_136492985));
	notech_ao4 i_135173660(.A(n_58401), .B(n_38997), .C(n_58477), .D(n_39925
		), .Z(n_136592986));
	notech_ao4 i_135073661(.A(n_58401), .B(n_38995), .C(n_58477), .D(n_39924
		), .Z(n_136692987));
	notech_ao4 i_134973662(.A(n_58401), .B(n_38993), .C(n_58477), .D(n_39923
		), .Z(n_136792988));
	notech_ao4 i_134873663(.A(n_58401), .B(n_38991), .C(n_58477), .D(n_39922
		), .Z(n_136892989));
	notech_ao4 i_134773664(.A(n_58401), .B(n_38989), .C(n_58477), .D(n_39921
		), .Z(n_136992990));
	notech_ao4 i_134673665(.A(n_58401), .B(n_38987), .C(n_58477), .D(n_39920
		), .Z(n_137092991));
	notech_ao4 i_134473667(.A(n_58401), .B(n_38983), .C(n_58477), .D(n_39918
		), .Z(n_137192992));
	notech_ao4 i_134373668(.A(n_58401), .B(n_38981), .C(n_58479), .D(n_39917
		), .Z(n_137292993));
	notech_ao4 i_134173670(.A(n_58401), .B(n_38977), .C(n_58479), .D(n_39915
		), .Z(n_137392994));
	notech_ao4 i_134073671(.A(n_58403), .B(n_38975), .C(n_58477), .D(n_39914
		), .Z(n_137492995));
	notech_ao4 i_133973672(.A(n_58401), .B(n_38973), .C(n_58477), .D(n_39913
		), .Z(n_137592996));
	notech_ao4 i_133873673(.A(n_58401), .B(n_38971), .C(n_58477), .D(n_39912
		), .Z(n_137692997));
	notech_ao4 i_133773674(.A(n_58401), .B(n_38969), .C(n_58477), .D(n_39911
		), .Z(n_137792998));
	notech_ao4 i_133673675(.A(n_58401), .B(n_38967), .C(n_58472), .D(n_39910
		), .Z(n_137892999));
	notech_ao4 i_133573676(.A(n_58389), .B(n_38965), .C(n_58465), .D(n_39909
		), .Z(n_137993000));
	notech_ao4 i_133473677(.A(n_58389), .B(n_38963), .C(n_58465), .D(n_39908
		), .Z(n_138093001));
	notech_ao4 i_133373678(.A(n_58389), .B(n_38961), .C(n_58465), .D(n_39907
		), .Z(n_138193002));
	notech_ao4 i_133273679(.A(n_58389), .B(n_38959), .C(n_58465), .D(n_39906
		), .Z(n_138293003));
	notech_ao4 i_133173680(.A(n_58389), .B(n_38957), .C(n_58465), .D(n_39905
		), .Z(n_138393004));
	notech_ao4 i_133073681(.A(n_58389), .B(n_38955), .C(n_58465), .D(n_39904
		), .Z(n_138493005));
	notech_ao4 i_132973682(.A(n_58389), .B(n_38953), .C(n_58465), .D(n_39903
		), .Z(n_138593006));
	notech_ao4 i_132873683(.A(n_58391), .B(n_38951), .C(n_58465), .D(n_39902
		), .Z(n_138693007));
	notech_ao4 i_132773684(.A(n_58391), .B(n_38949), .C(n_58467), .D(n_39901
		), .Z(n_138793008));
	notech_ao4 i_132673685(.A(n_58391), .B(n_38947), .C(n_58467), .D(n_39900
		), .Z(n_138893009));
	notech_ao4 i_132573686(.A(n_58391), .B(n_38945), .C(n_58467), .D(n_39899
		), .Z(n_138993010));
	notech_ao4 i_132473687(.A(n_58391), .B(n_38943), .C(n_58467), .D(n_39898
		), .Z(n_139093011));
	notech_ao4 i_132373688(.A(n_58391), .B(n_38941), .C(n_58467), .D(n_39897
		), .Z(n_139193012));
	notech_ao4 i_132273689(.A(n_58391), .B(n_38939), .C(n_58467), .D(n_39896
		), .Z(n_139293013));
	notech_ao4 i_132173690(.A(n_58389), .B(n_38937), .C(n_58467), .D(n_39895
		), .Z(n_139393014));
	notech_ao4 i_132073691(.A(n_58388), .B(n_38935), .C(n_58467), .D(n_39894
		), .Z(n_139493015));
	notech_ao4 i_131973692(.A(n_58388), .B(n_38933), .C(n_58464), .D(n_39893
		), .Z(n_139593016));
	notech_ao4 i_131873693(.A(n_58388), .B(n_38931), .C(n_58464), .D(n_39892
		), .Z(n_139693017));
	notech_ao4 i_131773694(.A(n_58388), .B(n_38929), .C(n_58464), .D(n_39891
		), .Z(n_139793018));
	notech_ao4 i_131673695(.A(n_58388), .B(n_38927), .C(n_58464), .D(n_39890
		), .Z(n_139893019));
	notech_ao4 i_131573696(.A(n_58388), .B(n_38925), .C(n_58464), .D(n_39889
		), .Z(n_139993020));
	notech_ao4 i_131473697(.A(n_58388), .B(n_38923), .C(n_58464), .D(n_39888
		), .Z(n_140093021));
	notech_ao4 i_131373698(.A(n_58389), .B(n_38921), .C(n_58464), .D(n_39887
		), .Z(n_140193022));
	notech_ao4 i_129873713(.A(n_58389), .B(n_38890), .C(n_58464), .D(n_39871
		), .Z(n_140293023));
	notech_ao4 i_129673715(.A(n_58389), .B(n_38886), .C(n_58465), .D(n_39869
		), .Z(n_140393024));
	notech_ao4 i_129573716(.A(n_58389), .B(n_38884), .C(n_58465), .D(n_39868
		), .Z(n_140493025));
	notech_ao4 i_129373718(.A(n_58389), .B(n_38879), .C(n_58465), .D(n_39865
		), .Z(n_140593026));
	notech_ao4 i_129273719(.A(n_58389), .B(n_38877), .C(n_58465), .D(n_39864
		), .Z(n_140693027));
	notech_ao4 i_129173720(.A(n_58389), .B(n_38875), .C(n_58465), .D(n_39863
		), .Z(n_140793028));
	notech_ao4 i_129073721(.A(n_58391), .B(n_38873), .C(n_58465), .D(n_39862
		), .Z(n_140893029));
	notech_nand3 i_16973207(.A(n_162393244), .B(n_162293243), .C(n_160493225
		), .Z(n_141093031));
	notech_ao4 i_16773209(.A(n_40209), .B(n_5299), .C(n_9089), .D(n_2218), .Z
		(n_155193172));
	notech_ao4 i_1273364(.A(n_38508), .B(n_2219), .C(n_5761), .D(n_1996), .Z
		(n_160393224));
	notech_nand2 i_71972664(.A(fpu), .B(n_38517), .Z(n_160493225));
	notech_and2 i_288992651(.A(lenpc1[7]), .B(n_58407), .Z(n_160793228));
	notech_or4 i_66272721(.A(n_251191358), .B(n_1249153), .C(n_261391460), .D
		(n_5674), .Z(n_160893229));
	notech_or2 i_66372720(.A(n_5304), .B(n_155193172), .Z(n_160993230));
	notech_ao3 i_3519(.A(int_excl[5]), .B(n_260791454), .C(n_2058), .Z(n_161193232
		));
	notech_and2 i_3525(.A(ififo_rvect3[0]), .B(n_162893249), .Z(n_161293233)
		);
	notech_and2 i_3530(.A(ififo_rvect3[1]), .B(n_162893249), .Z(n_161393234)
		);
	notech_and2 i_3531(.A(ififo_rvect3[2]), .B(n_162893249), .Z(n_161493235)
		);
	notech_and2 i_3532(.A(ififo_rvect3[3]), .B(n_162893249), .Z(n_161593236)
		);
	notech_and2 i_3533(.A(ififo_rvect3[4]), .B(n_162893249), .Z(n_161693237)
		);
	notech_and2 i_3534(.A(ififo_rvect3[5]), .B(n_162893249), .Z(n_161793238)
		);
	notech_and2 i_3535(.A(ififo_rvect3[6]), .B(n_162893249), .Z(n_161893239)
		);
	notech_and2 i_3536(.A(ififo_rvect3[7]), .B(n_162893249), .Z(n_161993240)
		);
	notech_ao3 i_3780(.A(n_1987), .B(n_38516), .C(n_1249153), .Z(n_162093241
		));
	notech_and3 i_3784(.A(db67), .B(n_41571), .C(n_141093031), .Z(n_162193242
		));
	notech_nao3 i_71772666(.A(n_1987), .B(n_38508), .C(n_5717), .Z(n_162293243
		));
	notech_nand3 i_71872665(.A(n_160393224), .B(\to_acu2_0[0] ), .C(\to_acu2_0[1] 
		), .Z(n_162393244));
	notech_ao3 i_3793(.A(n_59607), .B(in128[17]), .C(n_2849), .Z(n_162493245
		));
	notech_ao3 i_3799(.A(n_59596), .B(\to_acu2_0[3] ), .C(n_2849), .Z(n_162593246
		));
	notech_ao3 i_3801(.A(n_59596), .B(\to_acu2_0[7] ), .C(n_2849), .Z(n_162693247
		));
	notech_or4 i_3526(.A(intff), .B(trig_it), .C(n_38606), .D(n_40215), .Z(n_162793248
		));
	notech_nand2 i_210220(.A(trig_it), .B(n_38605), .Z(n_162893249));
	notech_xor2 i_35592652(.A(pfx_sz[2]), .B(n_170393324), .Z(n_163793258)
		);
	notech_xor2 i_35692653(.A(pfx_sz[3]), .B(n_170493325), .Z(n_163893259)
		);
	notech_xor2 i_35792654(.A(pfx_sz[4]), .B(n_170593326), .Z(n_163993260)
		);
	notech_xor2 i_36792655(.A(int_excl[1]), .B(int_excl[0]), .Z(n_164093261)
		);
	notech_xor2 i_36892656(.A(int_excl[3]), .B(n_1821), .Z(n_164193262));
	notech_ao4 i_4527781(.A(n_57481), .B(n_38504), .C(n_53788), .D(n_39605),
		 .Z(n_46387));
	notech_ao4 i_4127777(.A(n_57484), .B(n_38500), .C(n_53788), .D(n_39615),
		 .Z(n_46363));
	notech_ao4 i_4027776(.A(n_57484), .B(n_38499), .C(n_53727), .D(n_39619),
		 .Z(n_46357));
	notech_ao4 i_3927775(.A(n_57484), .B(n_38498), .C(n_53727), .D(n_39625),
		 .Z(n_46351));
	notech_ao4 i_3827774(.A(n_57484), .B(n_38497), .C(n_53727), .D(n_39632),
		 .Z(n_46345));
	notech_or2 i_327191(.A(n_5392), .B(n_168093301), .Z(n_49900));
	notech_and4 i_222716(.A(n_58835), .B(n_2833), .C(n_59596), .D(n_40105), 
		.Z(n_44589));
	notech_and4 i_129592667(.A(n_38325), .B(adz), .C(n_40184), .D(n_38326), 
		.Z(n_165293273));
	notech_xor2 i_34192668(.A(opz[1]), .B(opz[2]), .Z(n_165393274));
	notech_and3 i_129392669(.A(twobyte), .B(\to_acu2_0[16] ), .C(n_41571), .Z
		(n_165493275));
	notech_and4 i_129692670(.A(n_41571), .B(n_168193302), .C(n_1972), .D(n_165393274
		), .Z(n_165593276));
	notech_ao3 i_129492671(.A(opz[2]), .B(n_38325), .C(n_1810), .Z(n_165693277
		));
	notech_or4 i_323175(.A(n_165593276), .B(n_165493275), .C(n_165693277), .D
		(n_165293273), .Z(n_49828));
	notech_or4 i_130792672(.A(adz), .B(\to_acu2_0[73] ), .C(n_168393304), .D
		(n_168593306), .Z(n_165793278));
	notech_or4 i_130492673(.A(twobyte), .B(n_2812), .C(n_40121), .D(n_39117)
		, .Z(n_165893279));
	notech_nao3 i_130592674(.A(n_1972), .B(n_40105), .C(n_168293303), .Z(n_165993280
		));
	notech_or4 i_130692675(.A(n_1972), .B(n_168293303), .C(n_40105), .D(n_1810
		), .Z(n_166093281));
	notech_and4 i_223174(.A(n_165893279), .B(n_166093281), .C(n_165793278), 
		.D(n_165993280), .Z(n_49822));
	notech_or4 i_131692676(.A(n_1972), .B(n_168293303), .C(\to_acu2_0[73] ),
		 .D(n_40211), .Z(n_166193282));
	notech_nand3 i_34292677(.A(n_1810), .B(n_40185), .C(n_40183), .Z(n_166293283
		));
	notech_nao3 i_131592678(.A(n_59596), .B(n_1787), .C(n_2849), .Z(n_166393284
		));
	notech_nao3 i_131792679(.A(opz[0]), .B(n_166293283), .C(n_168293303), .Z
		(n_166493285));
	notech_nand3 i_123173(.A(n_166493285), .B(n_166393284), .C(n_166193282),
		 .Z(n_49816));
	notech_or4 i_134092680(.A(n_58835), .B(pc_req), .C(pg_fault), .D(n_166693287
		), .Z(n_166593286));
	notech_xor2 i_34792681(.A(n_38656), .B(idx_deco[1]), .Z(n_166693287));
	notech_nao3 i_133992682(.A(idx_deco[1]), .B(idx_deco[0]), .C(n_58394), .Z
		(n_166793288));
	notech_nand3 i_222702(.A(n_2056), .B(n_166793288), .C(n_166593286), .Z(n_41687
		));
	notech_or4 i_134392683(.A(n_58835), .B(pc_req), .C(pg_fault), .D(n_1994)
		, .Z(n_166893289));
	notech_nao3 i_134492684(.A(idx_deco[1]), .B(n_38656), .C(n_58394), .Z(n_166993290
		));
	notech_nand3 i_122701(.A(n_2056), .B(n_166993290), .C(n_166893289), .Z(n_41681
		));
	notech_or4 i_139192685(.A(n_58831), .B(pc_req), .C(pg_fault), .D(n_39866
		), .Z(n_167093291));
	notech_nao3 i_139292686(.A(inst_deco1[4]), .B(n_2847), .C(n_1995), .Z(n_167193292
		));
	notech_nand3 i_525656(.A(n_59695), .B(n_167193292), .C(n_167093291), .Z(n_45273
		));
	notech_ao4 i_226977(.A(n_39117), .B(n_170693327), .C(n_170793328), .D(n_40103
		), .Z(n_41904));
	notech_xor2 i_128092695(.A(int_excl[2]), .B(n_1801), .Z(n_168093301));
	notech_ao3 i_129092696(.A(n_40121), .B(n_40210), .C(n_2812), .Z(n_168193302
		));
	notech_nao3 i_17092697(.A(n_168193302), .B(n_59596), .C(n_2849), .Z(n_168293303
		));
	notech_nao3 i_20792698(.A(n_40185), .B(n_40183), .C(n_168293303), .Z(n_168393304
		));
	notech_nand3 i_29192700(.A(n_2819), .B(n_2816), .C(n_40211), .Z(n_168593306
		));
	notech_and2 i_295192718(.A(pfx_sz[0]), .B(pfx_sz[1]), .Z(n_170393324));
	notech_and3 i_1492719(.A(pfx_sz[0]), .B(pfx_sz[2]), .C(pfx_sz[1]), .Z(n_170493325
		));
	notech_and4 i_35992720(.A(pfx_sz[1]), .B(pfx_sz[0]), .C(pfx_sz[2]), .D(pfx_sz
		[3]), .Z(n_170593326));
	notech_nand2 i_140392721(.A(pfx_sz[0]), .B(n_40103), .Z(n_170693327));
	notech_nao3 i_73401(.A(n_18050174), .B(n_1568), .C(n_108292703), .Z(n_46591
		));
	notech_nao3 i_72360(.A(n_18050174), .B(n_1568), .C(n_108192702), .Z(\nbus_13550[1] 
		));
	notech_nao3 i_70966(.A(n_18050174), .B(n_1568), .C(n_17550169), .Z(\nbus_13541[0] 
		));
	notech_mux2 i_122086(.S(n_60686), .A(lenpc[0]), .B(lenpc1[0]), .Z(lenpc_out
		[0]));
	notech_mux2 i_222087(.S(n_60686), .A(lenpc[1]), .B(lenpc1[1]), .Z(lenpc_out
		[1]));
	notech_mux2 i_322088(.S(n_60680), .A(lenpc[2]), .B(lenpc1[2]), .Z(lenpc_out
		[2]));
	notech_mux2 i_422089(.S(n_60680), .A(lenpc[3]), .B(lenpc1[3]), .Z(lenpc_out
		[3]));
	notech_mux2 i_522090(.S(n_60680), .A(lenpc[4]), .B(lenpc1[4]), .Z(lenpc_out
		[4]));
	notech_mux2 i_622091(.S(n_60686), .A(lenpc[5]), .B(lenpc1[5]), .Z(lenpc_out
		[5]));
	notech_mux2 i_722092(.S(n_60686), .A(lenpc[6]), .B(lenpc1[6]), .Z(lenpc_out
		[6]));
	notech_mux2 i_822093(.S(n_60686), .A(lenpc[7]), .B(lenpc1[7]), .Z(lenpc_out
		[7]));
	notech_mux2 i_922094(.S(n_60686), .A(lenpc[8]), .B(lenpc1[8]), .Z(lenpc_out
		[8]));
	notech_mux2 i_1022095(.S(n_60686), .A(lenpc[9]), .B(lenpc1[9]), .Z(lenpc_out
		[9]));
	notech_mux2 i_1122096(.S(n_60686), .A(lenpc[10]), .B(lenpc1[10]), .Z(lenpc_out
		[10]));
	notech_mux2 i_1222097(.S(n_60686), .A(lenpc[11]), .B(lenpc1[11]), .Z(lenpc_out
		[11]));
	notech_mux2 i_1322098(.S(n_60680), .A(lenpc[12]), .B(lenpc1[12]), .Z(lenpc_out
		[12]));
	notech_mux2 i_1422099(.S(n_60680), .A(lenpc[13]), .B(lenpc1[13]), .Z(lenpc_out
		[13]));
	notech_mux2 i_1522100(.S(n_60680), .A(lenpc[14]), .B(lenpc1[14]), .Z(lenpc_out
		[14]));
	notech_mux2 i_1622101(.S(n_60680), .A(lenpc[15]), .B(lenpc1[15]), .Z(lenpc_out
		[15]));
	notech_mux2 i_1722102(.S(n_60680), .A(lenpc[16]), .B(lenpc1[16]), .Z(lenpc_out
		[16]));
	notech_mux2 i_1822103(.S(n_60680), .A(lenpc[17]), .B(lenpc1[17]), .Z(lenpc_out
		[17]));
	notech_mux2 i_1922104(.S(n_60680), .A(lenpc[18]), .B(lenpc1[18]), .Z(lenpc_out
		[18]));
	notech_mux2 i_2022105(.S(n_60680), .A(lenpc[19]), .B(lenpc1[19]), .Z(lenpc_out
		[19]));
	notech_mux2 i_2122106(.S(n_60680), .A(lenpc[20]), .B(lenpc1[20]), .Z(lenpc_out
		[20]));
	notech_mux2 i_2222107(.S(n_60680), .A(lenpc[21]), .B(lenpc1[21]), .Z(lenpc_out
		[21]));
	notech_mux2 i_2322108(.S(n_60680), .A(lenpc[22]), .B(lenpc1[22]), .Z(lenpc_out
		[22]));
	notech_mux2 i_2422109(.S(n_60680), .A(lenpc[23]), .B(lenpc1[23]), .Z(lenpc_out
		[23]));
	notech_mux2 i_2522110(.S(n_60680), .A(lenpc[24]), .B(lenpc1[24]), .Z(lenpc_out
		[24]));
	notech_mux2 i_2622111(.S(n_60686), .A(lenpc[25]), .B(lenpc1[25]), .Z(lenpc_out
		[25]));
	notech_mux2 i_2722112(.S(n_60691), .A(lenpc[26]), .B(lenpc1[26]), .Z(lenpc_out
		[26]));
	notech_mux2 i_2822113(.S(n_60691), .A(lenpc[27]), .B(lenpc1[27]), .Z(lenpc_out
		[27]));
	notech_mux2 i_2922114(.S(n_60691), .A(lenpc[28]), .B(lenpc1[28]), .Z(lenpc_out
		[28]));
	notech_mux2 i_3022115(.S(n_60691), .A(lenpc[29]), .B(lenpc1[29]), .Z(lenpc_out
		[29]));
	notech_mux2 i_3122116(.S(n_60691), .A(lenpc[30]), .B(lenpc1[30]), .Z(lenpc_out
		[30]));
	notech_mux2 i_3222117(.S(n_60691), .A(lenpc[31]), .B(lenpc1[31]), .Z(lenpc_out
		[31]));
	notech_mux2 i_123119(.S(n_60692), .A(reps0[0]), .B(reps1[0]), .Z(reps[0]
		));
	notech_mux2 i_223120(.S(n_60692), .A(reps0[1]), .B(reps1[1]), .Z(reps[1]
		));
	notech_mux2 i_323121(.S(n_60692), .A(reps0[2]), .B(reps1[2]), .Z(reps[2]
		));
	notech_mux2 i_123122(.S(n_60692), .A(opz0[0]), .B(opz1[0]), .Z(operand_size
		[0]));
	notech_mux2 i_223123(.S(n_60692), .A(opz0[1]), .B(opz1[1]), .Z(operand_size
		[1]));
	notech_mux2 i_323124(.S(n_60692), .A(opz0[2]), .B(opz1[2]), .Z(operand_size
		[2]));
	notech_mux2 i_125268(.S(n_60692), .A(inst_deco[0]), .B(inst_deco1[0]), .Z
		(to_vliw[0]));
	notech_mux2 i_225269(.S(n_60691), .A(inst_deco[1]), .B(inst_deco1[1]), .Z
		(to_vliw[1]));
	notech_mux2 i_325270(.S(n_60691), .A(inst_deco[2]), .B(inst_deco1[2]), .Z
		(to_vliw[2]));
	notech_mux2 i_425271(.S(n_60691), .A(inst_deco[3]), .B(inst_deco1[3]), .Z
		(to_vliw[3]));
	notech_mux2 i_525272(.S(n_60686), .A(inst_deco[4]), .B(inst_deco1[4]), .Z
		(to_vliw[4]));
	notech_mux2 i_625273(.S(n_60691), .A(inst_deco[5]), .B(inst_deco1[5]), .Z
		(to_vliw[5]));
	notech_mux2 i_725274(.S(n_60691), .A(inst_deco[6]), .B(inst_deco1[6]), .Z
		(to_vliw[6]));
	notech_mux2 i_825275(.S(n_60691), .A(inst_deco[7]), .B(inst_deco1[7]), .Z
		(to_vliw[7]));
	notech_mux2 i_925276(.S(n_60691), .A(inst_deco[8]), .B(inst_deco1[8]), .Z
		(to_vliw[8]));
	notech_mux2 i_1025277(.S(n_60691), .A(inst_deco[9]), .B(inst_deco1[9]), 
		.Z(to_vliw[9]));
	notech_mux2 i_1125278(.S(n_60691), .A(inst_deco[10]), .B(inst_deco1[10])
		, .Z(to_vliw[10]));
	notech_mux2 i_1225279(.S(n_60691), .A(inst_deco[11]), .B(inst_deco1[11])
		, .Z(to_vliw[11]));
	notech_mux2 i_1325280(.S(n_60691), .A(inst_deco[12]), .B(inst_deco1[12])
		, .Z(to_vliw[12]));
	notech_mux2 i_1425281(.S(n_60691), .A(inst_deco[13]), .B(inst_deco1[13])
		, .Z(to_vliw[13]));
	notech_mux2 i_1525282(.S(n_60680), .A(inst_deco[14]), .B(inst_deco1[14])
		, .Z(to_vliw[14]));
	notech_mux2 i_1625283(.S(n_60669), .A(inst_deco[15]), .B(inst_deco1[15])
		, .Z(to_vliw[15]));
	notech_mux2 i_1725284(.S(n_60669), .A(inst_deco[16]), .B(inst_deco1[16])
		, .Z(to_vliw[16]));
	notech_mux2 i_1825285(.S(n_60669), .A(inst_deco[17]), .B(inst_deco1[17])
		, .Z(to_vliw[17]));
	notech_mux2 i_1925286(.S(n_60669), .A(inst_deco[18]), .B(inst_deco1[18])
		, .Z(to_vliw[18]));
	notech_mux2 i_2025287(.S(n_60669), .A(inst_deco[19]), .B(inst_deco1[19])
		, .Z(to_vliw[19]));
	notech_mux2 i_2125288(.S(n_60669), .A(inst_deco[20]), .B(inst_deco1[20])
		, .Z(to_vliw[20]));
	notech_mux2 i_2225289(.S(n_60669), .A(inst_deco[21]), .B(inst_deco1[21])
		, .Z(to_vliw[21]));
	notech_mux2 i_2325290(.S(n_60674), .A(inst_deco[22]), .B(inst_deco1[22])
		, .Z(to_vliw[22]));
	notech_mux2 i_2425291(.S(n_60674), .A(inst_deco[23]), .B(inst_deco1[23])
		, .Z(to_vliw[23]));
	notech_mux2 i_2525292(.S(n_60674), .A(inst_deco[24]), .B(inst_deco1[24])
		, .Z(to_vliw[24]));
	notech_mux2 i_2625293(.S(n_60669), .A(inst_deco[25]), .B(inst_deco1[25])
		, .Z(to_vliw[25]));
	notech_mux2 i_2725294(.S(n_60669), .A(inst_deco[26]), .B(inst_deco1[26])
		, .Z(to_vliw[26]));
	notech_mux2 i_2825295(.S(n_60674), .A(inst_deco[27]), .B(inst_deco1[27])
		, .Z(to_vliw[27]));
	notech_mux2 i_2925296(.S(n_60668), .A(inst_deco[28]), .B(inst_deco1[28])
		, .Z(to_vliw[28]));
	notech_mux2 i_3025297(.S(n_60669), .A(inst_deco[29]), .B(inst_deco1[29])
		, .Z(to_vliw[29]));
	notech_mux2 i_3125298(.S(n_60669), .A(inst_deco[30]), .B(inst_deco1[30])
		, .Z(to_vliw[30]));
	notech_mux2 i_3225299(.S(n_60668), .A(inst_deco[31]), .B(inst_deco1[31])
		, .Z(to_vliw[31]));
	notech_mux2 i_3325300(.S(n_60668), .A(inst_deco[32]), .B(inst_deco1[32])
		, .Z(to_vliw[32]));
	notech_mux2 i_3425301(.S(n_60668), .A(inst_deco[33]), .B(inst_deco1[33])
		, .Z(to_vliw[33]));
	notech_mux2 i_3525302(.S(n_60669), .A(inst_deco[34]), .B(inst_deco1[34])
		, .Z(to_vliw[34]));
	notech_mux2 i_3625303(.S(n_60669), .A(inst_deco[35]), .B(inst_deco1[35])
		, .Z(to_vliw[35]));
	notech_mux2 i_3725304(.S(n_60669), .A(inst_deco[36]), .B(inst_deco1[36])
		, .Z(to_vliw[36]));
	notech_mux2 i_3825305(.S(n_60669), .A(inst_deco[37]), .B(inst_deco1[37])
		, .Z(to_vliw[37]));
	notech_mux2 i_3925306(.S(n_60669), .A(inst_deco[38]), .B(inst_deco1[38])
		, .Z(to_vliw[38]));
	notech_mux2 i_4025307(.S(n_60669), .A(inst_deco[39]), .B(inst_deco1[39])
		, .Z(to_vliw[39]));
	notech_mux2 i_4125308(.S(n_60669), .A(inst_deco[40]), .B(inst_deco1[40])
		, .Z(to_vliw[40]));
	notech_mux2 i_4225309(.S(n_60674), .A(inst_deco[41]), .B(inst_deco1[41])
		, .Z(to_vliw[41]));
	notech_mux2 i_4325310(.S(n_60679), .A(inst_deco[42]), .B(inst_deco1[42])
		, .Z(to_vliw[42]));
	notech_mux2 i_4425311(.S(n_60679), .A(inst_deco[43]), .B(inst_deco1[43])
		, .Z(to_vliw[43]));
	notech_mux2 i_4525312(.S(n_60679), .A(inst_deco[44]), .B(inst_deco1[44])
		, .Z(to_vliw[44]));
	notech_mux2 i_4625313(.S(n_60679), .A(inst_deco[45]), .B(inst_deco1[45])
		, .Z(to_vliw[45]));
	notech_mux2 i_4725314(.S(n_60679), .A(inst_deco[46]), .B(inst_deco1[46])
		, .Z(to_vliw[46]));
	notech_mux2 i_4825315(.S(n_60679), .A(inst_deco[47]), .B(inst_deco1[47])
		, .Z(to_vliw[47]));
	notech_mux2 i_4925316(.S(n_60679), .A(inst_deco[48]), .B(inst_deco1[48])
		, .Z(to_vliw[48]));
	notech_mux2 i_5025317(.S(n_60679), .A(inst_deco[49]), .B(inst_deco1[49])
		, .Z(to_vliw[49]));
	notech_mux2 i_5125318(.S(n_60679), .A(inst_deco[50]), .B(inst_deco1[50])
		, .Z(to_vliw[50]));
	notech_mux2 i_5225319(.S(n_60680), .A(inst_deco[51]), .B(inst_deco1[51])
		, .Z(to_vliw[51]));
	notech_mux2 i_5325320(.S(n_60679), .A(inst_deco[52]), .B(inst_deco1[52])
		, .Z(to_vliw[52]));
	notech_mux2 i_5425321(.S(n_60679), .A(inst_deco[53]), .B(inst_deco1[53])
		, .Z(to_vliw[53]));
	notech_mux2 i_5525322(.S(n_60679), .A(inst_deco[54]), .B(inst_deco1[54])
		, .Z(to_vliw[54]));
	notech_mux2 i_5625323(.S(n_60674), .A(inst_deco[55]), .B(inst_deco1[55])
		, .Z(to_vliw[55]));
	notech_mux2 i_5725324(.S(n_60674), .A(inst_deco[56]), .B(inst_deco1[56])
		, .Z(to_vliw[56]));
	notech_mux2 i_5825325(.S(n_60674), .A(inst_deco[57]), .B(inst_deco1[57])
		, .Z(to_vliw[57]));
	notech_mux2 i_5925326(.S(n_60674), .A(inst_deco[58]), .B(inst_deco1[58])
		, .Z(to_vliw[58]));
	notech_mux2 i_6025327(.S(n_60674), .A(inst_deco[59]), .B(inst_deco1[59])
		, .Z(to_vliw[59]));
	notech_mux2 i_6125328(.S(n_60674), .A(inst_deco[60]), .B(inst_deco1[60])
		, .Z(to_vliw[60]));
	notech_mux2 i_6225329(.S(n_60674), .A(inst_deco[61]), .B(inst_deco1[61])
		, .Z(to_vliw[61]));
	notech_mux2 i_6325330(.S(n_60679), .A(inst_deco[62]), .B(inst_deco1[62])
		, .Z(to_vliw[62]));
	notech_mux2 i_6425331(.S(n_60679), .A(inst_deco[63]), .B(inst_deco1[63])
		, .Z(to_vliw[63]));
	notech_mux2 i_6525332(.S(n_60679), .A(inst_deco[64]), .B(inst_deco1[64])
		, .Z(to_vliw[64]));
	notech_mux2 i_6625333(.S(n_60679), .A(inst_deco[65]), .B(inst_deco1[65])
		, .Z(to_vliw[65]));
	notech_mux2 i_6725334(.S(n_60679), .A(inst_deco[66]), .B(inst_deco1[66])
		, .Z(to_vliw[66]));
	notech_mux2 i_6825335(.S(n_60679), .A(inst_deco[67]), .B(inst_deco1[67])
		, .Z(to_vliw[67]));
	notech_mux2 i_6925336(.S(n_60708), .A(inst_deco[68]), .B(inst_deco1[68])
		, .Z(to_vliw[68]));
	notech_mux2 i_7025337(.S(n_60713), .A(inst_deco[69]), .B(inst_deco1[69])
		, .Z(to_vliw[69]));
	notech_mux2 i_7125338(.S(n_60713), .A(inst_deco[70]), .B(inst_deco1[70])
		, .Z(to_vliw[70]));
	notech_mux2 i_7225339(.S(n_60708), .A(inst_deco[71]), .B(inst_deco1[71])
		, .Z(to_vliw[71]));
	notech_mux2 i_7325340(.S(n_60708), .A(inst_deco[72]), .B(inst_deco1[72])
		, .Z(to_vliw[72]));
	notech_mux2 i_7425341(.S(n_60708), .A(inst_deco[73]), .B(inst_deco1[73])
		, .Z(to_vliw[73]));
	notech_mux2 i_7525342(.S(n_60713), .A(inst_deco[74]), .B(inst_deco1[74])
		, .Z(to_vliw[74]));
	notech_mux2 i_7625343(.S(n_60713), .A(inst_deco[75]), .B(inst_deco1[75])
		, .Z(to_vliw[75]));
	notech_mux2 i_7725344(.S(n_60713), .A(inst_deco[76]), .B(inst_deco1[76])
		, .Z(to_vliw[76]));
	notech_mux2 i_7825345(.S(n_60713), .A(inst_deco[77]), .B(inst_deco1[77])
		, .Z(to_vliw[77]));
	notech_mux2 i_7925346(.S(n_60713), .A(inst_deco[78]), .B(inst_deco1[78])
		, .Z(to_vliw[78]));
	notech_mux2 i_8025347(.S(n_60713), .A(inst_deco[79]), .B(inst_deco1[79])
		, .Z(to_vliw[79]));
	notech_mux2 i_8125348(.S(n_60713), .A(inst_deco[80]), .B(inst_deco1[80])
		, .Z(to_vliw[80]));
	notech_mux2 i_8225349(.S(n_60703), .A(inst_deco[81]), .B(inst_deco1[81])
		, .Z(to_vliw[81]));
	notech_mux2 i_8325350(.S(n_60703), .A(inst_deco[82]), .B(inst_deco1[82])
		, .Z(to_vliw[82]));
	notech_mux2 i_8425351(.S(n_60708), .A(inst_deco[83]), .B(inst_deco1[83])
		, .Z(to_vliw[83]));
	notech_mux2 i_8525352(.S(n_60703), .A(inst_deco[84]), .B(inst_deco1[84])
		, .Z(to_vliw[84]));
	notech_mux2 i_8625353(.S(n_60703), .A(inst_deco[85]), .B(inst_deco1[85])
		, .Z(to_vliw[85]));
	notech_mux2 i_8725354(.S(n_60703), .A(inst_deco[86]), .B(inst_deco1[86])
		, .Z(to_vliw[86]));
	notech_mux2 i_8825355(.S(n_60708), .A(inst_deco[87]), .B(inst_deco1[87])
		, .Z(to_vliw[87]));
	notech_mux2 i_8925356(.S(n_60708), .A(inst_deco[88]), .B(inst_deco1[88])
		, .Z(to_vliw[88]));
	notech_mux2 i_9025357(.S(n_60708), .A(inst_deco[89]), .B(inst_deco1[89])
		, .Z(to_vliw[89]));
	notech_mux2 i_9125358(.S(n_60708), .A(inst_deco[90]), .B(inst_deco1[90])
		, .Z(to_vliw[90]));
	notech_mux2 i_9225359(.S(n_60708), .A(inst_deco[91]), .B(inst_deco1[91])
		, .Z(to_vliw[91]));
	notech_mux2 i_9325360(.S(n_60708), .A(inst_deco[92]), .B(inst_deco1[92])
		, .Z(to_vliw[92]));
	notech_mux2 i_9425361(.S(n_60708), .A(inst_deco[93]), .B(inst_deco1[93])
		, .Z(to_vliw[93]));
	notech_mux2 i_9525362(.S(n_60713), .A(inst_deco[94]), .B(inst_deco1[94])
		, .Z(to_vliw[94]));
	notech_mux2 i_9625363(.S(n_60714), .A(inst_deco[95]), .B(inst_deco1[95])
		, .Z(to_vliw[95]));
	notech_mux2 i_9725364(.S(n_60714), .A(inst_deco[96]), .B(inst_deco1[96])
		, .Z(to_vliw[96]));
	notech_mux2 i_9825365(.S(n_60714), .A(inst_deco[97]), .B(inst_deco1[97])
		, .Z(to_vliw[97]));
	notech_mux2 i_9925366(.S(n_60714), .A(inst_deco[98]), .B(inst_deco1[98])
		, .Z(to_vliw[98]));
	notech_mux2 i_10025367(.S(n_60714), .A(inst_deco[99]), .B(inst_deco1[99]
		), .Z(to_vliw[99]));
	notech_mux2 i_10125368(.S(n_60714), .A(inst_deco[100]), .B(inst_deco1[
		100]), .Z(to_vliw[100]));
	notech_mux2 i_10225369(.S(n_60714), .A(inst_deco[101]), .B(inst_deco1[
		101]), .Z(to_vliw[101]));
	notech_mux2 i_10325370(.S(n_60714), .A(inst_deco[102]), .B(inst_deco1[
		102]), .Z(to_vliw[102]));
	notech_mux2 i_10425371(.S(n_60714), .A(inst_deco[103]), .B(inst_deco1[
		103]), .Z(to_vliw[103]));
	notech_mux2 i_10525372(.S(n_60714), .A(inst_deco[104]), .B(inst_deco1[
		104]), .Z(to_vliw[104]));
	notech_mux2 i_10625373(.S(n_60714), .A(inst_deco[105]), .B(inst_deco1[
		105]), .Z(to_vliw[105]));
	notech_mux2 i_10725374(.S(n_60714), .A(inst_deco[106]), .B(inst_deco1[
		106]), .Z(to_vliw[106]));
	notech_mux2 i_10825375(.S(n_60714), .A(inst_deco[107]), .B(inst_deco1[
		107]), .Z(to_vliw[107]));
	notech_mux2 i_10925376(.S(n_60713), .A(inst_deco[108]), .B(inst_deco1[
		108]), .Z(to_vliw[108]));
	notech_mux2 i_11025377(.S(n_60713), .A(inst_deco[109]), .B(inst_deco1[
		109]), .Z(to_vliw[109]));
	notech_mux2 i_11125378(.S(n_60713), .A(inst_deco[110]), .B(inst_deco1[
		110]), .Z(to_vliw[110]));
	notech_mux2 i_11225379(.S(n_60713), .A(inst_deco[111]), .B(inst_deco1[
		111]), .Z(to_vliw[111]));
	notech_mux2 i_11325380(.S(n_60713), .A(inst_deco[112]), .B(inst_deco1[
		112]), .Z(to_vliw[112]));
	notech_mux2 i_11425381(.S(n_60713), .A(inst_deco[113]), .B(inst_deco1[
		113]), .Z(to_vliw[113]));
	notech_mux2 i_11525382(.S(n_60713), .A(inst_deco[114]), .B(inst_deco1[
		114]), .Z(to_vliw[114]));
	notech_mux2 i_11625383(.S(n_60714), .A(inst_deco[115]), .B(inst_deco1[
		115]), .Z(to_vliw[115]));
	notech_mux2 i_11725384(.S(n_60714), .A(inst_deco[116]), .B(inst_deco1[
		116]), .Z(to_vliw[116]));
	notech_mux2 i_11825385(.S(n_60714), .A(inst_deco[117]), .B(inst_deco1[
		117]), .Z(to_vliw[117]));
	notech_mux2 i_11925386(.S(n_60713), .A(inst_deco[118]), .B(inst_deco1[
		118]), .Z(to_vliw[118]));
	notech_mux2 i_12025387(.S(n_60714), .A(inst_deco[119]), .B(inst_deco1[
		119]), .Z(to_vliw[119]));
	notech_mux2 i_12125388(.S(n_60714), .A(inst_deco[120]), .B(inst_deco1[
		120]), .Z(to_vliw[120]));
	notech_mux2 i_12225389(.S(n_60703), .A(inst_deco[121]), .B(inst_deco1[
		121]), .Z(to_vliw[121]));
	notech_mux2 i_12325390(.S(n_60697), .A(inst_deco[122]), .B(inst_deco1[
		122]), .Z(to_vliw[122]));
	notech_mux2 i_12425391(.S(n_60697), .A(inst_deco[123]), .B(inst_deco1[
		123]), .Z(to_vliw[123]));
	notech_mux2 i_12525392(.S(n_60697), .A(inst_deco[124]), .B(inst_deco1[
		124]), .Z(to_vliw[124]));
	notech_mux2 i_12625393(.S(n_60697), .A(inst_deco[125]), .B(inst_deco1[
		125]), .Z(to_vliw[125]));
	notech_mux2 i_12725394(.S(n_60697), .A(inst_deco[126]), .B(inst_deco1[
		126]), .Z(to_vliw[126]));
	notech_mux2 i_12825395(.S(n_60697), .A(inst_deco[127]), .B(inst_deco1[
		127]), .Z(to_vliw[127]));
	notech_mux2 i_125908(.S(n_60697), .A(to_acu0[0]), .B(to_acu1[0]), .Z(to_acu
		[0]));
	notech_mux2 i_225909(.S(n_60702), .A(to_acu0[1]), .B(to_acu1[1]), .Z(to_acu
		[1]));
	notech_mux2 i_325910(.S(n_60702), .A(to_acu0[2]), .B(to_acu1[2]), .Z(to_acu
		[2]));
	notech_mux2 i_425911(.S(n_60702), .A(to_acu0[3]), .B(to_acu1[3]), .Z(to_acu
		[3]));
	notech_mux2 i_525912(.S(n_60697), .A(to_acu0[4]), .B(to_acu1[4]), .Z(to_acu
		[4]));
	notech_mux2 i_625913(.S(n_60697), .A(to_acu0[5]), .B(to_acu1[5]), .Z(to_acu
		[5]));
	notech_mux2 i_725914(.S(n_60697), .A(to_acu0[6]), .B(to_acu1[6]), .Z(to_acu
		[6]));
	notech_mux2 i_825915(.S(n_60692), .A(to_acu0[7]), .B(to_acu1[7]), .Z(to_acu
		[7]));
	notech_mux2 i_925916(.S(n_60692), .A(to_acu0[8]), .B(to_acu1[8]), .Z(to_acu
		[8]));
	notech_mux2 i_1025917(.S(n_60692), .A(to_acu0[9]), .B(to_acu1[9]), .Z(to_acu
		[9]));
	notech_mux2 i_1125918(.S(n_60692), .A(to_acu0[10]), .B(to_acu1[10]), .Z(to_acu
		[10]));
	notech_mux2 i_1225919(.S(n_60692), .A(to_acu0[11]), .B(to_acu1[11]), .Z(to_acu
		[11]));
	notech_mux2 i_1325920(.S(n_60692), .A(to_acu0[12]), .B(to_acu1[12]), .Z(to_acu
		[12]));
	notech_mux2 i_1425921(.S(n_60692), .A(to_acu0[13]), .B(to_acu1[13]), .Z(to_acu
		[13]));
	notech_mux2 i_1525922(.S(n_60692), .A(to_acu0[14]), .B(to_acu1[14]), .Z(to_acu
		[14]));
	notech_mux2 i_1625923(.S(n_60697), .A(to_acu0[15]), .B(to_acu1[15]), .Z(to_acu
		[15]));
	notech_mux2 i_1725924(.S(n_60697), .A(to_acu0[16]), .B(to_acu1[16]), .Z(to_acu
		[16]));
	notech_mux2 i_1825925(.S(n_60692), .A(to_acu0[17]), .B(to_acu1[17]), .Z(to_acu
		[17]));
	notech_mux2 i_1925926(.S(n_60692), .A(to_acu0[18]), .B(to_acu1[18]), .Z(to_acu
		[18]));
	notech_mux2 i_2025927(.S(n_60692), .A(to_acu0[19]), .B(to_acu1[19]), .Z(to_acu
		[19]));
	notech_mux2 i_2125928(.S(n_60702), .A(to_acu0[20]), .B(to_acu1[20]), .Z(to_acu
		[20]));
	notech_mux2 i_2225929(.S(n_60703), .A(to_acu0[21]), .B(to_acu1[21]), .Z(to_acu
		[21]));
	notech_mux2 i_2325930(.S(n_60703), .A(to_acu0[22]), .B(to_acu1[22]), .Z(to_acu
		[22]));
	notech_mux2 i_2425931(.S(n_60703), .A(to_acu0[23]), .B(to_acu1[23]), .Z(to_acu
		[23]));
	notech_mux2 i_2525932(.S(n_60702), .A(to_acu0[24]), .B(to_acu1[24]), .Z(to_acu
		[24]));
	notech_mux2 i_2625933(.S(n_60703), .A(to_acu0[25]), .B(to_acu1[25]), .Z(to_acu
		[25]));
	notech_mux2 i_2725934(.S(n_60703), .A(to_acu0[26]), .B(to_acu1[26]), .Z(to_acu
		[26]));
	notech_mux2 i_2825935(.S(n_60703), .A(to_acu0[27]), .B(to_acu1[27]), .Z(to_acu
		[27]));
	notech_mux2 i_2925936(.S(n_60703), .A(to_acu0[28]), .B(to_acu1[28]), .Z(to_acu
		[28]));
	notech_mux2 i_3025937(.S(n_60703), .A(to_acu0[29]), .B(to_acu1[29]), .Z(to_acu
		[29]));
	notech_mux2 i_3125938(.S(n_60703), .A(to_acu0[30]), .B(to_acu1[30]), .Z(to_acu
		[30]));
	notech_mux2 i_3225939(.S(n_60703), .A(to_acu0[31]), .B(to_acu1[31]), .Z(to_acu
		[31]));
	notech_mux2 i_3325940(.S(n_60703), .A(to_acu0[32]), .B(to_acu1[32]), .Z(to_acu
		[32]));
	notech_mux2 i_3425941(.S(n_60703), .A(to_acu0[33]), .B(to_acu1[33]), .Z(to_acu
		[33]));
	notech_mux2 i_3525942(.S(n_60702), .A(to_acu0[34]), .B(to_acu1[34]), .Z(to_acu
		[34]));
	notech_mux2 i_3625943(.S(n_60702), .A(to_acu0[35]), .B(to_acu1[35]), .Z(to_acu
		[35]));
	notech_mux2 i_3725944(.S(n_60702), .A(to_acu0[36]), .B(to_acu1[36]), .Z(to_acu
		[36]));
	notech_mux2 i_3825945(.S(n_60702), .A(to_acu0[37]), .B(to_acu1[37]), .Z(to_acu
		[37]));
	notech_mux2 i_3925946(.S(n_60702), .A(to_acu0[38]), .B(to_acu1[38]), .Z(to_acu
		[38]));
	notech_mux2 i_4025947(.S(n_60702), .A(to_acu0[39]), .B(to_acu1[39]), .Z(to_acu
		[39]));
	notech_mux2 i_4125948(.S(n_60702), .A(to_acu0[40]), .B(to_acu1[40]), .Z(to_acu
		[40]));
	notech_mux2 i_4225949(.S(n_60702), .A(to_acu0[41]), .B(to_acu1[41]), .Z(to_acu
		[41]));
	notech_mux2 i_4325950(.S(n_60702), .A(to_acu0[42]), .B(to_acu1[42]), .Z(to_acu
		[42]));
	notech_mux2 i_4425951(.S(n_60702), .A(to_acu0[43]), .B(to_acu1[43]), .Z(to_acu
		[43]));
	notech_mux2 i_4525952(.S(n_60702), .A(to_acu0[44]), .B(to_acu1[44]), .Z(to_acu
		[44]));
	notech_mux2 i_4625953(.S(n_60702), .A(to_acu0[45]), .B(to_acu1[45]), .Z(to_acu
		[45]));
	notech_mux2 i_4725954(.S(n_60702), .A(to_acu0[46]), .B(to_acu1[46]), .Z(to_acu
		[46]));
	notech_mux2 i_4825955(.S(n_60668), .A(to_acu0[47]), .B(to_acu1[47]), .Z(to_acu
		[47]));
	notech_mux2 i_4925956(.S(n_60634), .A(to_acu0[48]), .B(to_acu1[48]), .Z(to_acu
		[48]));
	notech_mux2 i_5025957(.S(n_60634), .A(to_acu0[49]), .B(to_acu1[49]), .Z(to_acu
		[49]));
	notech_mux2 i_5125958(.S(n_60634), .A(to_acu0[50]), .B(to_acu1[50]), .Z(to_acu
		[50]));
	notech_mux2 i_5225959(.S(n_60634), .A(to_acu0[51]), .B(to_acu1[51]), .Z(to_acu
		[51]));
	notech_mux2 i_5325960(.S(n_60634), .A(to_acu0[52]), .B(to_acu1[52]), .Z(to_acu
		[52]));
	notech_mux2 i_5425961(.S(n_60634), .A(to_acu0[53]), .B(to_acu1[53]), .Z(to_acu
		[53]));
	notech_mux2 i_5525962(.S(n_60634), .A(to_acu0[54]), .B(to_acu1[54]), .Z(to_acu
		[54]));
	notech_mux2 i_5625963(.S(n_60635), .A(to_acu0[55]), .B(to_acu1[55]), .Z(to_acu
		[55]));
	notech_mux2 i_5725964(.S(n_60635), .A(to_acu0[56]), .B(to_acu1[56]), .Z(to_acu
		[56]));
	notech_mux2 i_5825965(.S(n_60635), .A(to_acu0[57]), .B(to_acu1[57]), .Z(to_acu
		[57]));
	notech_mux2 i_5925966(.S(n_60634), .A(to_acu0[58]), .B(to_acu1[58]), .Z(to_acu
		[58]));
	notech_mux2 i_6025967(.S(n_60635), .A(to_acu0[59]), .B(to_acu1[59]), .Z(to_acu
		[59]));
	notech_mux2 i_6125968(.S(n_60635), .A(to_acu0[60]), .B(to_acu1[60]), .Z(to_acu
		[60]));
	notech_mux2 i_6225969(.S(n_60634), .A(to_acu0[61]), .B(to_acu1[61]), .Z(to_acu
		[61]));
	notech_mux2 i_6325970(.S(n_60634), .A(to_acu0[62]), .B(to_acu1[62]), .Z(to_acu
		[62]));
	notech_mux2 i_6425971(.S(n_60634), .A(to_acu0[63]), .B(to_acu1[63]), .Z(to_acu
		[63]));
	notech_mux2 i_6525972(.S(n_60629), .A(to_acu0[64]), .B(to_acu1[64]), .Z(to_acu
		[64]));
	notech_mux2 i_6625973(.S(n_60629), .A(to_acu0[65]), .B(to_acu1[65]), .Z(to_acu
		[65]));
	notech_mux2 i_6725974(.S(n_60629), .A(to_acu0[66]), .B(to_acu1[66]), .Z(to_acu
		[66]));
	notech_mux2 i_6825975(.S(n_60634), .A(to_acu0[67]), .B(to_acu1[67]), .Z(to_acu
		[67]));
	notech_mux2 i_6925976(.S(n_60634), .A(to_acu0[68]), .B(to_acu1[68]), .Z(to_acu
		[68]));
	notech_mux2 i_7025977(.S(n_60634), .A(to_acu0[69]), .B(to_acu1[69]), .Z(to_acu
		[69]));
	notech_mux2 i_7125978(.S(n_60634), .A(to_acu0[70]), .B(to_acu1[70]), .Z(to_acu
		[70]));
	notech_mux2 i_7225979(.S(n_60634), .A(to_acu0[71]), .B(to_acu1[71]), .Z(to_acu
		[71]));
	notech_mux2 i_7325980(.S(n_60634), .A(to_acu0[72]), .B(to_acu1[72]), .Z(to_acu
		[72]));
	notech_mux2 i_7425981(.S(n_60634), .A(to_acu0[73]), .B(to_acu1[73]), .Z(to_acu
		[73]));
	notech_mux2 i_7525982(.S(n_60635), .A(to_acu0[74]), .B(to_acu1[74]), .Z(to_acu
		[74]));
	notech_mux2 i_7625983(.S(n_60640), .A(to_acu0[75]), .B(to_acu1[75]), .Z(to_acu
		[75]));
	notech_mux2 i_7725984(.S(n_60640), .A(to_acu0[76]), .B(to_acu1[76]), .Z(to_acu
		[76]));
	notech_mux2 i_7825985(.S(n_60640), .A(to_acu0[77]), .B(to_acu1[77]), .Z(to_acu
		[77]));
	notech_mux2 i_7925986(.S(n_60640), .A(to_acu0[78]), .B(to_acu1[78]), .Z(to_acu
		[78]));
	notech_mux2 i_8025987(.S(n_60640), .A(to_acu0[79]), .B(to_acu1[79]), .Z(to_acu
		[79]));
	notech_mux2 i_8125988(.S(n_60640), .A(to_acu0[80]), .B(to_acu1[80]), .Z(to_acu
		[80]));
	notech_mux2 i_8225989(.S(n_60640), .A(to_acu0[81]), .B(to_acu1[81]), .Z(to_acu
		[81]));
	notech_mux2 i_8325990(.S(n_60640), .A(to_acu0[82]), .B(to_acu1[82]), .Z(to_acu
		[82]));
	notech_mux2 i_8425991(.S(n_60645), .A(to_acu0[83]), .B(to_acu1[83]), .Z(to_acu
		[83]));
	notech_mux2 i_8525992(.S(n_60645), .A(to_acu0[84]), .B(to_acu1[84]), .Z(to_acu
		[84]));
	notech_mux2 i_8625993(.S(n_60640), .A(to_acu0[85]), .B(to_acu1[85]), .Z(to_acu
		[85]));
	notech_mux2 i_8725994(.S(n_60640), .A(to_acu0[86]), .B(to_acu1[86]), .Z(to_acu
		[86]));
	notech_mux2 i_8825995(.S(n_60640), .A(to_acu0[87]), .B(to_acu1[87]), .Z(to_acu
		[87]));
	notech_mux2 i_8925996(.S(n_60635), .A(to_acu0[88]), .B(to_acu1[88]), .Z(to_acu
		[88]));
	notech_mux2 i_9025997(.S(n_60635), .A(to_acu0[89]), .B(to_acu1[89]), .Z(to_acu
		[89]));
	notech_mux2 i_9125998(.S(n_60635), .A(to_acu0[90]), .B(to_acu1[90]), .Z(to_acu
		[90]));
	notech_mux2 i_9225999(.S(n_60635), .A(to_acu0[91]), .B(to_acu1[91]), .Z(to_acu
		[91]));
	notech_mux2 i_9326000(.S(n_60635), .A(to_acu0[92]), .B(to_acu1[92]), .Z(to_acu
		[92]));
	notech_mux2 i_9426001(.S(n_60635), .A(to_acu0[93]), .B(to_acu1[93]), .Z(to_acu
		[93]));
	notech_mux2 i_9526002(.S(n_60635), .A(to_acu0[94]), .B(to_acu1[94]), .Z(to_acu
		[94]));
	notech_mux2 i_9626003(.S(n_60635), .A(to_acu0[95]), .B(to_acu1[95]), .Z(to_acu
		[95]));
	notech_mux2 i_9726004(.S(n_60635), .A(to_acu0[96]), .B(to_acu1[96]), .Z(to_acu
		[96]));
	notech_mux2 i_9826005(.S(n_60640), .A(to_acu0[97]), .B(to_acu1[97]), .Z(to_acu
		[97]));
	notech_mux2 i_9926006(.S(n_60635), .A(to_acu0[98]), .B(to_acu1[98]), .Z(to_acu
		[98]));
	notech_mux2 i_10026007(.S(n_60635), .A(to_acu0[99]), .B(to_acu1[99]), .Z
		(to_acu[99]));
	notech_mux2 i_10126008(.S(n_60635), .A(to_acu0[100]), .B(to_acu1[100]), 
		.Z(to_acu[100]));
	notech_mux2 i_10226009(.S(n_60629), .A(to_acu0[101]), .B(to_acu1[101]), 
		.Z(to_acu[101]));
	notech_mux2 i_10326010(.S(n_60623), .A(to_acu0[102]), .B(to_acu1[102]), 
		.Z(to_acu[102]));
	notech_mux2 i_10426011(.S(n_60623), .A(to_acu0[103]), .B(to_acu1[103]), 
		.Z(to_acu[103]));
	notech_mux2 i_10526012(.S(n_60623), .A(to_acu0[104]), .B(to_acu1[104]), 
		.Z(to_acu[104]));
	notech_mux2 i_10626013(.S(n_60623), .A(to_acu0[105]), .B(to_acu1[105]), 
		.Z(to_acu[105]));
	notech_mux2 i_10726014(.S(n_60623), .A(to_acu0[106]), .B(to_acu1[106]), 
		.Z(to_acu[106]));
	notech_mux2 i_10826015(.S(n_60623), .A(to_acu0[107]), .B(to_acu1[107]), 
		.Z(to_acu[107]));
	notech_mux2 i_10926016(.S(n_60623), .A(to_acu0[108]), .B(to_acu1[108]), 
		.Z(to_acu[108]));
	notech_mux2 i_11026017(.S(n_60623), .A(to_acu0[109]), .B(to_acu1[109]), 
		.Z(to_acu[109]));
	notech_mux2 i_11126018(.S(n_60623), .A(to_acu0[110]), .B(to_acu1[110]), 
		.Z(to_acu[110]));
	notech_mux2 i_11226019(.S(n_60623), .A(to_acu0[111]), .B(to_acu1[111]), 
		.Z(to_acu[111]));
	notech_mux2 i_11326020(.S(n_60623), .A(to_acu0[112]), .B(to_acu1[112]), 
		.Z(to_acu[112]));
	notech_mux2 i_11426021(.S(n_60623), .A(to_acu0[113]), .B(to_acu1[113]), 
		.Z(to_acu[113]));
	notech_mux2 i_11526022(.S(n_60623), .A(to_acu0[114]), .B(to_acu1[114]), 
		.Z(to_acu[114]));
	notech_mux2 i_11626023(.S(n_60618), .A(to_acu0[115]), .B(to_acu1[115]), 
		.Z(to_acu[115]));
	notech_mux2 i_11726024(.S(n_60618), .A(to_acu0[116]), .B(to_acu1[116]), 
		.Z(to_acu[116]));
	notech_mux2 i_11826025(.S(n_60618), .A(to_acu0[117]), .B(to_acu1[117]), 
		.Z(to_acu[117]));
	notech_mux2 i_11926026(.S(n_60618), .A(to_acu0[118]), .B(to_acu1[118]), 
		.Z(to_acu[118]));
	notech_mux2 i_12026027(.S(n_60618), .A(to_acu0[119]), .B(to_acu1[119]), 
		.Z(to_acu[119]));
	notech_mux2 i_12126028(.S(n_60618), .A(to_acu0[120]), .B(to_acu1[120]), 
		.Z(to_acu[120]));
	notech_mux2 i_12226029(.S(n_60618), .A(to_acu0[121]), .B(to_acu1[121]), 
		.Z(to_acu[121]));
	notech_mux2 i_12326030(.S(n_60623), .A(to_acu0[122]), .B(to_acu1[122]), 
		.Z(to_acu[122]));
	notech_mux2 i_12426031(.S(n_60623), .A(to_acu0[123]), .B(to_acu1[123]), 
		.Z(to_acu[123]));
	notech_mux2 i_12526032(.S(n_60623), .A(to_acu0[124]), .B(to_acu1[124]), 
		.Z(to_acu[124]));
	notech_mux2 i_12626033(.S(n_60618), .A(to_acu0[125]), .B(to_acu1[125]), 
		.Z(to_acu[125]));
	notech_mux2 i_12726034(.S(n_60618), .A(to_acu0[126]), .B(to_acu1[126]), 
		.Z(to_acu[126]));
	notech_mux2 i_12826035(.S(n_60618), .A(to_acu0[127]), .B(to_acu1[127]), 
		.Z(to_acu[127]));
	notech_mux2 i_12926036(.S(n_60623), .A(to_acu0[128]), .B(to_acu1[128]), 
		.Z(to_acu[128]));
	notech_mux2 i_13026037(.S(n_60624), .A(to_acu0[129]), .B(to_acu1[129]), 
		.Z(to_acu[129]));
	notech_mux2 i_13126038(.S(n_60624), .A(to_acu0[130]), .B(to_acu1[130]), 
		.Z(to_acu[130]));
	notech_mux2 i_13226039(.S(n_60629), .A(to_acu0[131]), .B(to_acu1[131]), 
		.Z(to_acu[131]));
	notech_mux2 i_13326040(.S(n_60624), .A(to_acu0[132]), .B(to_acu1[132]), 
		.Z(to_acu[132]));
	notech_mux2 i_13426041(.S(n_60624), .A(to_acu0[133]), .B(to_acu1[133]), 
		.Z(to_acu[133]));
	notech_mux2 i_13526042(.S(n_60624), .A(to_acu0[134]), .B(to_acu1[134]), 
		.Z(to_acu[134]));
	notech_mux2 i_13626043(.S(n_60629), .A(to_acu0[135]), .B(to_acu1[135]), 
		.Z(to_acu[135]));
	notech_mux2 i_13726044(.S(n_60629), .A(to_acu0[136]), .B(to_acu1[136]), 
		.Z(to_acu[136]));
	notech_mux2 i_13826045(.S(n_60629), .A(to_acu0[137]), .B(to_acu1[137]), 
		.Z(to_acu[137]));
	notech_mux2 i_13926046(.S(n_60629), .A(to_acu0[138]), .B(to_acu1[138]), 
		.Z(to_acu[138]));
	notech_mux2 i_14026047(.S(n_60629), .A(to_acu0[139]), .B(to_acu1[139]), 
		.Z(to_acu[139]));
	notech_mux2 i_14126048(.S(n_60629), .A(to_acu0[140]), .B(to_acu1[140]), 
		.Z(to_acu[140]));
	notech_mux2 i_14226049(.S(n_60629), .A(to_acu0[141]), .B(to_acu1[141]), 
		.Z(to_acu[141]));
	notech_mux2 i_14326050(.S(n_60624), .A(to_acu0[142]), .B(to_acu1[142]), 
		.Z(to_acu[142]));
	notech_mux2 i_14426051(.S(n_60624), .A(to_acu0[143]), .B(to_acu1[143]), 
		.Z(to_acu[143]));
	notech_mux2 i_14526052(.S(n_60624), .A(to_acu0[144]), .B(to_acu1[144]), 
		.Z(to_acu[144]));
	notech_mux2 i_14626053(.S(n_60624), .A(to_acu0[145]), .B(to_acu1[145]), 
		.Z(to_acu[145]));
	notech_mux2 i_14726054(.S(n_60624), .A(to_acu0[146]), .B(to_acu1[146]), 
		.Z(to_acu[146]));
	notech_mux2 i_14826055(.S(n_60624), .A(to_acu0[147]), .B(to_acu1[147]), 
		.Z(to_acu[147]));
	notech_mux2 i_14926056(.S(n_60624), .A(to_acu0[148]), .B(to_acu1[148]), 
		.Z(to_acu[148]));
	notech_mux2 i_15026057(.S(n_60624), .A(to_acu0[149]), .B(to_acu1[149]), 
		.Z(to_acu[149]));
	notech_mux2 i_15126058(.S(n_60624), .A(to_acu0[150]), .B(to_acu1[150]), 
		.Z(to_acu[150]));
	notech_mux2 i_15226059(.S(n_60624), .A(to_acu0[151]), .B(to_acu1[151]), 
		.Z(to_acu[151]));
	notech_mux2 i_15326060(.S(n_60624), .A(to_acu0[152]), .B(to_acu1[152]), 
		.Z(to_acu[152]));
	notech_mux2 i_15426061(.S(n_60624), .A(to_acu0[153]), .B(to_acu1[153]), 
		.Z(to_acu[153]));
	notech_mux2 i_15526062(.S(n_60624), .A(to_acu0[154]), .B(to_acu1[154]), 
		.Z(to_acu[154]));
	notech_mux2 i_15626063(.S(n_60658), .A(to_acu0[155]), .B(to_acu1[155]), 
		.Z(to_acu[155]));
	notech_mux2 i_15726064(.S(n_60658), .A(to_acu0[156]), .B(to_acu1[156]), 
		.Z(to_acu[156]));
	notech_mux2 i_15826065(.S(n_60658), .A(to_acu0[157]), .B(to_acu1[157]), 
		.Z(to_acu[157]));
	notech_mux2 i_15926066(.S(n_60658), .A(to_acu0[158]), .B(to_acu1[158]), 
		.Z(to_acu[158]));
	notech_mux2 i_16026067(.S(n_60658), .A(to_acu0[159]), .B(to_acu1[159]), 
		.Z(to_acu[159]));
	notech_mux2 i_16126068(.S(n_60658), .A(to_acu0[160]), .B(to_acu1[160]), 
		.Z(to_acu[160]));
	notech_mux2 i_16226069(.S(n_60658), .A(to_acu0[161]), .B(to_acu1[161]), 
		.Z(to_acu[161]));
	notech_mux2 i_16326070(.S(n_60658), .A(to_acu0[162]), .B(to_acu1[162]), 
		.Z(to_acu[162]));
	notech_mux2 i_16426071(.S(n_60658), .A(to_acu0[163]), .B(to_acu1[163]), 
		.Z(to_acu[163]));
	notech_mux2 i_16526072(.S(n_60658), .A(to_acu0[164]), .B(to_acu1[164]), 
		.Z(to_acu[164]));
	notech_mux2 i_16626073(.S(n_60658), .A(to_acu0[165]), .B(to_acu1[165]), 
		.Z(to_acu[165]));
	notech_mux2 i_16726074(.S(n_60658), .A(to_acu0[166]), .B(to_acu1[166]), 
		.Z(to_acu[166]));
	notech_mux2 i_16826075(.S(n_60658), .A(to_acu0[167]), .B(to_acu1[167]), 
		.Z(to_acu[167]));
	notech_mux2 i_16926076(.S(n_60657), .A(to_acu0[168]), .B(to_acu1[168]), 
		.Z(to_acu[168]));
	notech_mux2 i_17026077(.S(n_60657), .A(to_acu0[169]), .B(to_acu1[169]), 
		.Z(to_acu[169]));
	notech_mux2 i_17126078(.S(n_60657), .A(to_acu0[170]), .B(to_acu1[170]), 
		.Z(to_acu[170]));
	notech_mux2 i_17226079(.S(n_60657), .A(to_acu0[171]), .B(to_acu1[171]), 
		.Z(to_acu[171]));
	notech_mux2 i_17326080(.S(n_60657), .A(to_acu0[172]), .B(to_acu1[172]), 
		.Z(to_acu[172]));
	notech_mux2 i_17426081(.S(n_60657), .A(to_acu0[173]), .B(to_acu1[173]), 
		.Z(to_acu[173]));
	notech_mux2 i_17526082(.S(n_60657), .A(to_acu0[174]), .B(to_acu1[174]), 
		.Z(to_acu[174]));
	notech_mux2 i_17626083(.S(n_60658), .A(to_acu0[175]), .B(to_acu1[175]), 
		.Z(to_acu[175]));
	notech_mux2 i_17726084(.S(n_60658), .A(to_acu0[176]), .B(to_acu1[176]), 
		.Z(to_acu[176]));
	notech_mux2 i_17826085(.S(n_60658), .A(to_acu0[177]), .B(to_acu1[177]), 
		.Z(to_acu[177]));
	notech_mux2 i_17926086(.S(n_60657), .A(to_acu0[178]), .B(to_acu1[178]), 
		.Z(to_acu[178]));
	notech_mux2 i_18026087(.S(n_60657), .A(to_acu0[179]), .B(to_acu1[179]), 
		.Z(to_acu[179]));
	notech_mux2 i_18126088(.S(n_60657), .A(to_acu0[180]), .B(to_acu1[180]), 
		.Z(to_acu[180]));
	notech_mux2 i_18226089(.S(n_60658), .A(to_acu0[181]), .B(to_acu1[181]), 
		.Z(to_acu[181]));
	notech_mux2 i_18326090(.S(n_60668), .A(to_acu0[182]), .B(to_acu1[182]), 
		.Z(to_acu[182]));
	notech_mux2 i_18426091(.S(n_60668), .A(to_acu0[183]), .B(to_acu1[183]), 
		.Z(to_acu[183]));
	notech_mux2 i_18526092(.S(n_60668), .A(to_acu0[184]), .B(to_acu1[184]), 
		.Z(to_acu[184]));
	notech_mux2 i_18626093(.S(n_60668), .A(to_acu0[185]), .B(to_acu1[185]), 
		.Z(to_acu[185]));
	notech_mux2 i_18726094(.S(n_60668), .A(to_acu0[186]), .B(to_acu1[186]), 
		.Z(to_acu[186]));
	notech_mux2 i_18826095(.S(n_60668), .A(to_acu0[187]), .B(to_acu1[187]), 
		.Z(to_acu[187]));
	notech_mux2 i_18926096(.S(n_60668), .A(to_acu0[188]), .B(to_acu1[188]), 
		.Z(to_acu[188]));
	notech_mux2 i_19026097(.S(n_60668), .A(to_acu0[189]), .B(to_acu1[189]), 
		.Z(to_acu[189]));
	notech_mux2 i_19126098(.S(n_60668), .A(to_acu0[190]), .B(to_acu1[190]), 
		.Z(to_acu[190]));
	notech_mux2 i_19226099(.S(n_60668), .A(to_acu0[191]), .B(to_acu1[191]), 
		.Z(to_acu[191]));
	notech_mux2 i_19326100(.S(n_60668), .A(to_acu0[192]), .B(to_acu1[192]), 
		.Z(to_acu[192]));
	notech_mux2 i_19426101(.S(n_60668), .A(to_acu0[193]), .B(to_acu1[193]), 
		.Z(to_acu[193]));
	notech_mux2 i_19526102(.S(n_60668), .A(to_acu0[194]), .B(to_acu1[194]), 
		.Z(to_acu[194]));
	notech_mux2 i_19626103(.S(n_60663), .A(to_acu0[195]), .B(to_acu1[195]), 
		.Z(to_acu[195]));
	notech_mux2 i_19726104(.S(n_60663), .A(to_acu0[196]), .B(to_acu1[196]), 
		.Z(to_acu[196]));
	notech_mux2 i_19826105(.S(n_60663), .A(to_acu0[197]), .B(to_acu1[197]), 
		.Z(to_acu[197]));
	notech_mux2 i_19926106(.S(n_60658), .A(to_acu0[198]), .B(to_acu1[198]), 
		.Z(to_acu[198]));
	notech_mux2 i_20026107(.S(n_60663), .A(to_acu0[199]), .B(to_acu1[199]), 
		.Z(to_acu[199]));
	notech_mux2 i_20126108(.S(n_60663), .A(to_acu0[200]), .B(to_acu1[200]), 
		.Z(to_acu[200]));
	notech_mux2 i_20226109(.S(n_60663), .A(to_acu0[201]), .B(to_acu1[201]), 
		.Z(to_acu[201]));
	notech_mux2 i_20326110(.S(n_60663), .A(to_acu0[202]), .B(to_acu1[202]), 
		.Z(to_acu[202]));
	notech_mux2 i_20426111(.S(n_60663), .A(to_acu0[203]), .B(to_acu1[203]), 
		.Z(to_acu[203]));
	notech_mux2 i_20526112(.S(n_60663), .A(to_acu0[204]), .B(to_acu1[204]), 
		.Z(to_acu[204]));
	notech_mux2 i_20626113(.S(n_60663), .A(to_acu0[205]), .B(to_acu1[205]), 
		.Z(to_acu[205]));
	notech_mux2 i_20726114(.S(n_60663), .A(to_acu0[206]), .B(to_acu1[206]), 
		.Z(to_acu[206]));
	notech_mux2 i_20826115(.S(n_60663), .A(to_acu0[207]), .B(to_acu1[207]), 
		.Z(to_acu[207]));
	notech_mux2 i_20926116(.S(n_60657), .A(to_acu0[208]), .B(to_acu1[208]), 
		.Z(to_acu[208]));
	notech_mux2 i_21026117(.S(n_60646), .A(to_acu0[209]), .B(to_acu1[209]), 
		.Z(to_acu[209]));
	notech_mux2 i_21126118(.S(n_60646), .A(to_acu0[210]), .B(to_acu1[210]), 
		.Z(to_acu[210]));
	notech_mux2 i_627212(.S(n_60646), .A(\over_seg0[5] ), .B(\over_seg1[5] )
		, .Z(over_seg[5]));
	notech_mux2 i_127609(.S(n_60645), .A(\imm0[0] ), .B(\imm1[0] ), .Z(immediate
		[0]));
	notech_mux2 i_227610(.S(n_60645), .A(\imm0[1] ), .B(\imm1[1] ), .Z(immediate
		[1]));
	notech_mux2 i_327611(.S(n_60645), .A(\imm0[2] ), .B(\imm1[2] ), .Z(immediate
		[2]));
	notech_mux2 i_427612(.S(n_60646), .A(\imm0[3] ), .B(\imm1[3] ), .Z(immediate
		[3]));
	notech_mux2 i_527613(.S(n_60646), .A(\imm0[4] ), .B(\imm1[4] ), .Z(immediate
		[4]));
	notech_mux2 i_627614(.S(n_60646), .A(\imm0[5] ), .B(\imm1[5] ), .Z(immediate
		[5]));
	notech_mux2 i_727615(.S(n_60646), .A(\imm0[6] ), .B(\imm1[6] ), .Z(immediate
		[6]));
	notech_mux2 i_827616(.S(n_60646), .A(\imm0[7] ), .B(\imm1[7] ), .Z(immediate
		[7]));
	notech_mux2 i_927617(.S(n_60646), .A(\imm0[8] ), .B(\imm1[8] ), .Z(immediate
		[8]));
	notech_mux2 i_1027618(.S(n_60646), .A(\imm0[9] ), .B(\imm1[9] ), .Z(immediate
		[9]));
	notech_mux2 i_1127619(.S(n_60645), .A(\imm0[10] ), .B(\imm1[10] ), .Z(immediate
		[10]));
	notech_mux2 i_1227620(.S(n_60645), .A(\imm0[11] ), .B(\imm1[11] ), .Z(immediate
		[11]));
	notech_mux2 i_1327621(.S(n_60645), .A(\imm0[12] ), .B(\imm1[12] ), .Z(immediate
		[12]));
	notech_mux2 i_1427622(.S(n_60645), .A(\imm0[13] ), .B(\imm1[13] ), .Z(immediate
		[13]));
	notech_mux2 i_1527623(.S(n_60645), .A(\imm0[14] ), .B(\imm1[14] ), .Z(immediate
		[14]));
	notech_mux2 i_1627624(.S(n_60645), .A(\imm0[15] ), .B(\imm1[15] ), .Z(immediate
		[15]));
	notech_mux2 i_1727625(.S(n_60645), .A(\imm0[16] ), .B(\imm1[16] ), .Z(immediate
		[16]));
	notech_mux2 i_1827626(.S(n_60645), .A(\imm0[17] ), .B(\imm1[17] ), .Z(immediate
		[17]));
	notech_mux2 i_1927627(.S(n_60645), .A(\imm0[18] ), .B(\imm1[18] ), .Z(immediate
		[18]));
	notech_mux2 i_2027628(.S(n_60645), .A(\imm0[19] ), .B(\imm1[19] ), .Z(immediate
		[19]));
	notech_mux2 i_2127629(.S(n_60645), .A(\imm0[20] ), .B(\imm1[20] ), .Z(immediate
		[20]));
	notech_mux2 i_2227630(.S(n_60645), .A(\imm0[21] ), .B(\imm1[21] ), .Z(immediate
		[21]));
	notech_mux2 i_2327631(.S(n_60645), .A(\imm0[22] ), .B(\imm1[22] ), .Z(immediate
		[22]));
	notech_mux2 i_2427632(.S(n_60646), .A(\imm0[23] ), .B(\imm1[23] ), .Z(immediate
		[23]));
	notech_mux2 i_2527633(.S(n_60652), .A(\imm0[24] ), .B(\imm1[24] ), .Z(immediate
		[24]));
	notech_mux2 i_2627634(.S(n_60652), .A(\imm0[25] ), .B(\imm1[25] ), .Z(immediate
		[25]));
	notech_mux2 i_2727635(.S(n_60652), .A(\imm0[26] ), .B(\imm1[26] ), .Z(immediate
		[26]));
	notech_mux2 i_2827636(.S(n_60652), .A(\imm0[27] ), .B(\imm1[27] ), .Z(immediate
		[27]));
	notech_mux2 i_2927637(.S(n_60652), .A(\imm0[28] ), .B(\imm1[28] ), .Z(immediate
		[28]));
	notech_mux2 i_3027638(.S(n_60652), .A(\imm0[29] ), .B(\imm1[29] ), .Z(immediate
		[29]));
	notech_mux2 i_3127639(.S(n_60657), .A(\imm0[30] ), .B(\imm1[30] ), .Z(immediate
		[30]));
	notech_mux2 i_3227640(.S(n_60657), .A(\imm0[31] ), .B(\imm1[31] ), .Z(immediate
		[31]));
	notech_mux2 i_3327641(.S(n_60657), .A(\imm0[32] ), .B(\imm1[32] ), .Z(immediate
		[32]));
	notech_mux2 i_3427642(.S(n_60657), .A(\imm0[33] ), .B(\imm1[33] ), .Z(immediate
		[33]));
	notech_mux2 i_3527643(.S(n_60657), .A(\imm0[34] ), .B(\imm1[34] ), .Z(immediate
		[34]));
	notech_mux2 i_3627644(.S(n_60657), .A(\imm0[35] ), .B(\imm1[35] ), .Z(immediate
		[35]));
	notech_mux2 i_3727645(.S(n_60657), .A(\imm0[36] ), .B(\imm1[36] ), .Z(immediate
		[36]));
	notech_mux2 i_3827646(.S(n_60646), .A(\imm0[37] ), .B(\imm1[37] ), .Z(immediate
		[37]));
	notech_mux2 i_3927647(.S(n_60646), .A(\imm0[38] ), .B(\imm1[38] ), .Z(immediate
		[38]));
	notech_mux2 i_4027648(.S(n_60646), .A(\imm0[39] ), .B(\imm1[39] ), .Z(immediate
		[39]));
	notech_mux2 i_4127649(.S(n_60646), .A(\imm0[40] ), .B(\imm1[40] ), .Z(immediate
		[40]));
	notech_mux2 i_4227650(.S(n_60646), .A(\imm0[41] ), .B(\imm1[41] ), .Z(immediate
		[41]));
	notech_mux2 i_4327651(.S(n_60646), .A(\imm0[42] ), .B(\imm1[42] ), .Z(immediate
		[42]));
	notech_mux2 i_4427652(.S(n_60646), .A(\imm0[43] ), .B(\imm1[43] ), .Z(immediate
		[43]));
	notech_mux2 i_4527653(.S(n_60652), .A(\imm0[44] ), .B(\imm1[44] ), .Z(immediate
		[44]));
	notech_mux2 i_4627654(.S(n_60652), .A(\imm0[45] ), .B(\imm1[45] ), .Z(immediate
		[45]));
	notech_mux2 i_4727655(.S(n_60652), .A(\imm0[46] ), .B(\imm1[46] ), .Z(immediate
		[46]));
	notech_mux2 i_4827656(.S(n_60652), .A(\imm0[47] ), .B(\imm1[47] ), .Z(immediate
		[47]));
	notech_or2 i_481(.A(n_2833), .B(pc_req), .Z(n_2872));
	notech_nand3 i_16075011(.A(n_3247), .B(n_59695), .C(n_22091849), .Z(\nbus_13538[0] 
		));
	notech_nand3 i_16175010(.A(n_3247), .B(n_59695), .C(n_21991848), .Z(\nbus_13549[0] 
		));
	notech_nand3 i_17175009(.A(n_59695), .B(n_21891847), .C(n_3247), .Z(\nbus_13539[0] 
		));
	notech_nao3 i_22175008(.A(n_18050174), .B(n_1568), .C(n_21791846), .Z(n_43061
		));
	notech_and2 i_430195(.A(cpl[0]), .B(cpl[1]), .Z(n_161751607));
	notech_ao4 i_6926187(.A(n_57484), .B(n_39225), .C(n_58672), .D(n_40186),
		 .Z(n_48806));
	notech_ao4 i_2026138(.A(n_57484), .B(n_39152), .C(n_58672), .D(n_40187),
		 .Z(n_48512));
	notech_ao4 i_2727827(.A(n_57484), .B(n_38558), .C(n_240991256), .D(n_58672
		), .Z(n_46767));
	notech_nand3 i_12825779(.A(n_59695), .B(n_3246), .C(n_130892929), .Z(n_46011
		));
	notech_nand3 i_12725778(.A(n_59695), .B(n_21391842), .C(n_131092931), .Z
		(n_46005));
	notech_nand3 i_12625777(.A(n_59695), .B(n_3246), .C(n_131192932), .Z(n_45999
		));
	notech_nand3 i_12525776(.A(n_59695), .B(n_21391842), .C(n_131292933), .Z
		(n_45993));
	notech_nand3 i_12425775(.A(n_59695), .B(n_21391842), .C(n_131392934), .Z
		(n_45987));
	notech_nand3 i_12325774(.A(n_59695), .B(n_21291841), .C(n_131592936), .Z
		(n_45981));
	notech_nand2 i_12225773(.A(n_59695), .B(n_131692937), .Z(n_45975));
	notech_nand3 i_12125772(.A(n_59695), .B(n_21391842), .C(n_131792938), .Z
		(n_45969));
	notech_nand3 i_12025771(.A(n_59695), .B(n_3246), .C(n_131892939), .Z(n_45963
		));
	notech_nand3 i_11925770(.A(n_59695), .B(n_3246), .C(n_131992940), .Z(n_45957
		));
	notech_nand3 i_11825769(.A(n_59695), .B(n_3246), .C(n_132092941), .Z(n_45951
		));
	notech_nand3 i_11725768(.A(n_59695), .B(n_21291841), .C(n_132192942), .Z
		(n_45945));
	notech_nand3 i_11325764(.A(n_59695), .B(n_2056), .C(n_132392944), .Z(n_45921
		));
	notech_nand2 i_11225763(.A(n_59693), .B(n_132592946), .Z(n_45915));
	notech_nand3 i_11125762(.A(n_59693), .B(n_3246), .C(n_132692947), .Z(n_45909
		));
	notech_nand2 i_11025761(.A(n_59693), .B(n_132792948), .Z(n_45903));
	notech_nand2 i_10925760(.A(n_59693), .B(n_132892949), .Z(n_45897));
	notech_nand3 i_10825759(.A(n_132992950), .B(n_16150155), .C(n_21191840),
		 .Z(n_45891));
	notech_nand3 i_10725758(.A(n_59693), .B(n_133092951), .C(n_126492885), .Z
		(n_45885));
	notech_nand2 i_10625757(.A(n_59693), .B(n_133292953), .Z(n_45879));
	notech_nand3 i_10525756(.A(n_59693), .B(n_21291841), .C(n_133392954), .Z
		(n_45873));
	notech_nand3 i_10425755(.A(n_59693), .B(n_21291841), .C(n_133492955), .Z
		(n_45867));
	notech_nand3 i_10325754(.A(n_59693), .B(n_21291841), .C(n_133592956), .Z
		(n_45861));
	notech_nand3 i_10225753(.A(n_59693), .B(n_21291841), .C(n_133692957), .Z
		(n_45855));
	notech_nand2 i_10125752(.A(n_59695), .B(n_133792958), .Z(n_45849));
	notech_nand3 i_9925750(.A(n_59693), .B(n_133892959), .C(n_1418), .Z(n_45837
		));
	notech_nand2 i_9625747(.A(n_59693), .B(n_133992960), .Z(n_45819));
	notech_nand2 i_9225743(.A(n_59693), .B(n_134092961), .Z(n_45795));
	notech_nand2 i_9125742(.A(n_59693), .B(n_134192962), .Z(n_45789));
	notech_nand2 i_9025741(.A(n_59693), .B(n_134292963), .Z(n_45783));
	notech_nand2 i_8925740(.A(n_59681), .B(n_134392964), .Z(n_45777));
	notech_nand3 i_8725738(.A(n_59681), .B(n_134492965), .C(n_123792858), .Z
		(n_45765));
	notech_or4 i_8225733(.A(pg_fault), .B(pc_req), .C(n_123492855), .D(n_38327
		), .Z(n_45735));
	notech_nand3 i_8125732(.A(n_59681), .B(n_134892969), .C(n_123192852), .Z
		(n_45729));
	notech_nand3 i_8025731(.A(n_59681), .B(n_21291841), .C(n_135092971), .Z(n_45723
		));
	notech_nand3 i_7925730(.A(n_59681), .B(n_21291841), .C(n_135192972), .Z(n_45717
		));
	notech_nand3 i_7825729(.A(n_59681), .B(n_21291841), .C(n_135292973), .Z(n_45711
		));
	notech_nand3 i_7725728(.A(n_59681), .B(n_21291841), .C(n_135392974), .Z(n_45705
		));
	notech_nand3 i_7625727(.A(n_59681), .B(n_21291841), .C(n_135492975), .Z(n_45699
		));
	notech_nand3 i_7525726(.A(n_59683), .B(n_21291841), .C(n_135592976), .Z(n_45693
		));
	notech_nand2 i_7425725(.A(n_59683), .B(n_135692977), .Z(n_45687));
	notech_nand3 i_7225723(.A(n_59683), .B(n_21391842), .C(n_135792978), .Z(n_45675
		));
	notech_nand3 i_7125722(.A(n_59683), .B(n_3246), .C(n_135892979), .Z(n_45669
		));
	notech_nand3 i_7025721(.A(n_59683), .B(n_3246), .C(n_135992980), .Z(n_45663
		));
	notech_nand3 i_6925720(.A(n_59681), .B(n_21391842), .C(n_136092981), .Z(n_45657
		));
	notech_nand3 i_6825719(.A(n_59683), .B(n_21391842), .C(n_136192982), .Z(n_45651
		));
	notech_nand3 i_6725718(.A(n_59683), .B(n_58425), .C(n_136292983), .Z(n_45645
		));
	notech_nand2 i_6625717(.A(n_59681), .B(n_136392984), .Z(n_45639));
	notech_nand3 i_6525716(.A(n_59680), .B(n_21291841), .C(n_136492985), .Z(n_45633
		));
	notech_nand2 i_6425715(.A(n_59680), .B(n_136592986), .Z(n_45627));
	notech_nand3 i_6325714(.A(n_59680), .B(n_58425), .C(n_136692987), .Z(n_45621
		));
	notech_nand3 i_6225713(.A(n_59680), .B(n_58425), .C(n_136792988), .Z(n_45615
		));
	notech_nand2 i_6125712(.A(n_59680), .B(n_136892989), .Z(n_45609));
	notech_nand2 i_6025711(.A(n_59680), .B(n_136992990), .Z(n_45603));
	notech_nand3 i_5925710(.A(n_59680), .B(n_58425), .C(n_137092991), .Z(n_45597
		));
	notech_nand3 i_5725708(.A(n_59680), .B(n_21391842), .C(n_137192992), .Z(n_45585
		));
	notech_nand3 i_5625707(.A(n_59681), .B(n_58416), .C(n_137292993), .Z(n_45579
		));
	notech_nand3 i_5425705(.A(n_59681), .B(n_21391842), .C(n_137392994), .Z(n_45567
		));
	notech_nand2 i_5325704(.A(n_59681), .B(n_137492995), .Z(n_45561));
	notech_nand2 i_5225703(.A(n_59681), .B(n_137592996), .Z(n_45555));
	notech_nand3 i_5125702(.A(n_59681), .B(n_58425), .C(n_137692997), .Z(n_45549
		));
	notech_nand2 i_5025701(.A(n_59681), .B(n_137792998), .Z(n_45543));
	notech_nand2 i_4925700(.A(n_59681), .B(n_137892999), .Z(n_45537));
	notech_nand3 i_4825699(.A(n_59681), .B(n_21391842), .C(n_137993000), .Z(n_45531
		));
	notech_nand3 i_4725698(.A(n_59683), .B(n_58425), .C(n_138093001), .Z(n_45525
		));
	notech_nand3 i_4625697(.A(n_59686), .B(n_58416), .C(n_138193002), .Z(n_45519
		));
	notech_nand2 i_4525696(.A(n_59686), .B(n_138293003), .Z(n_45513));
	notech_nand3 i_4425695(.A(n_59686), .B(n_58416), .C(n_138393004), .Z(n_45507
		));
	notech_nand3 i_4325694(.A(n_59686), .B(n_138493005), .C(n_21391842), .Z(n_45501
		));
	notech_nand2 i_4225693(.A(n_59686), .B(n_138593006), .Z(n_45495));
	notech_nand2 i_4125692(.A(n_59686), .B(n_138693007), .Z(n_45489));
	notech_nand2 i_4025691(.A(n_59686), .B(n_138793008), .Z(n_45483));
	notech_nand3 i_3925690(.A(n_59686), .B(n_58416), .C(n_138893009), .Z(n_45477
		));
	notech_nand3 i_3825689(.A(n_59688), .B(n_58416), .C(n_138993010), .Z(n_45471
		));
	notech_nand2 i_3725688(.A(n_59688), .B(n_139093011), .Z(n_45465));
	notech_nand2 i_3625687(.A(n_59688), .B(n_139193012), .Z(n_45459));
	notech_nand3 i_3525686(.A(n_59688), .B(n_58416), .C(n_139293013), .Z(n_45453
		));
	notech_nand3 i_3425685(.A(n_59686), .B(n_58416), .C(n_139393014), .Z(n_45447
		));
	notech_nand3 i_3325684(.A(n_59686), .B(n_58416), .C(n_139493015), .Z(n_45441
		));
	notech_nand2 i_3225683(.A(n_59688), .B(n_139593016), .Z(n_45435));
	notech_nand3 i_3125682(.A(n_59686), .B(n_58416), .C(n_139693017), .Z(n_45429
		));
	notech_nand3 i_3025681(.A(n_59686), .B(n_58416), .C(n_139793018), .Z(n_45423
		));
	notech_nand2 i_2925680(.A(n_59683), .B(n_139893019), .Z(n_45417));
	notech_nand2 i_2825679(.A(n_59683), .B(n_139993020), .Z(n_45411));
	notech_nand3 i_2725678(.A(n_59683), .B(n_58416), .C(n_140093021), .Z(n_45405
		));
	notech_nand3 i_2625677(.A(n_59683), .B(n_140193022), .C(n_58416), .Z(n_45399
		));
	notech_nand2 i_1025661(.A(n_59683), .B(n_140293023), .Z(n_45303));
	notech_nand3 i_825659(.A(n_59683), .B(n_58425), .C(n_140393024), .Z(n_45291
		));
	notech_nand3 i_725658(.A(n_59683), .B(n_3246), .C(n_140493025), .Z(n_45285
		));
	notech_nand3 i_425655(.A(n_59683), .B(n_58425), .C(n_140593026), .Z(n_45267
		));
	notech_nand3 i_325654(.A(n_59686), .B(n_58425), .C(n_140693027), .Z(n_45261
		));
	notech_nand3 i_225653(.A(n_59686), .B(n_140793028), .C(n_58425), .Z(n_45255
		));
	notech_nand2 i_125652(.A(n_140893029), .B(n_59686), .Z(n_45249));
	notech_ao4 i_223150(.A(n_58672), .B(n_40105), .C(n_57484), .D(n_39825), 
		.Z(n_42944));
	notech_ao4 i_123149(.A(n_58672), .B(n_40104), .C(n_57484), .D(n_39824), 
		.Z(n_42938));
	notech_and4 i_521(.A(n_59686), .B(n_2798), .C(n_2126), .D(n_2127), .Z(n_2869
		));
	notech_nao3 i_172(.A(n_1740), .B(n_2121), .C(n_2122), .Z(n_2867));
	notech_ao3 i_17(.A(n_1740), .B(n_2121), .C(n_2122), .Z(n_2864));
	notech_and2 i_498(.A(n_40174), .B(in128[9]), .Z(n_2856));
	notech_or2 i_484(.A(valid_len[2]), .B(valid_len[5]), .Z(n_2851));
	notech_ao3 i_3885(.A(n_40193), .B(n_59596), .C(n_2849), .Z(n_2850));
	notech_or4 i_6323(.A(fsm[2]), .B(fsm[0]), .C(n_2825), .D(fsm[1]), .Z(n_2849
		));
	notech_and2 i_5(.A(n_40193), .B(n_59596), .Z(n_2847));
	notech_or2 i_24(.A(ipg_fault), .B(n_2844), .Z(n_2845));
	notech_and2 i_6324(.A(n_60652), .B(n_38421), .Z(n_2844));
	notech_xor2 i_6335(.A(n_2835), .B(n_2840), .Z(n_2841));
	notech_xor2 i_215(.A(imm_sz[1]), .B(i_ptr[1]), .Z(n_2840));
	notech_xor2 i_15(.A(imm_sz[2]), .B(i_ptr[2]), .Z(n_2839));
	notech_nand2 i_6331(.A(i_ptr[3]), .B(n_39851), .Z(n_2838));
	notech_ao4 i_6332(.A(n_2097), .B(n_39852), .C(n_39860), .D(n_38653), .Z(n_2837
		));
	notech_ao4 i_2130159(.A(n_2835), .B(n_2094), .C(imm_sz[1]), .D(i_ptr[1])
		, .Z(n_2836));
	notech_nand2 i_75075(.A(n_162893249), .B(n_5392), .Z(\nbus_13566[0] ));
	notech_nand2 i_18973383(.A(n_162893249), .B(n_162793248), .Z(\nbus_13535[0] 
		));
	notech_mux2 i_828080(.S(n_162893249), .A(ififo_rvect4[7]), .B(ififo_rvect2
		[7]), .Z(n_46552));
	notech_mux2 i_728079(.S(n_162893249), .A(ififo_rvect4[6]), .B(ififo_rvect2
		[6]), .Z(n_46546));
	notech_mux2 i_628078(.S(n_162893249), .A(ififo_rvect4[5]), .B(ififo_rvect2
		[5]), .Z(n_46540));
	notech_mux2 i_528077(.S(n_162893249), .A(ififo_rvect4[4]), .B(ififo_rvect2
		[4]), .Z(n_46534));
	notech_mux2 i_428076(.S(n_162893249), .A(ififo_rvect4[3]), .B(ififo_rvect2
		[3]), .Z(n_46528));
	notech_mux2 i_328075(.S(n_162893249), .A(ififo_rvect4[2]), .B(ififo_rvect2
		[2]), .Z(n_46522));
	notech_mux2 i_228074(.S(n_162893249), .A(ififo_rvect4[1]), .B(ififo_rvect2
		[1]), .Z(n_46516));
	notech_mux2 i_128073(.S(n_55060), .A(ififo_rvect4[0]), .B(ififo_rvect2[0
		]), .Z(n_46510));
	notech_mux2 i_828040(.S(n_55060), .A(ififo_rvect3[7]), .B(ififo_rvect1[7
		]), .Z(n_41646));
	notech_mux2 i_728039(.S(n_55060), .A(ififo_rvect3[6]), .B(ififo_rvect1[6
		]), .Z(n_41640));
	notech_mux2 i_628038(.S(n_55060), .A(ififo_rvect3[5]), .B(ififo_rvect1[5
		]), .Z(n_41634));
	notech_mux2 i_528037(.S(n_55060), .A(ififo_rvect3[4]), .B(ififo_rvect1[4
		]), .Z(n_41628));
	notech_mux2 i_428036(.S(n_55060), .A(ififo_rvect3[3]), .B(ififo_rvect1[3
		]), .Z(n_41622));
	notech_mux2 i_328035(.S(n_55060), .A(ififo_rvect3[2]), .B(ififo_rvect1[2
		]), .Z(n_41616));
	notech_mux2 i_228034(.S(n_55060), .A(ififo_rvect3[1]), .B(ififo_rvect1[1
		]), .Z(n_41610));
	notech_mux2 i_128033(.S(n_55060), .A(ififo_rvect3[0]), .B(ififo_rvect1[0
		]), .Z(n_41604));
	notech_mux2 i_828048(.S(n_55060), .A(ififo_rvect2[7]), .B(ivect[7]), .Z(n_41864
		));
	notech_mux2 i_728047(.S(n_55060), .A(ififo_rvect2[6]), .B(ivect[6]), .Z(n_41858
		));
	notech_mux2 i_628046(.S(n_162893249), .A(ififo_rvect2[5]), .B(ivect[5]),
		 .Z(n_41852));
	notech_mux2 i_528045(.S(n_55060), .A(ififo_rvect2[4]), .B(ivect[4]), .Z(n_41846
		));
	notech_mux2 i_428044(.S(n_55060), .A(ififo_rvect2[3]), .B(ivect[3]), .Z(n_41840
		));
	notech_mux2 i_328043(.S(n_55060), .A(ififo_rvect2[2]), .B(ivect[2]), .Z(n_41834
		));
	notech_mux2 i_228042(.S(n_55060), .A(ififo_rvect2[1]), .B(ivect[1]), .Z(n_41828
		));
	notech_mux2 i_128041(.S(n_55060), .A(ififo_rvect2[0]), .B(ivect[0]), .Z(n_41822
		));
	notech_nand3 i_323229(.A(n_160993230), .B(n_160893229), .C(n_849150), .Z
		(n_41752));
	notech_ao4 i_10425499(.A(n_58672), .B(n_39965), .C(n_57484), .D(n_38835)
		, .Z(n_50550));
	notech_ao4 i_21126329(.A(n_58673), .B(n_40102), .C(n_57473), .D(n_39421)
		, .Z(n_49658));
	notech_ao4 i_21026328(.A(n_58673), .B(n_40101), .C(n_57462), .D(n_39420)
		, .Z(n_49652));
	notech_ao4 i_20926327(.A(n_58673), .B(n_40100), .C(n_57462), .D(n_39418)
		, .Z(n_49646));
	notech_ao4 i_20726325(.A(n_58673), .B(n_40098), .C(n_57462), .D(n_39415)
		, .Z(n_49634));
	notech_ao4 i_20626324(.A(n_58673), .B(n_40097), .C(n_57463), .D(n_39414)
		, .Z(n_49628));
	notech_ao4 i_20526323(.A(n_58673), .B(n_40096), .C(n_57462), .D(n_39412)
		, .Z(n_49622));
	notech_ao4 i_20226320(.A(n_58673), .B(n_40093), .C(n_57462), .D(n_39408)
		, .Z(n_49604));
	notech_ao4 i_19726315(.A(n_58673), .B(n_40088), .C(n_57462), .D(n_39400)
		, .Z(n_49574));
	notech_ao4 i_19626314(.A(n_58673), .B(n_40087), .C(n_57462), .D(n_39399)
		, .Z(n_49568));
	notech_ao4 i_19526313(.A(n_58673), .B(n_40086), .C(n_57462), .D(n_39397)
		, .Z(n_49562));
	notech_ao4 i_19426312(.A(n_58672), .B(n_40085), .C(n_57462), .D(n_39396)
		, .Z(n_49556));
	notech_ao4 i_19326311(.A(n_58667), .B(n_40084), .C(n_57463), .D(n_39394)
		, .Z(n_49550));
	notech_ao4 i_19226310(.A(n_58667), .B(n_40083), .C(n_57463), .D(n_39393)
		, .Z(n_49544));
	notech_ao4 i_19126309(.A(n_58667), .B(n_40082), .C(n_57463), .D(n_39391)
		, .Z(n_49538));
	notech_ao4 i_19026308(.A(n_58667), .B(n_40081), .C(n_57463), .D(n_39390)
		, .Z(n_49532));
	notech_ao4 i_18926307(.A(n_58667), .B(n_40080), .C(n_57463), .D(n_39388)
		, .Z(n_49526));
	notech_ao4 i_18826306(.A(n_58667), .B(n_40079), .C(n_57463), .D(n_39387)
		, .Z(n_49520));
	notech_ao4 i_18726305(.A(n_58667), .B(n_40078), .C(n_57463), .D(n_39385)
		, .Z(n_49514));
	notech_ao4 i_18626304(.A(n_58667), .B(n_40077), .C(n_57463), .D(n_39384)
		, .Z(n_49508));
	notech_ao4 i_18526303(.A(n_58667), .B(n_40076), .C(n_57463), .D(n_39382)
		, .Z(n_49502));
	notech_ao4 i_18426302(.A(n_58667), .B(n_40075), .C(n_57463), .D(n_39381)
		, .Z(n_49496));
	notech_ao4 i_18326301(.A(n_58672), .B(n_40074), .C(n_57462), .D(n_39379)
		, .Z(n_49490));
	notech_ao4 i_18226300(.A(n_58672), .B(n_40073), .C(n_57457), .D(n_39378)
		, .Z(n_49484));
	notech_ao4 i_18126299(.A(n_58672), .B(n_40072), .C(n_57457), .D(n_39376)
		, .Z(n_49478));
	notech_ao4 i_18026298(.A(n_58672), .B(n_40071), .C(n_57457), .D(n_39375)
		, .Z(n_49472));
	notech_ao4 i_17826296(.A(n_58672), .B(n_40069), .C(n_57457), .D(n_39372)
		, .Z(n_49460));
	notech_ao4 i_17726295(.A(n_58667), .B(n_40068), .C(n_57457), .D(n_39370)
		, .Z(n_49454));
	notech_ao4 i_17526293(.A(n_58667), .B(n_40066), .C(n_57457), .D(n_39367)
		, .Z(n_49442));
	notech_ao4 i_17226290(.A(n_58672), .B(n_40063), .C(n_57457), .D(n_39363)
		, .Z(n_49424));
	notech_ao4 i_17126289(.A(n_58672), .B(n_40062), .C(n_57457), .D(n_39361)
		, .Z(n_49418));
	notech_ao4 i_16326281(.A(n_58672), .B(n_40054), .C(n_57457), .D(n_39352)
		, .Z(n_49370));
	notech_ao4 i_16226280(.A(n_58673), .B(n_40053), .C(n_57457), .D(n_39351)
		, .Z(n_49364));
	notech_ao4 i_16126279(.A(n_58680), .B(n_40052), .C(n_57462), .D(n_39350)
		, .Z(n_49358));
	notech_ao4 i_16026278(.A(n_58680), .B(n_40051), .C(n_57462), .D(n_39349)
		, .Z(n_49352));
	notech_ao4 i_15926277(.A(n_58680), .B(n_40050), .C(n_57462), .D(n_39348)
		, .Z(n_49346));
	notech_ao4 i_15826276(.A(n_58680), .B(n_40049), .C(n_57462), .D(n_39347)
		, .Z(n_49340));
	notech_ao4 i_15726275(.A(n_58680), .B(n_40048), .C(n_57462), .D(n_39346)
		, .Z(n_49334));
	notech_ao4 i_15626274(.A(n_58680), .B(n_40047), .C(n_57457), .D(n_39345)
		, .Z(n_49328));
	notech_ao4 i_15526273(.A(n_58680), .B(n_40046), .C(n_57457), .D(n_39344)
		, .Z(n_49322));
	notech_ao4 i_15426272(.A(n_58680), .B(n_40045), .C(n_57462), .D(n_39343)
		, .Z(n_49316));
	notech_ao4 i_15326271(.A(n_58680), .B(n_40044), .C(n_57462), .D(n_39342)
		, .Z(n_49310));
	notech_ao4 i_15226270(.A(n_58680), .B(n_40043), .C(n_57462), .D(n_39341)
		, .Z(n_49304));
	notech_ao4 i_15126269(.A(n_58683), .B(n_40042), .C(n_57469), .D(n_39340)
		, .Z(n_49298));
	notech_ao4 i_15026268(.A(n_58683), .B(n_40041), .C(n_57469), .D(n_39339)
		, .Z(n_49292));
	notech_ao4 i_14926267(.A(n_58683), .B(n_40040), .C(n_57469), .D(n_39338)
		, .Z(n_49286));
	notech_ao4 i_14826266(.A(n_58683), .B(n_40039), .C(n_57469), .D(n_39337)
		, .Z(n_49280));
	notech_ao4 i_14626264(.A(n_58683), .B(n_40037), .C(n_57469), .D(n_39335)
		, .Z(n_49268));
	notech_ao4 i_14526263(.A(n_58680), .B(n_40036), .C(n_57469), .D(n_39334)
		, .Z(n_49262));
	notech_ao4 i_14426262(.A(n_58680), .B(n_40035), .C(n_57469), .D(n_39333)
		, .Z(n_49256));
	notech_ao4 i_14326261(.A(n_58680), .B(n_40034), .C(n_57469), .D(n_39332)
		, .Z(n_49250));
	notech_ao4 i_14226260(.A(n_58683), .B(n_40033), .C(n_57469), .D(n_39331)
		, .Z(n_49244));
	notech_ao4 i_14126259(.A(n_58683), .B(n_40032), .C(n_57469), .D(n_39330)
		, .Z(n_49238));
	notech_ao4 i_14026258(.A(n_58680), .B(n_40031), .C(n_57473), .D(n_39329)
		, .Z(n_49232));
	notech_ao4 i_13826256(.A(n_58678), .B(n_40029), .C(n_57473), .D(n_39327)
		, .Z(n_49220));
	notech_ao4 i_13726255(.A(n_58673), .B(n_40028), .C(n_57473), .D(n_39326)
		, .Z(n_49214));
	notech_ao4 i_13626254(.A(n_58678), .B(n_40027), .C(n_57473), .D(n_39324)
		, .Z(n_49208));
	notech_ao4 i_13526253(.A(n_58678), .B(n_40026), .C(n_57473), .D(n_39323)
		, .Z(n_49202));
	notech_ao4 i_13426252(.A(n_58678), .B(n_40025), .C(n_57469), .D(n_39321)
		, .Z(n_49196));
	notech_ao4 i_13326251(.A(n_58673), .B(n_40024), .C(n_57469), .D(n_39320)
		, .Z(n_49190));
	notech_ao4 i_13226250(.A(n_58673), .B(n_40023), .C(n_57473), .D(n_39318)
		, .Z(n_49184));
	notech_ao4 i_13126249(.A(n_58673), .B(n_40022), .C(n_57473), .D(n_39317)
		, .Z(n_49178));
	notech_ao4 i_13026248(.A(n_57473), .B(n_39315), .C(n_58673), .D(n_40021)
		, .Z(n_49172));
	notech_ao4 i_12926247(.A(n_58673), .B(n_40020), .C(n_57469), .D(n_39314)
		, .Z(n_49166));
	notech_ao4 i_12326241(.A(n_57463), .B(n_39306), .C(n_58678), .D(n_40014)
		, .Z(n_49130));
	notech_ao4 i_12226240(.A(n_57463), .B(n_39305), .C(n_58678), .D(n_40013)
		, .Z(n_49124));
	notech_ao4 i_12126239(.A(n_57475), .B(n_39304), .C(n_58678), .D(n_40012)
		, .Z(n_49118));
	notech_ao4 i_12026238(.A(n_58678), .B(n_40011), .C(n_57475), .D(n_39302)
		, .Z(n_49112));
	notech_ao4 i_11926237(.A(n_57475), .B(n_39301), .C(n_58678), .D(n_40010)
		, .Z(n_49106));
	notech_ao4 i_11826236(.A(n_58678), .B(n_40009), .C(n_57463), .D(n_39299)
		, .Z(n_49100));
	notech_ao4 i_11726235(.A(n_57463), .B(n_39298), .C(n_58678), .D(n_40008)
		, .Z(n_49094));
	notech_ao4 i_11626234(.A(n_57463), .B(n_39296), .C(n_58678), .D(n_40007)
		, .Z(n_49088));
	notech_ao4 i_11526233(.A(n_57463), .B(n_39295), .C(n_58678), .D(n_40006)
		, .Z(n_49082));
	notech_ao4 i_11426232(.A(n_57463), .B(n_39293), .C(n_58678), .D(n_40005)
		, .Z(n_49076));
	notech_ao4 i_11226230(.A(n_57469), .B(n_39290), .C(n_58723), .D(n_40003)
		, .Z(n_49064));
	notech_ao4 i_11126229(.A(n_57469), .B(n_39289), .C(n_58723), .D(n_40002)
		, .Z(n_49058));
	notech_ao4 i_11026228(.A(n_57469), .B(n_39287), .C(n_58723), .D(n_40001)
		, .Z(n_49052));
	notech_ao4 i_10926227(.A(n_57469), .B(n_39286), .C(n_58723), .D(n_40000)
		, .Z(n_49046));
	notech_ao4 i_10826226(.A(n_57469), .B(n_39284), .C(n_58723), .D(n_39999)
		, .Z(n_49040));
	notech_ao4 i_10626224(.A(n_57475), .B(n_39281), .C(n_58719), .D(n_39997)
		, .Z(n_49028));
	notech_ao4 i_10526223(.A(n_57475), .B(n_39280), .C(n_58719), .D(n_39996)
		, .Z(n_49022));
	notech_ao4 i_10426222(.A(n_57475), .B(n_39278), .C(n_58723), .D(n_39995)
		, .Z(n_49016));
	notech_ao4 i_10326221(.A(n_57469), .B(n_39277), .C(n_58723), .D(n_39994)
		, .Z(n_49010));
	notech_ao4 i_10226220(.A(n_57469), .B(n_39275), .C(n_58723), .D(n_39993)
		, .Z(n_49004));
	notech_ao4 i_9026208(.A(n_57490), .B(n_39257), .C(n_58725), .D(n_40201),
		 .Z(n_48932));
	notech_ao4 i_8926207(.A(n_57513), .B(n_39256), .C(n_58723), .D(n_40200),
		 .Z(n_48926));
	notech_ao4 i_8826206(.A(n_57513), .B(n_39254), .C(n_58725), .D(n_40199),
		 .Z(n_48920));
	notech_ao4 i_8426202(.A(n_57513), .B(n_39247), .C(n_58725), .D(n_40213),
		 .Z(n_48896));
	notech_ao4 i_8326201(.A(n_57513), .B(n_39246), .C(n_58725), .D(n_40177),
		 .Z(n_48890));
	notech_ao4 i_6426182(.A(n_58723), .B(n_40111), .C(n_57513), .D(n_39217),
		 .Z(n_48776));
	notech_ao4 i_6326181(.A(n_58723), .B(n_40165), .C(n_57513), .D(n_39216),
		 .Z(n_48770));
	notech_ao4 i_6226180(.A(n_58723), .B(n_40145), .C(n_57513), .D(n_39214),
		 .Z(n_48764));
	notech_ao4 i_6126179(.A(n_58723), .B(n_40112), .C(n_57513), .D(n_39213),
		 .Z(n_48758));
	notech_ao4 i_6026178(.A(n_58723), .B(n_40129), .C(n_57513), .D(n_39211),
		 .Z(n_48752));
	notech_ao4 i_5926177(.A(n_58719), .B(n_40122), .C(n_57513), .D(n_39210),
		 .Z(n_48746));
	notech_ao4 i_5826176(.A(n_58717), .B(n_40123), .C(n_57515), .D(n_39208),
		 .Z(n_48740));
	notech_ao4 i_5726175(.A(n_58717), .B(n_40120), .C(n_57515), .D(n_39207),
		 .Z(n_48734));
	notech_ao4 i_5626174(.A(n_58717), .B(n_40127), .C(n_57515), .D(n_39205),
		 .Z(n_48728));
	notech_ao4 i_5526173(.A(n_58719), .B(n_40128), .C(n_57515), .D(n_39204),
		 .Z(n_48722));
	notech_ao4 i_5426172(.A(n_58717), .B(n_40126), .C(n_57515), .D(n_39202),
		 .Z(n_48716));
	notech_ao4 i_5326171(.A(n_58717), .B(n_40124), .C(n_57513), .D(n_39201),
		 .Z(n_48710));
	notech_ao4 i_5226170(.A(n_58717), .B(n_40125), .C(n_57513), .D(n_39199),
		 .Z(n_48704));
	notech_ao4 i_5126169(.A(n_58717), .B(n_40121), .C(n_57513), .D(n_39198),
		 .Z(n_48698));
	notech_ao4 i_5026168(.A(n_58717), .B(n_40113), .C(n_57515), .D(n_39196),
		 .Z(n_48692));
	notech_ao4 i_4926167(.A(n_58717), .B(n_40131), .C(n_57513), .D(n_39195),
		 .Z(n_48686));
	notech_ao4 i_4826166(.A(n_58719), .B(n_40144), .C(n_57509), .D(n_39193),
		 .Z(n_48680));
	notech_ao4 i_4726165(.A(n_58719), .B(n_40142), .C(n_57507), .D(n_39192),
		 .Z(n_48674));
	notech_ao4 i_4626164(.A(n_58719), .B(n_40143), .C(n_57507), .D(n_39190),
		 .Z(n_48668));
	notech_ao4 i_4526163(.A(n_58719), .B(n_40141), .C(n_57509), .D(n_39189),
		 .Z(n_48662));
	notech_ao4 i_4426162(.A(n_58719), .B(n_40139), .C(n_57509), .D(n_39187),
		 .Z(n_48656));
	notech_ao4 i_4326161(.A(n_58719), .B(n_40140), .C(n_57509), .D(n_39186),
		 .Z(n_48650));
	notech_ao4 i_4226160(.A(n_58719), .B(n_40138), .C(n_57507), .D(n_39184),
		 .Z(n_48644));
	notech_ao4 i_4126159(.A(n_58719), .B(n_40136), .C(n_57507), .D(n_39183),
		 .Z(n_48638));
	notech_ao4 i_3926157(.A(n_58719), .B(n_40137), .C(n_57507), .D(n_39181),
		 .Z(n_48626));
	notech_ao4 i_3826156(.A(n_58719), .B(n_40134), .C(n_57507), .D(n_39179),
		 .Z(n_48620));
	notech_ao4 i_3726155(.A(n_58725), .B(n_40135), .C(n_57507), .D(n_39178),
		 .Z(n_48614));
	notech_ao4 i_3626154(.A(n_58730), .B(n_40132), .C(n_57509), .D(n_39176),
		 .Z(n_48608));
	notech_ao4 i_3526153(.A(n_58730), .B(n_40133), .C(n_57509), .D(n_39175),
		 .Z(n_48602));
	notech_ao4 i_3426152(.A(n_58730), .B(n_40114), .C(n_57509), .D(n_39173),
		 .Z(n_48596));
	notech_ao4 i_3326151(.A(n_58730), .B(n_40115), .C(n_57509), .D(n_39172),
		 .Z(n_48590));
	notech_ao4 i_3226150(.A(n_58730), .B(n_40116), .C(n_57509), .D(n_39170),
		 .Z(n_48584));
	notech_ao4 i_3126149(.A(n_58728), .B(n_40117), .C(n_57509), .D(n_39169),
		 .Z(n_48578));
	notech_ao4 i_3026148(.A(n_58728), .B(n_40118), .C(n_57509), .D(n_39167),
		 .Z(n_48572));
	notech_ao4 i_2226140(.A(n_58730), .B(n_40156), .C(n_57509), .D(n_39155),
		 .Z(n_48524));
	notech_ao4 i_2126139(.A(n_58730), .B(n_40155), .C(n_57509), .D(n_39154),
		 .Z(n_48518));
	notech_ao4 i_1926137(.A(n_58730), .B(n_40153), .C(n_57509), .D(n_39151),
		 .Z(n_48506));
	notech_ao4 i_1826136(.A(n_58734), .B(n_40152), .C(n_57520), .D(n_39149),
		 .Z(n_48500));
	notech_ao4 i_1726135(.A(n_58730), .B(n_40164), .C(n_57520), .D(n_39148),
		 .Z(n_48494));
	notech_ao4 i_1626134(.A(n_58734), .B(n_40149), .C(n_57520), .D(n_39146),
		 .Z(n_48488));
	notech_ao4 i_1226130(.A(n_58734), .B(n_40168), .C(n_57520), .D(n_39140),
		 .Z(n_48464));
	notech_ao4 i_1126129(.A(n_58734), .B(n_40169), .C(n_57520), .D(n_39139),
		 .Z(n_48458));
	notech_ao4 i_1026128(.A(n_58730), .B(n_40170), .C(n_57520), .D(n_39137),
		 .Z(n_48452));
	notech_ao4 i_826126(.A(n_58730), .B(n_40146), .C(n_57518), .D(n_39134), 
		.Z(n_48440));
	notech_ao4 i_726125(.A(n_58730), .B(n_40119), .C(n_57520), .D(n_39133), 
		.Z(n_48434));
	notech_ao4 i_626124(.A(n_58730), .B(n_40130), .C(n_57520), .D(n_39131), 
		.Z(n_48428));
	notech_ao4 i_426122(.A(n_58730), .B(n_40212), .C(n_57520), .D(n_39128), 
		.Z(n_48416));
	notech_ao4 i_226120(.A(n_58728), .B(n_40148), .C(n_57524), .D(n_39125), 
		.Z(n_48404));
	notech_ao4 i_17026499(.A(n_58725), .B(n_40061), .C(n_57524), .D(n_39749)
		, .Z(n_44092));
	notech_ao4 i_14726476(.A(n_58725), .B(n_40038), .C(n_57524), .D(n_39710)
		, .Z(n_43954));
	notech_ao4 i_13926468(.A(n_58725), .B(n_40030), .C(n_57524), .D(n_39695)
		, .Z(n_43906));
	notech_and2 i_6330(.A(imm_sz[0]), .B(i_ptr[0]), .Z(n_2835));
	notech_or4 i_12(.A(fsm[4]), .B(fsm[3]), .C(fsm[2]), .D(n_38659), .Z(n_2834
		));
	notech_or4 i_6340(.A(fsm[3]), .B(fsm[0]), .C(fsm[1]), .D(n_2830), .Z(n_2833
		));
	notech_nand2 i_504(.A(fsm[2]), .B(n_38664), .Z(n_2830));
	notech_or2 i_075012(.A(n_58831), .B(pc_req), .Z(n_2829));
	notech_or4 i_6338(.A(fsm[2]), .B(n_2825), .C(fsm[0]), .D(n_38661), .Z(n_2828
		));
	notech_or2 i_477(.A(fsm[4]), .B(fsm[3]), .Z(n_2825));
	notech_and3 i_434(.A(n_40211), .B(n_40120), .C(n_40121), .Z(n_2821));
	notech_and4 i_425(.A(n_2083), .B(n_40128), .C(n_40127), .D(n_40126), .Z(n_2819
		));
	notech_or2 i_294792731(.A(n_39117), .B(pfx_sz[0]), .Z(n_170793328));
	notech_and2 i_288892732(.A(lenpc1[6]), .B(n_58407), .Z(n_170893329));
	notech_ao3 i_294992733(.A(n_59602), .B(n_163793258), .C(n_2849), .Z(n_170993330
		));
	notech_ao3 i_295092734(.A(n_59602), .B(n_163893259), .C(n_2849), .Z(n_171093331
		));
	notech_ao3 i_295292735(.A(n_163993260), .B(n_59596), .C(n_2849), .Z(n_171193332
		));
	notech_ao3 i_3440(.A(n_59596), .B(in128[0]), .C(n_56589), .Z(n_171293333
		));
	notech_ao3 i_3513(.A(opz[2]), .B(n_59596), .C(n_56589), .Z(n_171393334)
		);
	notech_ao3 i_3515(.A(n_1740), .B(n_59596), .C(n_56589), .Z(n_171493335)
		);
	notech_nor2 i_3516(.A(n_5392), .B(int_excl[0]), .Z(n_171593336));
	notech_nor2 i_3517(.A(n_5392), .B(n_164093261), .Z(n_171693337));
	notech_nor2 i_3518(.A(n_5392), .B(n_164193262), .Z(n_171793338));
	notech_ao3 i_3537(.A(n_38415), .B(n_2844), .C(n_2872), .Z(n_171893339)
		);
	notech_ao3 i_3764(.A(n_59595), .B(n_40171), .C(n_56589), .Z(n_171993340)
		);
	notech_ao3 i_3792(.A(n_59595), .B(in128[16]), .C(n_56589), .Z(n_172093341
		));
	notech_ao3 i_3794(.A(n_59596), .B(in128[18]), .C(n_56589), .Z(n_172193342
		));
	notech_ao3 i_3795(.A(n_59595), .B(\to_acu2_0[0] ), .C(n_56589), .Z(n_172293343
		));
	notech_ao3 i_3798(.A(n_59595), .B(\to_acu2_0[2] ), .C(n_2849), .Z(n_172393344
		));
	notech_ao3 i_3800(.A(n_59595), .B(\to_acu2_0[4] ), .C(n_56589), .Z(n_172493345
		));
	notech_and4 i_423(.A(n_40125), .B(n_40124), .C(n_40123), .D(n_40122), .Z
		(n_2816));
	notech_reg term_f_reg(.CP(n_61914), .D(n_60652), .CD(n_61353), .Q(term_f
		));
	notech_reg db67_reg(.CP(n_61914), .D(n_30164), .CD(n_61353), .Q(db67));
	notech_mux2 i_35195(.S(n_46591), .A(db67), .B(n_251491361), .Z(n_30164)
		);
	notech_reg_set fpu_indrm_reg_0(.CP(n_61914), .D(n_30170), .SD(1'b1), .Q(\fpu_indrm[0] 
		));
	notech_mux2 i_35203(.S(\nbus_13559[0] ), .A(\fpu_indrm[0] ), .B(n_172293343
		), .Z(n_30170));
	notech_reg_set fpu_indrm_reg_2(.CP(n_61914), .D(n_30176), .SD(1'b1), .Q(\fpu_indrm[2] 
		));
	notech_mux2 i_35211(.S(\nbus_13559[0] ), .A(\fpu_indrm[2] ), .B(n_172393344
		), .Z(n_30176));
	notech_or4 i_65732(.A(n_2810), .B(n_2807), .C(n_2803), .D(n_2800), .Z(n_2812
		));
	notech_reg_set fpu_indrm_reg_3(.CP(n_61914), .D(n_30182), .SD(1'b1), .Q(\fpu_indrm[3] 
		));
	notech_mux2 i_35219(.S(\nbus_13559[0] ), .A(\fpu_indrm[3] ), .B(n_162593246
		), .Z(n_30182));
	notech_reg_set fpu_indrm_reg_4(.CP(n_61914), .D(n_30188), .SD(1'b1), .Q(\fpu_indrm[4] 
		));
	notech_mux2 i_35227(.S(\nbus_13559[0] ), .A(\fpu_indrm[4] ), .B(n_172493345
		), .Z(n_30188));
	notech_or4 i_411(.A(\to_acu2_0[79] ), .B(\to_acu2_0[47] ), .C(\to_acu2_0[45] 
		), .D(\to_acu2_0[46] ), .Z(n_2810));
	notech_reg_set fpu_indrm_reg_7(.CP(n_61914), .D(n_30194), .SD(1'b1), .Q(\fpu_indrm[7] 
		));
	notech_mux2 i_35235(.S(\nbus_13559[0] ), .A(\fpu_indrm[7] ), .B(n_162693247
		), .Z(n_30194));
	notech_reg_set fpu_modrm_reg_0(.CP(n_61914), .D(n_30200), .SD(1'b1), .Q(\fpu_modrm[0] 
		));
	notech_mux2 i_35243(.S(\nbus_13559[0] ), .A(\fpu_modrm[0] ), .B(n_172093341
		), .Z(n_30200));
	notech_reg_set fpu_modrm_reg_1(.CP(n_61914), .D(n_30206), .SD(1'b1), .Q(\fpu_modrm[1] 
		));
	notech_mux2 i_35251(.S(\nbus_13559[0] ), .A(\fpu_modrm[1] ), .B(n_162493245
		), .Z(n_30206));
	notech_or4 i_410(.A(\to_acu2_0[44] ), .B(\to_acu2_0[42] ), .C(\to_acu2_0[43] 
		), .D(\to_acu2_0[41] ), .Z(n_2807));
	notech_reg_set fpu_modrm_reg_2(.CP(n_61914), .D(n_30212), .SD(1'b1), .Q(\fpu_modrm[2] 
		));
	notech_mux2 i_35259(.S(\nbus_13559[0] ), .A(\fpu_modrm[2] ), .B(n_172193342
		), .Z(n_30212));
	notech_reg displc_reg_0(.CP(n_61914), .D(n_30218), .CD(n_61353), .Q(displc
		[0]));
	notech_mux2 i_35267(.S(n_3136), .A(n_252091367), .B(displc[0]), .Z(n_30218
		));
	notech_reg displc_reg_1(.CP(n_61912), .D(n_30224), .CD(n_61353), .Q(displc
		[1]));
	notech_mux2 i_35275(.S(n_3136), .A(n_162093241), .B(displc[1]), .Z(n_30224
		));
	notech_reg displc_reg_2(.CP(n_61912), .D(n_30230), .CD(n_61353), .Q(displc
		[2]));
	notech_mux2 i_35283(.S(n_3136), .A(n_162193242), .B(displc[2]), .Z(n_30230
		));
	notech_or4 i_409(.A(\to_acu2_0[38] ), .B(\to_acu2_0[40] ), .C(\to_acu2_0[36] 
		), .D(\to_acu2_0[37] ), .Z(n_2803));
	notech_reg sib_dec_reg(.CP(n_61912), .D(n_30236), .CD(n_61353), .Q(sib_dec
		));
	notech_mux2 i_35291(.S(n_3137), .A(n_41571), .B(sib_dec), .Z(n_30236));
	notech_reg mod_dec_reg(.CP(n_61912), .D(n_30242), .CD(n_61353), .Q(mod_dec
		));
	notech_mux2 i_35299(.S(n_3138), .A(n_171993340), .B(mod_dec), .Z(n_30242
		));
	notech_reg imm2_reg_0(.CP(n_61912), .D(n_30248), .CD(n_61353), .Q(\imm2[0] 
		));
	notech_mux2 i_35307(.S(n_54239), .A(\imm2[0] ), .B(n_44631), .Z(n_30248)
		);
	notech_nand3 i_408(.A(n_40133), .B(n_40132), .C(n_2079), .Z(n_2800));
	notech_reg imm2_reg_1(.CP(n_61914), .D(n_30254), .CD(n_61353), .Q(\imm2[1] 
		));
	notech_mux2 i_35315(.S(n_54239), .A(\imm2[1] ), .B(n_44637), .Z(n_30254)
		);
	notech_reg imm2_reg_2(.CP(n_61914), .D(n_30260), .CD(n_61353), .Q(\imm2[2] 
		));
	notech_mux2 i_35323(.S(n_54239), .A(\imm2[2] ), .B(n_44643), .Z(n_30260)
		);
	notech_nao3 i_157(.A(n_2120), .B(n_2864), .C(fpu), .Z(n_2798));
	notech_reg imm2_reg_3(.CP(n_61912), .D(n_30266), .CD(n_61353), .Q(\imm2[3] 
		));
	notech_mux2 i_35331(.S(n_54233), .A(\imm2[3] ), .B(n_44649), .Z(n_30266)
		);
	notech_ao4 i_223153(.A(n_57524), .B(n_38676), .C(n_58728), .D(n_38666), 
		.Z(n_2797));
	notech_reg imm2_reg_4(.CP(n_61912), .D(n_30272), .CD(n_61351), .Q(\imm2[4] 
		));
	notech_mux2 i_35339(.S(n_54233), .A(\imm2[4] ), .B(n_44655), .Z(n_30272)
		);
	notech_reg imm2_reg_5(.CP(n_61912), .D(n_30278), .CD(n_61351), .Q(\imm2[5] 
		));
	notech_mux2 i_35347(.S(n_54233), .A(\imm2[5] ), .B(n_44661), .Z(n_30278)
		);
	notech_ao4 i_323154(.A(n_57520), .B(n_38678), .C(n_38834), .D(n_38668), 
		.Z(n_2795));
	notech_reg imm2_reg_6(.CP(n_61917), .D(n_30284), .CD(n_61351), .Q(\imm2[6] 
		));
	notech_mux2 i_35355(.S(n_54239), .A(\imm2[6] ), .B(n_44667), .Z(n_30284)
		);
	notech_reg imm2_reg_7(.CP(n_61917), .D(n_30290), .CD(n_61351), .Q(\imm2[7] 
		));
	notech_mux2 i_35363(.S(n_54239), .A(\imm2[7] ), .B(n_44673), .Z(n_30290)
		);
	notech_ao4 i_70499(.A(n_58831), .B(n_40194), .C(n_1995), .D(n_39836), .Z
		(n_2793));
	notech_reg imm2_reg_8(.CP(n_61917), .D(n_30296), .CD(n_61351), .Q(\imm2[8] 
		));
	notech_mux2 i_35371(.S(n_54239), .A(\imm2[8] ), .B(n_44679), .Z(n_30296)
		);
	notech_reg imm2_reg_9(.CP(n_61917), .D(n_30302), .CD(n_61353), .Q(\imm2[9] 
		));
	notech_mux2 i_35379(.S(n_54239), .A(\imm2[9] ), .B(n_44685), .Z(n_30302)
		);
	notech_reg imm2_reg_10(.CP(n_61917), .D(n_30308), .CD(n_61353), .Q(\imm2[10] 
		));
	notech_mux2 i_35387(.S(n_54239), .A(\imm2[10] ), .B(n_44691), .Z(n_30308
		));
	notech_ao4 i_70503(.A(n_58831), .B(n_40192), .C(n_1995), .D(n_39837), .Z
		(n_2790));
	notech_reg imm2_reg_11(.CP(n_61917), .D(n_30314), .CD(n_61353), .Q(\imm2[11] 
		));
	notech_mux2 i_35395(.S(n_54239), .A(\imm2[11] ), .B(n_44697), .Z(n_30314
		));
	notech_reg imm2_reg_12(.CP(n_61917), .D(n_30320), .CD(n_61351), .Q(\imm2[12] 
		));
	notech_mux2 i_35403(.S(n_54239), .A(\imm2[12] ), .B(n_44703), .Z(n_30320
		));
	notech_reg imm2_reg_13(.CP(n_61917), .D(n_30326), .CD(n_61353), .Q(\imm2[13] 
		));
	notech_mux2 i_35411(.S(n_54233), .A(\imm2[13] ), .B(n_44709), .Z(n_30326
		));
	notech_ao4 i_70507(.A(n_58831), .B(n_40191), .C(n_1995), .D(n_39839), .Z
		(n_2787));
	notech_reg imm2_reg_14(.CP(n_61917), .D(n_30332), .CD(n_61356), .Q(\imm2[14] 
		));
	notech_mux2 i_35419(.S(n_54233), .A(\imm2[14] ), .B(n_44715), .Z(n_30332
		));
	notech_reg imm2_reg_15(.CP(n_61917), .D(n_30338), .CD(n_61356), .Q(\imm2[15] 
		));
	notech_mux2 i_35427(.S(n_54233), .A(\imm2[15] ), .B(n_2046), .Z(n_30338)
		);
	notech_reg imm2_reg_16(.CP(n_61917), .D(n_30344), .CD(n_61356), .Q(\imm2[16] 
		));
	notech_mux2 i_35435(.S(n_54233), .A(\imm2[16] ), .B(n_2045), .Z(n_30344)
		);
	notech_ao4 i_70511(.A(n_58831), .B(n_40190), .C(n_1995), .D(n_39840), .Z
		(n_2784));
	notech_reg imm2_reg_17(.CP(n_61914), .D(n_30350), .CD(n_61356), .Q(\imm2[17] 
		));
	notech_mux2 i_35443(.S(n_54233), .A(\imm2[17] ), .B(n_2044), .Z(n_30350)
		);
	notech_reg imm2_reg_18(.CP(n_61914), .D(n_30356), .CD(n_61356), .Q(\imm2[18] 
		));
	notech_mux2 i_35451(.S(n_54233), .A(\imm2[18] ), .B(n_2043), .Z(n_30356)
		);
	notech_reg imm2_reg_19(.CP(n_61914), .D(n_30362), .CD(n_61356), .Q(\imm2[19] 
		));
	notech_mux2 i_35459(.S(n_54233), .A(\imm2[19] ), .B(n_2042), .Z(n_30362)
		);
	notech_ao4 i_70515(.A(n_58831), .B(n_40189), .C(n_1995), .D(n_39842), .Z
		(n_278191628));
	notech_reg imm2_reg_20(.CP(n_61914), .D(n_30368), .CD(n_61356), .Q(\imm2[20] 
		));
	notech_mux2 i_35467(.S(n_54233), .A(\imm2[20] ), .B(n_44751), .Z(n_30368
		));
	notech_reg imm2_reg_21(.CP(n_61914), .D(n_30374), .CD(n_61356), .Q(\imm2[21] 
		));
	notech_mux2 i_35475(.S(n_54233), .A(\imm2[21] ), .B(n_44757), .Z(n_30374
		));
	notech_reg imm2_reg_22(.CP(n_61917), .D(n_30380), .CD(n_61356), .Q(\imm2[22] 
		));
	notech_mux2 i_35483(.S(n_54233), .A(\imm2[22] ), .B(n_44763), .Z(n_30380
		));
	notech_ao4 i_70519(.A(n_58831), .B(n_40188), .C(n_1995), .D(n_39844), .Z
		(n_277891625));
	notech_reg imm2_reg_23(.CP(n_61917), .D(n_30386), .CD(n_61356), .Q(\imm2[23] 
		));
	notech_mux2 i_35491(.S(n_54233), .A(\imm2[23] ), .B(n_44769), .Z(n_30386
		));
	notech_reg imm2_reg_24(.CP(n_61917), .D(n_30392), .CD(n_61356), .Q(\imm2[24] 
		));
	notech_mux2 i_35499(.S(n_54233), .A(\imm2[24] ), .B(n_44775), .Z(n_30392
		));
	notech_reg imm2_reg_25(.CP(n_61914), .D(n_30398), .CD(n_61353), .Q(\imm2[25] 
		));
	notech_mux2 i_35507(.S(n_54233), .A(\imm2[25] ), .B(n_44781), .Z(n_30398
		));
	notech_nand3 i_323151(.A(n_265391500), .B(n_59596), .C(n_277491621), .Z(n_277591622
		));
	notech_reg imm2_reg_26(.CP(n_61914), .D(n_30404), .CD(n_61353), .Q(\imm2[26] 
		));
	notech_mux2 i_35515(.S(n_54239), .A(\imm2[26] ), .B(n_44787), .Z(n_30404
		));
	notech_nand3 i_1519(.A(n_2124), .B(opz1[2]), .C(n_59596), .Z(n_277491621
		));
	notech_reg imm2_reg_27(.CP(n_61912), .D(n_30410), .CD(n_61353), .Q(\imm2[27] 
		));
	notech_mux2 i_35523(.S(n_54244), .A(\imm2[27] ), .B(n_44793), .Z(n_30410
		));
	notech_ao4 i_627224(.A(n_57520), .B(n_39122), .C(n_58725), .D(n_39118), 
		.Z(n_277391620));
	notech_reg imm2_reg_28(.CP(n_61907), .D(n_30416), .CD(n_61353), .Q(\imm2[28] 
		));
	notech_mux2 i_35531(.S(n_54244), .A(\imm2[28] ), .B(n_44799), .Z(n_30416
		));
	notech_reg imm2_reg_29(.CP(n_61907), .D(n_30422), .CD(n_61353), .Q(\imm2[29] 
		));
	notech_mux2 i_35539(.S(n_54244), .A(\imm2[29] ), .B(n_3248), .Z(n_30422)
		);
	notech_ao4 i_2026349(.A(n_57520), .B(n_39468), .C(n_58725), .D(n_40187),
		 .Z(n_277191618));
	notech_reg imm2_reg_30(.CP(n_61907), .D(n_30428), .CD(n_61356), .Q(\imm2[30] 
		));
	notech_mux2 i_35547(.S(n_54244), .A(\imm2[30] ), .B(n_44811), .Z(n_30428
		));
	notech_reg imm2_reg_31(.CP(n_61907), .D(n_30434), .CD(n_61356), .Q(\imm2[31] 
		));
	notech_mux2 i_35555(.S(n_54244), .A(\imm2[31] ), .B(n_44817), .Z(n_30434
		));
	notech_ao4 i_6926398(.A(n_57520), .B(n_39574), .C(n_58725), .D(n_40186),
		 .Z(n_276991616));
	notech_reg imm2_reg_32(.CP(n_61907), .D(n_30440), .CD(n_61356), .Q(\imm2[32] 
		));
	notech_mux2 i_35563(.S(n_54244), .A(\imm2[32] ), .B(n_44823), .Z(n_30440
		));
	notech_reg imm2_reg_33(.CP(n_61907), .D(n_30446), .CD(n_61356), .Q(\imm2[33] 
		));
	notech_mux2 i_35571(.S(n_54245), .A(\imm2[33] ), .B(n_44829), .Z(n_30446
		));
	notech_ao4 i_7126400(.A(n_57520), .B(n_39576), .C(n_58725), .D(n_40204),
		 .Z(n_276791614));
	notech_reg imm2_reg_34(.CP(n_61907), .D(n_30452), .CD(n_61356), .Q(\imm2[34] 
		));
	notech_mux2 i_35579(.S(n_54245), .A(\imm2[34] ), .B(n_44835), .Z(n_30452
		));
	notech_reg imm2_reg_35(.CP(n_61907), .D(n_30458), .CD(n_61346), .Q(\imm2[35] 
		));
	notech_mux2 i_35587(.S(n_54245), .A(\imm2[35] ), .B(n_44841), .Z(n_30458
		));
	notech_ao4 i_7226401(.A(n_57518), .B(n_39577), .C(n_58725), .D(n_40205),
		 .Z(n_276591612));
	notech_reg imm2_reg_36(.CP(n_61907), .D(n_30464), .CD(n_61346), .Q(\imm2[36] 
		));
	notech_mux2 i_35595(.S(n_54245), .A(\imm2[36] ), .B(n_44847), .Z(n_30464
		));
	notech_reg imm2_reg_37(.CP(n_61907), .D(n_30470), .CD(n_61346), .Q(\imm2[37] 
		));
	notech_mux2 i_35603(.S(n_54245), .A(\imm2[37] ), .B(n_44853), .Z(n_30470
		));
	notech_ao4 i_7326402(.A(n_57515), .B(n_39578), .C(n_58725), .D(n_40185),
		 .Z(n_276391610));
	notech_reg imm2_reg_38(.CP(n_61905), .D(n_30476), .CD(n_61346), .Q(\imm2[38] 
		));
	notech_mux2 i_35611(.S(n_54245), .A(\imm2[38] ), .B(n_44859), .Z(n_30476
		));
	notech_reg imm2_reg_39(.CP(n_61905), .D(n_30482), .CD(n_61346), .Q(\imm2[39] 
		));
	notech_mux2 i_35619(.S(n_54245), .A(\imm2[39] ), .B(n_44865), .Z(n_30482
		));
	notech_ao4 i_7426403(.A(n_57515), .B(n_39579), .C(n_58728), .D(n_40184),
		 .Z(n_276191608));
	notech_reg imm2_reg_40(.CP(n_61905), .D(n_30488), .CD(n_61346), .Q(\imm2[40] 
		));
	notech_mux2 i_35627(.S(n_54244), .A(\imm2[40] ), .B(n_44871), .Z(n_30488
		));
	notech_reg imm2_reg_41(.CP(n_61905), .D(n_30494), .CD(n_61346), .Q(\imm2[41] 
		));
	notech_mux2 i_35635(.S(n_54244), .A(\imm2[41] ), .B(n_44877), .Z(n_30494
		));
	notech_ao4 i_7526404(.A(n_57515), .B(n_39580), .C(n_58728), .D(n_40211),
		 .Z(n_275991606));
	notech_reg imm2_reg_42(.CP(n_61905), .D(n_30500), .CD(n_61346), .Q(\imm2[42] 
		));
	notech_mux2 i_35643(.S(n_54244), .A(\imm2[42] ), .B(n_44883), .Z(n_30500
		));
	notech_reg imm2_reg_43(.CP(n_61905), .D(n_30506), .CD(n_61346), .Q(\imm2[43] 
		));
	notech_mux2 i_35651(.S(n_54239), .A(\imm2[43] ), .B(n_44889), .Z(n_30506
		));
	notech_ao4 i_7626405(.A(n_57518), .B(n_39581), .C(n_58728), .D(n_40203),
		 .Z(n_275791604));
	notech_reg imm2_reg_44(.CP(n_61905), .D(n_30512), .CD(n_61346), .Q(\imm2[44] 
		));
	notech_mux2 i_35659(.S(n_54244), .A(\imm2[44] ), .B(n_44895), .Z(n_30512
		));
	notech_reg imm2_reg_45(.CP(n_61905), .D(n_30518), .CD(n_61346), .Q(\imm2[45] 
		));
	notech_mux2 i_35667(.S(n_54244), .A(\imm2[45] ), .B(n_44901), .Z(n_30518
		));
	notech_ao4 i_7726406(.A(n_57518), .B(n_39582), .C(n_58728), .D(n_40183),
		 .Z(n_275591602));
	notech_reg imm2_reg_46(.CP(n_61905), .D(n_30524), .CD(n_61344), .Q(\imm2[46] 
		));
	notech_mux2 i_35675(.S(n_54244), .A(\imm2[46] ), .B(n_44907), .Z(n_30524
		));
	notech_reg imm2_reg_47(.CP(n_61905), .D(n_30530), .CD(n_61344), .Q(\imm2[47] 
		));
	notech_mux2 i_35683(.S(n_54244), .A(\imm2[47] ), .B(n_44913), .Z(n_30530
		));
	notech_ao4 i_7826407(.A(n_57515), .B(n_39583), .C(n_58728), .D(n_40182),
		 .Z(n_275391600));
	notech_reg imm1_reg_0(.CP(n_61905), .D(n_30536), .CD(n_61344), .Q(\imm1[0] 
		));
	notech_mux2 i_35691(.S(n_57661), .A(\imm1[0] ), .B(n_38409), .Z(n_30536)
		);
	notech_reg imm1_reg_1(.CP(n_61912), .D(n_30542), .CD(n_61344), .Q(\imm1[1] 
		));
	notech_mux2 i_35699(.S(n_57661), .A(\imm1[1] ), .B(n_38410), .Z(n_30542)
		);
	notech_ao4 i_7926408(.A(n_57515), .B(n_39584), .C(n_58728), .D(n_40181),
		 .Z(n_275191598));
	notech_reg imm1_reg_2(.CP(n_61912), .D(n_30548), .CD(n_61344), .Q(\imm1[2] 
		));
	notech_mux2 i_35707(.S(n_57661), .A(\imm1[2] ), .B(n_38412), .Z(n_30548)
		);
	notech_reg imm1_reg_3(.CP(n_61912), .D(n_30554), .CD(n_61346), .Q(\imm1[3] 
		));
	notech_mux2 i_35715(.S(n_57655), .A(\imm1[3] ), .B(n_38413), .Z(n_30554)
		);
	notech_ao4 i_8026409(.A(n_57515), .B(n_39585), .C(n_58728), .D(n_40180),
		 .Z(n_274991596));
	notech_reg imm1_reg_4(.CP(n_61912), .D(n_30560), .CD(n_61346), .Q(\imm1[4] 
		));
	notech_mux2 i_35723(.S(n_57655), .A(\imm1[4] ), .B(n_38414), .Z(n_30560)
		);
	notech_reg imm1_reg_5(.CP(n_61912), .D(n_30566), .CD(n_61344), .Q(\imm1[5] 
		));
	notech_mux2 i_35731(.S(n_57655), .A(\imm1[5] ), .B(n_38416), .Z(n_30566)
		);
	notech_ao4 i_8126410(.A(n_57515), .B(n_39586), .C(n_58728), .D(n_40179),
		 .Z(n_274791594));
	notech_reg imm1_reg_6(.CP(n_61912), .D(n_30572), .CD(n_61344), .Q(\imm1[6] 
		));
	notech_mux2 i_35739(.S(n_57661), .A(\imm1[6] ), .B(n_38418), .Z(n_30572)
		);
	notech_reg imm1_reg_7(.CP(n_61912), .D(n_30578), .CD(n_61344), .Q(\imm1[7] 
		));
	notech_mux2 i_35747(.S(n_57661), .A(\imm1[7] ), .B(n_38419), .Z(n_30578)
		);
	notech_ao4 i_8226411(.A(n_57515), .B(n_39587), .C(n_58728), .D(n_40178),
		 .Z(n_274591592));
	notech_reg imm1_reg_8(.CP(n_61912), .D(n_30584), .CD(n_61351), .Q(\imm1[8] 
		));
	notech_mux2 i_35755(.S(n_57661), .A(\imm1[8] ), .B(n_38420), .Z(n_30584)
		);
	notech_reg imm1_reg_9(.CP(n_61912), .D(n_30590), .CD(n_61351), .Q(\imm1[9] 
		));
	notech_mux2 i_35763(.S(n_57661), .A(\imm1[9] ), .B(n_38422), .Z(n_30590)
		);
	notech_ao4 i_8326412(.A(n_57518), .B(n_39589), .C(n_58728), .D(n_40177),
		 .Z(n_274391590));
	notech_reg imm1_reg_10(.CP(n_61912), .D(n_30596), .CD(n_61351), .Q(\imm1[10] 
		));
	notech_mux2 i_35771(.S(n_57661), .A(\imm1[10] ), .B(n_38423), .Z(n_30596
		));
	notech_reg imm1_reg_11(.CP(n_61912), .D(n_30602), .CD(n_61351), .Q(\imm1[11] 
		));
	notech_mux2 i_35779(.S(n_57661), .A(\imm1[11] ), .B(n_38424), .Z(n_30602
		));
	notech_ao4 i_8426413(.A(n_57518), .B(n_39591), .C(n_58705), .D(n_40213),
		 .Z(n_274191588));
	notech_reg imm1_reg_12(.CP(n_61907), .D(n_30608), .CD(n_61351), .Q(\imm1[12] 
		));
	notech_mux2 i_35787(.S(n_57661), .A(\imm1[12] ), .B(n_38426), .Z(n_30608
		));
	notech_reg imm1_reg_13(.CP(n_61907), .D(n_30614), .CD(n_61351), .Q(\imm1[13] 
		));
	notech_mux2 i_35795(.S(n_57655), .A(\imm1[13] ), .B(n_38427), .Z(n_30614
		));
	notech_ao4 i_8526414(.A(n_58705), .B(n_40176), .C(n_57518), .D(n_39592),
		 .Z(n_273991586));
	notech_reg imm1_reg_14(.CP(n_61907), .D(n_30620), .CD(n_61351), .Q(\imm1[14] 
		));
	notech_mux2 i_35803(.S(n_57655), .A(\imm1[14] ), .B(n_38429), .Z(n_30620
		));
	notech_reg imm1_reg_15(.CP(n_61907), .D(n_30626), .CD(n_61351), .Q(\imm1[15] 
		));
	notech_mux2 i_35811(.S(n_57655), .A(\imm1[15] ), .B(n_38430), .Z(n_30626
		));
	notech_ao4 i_8626415(.A(n_57518), .B(n_39594), .C(n_58705), .D(n_40175),
		 .Z(n_273791584));
	notech_reg imm1_reg_16(.CP(n_61907), .D(n_30632), .CD(n_61351), .Q(\imm1[16] 
		));
	notech_mux2 i_35819(.S(n_57655), .A(\imm1[16] ), .B(n_38432), .Z(n_30632
		));
	notech_reg imm1_reg_17(.CP(n_61907), .D(n_30638), .CD(n_61351), .Q(\imm1[17] 
		));
	notech_mux2 i_35827(.S(n_57655), .A(\imm1[17] ), .B(n_38433), .Z(n_30638
		));
	notech_ao4 i_8726416(.A(n_57518), .B(n_39596), .C(n_58705), .D(n_40198),
		 .Z(n_273591582));
	notech_reg imm1_reg_18(.CP(n_61907), .D(n_30644), .CD(n_61351), .Q(\imm1[18] 
		));
	notech_mux2 i_35835(.S(n_57655), .A(\imm1[18] ), .B(n_38435), .Z(n_30644
		));
	notech_reg imm1_reg_19(.CP(n_61907), .D(n_30650), .CD(n_61346), .Q(\imm1[19] 
		));
	notech_mux2 i_35843(.S(n_57655), .A(\imm1[19] ), .B(n_38436), .Z(n_30650
		));
	notech_ao4 i_8826417(.A(n_57518), .B(n_39598), .C(n_58705), .D(n_40199),
		 .Z(n_273391580));
	notech_reg imm1_reg_20(.CP(n_61907), .D(n_30656), .CD(n_61346), .Q(\imm1[20] 
		));
	notech_mux2 i_35851(.S(n_57655), .A(\imm1[20] ), .B(n_38437), .Z(n_30656
		));
	notech_reg imm1_reg_21(.CP(n_61907), .D(n_30662), .CD(n_61346), .Q(\imm1[21] 
		));
	notech_mux2 i_35859(.S(n_57655), .A(\imm1[21] ), .B(n_38438), .Z(n_30662
		));
	notech_ao4 i_8926418(.A(n_57518), .B(n_39600), .C(n_58705), .D(n_40200),
		 .Z(n_273191578));
	notech_reg imm1_reg_22(.CP(n_61924), .D(n_30668), .CD(n_61346), .Q(\imm1[22] 
		));
	notech_mux2 i_35867(.S(n_57655), .A(\imm1[22] ), .B(n_38439), .Z(n_30668
		));
	notech_reg imm1_reg_23(.CP(n_61924), .D(n_30674), .CD(n_61346), .Q(\imm1[23] 
		));
	notech_mux2 i_35875(.S(n_57655), .A(\imm1[23] ), .B(n_38440), .Z(n_30674
		));
	notech_ao4 i_9026419(.A(n_57518), .B(n_39603), .C(n_58702), .D(n_40201),
		 .Z(n_272991576));
	notech_reg imm1_reg_24(.CP(n_61924), .D(n_30680), .CD(n_61351), .Q(\imm1[24] 
		));
	notech_mux2 i_35883(.S(n_57655), .A(\imm1[24] ), .B(n_38441), .Z(n_30680
		));
	notech_reg imm1_reg_25(.CP(n_61924), .D(n_30686), .CD(n_61351), .Q(\imm1[25] 
		));
	notech_mux2 i_35891(.S(n_57655), .A(\imm1[25] ), .B(n_38442), .Z(n_30686
		));
	notech_ao4 i_9126420(.A(n_57518), .B(n_39604), .C(n_58705), .D(n_40202),
		 .Z(n_272791574));
	notech_reg imm1_reg_26(.CP(n_61924), .D(n_30692), .CD(n_61351), .Q(\imm1[26] 
		));
	notech_mux2 i_35899(.S(n_57661), .A(\imm1[26] ), .B(n_38443), .Z(n_30692
		));
	notech_reg imm1_reg_27(.CP(n_61924), .D(n_30698), .CD(n_61346), .Q(\imm1[27] 
		));
	notech_mux2 i_35907(.S(n_57666), .A(\imm1[27] ), .B(n_38444), .Z(n_30698
		));
	notech_ao4 i_9226421(.A(n_57518), .B(n_39606), .C(n_58705), .D(n_40174),
		 .Z(n_272591572));
	notech_reg imm1_reg_28(.CP(n_61924), .D(n_30704), .CD(n_61346), .Q(\imm1[28] 
		));
	notech_mux2 i_35915(.S(n_57666), .A(\imm1[28] ), .B(n_38445), .Z(n_30704
		));
	notech_reg imm1_reg_29(.CP(n_61924), .D(n_30710), .CD(n_61356), .Q(\imm1[29] 
		));
	notech_mux2 i_35923(.S(n_57666), .A(\imm1[29] ), .B(n_38446), .Z(n_30710
		));
	notech_ao4 i_9326422(.A(n_57507), .B(n_39608), .C(n_58705), .D(n_40196),
		 .Z(n_272391570));
	notech_reg imm1_reg_30(.CP(n_61924), .D(n_30716), .CD(n_61363), .Q(\imm1[30] 
		));
	notech_mux2 i_35931(.S(n_57666), .A(\imm1[30] ), .B(n_38447), .Z(n_30716
		));
	notech_reg imm1_reg_31(.CP(n_61924), .D(n_30722), .CD(n_61363), .Q(\imm1[31] 
		));
	notech_mux2 i_35939(.S(n_57666), .A(\imm1[31] ), .B(n_38448), .Z(n_30722
		));
	notech_ao4 i_9426423(.A(n_57495), .B(n_39609), .C(n_58707), .D(n_40197),
		 .Z(n_272191568));
	notech_reg imm1_reg_32(.CP(n_61924), .D(n_30728), .CD(n_61363), .Q(\imm1[32] 
		));
	notech_mux2 i_35947(.S(n_57666), .A(\imm1[32] ), .B(n_38449), .Z(n_30728
		));
	notech_reg imm1_reg_33(.CP(n_61924), .D(n_30734), .CD(n_61363), .Q(\imm1[33] 
		));
	notech_mux2 i_35955(.S(n_57667), .A(\imm1[33] ), .B(n_38450), .Z(n_30734
		));
	notech_ao4 i_9526424(.A(n_57495), .B(n_39611), .C(n_58707), .D(n_40208),
		 .Z(n_271991566));
	notech_reg imm1_reg_34(.CP(n_61924), .D(n_30740), .CD(n_61363), .Q(\imm1[34] 
		));
	notech_mux2 i_35963(.S(n_57667), .A(\imm1[34] ), .B(n_38451), .Z(n_30740
		));
	notech_reg imm1_reg_35(.CP(n_61922), .D(n_30746), .CD(n_61363), .Q(\imm1[35] 
		));
	notech_mux2 i_35971(.S(n_57667), .A(\imm1[35] ), .B(n_38452), .Z(n_30746
		));
	notech_ao4 i_9626425(.A(n_57495), .B(n_39613), .C(n_58707), .D(n_40207),
		 .Z(n_271791564));
	notech_reg imm1_reg_36(.CP(n_61922), .D(n_30752), .CD(n_61363), .Q(\imm1[36] 
		));
	notech_mux2 i_35979(.S(n_57667), .A(\imm1[36] ), .B(n_38453), .Z(n_30752
		));
	notech_reg imm1_reg_37(.CP(n_61922), .D(n_30758), .CD(n_61363), .Q(\imm1[37] 
		));
	notech_mux2 i_35987(.S(n_57667), .A(\imm1[37] ), .B(n_38579), .Z(n_30758
		));
	notech_ao4 i_9726426(.A(n_57495), .B(n_39614), .C(n_58707), .D(n_40206),
		 .Z(n_271591562));
	notech_reg imm1_reg_38(.CP(n_61924), .D(n_30764), .CD(n_61363), .Q(\imm1[38] 
		));
	notech_mux2 i_35995(.S(n_57667), .A(\imm1[38] ), .B(n_38582), .Z(n_30764
		));
	notech_reg imm1_reg_39(.CP(n_61924), .D(n_30770), .CD(n_61363), .Q(\imm1[39] 
		));
	notech_mux2 i_36003(.S(n_57667), .A(\imm1[39] ), .B(n_38584), .Z(n_30770
		));
	notech_ao4 i_9826427(.A(n_57495), .B(n_39616), .C(n_58707), .D(n_40173),
		 .Z(n_271391560));
	notech_reg imm1_reg_40(.CP(n_61924), .D(n_30776), .CD(n_61363), .Q(\imm1[40] 
		));
	notech_mux2 i_36011(.S(n_57666), .A(\imm1[40] ), .B(n_38587), .Z(n_30776
		));
	notech_reg imm1_reg_41(.CP(n_61924), .D(n_30782), .CD(n_61363), .Q(\imm1[41] 
		));
	notech_mux2 i_36019(.S(n_57666), .A(\imm1[41] ), .B(n_38454), .Z(n_30782
		));
	notech_ao4 i_9926428(.A(n_57495), .B(n_39617), .C(n_58705), .D(n_40172),
		 .Z(n_271191558));
	notech_reg imm1_reg_42(.CP(n_61924), .D(n_30788), .CD(n_61363), .Q(\imm1[42] 
		));
	notech_mux2 i_36027(.S(n_57666), .A(\imm1[42] ), .B(n_38455), .Z(n_30788
		));
	notech_reg imm1_reg_43(.CP(n_61928), .D(n_30794), .CD(n_61363), .Q(\imm1[43] 
		));
	notech_mux2 i_36035(.S(n_57661), .A(\imm1[43] ), .B(n_38457), .Z(n_30794
		));
	notech_ao4 i_10026429(.A(n_57495), .B(n_39618), .C(n_58705), .D(n_39991)
		, .Z(n_270991556));
	notech_reg imm1_reg_44(.CP(n_61928), .D(n_30800), .CD(n_61361), .Q(\imm1[44] 
		));
	notech_mux2 i_36043(.S(n_57666), .A(\imm1[44] ), .B(n_38595), .Z(n_30800
		));
	notech_reg imm1_reg_45(.CP(n_61928), .D(n_30806), .CD(n_61363), .Q(\imm1[45] 
		));
	notech_mux2 i_36051(.S(n_57666), .A(\imm1[45] ), .B(n_38459), .Z(n_30806
		));
	notech_ao4 i_10126430(.A(n_57495), .B(n_39620), .C(n_58705), .D(n_39992)
		, .Z(n_270791554));
	notech_reg imm1_reg_46(.CP(n_61928), .D(n_30812), .CD(n_61363), .Q(\imm1[46] 
		));
	notech_mux2 i_36059(.S(n_57666), .A(\imm1[46] ), .B(n_38461), .Z(n_30812
		));
	notech_reg imm1_reg_47(.CP(n_61928), .D(n_30818), .CD(n_61363), .Q(\imm1[47] 
		));
	notech_mux2 i_36067(.S(n_57666), .A(\imm1[47] ), .B(n_38463), .Z(n_30818
		));
	notech_ao4 i_10226431(.A(n_57495), .B(n_39622), .C(n_58705), .D(n_39993)
		, .Z(n_270591552));
	notech_reg trig_it_reg(.CP(n_61928), .D(n_30824), .CD(n_61363), .Q(trig_it
		));
	notech_mux2 i_36075(.S(n_3139), .A(n_171893339), .B(trig_it), .Z(n_30824
		));
	notech_reg trig_itf_reg(.CP(n_61928), .D(trig_it), .CD(n_61363), .Q(trig_itf
		));
	notech_reg intf_reg(.CP(n_61928), .D(int_main), .CD(n_61363), .Q(intf)
		);
	notech_reg_set intff_reg(.CP(n_61928), .D(n_30834), .SD(1'b1), .Q(intff)
		);
	notech_mux2 i_36091(.S(n_61367), .A(intff), .B(intf), .Z(n_30834));
	notech_ao4 i_10326432(.A(n_57495), .B(n_39624), .C(n_58705), .D(n_39994)
		, .Z(n_270391550));
	notech_reg ififo_rvect4_reg_0(.CP(n_61928), .D(n_30840), .CD(n_61367), .Q
		(ififo_rvect4[0]));
	notech_mux2 i_36099(.S(\nbus_13535[0] ), .A(ififo_rvect4[0]), .B(n_161293233
		), .Z(n_30840));
	notech_reg ififo_rvect4_reg_1(.CP(n_61928), .D(n_30846), .CD(n_61367), .Q
		(ififo_rvect4[1]));
	notech_mux2 i_36107(.S(\nbus_13535[0] ), .A(ififo_rvect4[1]), .B(n_161393234
		), .Z(n_30846));
	notech_ao4 i_10426433(.A(n_57497), .B(n_39627), .C(n_58702), .D(n_39995)
		, .Z(n_270191548));
	notech_reg ififo_rvect4_reg_2(.CP(n_61928), .D(n_30852), .CD(n_61367), .Q
		(ififo_rvect4[2]));
	notech_mux2 i_36115(.S(\nbus_13535[0] ), .A(ififo_rvect4[2]), .B(n_161493235
		), .Z(n_30852));
	notech_reg ififo_rvect4_reg_3(.CP(n_61928), .D(n_30858), .CD(n_61367), .Q
		(ififo_rvect4[3]));
	notech_mux2 i_36123(.S(\nbus_13535[0] ), .A(ififo_rvect4[3]), .B(n_161593236
		), .Z(n_30858));
	notech_ao4 i_10526434(.A(n_57497), .B(n_39629), .C(n_58700), .D(n_39996)
		, .Z(n_269991546));
	notech_reg ififo_rvect4_reg_4(.CP(n_61928), .D(n_30864), .CD(n_61369), .Q
		(ififo_rvect4[4]));
	notech_mux2 i_36131(.S(\nbus_13535[0] ), .A(ififo_rvect4[4]), .B(n_161693237
		), .Z(n_30864));
	notech_reg ififo_rvect4_reg_5(.CP(n_61924), .D(n_30870), .CD(n_61369), .Q
		(ififo_rvect4[5]));
	notech_mux2 i_36139(.S(\nbus_13535[0] ), .A(ififo_rvect4[5]), .B(n_161793238
		), .Z(n_30870));
	notech_ao4 i_10626435(.A(n_57497), .B(n_39631), .C(n_58700), .D(n_39997)
		, .Z(n_269791544));
	notech_reg ififo_rvect4_reg_6(.CP(n_61924), .D(n_30876), .CD(n_61367), .Q
		(ififo_rvect4[6]));
	notech_mux2 i_36147(.S(\nbus_13535[0] ), .A(ififo_rvect4[6]), .B(n_161893239
		), .Z(n_30876));
	notech_reg ififo_rvect4_reg_7(.CP(n_61928), .D(n_30882), .CD(n_61367), .Q
		(ififo_rvect4[7]));
	notech_mux2 i_36155(.S(\nbus_13535[0] ), .A(ififo_rvect4[7]), .B(n_161993240
		), .Z(n_30882));
	notech_ao4 i_10726436(.A(n_57497), .B(n_39633), .C(n_58700), .D(n_39998)
		, .Z(n_269591542));
	notech_reg ififo_rvect3_reg_0(.CP(n_61928), .D(n_30888), .CD(n_61367), .Q
		(ififo_rvect3[0]));
	notech_mux2 i_36163(.S(\nbus_13535[0] ), .A(ififo_rvect3[0]), .B(n_46510
		), .Z(n_30888));
	notech_reg ififo_rvect3_reg_1(.CP(n_61928), .D(n_30894), .CD(n_61367), .Q
		(ififo_rvect3[1]));
	notech_mux2 i_36171(.S(\nbus_13535[0] ), .A(ififo_rvect3[1]), .B(n_46516
		), .Z(n_30894));
	notech_ao4 i_10826437(.A(n_57497), .B(n_39635), .C(n_58702), .D(n_39999)
		, .Z(n_269391540));
	notech_reg ififo_rvect3_reg_2(.CP(n_61928), .D(n_30900), .CD(n_61367), .Q
		(ififo_rvect3[2]));
	notech_mux2 i_36179(.S(\nbus_13535[0] ), .A(ififo_rvect3[2]), .B(n_46522
		), .Z(n_30900));
	notech_reg ififo_rvect3_reg_3(.CP(n_61928), .D(n_30906), .CD(n_61367), .Q
		(ififo_rvect3[3]));
	notech_mux2 i_36187(.S(\nbus_13535[0] ), .A(ififo_rvect3[3]), .B(n_46528
		), .Z(n_30906));
	notech_ao4 i_10926438(.A(n_57495), .B(n_39638), .C(n_58702), .D(n_40000)
		, .Z(n_269191538));
	notech_reg ififo_rvect3_reg_4(.CP(n_61922), .D(n_30912), .CD(n_61367), .Q
		(ififo_rvect3[4]));
	notech_mux2 i_36195(.S(\nbus_13535[0] ), .A(ififo_rvect3[4]), .B(n_46534
		), .Z(n_30912));
	notech_reg ififo_rvect3_reg_5(.CP(n_61919), .D(n_30918), .CD(n_61367), .Q
		(ififo_rvect3[5]));
	notech_mux2 i_36203(.S(\nbus_13535[0] ), .A(ififo_rvect3[5]), .B(n_46540
		), .Z(n_30918));
	notech_ao4 i_11026439(.A(n_57495), .B(n_39640), .C(n_58700), .D(n_40001)
		, .Z(n_268991536));
	notech_reg ififo_rvect3_reg_6(.CP(n_61919), .D(n_30924), .CD(n_61367), .Q
		(ififo_rvect3[6]));
	notech_mux2 i_36211(.S(\nbus_13535[0] ), .A(ififo_rvect3[6]), .B(n_46546
		), .Z(n_30924));
	notech_reg ififo_rvect3_reg_7(.CP(n_61919), .D(n_30930), .CD(n_61367), .Q
		(ififo_rvect3[7]));
	notech_mux2 i_36219(.S(\nbus_13535[0] ), .A(ififo_rvect3[7]), .B(n_46552
		), .Z(n_30930));
	notech_ao4 i_11126440(.A(n_57495), .B(n_39642), .C(n_58700), .D(n_40002)
		, .Z(n_268791534));
	notech_reg ififo_rvect2_reg_0(.CP(n_61919), .D(n_30936), .CD(n_61367), .Q
		(ififo_rvect2[0]));
	notech_mux2 i_36227(.S(n_55049), .A(ififo_rvect2[0]), .B(n_41604), .Z(n_30936
		));
	notech_reg ififo_rvect2_reg_1(.CP(n_61919), .D(n_30942), .CD(n_61367), .Q
		(ififo_rvect2[1]));
	notech_mux2 i_36235(.S(n_55049), .A(ififo_rvect2[1]), .B(n_41610), .Z(n_30942
		));
	notech_ao4 i_11226441(.A(n_57497), .B(n_39645), .C(n_58700), .D(n_40003)
		, .Z(n_268591532));
	notech_reg ififo_rvect2_reg_2(.CP(n_61919), .D(n_30948), .CD(n_61367), .Q
		(ififo_rvect2[2]));
	notech_mux2 i_36243(.S(n_55049), .A(ififo_rvect2[2]), .B(n_41616), .Z(n_30948
		));
	notech_reg ififo_rvect2_reg_3(.CP(n_61919), .D(n_30954), .CD(n_61367), .Q
		(ififo_rvect2[3]));
	notech_mux2 i_36251(.S(n_55049), .A(ififo_rvect2[3]), .B(n_41622), .Z(n_30954
		));
	notech_ao4 i_11426443(.A(n_57497), .B(n_39649), .C(n_58700), .D(n_40005)
		, .Z(n_268391530));
	notech_reg ififo_rvect2_reg_4(.CP(n_61919), .D(n_30960), .CD(n_61358), .Q
		(ififo_rvect2[4]));
	notech_mux2 i_36259(.S(n_55049), .A(ififo_rvect2[4]), .B(n_41628), .Z(n_30960
		));
	notech_reg ififo_rvect2_reg_5(.CP(n_61919), .D(n_30966), .CD(n_61358), .Q
		(ififo_rvect2[5]));
	notech_mux2 i_36267(.S(n_55049), .A(ififo_rvect2[5]), .B(n_41634), .Z(n_30966
		));
	notech_ao4 i_11526444(.A(n_57495), .B(n_39651), .C(n_58700), .D(n_40006)
		, .Z(n_268191528));
	notech_reg ififo_rvect2_reg_6(.CP(n_61919), .D(n_30972), .CD(n_61358), .Q
		(ififo_rvect2[6]));
	notech_mux2 i_36275(.S(n_55049), .A(ififo_rvect2[6]), .B(n_41640), .Z(n_30972
		));
	notech_reg ififo_rvect2_reg_7(.CP(n_61919), .D(n_30978), .CD(n_61358), .Q
		(ififo_rvect2[7]));
	notech_mux2 i_36283(.S(n_55049), .A(ififo_rvect2[7]), .B(n_41646), .Z(n_30978
		));
	notech_ao4 i_11626445(.A(n_57492), .B(n_39653), .C(n_58702), .D(n_40007)
		, .Z(n_267991526));
	notech_reg ififo_rvect1_reg_0(.CP(n_61917), .D(n_30984), .CD(n_61358), .Q
		(ififo_rvect1[0]));
	notech_mux2 i_36291(.S(n_55049), .A(ififo_rvect1[0]), .B(n_41822), .Z(n_30984
		));
	notech_reg ififo_rvect1_reg_1(.CP(n_61917), .D(n_30990), .CD(n_61358), .Q
		(ififo_rvect1[1]));
	notech_mux2 i_36299(.S(n_55049), .A(ififo_rvect1[1]), .B(n_41828), .Z(n_30990
		));
	notech_ao4 i_11726446(.A(n_57490), .B(n_39656), .C(n_58702), .D(n_40008)
		, .Z(n_267791524));
	notech_reg ififo_rvect1_reg_2(.CP(n_61917), .D(n_30996), .CD(n_61358), .Q
		(ififo_rvect1[2]));
	notech_mux2 i_36307(.S(n_55049), .A(ififo_rvect1[2]), .B(n_41834), .Z(n_30996
		));
	notech_reg ififo_rvect1_reg_3(.CP(n_61917), .D(n_31002), .CD(n_61358), .Q
		(ififo_rvect1[3]));
	notech_mux2 i_36315(.S(n_55049), .A(ififo_rvect1[3]), .B(n_41840), .Z(n_31002
		));
	notech_ao4 i_11926448(.A(n_57492), .B(n_39660), .C(n_58702), .D(n_40010)
		, .Z(n_267591522));
	notech_reg ififo_rvect1_reg_4(.CP(n_61917), .D(n_31008), .CD(n_61358), .Q
		(ififo_rvect1[4]));
	notech_mux2 i_36323(.S(n_55049), .A(ififo_rvect1[4]), .B(n_41846), .Z(n_31008
		));
	notech_reg ififo_rvect1_reg_5(.CP(n_61919), .D(n_31014), .CD(n_61358), .Q
		(ififo_rvect1[5]));
	notech_mux2 i_36331(.S(n_55049), .A(ififo_rvect1[5]), .B(n_41852), .Z(n_31014
		));
	notech_ao4 i_12126450(.A(n_57492), .B(n_39665), .C(n_58702), .D(n_40012)
		, .Z(n_267391520));
	notech_reg ififo_rvect1_reg_6(.CP(n_61919), .D(n_31020), .CD(n_61358), .Q
		(ififo_rvect1[6]));
	notech_mux2 i_36339(.S(n_55049), .A(ififo_rvect1[6]), .B(n_41858), .Z(n_31020
		));
	notech_reg ififo_rvect1_reg_7(.CP(n_61919), .D(n_31026), .CD(n_61358), .Q
		(ififo_rvect1[7]));
	notech_mux2 i_36347(.S(n_55049), .A(ififo_rvect1[7]), .B(n_41864), .Z(n_31026
		));
	notech_ao4 i_12226451(.A(n_57492), .B(n_39667), .C(n_58702), .D(n_40013)
		, .Z(n_267191518));
	notech_reg int_excl_reg_0(.CP(n_61917), .D(n_31032), .CD(n_61358), .Q(int_excl
		[0]));
	notech_mux2 i_36355(.S(\nbus_13566[0] ), .A(int_excl[0]), .B(n_171593336
		), .Z(n_31032));
	notech_reg int_excl_reg_1(.CP(n_61919), .D(n_31038), .CD(n_61356), .Q(int_excl
		[1]));
	notech_mux2 i_36363(.S(\nbus_13566[0] ), .A(int_excl[1]), .B(n_171693337
		), .Z(n_31038));
	notech_ao4 i_12326452(.A(n_57490), .B(n_39669), .C(n_58702), .D(n_40014)
		, .Z(n_266991516));
	notech_reg int_excl_reg_2(.CP(n_61922), .D(n_31044), .CD(n_61356), .Q(int_excl
		[2]));
	notech_mux2 i_36371(.S(\nbus_13566[0] ), .A(int_excl[2]), .B(n_49900), .Z
		(n_31044));
	notech_reg int_excl_reg_3(.CP(n_61922), .D(n_31050), .CD(n_61356), .Q(int_excl
		[3]));
	notech_mux2 i_36379(.S(\nbus_13566[0] ), .A(int_excl[3]), .B(n_171793338
		), .Z(n_31050));
	notech_ao4 i_12626455(.A(n_57490), .B(n_39672), .C(n_58702), .D(n_40017)
		, .Z(n_266791514));
	notech_reg int_excl_reg_4(.CP(n_61922), .D(n_31056), .CD(n_61358), .Q(int_excl
		[4]));
	notech_mux2 i_36387(.S(\nbus_13566[0] ), .A(int_excl[4]), .B(n_260991456
		), .Z(n_31056));
	notech_reg int_excl_reg_5(.CP(n_61922), .D(n_31062), .CD(n_61358), .Q(int_excl
		[5]));
	notech_mux2 i_36395(.S(\nbus_13566[0] ), .A(int_excl[5]), .B(n_161193232
		), .Z(n_31062));
	notech_ao4 i_13026459(.A(n_57490), .B(n_39678), .C(n_58702), .D(n_40021)
		, .Z(n_266591512));
	notech_reg fpu_reg(.CP(n_61922), .D(n_31068), .CD(n_61358), .Q(fpu));
	notech_mux2 i_36403(.S(n_3140), .A(n_171493335), .B(fpu), .Z(n_31068));
	notech_reg twobyte_reg(.CP(n_61922), .D(n_31074), .CD(n_61358), .Q(twobyte
		));
	notech_mux2 i_36411(.S(n_3141), .A(n_41571), .B(twobyte), .Z(n_31074));
	notech_ao4 i_13826467(.A(n_58702), .B(n_40029), .C(n_57490), .D(n_39694)
		, .Z(n_266391510));
	notech_reg opz_reg_0(.CP(n_61922), .D(n_31083), .CD(n_61358), .Q(opz[0])
		);
	notech_and4 i_36421(.A(n_59683), .B(n_2141), .C(n_18050174), .D(opz[0]),
		 .Z(n_31083));
	notech_reg opz_reg_1(.CP(n_61922), .D(n_31086), .CD(n_61361), .Q(opz[1])
		);
	notech_mux2 i_36427(.S(\nbus_13550[1] ), .A(opz[1]), .B(n_171393334), .Z
		(n_31086));
	notech_ao4 i_422121(.A(n_57490), .B(n_39831), .C(n_58702), .D(n_40190), 
		.Z(n_266191508));
	notech_reg_set opz_reg_2(.CP(n_61922), .D(n_31092), .SD(n_61361), .Q(opz
		[2]));
	notech_mux2 i_36435(.S(\nbus_13550[1] ), .A(opz[2]), .B(n_38647), .Z(n_31092
		));
	notech_reg imm_sz_reg_0(.CP(n_61922), .D(n_31098), .CD(n_61361), .Q(imm_sz
		[0]));
	notech_mux2 i_36443(.S(n_2091), .A(n_49816), .B(imm_sz[0]), .Z(n_31098)
		);
	notech_nand3 i_1425665(.A(n_59683), .B(n_265891505), .C(n_265791504), .Z
		(n_265991506));
	notech_reg imm_sz_reg_1(.CP(n_61922), .D(n_31104), .CD(n_61361), .Q(imm_sz
		[1]));
	notech_mux2 i_36451(.S(n_2091), .A(n_38649), .B(imm_sz[1]), .Z(n_31104)
		);
	notech_nao3 i_1386(.A(n_2847), .B(inst_deco1[13]), .C(n_1995), .Z(n_265891505
		));
	notech_reg imm_sz_reg_2(.CP(n_61919), .D(n_31110), .CD(n_61361), .Q(imm_sz
		[2]));
	notech_mux2 i_36459(.S(n_2091), .A(n_49828), .B(imm_sz[2]), .Z(n_31110)
		);
	notech_or4 i_1385(.A(n_58831), .B(pc_req), .C(pg_fault), .D(n_39875), .Z
		(n_265791504));
	notech_reg i_ptr_reg_0(.CP(n_61919), .D(n_31116), .CD(n_61361), .Q(i_ptr
		[0]));
	notech_mux2 i_36467(.S(n_2130), .A(n_38407), .B(i_ptr[0]), .Z(n_31116)
		);
	notech_nand3 i_323148(.A(n_265391500), .B(n_59596), .C(n_265591502), .Z(n_265691503
		));
	notech_reg i_ptr_reg_1(.CP(n_61919), .D(n_31122), .CD(n_61361), .Q(i_ptr
		[1]));
	notech_mux2 i_36475(.S(n_2130), .A(n_39303), .B(i_ptr[1]), .Z(n_31122)
		);
	notech_nand3 i_1383(.A(n_2124), .B(opz2[2]), .C(n_59596), .Z(n_265591502
		));
	notech_reg i_ptr_reg_2(.CP(n_61919), .D(n_31128), .CD(n_61361), .Q(i_ptr
		[2]));
	notech_mux2 i_36483(.S(n_2130), .A(n_41752), .B(i_ptr[2]), .Z(n_31128)
		);
	notech_nand2 i_204(.A(n_265391500), .B(n_59596), .Z(n_265491501));
	notech_reg i_ptr_reg_3(.CP(n_61919), .D(n_31137), .CD(n_61361), .Q(i_ptr
		[3]));
	notech_and2 i_36493(.A(n_2130), .B(i_ptr[3]), .Z(n_31137));
	notech_nao3 i_1381(.A(opz[2]), .B(n_59596), .C(n_58831), .Z(n_265391500)
		);
	notech_reg idx_deco_reg_0(.CP(n_61922), .D(n_31140), .CD(n_61361), .Q(idx_deco
		[0]));
	notech_mux2 i_36499(.S(n_3142), .A(n_41681), .B(idx_deco[0]), .Z(n_31140
		));
	notech_ao4 i_2027820(.A(n_57492), .B(n_38544), .C(n_2206), .D(n_58707), 
		.Z(n_265291499));
	notech_reg idx_deco_reg_1(.CP(n_61922), .D(n_31146), .CD(n_61361), .Q(idx_deco
		[1]));
	notech_mux2 i_36507(.S(n_3142), .A(n_41687), .B(idx_deco[1]), .Z(n_31146
		));
	notech_reg fsm_reg_0(.CP(n_61922), .D(n_31152), .CD(n_61361), .Q(fsm[0])
		);
	notech_mux2 i_36515(.S(n_3143), .A(n_38404), .B(fsm[0]), .Z(n_31152));
	notech_ao4 i_3027830(.A(n_1977), .B(n_58714), .C(n_57492), .D(n_38564), 
		.Z(n_265091497));
	notech_reg fsm_reg_1(.CP(n_61922), .D(n_31158), .CD(n_61361), .Q(fsm[1])
		);
	notech_mux2 i_36523(.S(n_3143), .A(n_38405), .B(fsm[1]), .Z(n_31158));
	notech_reg fsm_reg_2(.CP(n_61922), .D(n_31164), .CD(n_61361), .Q(fsm[2])
		);
	notech_mux2 i_36531(.S(n_3143), .A(n_38406), .B(fsm[2]), .Z(n_31164));
	notech_ao4 i_17026288(.A(n_58714), .B(n_40061), .C(n_57492), .D(n_39360)
		, .Z(n_264891495));
	notech_reg fsm_reg_3(.CP(n_61889), .D(n_31173), .CD(n_61358), .Q(fsm[3])
		);
	notech_and2 i_36541(.A(n_3143), .B(fsm[3]), .Z(n_31173));
	notech_reg fsm_reg_4(.CP(n_61889), .D(n_31179), .CD(n_61358), .Q(fsm[4])
		);
	notech_and2 i_36549(.A(n_3143), .B(fsm[4]), .Z(n_31179));
	notech_ao4 i_627218(.A(n_57492), .B(n_39120), .C(n_58714), .D(n_39118), 
		.Z(n_264691493));
	notech_reg repz_reg(.CP(n_61889), .D(n_31182), .CD(n_61361), .Q(repz));
	notech_mux2 i_36555(.S(n_43061), .A(repz), .B(n_171293333), .Z(n_31182)
		);
	notech_reg rep_reg(.CP(n_61889), .D(n_31188), .CD(n_61361), .Q(rep));
	notech_mux2 i_36563(.S(n_43061), .A(rep), .B(n_41571), .Z(n_31188));
	notech_ao4 i_12825523(.A(n_57492), .B(n_38871), .C(n_58714), .D(n_39989)
		, .Z(n_264491491));
	notech_reg reps2_reg_0(.CP(n_61889), .D(n_31194), .CD(n_61361), .Q(reps2
		[0]));
	notech_mux2 i_36571(.S(n_54244), .A(reps2[0]), .B(n_49757), .Z(n_31194)
		);
	notech_reg reps2_reg_1(.CP(n_61891), .D(n_31200), .CD(n_61361), .Q(reps2
		[1]));
	notech_mux2 i_36579(.S(n_54244), .A(reps2[1]), .B(n_49763), .Z(n_31200)
		);
	notech_ao4 i_123143(.A(n_57492), .B(n_38669), .C(n_39249), .D(n_40175), 
		.Z(n_264291489));
	notech_reg reps2_reg_2(.CP(n_61891), .D(n_31206), .CD(n_61361), .Q(reps2
		[2]));
	notech_mux2 i_36587(.S(n_54244), .A(reps2[2]), .B(n_49769), .Z(n_31206)
		);
	notech_reg reps1_reg_0(.CP(n_61891), .D(n_31212), .CD(n_61344), .Q(reps1
		[0]));
	notech_mux2 i_36595(.S(n_57666), .A(reps1[0]), .B(n_38401), .Z(n_31212)
		);
	notech_ao4 i_223144(.A(n_57492), .B(n_38671), .C(n_58714), .D(n_38666), 
		.Z(n_264091487));
	notech_reg reps1_reg_1(.CP(n_61889), .D(n_31218), .CD(n_61328), .Q(reps1
		[1]));
	notech_mux2 i_36603(.S(n_57666), .A(reps1[1]), .B(n_38402), .Z(n_31218)
		);
	notech_reg reps1_reg_2(.CP(n_61889), .D(n_31224), .CD(n_61328), .Q(reps1
		[2]));
	notech_mux2 i_36611(.S(n_57666), .A(reps1[2]), .B(n_38403), .Z(n_31224)
		);
	notech_ao4 i_323145(.A(n_57492), .B(n_38672), .C(n_38834), .D(n_38668), 
		.Z(n_263891485));
	notech_reg inst_deco2_reg_0(.CP(n_61889), .D(n_31230), .CD(n_61328), .Q(inst_deco2
		[0]));
	notech_mux2 i_36619(.S(n_54244), .A(inst_deco2[0]), .B(n_3443), .Z(n_31230
		));
	notech_reg inst_deco2_reg_1(.CP(n_61889), .D(n_31236), .CD(n_61328), .Q(inst_deco2
		[1]));
	notech_mux2 i_36627(.S(n_54244), .A(inst_deco2[1]), .B(n_3441), .Z(n_31236
		));
	notech_ao4 i_123110(.A(n_39117), .B(n_3134), .C(n_262891475), .D(n_39849
		), .Z(n_263691483));
	notech_reg inst_deco2_reg_2(.CP(n_61889), .D(n_31242), .CD(n_61328), .Q(inst_deco2
		[2]));
	notech_mux2 i_36635(.S(n_54222), .A(inst_deco2[2]), .B(n_3439), .Z(n_31242
		));
	notech_reg inst_deco2_reg_3(.CP(n_61889), .D(n_31248), .CD(n_61330), .Q(inst_deco2
		[3]));
	notech_mux2 i_36643(.S(n_54222), .A(inst_deco2[3]), .B(n_3437), .Z(n_31248
		));
	notech_ao4 i_223111(.A(n_39117), .B(n_263391480), .C(n_262891475), .D(n_39849
		), .Z(n_263491481));
	notech_reg inst_deco2_reg_4(.CP(n_61889), .D(n_31254), .CD(n_61330), .Q(inst_deco2
		[4]));
	notech_mux2 i_36651(.S(n_54222), .A(inst_deco2[4]), .B(n_3435), .Z(n_31254
		));
	notech_nor2 i_351(.A(ipg_fault), .B(n_263191478), .Z(n_263391480));
	notech_reg inst_deco2_reg_5(.CP(n_61889), .D(n_31260), .CD(n_61330), .Q(inst_deco2
		[5]));
	notech_mux2 i_36659(.S(n_54222), .A(inst_deco2[5]), .B(n_3433), .Z(n_31260
		));
	notech_reg inst_deco2_reg_6(.CP(n_61889), .D(n_31266), .CD(n_61328), .Q(inst_deco2
		[6]));
	notech_mux2 i_36667(.S(n_54222), .A(inst_deco2[6]), .B(n_3431), .Z(n_31266
		));
	notech_and2 i_1355(.A(n_1476), .B(n_2864), .Z(n_263191478));
	notech_reg inst_deco2_reg_7(.CP(n_61889), .D(n_31272), .CD(n_61330), .Q(inst_deco2
		[7]));
	notech_mux2 i_36675(.S(n_54222), .A(inst_deco2[7]), .B(n_3429), .Z(n_31272
		));
	notech_or2 i_349(.A(ipg_fault), .B(n_39117), .Z(n_263091477));
	notech_reg inst_deco2_reg_8(.CP(n_61889), .D(n_31278), .CD(n_61328), .Q(inst_deco2
		[8]));
	notech_mux2 i_36683(.S(n_54222), .A(inst_deco2[8]), .B(n_3427), .Z(n_31278
		));
	notech_nao3 i_350(.A(n_59602), .B(n_38661), .C(n_2834), .Z(n_262991476)
		);
	notech_reg inst_deco2_reg_9(.CP(n_61889), .D(n_31284), .CD(n_61328), .Q(inst_deco2
		[9]));
	notech_mux2 i_36691(.S(n_54227), .A(inst_deco2[9]), .B(n_3425), .Z(n_31284
		));
	notech_and3 i_1353(.A(n_58714), .B(n_263091477), .C(n_262991476), .Z(n_262891475
		));
	notech_reg inst_deco2_reg_10(.CP(n_61889), .D(n_31290), .CD(n_61328), .Q
		(inst_deco2[10]));
	notech_mux2 i_36699(.S(n_54227), .A(inst_deco2[10]), .B(n_3423), .Z(n_31290
		));
	notech_ao4 i_323112(.A(n_262691473), .B(n_2071), .C(n_2217), .D(n_2872),
		 .Z(n_262791474));
	notech_reg inst_deco2_reg_11(.CP(n_61891), .D(n_31296), .CD(n_61328), .Q
		(inst_deco2[11]));
	notech_mux2 i_36707(.S(n_54227), .A(inst_deco2[11]), .B(n_3421), .Z(n_31296
		));
	notech_ao4 i_348(.A(n_58712), .B(n_2844), .C(n_39117), .D(n_2845), .Z(n_262691473
		));
	notech_reg inst_deco2_reg_12(.CP(n_61891), .D(n_31302), .CD(n_61328), .Q
		(inst_deco2[12]));
	notech_mux2 i_36715(.S(n_54222), .A(inst_deco2[12]), .B(n_3419), .Z(n_31302
		));
	notech_reg inst_deco2_reg_13(.CP(n_61891), .D(n_31308), .CD(n_61328), .Q
		(inst_deco2[13]));
	notech_mux2 i_36723(.S(n_54227), .A(inst_deco2[13]), .B(n_3417), .Z(n_31308
		));
	notech_reg inst_deco2_reg_14(.CP(n_61891), .D(n_31314), .CD(n_61328), .Q
		(inst_deco2[14]));
	notech_mux2 i_36731(.S(n_54227), .A(inst_deco2[14]), .B(n_3415), .Z(n_31314
		));
	notech_reg inst_deco2_reg_15(.CP(n_61891), .D(n_31320), .CD(n_61328), .Q
		(inst_deco2[15]));
	notech_mux2 i_36739(.S(n_54222), .A(inst_deco2[15]), .B(n_3413), .Z(n_31320
		));
	notech_reg inst_deco2_reg_16(.CP(n_61895), .D(n_31326), .CD(n_61328), .Q
		(inst_deco2[16]));
	notech_mux2 i_36747(.S(n_54222), .A(inst_deco2[16]), .B(n_3411), .Z(n_31326
		));
	notech_and4 i_123227(.A(n_3130), .B(n_251091357), .C(n_250991356), .D(n_262091467
		), .Z(n_262191468));
	notech_reg inst_deco2_reg_17(.CP(n_61895), .D(n_31332), .CD(n_61328), .Q
		(inst_deco2[17]));
	notech_mux2 i_36755(.S(n_54222), .A(inst_deco2[17]), .B(n_3409), .Z(n_31332
		));
	notech_nand2 i_1335(.A(fpu), .B(n_39853), .Z(n_262091467));
	notech_reg inst_deco2_reg_18(.CP(n_61895), .D(n_31338), .CD(n_61328), .Q
		(inst_deco2[18]));
	notech_mux2 i_36763(.S(n_54221), .A(inst_deco2[18]), .B(n_3407), .Z(n_31338
		));
	notech_reg inst_deco2_reg_19(.CP(n_61891), .D(n_31344), .CD(n_61330), .Q
		(inst_deco2[19]));
	notech_mux2 i_36771(.S(n_54221), .A(inst_deco2[19]), .B(n_3405), .Z(n_31344
		));
	notech_reg inst_deco2_reg_20(.CP(n_61895), .D(n_31350), .CD(n_61334), .Q
		(inst_deco2[20]));
	notech_mux2 i_36779(.S(n_54221), .A(inst_deco2[20]), .B(n_3403), .Z(n_31350
		));
	notech_ao4 i_343(.A(n_3128), .B(n_3120), .C(n_250891355), .D(n_261391460
		), .Z(n_261791464));
	notech_reg inst_deco2_reg_21(.CP(n_61891), .D(n_31356), .CD(n_61330), .Q
		(inst_deco2[21]));
	notech_mux2 i_36787(.S(n_54222), .A(inst_deco2[21]), .B(n_3401), .Z(n_31356
		));
	notech_nor2 i_344(.A(n_2867), .B(n_261191458), .Z(n_261691463));
	notech_reg inst_deco2_reg_22(.CP(n_61891), .D(n_31362), .CD(n_61330), .Q
		(inst_deco2[22]));
	notech_mux2 i_36795(.S(n_54222), .A(inst_deco2[22]), .B(n_3399), .Z(n_31362
		));
	notech_and2 i_345(.A(n_2073), .B(n_261091457), .Z(n_261591462));
	notech_reg inst_deco2_reg_23(.CP(n_61891), .D(n_31368), .CD(n_61330), .Q
		(inst_deco2[23]));
	notech_mux2 i_36803(.S(n_54222), .A(inst_deco2[23]), .B(n_3397), .Z(n_31368
		));
	notech_reg inst_deco2_reg_24(.CP(n_61891), .D(n_31374), .CD(n_61334), .Q
		(inst_deco2[24]));
	notech_mux2 i_36811(.S(n_54222), .A(inst_deco2[24]), .B(n_3395), .Z(n_31374
		));
	notech_nor2 i_346(.A(n_2074), .B(\to_acu2_0[3] ), .Z(n_261391460));
	notech_reg inst_deco2_reg_25(.CP(n_61891), .D(n_31380), .CD(n_61334), .Q
		(inst_deco2[25]));
	notech_mux2 i_36819(.S(n_54222), .A(inst_deco2[25]), .B(n_3393), .Z(n_31380
		));
	notech_reg inst_deco2_reg_26(.CP(n_61891), .D(n_31386), .CD(n_61334), .Q
		(inst_deco2[26]));
	notech_mux2 i_36827(.S(n_54222), .A(inst_deco2[26]), .B(n_3391), .Z(n_31386
		));
	notech_ao3 i_1329(.A(n_2864), .B(n_251191358), .C(fpu), .Z(n_261191458)
		);
	notech_reg inst_deco2_reg_27(.CP(n_61891), .D(n_31392), .CD(n_61334), .Q
		(inst_deco2[27]));
	notech_mux2 i_36835(.S(n_54222), .A(inst_deco2[27]), .B(n_3389), .Z(n_31392
		));
	notech_or4 i_1327(.A(n_5717), .B(n_251191358), .C(n_38508), .D(n_40209),
		 .Z(n_261091457));
	notech_reg inst_deco2_reg_28(.CP(n_61891), .D(n_31398), .CD(n_61334), .Q
		(inst_deco2[28]));
	notech_mux2 i_36843(.S(n_54227), .A(inst_deco2[28]), .B(n_3387), .Z(n_31398
		));
	notech_nao3 i_527193(.A(n_260791454), .B(n_260891455), .C(n_5392), .Z(n_260991456
		));
	notech_reg inst_deco2_reg_29(.CP(n_61891), .D(n_31404), .CD(n_61330), .Q
		(inst_deco2[29]));
	notech_mux2 i_36851(.S(n_54232), .A(inst_deco2[29]), .B(n_3385), .Z(n_31404
		));
	notech_nand2 i_1275(.A(int_excl[4]), .B(n_1820), .Z(n_260891455));
	notech_reg inst_deco2_reg_30(.CP(n_61891), .D(n_31410), .CD(n_61330), .Q
		(inst_deco2[30]));
	notech_mux2 i_36859(.S(n_54232), .A(inst_deco2[30]), .B(n_3383), .Z(n_31410
		));
	notech_or2 i_169(.A(int_excl[4]), .B(n_1820), .Z(n_260791454));
	notech_reg inst_deco2_reg_31(.CP(n_61891), .D(n_31416), .CD(n_61330), .Q
		(inst_deco2[31]));
	notech_mux2 i_36867(.S(n_54232), .A(inst_deco2[31]), .B(n_3381), .Z(n_31416
		));
	notech_ao4 i_127737(.A(n_57492), .B(n_38456), .C(n_2225), .D(n_58714), .Z
		(n_260691453));
	notech_reg inst_deco2_reg_32(.CP(n_61889), .D(n_31422), .CD(n_61330), .Q
		(inst_deco2[32]));
	notech_mux2 i_36875(.S(n_54232), .A(inst_deco2[32]), .B(n_3379), .Z(n_31422
		));
	notech_reg inst_deco2_reg_33(.CP(n_61884), .D(n_31428), .CD(n_61330), .Q
		(inst_deco2[33]));
	notech_mux2 i_36883(.S(n_54232), .A(inst_deco2[33]), .B(n_3377), .Z(n_31428
		));
	notech_ao4 i_227738(.A(n_57492), .B(n_38458), .C(n_223393386), .D(n_58714
		), .Z(n_260491451));
	notech_reg inst_deco2_reg_34(.CP(n_61884), .D(n_31434), .CD(n_61330), .Q
		(inst_deco2[34]));
	notech_mux2 i_36891(.S(n_54232), .A(inst_deco2[34]), .B(n_3375), .Z(n_31434
		));
	notech_reg inst_deco2_reg_35(.CP(n_61884), .D(n_31440), .CD(n_61330), .Q
		(inst_deco2[35]));
	notech_mux2 i_36899(.S(n_54232), .A(inst_deco2[35]), .B(n_3373), .Z(n_31440
		));
	notech_ao4 i_327739(.A(n_57504), .B(n_38460), .C(n_224193378), .D(n_58714
		), .Z(n_260291449));
	notech_reg inst_deco2_reg_36(.CP(n_61884), .D(n_31446), .CD(n_61330), .Q
		(inst_deco2[36]));
	notech_mux2 i_36907(.S(n_54232), .A(inst_deco2[36]), .B(n_3371), .Z(n_31446
		));
	notech_reg inst_deco2_reg_37(.CP(n_61884), .D(n_31452), .CD(n_61330), .Q
		(inst_deco2[37]));
	notech_mux2 i_36915(.S(n_54233), .A(inst_deco2[37]), .B(n_3369), .Z(n_31452
		));
	notech_ao4 i_427740(.A(n_57504), .B(n_38462), .C(n_224993370), .D(n_58717
		), .Z(n_260091447));
	notech_reg inst_deco2_reg_38(.CP(n_61884), .D(n_31458), .CD(n_61330), .Q
		(inst_deco2[38]));
	notech_mux2 i_36923(.S(n_54233), .A(inst_deco2[38]), .B(n_3367), .Z(n_31458
		));
	notech_reg inst_deco2_reg_39(.CP(n_61884), .D(n_31464), .CD(n_61330), .Q
		(inst_deco2[39]));
	notech_mux2 i_36931(.S(n_54232), .A(inst_deco2[39]), .B(n_3365), .Z(n_31464
		));
	notech_ao4 i_527741(.A(n_57504), .B(n_38464), .C(n_225793362), .D(n_58717
		), .Z(n_259891445));
	notech_reg inst_deco2_reg_40(.CP(n_61884), .D(n_31470), .CD(n_61323), .Q
		(inst_deco2[40]));
	notech_mux2 i_36939(.S(n_54232), .A(inst_deco2[40]), .B(n_3363), .Z(n_31470
		));
	notech_reg inst_deco2_reg_41(.CP(n_61884), .D(n_31476), .CD(n_61323), .Q
		(inst_deco2[41]));
	notech_mux2 i_36947(.S(n_54232), .A(inst_deco2[41]), .B(n_3361), .Z(n_31476
		));
	notech_ao4 i_627742(.A(n_57504), .B(n_38465), .C(n_226593354), .D(n_58717
		), .Z(n_259691443));
	notech_reg inst_deco2_reg_42(.CP(n_61884), .D(n_31482), .CD(n_61323), .Q
		(inst_deco2[42]));
	notech_mux2 i_36955(.S(n_54227), .A(inst_deco2[42]), .B(n_3359), .Z(n_31482
		));
	notech_reg inst_deco2_reg_43(.CP(n_61884), .D(n_31488), .CD(n_61323), .Q
		(inst_deco2[43]));
	notech_mux2 i_36963(.S(n_54227), .A(inst_deco2[43]), .B(n_3357), .Z(n_31488
		));
	notech_ao4 i_727743(.A(n_57504), .B(n_38466), .C(n_227393346), .D(n_58717
		), .Z(n_259491441));
	notech_reg inst_deco2_reg_44(.CP(n_61884), .D(n_31494), .CD(n_61323), .Q
		(inst_deco2[44]));
	notech_mux2 i_36971(.S(n_54227), .A(inst_deco2[44]), .B(n_3355), .Z(n_31494
		));
	notech_reg inst_deco2_reg_45(.CP(n_61884), .D(n_31500), .CD(n_61323), .Q
		(inst_deco2[45]));
	notech_mux2 i_36979(.S(n_54227), .A(inst_deco2[45]), .B(n_3353), .Z(n_31500
		));
	notech_ao4 i_827744(.A(n_57504), .B(n_38467), .C(n_228191128), .D(n_58717
		), .Z(n_259291439));
	notech_reg inst_deco2_reg_46(.CP(n_61884), .D(n_31506), .CD(n_61323), .Q
		(inst_deco2[46]));
	notech_mux2 i_36987(.S(n_54227), .A(inst_deco2[46]), .B(n_3351), .Z(n_31506
		));
	notech_reg inst_deco2_reg_47(.CP(n_61881), .D(n_31512), .CD(n_61323), .Q
		(inst_deco2[47]));
	notech_mux2 i_36995(.S(n_54227), .A(inst_deco2[47]), .B(n_3349), .Z(n_31512
		));
	notech_ao4 i_927745(.A(n_57504), .B(n_38468), .C(n_228991136), .D(n_58714
		), .Z(n_259091437));
	notech_reg inst_deco2_reg_48(.CP(n_61881), .D(n_31518), .CD(n_61323), .Q
		(inst_deco2[48]));
	notech_mux2 i_37003(.S(n_54232), .A(inst_deco2[48]), .B(n_3347), .Z(n_31518
		));
	notech_reg inst_deco2_reg_49(.CP(n_61884), .D(n_31524), .CD(n_61323), .Q
		(inst_deco2[49]));
	notech_mux2 i_37011(.S(n_54232), .A(inst_deco2[49]), .B(n_3345), .Z(n_31524
		));
	notech_ao4 i_1027746(.A(n_57504), .B(n_38469), .C(n_229791144), .D(n_58714
		), .Z(n_258891435));
	notech_reg inst_deco2_reg_50(.CP(n_61884), .D(n_31530), .CD(n_61323), .Q
		(inst_deco2[50]));
	notech_mux2 i_37019(.S(n_54232), .A(inst_deco2[50]), .B(n_3343), .Z(n_31530
		));
	notech_reg inst_deco2_reg_51(.CP(n_61884), .D(n_31536), .CD(n_61320), .Q
		(inst_deco2[51]));
	notech_mux2 i_37027(.S(n_54232), .A(inst_deco2[51]), .B(n_3341), .Z(n_31536
		));
	notech_ao4 i_1127747(.A(n_57504), .B(n_38470), .C(n_230591152), .D(n_58714
		), .Z(n_258691433));
	notech_reg inst_deco2_reg_52(.CP(n_61884), .D(n_31542), .CD(n_61320), .Q
		(inst_deco2[52]));
	notech_mux2 i_37035(.S(n_54232), .A(inst_deco2[52]), .B(n_3339), .Z(n_31542
		));
	notech_reg inst_deco2_reg_53(.CP(n_61884), .D(n_31548), .CD(n_61320), .Q
		(inst_deco2[53]));
	notech_mux2 i_37043(.S(n_54232), .A(inst_deco2[53]), .B(n_3337), .Z(n_31548
		));
	notech_ao4 i_1227748(.A(n_57504), .B(n_38471), .C(n_231391160), .D(n_58714
		), .Z(n_258491431));
	notech_reg inst_deco2_reg_54(.CP(n_61886), .D(n_31554), .CD(n_61320), .Q
		(inst_deco2[54]));
	notech_mux2 i_37051(.S(n_54232), .A(inst_deco2[54]), .B(n_3335), .Z(n_31554
		));
	notech_reg inst_deco2_reg_55(.CP(n_61886), .D(n_31560), .CD(n_61320), .Q
		(inst_deco2[55]));
	notech_mux2 i_37059(.S(n_54245), .A(inst_deco2[55]), .B(n_3333), .Z(n_31560
		));
	notech_ao4 i_1327749(.A(n_57507), .B(n_38472), .C(n_232191168), .D(n_58714
		), .Z(n_258291429));
	notech_reg inst_deco2_reg_56(.CP(n_61886), .D(n_31566), .CD(n_61323), .Q
		(inst_deco2[56]));
	notech_mux2 i_37067(.S(n_54261), .A(inst_deco2[56]), .B(n_3331), .Z(n_31566
		));
	notech_reg inst_deco2_reg_57(.CP(n_61886), .D(n_31572), .CD(n_61323), .Q
		(inst_deco2[57]));
	notech_mux2 i_37075(.S(n_54266), .A(inst_deco2[57]), .B(n_3329), .Z(n_31572
		));
	notech_ao4 i_1427750(.A(n_57507), .B(n_38473), .C(n_232991176), .D(n_58712
		), .Z(n_258091427));
	notech_reg inst_deco2_reg_58(.CP(n_61886), .D(n_31578), .CD(n_61323), .Q
		(inst_deco2[58]));
	notech_mux2 i_37083(.S(n_54266), .A(inst_deco2[58]), .B(n_3327), .Z(n_31578
		));
	notech_reg inst_deco2_reg_59(.CP(n_61886), .D(n_31584), .CD(n_61323), .Q
		(inst_deco2[59]));
	notech_mux2 i_37091(.S(n_54261), .A(inst_deco2[59]), .B(n_3325), .Z(n_31584
		));
	notech_ao4 i_1527751(.A(n_57507), .B(n_38474), .C(n_233791184), .D(n_58707
		), .Z(n_257891425));
	notech_reg inst_deco2_reg_60(.CP(n_61889), .D(n_31590), .CD(n_61323), .Q
		(inst_deco2[60]));
	notech_mux2 i_37099(.S(n_54261), .A(inst_deco2[60]), .B(n_3323), .Z(n_31590
		));
	notech_reg inst_deco2_reg_61(.CP(n_61886), .D(n_31596), .CD(n_61325), .Q
		(inst_deco2[61]));
	notech_mux2 i_37107(.S(n_54261), .A(inst_deco2[61]), .B(n_3321), .Z(n_31596
		));
	notech_ao4 i_1627752(.A(n_57507), .B(n_38475), .C(n_2163), .D(n_58707), 
		.Z(n_257691423));
	notech_reg inst_deco2_reg_62(.CP(n_61886), .D(n_31602), .CD(n_61325), .Q
		(inst_deco2[62]));
	notech_mux2 i_37115(.S(n_54266), .A(inst_deco2[62]), .B(n_42534), .Z(n_31602
		));
	notech_reg inst_deco2_reg_63(.CP(n_61886), .D(n_31608), .CD(n_61325), .Q
		(inst_deco2[63]));
	notech_mux2 i_37123(.S(n_54266), .A(inst_deco2[63]), .B(n_42540), .Z(n_31608
		));
	notech_ao4 i_1727753(.A(n_57507), .B(n_38476), .C(n_2176), .D(n_58707), 
		.Z(n_257491421));
	notech_reg inst_deco2_reg_64(.CP(n_61886), .D(n_31614), .CD(n_61325), .Q
		(inst_deco2[64]));
	notech_mux2 i_37131(.S(n_54266), .A(inst_deco2[64]), .B(n_3317), .Z(n_31614
		));
	notech_reg inst_deco2_reg_65(.CP(n_61886), .D(n_31620), .CD(n_61325), .Q
		(inst_deco2[65]));
	notech_mux2 i_37139(.S(n_54266), .A(inst_deco2[65]), .B(n_42552), .Z(n_31620
		));
	notech_ao4 i_1827754(.A(n_57504), .B(n_38477), .C(n_2186), .D(n_58712), 
		.Z(n_257291419));
	notech_reg inst_deco2_reg_66(.CP(n_61886), .D(n_31626), .CD(n_61325), .Q
		(inst_deco2[66]));
	notech_mux2 i_37147(.S(n_54266), .A(inst_deco2[66]), .B(n_42558), .Z(n_31626
		));
	notech_reg inst_deco2_reg_67(.CP(n_61886), .D(n_31632), .CD(n_61328), .Q
		(inst_deco2[67]));
	notech_mux2 i_37155(.S(n_54266), .A(inst_deco2[67]), .B(n_3313), .Z(n_31632
		));
	notech_ao4 i_1927755(.A(n_57504), .B(n_38478), .C(n_2196), .D(n_58712), 
		.Z(n_257091417));
	notech_reg inst_deco2_reg_68(.CP(n_61886), .D(n_31638), .CD(n_61325), .Q
		(inst_deco2[68]));
	notech_mux2 i_37163(.S(n_54266), .A(inst_deco2[68]), .B(n_42570), .Z(n_31638
		));
	notech_reg inst_deco2_reg_69(.CP(n_61886), .D(n_31644), .CD(n_61325), .Q
		(inst_deco2[69]));
	notech_mux2 i_37171(.S(n_54256), .A(inst_deco2[69]), .B(n_42576), .Z(n_31644
		));
	notech_ao4 i_2027756(.A(n_57504), .B(n_38479), .C(n_2206), .D(n_58707), 
		.Z(n_256891415));
	notech_reg inst_deco2_reg_70(.CP(n_61886), .D(n_31650), .CD(n_61325), .Q
		(inst_deco2[70]));
	notech_mux2 i_37179(.S(n_54256), .A(inst_deco2[70]), .B(n_42582), .Z(n_31650
		));
	notech_reg inst_deco2_reg_71(.CP(n_61886), .D(n_31656), .CD(n_61325), .Q
		(inst_deco2[71]));
	notech_mux2 i_37187(.S(n_54261), .A(inst_deco2[71]), .B(n_42588), .Z(n_31656
		));
	notech_ao4 i_2127757(.A(n_57507), .B(n_38480), .C(n_234891195), .D(n_58707
		), .Z(n_256691413));
	notech_reg inst_deco2_reg_72(.CP(n_61886), .D(n_31662), .CD(n_61325), .Q
		(inst_deco2[72]));
	notech_mux2 i_37195(.S(n_54256), .A(inst_deco2[72]), .B(n_3307), .Z(n_31662
		));
	notech_reg inst_deco2_reg_73(.CP(n_61886), .D(n_31668), .CD(n_61325), .Q
		(inst_deco2[73]));
	notech_mux2 i_37203(.S(n_54256), .A(inst_deco2[73]), .B(n_42600), .Z(n_31668
		));
	notech_ao4 i_2227758(.A(n_57504), .B(n_38481), .C(n_235891205), .D(n_58707
		), .Z(n_256491411));
	notech_reg inst_deco2_reg_74(.CP(n_61886), .D(n_31674), .CD(n_61325), .Q
		(inst_deco2[74]));
	notech_mux2 i_37211(.S(n_54256), .A(inst_deco2[74]), .B(n_3304), .Z(n_31674
		));
	notech_reg inst_deco2_reg_75(.CP(n_61902), .D(n_31680), .CD(n_61323), .Q
		(inst_deco2[75]));
	notech_mux2 i_37219(.S(n_54261), .A(inst_deco2[75]), .B(n_42612), .Z(n_31680
		));
	notech_ao4 i_2327759(.A(n_57502), .B(n_38482), .C(n_236891215), .D(n_58707
		), .Z(n_256291409));
	notech_reg inst_deco2_reg_76(.CP(n_61902), .D(n_31686), .CD(n_61323), .Q
		(inst_deco2[76]));
	notech_mux2 i_37227(.S(n_54261), .A(inst_deco2[76]), .B(n_42618), .Z(n_31686
		));
	notech_reg inst_deco2_reg_77(.CP(n_61902), .D(n_31692), .CD(n_61325), .Q
		(inst_deco2[77]));
	notech_mux2 i_37235(.S(n_54261), .A(inst_deco2[77]), .B(n_42624), .Z(n_31692
		));
	notech_ao4 i_2427760(.A(n_57497), .B(n_38483), .C(n_237891225), .D(n_58707
		), .Z(n_256091407));
	notech_reg inst_deco2_reg_78(.CP(n_61900), .D(n_31698), .CD(n_61325), .Q
		(inst_deco2[78]));
	notech_mux2 i_37243(.S(n_54261), .A(inst_deco2[78]), .B(n_42630), .Z(n_31698
		));
	notech_reg inst_deco2_reg_79(.CP(n_61900), .D(n_31704), .CD(n_61325), .Q
		(inst_deco2[79]));
	notech_mux2 i_37251(.S(n_54261), .A(inst_deco2[79]), .B(n_42636), .Z(n_31704
		));
	notech_ao4 i_2527761(.A(n_57497), .B(n_38484), .C(n_238991236), .D(n_58712
		), .Z(n_255891405));
	notech_reg inst_deco2_reg_80(.CP(n_61902), .D(n_31710), .CD(n_61325), .Q
		(inst_deco2[80]));
	notech_mux2 i_37259(.S(n_54261), .A(inst_deco2[80]), .B(n_42642), .Z(n_31710
		));
	notech_reg inst_deco2_reg_81(.CP(n_61902), .D(n_31716), .CD(n_61325), .Q
		(inst_deco2[81]));
	notech_mux2 i_37267(.S(n_54261), .A(inst_deco2[81]), .B(n_42648), .Z(n_31716
		));
	notech_ao4 i_2627762(.A(n_57502), .B(n_38485), .C(n_239991246), .D(n_58712
		), .Z(n_255691403));
	notech_reg inst_deco2_reg_82(.CP(n_61902), .D(n_31722), .CD(n_61334), .Q
		(inst_deco2[82]));
	notech_mux2 i_37275(.S(n_54266), .A(inst_deco2[82]), .B(n_42654), .Z(n_31722
		));
	notech_reg inst_deco2_reg_83(.CP(n_61902), .D(n_31728), .CD(n_61341), .Q
		(inst_deco2[83]));
	notech_mux2 i_37283(.S(n_54267), .A(inst_deco2[83]), .B(n_42660), .Z(n_31728
		));
	notech_ao4 i_2727763(.A(n_57502), .B(n_38486), .C(n_240991256), .D(n_58712
		), .Z(n_255491401));
	notech_reg inst_deco2_reg_84(.CP(n_61902), .D(n_31734), .CD(n_61341), .Q
		(inst_deco2[84]));
	notech_mux2 i_37291(.S(n_54267), .A(inst_deco2[84]), .B(n_42666), .Z(n_31734
		));
	notech_reg inst_deco2_reg_85(.CP(n_61900), .D(n_31740), .CD(n_61341), .Q
		(inst_deco2[85]));
	notech_mux2 i_37299(.S(n_54267), .A(inst_deco2[85]), .B(n_42672), .Z(n_31740
		));
	notech_ao4 i_2827764(.A(n_57502), .B(n_38487), .C(n_241991266), .D(n_58712
		), .Z(n_255291399));
	notech_reg inst_deco2_reg_86(.CP(n_61900), .D(n_31746), .CD(n_61341), .Q
		(inst_deco2[86]));
	notech_mux2 i_37307(.S(n_54267), .A(inst_deco2[86]), .B(n_42678), .Z(n_31746
		));
	notech_reg inst_deco2_reg_87(.CP(n_61900), .D(n_31752), .CD(n_61341), .Q
		(inst_deco2[87]));
	notech_mux2 i_37315(.S(n_54267), .A(inst_deco2[87]), .B(n_42684), .Z(n_31752
		));
	notech_ao4 i_2927765(.A(n_57497), .B(n_38488), .C(n_242991276), .D(n_58712
		), .Z(n_255091397));
	notech_reg inst_deco2_reg_88(.CP(n_61900), .D(n_31758), .CD(n_61341), .Q
		(inst_deco2[88]));
	notech_mux2 i_37323(.S(n_54267), .A(inst_deco2[88]), .B(n_42690), .Z(n_31758
		));
	notech_reg inst_deco2_reg_89(.CP(n_61900), .D(n_31764), .CD(n_61341), .Q
		(inst_deco2[89]));
	notech_mux2 i_37331(.S(n_54267), .A(inst_deco2[89]), .B(n_42696), .Z(n_31764
		));
	notech_ao4 i_3027766(.A(n_1977), .B(n_58712), .C(n_57497), .D(n_38489), 
		.Z(n_254891395));
	notech_reg inst_deco2_reg_90(.CP(n_61900), .D(n_31770), .CD(n_61341), .Q
		(inst_deco2[90]));
	notech_mux2 i_37339(.S(n_54267), .A(inst_deco2[90]), .B(n_42702), .Z(n_31770
		));
	notech_reg inst_deco2_reg_91(.CP(n_61900), .D(n_31776), .CD(n_61341), .Q
		(inst_deco2[91]));
	notech_mux2 i_37347(.S(n_54267), .A(inst_deco2[91]), .B(n_42708), .Z(n_31776
		));
	notech_ao4 i_3127767(.A(n_57497), .B(n_38490), .C(n_243991286), .D(n_58712
		), .Z(n_254691393));
	notech_reg inst_deco2_reg_92(.CP(n_61900), .D(n_31782), .CD(n_61341), .Q
		(inst_deco2[92]));
	notech_mux2 i_37355(.S(n_54267), .A(inst_deco2[92]), .B(n_42714), .Z(n_31782
		));
	notech_reg inst_deco2_reg_93(.CP(n_61900), .D(n_31788), .CD(n_61339), .Q
		(inst_deco2[93]));
	notech_mux2 i_37363(.S(n_54267), .A(inst_deco2[93]), .B(n_42720), .Z(n_31788
		));
	notech_ao4 i_3227768(.A(n_57497), .B(n_38491), .C(n_245091297), .D(n_58712
		), .Z(n_254491391));
	notech_reg inst_deco2_reg_94(.CP(n_61900), .D(n_31794), .CD(n_61339), .Q
		(inst_deco2[94]));
	notech_mux2 i_37371(.S(n_54267), .A(inst_deco2[94]), .B(n_42726), .Z(n_31794
		));
	notech_reg inst_deco2_reg_95(.CP(n_61900), .D(n_31800), .CD(n_61339), .Q
		(inst_deco2[95]));
	notech_mux2 i_37379(.S(n_54267), .A(inst_deco2[95]), .B(n_42732), .Z(n_31800
		));
	notech_ao4 i_3327769(.A(n_57497), .B(n_38492), .C(n_53727), .D(n_39661),
		 .Z(n_254291389));
	notech_reg inst_deco2_reg_96(.CP(n_61905), .D(n_31806), .CD(n_61339), .Q
		(inst_deco2[96]));
	notech_mux2 i_37387(.S(n_54266), .A(inst_deco2[96]), .B(n_42738), .Z(n_31806
		));
	notech_reg inst_deco2_reg_97(.CP(n_61905), .D(n_31812), .CD(n_61339), .Q
		(inst_deco2[97]));
	notech_mux2 i_37395(.S(n_54266), .A(inst_deco2[97]), .B(n_42744), .Z(n_31812
		));
	notech_ao4 i_3427770(.A(n_57502), .B(n_38493), .C(n_53727), .D(n_39654),
		 .Z(n_254091387));
	notech_reg inst_deco2_reg_98(.CP(n_61905), .D(n_31818), .CD(n_61339), .Q
		(inst_deco2[98]));
	notech_mux2 i_37403(.S(n_54266), .A(inst_deco2[98]), .B(n_42750), .Z(n_31818
		));
	notech_reg inst_deco2_reg_99(.CP(n_61902), .D(n_31824), .CD(n_61339), .Q
		(inst_deco2[99]));
	notech_mux2 i_37411(.S(n_54266), .A(inst_deco2[99]), .B(n_42756), .Z(n_31824
		));
	notech_ao4 i_3527771(.A(n_57502), .B(n_38494), .C(n_53727), .D(n_39647),
		 .Z(n_253891385));
	notech_reg inst_deco2_reg_100(.CP(n_61905), .D(n_31830), .CD(n_61339), .Q
		(inst_deco2[100]));
	notech_mux2 i_37419(.S(n_54266), .A(inst_deco2[100]), .B(n_42762), .Z(n_31830
		));
	notech_reg inst_deco2_reg_101(.CP(n_61905), .D(n_31836), .CD(n_61339), .Q
		(inst_deco2[101]));
	notech_mux2 i_37427(.S(n_54266), .A(inst_deco2[101]), .B(n_42768), .Z(n_31836
		));
	notech_ao4 i_3627772(.A(n_57502), .B(n_38495), .C(n_53727), .D(n_39643),
		 .Z(n_253691383));
	notech_reg inst_deco2_reg_102(.CP(n_61905), .D(n_31842), .CD(n_61339), .Q
		(inst_deco2[102]));
	notech_mux2 i_37435(.S(n_54266), .A(inst_deco2[102]), .B(n_42774), .Z(n_31842
		));
	notech_reg inst_deco2_reg_103(.CP(n_61905), .D(n_31848), .CD(n_61339), .Q
		(inst_deco2[103]));
	notech_mux2 i_37443(.S(n_54267), .A(inst_deco2[103]), .B(n_42780), .Z(n_31848
		));
	notech_ao4 i_3727773(.A(n_57502), .B(n_38496), .C(n_53727), .D(n_39636),
		 .Z(n_253491381));
	notech_reg inst_deco2_reg_104(.CP(n_61905), .D(n_31854), .CD(n_61344), .Q
		(inst_deco2[104]));
	notech_mux2 i_37451(.S(n_54267), .A(inst_deco2[104]), .B(n_42786), .Z(n_31854
		));
	notech_reg inst_deco2_reg_105(.CP(n_61905), .D(n_31860), .CD(n_61344), .Q
		(inst_deco2[105]));
	notech_mux2 i_37459(.S(n_54267), .A(inst_deco2[105]), .B(n_42792), .Z(n_31860
		));
	notech_ao4 i_4227778(.A(n_57502), .B(n_38501), .C(n_53788), .D(n_39612),
		 .Z(n_253291379));
	notech_reg inst_deco2_reg_106(.CP(n_61902), .D(n_31866), .CD(n_61344), .Q
		(inst_deco2[106]));
	notech_mux2 i_37467(.S(n_54266), .A(inst_deco2[106]), .B(n_42798), .Z(n_31866
		));
	notech_reg inst_deco2_reg_107(.CP(n_61902), .D(n_31872), .CD(n_61344), .Q
		(inst_deco2[107]));
	notech_mux2 i_37475(.S(n_54267), .A(inst_deco2[107]), .B(n_42804), .Z(n_31872
		));
	notech_ao4 i_4327779(.A(n_57502), .B(n_38502), .C(n_53788), .D(n_39610),
		 .Z(n_253091377));
	notech_reg inst_deco2_reg_108(.CP(n_61902), .D(n_31878), .CD(n_61344), .Q
		(inst_deco2[108]));
	notech_mux2 i_37483(.S(n_54267), .A(inst_deco2[108]), .B(n_42810), .Z(n_31878
		));
	notech_reg inst_deco2_reg_109(.CP(n_61902), .D(n_31884), .CD(n_61344), .Q
		(inst_deco2[109]));
	notech_mux2 i_37491(.S(n_54250), .A(inst_deco2[109]), .B(n_42816), .Z(n_31884
		));
	notech_ao4 i_4427780(.A(n_57502), .B(n_38503), .C(n_53788), .D(n_39607),
		 .Z(n_252891375));
	notech_reg inst_deco2_reg_110(.CP(n_61902), .D(n_31890), .CD(n_61344), .Q
		(inst_deco2[110]));
	notech_mux2 i_37499(.S(n_54250), .A(inst_deco2[110]), .B(n_42822), .Z(n_31890
		));
	notech_reg inst_deco2_reg_111(.CP(n_61902), .D(n_31896), .CD(n_61344), .Q
		(inst_deco2[111]));
	notech_mux2 i_37507(.S(n_54250), .A(inst_deco2[111]), .B(n_42828), .Z(n_31896
		));
	notech_ao4 i_4627782(.A(n_57502), .B(n_38505), .C(n_53788), .D(n_39601),
		 .Z(n_252691373));
	notech_reg inst_deco2_reg_112(.CP(n_61902), .D(n_31902), .CD(n_61344), .Q
		(inst_deco2[112]));
	notech_mux2 i_37515(.S(n_54250), .A(inst_deco2[112]), .B(n_42834), .Z(n_31902
		));
	notech_reg inst_deco2_reg_113(.CP(n_61902), .D(n_31908), .CD(n_61344), .Q
		(inst_deco2[113]));
	notech_mux2 i_37523(.S(n_54250), .A(inst_deco2[113]), .B(n_42840), .Z(n_31908
		));
	notech_ao4 i_4727783(.A(n_57502), .B(n_38506), .C(n_53788), .D(n_39595),
		 .Z(n_252491371));
	notech_reg inst_deco2_reg_114(.CP(n_61902), .D(n_31914), .CD(n_61344), .Q
		(inst_deco2[114]));
	notech_mux2 i_37531(.S(n_54250), .A(inst_deco2[114]), .B(n_42846), .Z(n_31914
		));
	notech_reg inst_deco2_reg_115(.CP(n_61902), .D(n_31920), .CD(n_61341), .Q
		(inst_deco2[115]));
	notech_mux2 i_37539(.S(n_54250), .A(inst_deco2[115]), .B(n_42852), .Z(n_31920
		));
	notech_ao4 i_4827784(.A(n_57502), .B(n_38507), .C(n_53788), .D(n_39593),
		 .Z(n_252291369));
	notech_reg inst_deco2_reg_116(.CP(n_61902), .D(n_31926), .CD(n_61341), .Q
		(inst_deco2[116]));
	notech_mux2 i_37547(.S(n_54255), .A(inst_deco2[116]), .B(n_42858), .Z(n_31926
		));
	notech_reg inst_deco2_reg_117(.CP(n_61900), .D(n_31932), .CD(n_61341), .Q
		(inst_deco2[117]));
	notech_mux2 i_37555(.S(n_54255), .A(inst_deco2[117]), .B(n_42864), .Z(n_31932
		));
	notech_nand2 i_123167(.A(n_1980), .B(n_251891365), .Z(n_252091367));
	notech_reg inst_deco2_reg_118(.CP(n_61895), .D(n_31938), .CD(n_61341), .Q
		(inst_deco2[118]));
	notech_mux2 i_37563(.S(n_54255), .A(inst_deco2[118]), .B(n_42870), .Z(n_31938
		));
	notech_ao4 i_321(.A(n_5726), .B(n_251791364), .C(db67), .D(n_39117), .Z(n_251991366
		));
	notech_reg inst_deco2_reg_119(.CP(n_61895), .D(n_31944), .CD(n_61341), .Q
		(inst_deco2[119]));
	notech_mux2 i_37571(.S(n_54250), .A(inst_deco2[119]), .B(n_42876), .Z(n_31944
		));
	notech_nao3 i_1172(.A(n_1987), .B(\to_acu2_0[4] ), .C(n_251991366), .Z(n_251891365
		));
	notech_reg inst_deco2_reg_120(.CP(n_61895), .D(n_31950), .CD(n_61341), .Q
		(inst_deco2[120]));
	notech_mux2 i_37579(.S(n_54250), .A(inst_deco2[120]), .B(n_42882), .Z(n_31950
		));
	notech_and2 i_340(.A(n_2220), .B(n_251591362), .Z(n_251791364));
	notech_reg inst_deco2_reg_121(.CP(n_61895), .D(n_31956), .CD(n_61341), .Q
		(inst_deco2[121]));
	notech_mux2 i_37587(.S(n_54255), .A(inst_deco2[121]), .B(n_42888), .Z(n_31956
		));
	notech_reg inst_deco2_reg_122(.CP(n_61895), .D(n_31962), .CD(n_61341), .Q
		(inst_deco2[122]));
	notech_mux2 i_37595(.S(n_54245), .A(inst_deco2[122]), .B(n_42894), .Z(n_31962
		));
	notech_nao3 i_1169(.A(n_40212), .B(n_40147), .C(n_5717), .Z(n_251591362)
		);
	notech_reg inst_deco2_reg_123(.CP(n_61897), .D(n_31968), .CD(n_61341), .Q
		(inst_deco2[123]));
	notech_mux2 i_37603(.S(n_54245), .A(inst_deco2[123]), .B(n_42900), .Z(n_31968
		));
	notech_mux2 i_70618(.S(adz), .A(n_41571), .B(n_1781), .Z(n_251491361));
	notech_reg inst_deco2_reg_124(.CP(n_61897), .D(n_31974), .CD(n_61341), .Q
		(inst_deco2[124]));
	notech_mux2 i_37611(.S(n_54245), .A(inst_deco2[124]), .B(n_42906), .Z(n_31974
		));
	notech_reg inst_deco2_reg_125(.CP(n_61897), .D(n_31980), .CD(n_61336), .Q
		(inst_deco2[125]));
	notech_mux2 i_37619(.S(n_54245), .A(inst_deco2[125]), .B(n_42912), .Z(n_31980
		));
	notech_reg inst_deco2_reg_126(.CP(n_61897), .D(n_31986), .CD(n_61336), .Q
		(inst_deco2[126]));
	notech_mux2 i_37627(.S(n_54245), .A(inst_deco2[126]), .B(n_42918), .Z(n_31986
		));
	notech_mux2 i_31(.S(twobyte), .A(n_2214), .B(n_2957), .Z(n_251191358));
	notech_reg inst_deco2_reg_127(.CP(n_61897), .D(n_31992), .CD(n_61336), .Q
		(inst_deco2[127]));
	notech_mux2 i_37635(.S(n_54245), .A(inst_deco2[127]), .B(n_42924), .Z(n_31992
		));
	notech_or4 i_1140(.A(n_251191358), .B(n_5674), .C(n_250891355), .D(n_40209
		), .Z(n_251091357));
	notech_reg inst_deco1_reg_0(.CP(n_61895), .D(n_31998), .CD(n_61334), .Q(inst_deco1
		[0]));
	notech_mux2 i_37643(.S(n_57666), .A(inst_deco1[0]), .B(n_38998), .Z(n_31998
		));
	notech_or4 i_1139(.A(n_2958), .B(n_5304), .C(n_2220), .D(\to_acu2_0[4] )
		, .Z(n_250991356));
	notech_reg inst_deco1_reg_1(.CP(n_61895), .D(n_32004), .CD(n_61334), .Q(inst_deco1
		[1]));
	notech_mux2 i_37651(.S(n_57666), .A(inst_deco1[1]), .B(n_39000), .Z(n_32004
		));
	notech_or2 i_144(.A(db67), .B(n_39117), .Z(n_250891355));
	notech_reg inst_deco1_reg_2(.CP(n_61895), .D(n_32010), .CD(n_61336), .Q(inst_deco1
		[2]));
	notech_mux2 i_37659(.S(n_57644), .A(inst_deco1[2]), .B(n_39002), .Z(n_32010
		));
	notech_reg inst_deco1_reg_3(.CP(n_61895), .D(n_32016), .CD(n_61336), .Q(inst_deco1
		[3]));
	notech_mux2 i_37667(.S(n_57644), .A(inst_deco1[3]), .B(n_39004), .Z(n_32016
		));
	notech_nand3 i_210210(.A(\fpu_modrm[0] ), .B(\fpu_indrm[7] ), .C(n_3119)
		, .Z(n_250691353));
	notech_reg inst_deco1_reg_4(.CP(n_61895), .D(n_32022), .CD(n_61336), .Q(inst_deco1
		[4]));
	notech_mux2 i_37675(.S(n_57644), .A(inst_deco1[4]), .B(n_39006), .Z(n_32022
		));
	notech_reg inst_deco1_reg_5(.CP(n_61895), .D(n_32028), .CD(n_61336), .Q(inst_deco1
		[5]));
	notech_mux2 i_37683(.S(n_57644), .A(inst_deco1[5]), .B(n_39008), .Z(n_32028
		));
	notech_reg inst_deco1_reg_6(.CP(n_61895), .D(n_32034), .CD(n_61336), .Q(inst_deco1
		[6]));
	notech_mux2 i_37691(.S(n_57644), .A(inst_deco1[6]), .B(n_39010), .Z(n_32034
		));
	notech_and2 i_268(.A(n_3107), .B(in128[63]), .Z(n_250391350));
	notech_reg inst_deco1_reg_7(.CP(n_61895), .D(n_32040), .CD(n_61334), .Q(inst_deco1
		[7]));
	notech_mux2 i_37699(.S(n_57644), .A(inst_deco1[7]), .B(n_39012), .Z(n_32040
		));
	notech_reg inst_deco1_reg_8(.CP(n_61895), .D(n_32046), .CD(n_61334), .Q(inst_deco1
		[8]));
	notech_mux2 i_37707(.S(n_57644), .A(inst_deco1[8]), .B(n_39014), .Z(n_32046
		));
	notech_reg inst_deco1_reg_9(.CP(n_61895), .D(n_32052), .CD(n_61334), .Q(inst_deco1
		[9]));
	notech_mux2 i_37715(.S(n_57649), .A(inst_deco1[9]), .B(n_39016), .Z(n_32052
		));
	notech_and2 i_267(.A(n_3107), .B(in128[62]), .Z(n_250091347));
	notech_reg inst_deco1_reg_10(.CP(n_61895), .D(n_32058), .CD(n_61334), .Q
		(inst_deco1[10]));
	notech_mux2 i_37723(.S(n_57649), .A(inst_deco1[10]), .B(n_39018), .Z(n_32058
		));
	notech_reg inst_deco1_reg_11(.CP(n_61897), .D(n_32064), .CD(n_61334), .Q
		(inst_deco1[11]));
	notech_mux2 i_37731(.S(n_57649), .A(inst_deco1[11]), .B(n_39020), .Z(n_32064
		));
	notech_reg inst_deco1_reg_12(.CP(n_61900), .D(n_32070), .CD(n_61334), .Q
		(inst_deco1[12]));
	notech_mux2 i_37739(.S(n_57644), .A(inst_deco1[12]), .B(n_39022), .Z(n_32070
		));
	notech_and2 i_266(.A(n_3107), .B(in128[61]), .Z(n_249791344));
	notech_reg inst_deco1_reg_13(.CP(n_61897), .D(n_32076), .CD(n_61334), .Q
		(inst_deco1[13]));
	notech_mux2 i_37747(.S(n_57649), .A(inst_deco1[13]), .B(n_39024), .Z(n_32076
		));
	notech_reg inst_deco1_reg_14(.CP(n_61897), .D(n_32082), .CD(n_61334), .Q
		(inst_deco1[14]));
	notech_mux2 i_37755(.S(n_57649), .A(inst_deco1[14]), .B(n_39026), .Z(n_32082
		));
	notech_reg inst_deco1_reg_15(.CP(n_61897), .D(n_32088), .CD(n_61334), .Q
		(inst_deco1[15]));
	notech_mux2 i_37763(.S(n_57644), .A(inst_deco1[15]), .B(n_39028), .Z(n_32088
		));
	notech_and2 i_265(.A(n_3107), .B(in128[60]), .Z(n_249491341));
	notech_reg inst_deco1_reg_16(.CP(n_61900), .D(n_32094), .CD(n_61334), .Q
		(inst_deco1[16]));
	notech_mux2 i_37771(.S(n_57644), .A(inst_deco1[16]), .B(n_39030), .Z(n_32094
		));
	notech_reg inst_deco1_reg_17(.CP(n_61900), .D(n_32100), .CD(n_61334), .Q
		(inst_deco1[17]));
	notech_mux2 i_37779(.S(n_57644), .A(inst_deco1[17]), .B(n_39031), .Z(n_32100
		));
	notech_reg inst_deco1_reg_18(.CP(n_61900), .D(n_32106), .CD(n_61339), .Q
		(inst_deco1[18]));
	notech_mux2 i_37787(.S(n_57643), .A(inst_deco1[18]), .B(n_39032), .Z(n_32106
		));
	notech_and2 i_264(.A(n_3107), .B(in128[59]), .Z(n_249191338));
	notech_reg inst_deco1_reg_19(.CP(n_61900), .D(n_32112), .CD(n_61339), .Q
		(inst_deco1[19]));
	notech_mux2 i_37795(.S(n_57643), .A(inst_deco1[19]), .B(n_39033), .Z(n_32112
		));
	notech_reg inst_deco1_reg_20(.CP(n_61900), .D(n_32118), .CD(n_61339), .Q
		(inst_deco1[20]));
	notech_mux2 i_37803(.S(n_57643), .A(inst_deco1[20]), .B(n_39034), .Z(n_32118
		));
	notech_reg inst_deco1_reg_21(.CP(n_61897), .D(n_32124), .CD(n_61336), .Q
		(inst_deco1[21]));
	notech_mux2 i_37811(.S(n_57644), .A(inst_deco1[21]), .B(n_39035), .Z(n_32124
		));
	notech_and2 i_263(.A(n_3107), .B(in128[58]), .Z(n_248891335));
	notech_reg inst_deco1_reg_22(.CP(n_61897), .D(n_32130), .CD(n_61339), .Q
		(inst_deco1[22]));
	notech_mux2 i_37819(.S(n_57644), .A(inst_deco1[22]), .B(n_39036), .Z(n_32130
		));
	notech_reg inst_deco1_reg_23(.CP(n_61897), .D(n_32136), .CD(n_61339), .Q
		(inst_deco1[23]));
	notech_mux2 i_37827(.S(n_57644), .A(inst_deco1[23]), .B(n_39037), .Z(n_32136
		));
	notech_reg inst_deco1_reg_24(.CP(n_61897), .D(n_32142), .CD(n_61339), .Q
		(inst_deco1[24]));
	notech_mux2 i_37835(.S(n_57644), .A(inst_deco1[24]), .B(n_39038), .Z(n_32142
		));
	notech_and2 i_262(.A(n_3107), .B(in128[57]), .Z(n_248591332));
	notech_reg inst_deco1_reg_25(.CP(n_61897), .D(n_32148), .CD(n_61339), .Q
		(inst_deco1[25]));
	notech_mux2 i_37843(.S(n_57644), .A(inst_deco1[25]), .B(n_39040), .Z(n_32148
		));
	notech_reg inst_deco1_reg_26(.CP(n_61897), .D(n_32154), .CD(n_61339), .Q
		(inst_deco1[26]));
	notech_mux2 i_37851(.S(n_57644), .A(inst_deco1[26]), .B(n_39042), .Z(n_32154
		));
	notech_reg inst_deco1_reg_27(.CP(n_61897), .D(n_32160), .CD(n_61339), .Q
		(inst_deco1[27]));
	notech_mux2 i_37859(.S(n_57644), .A(inst_deco1[27]), .B(n_39044), .Z(n_32160
		));
	notech_and2 i_261(.A(n_3107), .B(in128[56]), .Z(n_248291329));
	notech_reg inst_deco1_reg_28(.CP(n_61897), .D(n_32166), .CD(n_61336), .Q
		(inst_deco1[28]));
	notech_mux2 i_37867(.S(n_57649), .A(inst_deco1[28]), .B(n_39046), .Z(n_32166
		));
	notech_or2 i_1098(.A(n_3107), .B(n_3095), .Z(n_248191328));
	notech_reg inst_deco1_reg_29(.CP(n_61897), .D(n_32172), .CD(n_61336), .Q
		(inst_deco1[29]));
	notech_mux2 i_37875(.S(n_57654), .A(inst_deco1[29]), .B(n_39048), .Z(n_32172
		));
	notech_reg inst_deco1_reg_30(.CP(n_61897), .D(n_32178), .CD(n_61336), .Q
		(inst_deco1[30]));
	notech_mux2 i_37883(.S(n_57654), .A(inst_deco1[30]), .B(n_39050), .Z(n_32178
		));
	notech_reg inst_deco1_reg_31(.CP(n_61897), .D(n_32184), .CD(n_61336), .Q
		(inst_deco1[31]));
	notech_mux2 i_37891(.S(n_57654), .A(inst_deco1[31]), .B(n_39052), .Z(n_32184
		));
	notech_and2 i_260(.A(n_3095), .B(in128[47]), .Z(n_247891325));
	notech_reg inst_deco1_reg_32(.CP(n_61928), .D(n_32190), .CD(n_61336), .Q
		(inst_deco1[32]));
	notech_mux2 i_37899(.S(n_57654), .A(inst_deco1[32]), .B(n_39054), .Z(n_32190
		));
	notech_and3 i_185(.A(n_2915), .B(n_2914), .C(n_245491301), .Z(n_247791324
		));
	notech_reg inst_deco1_reg_33(.CP(n_61960), .D(n_32196), .CD(n_61336), .Q
		(inst_deco1[33]));
	notech_mux2 i_37907(.S(n_57654), .A(inst_deco1[33]), .B(n_39056), .Z(n_32196
		));
	notech_reg inst_deco1_reg_34(.CP(n_61960), .D(n_32202), .CD(n_61336), .Q
		(inst_deco1[34]));
	notech_mux2 i_37915(.S(n_57654), .A(inst_deco1[34]), .B(n_39058), .Z(n_32202
		));
	notech_reg inst_deco1_reg_35(.CP(n_61960), .D(n_32208), .CD(n_61336), .Q
		(inst_deco1[35]));
	notech_mux2 i_37923(.S(n_57654), .A(inst_deco1[35]), .B(n_39060), .Z(n_32208
		));
	notech_and2 i_259(.A(n_3095), .B(in128[46]), .Z(n_247491321));
	notech_reg inst_deco1_reg_36(.CP(n_61960), .D(n_32214), .CD(n_61336), .Q
		(inst_deco1[36]));
	notech_mux2 i_37931(.S(n_57654), .A(inst_deco1[36]), .B(n_39062), .Z(n_32214
		));
	notech_reg inst_deco1_reg_37(.CP(n_61960), .D(n_32220), .CD(n_61336), .Q
		(inst_deco1[37]));
	notech_mux2 i_37939(.S(n_57655), .A(inst_deco1[37]), .B(n_39064), .Z(n_32220
		));
	notech_reg inst_deco1_reg_38(.CP(n_61960), .D(n_32226), .CD(n_61336), .Q
		(inst_deco1[38]));
	notech_mux2 i_37947(.S(n_57655), .A(inst_deco1[38]), .B(n_39066), .Z(n_32226
		));
	notech_and2 i_258(.A(n_3095), .B(in128[45]), .Z(n_247191318));
	notech_reg inst_deco1_reg_39(.CP(n_61960), .D(n_32232), .CD(n_61399), .Q
		(inst_deco1[39]));
	notech_mux2 i_37955(.S(n_57654), .A(inst_deco1[39]), .B(n_39068), .Z(n_32232
		));
	notech_reg inst_deco1_reg_40(.CP(n_61960), .D(n_32238), .CD(n_61399), .Q
		(inst_deco1[40]));
	notech_mux2 i_37963(.S(n_57654), .A(inst_deco1[40]), .B(n_39071), .Z(n_32238
		));
	notech_reg inst_deco1_reg_41(.CP(n_61960), .D(n_32244), .CD(n_61399), .Q
		(inst_deco1[41]));
	notech_mux2 i_37971(.S(n_57654), .A(inst_deco1[41]), .B(n_39073), .Z(n_32244
		));
	notech_and2 i_257(.A(n_3095), .B(in128[44]), .Z(n_246891315));
	notech_reg inst_deco1_reg_42(.CP(n_61960), .D(n_32250), .CD(n_61399), .Q
		(inst_deco1[42]));
	notech_mux2 i_37979(.S(n_57649), .A(inst_deco1[42]), .B(n_39075), .Z(n_32250
		));
	notech_reg inst_deco1_reg_43(.CP(n_61960), .D(n_32256), .CD(n_61399), .Q
		(inst_deco1[43]));
	notech_mux2 i_37987(.S(n_57649), .A(inst_deco1[43]), .B(n_39076), .Z(n_32256
		));
	notech_reg inst_deco1_reg_44(.CP(n_61956), .D(n_32262), .CD(n_61400), .Q
		(inst_deco1[44]));
	notech_mux2 i_37995(.S(n_57649), .A(inst_deco1[44]), .B(n_39078), .Z(n_32262
		));
	notech_and2 i_256(.A(n_3095), .B(in128[43]), .Z(n_246591312));
	notech_reg inst_deco1_reg_45(.CP(n_61956), .D(n_32268), .CD(n_61400), .Q
		(inst_deco1[45]));
	notech_mux2 i_38003(.S(n_57649), .A(inst_deco1[45]), .B(n_39080), .Z(n_32268
		));
	notech_reg inst_deco1_reg_46(.CP(n_61956), .D(n_32274), .CD(n_61400), .Q
		(inst_deco1[46]));
	notech_mux2 i_38011(.S(n_57649), .A(inst_deco1[46]), .B(n_39082), .Z(n_32274
		));
	notech_reg inst_deco1_reg_47(.CP(n_61956), .D(n_32280), .CD(n_61400), .Q
		(inst_deco1[47]));
	notech_mux2 i_38019(.S(n_57649), .A(inst_deco1[47]), .B(n_39084), .Z(n_32280
		));
	notech_and2 i_255(.A(n_3095), .B(in128[42]), .Z(n_246291309));
	notech_reg inst_deco1_reg_48(.CP(n_61956), .D(n_32286), .CD(n_61400), .Q
		(inst_deco1[48]));
	notech_mux2 i_38027(.S(n_57654), .A(inst_deco1[48]), .B(n_39086), .Z(n_32286
		));
	notech_reg inst_deco1_reg_49(.CP(n_61960), .D(n_32292), .CD(n_61399), .Q
		(inst_deco1[49]));
	notech_mux2 i_38035(.S(n_57654), .A(inst_deco1[49]), .B(n_39088), .Z(n_32292
		));
	notech_reg inst_deco1_reg_50(.CP(n_61960), .D(n_32298), .CD(n_61395), .Q
		(inst_deco1[50]));
	notech_mux2 i_38043(.S(n_57654), .A(inst_deco1[50]), .B(n_39089), .Z(n_32298
		));
	notech_and2 i_254(.A(n_3095), .B(in128[41]), .Z(n_245991306));
	notech_reg inst_deco1_reg_51(.CP(n_61960), .D(n_32304), .CD(n_61395), .Q
		(inst_deco1[51]));
	notech_mux2 i_38051(.S(n_57654), .A(inst_deco1[51]), .B(n_39091), .Z(n_32304
		));
	notech_reg inst_deco1_reg_52(.CP(n_61956), .D(n_32310), .CD(n_61395), .Q
		(inst_deco1[52]));
	notech_mux2 i_38059(.S(n_57654), .A(inst_deco1[52]), .B(n_39093), .Z(n_32310
		));
	notech_reg inst_deco1_reg_53(.CP(n_61956), .D(n_32316), .CD(n_61395), .Q
		(inst_deco1[53]));
	notech_mux2 i_38067(.S(n_57654), .A(inst_deco1[53]), .B(n_39095), .Z(n_32316
		));
	notech_and2 i_253(.A(n_3095), .B(in128[40]), .Z(n_245691303));
	notech_reg inst_deco1_reg_54(.CP(n_61962), .D(n_32322), .CD(n_61395), .Q
		(inst_deco1[54]));
	notech_mux2 i_38075(.S(n_57654), .A(inst_deco1[54]), .B(n_39097), .Z(n_32322
		));
	notech_or2 i_1064(.A(n_247791324), .B(n_3095), .Z(n_245591302));
	notech_reg inst_deco1_reg_55(.CP(n_61962), .D(n_32328), .CD(n_61399), .Q
		(inst_deco1[55]));
	notech_mux2 i_38083(.S(n_57667), .A(inst_deco1[55]), .B(n_39099), .Z(n_32328
		));
	notech_nand2 i_1062(.A(n_245391300), .B(n_39860), .Z(n_245491301));
	notech_reg inst_deco1_reg_56(.CP(n_61962), .D(n_32334), .CD(n_61399), .Q
		(inst_deco1[56]));
	notech_mux2 i_38091(.S(n_57683), .A(inst_deco1[56]), .B(n_39101), .Z(n_32334
		));
	notech_nand2 i_830092(.A(imm_sz[0]), .B(n_39859), .Z(n_245391300));
	notech_reg inst_deco1_reg_57(.CP(n_61962), .D(n_32340), .CD(n_61399), .Q
		(inst_deco1[57]));
	notech_mux2 i_38099(.S(n_57688), .A(inst_deco1[57]), .B(n_39103), .Z(n_32340
		));
	notech_nao3 i_250(.A(n_2175), .B(in128[39]), .C(n_2898), .Z(n_245291299)
		);
	notech_reg inst_deco1_reg_58(.CP(n_61962), .D(n_32346), .CD(n_61395), .Q
		(inst_deco1[58]));
	notech_mux2 i_38107(.S(n_57688), .A(inst_deco1[58]), .B(n_39105), .Z(n_32346
		));
	notech_ao4 i_251(.A(n_2929), .B(n_40046), .C(n_2928), .D(n_40062), .Z(n_245191298
		));
	notech_reg inst_deco1_reg_59(.CP(n_61962), .D(n_32352), .CD(n_61399), .Q
		(inst_deco1[59]));
	notech_mux2 i_38115(.S(n_57683), .A(inst_deco1[59]), .B(n_39107), .Z(n_32352
		));
	notech_and4 i_1059(.A(n_245191298), .B(n_3091), .C(n_3090), .D(n_245291299
		), .Z(n_245091297));
	notech_reg inst_deco1_reg_60(.CP(n_61962), .D(n_32358), .CD(n_61400), .Q
		(inst_deco1[60]));
	notech_mux2 i_38123(.S(n_57683), .A(inst_deco1[60]), .B(n_39109), .Z(n_32358
		));
	notech_reg inst_deco1_reg_61(.CP(n_61962), .D(n_32364), .CD(n_61404), .Q
		(inst_deco1[61]));
	notech_mux2 i_38131(.S(n_57683), .A(inst_deco1[61]), .B(n_39111), .Z(n_32364
		));
	notech_reg inst_deco1_reg_62(.CP(n_61962), .D(n_32370), .CD(n_61400), .Q
		(inst_deco1[62]));
	notech_mux2 i_38139(.S(n_57688), .A(inst_deco1[62]), .B(n_39113), .Z(n_32370
		));
	notech_reg inst_deco1_reg_63(.CP(n_61962), .D(n_32376), .CD(n_61400), .Q
		(inst_deco1[63]));
	notech_mux2 i_38147(.S(n_57688), .A(inst_deco1[63]), .B(n_39115), .Z(n_32376
		));
	notech_reg inst_deco1_reg_64(.CP(n_61962), .D(n_32382), .CD(n_61400), .Q
		(inst_deco1[64]));
	notech_mux2 i_38155(.S(n_57688), .A(inst_deco1[64]), .B(n_39119), .Z(n_32382
		));
	notech_reg inst_deco1_reg_65(.CP(n_61960), .D(n_32388), .CD(n_61404), .Q
		(inst_deco1[65]));
	notech_mux2 i_38163(.S(n_57688), .A(inst_deco1[65]), .B(n_39121), .Z(n_32388
		));
	notech_reg inst_deco1_reg_66(.CP(n_61960), .D(n_32394), .CD(n_61404), .Q
		(inst_deco1[66]));
	notech_mux2 i_38171(.S(n_57688), .A(inst_deco1[66]), .B(n_39123), .Z(n_32394
		));
	notech_reg inst_deco1_reg_67(.CP(n_61960), .D(n_32400), .CD(n_61404), .Q
		(inst_deco1[67]));
	notech_mux2 i_38179(.S(n_57688), .A(inst_deco1[67]), .B(n_39126), .Z(n_32400
		));
	notech_reg inst_deco1_reg_68(.CP(n_61960), .D(n_32406), .CD(n_61404), .Q
		(inst_deco1[68]));
	notech_mux2 i_38187(.S(n_57688), .A(inst_deco1[68]), .B(n_39129), .Z(n_32406
		));
	notech_nao3 i_247(.A(n_2175), .B(in128[38]), .C(n_2898), .Z(n_244191288)
		);
	notech_reg inst_deco1_reg_69(.CP(n_61960), .D(n_32412), .CD(n_61404), .Q
		(inst_deco1[69]));
	notech_mux2 i_38195(.S(n_57678), .A(inst_deco1[69]), .B(n_39132), .Z(n_32412
		));
	notech_ao4 i_248(.A(n_2929), .B(n_40045), .C(n_2928), .D(n_40061), .Z(n_244091287
		));
	notech_reg inst_deco1_reg_70(.CP(n_61962), .D(n_32418), .CD(n_61400), .Q
		(inst_deco1[70]));
	notech_mux2 i_38203(.S(n_57678), .A(inst_deco1[70]), .B(n_39135), .Z(n_32418
		));
	notech_and4 i_1047(.A(n_244091287), .B(n_3086), .C(n_3085), .D(n_244191288
		), .Z(n_243991286));
	notech_reg inst_deco1_reg_71(.CP(n_61962), .D(n_32424), .CD(n_61400), .Q
		(inst_deco1[71]));
	notech_mux2 i_38211(.S(n_57683), .A(inst_deco1[71]), .B(n_39138), .Z(n_32424
		));
	notech_reg inst_deco1_reg_72(.CP(n_61962), .D(n_32430), .CD(n_61400), .Q
		(inst_deco1[72]));
	notech_mux2 i_38219(.S(n_57678), .A(inst_deco1[72]), .B(n_39141), .Z(n_32430
		));
	notech_reg inst_deco1_reg_73(.CP(n_61960), .D(n_32436), .CD(n_61400), .Q
		(inst_deco1[73]));
	notech_mux2 i_38227(.S(n_57678), .A(inst_deco1[73]), .B(n_39144), .Z(n_32436
		));
	notech_reg inst_deco1_reg_74(.CP(n_61962), .D(n_32442), .CD(n_61400), .Q
		(inst_deco1[74]));
	notech_mux2 i_38235(.S(n_57678), .A(inst_deco1[74]), .B(n_39147), .Z(n_32442
		));
	notech_reg inst_deco1_reg_75(.CP(n_61956), .D(n_32448), .CD(n_61400), .Q
		(inst_deco1[75]));
	notech_mux2 i_38243(.S(n_57683), .A(inst_deco1[75]), .B(n_39150), .Z(n_32448
		));
	notech_reg inst_deco1_reg_76(.CP(n_61954), .D(n_32454), .CD(n_61400), .Q
		(inst_deco1[76]));
	notech_mux2 i_38251(.S(n_57683), .A(inst_deco1[76]), .B(n_39153), .Z(n_32454
		));
	notech_reg inst_deco1_reg_77(.CP(n_61954), .D(n_32460), .CD(n_61400), .Q
		(inst_deco1[77]));
	notech_mux2 i_38259(.S(n_57683), .A(inst_deco1[77]), .B(n_39156), .Z(n_32460
		));
	notech_reg inst_deco1_reg_78(.CP(n_61954), .D(n_32466), .CD(n_61400), .Q
		(inst_deco1[78]));
	notech_mux2 i_38267(.S(n_57683), .A(inst_deco1[78]), .B(n_39159), .Z(n_32466
		));
	notech_nao3 i_238(.A(n_2175), .B(in128[36]), .C(n_2898), .Z(n_243191278)
		);
	notech_reg inst_deco1_reg_79(.CP(n_61954), .D(n_32472), .CD(n_61400), .Q
		(inst_deco1[79]));
	notech_mux2 i_38275(.S(n_57683), .A(inst_deco1[79]), .B(n_39162), .Z(n_32472
		));
	notech_ao4 i_239(.A(n_2929), .B(n_40043), .C(n_2928), .D(n_40059), .Z(n_243091277
		));
	notech_reg inst_deco1_reg_80(.CP(n_61954), .D(n_32478), .CD(n_61400), .Q
		(inst_deco1[80]));
	notech_mux2 i_38283(.S(n_57683), .A(inst_deco1[80]), .B(n_39165), .Z(n_32478
		));
	notech_and4 i_1035(.A(n_243091277), .B(n_3081), .C(n_3080), .D(n_243191278
		), .Z(n_242991276));
	notech_reg inst_deco1_reg_81(.CP(n_61954), .D(n_32484), .CD(n_61393), .Q
		(inst_deco1[81]));
	notech_mux2 i_38291(.S(n_57683), .A(inst_deco1[81]), .B(n_39168), .Z(n_32484
		));
	notech_reg inst_deco1_reg_82(.CP(n_61954), .D(n_32490), .CD(n_61393), .Q
		(inst_deco1[82]));
	notech_mux2 i_38299(.S(n_57688), .A(inst_deco1[82]), .B(n_39171), .Z(n_32490
		));
	notech_reg inst_deco1_reg_83(.CP(n_61954), .D(n_32496), .CD(n_61393), .Q
		(inst_deco1[83]));
	notech_mux2 i_38307(.S(n_57689), .A(inst_deco1[83]), .B(n_39174), .Z(n_32496
		));
	notech_reg inst_deco1_reg_84(.CP(n_61954), .D(n_32502), .CD(n_61393), .Q
		(inst_deco1[84]));
	notech_mux2 i_38315(.S(n_57689), .A(inst_deco1[84]), .B(n_39177), .Z(n_32502
		));
	notech_reg inst_deco1_reg_85(.CP(n_61954), .D(n_32508), .CD(n_61393), .Q
		(inst_deco1[85]));
	notech_mux2 i_38323(.S(n_57689), .A(inst_deco1[85]), .B(n_39180), .Z(n_32508
		));
	notech_reg inst_deco1_reg_86(.CP(n_61954), .D(n_32514), .CD(n_61393), .Q
		(inst_deco1[86]));
	notech_mux2 i_38331(.S(n_57689), .A(inst_deco1[86]), .B(n_39182), .Z(n_32514
		));
	notech_reg inst_deco1_reg_87(.CP(n_61951), .D(n_32520), .CD(n_61393), .Q
		(inst_deco1[87]));
	notech_mux2 i_38339(.S(n_57689), .A(inst_deco1[87]), .B(n_39185), .Z(n_32520
		));
	notech_reg inst_deco1_reg_88(.CP(n_61951), .D(n_32526), .CD(n_61393), .Q
		(inst_deco1[88]));
	notech_mux2 i_38347(.S(n_57689), .A(inst_deco1[88]), .B(n_39188), .Z(n_32526
		));
	notech_nao3 i_235(.A(n_2175), .B(in128[35]), .C(n_2898), .Z(n_242191268)
		);
	notech_reg inst_deco1_reg_89(.CP(n_61951), .D(n_32532), .CD(n_61393), .Q
		(inst_deco1[89]));
	notech_mux2 i_38355(.S(n_57689), .A(inst_deco1[89]), .B(n_39191), .Z(n_32532
		));
	notech_ao4 i_236(.A(n_2929), .B(n_40042), .C(n_2928), .D(n_40058), .Z(n_242091267
		));
	notech_reg inst_deco1_reg_90(.CP(n_61951), .D(n_32538), .CD(n_61393), .Q
		(inst_deco1[90]));
	notech_mux2 i_38363(.S(n_57689), .A(inst_deco1[90]), .B(n_39194), .Z(n_32538
		));
	notech_and4 i_1023(.A(n_242091267), .B(n_3076), .C(n_3075), .D(n_242191268
		), .Z(n_241991266));
	notech_reg inst_deco1_reg_91(.CP(n_61951), .D(n_32544), .CD(n_61393), .Q
		(inst_deco1[91]));
	notech_mux2 i_38371(.S(n_57689), .A(inst_deco1[91]), .B(n_39197), .Z(n_32544
		));
	notech_reg inst_deco1_reg_92(.CP(n_61951), .D(n_32550), .CD(n_61390), .Q
		(inst_deco1[92]));
	notech_mux2 i_38379(.S(n_57689), .A(inst_deco1[92]), .B(n_39200), .Z(n_32550
		));
	notech_reg inst_deco1_reg_93(.CP(n_61951), .D(n_32556), .CD(n_61390), .Q
		(inst_deco1[93]));
	notech_mux2 i_38387(.S(n_57689), .A(inst_deco1[93]), .B(n_39203), .Z(n_32556
		));
	notech_reg inst_deco1_reg_94(.CP(n_61951), .D(n_32562), .CD(n_61390), .Q
		(inst_deco1[94]));
	notech_mux2 i_38395(.S(n_57689), .A(inst_deco1[94]), .B(n_39206), .Z(n_32562
		));
	notech_reg inst_deco1_reg_95(.CP(n_61951), .D(n_32568), .CD(n_61390), .Q
		(inst_deco1[95]));
	notech_mux2 i_38403(.S(n_57689), .A(inst_deco1[95]), .B(n_39209), .Z(n_32568
		));
	notech_reg inst_deco1_reg_96(.CP(n_61951), .D(n_32574), .CD(n_61390), .Q
		(inst_deco1[96]));
	notech_mux2 i_38411(.S(n_57688), .A(inst_deco1[96]), .B(n_39212), .Z(n_32574
		));
	notech_reg inst_deco1_reg_97(.CP(n_61956), .D(n_32580), .CD(n_61393), .Q
		(inst_deco1[97]));
	notech_mux2 i_38419(.S(n_57688), .A(inst_deco1[97]), .B(n_39215), .Z(n_32580
		));
	notech_reg inst_deco1_reg_98(.CP(n_61956), .D(n_32586), .CD(n_61393), .Q
		(inst_deco1[98]));
	notech_mux2 i_38427(.S(n_57688), .A(inst_deco1[98]), .B(n_39218), .Z(n_32586
		));
	notech_nao3 i_232(.A(n_2175), .B(in128[34]), .C(n_2898), .Z(n_241191258)
		);
	notech_reg inst_deco1_reg_99(.CP(n_61956), .D(n_32592), .CD(n_61390), .Q
		(inst_deco1[99]));
	notech_mux2 i_38435(.S(n_57688), .A(inst_deco1[99]), .B(n_39221), .Z(n_32592
		));
	notech_ao4 i_233(.A(n_2929), .B(n_40041), .C(n_2928), .D(n_40057), .Z(n_241091257
		));
	notech_reg inst_deco1_reg_100(.CP(n_61956), .D(n_32598), .CD(n_61390), .Q
		(inst_deco1[100]));
	notech_mux2 i_38443(.S(n_57688), .A(inst_deco1[100]), .B(n_39224), .Z(n_32598
		));
	notech_and4 i_1011(.A(n_241091257), .B(n_3071), .C(n_3070), .D(n_241191258
		), .Z(n_240991256));
	notech_reg inst_deco1_reg_101(.CP(n_61956), .D(n_32604), .CD(n_61390), .Q
		(inst_deco1[101]));
	notech_mux2 i_38451(.S(n_57688), .A(inst_deco1[101]), .B(n_39227), .Z(n_32604
		));
	notech_reg inst_deco1_reg_102(.CP(n_61956), .D(n_32610), .CD(n_61395), .Q
		(inst_deco1[102]));
	notech_mux2 i_38459(.S(n_57688), .A(inst_deco1[102]), .B(n_39230), .Z(n_32610
		));
	notech_reg inst_deco1_reg_103(.CP(n_61956), .D(n_32616), .CD(n_61395), .Q
		(inst_deco1[103]));
	notech_mux2 i_38467(.S(n_57689), .A(inst_deco1[103]), .B(n_39069), .Z(n_32616
		));
	notech_reg inst_deco1_reg_104(.CP(n_61956), .D(n_32622), .CD(n_61395), .Q
		(inst_deco1[104]));
	notech_mux2 i_38475(.S(n_57689), .A(inst_deco1[104]), .B(n_39233), .Z(n_32622
		));
	notech_reg inst_deco1_reg_105(.CP(n_61956), .D(n_32628), .CD(n_61395), .Q
		(inst_deco1[105]));
	notech_mux2 i_38483(.S(n_57689), .A(inst_deco1[105]), .B(n_39236), .Z(n_32628
		));
	notech_reg inst_deco1_reg_106(.CP(n_61956), .D(n_32634), .CD(n_61395), .Q
		(inst_deco1[106]));
	notech_mux2 i_38491(.S(n_57688), .A(inst_deco1[106]), .B(n_39239), .Z(n_32634
		));
	notech_reg inst_deco1_reg_107(.CP(n_61956), .D(n_32640), .CD(n_61395), .Q
		(inst_deco1[107]));
	notech_mux2 i_38499(.S(n_57689), .A(inst_deco1[107]), .B(n_39242), .Z(n_32640
		));
	notech_reg inst_deco1_reg_108(.CP(n_61954), .D(n_32646), .CD(n_61395), .Q
		(inst_deco1[108]));
	notech_mux2 i_38507(.S(n_57689), .A(inst_deco1[108]), .B(n_39245), .Z(n_32646
		));
	notech_nao3 i_229(.A(n_2175), .B(in128[33]), .C(n_2898), .Z(n_240191248)
		);
	notech_reg inst_deco1_reg_109(.CP(n_61954), .D(n_32652), .CD(n_61395), .Q
		(inst_deco1[109]));
	notech_mux2 i_38515(.S(n_57672), .A(inst_deco1[109]), .B(n_39248), .Z(n_32652
		));
	notech_ao4 i_230(.A(n_2929), .B(n_40040), .C(n_2928), .D(n_40056), .Z(n_240091247
		));
	notech_reg inst_deco1_reg_110(.CP(n_61954), .D(n_32658), .CD(n_61395), .Q
		(inst_deco1[110]));
	notech_mux2 i_38523(.S(n_57672), .A(inst_deco1[110]), .B(n_39252), .Z(n_32658
		));
	notech_and4 i_999(.A(n_240091247), .B(n_3066), .C(n_3065), .D(n_240191248
		), .Z(n_239991246));
	notech_reg inst_deco1_reg_111(.CP(n_61954), .D(n_32664), .CD(n_61395), .Q
		(inst_deco1[111]));
	notech_mux2 i_38531(.S(n_57672), .A(inst_deco1[111]), .B(n_39255), .Z(n_32664
		));
	notech_reg inst_deco1_reg_112(.CP(n_61954), .D(n_32670), .CD(n_61395), .Q
		(inst_deco1[112]));
	notech_mux2 i_38539(.S(n_57672), .A(inst_deco1[112]), .B(n_39258), .Z(n_32670
		));
	notech_reg inst_deco1_reg_113(.CP(n_61954), .D(n_32676), .CD(n_61393), .Q
		(inst_deco1[113]));
	notech_mux2 i_38547(.S(n_57672), .A(inst_deco1[113]), .B(n_39261), .Z(n_32676
		));
	notech_reg inst_deco1_reg_114(.CP(n_61956), .D(n_32682), .CD(n_61393), .Q
		(inst_deco1[114]));
	notech_mux2 i_38555(.S(n_57672), .A(inst_deco1[114]), .B(n_39264), .Z(n_32682
		));
	notech_reg inst_deco1_reg_115(.CP(n_61954), .D(n_32688), .CD(n_61393), .Q
		(inst_deco1[115]));
	notech_mux2 i_38563(.S(n_57672), .A(inst_deco1[115]), .B(n_39267), .Z(n_32688
		));
	notech_reg inst_deco1_reg_116(.CP(n_61954), .D(n_32694), .CD(n_61393), .Q
		(inst_deco1[116]));
	notech_mux2 i_38571(.S(n_57677), .A(inst_deco1[116]), .B(n_39270), .Z(n_32694
		));
	notech_reg inst_deco1_reg_117(.CP(n_61954), .D(n_32700), .CD(n_61393), .Q
		(inst_deco1[117]));
	notech_mux2 i_38579(.S(n_57677), .A(inst_deco1[117]), .B(n_39273), .Z(n_32700
		));
	notech_reg inst_deco1_reg_118(.CP(n_61970), .D(n_32706), .CD(n_61395), .Q
		(inst_deco1[118]));
	notech_mux2 i_38587(.S(n_57677), .A(inst_deco1[118]), .B(n_39276), .Z(n_32706
		));
	notech_nao3 i_225(.A(n_2175), .B(in128[32]), .C(n_2898), .Z(n_239191238)
		);
	notech_reg inst_deco1_reg_119(.CP(n_61970), .D(n_32712), .CD(n_61395), .Q
		(inst_deco1[119]));
	notech_mux2 i_38595(.S(n_57672), .A(inst_deco1[119]), .B(n_39279), .Z(n_32712
		));
	notech_ao4 i_227(.A(n_2929), .B(n_40039), .C(n_2928), .D(n_40055), .Z(n_239091237
		));
	notech_reg inst_deco1_reg_120(.CP(n_61970), .D(n_32718), .CD(n_61395), .Q
		(inst_deco1[120]));
	notech_mux2 i_38603(.S(n_57672), .A(inst_deco1[120]), .B(n_39282), .Z(n_32718
		));
	notech_and4 i_987(.A(n_239091237), .B(n_3061), .C(n_3057), .D(n_239191238
		), .Z(n_238991236));
	notech_reg inst_deco1_reg_121(.CP(n_61970), .D(n_32724), .CD(n_61393), .Q
		(inst_deco1[121]));
	notech_mux2 i_38611(.S(n_57677), .A(inst_deco1[121]), .B(n_39285), .Z(n_32724
		));
	notech_reg inst_deco1_reg_122(.CP(n_61970), .D(n_32730), .CD(n_61393), .Q
		(inst_deco1[122]));
	notech_mux2 i_38619(.S(n_57667), .A(inst_deco1[122]), .B(n_39288), .Z(n_32730
		));
	notech_reg inst_deco1_reg_123(.CP(n_61970), .D(n_32736), .CD(n_61404), .Q
		(inst_deco1[123]));
	notech_mux2 i_38627(.S(n_57667), .A(inst_deco1[123]), .B(n_39291), .Z(n_32736
		));
	notech_reg inst_deco1_reg_124(.CP(n_61970), .D(n_32742), .CD(n_61410), .Q
		(inst_deco1[124]));
	notech_mux2 i_38635(.S(n_57667), .A(inst_deco1[124]), .B(n_39294), .Z(n_32742
		));
	notech_reg inst_deco1_reg_125(.CP(n_61970), .D(n_32748), .CD(n_61410), .Q
		(inst_deco1[125]));
	notech_mux2 i_38643(.S(n_57667), .A(inst_deco1[125]), .B(n_39297), .Z(n_32748
		));
	notech_reg inst_deco1_reg_126(.CP(n_61970), .D(n_32754), .CD(n_61410), .Q
		(inst_deco1[126]));
	notech_mux2 i_38651(.S(n_57667), .A(inst_deco1[126]), .B(n_39300), .Z(n_32754
		));
	notech_reg inst_deco1_reg_127(.CP(n_61970), .D(n_32760), .CD(n_61410), .Q
		(inst_deco1[127]));
	notech_mux2 i_38659(.S(n_57667), .A(inst_deco1[127]), .B(n_38400), .Z(n_32760
		));
	notech_reg overgs_reg(.CP(n_61970), .D(n_32766), .CD(n_61410), .Q(overgs
		));
	notech_mux2 i_38667(.S(n_3144), .A(n_41571), .B(overgs), .Z(n_32766));
	notech_ao3 i_976(.A(n_245391300), .B(n_39860), .C(n_2884), .Z(n_238191228
		));
	notech_reg over_seg2_reg_5(.CP(n_61970), .D(n_32772), .CD(n_61410), .Q(\over_seg2[5] 
		));
	notech_mux2 i_38675(.S(n_54245), .A(\over_seg2[5] ), .B(n_46109), .Z(n_32772
		));
	notech_nao3 i_221(.A(n_2175), .B(in128[31]), .C(n_2898), .Z(n_238091227)
		);
	notech_reg over_seg1_reg_5(.CP(n_61970), .D(n_32778), .CD(n_61410), .Q(\over_seg1[5] 
		));
	notech_mux2 i_38683(.S(n_57667), .A(\over_seg1[5] ), .B(n_38399), .Z(n_32778
		));
	notech_ao4 i_222(.A(n_2928), .B(n_40054), .C(n_2929), .D(n_40038), .Z(n_237991226
		));
	notech_reg to_acu2_reg_0(.CP(n_61970), .D(n_32784), .CD(n_61410), .Q(to_acu2
		[0]));
	notech_mux2 i_38691(.S(n_54250), .A(to_acu2[0]), .B(n_3547), .Z(n_32784)
		);
	notech_and4 i_973(.A(n_237991226), .B(n_237191218), .C(n_238091227), .D(n_3053
		), .Z(n_237891225));
	notech_reg to_acu2_reg_1(.CP(n_61967), .D(n_32790), .CD(n_61410), .Q(to_acu2
		[1]));
	notech_mux2 i_38699(.S(n_54250), .A(to_acu2[1]), .B(n_3810), .Z(n_32790)
		);
	notech_reg to_acu2_reg_2(.CP(n_61967), .D(n_32796), .CD(n_61410), .Q(to_acu2
		[2]));
	notech_mux2 i_38707(.S(n_54250), .A(to_acu2[2]), .B(n_3545), .Z(n_32796)
		);
	notech_reg to_acu2_reg_3(.CP(n_61970), .D(n_32802), .CD(n_61409), .Q(to_acu2
		[3]));
	notech_mux2 i_38715(.S(n_54245), .A(to_acu2[3]), .B(n_3807), .Z(n_32802)
		);
	notech_reg to_acu2_reg_4(.CP(n_61970), .D(n_32808), .CD(n_61409), .Q(to_acu2
		[4]));
	notech_mux2 i_38723(.S(n_54245), .A(to_acu2[4]), .B(n_3543), .Z(n_32808)
		);
	notech_or2 i_964(.A(n_2922), .B(n_40030), .Z(n_237491221));
	notech_reg to_acu2_reg_5(.CP(n_61970), .D(n_32814), .CD(n_61409), .Q(to_acu2
		[5]));
	notech_mux2 i_38731(.S(n_54245), .A(to_acu2[5]), .B(n_3804), .Z(n_32814)
		);
	notech_reg to_acu2_reg_6(.CP(n_61970), .D(n_32820), .CD(n_61409), .Q(to_acu2
		[6]));
	notech_mux2 i_38739(.S(n_54255), .A(to_acu2[6]), .B(n_3802), .Z(n_32820)
		);
	notech_reg to_acu2_reg_7(.CP(n_61970), .D(n_32826), .CD(n_61409), .Q(to_acu2
		[7]));
	notech_mux2 i_38747(.S(n_54256), .A(to_acu2[7]), .B(n_3800), .Z(n_32826)
		);
	notech_or2 i_966(.A(n_2921), .B(n_40022), .Z(n_237191218));
	notech_reg to_acu2_reg_8(.CP(n_61972), .D(n_32832), .CD(n_61409), .Q(to_acu2
		[8]));
	notech_mux2 i_38755(.S(n_54256), .A(to_acu2[8]), .B(n_3541), .Z(n_32832)
		);
	notech_nao3 i_216(.A(n_2175), .B(in128[30]), .C(n_53815), .Z(n_237091217
		));
	notech_reg to_acu2_reg_9(.CP(n_61972), .D(n_32838), .CD(n_61409), .Q(to_acu2
		[9]));
	notech_mux2 i_38763(.S(n_54256), .A(to_acu2[9]), .B(n_3797), .Z(n_32838)
		);
	notech_ao4 i_218(.A(n_2928), .B(n_40053), .C(n_2929), .D(n_40037), .Z(n_236991216
		));
	notech_reg to_acu2_reg_10(.CP(n_61972), .D(n_32844), .CD(n_61409), .Q(to_acu2
		[10]));
	notech_mux2 i_38771(.S(n_54256), .A(to_acu2[10]), .B(n_3795), .Z(n_32844
		));
	notech_and4 i_955(.A(n_236991216), .B(n_236191208), .C(n_237091217), .D(n_3048
		), .Z(n_236891215));
	notech_reg to_acu2_reg_11(.CP(n_61972), .D(n_32850), .CD(n_61409), .Q(to_acu2
		[11]));
	notech_mux2 i_38779(.S(n_54256), .A(to_acu2[11]), .B(n_3793), .Z(n_32850
		));
	notech_reg to_acu2_reg_12(.CP(n_61972), .D(n_32856), .CD(n_61409), .Q(to_acu2
		[12]));
	notech_mux2 i_38787(.S(n_54256), .A(to_acu2[12]), .B(n_3539), .Z(n_32856
		));
	notech_reg to_acu2_reg_13(.CP(n_61972), .D(n_32862), .CD(n_61409), .Q(to_acu2
		[13]));
	notech_mux2 i_38795(.S(n_54256), .A(to_acu2[13]), .B(n_3537), .Z(n_32862
		));
	notech_reg to_acu2_reg_14(.CP(n_61972), .D(n_32868), .CD(n_61412), .Q(to_acu2
		[14]));
	notech_mux2 i_38803(.S(n_54256), .A(to_acu2[14]), .B(n_3535), .Z(n_32868
		));
	notech_or2 i_946(.A(n_2922), .B(n_40029), .Z(n_236491211));
	notech_reg to_acu2_reg_15(.CP(n_61972), .D(n_32874), .CD(n_61412), .Q(to_acu2
		[15]));
	notech_mux2 i_38811(.S(n_54256), .A(to_acu2[15]), .B(n_3788), .Z(n_32874
		));
	notech_reg to_acu2_reg_16(.CP(n_61972), .D(n_32880), .CD(n_61412), .Q(to_acu2
		[16]));
	notech_mux2 i_38819(.S(n_54256), .A(to_acu2[16]), .B(n_3786), .Z(n_32880
		));
	notech_reg to_acu2_reg_17(.CP(n_61972), .D(n_32886), .CD(n_61412), .Q(to_acu2
		[17]));
	notech_mux2 i_38827(.S(n_54256), .A(to_acu2[17]), .B(n_3784), .Z(n_32886
		));
	notech_or2 i_948(.A(n_2921), .B(n_40021), .Z(n_236191208));
	notech_reg to_acu2_reg_18(.CP(n_61972), .D(n_32892), .CD(n_61412), .Q(to_acu2
		[18]));
	notech_mux2 i_38835(.S(n_54256), .A(to_acu2[18]), .B(n_3782), .Z(n_32892
		));
	notech_nao3 i_211(.A(n_2175), .B(in128[29]), .C(n_53815), .Z(n_236091207
		));
	notech_reg to_acu2_reg_19(.CP(n_61972), .D(n_32898), .CD(n_61412), .Q(to_acu2
		[19]));
	notech_mux2 i_38843(.S(n_54256), .A(to_acu2[19]), .B(n_2033), .Z(n_32898
		));
	notech_ao4 i_212(.A(n_2928), .B(n_40052), .C(n_2929), .D(n_40036), .Z(n_235991206
		));
	notech_reg to_acu2_reg_20(.CP(n_61972), .D(n_32904), .CD(n_61412), .Q(to_acu2
		[20]));
	notech_mux2 i_38851(.S(n_54255), .A(to_acu2[20]), .B(n_3780), .Z(n_32904
		));
	notech_and4 i_943(.A(n_235991206), .B(n_235191198), .C(n_236091207), .D(n_3043
		), .Z(n_235891205));
	notech_reg to_acu2_reg_21(.CP(n_61972), .D(n_32910), .CD(n_61412), .Q(to_acu2
		[21]));
	notech_mux2 i_38859(.S(n_54255), .A(to_acu2[21]), .B(n_3778), .Z(n_32910
		));
	notech_reg to_acu2_reg_22(.CP(n_61970), .D(n_32916), .CD(n_61412), .Q(to_acu2
		[22]));
	notech_mux2 i_38867(.S(n_54255), .A(to_acu2[22]), .B(n_3533), .Z(n_32916
		));
	notech_reg to_acu2_reg_23(.CP(n_61972), .D(n_32922), .CD(n_61412), .Q(to_acu2
		[23]));
	notech_mux2 i_38875(.S(n_54255), .A(to_acu2[23]), .B(n_3531), .Z(n_32922
		));
	notech_reg to_acu2_reg_24(.CP(n_61972), .D(n_32928), .CD(n_61412), .Q(to_acu2
		[24]));
	notech_mux2 i_38883(.S(n_54255), .A(to_acu2[24]), .B(n_3529), .Z(n_32928
		));
	notech_or2 i_934(.A(n_2922), .B(n_40028), .Z(n_235491201));
	notech_reg to_acu2_reg_25(.CP(n_61972), .D(n_32934), .CD(n_61410), .Q(to_acu2
		[25]));
	notech_mux2 i_38891(.S(n_54255), .A(to_acu2[25]), .B(n_3527), .Z(n_32934
		));
	notech_reg to_acu2_reg_26(.CP(n_61972), .D(n_32940), .CD(n_61410), .Q(to_acu2
		[26]));
	notech_mux2 i_38899(.S(n_54255), .A(to_acu2[26]), .B(n_3525), .Z(n_32940
		));
	notech_reg to_acu2_reg_27(.CP(n_61972), .D(n_32946), .CD(n_61410), .Q(to_acu2
		[27]));
	notech_mux2 i_38907(.S(n_54255), .A(to_acu2[27]), .B(n_3523), .Z(n_32946
		));
	notech_or2 i_936(.A(n_2921), .B(n_40020), .Z(n_235191198));
	notech_reg to_acu2_reg_28(.CP(n_61972), .D(n_32952), .CD(n_61410), .Q(to_acu2
		[28]));
	notech_mux2 i_38915(.S(n_54255), .A(to_acu2[28]), .B(n_3521), .Z(n_32952
		));
	notech_nao3 i_205(.A(n_2175), .B(in128[28]), .C(n_53815), .Z(n_235091197
		));
	notech_reg to_acu2_reg_29(.CP(n_61967), .D(n_32958), .CD(n_61410), .Q(to_acu2
		[29]));
	notech_mux2 i_38923(.S(n_54255), .A(to_acu2[29]), .B(n_3769), .Z(n_32958
		));
	notech_ao4 i_206(.A(n_2928), .B(n_40051), .C(n_2929), .D(n_40035), .Z(n_234991196
		));
	notech_reg to_acu2_reg_30(.CP(n_61965), .D(n_32964), .CD(n_61410), .Q(to_acu2
		[30]));
	notech_mux2 i_38931(.S(n_54255), .A(to_acu2[30]), .B(n_3767), .Z(n_32964
		));
	notech_and4 i_931(.A(n_234991196), .B(n_234191188), .C(n_235091197), .D(n_3038
		), .Z(n_234891195));
	notech_reg to_acu2_reg_31(.CP(n_61965), .D(n_32970), .CD(n_61410), .Q(to_acu2
		[31]));
	notech_mux2 i_38939(.S(n_54255), .A(to_acu2[31]), .B(n_3765), .Z(n_32970
		));
	notech_reg to_acu2_reg_32(.CP(n_61965), .D(n_32976), .CD(n_61410), .Q(to_acu2
		[32]));
	notech_mux2 i_38947(.S(n_54255), .A(to_acu2[32]), .B(n_3763), .Z(n_32976
		));
	notech_reg to_acu2_reg_33(.CP(n_61965), .D(n_32982), .CD(n_61410), .Q(to_acu2
		[33]));
	notech_mux2 i_38955(.S(n_54187), .A(to_acu2[33]), .B(n_3761), .Z(n_32982
		));
	notech_reg to_acu2_reg_34(.CP(n_61965), .D(n_32988), .CD(n_61410), .Q(to_acu2
		[34]));
	notech_mux2 i_38963(.S(n_54187), .A(to_acu2[34]), .B(n_3759), .Z(n_32988
		));
	notech_or2 i_922(.A(n_2922), .B(n_40027), .Z(n_234491191));
	notech_reg to_acu2_reg_35(.CP(n_61965), .D(n_32994), .CD(n_61405), .Q(to_acu2
		[35]));
	notech_mux2 i_38971(.S(n_54187), .A(to_acu2[35]), .B(n_3757), .Z(n_32994
		));
	notech_reg to_acu2_reg_36(.CP(n_61965), .D(n_33000), .CD(n_61405), .Q(to_acu2
		[36]));
	notech_mux2 i_38979(.S(n_54187), .A(to_acu2[36]), .B(n_3755), .Z(n_33000
		));
	notech_reg to_acu2_reg_37(.CP(n_61965), .D(n_33006), .CD(n_61405), .Q(to_acu2
		[37]));
	notech_mux2 i_38987(.S(n_54187), .A(to_acu2[37]), .B(n_3753), .Z(n_33006
		));
	notech_or2 i_924(.A(n_2921), .B(n_40019), .Z(n_234191188));
	notech_reg to_acu2_reg_38(.CP(n_61965), .D(n_33012), .CD(n_61404), .Q(to_acu2
		[38]));
	notech_mux2 i_38995(.S(n_54187), .A(to_acu2[38]), .B(n_3751), .Z(n_33012
		));
	notech_or4 i_201(.A(n_2887), .B(n_39845), .C(n_2885), .D(n_40013), .Z(n_234091187
		));
	notech_reg to_acu2_reg_39(.CP(n_61965), .D(n_33022), .CD(n_61404), .Q(to_acu2
		[39]));
	notech_ao3 i_39007(.A(to_acu2[39]), .B(1'b1), .C(n_54188), .Z(n_33022)
		);
	notech_reg to_acu2_reg_40(.CP(n_61965), .D(n_33024), .CD(n_61405), .Q(to_acu2
		[40]));
	notech_mux2 i_39011(.S(n_54188), .A(to_acu2[40]), .B(n_3749), .Z(n_33024
		));
	notech_reg to_acu2_reg_41(.CP(n_61962), .D(n_33030), .CD(n_61405), .Q(to_acu2
		[41]));
	notech_mux2 i_39019(.S(n_54188), .A(to_acu2[41]), .B(n_3747), .Z(n_33030
		));
	notech_and4 i_918(.A(n_3035), .B(n_234091187), .C(n_233391180), .D(n_3033
		), .Z(n_233791184));
	notech_reg to_acu2_reg_42(.CP(n_61962), .D(n_33036), .CD(n_61405), .Q(to_acu2
		[42]));
	notech_mux2 i_39027(.S(n_54188), .A(to_acu2[42]), .B(n_3745), .Z(n_33036
		));
	notech_nao3 i_915(.A(n_2156), .B(in128[22]), .C(n_53815), .Z(n_233691183
		));
	notech_reg to_acu2_reg_43(.CP(n_61962), .D(n_33042), .CD(n_61405), .Q(to_acu2
		[43]));
	notech_mux2 i_39035(.S(n_54188), .A(to_acu2[43]), .B(n_3743), .Z(n_33042
		));
	notech_reg to_acu2_reg_44(.CP(n_61962), .D(n_33048), .CD(n_61405), .Q(to_acu2
		[44]));
	notech_mux2 i_39043(.S(n_54188), .A(to_acu2[44]), .B(n_3741), .Z(n_33048
		));
	notech_reg to_acu2_reg_45(.CP(n_61962), .D(n_33054), .CD(n_61404), .Q(to_acu2
		[45]));
	notech_mux2 i_39051(.S(n_54188), .A(to_acu2[45]), .B(n_3739), .Z(n_33054
		));
	notech_nao3 i_913(.A(n_2894), .B(in128[46]), .C(n_2885), .Z(n_233391180)
		);
	notech_reg to_acu2_reg_46(.CP(n_61965), .D(n_33060), .CD(n_61404), .Q(to_acu2
		[46]));
	notech_mux2 i_39059(.S(n_54187), .A(to_acu2[46]), .B(n_3737), .Z(n_33060
		));
	notech_or4 i_196(.A(n_2887), .B(n_39845), .C(n_2885), .D(n_40012), .Z(n_233291179
		));
	notech_reg to_acu2_reg_47(.CP(n_61965), .D(n_33066), .CD(n_61404), .Q(to_acu2
		[47]));
	notech_mux2 i_39067(.S(n_54187), .A(to_acu2[47]), .B(n_3735), .Z(n_33066
		));
	notech_reg to_acu2_reg_48(.CP(n_61965), .D(n_33072), .CD(n_61404), .Q(to_acu2
		[48]));
	notech_mux2 i_39075(.S(n_54187), .A(to_acu2[48]), .B(n_3733), .Z(n_33072
		));
	notech_reg to_acu2_reg_49(.CP(n_61965), .D(n_33078), .CD(n_61404), .Q(to_acu2
		[49]));
	notech_mux2 i_39083(.S(n_54182), .A(to_acu2[49]), .B(n_3731), .Z(n_33078
		));
	notech_and4 i_908(.A(n_3030), .B(n_233291179), .C(n_232591172), .D(n_3028
		), .Z(n_232991176));
	notech_reg to_acu2_reg_50(.CP(n_61965), .D(n_33084), .CD(n_61404), .Q(to_acu2
		[50]));
	notech_mux2 i_39091(.S(n_54187), .A(to_acu2[50]), .B(n_3729), .Z(n_33084
		));
	notech_nao3 i_905(.A(n_2156), .B(in128[21]), .C(n_53815), .Z(n_232891175
		));
	notech_reg to_acu2_reg_51(.CP(n_61967), .D(n_33090), .CD(n_61404), .Q(to_acu2
		[51]));
	notech_mux2 i_39099(.S(n_54187), .A(to_acu2[51]), .B(n_3727), .Z(n_33090
		));
	notech_reg to_acu2_reg_52(.CP(n_61967), .D(n_33096), .CD(n_61404), .Q(to_acu2
		[52]));
	notech_mux2 i_39107(.S(n_54187), .A(to_acu2[52]), .B(n_3725), .Z(n_33096
		));
	notech_reg to_acu2_reg_53(.CP(n_61967), .D(n_33102), .CD(n_61404), .Q(to_acu2
		[53]));
	notech_mux2 i_39115(.S(n_54187), .A(to_acu2[53]), .B(n_3723), .Z(n_33102
		));
	notech_nao3 i_903(.A(n_2894), .B(in128[45]), .C(n_2885), .Z(n_232591172)
		);
	notech_reg to_acu2_reg_54(.CP(n_61967), .D(n_33108), .CD(n_61404), .Q(to_acu2
		[54]));
	notech_mux2 i_39123(.S(n_54187), .A(to_acu2[54]), .B(n_3721), .Z(n_33108
		));
	notech_or4 i_192(.A(n_2887), .B(n_39845), .C(n_2885), .D(n_40011), .Z(n_232491171
		));
	notech_reg to_acu2_reg_55(.CP(n_61967), .D(n_33114), .CD(n_61404), .Q(to_acu2
		[55]));
	notech_mux2 i_39131(.S(n_54187), .A(to_acu2[55]), .B(n_3719), .Z(n_33114
		));
	notech_reg to_acu2_reg_56(.CP(n_61967), .D(n_33120), .CD(n_61409), .Q(to_acu2
		[56]));
	notech_mux2 i_39139(.S(n_54187), .A(to_acu2[56]), .B(n_3717), .Z(n_33120
		));
	notech_reg to_acu2_reg_57(.CP(n_61967), .D(n_33126), .CD(n_61409), .Q(to_acu2
		[57]));
	notech_mux2 i_39147(.S(n_54187), .A(to_acu2[57]), .B(n_3715), .Z(n_33126
		));
	notech_and4 i_898(.A(n_3025), .B(n_232491171), .C(n_231791164), .D(n_3023
		), .Z(n_232191168));
	notech_reg to_acu2_reg_58(.CP(n_61967), .D(n_33132), .CD(n_61409), .Q(to_acu2
		[58]));
	notech_mux2 i_39155(.S(n_54187), .A(to_acu2[58]), .B(n_3713), .Z(n_33132
		));
	notech_nao3 i_895(.A(n_2156), .B(in128[20]), .C(n_53815), .Z(n_232091167
		));
	notech_reg to_acu2_reg_59(.CP(n_61967), .D(n_33138), .CD(n_61405), .Q(to_acu2
		[59]));
	notech_mux2 i_39163(.S(n_54188), .A(to_acu2[59]), .B(n_3711), .Z(n_33138
		));
	notech_reg to_acu2_reg_60(.CP(n_61967), .D(n_33144), .CD(n_61409), .Q(to_acu2
		[60]));
	notech_mux2 i_39171(.S(n_54171), .A(to_acu2[60]), .B(n_3709), .Z(n_33144
		));
	notech_reg to_acu2_reg_61(.CP(n_61967), .D(n_33150), .CD(n_61409), .Q(to_acu2
		[61]));
	notech_mux2 i_39179(.S(n_54171), .A(to_acu2[61]), .B(n_3707), .Z(n_33150
		));
	notech_nao3 i_893(.A(n_2894), .B(in128[44]), .C(n_2885), .Z(n_231791164)
		);
	notech_reg to_acu2_reg_62(.CP(n_61965), .D(n_33156), .CD(n_61409), .Q(to_acu2
		[62]));
	notech_mux2 i_39187(.S(n_54171), .A(to_acu2[62]), .B(n_3705), .Z(n_33156
		));
	notech_or4 i_176(.A(n_2887), .B(n_39845), .C(n_2885), .D(n_40010), .Z(n_231691163
		));
	notech_reg to_acu2_reg_63(.CP(n_61967), .D(n_33162), .CD(n_61409), .Q(to_acu2
		[63]));
	notech_mux2 i_39195(.S(n_54171), .A(to_acu2[63]), .B(n_3703), .Z(n_33162
		));
	notech_reg to_acu2_reg_64(.CP(n_61965), .D(n_33168), .CD(n_61409), .Q(to_acu2
		[64]));
	notech_mux2 i_39203(.S(n_54171), .A(to_acu2[64]), .B(n_3519), .Z(n_33168
		));
	notech_reg to_acu2_reg_65(.CP(n_61965), .D(n_33174), .CD(n_61409), .Q(to_acu2
		[65]));
	notech_mux2 i_39211(.S(n_54171), .A(to_acu2[65]), .B(n_3517), .Z(n_33174
		));
	notech_and4 i_888(.A(n_3020), .B(n_231691163), .C(n_230991156), .D(n_3018
		), .Z(n_231391160));
	notech_reg to_acu2_reg_66(.CP(n_61965), .D(n_33180), .CD(n_61405), .Q(to_acu2
		[66]));
	notech_mux2 i_39219(.S(n_54171), .A(to_acu2[66]), .B(n_3515), .Z(n_33180
		));
	notech_nao3 i_885(.A(n_2156), .B(in128[19]), .C(n_53815), .Z(n_231291159
		));
	notech_reg to_acu2_reg_67(.CP(n_61967), .D(n_33186), .CD(n_61405), .Q(to_acu2
		[67]));
	notech_mux2 i_39227(.S(n_54198), .A(to_acu2[67]), .B(n_3513), .Z(n_33186
		));
	notech_reg to_acu2_reg_68(.CP(n_61967), .D(n_33192), .CD(n_61405), .Q(to_acu2
		[68]));
	notech_mux2 i_39235(.S(n_54198), .A(to_acu2[68]), .B(n_2034), .Z(n_33192
		));
	notech_reg to_acu2_reg_69(.CP(n_61967), .D(n_33198), .CD(n_61405), .Q(to_acu2
		[69]));
	notech_mux2 i_39243(.S(n_54198), .A(to_acu2[69]), .B(n_3511), .Z(n_33198
		));
	notech_nao3 i_883(.A(n_2894), .B(in128[43]), .C(n_53797), .Z(n_230991156
		));
	notech_reg to_acu2_reg_70(.CP(n_61967), .D(n_33204), .CD(n_61405), .Q(to_acu2
		[70]));
	notech_mux2 i_39251(.S(n_54171), .A(to_acu2[70]), .B(n_2039), .Z(n_33204
		));
	notech_or4 i_173(.A(n_2887), .B(n_39845), .C(n_53797), .D(n_40009), .Z(n_230891155
		));
	notech_reg to_acu2_reg_71(.CP(n_61967), .D(n_33210), .CD(n_61405), .Q(to_acu2
		[71]));
	notech_mux2 i_39259(.S(n_54171), .A(to_acu2[71]), .B(n_2010), .Z(n_33210
		));
	notech_reg to_acu2_reg_72(.CP(n_61935), .D(n_33216), .CD(n_61405), .Q(to_acu2
		[72]));
	notech_mux2 i_39267(.S(n_54198), .A(to_acu2[72]), .B(n_2035), .Z(n_33216
		));
	notech_reg to_acu2_reg_73(.CP(n_61935), .D(n_33222), .CD(n_61405), .Q(to_acu2
		[73]));
	notech_mux2 i_39275(.S(n_54188), .A(to_acu2[73]), .B(n_2013), .Z(n_33222
		));
	notech_and4 i_878(.A(n_3015), .B(n_230891155), .C(n_230191148), .D(n_3013
		), .Z(n_230591152));
	notech_reg to_acu2_reg_74(.CP(n_61935), .D(n_33228), .CD(n_61405), .Q(to_acu2
		[74]));
	notech_mux2 i_39283(.S(n_54188), .A(to_acu2[74]), .B(n_2007), .Z(n_33228
		));
	notech_nao3 i_875(.A(n_2156), .B(in128[18]), .C(n_53815), .Z(n_230491151
		));
	notech_reg to_acu2_reg_75(.CP(n_61935), .D(n_33234), .CD(n_61405), .Q(to_acu2
		[75]));
	notech_mux2 i_39291(.S(n_54188), .A(to_acu2[75]), .B(n_2040), .Z(n_33234
		));
	notech_reg to_acu2_reg_76(.CP(n_61935), .D(n_33240), .CD(n_61405), .Q(to_acu2
		[76]));
	notech_mux2 i_39299(.S(n_54188), .A(to_acu2[76]), .B(n_2036), .Z(n_33240
		));
	notech_reg to_acu2_reg_77(.CP(n_61938), .D(n_33246), .CD(n_61390), .Q(to_acu2
		[77]));
	notech_mux2 i_39307(.S(n_54188), .A(to_acu2[77]), .B(n_2054), .Z(n_33246
		));
	notech_nao3 i_873(.A(n_2894), .B(in128[42]), .C(n_53797), .Z(n_230191148
		));
	notech_reg to_acu2_reg_78(.CP(n_61938), .D(n_33252), .CD(n_61374), .Q(to_acu2
		[78]));
	notech_mux2 i_39315(.S(n_54188), .A(to_acu2[78]), .B(n_2037), .Z(n_33252
		));
	notech_or4 i_165(.A(n_53824), .B(n_39845), .C(n_53797), .D(n_40008), .Z(n_230091147
		));
	notech_reg to_acu2_reg_79(.CP(n_61938), .D(n_33258), .CD(n_61374), .Q(to_acu2
		[79]));
	notech_mux2 i_39323(.S(n_54188), .A(to_acu2[79]), .B(n_2038), .Z(n_33258
		));
	notech_reg to_acu2_reg_80(.CP(n_61935), .D(n_33264), .CD(n_61374), .Q(to_acu2
		[80]));
	notech_mux2 i_39331(.S(n_54171), .A(to_acu2[80]), .B(n_2041), .Z(n_33264
		));
	notech_reg to_acu2_reg_81(.CP(n_61938), .D(n_33270), .CD(n_61374), .Q(to_acu2
		[81]));
	notech_mux2 i_39339(.S(n_54171), .A(to_acu2[81]), .B(n_2048), .Z(n_33270
		));
	notech_and4 i_868(.A(n_3010), .B(n_230091147), .C(n_229391140), .D(n_3008
		), .Z(n_229791144));
	notech_reg to_acu2_reg_82(.CP(n_61935), .D(n_33276), .CD(n_61374), .Q(to_acu2
		[82]));
	notech_mux2 i_39347(.S(n_54171), .A(to_acu2[82]), .B(n_2047), .Z(n_33276
		));
	notech_nao3 i_865(.A(n_2156), .B(in128[17]), .C(n_53815), .Z(n_229691143
		));
	notech_reg to_acu2_reg_83(.CP(n_61935), .D(n_33282), .CD(n_61377), .Q(to_acu2
		[83]));
	notech_mux2 i_39355(.S(n_54188), .A(to_acu2[83]), .B(n_2002), .Z(n_33282
		));
	notech_reg to_acu2_reg_84(.CP(n_61935), .D(n_33288), .CD(n_61377), .Q(to_acu2
		[84]));
	notech_mux2 i_39363(.S(n_54188), .A(to_acu2[84]), .B(n_47603), .Z(n_33288
		));
	notech_reg to_acu2_reg_85(.CP(n_61935), .D(n_33294), .CD(n_61377), .Q(to_acu2
		[85]));
	notech_mux2 i_39371(.S(n_54188), .A(to_acu2[85]), .B(n_2027), .Z(n_33294
		));
	notech_nao3 i_863(.A(n_2894), .B(in128[41]), .C(n_53797), .Z(n_229391140
		));
	notech_reg to_acu2_reg_86(.CP(n_61935), .D(n_33300), .CD(n_61377), .Q(to_acu2
		[86]));
	notech_mux2 i_39379(.S(n_54176), .A(to_acu2[86]), .B(n_2053), .Z(n_33300
		));
	notech_or4 i_160(.A(n_53824), .B(n_39845), .C(n_53797), .D(n_40007), .Z(n_229291139
		));
	notech_reg to_acu2_reg_87(.CP(n_61935), .D(n_33306), .CD(n_61377), .Q(to_acu2
		[87]));
	notech_mux2 i_39387(.S(n_54176), .A(to_acu2[87]), .B(n_2052), .Z(n_33306
		));
	notech_reg to_acu2_reg_88(.CP(n_61935), .D(n_33312), .CD(n_61374), .Q(to_acu2
		[88]));
	notech_mux2 i_39395(.S(n_54176), .A(to_acu2[88]), .B(n_2051), .Z(n_33312
		));
	notech_reg to_acu2_reg_89(.CP(n_61935), .D(n_33318), .CD(n_61374), .Q(to_acu2
		[89]));
	notech_mux2 i_39403(.S(n_54176), .A(to_acu2[89]), .B(n_2050), .Z(n_33318
		));
	notech_and4 i_858(.A(n_3005), .B(n_229291139), .C(n_228591132), .D(n_3003
		), .Z(n_228991136));
	notech_reg to_acu2_reg_90(.CP(n_61935), .D(n_33324), .CD(n_61374), .Q(to_acu2
		[90]));
	notech_mux2 i_39411(.S(n_54176), .A(to_acu2[90]), .B(n_2049), .Z(n_33324
		));
	notech_nao3 i_855(.A(n_2156), .B(in128[16]), .C(n_53815), .Z(n_228891135
		));
	notech_reg to_acu2_reg_91(.CP(n_61935), .D(n_33330), .CD(n_61374), .Q(to_acu2
		[91]));
	notech_mux2 i_39419(.S(n_54176), .A(to_acu2[91]), .B(n_2016), .Z(n_33330
		));
	notech_reg to_acu2_reg_92(.CP(n_61935), .D(n_33336), .CD(n_61374), .Q(to_acu2
		[92]));
	notech_mux2 i_39427(.S(n_54176), .A(to_acu2[92]), .B(n_2014), .Z(n_33336
		));
	notech_reg to_acu2_reg_93(.CP(n_61938), .D(n_33342), .CD(n_61374), .Q(to_acu2
		[93]));
	notech_mux2 i_39435(.S(n_54176), .A(to_acu2[93]), .B(n_2032), .Z(n_33342
		));
	notech_nao3 i_853(.A(n_2894), .B(in128[40]), .C(n_53797), .Z(n_228591132
		));
	notech_reg to_acu2_reg_94(.CP(n_61938), .D(n_33348), .CD(n_61374), .Q(to_acu2
		[94]));
	notech_mux2 i_39443(.S(n_54176), .A(to_acu2[94]), .B(n_1998), .Z(n_33348
		));
	notech_nand2 i_158(.A(n_2914), .B(in128[23]), .Z(n_228491131));
	notech_reg to_acu2_reg_95(.CP(n_61938), .D(n_33354), .CD(n_61374), .Q(to_acu2
		[95]));
	notech_mux2 i_39451(.S(n_54177), .A(to_acu2[95]), .B(n_2000), .Z(n_33354
		));
	notech_reg to_acu2_reg_96(.CP(n_61938), .D(n_33360), .CD(n_61374), .Q(to_acu2
		[96]));
	notech_mux2 i_39459(.S(n_54176), .A(to_acu2[96]), .B(n_2004), .Z(n_33360
		));
	notech_reg to_acu2_reg_97(.CP(n_61938), .D(n_33366), .CD(n_61374), .Q(to_acu2
		[97]));
	notech_mux2 i_39467(.S(n_54176), .A(to_acu2[97]), .B(n_2015), .Z(n_33366
		));
	notech_and4 i_848(.A(n_3000), .B(n_228491131), .C(n_227791124), .D(n_2998
		), .Z(n_228191128));
	notech_reg to_acu2_reg_98(.CP(n_61940), .D(n_33372), .CD(n_61374), .Q(to_acu2
		[98]));
	notech_mux2 i_39475(.S(n_54176), .A(to_acu2[98]), .B(n_1999), .Z(n_33372
		));
	notech_or4 i_842(.A(n_2154), .B(n_2153), .C(n_39845), .D(n_40006), .Z(n_228091127
		));
	notech_reg to_acu2_reg_99(.CP(n_61940), .D(n_33378), .CD(n_61377), .Q(to_acu2
		[99]));
	notech_mux2 i_39483(.S(n_54171), .A(to_acu2[99]), .B(n_2028), .Z(n_33378
		));
	notech_reg to_acu2_reg_100(.CP(n_61940), .D(n_33384), .CD(n_61379), .Q(to_acu2
		[100]));
	notech_mux2 i_39491(.S(n_54171), .A(to_acu2[100]), .B(n_2005), .Z(n_33384
		));
	notech_reg to_acu2_reg_101(.CP(n_61940), .D(n_33390), .CD(n_61377), .Q(to_acu2
		[101]));
	notech_mux2 i_39499(.S(n_54176), .A(to_acu2[101]), .B(n_2011), .Z(n_33390
		));
	notech_nao3 i_843(.A(n_53824), .B(in128[39]), .C(n_39845), .Z(n_227791124
		));
	notech_reg to_acu2_reg_102(.CP(n_61940), .D(n_33396), .CD(n_61377), .Q(to_acu2
		[102]));
	notech_mux2 i_39507(.S(n_54171), .A(to_acu2[102]), .B(n_2006), .Z(n_33396
		));
	notech_nand2 i_143(.A(n_2914), .B(in128[22]), .Z(n_227691123));
	notech_reg to_acu2_reg_103(.CP(n_61938), .D(n_33402), .CD(n_61377), .Q(to_acu2
		[103]));
	notech_mux2 i_39515(.S(n_54171), .A(to_acu2[103]), .B(n_2026), .Z(n_33402
		));
	notech_reg to_acu2_reg_104(.CP(n_61938), .D(n_33408), .CD(n_61379), .Q(to_acu2
		[104]));
	notech_mux2 i_39523(.S(n_54171), .A(to_acu2[104]), .B(n_2001), .Z(n_33408
		));
	notech_reg to_acu2_reg_105(.CP(n_61938), .D(n_33414), .CD(n_61379), .Q(to_acu2
		[105]));
	notech_mux2 i_39531(.S(n_54176), .A(to_acu2[105]), .B(n_2018), .Z(n_33414
		));
	notech_and4 i_838(.A(n_2995), .B(n_227691123), .C(n_226993350), .D(n_2993
		), .Z(n_227393346));
	notech_reg to_acu2_reg_106(.CP(n_61938), .D(n_33420), .CD(n_61379), .Q(to_acu2
		[106]));
	notech_mux2 i_39539(.S(n_54176), .A(to_acu2[106]), .B(n_2031), .Z(n_33420
		));
	notech_or4 i_832(.A(n_2154), .B(n_2153), .C(n_39845), .D(n_40005), .Z(n_227293347
		));
	notech_reg to_acu2_reg_107(.CP(n_61938), .D(n_33426), .CD(n_61379), .Q(to_acu2
		[107]));
	notech_mux2 i_39547(.S(n_54176), .A(to_acu2[107]), .B(n_1997), .Z(n_33426
		));
	notech_reg to_acu2_reg_108(.CP(n_61938), .D(n_33432), .CD(n_61379), .Q(to_acu2
		[108]));
	notech_mux2 i_39555(.S(n_54176), .A(to_acu2[108]), .B(n_2017), .Z(n_33432
		));
	notech_reg to_acu2_reg_109(.CP(n_61938), .D(n_33438), .CD(n_61377), .Q(to_acu2
		[109]));
	notech_mux2 i_39563(.S(n_54176), .A(to_acu2[109]), .B(n_2003), .Z(n_33438
		));
	notech_nao3 i_833(.A(n_53824), .B(in128[38]), .C(n_39845), .Z(n_226993350
		));
	notech_reg to_acu2_reg_110(.CP(n_61938), .D(n_33444), .CD(n_61377), .Q(to_acu2
		[110]));
	notech_mux2 i_39571(.S(n_54176), .A(to_acu2[110]), .B(n_2030), .Z(n_33444
		));
	notech_nand2 i_137(.A(n_2914), .B(in128[21]), .Z(n_226893351));
	notech_reg to_acu2_reg_111(.CP(n_61938), .D(n_33450), .CD(n_61377), .Q(to_acu2
		[111]));
	notech_mux2 i_39579(.S(n_54176), .A(to_acu2[111]), .B(n_2029), .Z(n_33450
		));
	notech_reg to_acu2_reg_112(.CP(n_61938), .D(n_33456), .CD(n_61377), .Q(to_acu2
		[112]));
	notech_mux2 i_39587(.S(n_54177), .A(to_acu2[112]), .B(n_3492), .Z(n_33456
		));
	notech_reg to_acu2_reg_113(.CP(n_61938), .D(n_33462), .CD(n_61377), .Q(to_acu2
		[113]));
	notech_mux2 i_39595(.S(n_54182), .A(to_acu2[113]), .B(n_2009), .Z(n_33462
		));
	notech_and4 i_828(.A(n_2990), .B(n_226893351), .C(n_226193358), .D(n_2988
		), .Z(n_226593354));
	notech_reg to_acu2_reg_114(.CP(n_61935), .D(n_33468), .CD(n_61377), .Q(to_acu2
		[114]));
	notech_mux2 i_39603(.S(n_54182), .A(to_acu2[114]), .B(n_2019), .Z(n_33468
		));
	notech_or4 i_822(.A(n_2154), .B(n_2153), .C(n_53806), .D(n_40004), .Z(n_226493355
		));
	notech_reg to_acu2_reg_115(.CP(n_61930), .D(n_33474), .CD(n_61377), .Q(to_acu2
		[115]));
	notech_mux2 i_39611(.S(n_54182), .A(to_acu2[115]), .B(n_2024), .Z(n_33474
		));
	notech_reg to_acu2_reg_116(.CP(n_61930), .D(n_33480), .CD(n_61377), .Q(to_acu2
		[116]));
	notech_mux2 i_39619(.S(n_54177), .A(to_acu2[116]), .B(n_2025), .Z(n_33480
		));
	notech_reg to_acu2_reg_117(.CP(n_61930), .D(n_33486), .CD(n_61377), .Q(to_acu2
		[117]));
	notech_mux2 i_39627(.S(n_54177), .A(to_acu2[117]), .B(n_3695), .Z(n_33486
		));
	notech_nao3 i_823(.A(n_53824), .B(in128[37]), .C(n_53806), .Z(n_226193358
		));
	notech_reg to_acu2_reg_118(.CP(n_61930), .D(n_33492), .CD(n_61377), .Q(to_acu2
		[118]));
	notech_mux2 i_39635(.S(n_54182), .A(to_acu2[118]), .B(n_2020), .Z(n_33492
		));
	notech_nand2 i_133(.A(n_2914), .B(in128[20]), .Z(n_226093359));
	notech_reg to_acu2_reg_119(.CP(n_61930), .D(n_33498), .CD(n_61377), .Q(to_acu2
		[119]));
	notech_mux2 i_39643(.S(n_54182), .A(to_acu2[119]), .B(n_3693), .Z(n_33498
		));
	notech_reg to_acu2_reg_120(.CP(n_61930), .D(n_33504), .CD(n_61369), .Q(to_acu2
		[120]));
	notech_mux2 i_39651(.S(n_54182), .A(to_acu2[120]), .B(n_2023), .Z(n_33504
		));
	notech_reg to_acu2_reg_121(.CP(n_61933), .D(n_33510), .CD(n_61369), .Q(to_acu2
		[121]));
	notech_mux2 i_39659(.S(n_54182), .A(to_acu2[121]), .B(n_2022), .Z(n_33510
		));
	notech_and4 i_818(.A(n_2985), .B(n_226093359), .C(n_225393366), .D(n_2983
		), .Z(n_225793362));
	notech_reg to_acu2_reg_122(.CP(n_61930), .D(n_33516), .CD(n_61369), .Q(to_acu2
		[122]));
	notech_mux2 i_39667(.S(n_54182), .A(to_acu2[122]), .B(n_2012), .Z(n_33516
		));
	notech_or4 i_812(.A(n_2154), .B(n_2153), .C(n_53806), .D(n_40003), .Z(n_225693363
		));
	notech_reg to_acu2_reg_123(.CP(n_61930), .D(n_33522), .CD(n_61369), .Q(to_acu2
		[123]));
	notech_mux2 i_39675(.S(n_54182), .A(to_acu2[123]), .B(n_3490), .Z(n_33522
		));
	notech_reg to_acu2_reg_124(.CP(n_61930), .D(n_33528), .CD(n_61369), .Q(to_acu2
		[124]));
	notech_mux2 i_39683(.S(n_54182), .A(to_acu2[124]), .B(n_3488), .Z(n_33528
		));
	notech_reg to_acu2_reg_125(.CP(n_61930), .D(n_33534), .CD(n_61372), .Q(to_acu2
		[125]));
	notech_mux2 i_39691(.S(n_54182), .A(to_acu2[125]), .B(n_2021), .Z(n_33534
		));
	notech_nao3 i_813(.A(n_53824), .B(in128[36]), .C(n_53806), .Z(n_225393366
		));
	notech_reg to_acu2_reg_126(.CP(n_61930), .D(n_33540), .CD(n_61372), .Q(to_acu2
		[126]));
	notech_mux2 i_39699(.S(n_54177), .A(to_acu2[126]), .B(n_3485), .Z(n_33540
		));
	notech_nand2 i_73(.A(n_2914), .B(in128[19]), .Z(n_225293367));
	notech_reg to_acu2_reg_127(.CP(n_61930), .D(n_33546), .CD(n_61372), .Q(to_acu2
		[127]));
	notech_mux2 i_39707(.S(n_54177), .A(to_acu2[127]), .B(n_3483), .Z(n_33546
		));
	notech_reg to_acu2_reg_128(.CP(n_61930), .D(n_33552), .CD(n_61369), .Q(to_acu2
		[128]));
	notech_mux2 i_39715(.S(n_54177), .A(to_acu2[128]), .B(n_3687), .Z(n_33552
		));
	notech_reg to_acu2_reg_129(.CP(n_61930), .D(n_33558), .CD(n_61369), .Q(to_acu2
		[129]));
	notech_mux2 i_39723(.S(n_54177), .A(to_acu2[129]), .B(n_2008), .Z(n_33558
		));
	notech_and4 i_808(.A(n_2980), .B(n_225293367), .C(n_224593374), .D(n_2978
		), .Z(n_224993370));
	notech_reg to_acu2_reg_130(.CP(n_61930), .D(n_33564), .CD(n_61369), .Q(to_acu2
		[130]));
	notech_mux2 i_39731(.S(n_54177), .A(to_acu2[130]), .B(n_3685), .Z(n_33564
		));
	notech_or4 i_802(.A(n_2154), .B(n_2153), .C(n_53806), .D(n_40002), .Z(n_224893371
		));
	notech_reg to_acu2_reg_131(.CP(n_61930), .D(n_33570), .CD(n_61369), .Q(to_acu2
		[131]));
	notech_mux2 i_39739(.S(n_54177), .A(to_acu2[131]), .B(n_3683), .Z(n_33570
		));
	notech_reg to_acu2_reg_132(.CP(n_61930), .D(n_33576), .CD(n_61369), .Q(to_acu2
		[132]));
	notech_mux2 i_39747(.S(n_54177), .A(to_acu2[132]), .B(n_3681), .Z(n_33576
		));
	notech_reg to_acu2_reg_133(.CP(n_61930), .D(n_33582), .CD(n_61369), .Q(to_acu2
		[133]));
	notech_mux2 i_39755(.S(n_54177), .A(to_acu2[133]), .B(n_3679), .Z(n_33582
		));
	notech_nao3 i_803(.A(n_53824), .B(in128[35]), .C(n_53806), .Z(n_224593374
		));
	notech_reg to_acu2_reg_134(.CP(n_61930), .D(n_33588), .CD(n_61369), .Q(to_acu2
		[134]));
	notech_mux2 i_39763(.S(n_54177), .A(to_acu2[134]), .B(n_3677), .Z(n_33588
		));
	notech_nand2 i_62(.A(n_2914), .B(in128[18]), .Z(n_224493375));
	notech_reg to_acu2_reg_135(.CP(n_61930), .D(n_33594), .CD(n_61369), .Q(to_acu2
		[135]));
	notech_mux2 i_39771(.S(n_54177), .A(to_acu2[135]), .B(n_3675), .Z(n_33594
		));
	notech_reg to_acu2_reg_136(.CP(n_61933), .D(n_33600), .CD(n_61369), .Q(to_acu2
		[136]));
	notech_mux2 i_39779(.S(n_54177), .A(to_acu2[136]), .B(n_3673), .Z(n_33600
		));
	notech_reg to_acu2_reg_137(.CP(n_61933), .D(n_33606), .CD(n_61369), .Q(to_acu2
		[137]));
	notech_mux2 i_39787(.S(n_54177), .A(to_acu2[137]), .B(n_3249), .Z(n_33606
		));
	notech_and4 i_798(.A(n_2975), .B(n_224493375), .C(n_223793382), .D(n_2973
		), .Z(n_224193378));
	notech_reg to_acu2_reg_138(.CP(n_61933), .D(n_33612), .CD(n_61369), .Q(to_acu2
		[138]));
	notech_mux2 i_39795(.S(n_54177), .A(to_acu2[138]), .B(n_3481), .Z(n_33612
		));
	notech_or4 i_792(.A(n_2154), .B(n_2153), .C(n_53806), .D(n_40001), .Z(n_224093379
		));
	notech_reg to_acu2_reg_139(.CP(n_61933), .D(n_33618), .CD(n_61369), .Q(to_acu2
		[139]));
	notech_mux2 i_39803(.S(n_54198), .A(to_acu2[139]), .B(n_3671), .Z(n_33618
		));
	notech_reg to_acu2_reg_140(.CP(n_61933), .D(n_33624), .CD(n_61369), .Q(to_acu2
		[140]));
	notech_mux2 i_39811(.S(n_54211), .A(to_acu2[140]), .B(n_3669), .Z(n_33624
		));
	notech_reg to_acu2_reg_141(.CP(n_61935), .D(n_33630), .CD(n_61372), .Q(to_acu2
		[141]));
	notech_mux2 i_39819(.S(n_54211), .A(to_acu2[141]), .B(n_3667), .Z(n_33630
		));
	notech_nao3 i_793(.A(n_53824), .B(in128[34]), .C(n_53806), .Z(n_223793382
		));
	notech_reg to_acu2_reg_142(.CP(n_61935), .D(n_33636), .CD(n_61372), .Q(to_acu2
		[142]));
	notech_mux2 i_39827(.S(n_54211), .A(to_acu2[142]), .B(n_3665), .Z(n_33636
		));
	notech_nand2 i_59(.A(n_2914), .B(in128[17]), .Z(n_223693383));
	notech_reg to_acu2_reg_143(.CP(n_61933), .D(n_33642), .CD(n_61372), .Q(to_acu2
		[143]));
	notech_mux2 i_39835(.S(n_54211), .A(to_acu2[143]), .B(n_3663), .Z(n_33642
		));
	notech_reg to_acu2_reg_144(.CP(n_61933), .D(n_33648), .CD(n_61372), .Q(to_acu2
		[144]));
	notech_mux2 i_39843(.S(n_54211), .A(to_acu2[144]), .B(n_3661), .Z(n_33648
		));
	notech_reg to_acu2_reg_145(.CP(n_61933), .D(n_33654), .CD(n_61372), .Q(to_acu2
		[145]));
	notech_mux2 i_39851(.S(n_54211), .A(to_acu2[145]), .B(n_3659), .Z(n_33654
		));
	notech_and4 i_788(.A(n_2970), .B(n_223693383), .C(n_2229), .D(n_2968), .Z
		(n_223393386));
	notech_reg to_acu2_reg_146(.CP(n_61933), .D(n_33660), .CD(n_61374), .Q(to_acu2
		[146]));
	notech_mux2 i_39859(.S(n_54211), .A(to_acu2[146]), .B(n_3479), .Z(n_33660
		));
	notech_or4 i_782(.A(n_2154), .B(n_2153), .C(n_53806), .D(n_40000), .Z(n_223293387
		));
	notech_reg to_acu2_reg_147(.CP(n_61933), .D(n_33666), .CD(n_61374), .Q(to_acu2
		[147]));
	notech_mux2 i_39867(.S(n_54211), .A(to_acu2[147]), .B(n_3657), .Z(n_33666
		));
	notech_reg to_acu2_reg_148(.CP(n_61933), .D(n_33672), .CD(n_61374), .Q(to_acu2
		[148]));
	notech_mux2 i_39875(.S(n_54211), .A(to_acu2[148]), .B(n_3655), .Z(n_33672
		));
	notech_reg to_acu2_reg_149(.CP(n_61933), .D(n_33678), .CD(n_61372), .Q(to_acu2
		[149]));
	notech_mux2 i_39883(.S(n_54211), .A(to_acu2[149]), .B(n_3653), .Z(n_33678
		));
	notech_nao3 i_783(.A(n_53824), .B(in128[33]), .C(n_39845), .Z(n_2229));
	notech_reg to_acu2_reg_150(.CP(n_61933), .D(n_33684), .CD(n_61374), .Q(to_acu2
		[150]));
	notech_mux2 i_39891(.S(n_54211), .A(to_acu2[150]), .B(n_3651), .Z(n_33684
		));
	notech_nand2 i_56(.A(n_2914), .B(in128[16]), .Z(n_2228));
	notech_reg to_acu2_reg_151(.CP(n_61933), .D(n_33690), .CD(n_61372), .Q(to_acu2
		[151]));
	notech_mux2 i_39899(.S(n_54211), .A(to_acu2[151]), .B(n_3649), .Z(n_33690
		));
	notech_reg to_acu2_reg_152(.CP(n_61933), .D(n_33696), .CD(n_61372), .Q(to_acu2
		[152]));
	notech_mux2 i_39907(.S(n_54211), .A(to_acu2[152]), .B(n_3647), .Z(n_33696
		));
	notech_reg to_acu2_reg_153(.CP(n_61933), .D(n_33702), .CD(n_61372), .Q(to_acu2
		[153]));
	notech_mux2 i_39915(.S(n_54210), .A(to_acu2[153]), .B(n_3645), .Z(n_33702
		));
	notech_and4 i_778(.A(n_2965), .B(n_2228), .C(n_2221), .D(n_2963), .Z(n_2225
		));
	notech_reg to_acu2_reg_154(.CP(n_61933), .D(n_33708), .CD(n_61372), .Q(to_acu2
		[154]));
	notech_mux2 i_39923(.S(n_54210), .A(to_acu2[154]), .B(n_3643), .Z(n_33708
		));
	notech_or4 i_772(.A(n_53806), .B(n_2154), .C(n_2153), .D(n_39999), .Z(n_2224
		));
	notech_reg to_acu2_reg_155(.CP(n_61933), .D(n_33714), .CD(n_61372), .Q(to_acu2
		[155]));
	notech_mux2 i_39931(.S(n_54210), .A(to_acu2[155]), .B(n_3641), .Z(n_33714
		));
	notech_reg to_acu2_reg_156(.CP(n_61933), .D(n_33720), .CD(n_61372), .Q(to_acu2
		[156]));
	notech_mux2 i_39939(.S(n_54210), .A(to_acu2[156]), .B(n_3639), .Z(n_33720
		));
	notech_reg to_acu2_reg_157(.CP(n_61949), .D(n_33726), .CD(n_61372), .Q(to_acu2
		[157]));
	notech_mux2 i_39947(.S(n_54210), .A(to_acu2[157]), .B(n_3637), .Z(n_33726
		));
	notech_nao3 i_773(.A(n_53824), .B(in128[32]), .C(n_53806), .Z(n_2221));
	notech_reg to_acu2_reg_158(.CP(n_61949), .D(n_33732), .CD(n_61372), .Q(to_acu2
		[158]));
	notech_mux2 i_39955(.S(n_54210), .A(to_acu2[158]), .B(n_3635), .Z(n_33732
		));
	notech_nao3 i_135(.A(n_40212), .B(n_40147), .C(n_2219), .Z(n_2220));
	notech_reg to_acu2_reg_159(.CP(n_61949), .D(n_33738), .CD(n_61372), .Q(to_acu2
		[159]));
	notech_mux2 i_39963(.S(n_54210), .A(to_acu2[159]), .B(n_3633), .Z(n_33738
		));
	notech_and4 i_705(.A(n_39992), .B(\to_acu2_0[7] ), .C(in128[18]), .D(in128
		[16]), .Z(n_2219));
	notech_reg to_acu2_reg_160(.CP(n_61946), .D(n_33744), .CD(n_61372), .Q(to_acu2
		[160]));
	notech_mux2 i_39971(.S(n_54211), .A(to_acu2[160]), .B(n_3631), .Z(n_33744
		));
	notech_and2 i_209(.A(n_40212), .B(n_40147), .Z(n_2218));
	notech_reg to_acu2_reg_161(.CP(n_61949), .D(n_33750), .CD(n_61372), .Q(to_acu2
		[161]));
	notech_mux2 i_39979(.S(n_54211), .A(to_acu2[161]), .B(n_3629), .Z(n_33750
		));
	notech_or4 i_6351(.A(int_excl[5]), .B(n_260791454), .C(n_2142), .D(n_2882
		), .Z(n_2217));
	notech_reg to_acu2_reg_162(.CP(n_61949), .D(n_33756), .CD(n_61379), .Q(to_acu2
		[162]));
	notech_mux2 i_39987(.S(n_54211), .A(to_acu2[162]), .B(n_3627), .Z(n_33756
		));
	notech_reg to_acu2_reg_163(.CP(n_61949), .D(n_33762), .CD(n_61388), .Q(to_acu2
		[163]));
	notech_mux2 i_39995(.S(n_54210), .A(to_acu2[163]), .B(n_3477), .Z(n_33762
		));
	notech_reg to_acu2_reg_164(.CP(n_61949), .D(n_33768), .CD(n_61388), .Q(to_acu2
		[164]));
	notech_mux2 i_40003(.S(n_54211), .A(to_acu2[164]), .B(n_3475), .Z(n_33768
		));
	notech_and3 i_65834(.A(n_2210), .B(n_2950), .C(n_2077), .Z(n_2214));
	notech_reg to_acu2_reg_165(.CP(n_61949), .D(n_33774), .CD(n_61388), .Q(to_acu2
		[165]));
	notech_mux2 i_40011(.S(n_54211), .A(to_acu2[165]), .B(n_3473), .Z(n_33774
		));
	notech_reg to_acu2_reg_166(.CP(n_61949), .D(n_33780), .CD(n_61388), .Q(to_acu2
		[166]));
	notech_mux2 i_40019(.S(n_54216), .A(to_acu2[166]), .B(n_3471), .Z(n_33780
		));
	notech_nand2 i_387(.A(n_2211), .B(\to_acu2_0[26] ), .Z(n_2212));
	notech_reg to_acu2_reg_167(.CP(n_61946), .D(n_33786), .CD(n_61388), .Q(to_acu2
		[167]));
	notech_mux2 i_40027(.S(n_54221), .A(to_acu2[167]), .B(n_3469), .Z(n_33786
		));
	notech_nand2 i_693(.A(n_40159), .B(n_40186), .Z(n_2211));
	notech_reg to_acu2_reg_168(.CP(n_61946), .D(n_33792), .CD(n_61388), .Q(to_acu2
		[168]));
	notech_mux2 i_40035(.S(n_54221), .A(to_acu2[168]), .B(n_3467), .Z(n_33792
		));
	notech_nand2 i_386(.A(\to_acu2_0[18] ), .B(\to_acu2_0[17] ), .Z(n_2210)
		);
	notech_reg to_acu2_reg_169(.CP(n_61946), .D(n_33798), .CD(n_61388), .Q(to_acu2
		[169]));
	notech_mux2 i_40043(.S(n_54221), .A(to_acu2[169]), .B(n_3250), .Z(n_33798
		));
	notech_nand2 i_687(.A(n_40150), .B(n_40149), .Z(n_2209));
	notech_reg to_acu2_reg_170(.CP(n_61946), .D(n_33804), .CD(n_61388), .Q(to_acu2
		[170]));
	notech_mux2 i_40051(.S(n_54221), .A(to_acu2[170]), .B(n_3619), .Z(n_33804
		));
	notech_nao3 i_51(.A(n_2175), .B(in128[27]), .C(n_2898), .Z(n_2208));
	notech_reg to_acu2_reg_171(.CP(n_61946), .D(n_33810), .CD(n_61388), .Q(to_acu2
		[171]));
	notech_mux2 i_40059(.S(n_54221), .A(to_acu2[171]), .B(n_3617), .Z(n_33810
		));
	notech_ao4 i_52(.A(n_2928), .B(n_40050), .C(n_2929), .D(n_40034), .Z(n_2207
		));
	notech_reg to_acu2_reg_172(.CP(n_61946), .D(n_33816), .CD(n_61388), .Q(to_acu2
		[172]));
	notech_mux2 i_40067(.S(n_54221), .A(to_acu2[172]), .B(n_3465), .Z(n_33816
		));
	notech_and4 i_637(.A(n_2207), .B(n_2199), .C(n_2208), .D(n_2944), .Z(n_2206
		));
	notech_reg to_acu2_reg_173(.CP(n_61946), .D(n_33822), .CD(n_61385), .Q(to_acu2
		[173]));
	notech_mux2 i_40075(.S(n_54221), .A(to_acu2[173]), .B(n_3463), .Z(n_33822
		));
	notech_reg to_acu2_reg_174(.CP(n_61946), .D(n_33828), .CD(n_61385), .Q(to_acu2
		[174]));
	notech_mux2 i_40083(.S(n_54221), .A(to_acu2[174]), .B(n_3613), .Z(n_33828
		));
	notech_reg to_acu2_reg_175(.CP(n_61946), .D(n_33834), .CD(n_61385), .Q(to_acu2
		[175]));
	notech_mux2 i_40091(.S(n_54221), .A(to_acu2[175]), .B(n_3461), .Z(n_33834
		));
	notech_reg to_acu2_reg_176(.CP(n_61946), .D(n_33840), .CD(n_61385), .Q(to_acu2
		[176]));
	notech_mux2 i_40099(.S(n_54221), .A(to_acu2[176]), .B(n_3610), .Z(n_33840
		));
	notech_or2 i_628(.A(n_2922), .B(n_40026), .Z(n_2202));
	notech_reg to_acu2_reg_177(.CP(n_61946), .D(n_33846), .CD(n_61385), .Q(to_acu2
		[177]));
	notech_mux2 i_40107(.S(n_54221), .A(to_acu2[177]), .B(n_3608), .Z(n_33846
		));
	notech_reg to_acu2_reg_178(.CP(n_61951), .D(n_33852), .CD(n_61385), .Q(to_acu2
		[178]));
	notech_mux2 i_40115(.S(n_54221), .A(to_acu2[178]), .B(n_3459), .Z(n_33852
		));
	notech_reg to_acu2_reg_179(.CP(n_61951), .D(n_33858), .CD(n_61385), .Q(to_acu2
		[179]));
	notech_mux2 i_40123(.S(n_54221), .A(to_acu2[179]), .B(n_3605), .Z(n_33858
		));
	notech_or2 i_630(.A(n_2921), .B(n_40018), .Z(n_2199));
	notech_reg to_acu2_reg_180(.CP(n_61951), .D(n_33864), .CD(n_61385), .Q(to_acu2
		[180]));
	notech_mux2 i_40131(.S(n_54216), .A(to_acu2[180]), .B(n_3603), .Z(n_33864
		));
	notech_nao3 i_48(.A(n_2175), .B(in128[26]), .C(n_53815), .Z(n_2198));
	notech_reg to_acu2_reg_181(.CP(n_61951), .D(n_33870), .CD(n_61385), .Q(to_acu2
		[181]));
	notech_mux2 i_40139(.S(n_54216), .A(to_acu2[181]), .B(n_3601), .Z(n_33870
		));
	notech_ao4 i_49(.A(n_2928), .B(n_40049), .C(n_2929), .D(n_40033), .Z(n_2197
		));
	notech_reg to_acu2_reg_182(.CP(n_61951), .D(n_33876), .CD(n_61385), .Q(to_acu2
		[182]));
	notech_mux2 i_40147(.S(n_54216), .A(to_acu2[182]), .B(n_3599), .Z(n_33876
		));
	notech_and4 i_625(.A(n_2197), .B(n_2189), .C(n_2198), .D(n_2939), .Z(n_2196
		));
	notech_reg to_acu2_reg_183(.CP(n_61951), .D(n_33882), .CD(n_61385), .Q(to_acu2
		[183]));
	notech_mux2 i_40155(.S(n_54216), .A(to_acu2[183]), .B(n_3597), .Z(n_33882
		));
	notech_reg to_acu2_reg_184(.CP(n_61951), .D(n_33888), .CD(n_61390), .Q(to_acu2
		[184]));
	notech_mux2 i_40163(.S(n_54216), .A(to_acu2[184]), .B(n_3595), .Z(n_33888
		));
	notech_reg to_acu2_reg_185(.CP(n_61951), .D(n_33894), .CD(n_61390), .Q(to_acu2
		[185]));
	notech_mux2 i_40171(.S(n_54216), .A(to_acu2[185]), .B(n_3593), .Z(n_33894
		));
	notech_reg to_acu2_reg_186(.CP(n_61951), .D(n_33900), .CD(n_61390), .Q(to_acu2
		[186]));
	notech_mux2 i_40179(.S(n_54216), .A(to_acu2[186]), .B(n_3591), .Z(n_33900
		));
	notech_or2 i_616(.A(n_2922), .B(n_40025), .Z(n_2192));
	notech_reg to_acu2_reg_187(.CP(n_61951), .D(n_33906), .CD(n_61390), .Q(to_acu2
		[187]));
	notech_mux2 i_40187(.S(n_54216), .A(to_acu2[187]), .B(n_3589), .Z(n_33906
		));
	notech_reg to_acu2_reg_188(.CP(n_61949), .D(n_33912), .CD(n_61390), .Q(to_acu2
		[188]));
	notech_mux2 i_40195(.S(n_54221), .A(to_acu2[188]), .B(n_3587), .Z(n_33912
		));
	notech_reg to_acu2_reg_189(.CP(n_61949), .D(n_33918), .CD(n_61390), .Q(to_acu2
		[189]));
	notech_mux2 i_40203(.S(n_54221), .A(to_acu2[189]), .B(n_3585), .Z(n_33918
		));
	notech_or2 i_618(.A(n_2921), .B(n_40017), .Z(n_2189));
	notech_reg to_acu2_reg_190(.CP(n_61949), .D(n_33924), .CD(n_61390), .Q(to_acu2
		[190]));
	notech_mux2 i_40211(.S(n_54216), .A(to_acu2[190]), .B(n_3583), .Z(n_33924
		));
	notech_nao3 i_45(.A(n_2175), .B(in128[25]), .C(n_53815), .Z(n_2188));
	notech_reg to_acu2_reg_191(.CP(n_61949), .D(n_33930), .CD(n_61390), .Q(to_acu2
		[191]));
	notech_mux2 i_40219(.S(n_54216), .A(to_acu2[191]), .B(n_3581), .Z(n_33930
		));
	notech_ao4 i_46(.A(n_2928), .B(n_40048), .C(n_2929), .D(n_40032), .Z(n_2187
		));
	notech_reg to_acu2_reg_192(.CP(n_61949), .D(n_33936), .CD(n_61390), .Q(to_acu2
		[192]));
	notech_mux2 i_40227(.S(n_54216), .A(to_acu2[192]), .B(n_3579), .Z(n_33936
		));
	notech_and4 i_613(.A(n_2187), .B(n_2179), .C(n_2188), .D(n_2934), .Z(n_2186
		));
	notech_reg to_acu2_reg_193(.CP(n_61949), .D(n_33942), .CD(n_61390), .Q(to_acu2
		[193]));
	notech_mux2 i_40235(.S(n_54199), .A(to_acu2[193]), .B(n_3577), .Z(n_33942
		));
	notech_reg to_acu2_reg_194(.CP(n_61949), .D(n_33948), .CD(n_61390), .Q(to_acu2
		[194]));
	notech_mux2 i_40243(.S(n_54199), .A(to_acu2[194]), .B(n_3575), .Z(n_33948
		));
	notech_reg to_acu2_reg_195(.CP(n_61949), .D(n_33954), .CD(n_61388), .Q(to_acu2
		[195]));
	notech_mux2 i_40251(.S(n_54199), .A(to_acu2[195]), .B(n_3573), .Z(n_33954
		));
	notech_reg to_acu2_reg_196(.CP(n_61949), .D(n_33960), .CD(n_61388), .Q(to_acu2
		[196]));
	notech_mux2 i_40259(.S(n_54199), .A(to_acu2[196]), .B(n_3571), .Z(n_33960
		));
	notech_or2 i_604(.A(n_2922), .B(n_40024), .Z(n_2182));
	notech_reg to_acu2_reg_197(.CP(n_61949), .D(n_33966), .CD(n_61388), .Q(to_acu2
		[197]));
	notech_mux2 i_40267(.S(n_54199), .A(to_acu2[197]), .B(n_3457), .Z(n_33966
		));
	notech_reg to_acu2_reg_198(.CP(n_61949), .D(n_33972), .CD(n_61388), .Q(to_acu2
		[198]));
	notech_mux2 i_40275(.S(n_54199), .A(to_acu2[198]), .B(n_3455), .Z(n_33972
		));
	notech_reg to_acu2_reg_199(.CP(n_61946), .D(n_33978), .CD(n_61388), .Q(to_acu2
		[199]));
	notech_mux2 i_40283(.S(n_54199), .A(to_acu2[199]), .B(n_3453), .Z(n_33978
		));
	notech_or2 i_606(.A(n_2921), .B(n_40016), .Z(n_2179));
	notech_reg to_acu2_reg_200(.CP(n_61940), .D(n_33984), .CD(n_61388), .Q(to_acu2
		[200]));
	notech_mux2 i_40291(.S(n_54199), .A(to_acu2[200]), .B(n_3451), .Z(n_33984
		));
	notech_nao3 i_42(.A(n_2175), .B(in128[24]), .C(n_53815), .Z(n_2178));
	notech_reg to_acu2_reg_201(.CP(n_61944), .D(n_33990), .CD(n_61388), .Q(to_acu2
		[201]));
	notech_mux2 i_40299(.S(n_54199), .A(to_acu2[201]), .B(n_3565), .Z(n_33990
		));
	notech_ao4 i_43(.A(n_2928), .B(n_40047), .C(n_2929), .D(n_40031), .Z(n_2177
		));
	notech_reg to_acu2_reg_202(.CP(n_61940), .D(n_33996), .CD(n_61388), .Q(to_acu2
		[202]));
	notech_mux2 i_40307(.S(n_54199), .A(to_acu2[202]), .B(n_3449), .Z(n_33996
		));
	notech_and4 i_601(.A(n_2177), .B(n_2168), .C(n_2178), .D(n_2926), .Z(n_2176
		));
	notech_reg to_acu2_reg_203(.CP(n_61940), .D(n_34002), .CD(n_61388), .Q(to_acu2
		[203]));
	notech_mux2 i_40315(.S(n_54199), .A(to_acu2[203]), .B(n_3447), .Z(n_34002
		));
	notech_or2 i_600(.A(n_2884), .B(n_2900), .Z(n_2175));
	notech_reg to_acu2_reg_204(.CP(n_61940), .D(n_34008), .CD(n_61388), .Q(to_acu2
		[204]));
	notech_mux2 i_40323(.S(n_54199), .A(to_acu2[204]), .B(n_3561), .Z(n_34008
		));
	notech_reg to_acu2_reg_205(.CP(n_61944), .D(n_34014), .CD(n_61383), .Q(to_acu2
		[205]));
	notech_mux2 i_40331(.S(n_54199), .A(to_acu2[205]), .B(n_3559), .Z(n_34014
		));
	notech_reg to_acu2_reg_206(.CP(n_61944), .D(n_34020), .CD(n_61383), .Q(to_acu2
		[206]));
	notech_mux2 i_40339(.S(n_54198), .A(to_acu2[206]), .B(n_3557), .Z(n_34020
		));
	notech_reg to_acu2_reg_207(.CP(n_61944), .D(n_34026), .CD(n_61383), .Q(to_acu2
		[207]));
	notech_mux2 i_40347(.S(n_54198), .A(to_acu2[207]), .B(n_3445), .Z(n_34026
		));
	notech_or2 i_591(.A(n_2922), .B(n_40023), .Z(n_2171));
	notech_reg to_acu2_reg_208(.CP(n_61944), .D(n_34032), .CD(n_61379), .Q(to_acu2
		[208]));
	notech_mux2 i_40355(.S(n_54198), .A(to_acu2[208]), .B(n_3554), .Z(n_34032
		));
	notech_reg to_acu2_reg_209(.CP(n_61944), .D(n_34038), .CD(n_61379), .Q(to_acu2
		[209]));
	notech_mux2 i_40363(.S(n_54198), .A(to_acu2[209]), .B(n_3552), .Z(n_34038
		));
	notech_reg to_acu2_reg_210(.CP(n_61940), .D(n_34044), .CD(n_61383), .Q(to_acu2
		[210]));
	notech_mux2 i_40371(.S(n_54198), .A(to_acu2[210]), .B(n_48359), .Z(n_34044
		));
	notech_or2 i_593(.A(n_2921), .B(n_40015), .Z(n_2168));
	notech_reg to_acu1_reg_0(.CP(n_61940), .D(n_34050), .CD(n_61383), .Q(to_acu1
		[0]));
	notech_mux2 i_40379(.S(n_57672), .A(to_acu1[0]), .B(n_38878), .Z(n_34050
		));
	notech_or2 i_590(.A(n_2915), .B(n_2884), .Z(n_2167));
	notech_reg to_acu1_reg_1(.CP(n_61940), .D(n_34056), .CD(n_61383), .Q(to_acu1
		[1]));
	notech_mux2 i_40387(.S(n_57672), .A(to_acu1[1]), .B(n_39425), .Z(n_34056
		));
	notech_or4 i_40(.A(n_53824), .B(n_53806), .C(n_2885), .D(n_40014), .Z(n_2166
		));
	notech_reg to_acu1_reg_2(.CP(n_61940), .D(n_34062), .CD(n_61383), .Q(to_acu1
		[2]));
	notech_mux2 i_40395(.S(n_57672), .A(to_acu1[2]), .B(n_38880), .Z(n_34062
		));
	notech_reg to_acu1_reg_3(.CP(n_61940), .D(n_34068), .CD(n_61383), .Q(to_acu1
		[3]));
	notech_mux2 i_40403(.S(n_57667), .A(to_acu1[3]), .B(n_39429), .Z(n_34068
		));
	notech_reg to_acu1_reg_4(.CP(n_61940), .D(n_34074), .CD(n_61379), .Q(to_acu1
		[4]));
	notech_mux2 i_40411(.S(n_57667), .A(to_acu1[4]), .B(n_38881), .Z(n_34074
		));
	notech_and4 i_586(.A(n_2919), .B(n_2166), .C(n_2157), .D(n_2909), .Z(n_2163
		));
	notech_reg to_acu1_reg_5(.CP(n_61940), .D(n_34080), .CD(n_61379), .Q(to_acu1
		[5]));
	notech_mux2 i_40419(.S(n_57667), .A(to_acu1[5]), .B(n_39434), .Z(n_34080
		));
	notech_nao3 i_584(.A(n_53797), .B(n_39860), .C(imm_sz[1]), .Z(n_2162));
	notech_reg to_acu1_reg_6(.CP(n_61940), .D(n_34086), .CD(n_61379), .Q(to_acu1
		[6]));
	notech_mux2 i_40427(.S(n_57677), .A(to_acu1[6]), .B(n_39436), .Z(n_34086
		));
	notech_or2 i_583(.A(imm_sz[1]), .B(imm_sz[2]), .Z(n_2161));
	notech_reg to_acu1_reg_7(.CP(n_61940), .D(n_34092), .CD(n_61379), .Q(to_acu1
		[7]));
	notech_mux2 i_40435(.S(n_57678), .A(to_acu1[7]), .B(n_39439), .Z(n_34092
		));
	notech_nao3 i_579(.A(n_2156), .B(in128[23]), .C(n_53815), .Z(n_2160));
	notech_reg to_acu1_reg_8(.CP(n_61940), .D(n_34098), .CD(n_61379), .Q(to_acu1
		[8]));
	notech_mux2 i_40443(.S(n_57678), .A(to_acu1[8]), .B(n_38883), .Z(n_34098
		));
	notech_reg to_acu1_reg_9(.CP(n_61940), .D(n_34104), .CD(n_61379), .Q(to_acu1
		[9]));
	notech_mux2 i_40451(.S(n_57678), .A(to_acu1[9]), .B(n_39443), .Z(n_34104
		));
	notech_reg to_acu1_reg_10(.CP(n_61946), .D(n_34110), .CD(n_61379), .Q(to_acu1
		[10]));
	notech_mux2 i_40459(.S(n_57678), .A(to_acu1[10]), .B(n_39446), .Z(n_34110
		));
	notech_nao3 i_577(.A(n_2894), .B(in128[47]), .C(n_53797), .Z(n_2157));
	notech_reg to_acu1_reg_11(.CP(n_61946), .D(n_34116), .CD(n_61379), .Q(to_acu1
		[11]));
	notech_mux2 i_40467(.S(n_57678), .A(to_acu1[11]), .B(n_39448), .Z(n_34116
		));
	notech_nand2 i_575(.A(n_53797), .B(n_39843), .Z(n_2156));
	notech_reg to_acu1_reg_12(.CP(n_61944), .D(n_34122), .CD(n_61379), .Q(to_acu1
		[12]));
	notech_mux2 i_40475(.S(n_57678), .A(to_acu1[12]), .B(n_38885), .Z(n_34122
		));
	notech_nor2 i_630049(.A(imm_sz[0]), .B(n_2161), .Z(n_2155));
	notech_reg to_acu1_reg_13(.CP(n_61944), .D(n_34128), .CD(n_61379), .Q(to_acu1
		[13]));
	notech_mux2 i_40483(.S(n_57678), .A(to_acu1[13]), .B(n_38887), .Z(n_34128
		));
	notech_nor2 i_568(.A(displc[0]), .B(n_2886), .Z(n_2154));
	notech_reg to_acu1_reg_14(.CP(n_61944), .D(n_34134), .CD(n_61379), .Q(to_acu1
		[14]));
	notech_mux2 i_40491(.S(n_57678), .A(to_acu1[14]), .B(n_38889), .Z(n_34134
		));
	notech_and2 i_567(.A(displc[0]), .B(n_2886), .Z(n_2153));
	notech_reg to_acu1_reg_15(.CP(n_61946), .D(n_34140), .CD(n_61385), .Q(to_acu1
		[15]));
	notech_mux2 i_40499(.S(n_57678), .A(to_acu1[15]), .B(n_39457), .Z(n_34140
		));
	notech_reg to_acu1_reg_16(.CP(n_61946), .D(n_34146), .CD(n_61385), .Q(to_acu1
		[16]));
	notech_mux2 i_40507(.S(n_57678), .A(to_acu1[16]), .B(n_39459), .Z(n_34146
		));
	notech_reg to_acu1_reg_17(.CP(n_61946), .D(n_34152), .CD(n_61385), .Q(to_acu1
		[17]));
	notech_mux2 i_40515(.S(n_57678), .A(to_acu1[17]), .B(n_39462), .Z(n_34152
		));
	notech_reg to_acu1_reg_18(.CP(n_61946), .D(n_34158), .CD(n_61383), .Q(to_acu1
		[18]));
	notech_mux2 i_40523(.S(n_57678), .A(to_acu1[18]), .B(n_39464), .Z(n_34158
		));
	notech_reg to_acu1_reg_19(.CP(n_61946), .D(n_34164), .CD(n_61385), .Q(to_acu1
		[19]));
	notech_mux2 i_40531(.S(n_57678), .A(to_acu1[19]), .B(n_39467), .Z(n_34164
		));
	notech_reg to_acu1_reg_20(.CP(n_61944), .D(n_34170), .CD(n_61385), .Q(to_acu1
		[20]));
	notech_mux2 i_40539(.S(n_57677), .A(to_acu1[20]), .B(n_39469), .Z(n_34170
		));
	notech_reg to_acu1_reg_21(.CP(n_61944), .D(n_34176), .CD(n_61385), .Q(to_acu1
		[21]));
	notech_mux2 i_40547(.S(n_57677), .A(to_acu1[21]), .B(n_39472), .Z(n_34176
		));
	notech_and2 i_353(.A(n_40178), .B(n_39861), .Z(n_2146));
	notech_reg to_acu1_reg_22(.CP(n_61944), .D(n_34182), .CD(n_61385), .Q(to_acu1
		[22]));
	notech_mux2 i_40555(.S(n_57677), .A(to_acu1[22]), .B(n_38891), .Z(n_34182
		));
	notech_reg to_acu1_reg_23(.CP(n_61944), .D(n_34188), .CD(n_61385), .Q(to_acu1
		[23]));
	notech_mux2 i_40563(.S(n_57677), .A(to_acu1[23]), .B(n_38893), .Z(n_34188
		));
	notech_reg to_acu1_reg_24(.CP(n_61944), .D(n_34194), .CD(n_61385), .Q(to_acu1
		[24]));
	notech_mux2 i_40571(.S(n_57677), .A(to_acu1[24]), .B(n_38895), .Z(n_34194
		));
	notech_nor2 i_557(.A(imm_sz[0]), .B(imm_sz[2]), .Z(n_2143));
	notech_reg to_acu1_reg_25(.CP(n_61944), .D(n_34200), .CD(n_61383), .Q(to_acu1
		[25]));
	notech_mux2 i_40579(.S(n_57677), .A(to_acu1[25]), .B(n_38897), .Z(n_34200
		));
	notech_and4 i_389(.A(n_38625), .B(n_38624), .C(n_2878), .D(n_2877), .Z(n_2142
		));
	notech_reg to_acu1_reg_26(.CP(n_61944), .D(n_34206), .CD(n_61383), .Q(to_acu1
		[26]));
	notech_mux2 i_40587(.S(n_57677), .A(to_acu1[26]), .B(n_38898), .Z(n_34206
		));
	notech_nao3 i_140(.A(n_40193), .B(n_59607), .C(n_2833), .Z(n_2141));
	notech_reg to_acu1_reg_27(.CP(n_61944), .D(n_34212), .CD(n_61383), .Q(to_acu1
		[27]));
	notech_mux2 i_40595(.S(n_57677), .A(to_acu1[27]), .B(n_38900), .Z(n_34212
		));
	notech_ao4 i_37(.A(n_58712), .B(n_2873), .C(n_2136), .D(pc_req), .Z(n_2140
		));
	notech_reg to_acu1_reg_28(.CP(n_61944), .D(n_34218), .CD(n_61383), .Q(to_acu1
		[28]));
	notech_mux2 i_40603(.S(n_57677), .A(to_acu1[28]), .B(n_38902), .Z(n_34218
		));
	notech_reg to_acu1_reg_29(.CP(n_61944), .D(n_34224), .CD(n_61383), .Q(to_acu1
		[29]));
	notech_mux2 i_40611(.S(n_57677), .A(to_acu1[29]), .B(n_39488), .Z(n_34224
		));
	notech_ao3 i_3230191(.A(n_2117), .B(n_39990), .C(n_2114), .Z(n_2138));
	notech_reg to_acu1_reg_30(.CP(n_61944), .D(n_34230), .CD(n_61383), .Q(to_acu1
		[30]));
	notech_mux2 i_40619(.S(n_57677), .A(to_acu1[30]), .B(n_39491), .Z(n_34230
		));
	notech_reg to_acu1_reg_31(.CP(n_61881), .D(n_34236), .CD(n_61383), .Q(to_acu1
		[31]));
	notech_mux2 i_40627(.S(n_57677), .A(to_acu1[31]), .B(n_39493), .Z(n_34236
		));
	notech_mux2 i_38(.S(n_5408), .A(n_2134), .B(n_2132), .Z(n_2136));
	notech_reg to_acu1_reg_32(.CP(n_61814), .D(n_34242), .CD(n_61383), .Q(to_acu1
		[32]));
	notech_mux2 i_40635(.S(n_57677), .A(to_acu1[32]), .B(n_39496), .Z(n_34242
		));
	notech_reg to_acu1_reg_33(.CP(n_61814), .D(n_34248), .CD(n_61383), .Q(to_acu1
		[33]));
	notech_mux2 i_40643(.S(n_57609), .A(to_acu1[33]), .B(n_39498), .Z(n_34248
		));
	notech_and2 i_4231(.A(n_5415), .B(n_2071), .Z(n_2134));
	notech_reg to_acu1_reg_34(.CP(n_61814), .D(n_34254), .CD(n_61383), .Q(to_acu1
		[34]));
	notech_mux2 i_40651(.S(n_57609), .A(to_acu1[34]), .B(n_39501), .Z(n_34254
		));
	notech_reg to_acu1_reg_35(.CP(n_61814), .D(n_34260), .CD(n_61383), .Q(to_acu1
		[35]));
	notech_mux2 i_40659(.S(n_57609), .A(to_acu1[35]), .B(n_39503), .Z(n_34260
		));
	notech_nor2 i_65890(.A(n_2834), .B(n_38661), .Z(n_2132));
	notech_reg to_acu1_reg_36(.CP(n_61814), .D(n_34266), .CD(n_61253), .Q(to_acu1
		[36]));
	notech_mux2 i_40667(.S(n_57609), .A(to_acu1[36]), .B(n_39506), .Z(n_34266
		));
	notech_reg to_acu1_reg_37(.CP(n_61814), .D(n_34272), .CD(n_61253), .Q(to_acu1
		[37]));
	notech_mux2 i_40675(.S(n_57609), .A(to_acu1[37]), .B(n_39508), .Z(n_34272
		));
	notech_and4 i_70866(.A(n_2869), .B(n_58465), .C(n_2129), .D(n_2128), .Z(n_2130
		));
	notech_reg to_acu1_reg_38(.CP(n_61814), .D(n_34278), .CD(n_61253), .Q(to_acu1
		[38]));
	notech_mux2 i_40683(.S(n_57609), .A(to_acu1[38]), .B(n_39511), .Z(n_34278
		));
	notech_nand3 i_2516(.A(n_2124), .B(n_59607), .C(n_40193), .Z(n_2129));
	notech_reg to_acu1_reg_39(.CP(n_61814), .D(n_34284), .CD(n_61253), .Q(to_acu1
		[39]));
	notech_mux2 i_40691(.S(n_57610), .A(to_acu1[39]), .B(n_130392924), .Z(n_34284
		));
	notech_nand3 i_2843(.A(fpu), .B(n_2120), .C(n_2072), .Z(n_2128));
	notech_reg to_acu1_reg_40(.CP(n_61814), .D(n_34290), .CD(n_61253), .Q(to_acu1
		[40]));
	notech_mux2 i_40699(.S(n_57610), .A(to_acu1[40]), .B(n_39514), .Z(n_34290
		));
	notech_nand2 i_519(.A(n_2120), .B(n_2867), .Z(n_2127));
	notech_reg to_acu1_reg_41(.CP(n_61814), .D(n_34296), .CD(n_61253), .Q(to_acu1
		[41]));
	notech_mux2 i_40707(.S(n_57610), .A(to_acu1[41]), .B(n_39517), .Z(n_34296
		));
	notech_or4 i_517(.A(n_2834), .B(pg_fault), .C(pc_req), .D(fsm[1]), .Z(n_2126
		));
	notech_reg to_acu1_reg_42(.CP(n_61814), .D(n_34302), .CD(n_61253), .Q(to_acu1
		[42]));
	notech_mux2 i_40715(.S(n_57610), .A(to_acu1[42]), .B(n_39519), .Z(n_34302
		));
	notech_nand2 i_164(.A(n_1740), .B(n_2121), .Z(n_2125));
	notech_reg to_acu1_reg_43(.CP(n_61814), .D(n_34308), .CD(n_61253), .Q(to_acu1
		[43]));
	notech_mux2 i_40723(.S(n_57610), .A(to_acu1[43]), .B(n_39522), .Z(n_34308
		));
	notech_nand2 i_506(.A(n_38510), .B(n_2833), .Z(n_2124));
	notech_reg to_acu1_reg_44(.CP(n_61814), .D(n_34314), .CD(n_61253), .Q(to_acu1
		[44]));
	notech_mux2 i_40731(.S(n_57610), .A(to_acu1[44]), .B(n_39524), .Z(n_34314
		));
	notech_and2 i_213(.A(fpu), .B(n_2120), .Z(n_2123));
	notech_reg to_acu1_reg_45(.CP(n_61810), .D(n_34320), .CD(n_61253), .Q(to_acu1
		[45]));
	notech_mux2 i_40739(.S(n_57610), .A(to_acu1[45]), .B(n_39527), .Z(n_34320
		));
	notech_ao3 i_494(.A(n_40171), .B(\to_acu2_0[62] ), .C(twobyte), .Z(n_2122
		));
	notech_reg to_acu1_reg_46(.CP(n_61810), .D(n_34326), .CD(n_61253), .Q(to_acu1
		[46]));
	notech_mux2 i_40747(.S(n_57609), .A(to_acu1[46]), .B(n_39529), .Z(n_34326
		));
	notech_nao3 i_493(.A(n_40171), .B(\to_acu2_0[69] ), .C(twobyte), .Z(n_2121
		));
	notech_reg to_acu1_reg_47(.CP(n_61810), .D(n_34332), .CD(n_61249), .Q(to_acu1
		[47]));
	notech_mux2 i_40755(.S(n_57609), .A(to_acu1[47]), .B(n_39532), .Z(n_34332
		));
	notech_and4 i_28(.A(n_2119), .B(n_2850), .C(n_1476), .D(n_39847), .Z(n_2120
		));
	notech_reg to_acu1_reg_48(.CP(n_61814), .D(n_34338), .CD(n_61253), .Q(to_acu1
		[48]));
	notech_mux2 i_40763(.S(n_57609), .A(to_acu1[48]), .B(n_39534), .Z(n_34338
		));
	notech_or4 i_20(.A(valid_len[3]), .B(valid_len[4]), .C(n_2118), .D(n_2851
		), .Z(n_2119));
	notech_reg to_acu1_reg_49(.CP(n_61814), .D(n_34344), .CD(n_61249), .Q(to_acu1
		[49]));
	notech_mux2 i_40771(.S(n_57604), .A(to_acu1[49]), .B(n_39537), .Z(n_34344
		));
	notech_and2 i_479(.A(valid_len[0]), .B(valid_len[1]), .Z(n_2118));
	notech_reg to_acu1_reg_50(.CP(n_61814), .D(n_34350), .CD(n_61249), .Q(to_acu1
		[50]));
	notech_mux2 i_40779(.S(n_57609), .A(to_acu1[50]), .B(n_39539), .Z(n_34350
		));
	notech_nand2 i_473(.A(n_2838), .B(valid_len[4]), .Z(n_2117));
	notech_reg to_acu1_reg_51(.CP(n_61814), .D(n_34356), .CD(n_61249), .Q(to_acu1
		[51]));
	notech_mux2 i_40787(.S(n_57609), .A(to_acu1[51]), .B(n_39542), .Z(n_34356
		));
	notech_reg to_acu1_reg_52(.CP(n_61814), .D(n_34362), .CD(n_61253), .Q(to_acu1
		[52]));
	notech_mux2 i_40795(.S(n_57609), .A(to_acu1[52]), .B(n_39544), .Z(n_34362
		));
	notech_reg to_acu1_reg_53(.CP(n_61816), .D(n_34368), .CD(n_61253), .Q(to_acu1
		[53]));
	notech_mux2 i_40803(.S(n_57609), .A(to_acu1[53]), .B(n_39546), .Z(n_34368
		));
	notech_ao4 i_474(.A(n_2111), .B(n_2110), .C(valid_len[4]), .D(n_2838), .Z
		(n_2114));
	notech_reg to_acu1_reg_54(.CP(n_61816), .D(n_34374), .CD(n_61253), .Q(to_acu1
		[54]));
	notech_mux2 i_40811(.S(n_57609), .A(to_acu1[54]), .B(n_39548), .Z(n_34374
		));
	notech_reg to_acu1_reg_55(.CP(n_61816), .D(n_34380), .CD(n_61253), .Q(to_acu1
		[55]));
	notech_mux2 i_40819(.S(n_57609), .A(to_acu1[55]), .B(n_39550), .Z(n_34380
		));
	notech_reg to_acu1_reg_56(.CP(n_61816), .D(n_34386), .CD(n_61253), .Q(to_acu1
		[56]));
	notech_mux2 i_40827(.S(n_57609), .A(to_acu1[56]), .B(n_39552), .Z(n_34386
		));
	notech_ao4 i_472(.A(n_2107), .B(n_2106), .C(valid_len[3]), .D(n_9538), .Z
		(n_2111));
	notech_reg to_acu1_reg_57(.CP(n_61816), .D(n_34392), .CD(n_61255), .Q(to_acu1
		[57]));
	notech_mux2 i_40835(.S(n_57609), .A(to_acu1[57]), .B(n_39554), .Z(n_34392
		));
	notech_and2 i_469(.A(n_9538), .B(valid_len[3]), .Z(n_2110));
	notech_reg to_acu1_reg_58(.CP(n_61819), .D(n_34398), .CD(n_61255), .Q(to_acu1
		[58]));
	notech_mux2 i_40843(.S(n_57609), .A(to_acu1[58]), .B(n_39556), .Z(n_34398
		));
	notech_reg to_acu1_reg_59(.CP(n_61819), .D(n_34404), .CD(n_61255), .Q(to_acu1
		[59]));
	notech_mux2 i_40851(.S(n_57610), .A(to_acu1[59]), .B(n_39558), .Z(n_34404
		));
	notech_reg to_acu1_reg_60(.CP(n_61819), .D(n_34410), .CD(n_61255), .Q(to_acu1
		[60]));
	notech_mux2 i_40859(.S(n_57593), .A(to_acu1[60]), .B(n_39560), .Z(n_34410
		));
	notech_ao4 i_468(.A(valid_len[2]), .B(n_38328), .C(n_2104), .D(n_2103), 
		.Z(n_2107));
	notech_reg to_acu1_reg_61(.CP(n_61816), .D(n_34416), .CD(n_61255), .Q(to_acu1
		[61]));
	notech_mux2 i_40867(.S(n_57593), .A(to_acu1[61]), .B(n_39562), .Z(n_34416
		));
	notech_and2 i_467(.A(valid_len[2]), .B(n_38328), .Z(n_2106));
	notech_reg to_acu1_reg_62(.CP(n_61816), .D(n_34422), .CD(n_61258), .Q(to_acu1
		[62]));
	notech_mux2 i_40875(.S(n_57593), .A(to_acu1[62]), .B(n_39564), .Z(n_34422
		));
	notech_or2 i_395(.A(valid_len[1]), .B(n_39850), .Z(n_2105));
	notech_reg to_acu1_reg_63(.CP(n_61816), .D(n_34428), .CD(n_61258), .Q(to_acu1
		[63]));
	notech_mux2 i_40883(.S(n_57593), .A(to_acu1[63]), .B(n_39566), .Z(n_34428
		));
	notech_ao3 i_464(.A(valid_len[0]), .B(n_2105), .C(n_1741), .Z(n_2104));
	notech_reg to_acu1_reg_64(.CP(n_61816), .D(n_34434), .CD(n_61255), .Q(to_acu1
		[64]));
	notech_mux2 i_40891(.S(n_57593), .A(to_acu1[64]), .B(n_38904), .Z(n_34434
		));
	notech_and2 i_462(.A(valid_len[1]), .B(n_39850), .Z(n_2103));
	notech_reg to_acu1_reg_65(.CP(n_61816), .D(n_34440), .CD(n_61255), .Q(to_acu1
		[65]));
	notech_mux2 i_40899(.S(n_57593), .A(to_acu1[65]), .B(n_38906), .Z(n_34440
		));
	notech_reg to_acu1_reg_66(.CP(n_61816), .D(n_34446), .CD(n_61255), .Q(to_acu1
		[66]));
	notech_mux2 i_40907(.S(n_57593), .A(to_acu1[66]), .B(n_38908), .Z(n_34446
		));
	notech_reg to_acu1_reg_67(.CP(n_61816), .D(n_34452), .CD(n_61255), .Q(to_acu1
		[67]));
	notech_mux2 i_40915(.S(n_57620), .A(to_acu1[67]), .B(n_38910), .Z(n_34452
		));
	notech_reg to_acu1_reg_68(.CP(n_61816), .D(n_34458), .CD(n_61255), .Q(to_acu1
		[68]));
	notech_mux2 i_40923(.S(n_57620), .A(to_acu1[68]), .B(n_39573), .Z(n_34458
		));
	notech_reg to_acu1_reg_69(.CP(n_61816), .D(n_34464), .CD(n_61255), .Q(to_acu1
		[69]));
	notech_mux2 i_40931(.S(n_57620), .A(to_acu1[69]), .B(n_38912), .Z(n_34464
		));
	notech_reg to_acu1_reg_70(.CP(n_61816), .D(n_34470), .CD(n_61255), .Q(to_acu1
		[70]));
	notech_mux2 i_40939(.S(n_57593), .A(to_acu1[70]), .B(n_39500), .Z(n_34470
		));
	notech_and2 i_370(.A(n_39860), .B(n_38653), .Z(n_2097));
	notech_reg to_acu1_reg_71(.CP(n_61816), .D(n_34476), .CD(n_61253), .Q(to_acu1
		[71]));
	notech_mux2 i_40947(.S(n_57593), .A(to_acu1[71]), .B(n_39505), .Z(n_34476
		));
	notech_reg to_acu1_reg_72(.CP(n_61816), .D(n_34482), .CD(n_61255), .Q(to_acu1
		[72]));
	notech_mux2 i_40955(.S(n_57620), .A(to_acu1[72]), .B(n_39510), .Z(n_34482
		));
	notech_reg to_acu1_reg_73(.CP(n_61816), .D(n_34488), .CD(n_61255), .Q(to_acu1
		[73]));
	notech_mux2 i_40963(.S(n_57610), .A(to_acu1[73]), .B(n_39513), .Z(n_34488
		));
	notech_and2 i_369(.A(imm_sz[1]), .B(i_ptr[1]), .Z(n_2094));
	notech_reg to_acu1_reg_74(.CP(n_61810), .D(n_34494), .CD(n_61255), .Q(to_acu1
		[74]));
	notech_mux2 i_40971(.S(n_57610), .A(to_acu1[74]), .B(n_39516), .Z(n_34494
		));
	notech_reg to_acu1_reg_75(.CP(n_61808), .D(n_34500), .CD(n_61255), .Q(to_acu1
		[75]));
	notech_mux2 i_40979(.S(n_57610), .A(to_acu1[75]), .B(n_39521), .Z(n_34500
		));
	notech_reg to_acu1_reg_76(.CP(n_61808), .D(n_34506), .CD(n_61255), .Q(to_acu1
		[76]));
	notech_mux2 i_40987(.S(n_57610), .A(to_acu1[76]), .B(n_39526), .Z(n_34506
		));
	notech_and4 i_75034(.A(n_59686), .B(n_2141), .C(n_18050174), .D(n_2089),
		 .Z(n_2091));
	notech_reg to_acu1_reg_77(.CP(n_61808), .D(n_34512), .CD(n_61255), .Q(to_acu1
		[77]));
	notech_mux2 i_40995(.S(n_57610), .A(to_acu1[77]), .B(n_39531), .Z(n_34512
		));
	notech_and4 i_34(.A(n_2081), .B(n_2080), .C(n_2088), .D(n_2085), .Z(n_2090
		));
	notech_reg to_acu1_reg_78(.CP(n_61808), .D(n_34518), .CD(n_61247), .Q(to_acu1
		[78]));
	notech_mux2 i_41003(.S(n_57610), .A(to_acu1[78]), .B(n_39536), .Z(n_34518
		));
	notech_or2 i_442(.A(n_2798), .B(n_2090), .Z(n_2089));
	notech_reg to_acu1_reg_79(.CP(n_61808), .D(n_34524), .CD(n_61247), .Q(to_acu1
		[79]));
	notech_mux2 i_41011(.S(n_57610), .A(to_acu1[79]), .B(n_39541), .Z(n_34524
		));
	notech_nand2 i_438(.A(twobyte), .B(n_2087), .Z(n_2088));
	notech_reg to_acu1_reg_80(.CP(n_61808), .D(n_34530), .CD(n_61247), .Q(to_acu1
		[80]));
	notech_mux2 i_41019(.S(n_57593), .A(to_acu1[80]), .B(n_38914), .Z(n_34530
		));
	notech_nand2 i_35(.A(n_40164), .B(n_40179), .Z(n_2087));
	notech_reg to_acu1_reg_81(.CP(n_61808), .D(n_34536), .CD(n_61247), .Q(to_acu1
		[81]));
	notech_mux2 i_41027(.S(n_57593), .A(to_acu1[81]), .B(n_38916), .Z(n_34536
		));
	notech_nao3 i_36(.A(n_1810), .B(n_2821), .C(n_1972), .Z(n_2086));
	notech_reg to_acu1_reg_82(.CP(n_61808), .D(n_34542), .CD(n_61247), .Q(to_acu1
		[82]));
	notech_mux2 i_41035(.S(n_57593), .A(to_acu1[82]), .B(n_39588), .Z(n_34542
		));
	notech_nao3 i_437(.A(n_40210), .B(n_2086), .C(n_2812), .Z(n_2085));
	notech_reg to_acu1_reg_83(.CP(n_61808), .D(n_34548), .CD(n_61247), .Q(to_acu1
		[83]));
	notech_mux2 i_41043(.S(n_57610), .A(to_acu1[83]), .B(n_39590), .Z(n_34548
		));
	notech_nand2 i_430(.A(n_1973), .B(n_40211), .Z(n_2084));
	notech_reg to_acu1_reg_84(.CP(n_61808), .D(n_34554), .CD(n_61247), .Q(to_acu1
		[84]));
	notech_mux2 i_41051(.S(n_57610), .A(to_acu1[84]), .B(n_38918), .Z(n_34554
		));
	notech_nand2 i_418(.A(\to_acu2_0[5] ), .B(\to_acu2_0[59] ), .Z(n_2083)
		);
	notech_reg to_acu1_reg_85(.CP(n_61808), .D(n_34560), .CD(n_61247), .Q(to_acu1
		[85]));
	notech_mux2 i_41059(.S(n_57610), .A(to_acu1[85]), .B(n_38920), .Z(n_34560
		));
	notech_nand2 i_354(.A(n_40181), .B(n_40145), .Z(n_2082));
	notech_reg to_acu1_reg_86(.CP(n_61805), .D(n_34566), .CD(n_61247), .Q(to_acu1
		[86]));
	notech_mux2 i_41067(.S(n_57598), .A(to_acu1[86]), .B(n_38922), .Z(n_34566
		));
	notech_nand3 i_416(.A(n_40164), .B(twobyte), .C(n_2082), .Z(n_2081));
	notech_reg to_acu1_reg_87(.CP(n_61805), .D(n_34572), .CD(n_61247), .Q(to_acu1
		[87]));
	notech_mux2 i_41075(.S(n_57598), .A(to_acu1[87]), .B(n_39597), .Z(n_34572
		));
	notech_nand2 i_415(.A(n_2812), .B(n_40210), .Z(n_2080));
	notech_reg to_acu1_reg_88(.CP(n_61805), .D(n_34578), .CD(n_61247), .Q(to_acu1
		[88]));
	notech_mux2 i_41083(.S(n_57598), .A(to_acu1[88]), .B(n_39599), .Z(n_34578
		));
	notech_nand2 i_396(.A(\to_acu2_0[48] ), .B(\to_acu2_0[5] ), .Z(n_2079)
		);
	notech_reg to_acu1_reg_89(.CP(n_61805), .D(n_34584), .CD(n_61244), .Q(to_acu1
		[89]));
	notech_mux2 i_41091(.S(n_57598), .A(to_acu1[89]), .B(n_39602), .Z(n_34584
		));
	notech_nand3 i_388(.A(\to_acu2_0[23] ), .B(\to_acu2_0[21] ), .C(\to_acu2_0[22] 
		), .Z(n_2078));
	notech_reg to_acu1_reg_90(.CP(n_61805), .D(n_34590), .CD(n_61244), .Q(to_acu1
		[90]));
	notech_mux2 i_41099(.S(n_57598), .A(to_acu1[90]), .B(n_38924), .Z(n_34590
		));
	notech_nand2 i_385(.A(n_2209), .B(\to_acu2_0[13] ), .Z(n_2077));
	notech_reg to_acu1_reg_91(.CP(n_61805), .D(n_34596), .CD(n_61244), .Q(to_acu1
		[91]));
	notech_mux2 i_41107(.S(n_57598), .A(to_acu1[91]), .B(n_38926), .Z(n_34596
		));
	notech_or4 i_372(.A(\to_acu2_0[9] ), .B(\to_acu2_0[10] ), .C(\to_acu2_0[11] 
		), .D(\to_acu2_0[8] ), .Z(n_2076));
	notech_reg to_acu1_reg_92(.CP(n_61805), .D(n_34602), .CD(n_61244), .Q(to_acu1
		[92]));
	notech_mux2 i_41115(.S(n_57598), .A(to_acu1[92]), .B(n_38928), .Z(n_34602
		));
	notech_reg to_acu1_reg_93(.CP(n_61805), .D(n_34608), .CD(n_61244), .Q(to_acu1
		[93]));
	notech_mux2 i_41123(.S(n_57598), .A(to_acu1[93]), .B(n_38930), .Z(n_34608
		));
	notech_and4 i_1130055(.A(n_40173), .B(n_57713), .C(n_40172), .D(n_2856),
		 .Z(n_2074));
	notech_reg to_acu1_reg_94(.CP(n_61805), .D(n_34614), .CD(n_61244), .Q(to_acu1
		[94]));
	notech_mux2 i_41131(.S(n_57598), .A(to_acu1[94]), .B(n_38932), .Z(n_34614
		));
	notech_nao3 i_138(.A(n_5717), .B(n_2220), .C(n_251191358), .Z(n_2073));
	notech_reg to_acu1_reg_95(.CP(n_61805), .D(n_34620), .CD(n_61244), .Q(to_acu1
		[95]));
	notech_mux2 i_41139(.S(n_57599), .A(to_acu1[95]), .B(n_38934), .Z(n_34620
		));
	notech_or4 i_71544(.A(db67), .B(\to_acu2_0[3] ), .C(\to_acu2_0[4] ), .D(n_2074
		), .Z(n_2072));
	notech_reg to_acu1_reg_96(.CP(n_61810), .D(n_34626), .CD(n_61244), .Q(to_acu1
		[96]));
	notech_mux2 i_41147(.S(n_57598), .A(to_acu1[96]), .B(n_38936), .Z(n_34626
		));
	notech_nand2 i_6325(.A(idx_deco[1]), .B(idx_deco[0]), .Z(n_2071));
	notech_reg to_acu1_reg_97(.CP(n_61810), .D(n_34632), .CD(n_61244), .Q(to_acu1
		[97]));
	notech_mux2 i_41155(.S(n_57598), .A(to_acu1[97]), .B(n_38938), .Z(n_34632
		));
	notech_ao3 i_42073378(.A(in128[1]), .B(in128[2]), .C(n_58712), .Z(n_49757
		));
	notech_reg to_acu1_reg_98(.CP(n_61810), .D(n_34638), .CD(n_61244), .Q(to_acu1
		[98]));
	notech_mux2 i_41163(.S(n_57598), .A(to_acu1[98]), .B(n_38940), .Z(n_34638
		));
	notech_reg to_acu1_reg_99(.CP(n_61810), .D(n_34644), .CD(n_61249), .Q(to_acu1
		[99]));
	notech_mux2 i_41171(.S(n_57593), .A(to_acu1[99]), .B(n_38942), .Z(n_34644
		));
	notech_reg to_acu1_reg_100(.CP(n_61810), .D(n_34650), .CD(n_61249), .Q(to_acu1
		[100]));
	notech_mux2 i_41179(.S(n_57593), .A(to_acu1[100]), .B(n_38944), .Z(n_34650
		));
	notech_reg to_acu1_reg_101(.CP(n_61810), .D(n_34656), .CD(n_61249), .Q(to_acu1
		[101]));
	notech_mux2 i_41187(.S(n_57598), .A(to_acu1[101]), .B(n_39621), .Z(n_34656
		));
	notech_and3 i_94472439(.A(n_251091357), .B(n_250991356), .C(n_849150), .Z
		(n_2067));
	notech_reg to_acu1_reg_102(.CP(n_61810), .D(n_34662), .CD(n_61249), .Q(to_acu1
		[102]));
	notech_mux2 i_41195(.S(n_57593), .A(to_acu1[102]), .B(n_39623), .Z(n_34662
		));
	notech_reg to_acu1_reg_103(.CP(n_61810), .D(n_34668), .CD(n_61249), .Q(to_acu1
		[103]));
	notech_mux2 i_41203(.S(n_57593), .A(to_acu1[103]), .B(n_39626), .Z(n_34668
		));
	notech_reg to_acu1_reg_104(.CP(n_61810), .D(n_34674), .CD(n_61249), .Q(to_acu1
		[104]));
	notech_mux2 i_41211(.S(n_57593), .A(to_acu1[104]), .B(n_39628), .Z(n_34674
		));
	notech_reg to_acu1_reg_105(.CP(n_61810), .D(n_34680), .CD(n_61249), .Q(to_acu1
		[105]));
	notech_mux2 i_41219(.S(n_57598), .A(to_acu1[105]), .B(n_39630), .Z(n_34680
		));
	notech_reg to_acu1_reg_106(.CP(n_61810), .D(n_34686), .CD(n_61249), .Q(to_acu1
		[106]));
	notech_mux2 i_41227(.S(n_57598), .A(to_acu1[106]), .B(n_38946), .Z(n_34686
		));
	notech_ao4 i_1173365(.A(n_5304), .B(n_2073), .C(n_3813), .D(n_2062), .Z(n_849150
		));
	notech_reg to_acu1_reg_107(.CP(n_61808), .D(n_34692), .CD(n_61249), .Q(to_acu1
		[107]));
	notech_mux2 i_41235(.S(n_57598), .A(to_acu1[107]), .B(n_39634), .Z(n_34692
		));
	notech_nand3 i_95072433(.A(db67), .B(fpu), .C(n_41571), .Z(n_2062));
	notech_reg to_acu1_reg_108(.CP(n_61808), .D(n_34698), .CD(n_61249), .Q(to_acu1
		[108]));
	notech_mux2 i_41243(.S(n_57598), .A(to_acu1[108]), .B(n_39637), .Z(n_34698
		));
	notech_or4 i_16473212(.A(n_56589), .B(db67), .C(pc_req), .D(\to_acu2_0[4] 
		), .Z(n_1249153));
	notech_reg to_acu1_reg_109(.CP(n_61808), .D(n_34704), .CD(n_61249), .Q(to_acu1
		[109]));
	notech_mux2 i_41251(.S(n_57598), .A(to_acu1[109]), .B(n_39639), .Z(n_34704
		));
	notech_reg to_acu1_reg_110(.CP(n_61808), .D(n_34710), .CD(n_61247), .Q(to_acu1
		[110]));
	notech_mux2 i_41259(.S(n_57598), .A(to_acu1[110]), .B(n_39641), .Z(n_34710
		));
	notech_ao4 i_97072418(.A(n_2928), .B(n_40060), .C(n_2929), .D(n_40044), 
		.Z(n_2060));
	notech_reg to_acu1_reg_111(.CP(n_61808), .D(n_34716), .CD(n_61247), .Q(to_acu1
		[111]));
	notech_mux2 i_41267(.S(n_57598), .A(to_acu1[111]), .B(n_39644), .Z(n_34716
		));
	notech_reg to_acu1_reg_112(.CP(n_61810), .D(n_34722), .CD(n_61247), .Q(to_acu1
		[112]));
	notech_mux2 i_41275(.S(n_57599), .A(to_acu1[112]), .B(n_38948), .Z(n_34722
		));
	notech_ao4 i_97272416(.A(n_2922), .B(n_40036), .C(n_2923), .D(n_40052), 
		.Z(n_1993));
	notech_reg to_acu1_reg_113(.CP(n_61810), .D(n_34728), .CD(n_61247), .Q(to_acu1
		[113]));
	notech_mux2 i_41283(.S(n_57604), .A(to_acu1[113]), .B(n_39648), .Z(n_34728
		));
	notech_ao4 i_97372415(.A(n_2921), .B(n_40028), .C(n_3060), .D(n_40020), 
		.Z(n_1992));
	notech_reg to_acu1_reg_114(.CP(n_61810), .D(n_34734), .CD(n_61247), .Q(to_acu1
		[114]));
	notech_mux2 i_41291(.S(n_57604), .A(to_acu1[114]), .B(n_39650), .Z(n_34734
		));
	notech_nao3 i_97572413(.A(n_38431), .B(n_38428), .C(n_3120), .Z(n_1991)
		);
	notech_reg to_acu1_reg_115(.CP(n_61808), .D(n_34740), .CD(n_61249), .Q(to_acu1
		[115]));
	notech_mux2 i_41299(.S(n_57604), .A(to_acu1[115]), .B(n_39652), .Z(n_34740
		));
	notech_reg to_acu1_reg_116(.CP(n_61808), .D(n_34746), .CD(n_61249), .Q(to_acu1
		[116]));
	notech_mux2 i_41307(.S(n_57599), .A(to_acu1[116]), .B(n_39655), .Z(n_34746
		));
	notech_reg to_acu1_reg_117(.CP(n_61826), .D(n_34752), .CD(n_61249), .Q(to_acu1
		[117]));
	notech_mux2 i_41315(.S(n_57599), .A(to_acu1[117]), .B(n_39657), .Z(n_34752
		));
	notech_reg to_acu1_reg_118(.CP(n_61826), .D(n_34758), .CD(n_61247), .Q(to_acu1
		[118]));
	notech_mux2 i_41323(.S(n_57604), .A(to_acu1[118]), .B(n_39659), .Z(n_34758
		));
	notech_reg to_acu1_reg_119(.CP(n_61826), .D(n_34764), .CD(n_61247), .Q(to_acu1
		[119]));
	notech_mux2 i_41331(.S(n_57604), .A(to_acu1[119]), .B(n_39662), .Z(n_34764
		));
	notech_nao3 i_873368(.A(n_2175), .B(in128[37]), .C(n_53815), .Z(n_1985)
		);
	notech_reg to_acu1_reg_120(.CP(n_61826), .D(n_34770), .CD(n_61258), .Q(to_acu1
		[120]));
	notech_mux2 i_41339(.S(n_57604), .A(to_acu1[120]), .B(n_39664), .Z(n_34770
		));
	notech_reg to_acu1_reg_121(.CP(n_61826), .D(n_34776), .CD(n_61265), .Q(to_acu1
		[121]));
	notech_mux2 i_41347(.S(n_57604), .A(to_acu1[121]), .B(n_39666), .Z(n_34776
		));
	notech_reg to_acu1_reg_122(.CP(n_61826), .D(n_34782), .CD(n_61265), .Q(to_acu1
		[122]));
	notech_mux2 i_41355(.S(n_57604), .A(to_acu1[122]), .B(n_39668), .Z(n_34782
		));
	notech_or4 i_66172722(.A(n_5674), .B(n_251191358), .C(n_5726), .D(n_5717
		), .Z(n_1982));
	notech_reg to_acu1_reg_123(.CP(n_61826), .D(n_34788), .CD(n_61265), .Q(to_acu1
		[123]));
	notech_mux2 i_41363(.S(n_57604), .A(to_acu1[123]), .B(n_38950), .Z(n_34788
		));
	notech_nand2 i_66072723(.A(fpu), .B(n_39826), .Z(n_1980));
	notech_reg to_acu1_reg_124(.CP(n_61826), .D(n_34794), .CD(n_61265), .Q(to_acu1
		[124]));
	notech_mux2 i_41371(.S(n_57604), .A(to_acu1[124]), .B(n_38952), .Z(n_34794
		));
	notech_or4 i_65972724(.A(n_1249153), .B(n_251191358), .C(n_5674), .D(n_38516
		), .Z(n_1979));
	notech_reg to_acu1_reg_125(.CP(n_61826), .D(n_34800), .CD(n_61265), .Q(to_acu1
		[125]));
	notech_mux2 i_41379(.S(n_57604), .A(to_acu1[125]), .B(n_38954), .Z(n_34800
		));
	notech_reg to_acu1_reg_126(.CP(n_61826), .D(n_34806), .CD(n_61265), .Q(to_acu1
		[126]));
	notech_mux2 i_41387(.S(n_57599), .A(to_acu1[126]), .B(n_38956), .Z(n_34806
		));
	notech_and4 i_72272661(.A(n_2060), .B(n_1993), .C(n_1992), .D(n_1985), .Z
		(n_1977));
	notech_reg to_acu1_reg_127(.CP(n_61826), .D(n_34812), .CD(n_61265), .Q(to_acu1
		[127]));
	notech_mux2 i_41395(.S(n_57599), .A(to_acu1[127]), .B(n_38958), .Z(n_34812
		));
	notech_reg to_acu1_reg_128(.CP(n_61824), .D(n_34818), .CD(n_61265), .Q(to_acu1
		[128]));
	notech_mux2 i_41403(.S(n_57599), .A(to_acu1[128]), .B(n_39675), .Z(n_34818
		));
	notech_reg to_acu1_reg_129(.CP(n_61824), .D(n_34824), .CD(n_61265), .Q(to_acu1
		[129]));
	notech_mux2 i_41411(.S(n_57599), .A(to_acu1[129]), .B(n_39677), .Z(n_34824
		));
	notech_reg to_acu1_reg_130(.CP(n_61824), .D(n_34830), .CD(n_61265), .Q(to_acu1
		[130]));
	notech_mux2 i_41419(.S(n_57599), .A(to_acu1[130]), .B(n_39679), .Z(n_34830
		));
	notech_reg to_acu1_reg_131(.CP(n_61824), .D(n_34836), .CD(n_61265), .Q(to_acu1
		[131]));
	notech_mux2 i_41427(.S(n_57599), .A(to_acu1[131]), .B(n_39681), .Z(n_34836
		));
	notech_reg to_acu1_reg_132(.CP(n_61824), .D(n_34842), .CD(n_61263), .Q(to_acu1
		[132]));
	notech_mux2 i_41435(.S(n_57599), .A(to_acu1[132]), .B(n_39683), .Z(n_34842
		));
	notech_reg to_acu1_reg_133(.CP(n_61826), .D(n_34848), .CD(n_61263), .Q(to_acu1
		[133]));
	notech_mux2 i_41443(.S(n_57599), .A(to_acu1[133]), .B(n_39685), .Z(n_34848
		));
	notech_reg to_acu1_reg_134(.CP(n_61826), .D(n_34854), .CD(n_61263), .Q(to_acu1
		[134]));
	notech_mux2 i_41451(.S(n_57599), .A(to_acu1[134]), .B(n_39687), .Z(n_34854
		));
	notech_reg to_acu1_reg_135(.CP(n_61824), .D(n_34860), .CD(n_61263), .Q(to_acu1
		[135]));
	notech_mux2 i_41459(.S(n_57599), .A(to_acu1[135]), .B(n_39689), .Z(n_34860
		));
	notech_reg to_acu1_reg_136(.CP(n_61824), .D(n_34866), .CD(n_61263), .Q(to_acu1
		[136]));
	notech_mux2 i_41467(.S(n_57599), .A(to_acu1[136]), .B(n_39691), .Z(n_34866
		));
	notech_reg to_acu1_reg_137(.CP(n_61824), .D(n_34872), .CD(n_61263), .Q(to_acu1
		[137]));
	notech_mux2 i_41475(.S(n_57599), .A(to_acu1[137]), .B(n_39693), .Z(n_34872
		));
	notech_reg to_acu1_reg_138(.CP(n_61830), .D(n_34878), .CD(n_61265), .Q(to_acu1
		[138]));
	notech_mux2 i_41483(.S(n_57599), .A(to_acu1[138]), .B(n_38960), .Z(n_34878
		));
	notech_reg to_acu1_reg_139(.CP(n_61830), .D(n_34884), .CD(n_61263), .Q(to_acu1
		[139]));
	notech_mux2 i_41491(.S(n_57620), .A(to_acu1[139]), .B(n_39696), .Z(n_34884
		));
	notech_reg to_acu1_reg_140(.CP(n_61830), .D(n_34890), .CD(n_61263), .Q(to_acu1
		[140]));
	notech_mux2 i_41499(.S(n_57633), .A(to_acu1[140]), .B(n_39698), .Z(n_34890
		));
	notech_reg to_acu1_reg_141(.CP(n_61830), .D(n_34896), .CD(n_61263), .Q(to_acu1
		[141]));
	notech_mux2 i_41507(.S(n_57633), .A(to_acu1[141]), .B(n_39700), .Z(n_34896
		));
	notech_reg to_acu1_reg_142(.CP(n_61830), .D(n_34902), .CD(n_61269), .Q(to_acu1
		[142]));
	notech_mux2 i_41515(.S(n_57633), .A(to_acu1[142]), .B(n_39702), .Z(n_34902
		));
	notech_reg to_acu1_reg_143(.CP(n_61830), .D(n_34908), .CD(n_61269), .Q(to_acu1
		[143]));
	notech_mux2 i_41523(.S(n_57633), .A(to_acu1[143]), .B(n_39704), .Z(n_34908
		));
	notech_reg to_acu1_reg_144(.CP(n_61830), .D(n_34914), .CD(n_61269), .Q(to_acu1
		[144]));
	notech_mux2 i_41531(.S(n_57633), .A(to_acu1[144]), .B(n_39706), .Z(n_34914
		));
	notech_reg to_acu1_reg_145(.CP(n_61830), .D(n_34920), .CD(n_61269), .Q(to_acu1
		[145]));
	notech_mux2 i_41539(.S(n_57633), .A(to_acu1[145]), .B(n_39708), .Z(n_34920
		));
	notech_reg to_acu1_reg_146(.CP(n_61830), .D(n_34926), .CD(n_61269), .Q(to_acu1
		[146]));
	notech_mux2 i_41547(.S(n_57633), .A(to_acu1[146]), .B(n_38962), .Z(n_34926
		));
	notech_reg to_acu1_reg_147(.CP(n_61830), .D(n_34932), .CD(n_61269), .Q(to_acu1
		[147]));
	notech_mux2 i_41555(.S(n_57633), .A(to_acu1[147]), .B(n_39711), .Z(n_34932
		));
	notech_reg to_acu1_reg_148(.CP(n_61830), .D(n_34938), .CD(n_61269), .Q(to_acu1
		[148]));
	notech_mux2 i_41563(.S(n_57633), .A(to_acu1[148]), .B(n_39713), .Z(n_34938
		));
	notech_reg to_acu1_reg_149(.CP(n_61826), .D(n_34944), .CD(n_61269), .Q(to_acu1
		[149]));
	notech_mux2 i_41571(.S(n_57633), .A(to_acu1[149]), .B(n_39715), .Z(n_34944
		));
	notech_reg to_acu1_reg_150(.CP(n_61826), .D(n_34950), .CD(n_61269), .Q(to_acu1
		[150]));
	notech_mux2 i_41579(.S(n_57633), .A(to_acu1[150]), .B(n_39717), .Z(n_34950
		));
	notech_reg to_acu1_reg_151(.CP(n_61826), .D(n_34956), .CD(n_61269), .Q(to_acu1
		[151]));
	notech_mux2 i_41587(.S(n_57633), .A(to_acu1[151]), .B(n_39719), .Z(n_34956
		));
	notech_reg to_acu1_reg_152(.CP(n_61826), .D(n_34962), .CD(n_61269), .Q(to_acu1
		[152]));
	notech_mux2 i_41595(.S(n_57633), .A(to_acu1[152]), .B(n_39721), .Z(n_34962
		));
	notech_reg to_acu1_reg_153(.CP(n_61826), .D(n_34968), .CD(n_61265), .Q(to_acu1
		[153]));
	notech_mux2 i_41603(.S(n_57632), .A(to_acu1[153]), .B(n_39723), .Z(n_34968
		));
	notech_reg to_acu1_reg_154(.CP(n_61830), .D(n_34974), .CD(n_61265), .Q(to_acu1
		[154]));
	notech_mux2 i_41611(.S(n_57632), .A(to_acu1[154]), .B(n_39725), .Z(n_34974
		));
	notech_reg to_acu1_reg_155(.CP(n_61830), .D(n_34980), .CD(n_61265), .Q(to_acu1
		[155]));
	notech_mux2 i_41619(.S(n_57632), .A(to_acu1[155]), .B(n_39727), .Z(n_34980
		));
	notech_reg to_acu1_reg_156(.CP(n_61830), .D(n_34986), .CD(n_61265), .Q(to_acu1
		[156]));
	notech_mux2 i_41627(.S(n_57632), .A(to_acu1[156]), .B(n_39729), .Z(n_34986
		));
	notech_reg to_acu1_reg_157(.CP(n_61830), .D(n_34992), .CD(n_61265), .Q(to_acu1
		[157]));
	notech_mux2 i_41635(.S(n_57632), .A(to_acu1[157]), .B(n_39731), .Z(n_34992
		));
	notech_reg to_acu1_reg_158(.CP(n_61830), .D(n_34998), .CD(n_61269), .Q(to_acu1
		[158]));
	notech_mux2 i_41643(.S(n_57632), .A(to_acu1[158]), .B(n_39733), .Z(n_34998
		));
	notech_reg to_acu1_reg_159(.CP(n_61824), .D(n_35004), .CD(n_61269), .Q(to_acu1
		[159]));
	notech_mux2 i_41651(.S(n_57632), .A(to_acu1[159]), .B(n_39735), .Z(n_35004
		));
	notech_reg to_acu1_reg_160(.CP(n_61819), .D(n_35010), .CD(n_61269), .Q(to_acu1
		[160]));
	notech_mux2 i_41659(.S(n_57633), .A(to_acu1[160]), .B(n_39737), .Z(n_35010
		));
	notech_reg to_acu1_reg_161(.CP(n_61821), .D(n_35016), .CD(n_61265), .Q(to_acu1
		[161]));
	notech_mux2 i_41667(.S(n_57633), .A(to_acu1[161]), .B(n_39739), .Z(n_35016
		));
	notech_reg to_acu1_reg_162(.CP(n_61819), .D(n_35022), .CD(n_61269), .Q(to_acu1
		[162]));
	notech_mux2 i_41675(.S(n_57633), .A(to_acu1[162]), .B(n_39741), .Z(n_35022
		));
	notech_reg to_acu1_reg_163(.CP(n_61819), .D(n_35028), .CD(n_61258), .Q(to_acu1
		[163]));
	notech_mux2 i_41683(.S(n_57632), .A(to_acu1[163]), .B(n_38964), .Z(n_35028
		));
	notech_reg to_acu1_reg_164(.CP(n_61819), .D(n_35034), .CD(n_61260), .Q(to_acu1
		[164]));
	notech_mux2 i_41691(.S(n_57633), .A(to_acu1[164]), .B(n_38966), .Z(n_35034
		));
	notech_reg to_acu1_reg_165(.CP(n_61821), .D(n_35040), .CD(n_61258), .Q(to_acu1
		[165]));
	notech_mux2 i_41699(.S(n_57633), .A(to_acu1[165]), .B(n_38968), .Z(n_35040
		));
	notech_reg to_acu1_reg_166(.CP(n_61821), .D(n_35046), .CD(n_61258), .Q(to_acu1
		[166]));
	notech_mux2 i_41707(.S(n_57638), .A(to_acu1[166]), .B(n_38970), .Z(n_35046
		));
	notech_reg to_acu1_reg_167(.CP(n_61821), .D(n_35052), .CD(n_61258), .Q(to_acu1
		[167]));
	notech_mux2 i_41715(.S(n_57643), .A(to_acu1[167]), .B(n_38972), .Z(n_35052
		));
	notech_reg to_acu1_reg_168(.CP(n_61821), .D(n_35058), .CD(n_61260), .Q(to_acu1
		[168]));
	notech_mux2 i_41723(.S(n_57643), .A(to_acu1[168]), .B(n_38974), .Z(n_35058
		));
	notech_reg to_acu1_reg_169(.CP(n_61821), .D(n_35064), .CD(n_61260), .Q(to_acu1
		[169]));
	notech_mux2 i_41731(.S(n_57643), .A(to_acu1[169]), .B(n_38398), .Z(n_35064
		));
	notech_reg to_acu1_reg_170(.CP(n_61819), .D(n_35070), .CD(n_61260), .Q(to_acu1
		[170]));
	notech_mux2 i_41739(.S(n_57643), .A(to_acu1[170]), .B(n_39750), .Z(n_35070
		));
	notech_reg to_acu1_reg_171(.CP(n_61819), .D(n_35076), .CD(n_61260), .Q(to_acu1
		[171]));
	notech_mux2 i_41747(.S(n_57643), .A(to_acu1[171]), .B(n_39752), .Z(n_35076
		));
	notech_reg to_acu1_reg_172(.CP(n_61819), .D(n_35082), .CD(n_61260), .Q(to_acu1
		[172]));
	notech_mux2 i_41755(.S(n_57643), .A(to_acu1[172]), .B(n_38976), .Z(n_35082
		));
	notech_reg to_acu1_reg_173(.CP(n_61819), .D(n_35088), .CD(n_61258), .Q(to_acu1
		[173]));
	notech_mux2 i_41763(.S(n_57643), .A(to_acu1[173]), .B(n_38978), .Z(n_35088
		));
	notech_reg to_acu1_reg_174(.CP(n_61819), .D(n_35094), .CD(n_61258), .Q(to_acu1
		[174]));
	notech_mux2 i_41771(.S(n_57643), .A(to_acu1[174]), .B(n_39756), .Z(n_35094
		));
	notech_reg to_acu1_reg_175(.CP(n_61819), .D(n_35100), .CD(n_61258), .Q(to_acu1
		[175]));
	notech_mux2 i_41779(.S(n_57643), .A(to_acu1[175]), .B(n_38980), .Z(n_35100
		));
	notech_reg to_acu1_reg_176(.CP(n_61819), .D(n_35106), .CD(n_61258), .Q(to_acu1
		[176]));
	notech_mux2 i_41787(.S(n_57643), .A(to_acu1[176]), .B(n_39759), .Z(n_35106
		));
	notech_reg to_acu1_reg_177(.CP(n_61819), .D(n_35112), .CD(n_61258), .Q(to_acu1
		[177]));
	notech_mux2 i_41795(.S(n_57643), .A(to_acu1[177]), .B(n_39761), .Z(n_35112
		));
	notech_reg to_acu1_reg_178(.CP(n_61819), .D(n_35118), .CD(n_61258), .Q(to_acu1
		[178]));
	notech_mux2 i_41803(.S(n_57643), .A(to_acu1[178]), .B(n_38982), .Z(n_35118
		));
	notech_reg to_acu1_reg_179(.CP(n_61819), .D(n_35124), .CD(n_61258), .Q(to_acu1
		[179]));
	notech_mux2 i_41811(.S(n_57643), .A(to_acu1[179]), .B(n_39764), .Z(n_35124
		));
	notech_reg to_acu1_reg_180(.CP(n_61819), .D(n_35130), .CD(n_61258), .Q(to_acu1
		[180]));
	notech_mux2 i_41819(.S(n_57638), .A(to_acu1[180]), .B(n_39766), .Z(n_35130
		));
	notech_reg to_acu1_reg_181(.CP(n_61824), .D(n_35136), .CD(n_61258), .Q(to_acu1
		[181]));
	notech_mux2 i_41827(.S(n_57638), .A(to_acu1[181]), .B(n_39768), .Z(n_35136
		));
	notech_reg to_acu1_reg_182(.CP(n_61824), .D(n_35142), .CD(n_61258), .Q(to_acu1
		[182]));
	notech_mux2 i_41835(.S(n_57638), .A(to_acu1[182]), .B(n_39770), .Z(n_35142
		));
	notech_reg to_acu1_reg_183(.CP(n_61824), .D(n_35148), .CD(n_61258), .Q(to_acu1
		[183]));
	notech_mux2 i_41843(.S(n_57638), .A(to_acu1[183]), .B(n_39772), .Z(n_35148
		));
	notech_reg to_acu1_reg_184(.CP(n_61821), .D(n_35154), .CD(n_61263), .Q(to_acu1
		[184]));
	notech_mux2 i_41851(.S(n_57638), .A(to_acu1[184]), .B(n_39774), .Z(n_35154
		));
	notech_reg to_acu1_reg_185(.CP(n_61824), .D(n_35160), .CD(n_61263), .Q(to_acu1
		[185]));
	notech_mux2 i_41859(.S(n_57638), .A(to_acu1[185]), .B(n_39776), .Z(n_35160
		));
	notech_reg to_acu1_reg_186(.CP(n_61824), .D(n_35166), .CD(n_61263), .Q(to_acu1
		[186]));
	notech_mux2 i_41867(.S(n_57638), .A(to_acu1[186]), .B(n_39778), .Z(n_35166
		));
	notech_reg to_acu1_reg_187(.CP(n_61824), .D(n_35172), .CD(n_61260), .Q(to_acu1
		[187]));
	notech_mux2 i_41875(.S(n_57638), .A(to_acu1[187]), .B(n_39780), .Z(n_35172
		));
	notech_reg to_acu1_reg_188(.CP(n_61824), .D(n_35178), .CD(n_61263), .Q(to_acu1
		[188]));
	notech_mux2 i_41883(.S(n_57643), .A(to_acu1[188]), .B(n_39782), .Z(n_35178
		));
	notech_reg to_acu1_reg_189(.CP(n_61824), .D(n_35184), .CD(n_61263), .Q(to_acu1
		[189]));
	notech_mux2 i_41891(.S(n_57643), .A(to_acu1[189]), .B(n_39784), .Z(n_35184
		));
	notech_reg to_acu1_reg_190(.CP(n_61824), .D(n_35190), .CD(n_61263), .Q(to_acu1
		[190]));
	notech_mux2 i_41899(.S(n_57638), .A(to_acu1[190]), .B(n_39786), .Z(n_35190
		));
	notech_reg to_acu1_reg_191(.CP(n_61821), .D(n_35196), .CD(n_61263), .Q(to_acu1
		[191]));
	notech_mux2 i_41907(.S(n_57638), .A(to_acu1[191]), .B(n_39788), .Z(n_35196
		));
	notech_reg to_acu1_reg_192(.CP(n_61821), .D(n_35202), .CD(n_61263), .Q(to_acu1
		[192]));
	notech_mux2 i_41915(.S(n_57638), .A(to_acu1[192]), .B(n_39790), .Z(n_35202
		));
	notech_reg to_acu1_reg_193(.CP(n_61821), .D(n_35208), .CD(n_61263), .Q(to_acu1
		[193]));
	notech_mux2 i_41923(.S(n_57621), .A(to_acu1[193]), .B(n_39792), .Z(n_35208
		));
	notech_reg to_acu1_reg_194(.CP(n_61821), .D(n_35214), .CD(n_61260), .Q(to_acu1
		[194]));
	notech_mux2 i_41931(.S(n_57621), .A(to_acu1[194]), .B(n_39794), .Z(n_35214
		));
	notech_reg to_acu1_reg_195(.CP(n_61821), .D(n_35220), .CD(n_61260), .Q(to_acu1
		[195]));
	notech_mux2 i_41939(.S(n_57621), .A(to_acu1[195]), .B(n_39796), .Z(n_35220
		));
	notech_reg to_acu1_reg_196(.CP(n_61821), .D(n_35226), .CD(n_61260), .Q(to_acu1
		[196]));
	notech_mux2 i_41947(.S(n_57621), .A(to_acu1[196]), .B(n_39798), .Z(n_35226
		));
	notech_reg to_acu1_reg_197(.CP(n_61821), .D(n_35232), .CD(n_61260), .Q(to_acu1
		[197]));
	notech_mux2 i_41955(.S(n_57621), .A(to_acu1[197]), .B(n_38984), .Z(n_35232
		));
	notech_reg to_acu1_reg_198(.CP(n_61821), .D(n_35238), .CD(n_61260), .Q(to_acu1
		[198]));
	notech_mux2 i_41963(.S(n_57621), .A(to_acu1[198]), .B(n_38986), .Z(n_35238
		));
	notech_reg to_acu1_reg_199(.CP(n_61821), .D(n_35244), .CD(n_61260), .Q(to_acu1
		[199]));
	notech_mux2 i_41971(.S(n_57621), .A(to_acu1[199]), .B(n_38988), .Z(n_35244
		));
	notech_reg to_acu1_reg_200(.CP(n_61821), .D(n_35250), .CD(n_61260), .Q(to_acu1
		[200]));
	notech_mux2 i_41979(.S(n_57621), .A(to_acu1[200]), .B(n_38990), .Z(n_35250
		));
	notech_reg to_acu1_reg_201(.CP(n_61821), .D(n_35256), .CD(n_61260), .Q(to_acu1
		[201]));
	notech_mux2 i_41987(.S(n_57621), .A(to_acu1[201]), .B(n_39804), .Z(n_35256
		));
	notech_reg to_acu1_reg_202(.CP(n_61789), .D(n_35262), .CD(n_61260), .Q(to_acu1
		[202]));
	notech_mux2 i_41995(.S(n_57621), .A(to_acu1[202]), .B(n_38992), .Z(n_35262
		));
	notech_reg to_acu1_reg_203(.CP(n_61789), .D(n_35268), .CD(n_61260), .Q(to_acu1
		[203]));
	notech_mux2 i_42003(.S(n_57621), .A(to_acu1[203]), .B(n_38994), .Z(n_35268
		));
	notech_reg to_acu1_reg_204(.CP(n_61789), .D(n_35274), .CD(n_61260), .Q(to_acu1
		[204]));
	notech_mux2 i_42011(.S(n_57621), .A(to_acu1[204]), .B(n_39808), .Z(n_35274
		));
	notech_reg to_acu1_reg_205(.CP(n_61789), .D(n_35280), .CD(n_61244), .Q(to_acu1
		[205]));
	notech_mux2 i_42019(.S(n_57621), .A(to_acu1[205]), .B(n_39810), .Z(n_35280
		));
	notech_reg to_acu1_reg_206(.CP(n_61789), .D(n_35286), .CD(n_61228), .Q(to_acu1
		[206]));
	notech_mux2 i_42027(.S(n_57620), .A(to_acu1[206]), .B(n_39812), .Z(n_35286
		));
	notech_reg to_acu1_reg_207(.CP(n_61789), .D(n_35292), .CD(n_61228), .Q(to_acu1
		[207]));
	notech_mux2 i_42035(.S(n_57620), .A(to_acu1[207]), .B(n_38996), .Z(n_35292
		));
	notech_reg to_acu1_reg_208(.CP(n_61789), .D(n_35298), .CD(n_61228), .Q(to_acu1
		[208]));
	notech_mux2 i_42043(.S(n_57620), .A(to_acu1[208]), .B(n_39815), .Z(n_35298
		));
	notech_reg to_acu1_reg_209(.CP(n_61789), .D(n_35304), .CD(n_61226), .Q(to_acu1
		[209]));
	notech_mux2 i_42051(.S(n_57620), .A(to_acu1[209]), .B(n_39817), .Z(n_35304
		));
	notech_reg to_acu1_reg_210(.CP(n_61789), .D(n_35310), .CD(n_61228), .Q(to_acu1
		[210]));
	notech_mux2 i_42059(.S(n_57620), .A(to_acu1[210]), .B(n_39819), .Z(n_35310
		));
	notech_reg iack_reg(.CP(n_61789), .D(n_38408), .CD(n_61228), .Q(iack));
	notech_reg imm0_reg_0(.CP(n_61787), .D(n_35318), .CD(n_61228), .Q(\imm0[0] 
		));
	notech_mux2 i_42071(.S(n_55013), .A(\imm0[0] ), .B(n_39368), .Z(n_35318)
		);
	notech_reg imm0_reg_1(.CP(n_61787), .D(n_35324), .CD(n_61228), .Q(\imm0[1] 
		));
	notech_mux2 i_42079(.S(n_55013), .A(\imm0[1] ), .B(n_38872), .Z(n_35324)
		);
	notech_reg imm0_reg_2(.CP(n_61787), .D(n_35330), .CD(n_61228), .Q(\imm0[2] 
		));
	notech_mux2 i_42087(.S(n_54983), .A(\imm0[2] ), .B(n_38874), .Z(n_35330)
		);
	notech_reg imm0_reg_3(.CP(n_61787), .D(n_35336), .CD(n_61228), .Q(\imm0[3] 
		));
	notech_mux2 i_42095(.S(n_54983), .A(\imm0[3] ), .B(n_39371), .Z(n_35336)
		);
	notech_reg imm0_reg_4(.CP(n_61787), .D(n_35342), .CD(n_61226), .Q(\imm0[4] 
		));
	notech_mux2 i_42103(.S(n_55013), .A(\imm0[4] ), .B(n_38876), .Z(n_35342)
		);
	notech_reg imm0_reg_5(.CP(n_61787), .D(n_35348), .CD(n_61226), .Q(\imm0[5] 
		));
	notech_mux2 i_42111(.S(n_55013), .A(\imm0[5] ), .B(n_39374), .Z(n_35348)
		);
	notech_reg imm0_reg_6(.CP(n_61787), .D(n_35354), .CD(n_61226), .Q(\imm0[6] 
		));
	notech_mux2 i_42119(.S(n_55013), .A(\imm0[6] ), .B(n_39377), .Z(n_35354)
		);
	notech_reg imm0_reg_7(.CP(n_61787), .D(n_35360), .CD(n_61226), .Q(\imm0[7] 
		));
	notech_mux2 i_42127(.S(n_55013), .A(\imm0[7] ), .B(n_39380), .Z(n_35360)
		);
	notech_reg imm0_reg_8(.CP(n_61787), .D(n_35366), .CD(n_61226), .Q(\imm0[8] 
		));
	notech_mux2 i_42135(.S(n_54983), .A(\imm0[8] ), .B(n_39383), .Z(n_35366)
		);
	notech_reg imm0_reg_9(.CP(n_61787), .D(n_35372), .CD(n_61226), .Q(\imm0[9] 
		));
	notech_mux2 i_42143(.S(n_54983), .A(\imm0[9] ), .B(n_39386), .Z(n_35372)
		);
	notech_reg imm0_reg_10(.CP(n_61787), .D(n_35378), .CD(n_61226), .Q(\imm0[10] 
		));
	notech_mux2 i_42151(.S(n_54983), .A(\imm0[10] ), .B(n_39389), .Z(n_35378
		));
	notech_reg imm0_reg_11(.CP(n_61792), .D(n_35384), .CD(n_61226), .Q(\imm0[11] 
		));
	notech_mux2 i_42159(.S(n_54983), .A(\imm0[11] ), .B(n_39392), .Z(n_35384
		));
	notech_reg imm0_reg_12(.CP(n_61792), .D(n_35390), .CD(n_61226), .Q(\imm0[12] 
		));
	notech_mux2 i_42167(.S(n_54983), .A(\imm0[12] ), .B(n_39395), .Z(n_35390
		));
	notech_reg imm0_reg_13(.CP(n_61792), .D(n_35396), .CD(n_61226), .Q(\imm0[13] 
		));
	notech_mux2 i_42175(.S(n_54983), .A(\imm0[13] ), .B(n_39398), .Z(n_35396
		));
	notech_reg imm0_reg_14(.CP(n_61792), .D(n_35402), .CD(n_61226), .Q(\imm0[14] 
		));
	notech_mux2 i_42183(.S(n_54983), .A(\imm0[14] ), .B(n_39401), .Z(n_35402
		));
	notech_reg imm0_reg_15(.CP(n_61792), .D(n_35408), .CD(n_61231), .Q(\imm0[15] 
		));
	notech_mux2 i_42191(.S(n_54983), .A(\imm0[15] ), .B(n_39404), .Z(n_35408
		));
	notech_reg imm0_reg_16(.CP(n_61792), .D(n_35414), .CD(n_61231), .Q(\imm0[16] 
		));
	notech_mux2 i_42199(.S(n_55013), .A(\imm0[16] ), .B(n_39407), .Z(n_35414
		));
	notech_reg imm0_reg_17(.CP(n_61792), .D(n_35420), .CD(n_61231), .Q(\imm0[17] 
		));
	notech_mux2 i_42207(.S(n_55017), .A(\imm0[17] ), .B(n_39410), .Z(n_35420
		));
	notech_reg imm0_reg_18(.CP(n_61792), .D(n_35426), .CD(n_61231), .Q(\imm0[18] 
		));
	notech_mux2 i_42215(.S(n_55017), .A(\imm0[18] ), .B(n_39413), .Z(n_35426
		));
	notech_reg imm0_reg_19(.CP(n_61792), .D(n_35432), .CD(n_61231), .Q(\imm0[19] 
		));
	notech_mux2 i_42223(.S(n_55017), .A(\imm0[19] ), .B(n_38396), .Z(n_35432
		));
	notech_reg imm0_reg_20(.CP(n_61792), .D(n_35438), .CD(n_61231), .Q(\imm0[20] 
		));
	notech_mux2 i_42231(.S(n_55017), .A(\imm0[20] ), .B(n_39416), .Z(n_35438
		));
	notech_reg imm0_reg_21(.CP(n_61792), .D(n_35444), .CD(n_61231), .Q(\imm0[21] 
		));
	notech_mux2 i_42239(.S(n_55017), .A(\imm0[21] ), .B(n_39419), .Z(n_35444
		));
	notech_reg imm0_reg_22(.CP(n_61789), .D(n_35450), .CD(n_61231), .Q(\imm0[22] 
		));
	notech_mux2 i_42247(.S(n_55017), .A(\imm0[22] ), .B(n_39422), .Z(n_35450
		));
	notech_reg imm0_reg_23(.CP(n_61789), .D(n_35456), .CD(n_61231), .Q(\imm0[23] 
		));
	notech_mux2 i_42255(.S(n_55017), .A(\imm0[23] ), .B(n_39424), .Z(n_35456
		));
	notech_reg imm0_reg_24(.CP(n_61789), .D(n_35462), .CD(n_61231), .Q(\imm0[24] 
		));
	notech_mux2 i_42263(.S(n_55017), .A(\imm0[24] ), .B(n_39427), .Z(n_35462
		));
	notech_reg imm0_reg_25(.CP(n_61789), .D(n_35468), .CD(n_61231), .Q(\imm0[25] 
		));
	notech_mux2 i_42271(.S(n_55013), .A(\imm0[25] ), .B(n_39431), .Z(n_35468
		));
	notech_reg imm0_reg_26(.CP(n_61789), .D(n_35474), .CD(n_61228), .Q(\imm0[26] 
		));
	notech_mux2 i_42279(.S(n_55013), .A(\imm0[26] ), .B(n_39821), .Z(n_35474
		));
	notech_reg imm0_reg_27(.CP(n_61792), .D(n_35480), .CD(n_61228), .Q(\imm0[27] 
		));
	notech_mux2 i_42287(.S(n_55013), .A(\imm0[27] ), .B(n_39433), .Z(n_35480
		));
	notech_reg imm0_reg_28(.CP(n_61792), .D(n_35486), .CD(n_61228), .Q(\imm0[28] 
		));
	notech_mux2 i_42295(.S(n_55013), .A(\imm0[28] ), .B(n_39438), .Z(n_35486
		));
	notech_reg imm0_reg_29(.CP(n_61789), .D(n_35492), .CD(n_61228), .Q(\imm0[29] 
		));
	notech_mux2 i_42303(.S(n_55013), .A(\imm0[29] ), .B(n_38397), .Z(n_35492
		));
	notech_reg imm0_reg_30(.CP(n_61789), .D(n_35498), .CD(n_61228), .Q(\imm0[30] 
		));
	notech_mux2 i_42311(.S(n_55013), .A(\imm0[30] ), .B(n_39441), .Z(n_35498
		));
	notech_reg imm0_reg_31(.CP(n_61789), .D(n_35504), .CD(n_61228), .Q(\imm0[31] 
		));
	notech_mux2 i_42319(.S(n_55013), .A(\imm0[31] ), .B(n_39445), .Z(n_35504
		));
	notech_reg imm0_reg_32(.CP(n_61787), .D(n_35510), .CD(n_61231), .Q(\imm0[32] 
		));
	notech_mux2 i_42327(.S(n_55013), .A(\imm0[32] ), .B(n_39450), .Z(n_35510
		));
	notech_reg imm0_reg_33(.CP(n_61782), .D(n_35516), .CD(n_61228), .Q(\imm0[33] 
		));
	notech_mux2 i_42335(.S(n_54998), .A(\imm0[33] ), .B(n_39452), .Z(n_35516
		));
	notech_reg imm0_reg_34(.CP(n_61782), .D(n_35522), .CD(n_61228), .Q(\imm0[34] 
		));
	notech_mux2 i_42343(.S(n_54998), .A(\imm0[34] ), .B(n_39454), .Z(n_35522
		));
	notech_reg imm0_reg_35(.CP(n_61782), .D(n_35528), .CD(n_61228), .Q(\imm0[35] 
		));
	notech_mux2 i_42351(.S(n_54998), .A(\imm0[35] ), .B(n_39456), .Z(n_35528
		));
	notech_reg imm0_reg_36(.CP(n_61782), .D(n_35534), .CD(n_61221), .Q(\imm0[36] 
		));
	notech_mux2 i_42359(.S(n_54998), .A(\imm0[36] ), .B(n_39461), .Z(n_35534
		));
	notech_reg imm0_reg_37(.CP(n_61782), .D(n_35540), .CD(n_61221), .Q(\imm0[37] 
		));
	notech_mux2 i_42367(.S(n_55003), .A(\imm0[37] ), .B(n_39466), .Z(n_35540
		));
	notech_reg imm0_reg_38(.CP(n_61784), .D(n_35546), .CD(n_61221), .Q(\imm0[38] 
		));
	notech_mux2 i_42375(.S(n_55003), .A(\imm0[38] ), .B(n_39471), .Z(n_35546
		));
	notech_reg imm0_reg_39(.CP(n_61784), .D(n_35552), .CD(n_61221), .Q(\imm0[39] 
		));
	notech_mux2 i_42383(.S(n_54998), .A(\imm0[39] ), .B(n_39474), .Z(n_35552
		));
	notech_reg imm0_reg_40(.CP(n_61784), .D(n_35558), .CD(n_61221), .Q(\imm0[40] 
		));
	notech_mux2 i_42391(.S(n_55003), .A(\imm0[40] ), .B(n_39476), .Z(n_35558
		));
	notech_reg imm0_reg_41(.CP(n_61782), .D(n_35564), .CD(n_61223), .Q(\imm0[41] 
		));
	notech_mux2 i_42399(.S(n_54998), .A(\imm0[41] ), .B(n_39478), .Z(n_35564
		));
	notech_reg imm0_reg_42(.CP(n_61782), .D(n_35570), .CD(n_61223), .Q(\imm0[42] 
		));
	notech_mux2 i_42407(.S(n_54998), .A(\imm0[42] ), .B(n_39480), .Z(n_35570
		));
	notech_reg imm0_reg_43(.CP(n_61782), .D(n_35576), .CD(n_61223), .Q(\imm0[43] 
		));
	notech_mux2 i_42415(.S(n_54998), .A(\imm0[43] ), .B(n_39482), .Z(n_35576
		));
	notech_reg imm0_reg_44(.CP(n_61782), .D(n_35582), .CD(n_61221), .Q(\imm0[44] 
		));
	notech_mux2 i_42423(.S(n_54998), .A(\imm0[44] ), .B(n_39484), .Z(n_35582
		));
	notech_reg imm0_reg_45(.CP(n_61782), .D(n_35588), .CD(n_61221), .Q(\imm0[45] 
		));
	notech_mux2 i_42431(.S(n_54998), .A(\imm0[45] ), .B(n_39486), .Z(n_35588
		));
	notech_reg imm0_reg_46(.CP(n_61782), .D(n_35594), .CD(n_61221), .Q(\imm0[46] 
		));
	notech_mux2 i_42439(.S(n_54998), .A(\imm0[46] ), .B(n_39490), .Z(n_35594
		));
	notech_reg imm0_reg_47(.CP(n_61782), .D(n_35600), .CD(n_61221), .Q(\imm0[47] 
		));
	notech_mux2 i_42447(.S(n_54998), .A(\imm0[47] ), .B(n_39495), .Z(n_35600
		));
	notech_reg opz2_reg_0(.CP(n_61782), .D(n_35606), .CD(n_61221), .Q(opz2[0
		]));
	notech_mux2 i_42455(.S(n_54198), .A(opz2[0]), .B(n_3201), .Z(n_35606));
	notech_reg opz2_reg_1(.CP(n_61782), .D(n_35612), .CD(n_61221), .Q(opz2[1
		]));
	notech_mux2 i_42463(.S(n_54198), .A(opz2[1]), .B(n_3199), .Z(n_35612));
	notech_reg_set opz2_reg_2(.CP(n_61782), .D(n_35618), .SD(n_61221), .Q(opz2
		[2]));
	notech_mux2 i_42471(.S(n_54198), .A(opz2[2]), .B(n_265491501), .Z(n_35618
		));
	notech_reg opz1_reg_0(.CP(n_61782), .D(n_35624), .CD(n_61221), .Q(opz1[0
		]));
	notech_mux2 i_42479(.S(n_57620), .A(opz1[0]), .B(n_39362), .Z(n_35624)
		);
	notech_reg opz1_reg_1(.CP(n_61782), .D(n_35630), .CD(n_61221), .Q(opz1[1
		]));
	notech_mux2 i_42487(.S(n_57620), .A(opz1[1]), .B(n_39365), .Z(n_35630)
		);
	notech_reg_set opz1_reg_2(.CP(n_61782), .D(n_35636), .SD(n_61221), .Q(opz1
		[2]));
	notech_mux2 i_42495(.S(n_57620), .A(opz1[2]), .B(n_265691503), .Z(n_35636
		));
	notech_reg_set inst_deco_reg_0(.CP(n_61784), .D(n_35642), .SD(n_61221), 
		.Q(inst_deco[0]));
	notech_mux2 i_42503(.S(n_58446), .A(n_45249), .B(inst_deco[0]), .Z(n_35642
		));
	notech_reg_set inst_deco_reg_1(.CP(n_61787), .D(n_35648), .SD(n_61221), 
		.Q(inst_deco[1]));
	notech_mux2 i_42511(.S(n_58446), .A(n_45255), .B(inst_deco[1]), .Z(n_35648
		));
	notech_reg_set inst_deco_reg_2(.CP(n_61784), .D(n_35654), .SD(n_61221), 
		.Q(inst_deco[2]));
	notech_mux2 i_42519(.S(n_58446), .A(n_45261), .B(inst_deco[2]), .Z(n_35654
		));
	notech_reg_set inst_deco_reg_3(.CP(n_61784), .D(n_35660), .SD(n_61223), 
		.Q(inst_deco[3]));
	notech_mux2 i_42527(.S(n_58446), .A(n_45267), .B(inst_deco[3]), .Z(n_35660
		));
	notech_reg_set inst_deco_reg_4(.CP(n_61784), .D(n_35666), .SD(n_61226), 
		.Q(inst_deco[4]));
	notech_mux2 i_42535(.S(n_58446), .A(n_45273), .B(inst_deco[4]), .Z(n_35666
		));
	notech_reg_set inst_deco_reg_5(.CP(n_61787), .D(n_35672), .SD(n_61223), 
		.Q(inst_deco[5]));
	notech_mux2 i_42543(.S(n_58446), .A(n_3235), .B(inst_deco[5]), .Z(n_35672
		));
	notech_reg_set inst_deco_reg_6(.CP(n_61787), .D(n_35678), .SD(n_61223), 
		.Q(inst_deco[6]));
	notech_mux2 i_42551(.S(n_58446), .A(n_45285), .B(inst_deco[6]), .Z(n_35678
		));
	notech_reg_set inst_deco_reg_7(.CP(n_61787), .D(n_35684), .SD(n_61223), 
		.Q(inst_deco[7]));
	notech_mux2 i_42559(.S(n_58446), .A(n_45291), .B(inst_deco[7]), .Z(n_35684
		));
	notech_reg_set inst_deco_reg_8(.CP(n_61787), .D(n_35690), .SD(n_61226), 
		.Q(inst_deco[8]));
	notech_mux2 i_42567(.S(n_58446), .A(n_3234), .B(inst_deco[8]), .Z(n_35690
		));
	notech_reg_set inst_deco_reg_9(.CP(n_61787), .D(n_35696), .SD(n_61226), 
		.Q(inst_deco[9]));
	notech_mux2 i_42575(.S(n_58446), .A(n_45303), .B(inst_deco[9]), .Z(n_35696
		));
	notech_reg_set inst_deco_reg_10(.CP(n_61784), .D(n_35702), .SD(n_61226),
		 .Q(inst_deco[10]));
	notech_mux2 i_42583(.S(n_58446), .A(n_3233), .B(inst_deco[10]), .Z(n_35702
		));
	notech_reg_set inst_deco_reg_11(.CP(n_61784), .D(n_35708), .SD(n_61226),
		 .Q(inst_deco[11]));
	notech_mux2 i_42591(.S(n_58446), .A(n_3232), .B(inst_deco[11]), .Z(n_35708
		));
	notech_reg_set inst_deco_reg_12(.CP(n_61784), .D(n_35714), .SD(n_61226),
		 .Q(inst_deco[12]));
	notech_mux2 i_42599(.S(n_58446), .A(n_3231), .B(inst_deco[12]), .Z(n_35714
		));
	notech_reg_set inst_deco_reg_13(.CP(n_61784), .D(n_35720), .SD(n_61223),
		 .Q(inst_deco[13]));
	notech_mux2 i_42607(.S(n_58446), .A(n_265991506), .B(inst_deco[13]), .Z(n_35720
		));
	notech_reg_set inst_deco_reg_14(.CP(n_61784), .D(n_35726), .SD(n_61223),
		 .Q(inst_deco[14]));
	notech_mux2 i_42615(.S(n_58446), .A(n_3230), .B(inst_deco[14]), .Z(n_35726
		));
	notech_reg_set inst_deco_reg_15(.CP(n_61784), .D(n_35732), .SD(n_61223),
		 .Q(inst_deco[15]));
	notech_mux2 i_42623(.S(n_58446), .A(n_3229), .B(inst_deco[15]), .Z(n_35732
		));
	notech_reg_set inst_deco_reg_16(.CP(n_61784), .D(n_35738), .SD(n_61223),
		 .Q(inst_deco[16]));
	notech_mux2 i_42631(.S(n_58444), .A(n_3228), .B(inst_deco[16]), .Z(n_35738
		));
	notech_reg_set inst_deco_reg_17(.CP(n_61784), .D(n_35744), .SD(n_61223),
		 .Q(inst_deco[17]));
	notech_mux2 i_42639(.S(n_58444), .A(n_3227), .B(inst_deco[17]), .Z(n_35744
		));
	notech_reg_set inst_deco_reg_18(.CP(n_61784), .D(n_35750), .SD(n_61223),
		 .Q(inst_deco[18]));
	notech_mux2 i_42647(.S(n_58444), .A(n_3226), .B(inst_deco[18]), .Z(n_35750
		));
	notech_reg_set inst_deco_reg_19(.CP(n_61784), .D(n_35756), .SD(n_61223),
		 .Q(inst_deco[19]));
	notech_mux2 i_42655(.S(n_58444), .A(n_3225), .B(inst_deco[19]), .Z(n_35756
		));
	notech_reg_set inst_deco_reg_20(.CP(n_61784), .D(n_35762), .SD(n_61223),
		 .Q(inst_deco[20]));
	notech_mux2 i_42663(.S(n_58444), .A(n_3224), .B(inst_deco[20]), .Z(n_35762
		));
	notech_reg_set inst_deco_reg_21(.CP(n_61800), .D(n_35768), .SD(n_61223),
		 .Q(inst_deco[21]));
	notech_mux2 i_42671(.S(n_58444), .A(n_3223), .B(inst_deco[21]), .Z(n_35768
		));
	notech_reg_set inst_deco_reg_22(.CP(n_61800), .D(n_35774), .SD(n_61223),
		 .Q(inst_deco[22]));
	notech_mux2 i_42679(.S(n_58444), .A(n_3222), .B(inst_deco[22]), .Z(n_35774
		));
	notech_reg_set inst_deco_reg_23(.CP(n_61800), .D(n_35780), .SD(n_61223),
		 .Q(inst_deco[23]));
	notech_mux2 i_42687(.S(n_58444), .A(n_3221), .B(inst_deco[23]), .Z(n_35780
		));
	notech_reg_set inst_deco_reg_24(.CP(n_61800), .D(n_35786), .SD(n_61231),
		 .Q(inst_deco[24]));
	notech_mux2 i_42695(.S(n_58444), .A(n_3220), .B(inst_deco[24]), .Z(n_35786
		));
	notech_reg_set inst_deco_reg_25(.CP(n_61800), .D(n_35792), .SD(n_61239),
		 .Q(inst_deco[25]));
	notech_mux2 i_42703(.S(n_58444), .A(n_45399), .B(inst_deco[25]), .Z(n_35792
		));
	notech_reg_set inst_deco_reg_26(.CP(n_61803), .D(n_35798), .SD(n_61239),
		 .Q(inst_deco[26]));
	notech_mux2 i_42711(.S(n_58444), .A(n_45405), .B(inst_deco[26]), .Z(n_35798
		));
	notech_reg_set inst_deco_reg_27(.CP(n_61803), .D(n_35804), .SD(n_61239),
		 .Q(inst_deco[27]));
	notech_mux2 i_42719(.S(n_58444), .A(n_45411), .B(inst_deco[27]), .Z(n_35804
		));
	notech_reg_set inst_deco_reg_28(.CP(n_61803), .D(n_35810), .SD(n_61239),
		 .Q(inst_deco[28]));
	notech_mux2 i_42727(.S(n_58444), .A(n_45417), .B(inst_deco[28]), .Z(n_35810
		));
	notech_reg_set inst_deco_reg_29(.CP(n_61803), .D(n_35816), .SD(n_61239),
		 .Q(inst_deco[29]));
	notech_mux2 i_42735(.S(n_58444), .A(n_45423), .B(inst_deco[29]), .Z(n_35816
		));
	notech_reg_set inst_deco_reg_30(.CP(n_61803), .D(n_35822), .SD(n_61242),
		 .Q(inst_deco[30]));
	notech_mux2 i_42743(.S(n_58444), .A(n_45429), .B(inst_deco[30]), .Z(n_35822
		));
	notech_reg_set inst_deco_reg_31(.CP(n_61800), .D(n_35828), .SD(n_61242),
		 .Q(inst_deco[31]));
	notech_mux2 i_42751(.S(n_58444), .A(n_45435), .B(inst_deco[31]), .Z(n_35828
		));
	notech_reg_set inst_deco_reg_32(.CP(n_61800), .D(n_35834), .SD(n_61242),
		 .Q(inst_deco[32]));
	notech_mux2 i_42759(.S(n_58451), .A(n_45441), .B(inst_deco[32]), .Z(n_35834
		));
	notech_reg_set inst_deco_reg_33(.CP(n_61800), .D(n_35840), .SD(n_61239),
		 .Q(inst_deco[33]));
	notech_mux2 i_42767(.S(n_58451), .A(n_45447), .B(inst_deco[33]), .Z(n_35840
		));
	notech_reg_set inst_deco_reg_34(.CP(n_61800), .D(n_35846), .SD(n_61242),
		 .Q(inst_deco[34]));
	notech_mux2 i_42775(.S(n_58451), .A(n_45453), .B(inst_deco[34]), .Z(n_35846
		));
	notech_reg_set inst_deco_reg_35(.CP(n_61800), .D(n_35852), .SD(n_61239),
		 .Q(inst_deco[35]));
	notech_mux2 i_42783(.S(n_58451), .A(n_45459), .B(inst_deco[35]), .Z(n_35852
		));
	notech_reg_set inst_deco_reg_36(.CP(n_61800), .D(n_35858), .SD(n_61239),
		 .Q(inst_deco[36]));
	notech_mux2 i_42791(.S(n_58451), .A(n_45465), .B(inst_deco[36]), .Z(n_35858
		));
	notech_reg_set inst_deco_reg_37(.CP(n_61800), .D(n_35864), .SD(n_61239),
		 .Q(inst_deco[37]));
	notech_mux2 i_42799(.S(n_58451), .A(n_45471), .B(inst_deco[37]), .Z(n_35864
		));
	notech_reg_set inst_deco_reg_38(.CP(n_61800), .D(n_35870), .SD(n_61239),
		 .Q(inst_deco[38]));
	notech_mux2 i_42807(.S(n_58451), .A(n_45477), .B(inst_deco[38]), .Z(n_35870
		));
	notech_reg_set inst_deco_reg_39(.CP(n_61800), .D(n_35876), .SD(n_61239),
		 .Q(inst_deco[39]));
	notech_mux2 i_42815(.S(n_58451), .A(n_45483), .B(inst_deco[39]), .Z(n_35876
		));
	notech_reg_set inst_deco_reg_40(.CP(n_61800), .D(n_35882), .SD(n_61239),
		 .Q(inst_deco[40]));
	notech_mux2 i_42823(.S(n_58451), .A(n_45489), .B(inst_deco[40]), .Z(n_35882
		));
	notech_reg_set inst_deco_reg_41(.CP(n_61800), .D(n_35888), .SD(n_61239),
		 .Q(inst_deco[41]));
	notech_mux2 i_42831(.S(n_58451), .A(n_45495), .B(inst_deco[41]), .Z(n_35888
		));
	notech_reg_set inst_deco_reg_42(.CP(n_61805), .D(n_35894), .SD(n_61239),
		 .Q(inst_deco[42]));
	notech_mux2 i_42839(.S(n_58451), .A(n_45501), .B(inst_deco[42]), .Z(n_35894
		));
	notech_reg_set inst_deco_reg_43(.CP(n_61805), .D(n_35900), .SD(n_61239),
		 .Q(inst_deco[43]));
	notech_mux2 i_42847(.S(n_58451), .A(n_45507), .B(inst_deco[43]), .Z(n_35900
		));
	notech_reg_set inst_deco_reg_44(.CP(n_61805), .D(n_35906), .SD(n_61239),
		 .Q(inst_deco[44]));
	notech_mux2 i_42855(.S(n_58451), .A(n_45513), .B(inst_deco[44]), .Z(n_35906
		));
	notech_reg_set inst_deco_reg_45(.CP(n_61803), .D(n_35912), .SD(n_61239),
		 .Q(inst_deco[45]));
	notech_mux2 i_42863(.S(n_58451), .A(n_45519), .B(inst_deco[45]), .Z(n_35912
		));
	notech_reg_set inst_deco_reg_46(.CP(n_61803), .D(n_35918), .SD(n_61244),
		 .Q(inst_deco[46]));
	notech_mux2 i_42871(.S(n_58451), .A(n_45525), .B(inst_deco[46]), .Z(n_35918
		));
	notech_reg_set inst_deco_reg_47(.CP(n_61805), .D(n_35924), .SD(n_61244),
		 .Q(inst_deco[47]));
	notech_mux2 i_42879(.S(n_58451), .A(n_45531), .B(inst_deco[47]), .Z(n_35924
		));
	notech_reg_set inst_deco_reg_48(.CP(n_61805), .D(n_35930), .SD(n_61242),
		 .Q(inst_deco[48]));
	notech_mux2 i_42887(.S(n_58449), .A(n_45537), .B(inst_deco[48]), .Z(n_35930
		));
	notech_reg_set inst_deco_reg_49(.CP(n_61805), .D(n_35936), .SD(n_61242),
		 .Q(inst_deco[49]));
	notech_mux2 i_42895(.S(n_58449), .A(n_45543), .B(inst_deco[49]), .Z(n_35936
		));
	notech_reg_set inst_deco_reg_50(.CP(n_61805), .D(n_35942), .SD(n_61242),
		 .Q(inst_deco[50]));
	notech_mux2 i_42903(.S(n_58449), .A(n_45549), .B(inst_deco[50]), .Z(n_35942
		));
	notech_reg_set inst_deco_reg_51(.CP(n_61805), .D(n_35948), .SD(n_61244),
		 .Q(inst_deco[51]));
	notech_mux2 i_42911(.S(n_58449), .A(n_45555), .B(inst_deco[51]), .Z(n_35948
		));
	notech_reg_set inst_deco_reg_52(.CP(n_61803), .D(n_35954), .SD(n_61244),
		 .Q(inst_deco[52]));
	notech_mux2 i_42919(.S(n_58449), .A(n_45561), .B(inst_deco[52]), .Z(n_35954
		));
	notech_reg_set inst_deco_reg_53(.CP(n_61803), .D(n_35960), .SD(n_61244),
		 .Q(inst_deco[53]));
	notech_mux2 i_42927(.S(n_58449), .A(n_45567), .B(inst_deco[53]), .Z(n_35960
		));
	notech_reg_set inst_deco_reg_54(.CP(n_61803), .D(n_35966), .SD(n_61244),
		 .Q(inst_deco[54]));
	notech_mux2 i_42935(.S(n_58449), .A(n_3219), .B(inst_deco[54]), .Z(n_35966
		));
	notech_reg_set inst_deco_reg_55(.CP(n_61803), .D(n_35972), .SD(n_61244),
		 .Q(inst_deco[55]));
	notech_mux2 i_42943(.S(n_58449), .A(n_45579), .B(inst_deco[55]), .Z(n_35972
		));
	notech_reg_set inst_deco_reg_56(.CP(n_61803), .D(n_35978), .SD(n_61242),
		 .Q(inst_deco[56]));
	notech_mux2 i_42951(.S(n_58449), .A(n_45585), .B(inst_deco[56]), .Z(n_35978
		));
	notech_reg_set inst_deco_reg_57(.CP(n_61803), .D(n_35984), .SD(n_61242),
		 .Q(inst_deco[57]));
	notech_mux2 i_42959(.S(n_58449), .A(n_3218), .B(inst_deco[57]), .Z(n_35984
		));
	notech_reg_set inst_deco_reg_58(.CP(n_61803), .D(n_35990), .SD(n_61242),
		 .Q(inst_deco[58]));
	notech_mux2 i_42967(.S(n_58449), .A(n_45597), .B(inst_deco[58]), .Z(n_35990
		));
	notech_reg_set inst_deco_reg_59(.CP(n_61803), .D(n_35996), .SD(n_61242),
		 .Q(inst_deco[59]));
	notech_mux2 i_42975(.S(n_58449), .A(n_45603), .B(inst_deco[59]), .Z(n_35996
		));
	notech_reg_set inst_deco_reg_60(.CP(n_61803), .D(n_36002), .SD(n_61242),
		 .Q(inst_deco[60]));
	notech_mux2 i_42983(.S(n_58449), .A(n_45609), .B(inst_deco[60]), .Z(n_36002
		));
	notech_reg_set inst_deco_reg_61(.CP(n_61803), .D(n_36008), .SD(n_61242),
		 .Q(inst_deco[61]));
	notech_mux2 i_42991(.S(n_58449), .A(n_45615), .B(inst_deco[61]), .Z(n_36008
		));
	notech_reg_set inst_deco_reg_62(.CP(n_61803), .D(n_36014), .SD(n_61242),
		 .Q(inst_deco[62]));
	notech_mux2 i_42999(.S(n_58449), .A(n_45621), .B(inst_deco[62]), .Z(n_36014
		));
	notech_reg_set inst_deco_reg_63(.CP(n_61800), .D(n_36020), .SD(n_61242),
		 .Q(inst_deco[63]));
	notech_mux2 i_43007(.S(n_58449), .A(n_45627), .B(inst_deco[63]), .Z(n_36020
		));
	notech_reg_set inst_deco_reg_64(.CP(n_61794), .D(n_36026), .SD(n_61242),
		 .Q(inst_deco[64]));
	notech_mux2 i_43015(.S(n_58436), .A(n_45633), .B(inst_deco[64]), .Z(n_36026
		));
	notech_reg_set inst_deco_reg_65(.CP(n_61794), .D(n_36032), .SD(n_61242),
		 .Q(inst_deco[65]));
	notech_mux2 i_43023(.S(n_58436), .A(n_45639), .B(inst_deco[65]), .Z(n_36032
		));
	notech_reg_set inst_deco_reg_66(.CP(n_61794), .D(n_36038), .SD(n_61242),
		 .Q(inst_deco[66]));
	notech_mux2 i_43031(.S(n_58436), .A(n_45645), .B(inst_deco[66]), .Z(n_36038
		));
	notech_reg_set inst_deco_reg_67(.CP(n_61794), .D(n_36044), .SD(n_61233),
		 .Q(inst_deco[67]));
	notech_mux2 i_43039(.S(n_58436), .A(n_45651), .B(inst_deco[67]), .Z(n_36044
		));
	notech_reg_set inst_deco_reg_68(.CP(n_61794), .D(n_36050), .SD(n_61233),
		 .Q(inst_deco[68]));
	notech_mux2 i_43047(.S(n_58436), .A(n_45657), .B(inst_deco[68]), .Z(n_36050
		));
	notech_reg_set inst_deco_reg_69(.CP(n_61794), .D(n_36056), .SD(n_61233),
		 .Q(inst_deco[69]));
	notech_mux2 i_43055(.S(n_58436), .A(n_45663), .B(inst_deco[69]), .Z(n_36056
		));
	notech_reg_set inst_deco_reg_70(.CP(n_61794), .D(n_36062), .SD(n_61233),
		 .Q(inst_deco[70]));
	notech_mux2 i_43063(.S(n_58436), .A(n_45669), .B(inst_deco[70]), .Z(n_36062
		));
	notech_reg_set inst_deco_reg_71(.CP(n_61794), .D(n_36068), .SD(n_61233),
		 .Q(inst_deco[71]));
	notech_mux2 i_43071(.S(n_58436), .A(n_45675), .B(inst_deco[71]), .Z(n_36068
		));
	notech_reg_set inst_deco_reg_72(.CP(n_61794), .D(n_36074), .SD(n_61233),
		 .Q(inst_deco[72]));
	notech_mux2 i_43079(.S(n_58436), .A(n_3217), .B(inst_deco[72]), .Z(n_36074
		));
	notech_reg_set inst_deco_reg_73(.CP(n_61794), .D(n_36080), .SD(n_61233),
		 .Q(inst_deco[73]));
	notech_mux2 i_43087(.S(n_58436), .A(n_45687), .B(inst_deco[73]), .Z(n_36080
		));
	notech_reg_set inst_deco_reg_74(.CP(n_61794), .D(n_36086), .SD(n_61233),
		 .Q(inst_deco[74]));
	notech_mux2 i_43095(.S(n_58436), .A(n_45693), .B(inst_deco[74]), .Z(n_36086
		));
	notech_reg_set inst_deco_reg_75(.CP(n_61792), .D(n_36092), .SD(n_61233),
		 .Q(inst_deco[75]));
	notech_mux2 i_43103(.S(n_58436), .A(n_45699), .B(inst_deco[75]), .Z(n_36092
		));
	notech_reg_set inst_deco_reg_76(.CP(n_61792), .D(n_36098), .SD(n_61233),
		 .Q(inst_deco[76]));
	notech_mux2 i_43111(.S(n_58436), .A(n_45705), .B(inst_deco[76]), .Z(n_36098
		));
	notech_reg_set inst_deco_reg_77(.CP(n_61792), .D(n_36104), .SD(n_61233),
		 .Q(inst_deco[77]));
	notech_mux2 i_43119(.S(n_58436), .A(n_45711), .B(inst_deco[77]), .Z(n_36104
		));
	notech_reg_set inst_deco_reg_78(.CP(n_61792), .D(n_36110), .SD(n_61231),
		 .Q(inst_deco[78]));
	notech_mux2 i_43127(.S(n_58436), .A(n_45717), .B(inst_deco[78]), .Z(n_36110
		));
	notech_reg_set inst_deco_reg_79(.CP(n_61792), .D(n_36116), .SD(n_61231),
		 .Q(inst_deco[79]));
	notech_mux2 i_43135(.S(n_58436), .A(n_45723), .B(inst_deco[79]), .Z(n_36116
		));
	notech_reg_set inst_deco_reg_80(.CP(n_61794), .D(n_36122), .SD(n_61231),
		 .Q(inst_deco[80]));
	notech_mux2 i_43143(.S(n_58434), .A(n_45729), .B(inst_deco[80]), .Z(n_36122
		));
	notech_reg_set inst_deco_reg_81(.CP(n_61794), .D(n_36128), .SD(n_61231),
		 .Q(inst_deco[81]));
	notech_mux2 i_43151(.S(n_58434), .A(n_45735), .B(inst_deco[81]), .Z(n_36128
		));
	notech_reg_set inst_deco_reg_82(.CP(n_61794), .D(n_36134), .SD(n_61231),
		 .Q(inst_deco[82]));
	notech_mux2 i_43159(.S(n_58434), .A(n_3216), .B(inst_deco[82]), .Z(n_36134
		));
	notech_reg_set inst_deco_reg_83(.CP(n_61794), .D(n_36140), .SD(n_61233),
		 .Q(inst_deco[83]));
	notech_mux2 i_43167(.S(n_58434), .A(n_3215), .B(inst_deco[83]), .Z(n_36140
		));
	notech_reg_set inst_deco_reg_84(.CP(n_61794), .D(n_36146), .SD(n_61233),
		 .Q(inst_deco[84]));
	notech_mux2 i_43175(.S(n_58434), .A(n_3214), .B(inst_deco[84]), .Z(n_36146
		));
	notech_reg_set inst_deco_reg_85(.CP(n_61798), .D(n_36152), .SD(n_61233),
		 .Q(inst_deco[85]));
	notech_mux2 i_43183(.S(n_58434), .A(n_3213), .B(inst_deco[85]), .Z(n_36152
		));
	notech_reg_set inst_deco_reg_86(.CP(n_61798), .D(n_36158), .SD(n_61233),
		 .Q(inst_deco[86]));
	notech_mux2 i_43191(.S(n_58434), .A(n_45765), .B(inst_deco[86]), .Z(n_36158
		));
	notech_reg_set inst_deco_reg_87(.CP(n_61798), .D(n_36164), .SD(n_61233),
		 .Q(inst_deco[87]));
	notech_mux2 i_43199(.S(n_58434), .A(n_3212), .B(inst_deco[87]), .Z(n_36164
		));
	notech_reg_set inst_deco_reg_88(.CP(n_61798), .D(n_36170), .SD(n_61237),
		 .Q(inst_deco[88]));
	notech_mux2 i_43207(.S(n_58434), .A(n_45777), .B(inst_deco[88]), .Z(n_36170
		));
	notech_reg_set inst_deco_reg_89(.CP(n_61798), .D(n_36176), .SD(n_61237),
		 .Q(inst_deco[89]));
	notech_mux2 i_43215(.S(n_58434), .A(n_45783), .B(inst_deco[89]), .Z(n_36176
		));
	notech_reg_set inst_deco_reg_90(.CP(n_61798), .D(n_36182), .SD(n_61237),
		 .Q(inst_deco[90]));
	notech_mux2 i_43223(.S(n_58434), .A(n_45789), .B(inst_deco[90]), .Z(n_36182
		));
	notech_reg_set inst_deco_reg_91(.CP(n_61800), .D(n_36188), .SD(n_61237),
		 .Q(inst_deco[91]));
	notech_mux2 i_43231(.S(n_58434), .A(n_45795), .B(inst_deco[91]), .Z(n_36188
		));
	notech_reg_set inst_deco_reg_92(.CP(n_61798), .D(n_36194), .SD(n_61237),
		 .Q(inst_deco[92]));
	notech_mux2 i_43239(.S(n_58434), .A(n_3211), .B(inst_deco[92]), .Z(n_36194
		));
	notech_reg_set inst_deco_reg_93(.CP(n_61798), .D(n_36200), .SD(n_61237),
		 .Q(inst_deco[93]));
	notech_mux2 i_43247(.S(n_58434), .A(n_3210), .B(inst_deco[93]), .Z(n_36200
		));
	notech_reg_set inst_deco_reg_94(.CP(n_61798), .D(n_36206), .SD(n_61239),
		 .Q(inst_deco[94]));
	notech_mux2 i_43255(.S(n_58434), .A(n_3209), .B(inst_deco[94]), .Z(n_36206
		));
	notech_reg_set inst_deco_reg_95(.CP(n_61798), .D(n_36212), .SD(n_61237),
		 .Q(inst_deco[95]));
	notech_mux2 i_43263(.S(n_58434), .A(n_45819), .B(inst_deco[95]), .Z(n_36212
		));
	notech_reg_set inst_deco_reg_96(.CP(n_61798), .D(n_36218), .SD(n_61237),
		 .Q(inst_deco[96]));
	notech_mux2 i_43271(.S(n_58441), .A(n_3208), .B(inst_deco[96]), .Z(n_36218
		));
	notech_reg_set inst_deco_reg_97(.CP(n_61798), .D(n_36224), .SD(n_61237),
		 .Q(inst_deco[97]));
	notech_mux2 i_43279(.S(n_58441), .A(n_3207), .B(inst_deco[97]), .Z(n_36224
		));
	notech_reg_set inst_deco_reg_98(.CP(n_61798), .D(n_36230), .SD(n_61237),
		 .Q(inst_deco[98]));
	notech_mux2 i_43287(.S(n_58441), .A(n_45837), .B(inst_deco[98]), .Z(n_36230
		));
	notech_reg_set inst_deco_reg_99(.CP(n_61794), .D(n_36236), .SD(n_61237),
		 .Q(inst_deco[99]));
	notech_mux2 i_43295(.S(n_58441), .A(n_3206), .B(inst_deco[99]), .Z(n_36236
		));
	notech_reg_set inst_deco_reg_100(.CP(n_61794), .D(n_36242), .SD(n_61237)
		, .Q(inst_deco[100]));
	notech_mux2 i_43303(.S(n_58441), .A(n_45849), .B(inst_deco[100]), .Z(n_36242
		));
	notech_reg_set inst_deco_reg_101(.CP(n_61798), .D(n_36248), .SD(n_61237)
		, .Q(inst_deco[101]));
	notech_mux2 i_43311(.S(n_58441), .A(n_45855), .B(inst_deco[101]), .Z(n_36248
		));
	notech_reg_set inst_deco_reg_102(.CP(n_61798), .D(n_36254), .SD(n_61233)
		, .Q(inst_deco[102]));
	notech_mux2 i_43319(.S(n_58441), .A(n_45861), .B(inst_deco[102]), .Z(n_36254
		));
	notech_reg_set inst_deco_reg_103(.CP(n_61798), .D(n_36260), .SD(n_61233)
		, .Q(inst_deco[103]));
	notech_mux2 i_43327(.S(n_58441), .A(n_45867), .B(inst_deco[103]), .Z(n_36260
		));
	notech_reg_set inst_deco_reg_104(.CP(n_61798), .D(n_36266), .SD(n_61237)
		, .Q(inst_deco[104]));
	notech_mux2 i_43335(.S(n_58441), .A(n_45873), .B(inst_deco[104]), .Z(n_36266
		));
	notech_reg_set inst_deco_reg_105(.CP(n_61798), .D(n_36272), .SD(n_61237)
		, .Q(inst_deco[105]));
	notech_mux2 i_43343(.S(n_58441), .A(n_45879), .B(inst_deco[105]), .Z(n_36272
		));
	notech_reg_set inst_deco_reg_106(.CP(n_61830), .D(n_36278), .SD(n_61237)
		, .Q(inst_deco[106]));
	notech_mux2 i_43351(.S(n_58441), .A(n_45885), .B(inst_deco[106]), .Z(n_36278
		));
	notech_reg_set inst_deco_reg_107(.CP(n_61865), .D(n_36284), .SD(n_61237)
		, .Q(inst_deco[107]));
	notech_mux2 i_43359(.S(n_58441), .A(n_45891), .B(inst_deco[107]), .Z(n_36284
		));
	notech_reg_set inst_deco_reg_108(.CP(n_61865), .D(n_36290), .SD(n_61237)
		, .Q(inst_deco[108]));
	notech_mux2 i_43367(.S(n_58441), .A(n_45897), .B(inst_deco[108]), .Z(n_36290
		));
	notech_reg_set inst_deco_reg_109(.CP(n_61865), .D(n_36296), .SD(n_61304)
		, .Q(inst_deco[109]));
	notech_mux2 i_43375(.S(n_58441), .A(n_45903), .B(inst_deco[109]), .Z(n_36296
		));
	notech_reg_set inst_deco_reg_110(.CP(n_61865), .D(n_36302), .SD(n_61304)
		, .Q(inst_deco[110]));
	notech_mux2 i_43383(.S(n_58441), .A(n_45909), .B(inst_deco[110]), .Z(n_36302
		));
	notech_reg_set inst_deco_reg_111(.CP(n_61865), .D(n_36308), .SD(n_61304)
		, .Q(inst_deco[111]));
	notech_mux2 i_43391(.S(n_58441), .A(n_45915), .B(inst_deco[111]), .Z(n_36308
		));
	notech_reg_set inst_deco_reg_112(.CP(n_61865), .D(n_36314), .SD(n_61304)
		, .Q(inst_deco[112]));
	notech_mux2 i_43399(.S(n_58439), .A(n_45921), .B(inst_deco[112]), .Z(n_36314
		));
	notech_reg_set inst_deco_reg_113(.CP(n_61865), .D(n_36320), .SD(n_61304)
		, .Q(inst_deco[113]));
	notech_mux2 i_43407(.S(n_58439), .A(n_39358), .B(inst_deco[113]), .Z(n_36320
		));
	notech_reg_set inst_deco_reg_114(.CP(n_61865), .D(n_36326), .SD(n_61304)
		, .Q(inst_deco[114]));
	notech_mux2 i_43415(.S(n_58439), .A(n_3204), .B(inst_deco[114]), .Z(n_36326
		));
	notech_reg_set inst_deco_reg_115(.CP(n_61865), .D(n_36332), .SD(n_61304)
		, .Q(inst_deco[115]));
	notech_mux2 i_43423(.S(n_58439), .A(n_3203), .B(inst_deco[115]), .Z(n_36332
		));
	notech_reg_set inst_deco_reg_116(.CP(n_61865), .D(n_36338), .SD(n_61304)
		, .Q(inst_deco[116]));
	notech_mux2 i_43431(.S(n_58439), .A(n_45945), .B(inst_deco[116]), .Z(n_36338
		));
	notech_reg_set inst_deco_reg_117(.CP(n_61865), .D(n_36344), .SD(n_61304)
		, .Q(inst_deco[117]));
	notech_mux2 i_43439(.S(n_58439), .A(n_45951), .B(inst_deco[117]), .Z(n_36344
		));
	notech_reg_set inst_deco_reg_118(.CP(n_61863), .D(n_36350), .SD(n_61304)
		, .Q(inst_deco[118]));
	notech_mux2 i_43447(.S(n_58439), .A(n_45957), .B(inst_deco[118]), .Z(n_36350
		));
	notech_reg_set inst_deco_reg_119(.CP(n_61865), .D(n_36356), .SD(n_61304)
		, .Q(inst_deco[119]));
	notech_mux2 i_43455(.S(n_58439), .A(n_45963), .B(inst_deco[119]), .Z(n_36356
		));
	notech_reg_set inst_deco_reg_120(.CP(n_61863), .D(n_36362), .SD(n_61302)
		, .Q(inst_deco[120]));
	notech_mux2 i_43463(.S(n_58439), .A(n_45969), .B(inst_deco[120]), .Z(n_36362
		));
	notech_reg_set inst_deco_reg_121(.CP(n_61863), .D(n_36368), .SD(n_61302)
		, .Q(inst_deco[121]));
	notech_mux2 i_43471(.S(n_58439), .A(n_45975), .B(inst_deco[121]), .Z(n_36368
		));
	notech_reg_set inst_deco_reg_122(.CP(n_61863), .D(n_36374), .SD(n_61302)
		, .Q(inst_deco[122]));
	notech_mux2 i_43479(.S(n_58439), .A(n_45981), .B(inst_deco[122]), .Z(n_36374
		));
	notech_reg_set inst_deco_reg_123(.CP(n_61865), .D(n_36380), .SD(n_61302)
		, .Q(inst_deco[123]));
	notech_mux2 i_43487(.S(n_58439), .A(n_45987), .B(inst_deco[123]), .Z(n_36380
		));
	notech_reg_set inst_deco_reg_124(.CP(n_61865), .D(n_36386), .SD(n_61302)
		, .Q(inst_deco[124]));
	notech_mux2 i_43495(.S(n_58439), .A(n_45993), .B(inst_deco[124]), .Z(n_36386
		));
	notech_reg_set inst_deco_reg_125(.CP(n_61865), .D(n_36392), .SD(n_61304)
		, .Q(inst_deco[125]));
	notech_mux2 i_43503(.S(n_58439), .A(n_45999), .B(inst_deco[125]), .Z(n_36392
		));
	notech_reg_set inst_deco_reg_126(.CP(n_61865), .D(n_36398), .SD(n_61304)
		, .Q(inst_deco[126]));
	notech_mux2 i_43511(.S(n_58439), .A(n_46005), .B(inst_deco[126]), .Z(n_36398
		));
	notech_reg_set inst_deco_reg_127(.CP(n_61865), .D(n_36404), .SD(n_61304)
		, .Q(inst_deco[127]));
	notech_mux2 i_43519(.S(n_58439), .A(n_46011), .B(inst_deco[127]), .Z(n_36404
		));
	notech_reg pfx_sz_reg_0(.CP(n_61868), .D(n_36410), .CD(n_61302), .Q(pfx_sz
		[0]));
	notech_mux2 i_43527(.S(\nbus_13541[0] ), .A(pfx_sz[0]), .B(n_38411), .Z(n_36410
		));
	notech_reg pfx_sz_reg_1(.CP(n_61868), .D(n_36416), .CD(n_61302), .Q(pfx_sz
		[1]));
	notech_mux2 i_43535(.S(\nbus_13541[0] ), .A(pfx_sz[1]), .B(n_39827), .Z(n_36416
		));
	notech_reg pfx_sz_reg_2(.CP(n_61868), .D(n_36422), .CD(n_61307), .Q(pfx_sz
		[2]));
	notech_mux2 i_43543(.S(\nbus_13541[0] ), .A(pfx_sz[2]), .B(n_170993330),
		 .Z(n_36422));
	notech_reg pfx_sz_reg_3(.CP(n_61868), .D(n_36428), .CD(n_61307), .Q(pfx_sz
		[3]));
	notech_mux2 i_43551(.S(\nbus_13541[0] ), .A(pfx_sz[3]), .B(n_171093331),
		 .Z(n_36428));
	notech_reg pfx_sz_reg_4(.CP(n_61868), .D(n_36434), .CD(n_61307), .Q(pfx_sz
		[4]));
	notech_mux2 i_43559(.S(\nbus_13541[0] ), .A(pfx_sz[4]), .B(n_171193332),
		 .Z(n_36434));
	notech_reg lenpc2_reg_0(.CP(n_61870), .D(n_36440), .CD(n_61307), .Q(lenpc2
		[0]));
	notech_mux2 i_43567(.S(n_54198), .A(lenpc2[0]), .B(n_3244), .Z(n_36440)
		);
	notech_reg lenpc2_reg_1(.CP(n_61870), .D(n_36446), .CD(n_61307), .Q(lenpc2
		[1]));
	notech_mux2 i_43575(.S(n_54198), .A(lenpc2[1]), .B(n_3242), .Z(n_36446)
		);
	notech_reg lenpc2_reg_2(.CP(n_61868), .D(n_36452), .CD(n_61307), .Q(lenpc2
		[2]));
	notech_mux2 i_43583(.S(n_54198), .A(lenpc2[2]), .B(n_45035), .Z(n_36452)
		);
	notech_reg lenpc2_reg_3(.CP(n_61868), .D(n_36458), .CD(n_61307), .Q(lenpc2
		[3]));
	notech_mux2 i_43591(.S(n_54198), .A(lenpc2[3]), .B(n_2057), .Z(n_36458)
		);
	notech_reg lenpc2_reg_4(.CP(n_61868), .D(n_36464), .CD(n_61307), .Q(lenpc2
		[4]));
	notech_mux2 i_43599(.S(n_54198), .A(lenpc2[4]), .B(n_3239), .Z(n_36464)
		);
	notech_reg lenpc2_reg_5(.CP(n_61868), .D(n_36470), .CD(n_61307), .Q(lenpc2
		[5]));
	notech_mux2 i_43607(.S(n_54199), .A(lenpc2[5]), .B(n_3237), .Z(n_36470)
		);
	notech_reg lenpc2_reg_6(.CP(n_61868), .D(n_36480), .CD(n_61307), .Q(lenpc2
		[6]));
	notech_ao3 i_43619(.A(lenpc2[6]), .B(1'b1), .C(n_54210), .Z(n_36480));
	notech_reg lenpc2_reg_7(.CP(n_61868), .D(n_36486), .CD(n_61307), .Q(lenpc2
		[7]));
	notech_ao3 i_43627(.A(lenpc2[7]), .B(1'b1), .C(n_54210), .Z(n_36486));
	notech_reg lenpc2_reg_8(.CP(n_61868), .D(n_36492), .CD(n_61304), .Q(lenpc2
		[8]));
	notech_ao3 i_43635(.A(lenpc2[8]), .B(1'b1), .C(n_54210), .Z(n_36492));
	notech_reg lenpc2_reg_9(.CP(n_61865), .D(n_36498), .CD(n_61307), .Q(lenpc2
		[9]));
	notech_ao3 i_43643(.A(lenpc2[9]), .B(1'b1), .C(n_54205), .Z(n_36498));
	notech_reg lenpc2_reg_10(.CP(n_61868), .D(n_36504), .CD(n_61304), .Q(lenpc2
		[10]));
	notech_ao3 i_43651(.A(lenpc2[10]), .B(1'b1), .C(n_54205), .Z(n_36504));
	notech_reg lenpc2_reg_11(.CP(n_61868), .D(n_36510), .CD(n_61304), .Q(lenpc2
		[11]));
	notech_ao3 i_43659(.A(lenpc2[11]), .B(1'b1), .C(n_54205), .Z(n_36510));
	notech_reg lenpc2_reg_12(.CP(n_61868), .D(n_36516), .CD(n_61304), .Q(lenpc2
		[12]));
	notech_ao3 i_43667(.A(lenpc2[12]), .B(1'b1), .C(n_54210), .Z(n_36516));
	notech_reg lenpc2_reg_13(.CP(n_61868), .D(n_36522), .CD(n_61307), .Q(lenpc2
		[13]));
	notech_ao3 i_43675(.A(lenpc2[13]), .B(1'b1), .C(n_54210), .Z(n_36522));
	notech_reg lenpc2_reg_14(.CP(n_61868), .D(n_36528), .CD(n_61307), .Q(lenpc2
		[14]));
	notech_ao3 i_43683(.A(lenpc2[14]), .B(1'b1), .C(n_54210), .Z(n_36528));
	notech_reg lenpc2_reg_15(.CP(n_61868), .D(n_36534), .CD(n_61307), .Q(lenpc2
		[15]));
	notech_ao3 i_43691(.A(lenpc2[15]), .B(1'b1), .C(n_54210), .Z(n_36534));
	notech_reg lenpc2_reg_16(.CP(n_61863), .D(n_36540), .CD(n_61307), .Q(lenpc2
		[16]));
	notech_ao3 i_43699(.A(lenpc2[16]), .B(1'b1), .C(n_54210), .Z(n_36540));
	notech_reg lenpc2_reg_17(.CP(n_61859), .D(n_36546), .CD(n_61307), .Q(lenpc2
		[17]));
	notech_ao3 i_43707(.A(lenpc2[17]), .B(1'b1), .C(n_54210), .Z(n_36546));
	notech_reg lenpc2_reg_18(.CP(n_61859), .D(n_36552), .CD(n_61298), .Q(lenpc2
		[18]));
	notech_ao3 i_43715(.A(lenpc2[18]), .B(1'b1), .C(n_54210), .Z(n_36552));
	notech_reg lenpc2_reg_19(.CP(n_61859), .D(n_36558), .CD(n_61298), .Q(lenpc2
		[19]));
	notech_ao3 i_43723(.A(lenpc2[19]), .B(1'b1), .C(n_54199), .Z(n_36558));
	notech_reg lenpc2_reg_20(.CP(n_61859), .D(n_36564), .CD(n_61298), .Q(lenpc2
		[20]));
	notech_ao3 i_43731(.A(lenpc2[20]), .B(1'b1), .C(n_54205), .Z(n_36564));
	notech_reg lenpc2_reg_21(.CP(n_61859), .D(n_36570), .CD(n_61296), .Q(lenpc2
		[21]));
	notech_ao3 i_43739(.A(lenpc2[21]), .B(1'b1), .C(n_54205), .Z(n_36570));
	notech_reg lenpc2_reg_22(.CP(n_61859), .D(n_36576), .CD(n_61296), .Q(lenpc2
		[22]));
	notech_ao3 i_43747(.A(lenpc2[22]), .B(1'b1), .C(n_54199), .Z(n_36576));
	notech_reg lenpc2_reg_23(.CP(n_61859), .D(n_36582), .CD(n_61298), .Q(lenpc2
		[23]));
	notech_ao3 i_43755(.A(lenpc2[23]), .B(1'b1), .C(n_54199), .Z(n_36582));
	notech_reg lenpc2_reg_24(.CP(n_61859), .D(n_36588), .CD(n_61298), .Q(lenpc2
		[24]));
	notech_ao3 i_43763(.A(lenpc2[24]), .B(1'b1), .C(n_54199), .Z(n_36588));
	notech_reg lenpc2_reg_25(.CP(n_61859), .D(n_36594), .CD(n_61298), .Q(lenpc2
		[25]));
	notech_ao3 i_43771(.A(lenpc2[25]), .B(1'b1), .C(n_54205), .Z(n_36594));
	notech_reg lenpc2_reg_26(.CP(n_61859), .D(n_36600), .CD(n_61298), .Q(lenpc2
		[26]));
	notech_ao3 i_43779(.A(lenpc2[26]), .B(1'b1), .C(n_54205), .Z(n_36600));
	notech_reg lenpc2_reg_27(.CP(n_61857), .D(n_36606), .CD(n_61298), .Q(lenpc2
		[27]));
	notech_ao3 i_43787(.A(lenpc2[27]), .B(1'b1), .C(n_54205), .Z(n_36606));
	notech_reg lenpc2_reg_28(.CP(n_61857), .D(n_36612), .CD(n_61296), .Q(lenpc2
		[28]));
	notech_ao3 i_43795(.A(lenpc2[28]), .B(1'b1), .C(n_54205), .Z(n_36612));
	notech_reg lenpc2_reg_29(.CP(n_61857), .D(n_36618), .CD(n_61296), .Q(lenpc2
		[29]));
	notech_ao3 i_43803(.A(lenpc2[29]), .B(1'b1), .C(n_54205), .Z(n_36618));
	notech_reg lenpc2_reg_30(.CP(n_61857), .D(n_36624), .CD(n_61296), .Q(lenpc2
		[30]));
	notech_ao3 i_43811(.A(lenpc2[30]), .B(1'b1), .C(n_54205), .Z(n_36624));
	notech_reg lenpc2_reg_31(.CP(n_61857), .D(n_36630), .CD(n_61296), .Q(lenpc2
		[31]));
	notech_ao3 i_43819(.A(lenpc2[31]), .B(1'b1), .C(n_54205), .Z(n_36630));
	notech_reg lenpc1_reg_0(.CP(n_61857), .D(n_36632), .CD(n_61296), .Q(lenpc1
		[0]));
	notech_mux2 i_43823(.S(n_57620), .A(lenpc1[0]), .B(n_39313), .Z(n_36632)
		);
	notech_reg lenpc1_reg_1(.CP(n_61857), .D(n_36638), .CD(n_61296), .Q(lenpc1
		[1]));
	notech_mux2 i_43831(.S(n_57620), .A(lenpc1[1]), .B(n_39316), .Z(n_36638)
		);
	notech_reg lenpc1_reg_2(.CP(n_61857), .D(n_36644), .CD(n_61296), .Q(lenpc1
		[2]));
	notech_mux2 i_43839(.S(n_57620), .A(lenpc1[2]), .B(n_39319), .Z(n_36644)
		);
	notech_reg lenpc1_reg_3(.CP(n_61857), .D(n_36650), .CD(n_61296), .Q(lenpc1
		[3]));
	notech_mux2 i_43847(.S(n_57620), .A(lenpc1[3]), .B(n_38395), .Z(n_36650)
		);
	notech_reg lenpc1_reg_4(.CP(n_61857), .D(n_36656), .CD(n_61296), .Q(lenpc1
		[4]));
	notech_mux2 i_43855(.S(n_57620), .A(lenpc1[4]), .B(n_39322), .Z(n_36656)
		);
	notech_reg lenpc1_reg_5(.CP(n_61857), .D(n_36662), .CD(n_61296), .Q(lenpc1
		[5]));
	notech_mux2 i_43863(.S(n_57621), .A(lenpc1[5]), .B(n_39325), .Z(n_36662)
		);
	notech_reg lenpc1_reg_6(.CP(n_61863), .D(n_36668), .CD(n_61296), .Q(lenpc1
		[6]));
	notech_mux2 i_43871(.S(n_57632), .A(lenpc1[6]), .B(n_44398), .Z(n_36668)
		);
	notech_reg lenpc1_reg_7(.CP(n_61863), .D(n_36674), .CD(n_61302), .Q(lenpc1
		[7]));
	notech_mux2 i_43879(.S(n_57632), .A(lenpc1[7]), .B(n_44404), .Z(n_36674)
		);
	notech_reg lenpc1_reg_8(.CP(n_61863), .D(n_36680), .CD(n_61302), .Q(lenpc1
		[8]));
	notech_mux2 i_43887(.S(n_57632), .A(lenpc1[8]), .B(n_44410), .Z(n_36680)
		);
	notech_reg lenpc1_reg_9(.CP(n_61863), .D(n_36686), .CD(n_61302), .Q(lenpc1
		[9]));
	notech_mux2 i_43895(.S(n_57627), .A(lenpc1[9]), .B(n_44416), .Z(n_36686)
		);
	notech_reg lenpc1_reg_10(.CP(n_61863), .D(n_36692), .CD(n_61302), .Q(lenpc1
		[10]));
	notech_mux2 i_43903(.S(n_57627), .A(lenpc1[10]), .B(n_44422), .Z(n_36692
		));
	notech_reg lenpc1_reg_11(.CP(n_61863), .D(n_36698), .CD(n_61302), .Q(lenpc1
		[11]));
	notech_mux2 i_43911(.S(n_57627), .A(lenpc1[11]), .B(n_44428), .Z(n_36698
		));
	notech_reg lenpc1_reg_12(.CP(n_61863), .D(n_36704), .CD(n_61302), .Q(lenpc1
		[12]));
	notech_mux2 i_43919(.S(n_57632), .A(lenpc1[12]), .B(n_44434), .Z(n_36704
		));
	notech_reg lenpc1_reg_13(.CP(n_61863), .D(n_36710), .CD(n_61302), .Q(lenpc1
		[13]));
	notech_mux2 i_43927(.S(n_57632), .A(lenpc1[13]), .B(n_44440), .Z(n_36710
		));
	notech_reg lenpc1_reg_14(.CP(n_61863), .D(n_36716), .CD(n_61302), .Q(lenpc1
		[14]));
	notech_mux2 i_43935(.S(n_57632), .A(lenpc1[14]), .B(n_44446), .Z(n_36716
		));
	notech_reg lenpc1_reg_15(.CP(n_61863), .D(n_36722), .CD(n_61302), .Q(lenpc1
		[15]));
	notech_mux2 i_43943(.S(n_57632), .A(lenpc1[15]), .B(n_44452), .Z(n_36722
		));
	notech_reg lenpc1_reg_16(.CP(n_61863), .D(n_36728), .CD(n_61302), .Q(lenpc1
		[16]));
	notech_mux2 i_43951(.S(n_57632), .A(lenpc1[16]), .B(n_44458), .Z(n_36728
		));
	notech_reg lenpc1_reg_17(.CP(n_61859), .D(n_36734), .CD(n_61302), .Q(lenpc1
		[17]));
	notech_mux2 i_43959(.S(n_57632), .A(lenpc1[17]), .B(n_44464), .Z(n_36734
		));
	notech_reg lenpc1_reg_18(.CP(n_61859), .D(n_36740), .CD(n_61298), .Q(lenpc1
		[18]));
	notech_mux2 i_43967(.S(n_57632), .A(lenpc1[18]), .B(n_44470), .Z(n_36740
		));
	notech_reg lenpc1_reg_19(.CP(n_61859), .D(n_36746), .CD(n_61298), .Q(lenpc1
		[19]));
	notech_mux2 i_43975(.S(n_57621), .A(lenpc1[19]), .B(n_44476), .Z(n_36746
		));
	notech_reg lenpc1_reg_20(.CP(n_61859), .D(n_36752), .CD(n_61298), .Q(lenpc1
		[20]));
	notech_mux2 i_43983(.S(n_57627), .A(lenpc1[20]), .B(n_44482), .Z(n_36752
		));
	notech_reg lenpc1_reg_21(.CP(n_61859), .D(n_36758), .CD(n_61298), .Q(lenpc1
		[21]));
	notech_mux2 i_43991(.S(n_57627), .A(lenpc1[21]), .B(n_110792728), .Z(n_36758
		));
	notech_reg lenpc1_reg_22(.CP(n_61863), .D(n_36764), .CD(n_61298), .Q(lenpc1
		[22]));
	notech_mux2 i_43999(.S(n_57621), .A(lenpc1[22]), .B(n_110892729), .Z(n_36764
		));
	notech_reg lenpc1_reg_23(.CP(n_61863), .D(n_36770), .CD(n_61298), .Q(lenpc1
		[23]));
	notech_mux2 i_44007(.S(n_57621), .A(lenpc1[23]), .B(n_110992730), .Z(n_36770
		));
	notech_reg lenpc1_reg_24(.CP(n_61859), .D(n_36776), .CD(n_61298), .Q(lenpc1
		[24]));
	notech_mux2 i_44015(.S(n_57621), .A(lenpc1[24]), .B(n_111092731), .Z(n_36776
		));
	notech_reg lenpc1_reg_25(.CP(n_61859), .D(n_36782), .CD(n_61298), .Q(lenpc1
		[25]));
	notech_mux2 i_44023(.S(n_57627), .A(lenpc1[25]), .B(n_111192732), .Z(n_36782
		));
	notech_reg lenpc1_reg_26(.CP(n_61859), .D(n_36788), .CD(n_61298), .Q(lenpc1
		[26]));
	notech_mux2 i_44031(.S(n_57627), .A(lenpc1[26]), .B(n_111292733), .Z(n_36788
		));
	notech_reg lenpc1_reg_27(.CP(n_61879), .D(n_36794), .CD(n_61298), .Q(lenpc1
		[27]));
	notech_mux2 i_44039(.S(n_57627), .A(lenpc1[27]), .B(n_44524), .Z(n_36794
		));
	notech_reg lenpc1_reg_28(.CP(n_61879), .D(n_36800), .CD(n_61307), .Q(lenpc1
		[28]));
	notech_mux2 i_44047(.S(n_57627), .A(lenpc1[28]), .B(n_44530), .Z(n_36800
		));
	notech_reg lenpc1_reg_29(.CP(n_61879), .D(n_36806), .CD(n_61318), .Q(lenpc1
		[29]));
	notech_mux2 i_44055(.S(n_57627), .A(lenpc1[29]), .B(n_44536), .Z(n_36806
		));
	notech_reg lenpc1_reg_30(.CP(n_61879), .D(n_36812), .CD(n_61318), .Q(lenpc1
		[30]));
	notech_mux2 i_44063(.S(n_57627), .A(lenpc1[30]), .B(n_44542), .Z(n_36812
		));
	notech_reg lenpc1_reg_31(.CP(n_61879), .D(n_36818), .CD(n_61318), .Q(lenpc1
		[31]));
	notech_mux2 i_44071(.S(n_57627), .A(lenpc1[31]), .B(n_44548), .Z(n_36818
		));
	notech_reg to_acu0_reg_0(.CP(n_61879), .D(n_36824), .CD(n_61318), .Q(to_acu0
		[0]));
	notech_mux2 i_44079(.S(n_54998), .A(to_acu0[0]), .B(n_38521), .Z(n_36824
		));
	notech_reg to_acu0_reg_1(.CP(n_61879), .D(n_36830), .CD(n_61318), .Q(to_acu0
		[1]));
	notech_mux2 i_44087(.S(n_55003), .A(to_acu0[1]), .B(n_38523), .Z(n_36830
		));
	notech_reg to_acu0_reg_2(.CP(n_61879), .D(n_36836), .CD(n_61318), .Q(to_acu0
		[2]));
	notech_mux2 i_44095(.S(n_55003), .A(to_acu0[2]), .B(n_38525), .Z(n_36836
		));
	notech_reg to_acu0_reg_3(.CP(n_61879), .D(n_36842), .CD(n_61318), .Q(to_acu0
		[3]));
	notech_mux2 i_44103(.S(n_54983), .A(to_acu0[3]), .B(n_38527), .Z(n_36842
		));
	notech_reg to_acu0_reg_4(.CP(n_61879), .D(n_36848), .CD(n_61318), .Q(to_acu0
		[4]));
	notech_mux2 i_44111(.S(n_55003), .A(to_acu0[4]), .B(n_38529), .Z(n_36848
		));
	notech_reg to_acu0_reg_5(.CP(n_61879), .D(n_36854), .CD(n_61318), .Q(to_acu0
		[5]));
	notech_mux2 i_44119(.S(n_55003), .A(to_acu0[5]), .B(n_38531), .Z(n_36854
		));
	notech_reg to_acu0_reg_6(.CP(n_61875), .D(n_36860), .CD(n_61318), .Q(to_acu0
		[6]));
	notech_mux2 i_44127(.S(n_54983), .A(to_acu0[6]), .B(n_38533), .Z(n_36860
		));
	notech_reg to_acu0_reg_7(.CP(n_61875), .D(n_36866), .CD(n_61314), .Q(to_acu0
		[7]));
	notech_mux2 i_44135(.S(n_54983), .A(to_acu0[7]), .B(n_38535), .Z(n_36866
		));
	notech_reg to_acu0_reg_8(.CP(n_61875), .D(n_36872), .CD(n_61314), .Q(to_acu0
		[8]));
	notech_mux2 i_44143(.S(n_54983), .A(to_acu0[8]), .B(n_38537), .Z(n_36872
		));
	notech_reg to_acu0_reg_9(.CP(n_61875), .D(n_36878), .CD(n_61314), .Q(to_acu0
		[9]));
	notech_mux2 i_44151(.S(n_54983), .A(to_acu0[9]), .B(n_38539), .Z(n_36878
		));
	notech_ao4 i_129473717(.A(n_58394), .B(n_38882), .C(n_58465), .D(n_39867
		), .Z(n_1621));
	notech_reg to_acu0_reg_10(.CP(n_61875), .D(n_36884), .CD(n_61314), .Q(to_acu0
		[10]));
	notech_mux2 i_44159(.S(n_55003), .A(to_acu0[10]), .B(n_38541), .Z(n_36884
		));
	notech_ao4 i_129773714(.A(n_58394), .B(n_38888), .C(n_58467), .D(n_39870
		), .Z(n_1620));
	notech_reg to_acu0_reg_11(.CP(n_61875), .D(n_36890), .CD(n_61314), .Q(to_acu0
		[11]));
	notech_mux2 i_44167(.S(n_55003), .A(to_acu0[11]), .B(n_38543), .Z(n_36890
		));
	notech_ao4 i_129973712(.A(n_58394), .B(n_38892), .C(n_58470), .D(n_39872
		), .Z(n_1619));
	notech_reg to_acu0_reg_12(.CP(n_61879), .D(n_36896), .CD(n_61314), .Q(to_acu0
		[12]));
	notech_mux2 i_44175(.S(n_55003), .A(to_acu0[12]), .B(n_38545), .Z(n_36896
		));
	notech_ao4 i_130073711(.A(n_58394), .B(n_38894), .C(n_58470), .D(n_39873
		), .Z(n_1618));
	notech_reg to_acu0_reg_13(.CP(n_61875), .D(n_36902), .CD(n_61314), .Q(to_acu0
		[13]));
	notech_mux2 i_44183(.S(n_55003), .A(to_acu0[13]), .B(n_38547), .Z(n_36902
		));
	notech_ao4 i_130173710(.A(n_58394), .B(n_38896), .C(n_58470), .D(n_39874
		), .Z(n_1617));
	notech_reg to_acu0_reg_14(.CP(n_61875), .D(n_36908), .CD(n_61314), .Q(to_acu0
		[14]));
	notech_mux2 i_44191(.S(n_55003), .A(to_acu0[14]), .B(n_38549), .Z(n_36908
		));
	notech_ao4 i_130273709(.A(n_58396), .B(n_38899), .C(n_58470), .D(n_39876
		), .Z(n_1616));
	notech_reg to_acu0_reg_15(.CP(n_61875), .D(n_36914), .CD(n_61314), .Q(to_acu0
		[15]));
	notech_mux2 i_44199(.S(n_55003), .A(to_acu0[15]), .B(n_38551), .Z(n_36914
		));
	notech_ao4 i_130373708(.A(n_58396), .B(n_38901), .C(n_58470), .D(n_39877
		), .Z(n_1615));
	notech_reg to_acu0_reg_16(.CP(n_61881), .D(n_36920), .CD(n_61314), .Q(to_acu0
		[16]));
	notech_mux2 i_44207(.S(n_55003), .A(to_acu0[16]), .B(n_38553), .Z(n_36920
		));
	notech_ao4 i_130473707(.A(n_58396), .B(n_38903), .C(n_58470), .D(n_39878
		), .Z(n_1614));
	notech_reg to_acu0_reg_17(.CP(n_61881), .D(n_36926), .CD(n_61314), .Q(to_acu0
		[17]));
	notech_mux2 i_44215(.S(n_55003), .A(to_acu0[17]), .B(n_38555), .Z(n_36926
		));
	notech_ao4 i_130573706(.A(n_58396), .B(n_38905), .C(n_58470), .D(n_39879
		), .Z(n_1613));
	notech_reg to_acu0_reg_18(.CP(n_61881), .D(n_36932), .CD(n_61320), .Q(to_acu0
		[18]));
	notech_mux2 i_44223(.S(n_55017), .A(to_acu0[18]), .B(n_38557), .Z(n_36932
		));
	notech_ao4 i_130673705(.A(n_58394), .B(n_38907), .C(n_58470), .D(n_39880
		), .Z(n_1612));
	notech_reg to_acu0_reg_19(.CP(n_61881), .D(n_36938), .CD(n_61320), .Q(to_acu0
		[19]));
	notech_mux2 i_44231(.S(n_55031), .A(to_acu0[19]), .B(n_38340), .Z(n_36938
		));
	notech_ao4 i_130773704(.A(n_58394), .B(n_38909), .C(n_58472), .D(n_39881
		), .Z(n_1611));
	notech_reg to_acu0_reg_20(.CP(n_61881), .D(n_36944), .CD(n_61320), .Q(to_acu0
		[20]));
	notech_mux2 i_44239(.S(n_55031), .A(to_acu0[20]), .B(n_38559), .Z(n_36944
		));
	notech_ao4 i_130873703(.A(n_58396), .B(n_38911), .C(n_58472), .D(n_39882
		), .Z(n_1610));
	notech_reg to_acu0_reg_21(.CP(n_61881), .D(n_36950), .CD(n_61320), .Q(to_acu0
		[21]));
	notech_mux2 i_44247(.S(n_55031), .A(to_acu0[21]), .B(n_38561), .Z(n_36950
		));
	notech_ao4 i_130973702(.A(n_58394), .B(n_38913), .C(n_58472), .D(n_39883
		), .Z(n_1609));
	notech_reg to_acu0_reg_22(.CP(n_61881), .D(n_36956), .CD(n_61320), .Q(to_acu0
		[22]));
	notech_mux2 i_44255(.S(n_55031), .A(to_acu0[22]), .B(n_38563), .Z(n_36956
		));
	notech_ao4 i_131073701(.A(n_58391), .B(n_38915), .C(n_58472), .D(n_39884
		), .Z(n_1608));
	notech_reg to_acu0_reg_23(.CP(n_61881), .D(n_36962), .CD(n_61320), .Q(to_acu0
		[23]));
	notech_mux2 i_44263(.S(n_55031), .A(to_acu0[23]), .B(n_38565), .Z(n_36962
		));
	notech_ao4 i_131173700(.A(n_58391), .B(n_38917), .C(n_58470), .D(n_39885
		), .Z(n_1607));
	notech_reg to_acu0_reg_24(.CP(n_61881), .D(n_36968), .CD(n_61320), .Q(to_acu0
		[24]));
	notech_mux2 i_44271(.S(n_55031), .A(to_acu0[24]), .B(n_38567), .Z(n_36968
		));
	notech_ao4 i_131273699(.A(n_58391), .B(n_38919), .C(n_58470), .D(n_39886
		), .Z(n_1606));
	notech_reg to_acu0_reg_25(.CP(n_61881), .D(n_36974), .CD(n_61320), .Q(to_acu0
		[25]));
	notech_mux2 i_44279(.S(n_55031), .A(to_acu0[25]), .B(n_38569), .Z(n_36974
		));
	notech_ao4 i_134273669(.A(n_58391), .B(n_38979), .C(n_58472), .D(n_39916
		), .Z(n_1605));
	notech_reg to_acu0_reg_26(.CP(n_61881), .D(n_36980), .CD(n_61320), .Q(to_acu0
		[26]));
	notech_mux2 i_44287(.S(n_55031), .A(to_acu0[26]), .B(n_38571), .Z(n_36980
		));
	notech_ao4 i_134573666(.A(n_58391), .B(n_38985), .C(n_58472), .D(n_39919
		), .Z(n_1604));
	notech_reg to_acu0_reg_27(.CP(n_61879), .D(n_36986), .CD(n_61320), .Q(to_acu0
		[27]));
	notech_mux2 i_44295(.S(n_55026), .A(to_acu0[27]), .B(n_38573), .Z(n_36986
		));
	notech_ao4 i_136073651(.A(n_58391), .B(n_39015), .C(n_58467), .D(n_39934
		), .Z(n_1603));
	notech_reg to_acu0_reg_28(.CP(n_61879), .D(n_36992), .CD(n_61320), .Q(to_acu0
		[28]));
	notech_mux2 i_44303(.S(n_55031), .A(to_acu0[28]), .B(n_38575), .Z(n_36992
		));
	notech_reg to_acu0_reg_29(.CP(n_61879), .D(n_36998), .CD(n_61318), .Q(to_acu0
		[29]));
	notech_mux2 i_44311(.S(n_55026), .A(to_acu0[29]), .B(n_38577), .Z(n_36998
		));
	notech_ao4 i_137373638(.A(n_58467), .B(n_39944), .C(n_2056), .D(n_38627)
		, .Z(n_1601));
	notech_reg to_acu0_reg_30(.CP(n_61879), .D(n_37004), .CD(n_61318), .Q(to_acu0
		[30]));
	notech_mux2 i_44319(.S(n_55026), .A(to_acu0[30]), .B(n_38581), .Z(n_37004
		));
	notech_reg to_acu0_reg_31(.CP(n_61879), .D(n_37010), .CD(n_61318), .Q(to_acu0
		[31]));
	notech_mux2 i_44327(.S(n_55031), .A(to_acu0[31]), .B(n_38586), .Z(n_37010
		));
	notech_ao4 i_137573636(.A(n_58467), .B(n_39945), .C(n_2056), .D(n_38628)
		, .Z(n_1599));
	notech_reg to_acu0_reg_32(.CP(n_61881), .D(n_37016), .CD(n_61318), .Q(to_acu0
		[32]));
	notech_mux2 i_44335(.S(n_55031), .A(to_acu0[32]), .B(n_38589), .Z(n_37016
		));
	notech_reg to_acu0_reg_33(.CP(n_61881), .D(n_37022), .CD(n_61318), .Q(to_acu0
		[33]));
	notech_mux2 i_44343(.S(n_55031), .A(to_acu0[33]), .B(n_38591), .Z(n_37022
		));
	notech_ao4 i_137773634(.A(n_58467), .B(n_39946), .C(n_2056), .D(n_38630)
		, .Z(n_1597));
	notech_reg to_acu0_reg_34(.CP(n_61881), .D(n_37028), .CD(n_61320), .Q(to_acu0
		[34]));
	notech_mux2 i_44351(.S(n_55031), .A(to_acu0[34]), .B(n_38593), .Z(n_37028
		));
	notech_reg to_acu0_reg_35(.CP(n_61879), .D(n_37034), .CD(n_61320), .Q(to_acu0
		[35]));
	notech_mux2 i_44359(.S(n_55031), .A(to_acu0[35]), .B(n_38597), .Z(n_37034
		));
	notech_ao4 i_137973632(.A(n_58467), .B(n_39947), .C(n_2056), .D(n_38631)
		, .Z(n_1595));
	notech_reg to_acu0_reg_36(.CP(n_61881), .D(n_37040), .CD(n_61318), .Q(to_acu0
		[36]));
	notech_mux2 i_44367(.S(\nbus_13539[0] ), .A(to_acu0[36]), .B(n_38599), .Z
		(n_37040));
	notech_reg to_acu0_reg_37(.CP(n_61875), .D(n_37046), .CD(n_61318), .Q(to_acu0
		[37]));
	notech_mux2 i_44375(.S(\nbus_13539[0] ), .A(to_acu0[37]), .B(n_38601), .Z
		(n_37046));
	notech_ao4 i_138373628(.A(n_58467), .B(n_39949), .C(n_2056), .D(n_38634)
		, .Z(n_1593));
	notech_reg to_acu0_reg_38(.CP(n_61870), .D(n_37052), .CD(n_61318), .Q(to_acu0
		[38]));
	notech_mux2 i_44383(.S(\nbus_13539[0] ), .A(to_acu0[38]), .B(n_38603), .Z
		(n_37052));
	notech_ao4 i_138873623(.A(n_58391), .B(n_39047), .C(n_58467), .D(n_39954
		), .Z(n_1592));
	notech_reg to_acu0_reg_39(.CP(n_61870), .D(n_37058), .CD(n_61309), .Q(to_acu0
		[39]));
	notech_mux2 i_44391(.S(\nbus_13539[0] ), .A(to_acu0[39]), .B(n_43312), .Z
		(n_37058));
	notech_ao4 i_138973622(.A(n_58394), .B(n_39049), .C(n_58467), .D(n_39955
		), .Z(n_1591));
	notech_reg to_acu0_reg_40(.CP(n_61870), .D(n_37064), .CD(n_61309), .Q(to_acu0
		[40]));
	notech_mux2 i_44399(.S(\nbus_13539[0] ), .A(to_acu0[40]), .B(n_38604), .Z
		(n_37064));
	notech_ao4 i_139073621(.A(n_58394), .B(n_39051), .C(n_58470), .D(n_39956
		), .Z(n_1590));
	notech_reg to_acu0_reg_41(.CP(n_61870), .D(n_37070), .CD(n_61309), .Q(to_acu0
		[41]));
	notech_mux2 i_44407(.S(\nbus_13539[0] ), .A(to_acu0[41]), .B(n_38607), .Z
		(n_37070));
	notech_ao4 i_139273619(.A(n_58394), .B(n_39055), .C(n_58470), .D(n_39958
		), .Z(n_1589));
	notech_reg to_acu0_reg_42(.CP(n_61870), .D(n_37076), .CD(n_61309), .Q(to_acu0
		[42]));
	notech_mux2 i_44415(.S(\nbus_13539[0] ), .A(to_acu0[42]), .B(n_38608), .Z
		(n_37076));
	notech_ao4 i_139373618(.A(n_58394), .B(n_39057), .C(n_58470), .D(n_39959
		), .Z(n_1588));
	notech_reg to_acu0_reg_43(.CP(n_61873), .D(n_37082), .CD(n_61309), .Q(to_acu0
		[43]));
	notech_mux2 i_44423(.S(\nbus_13539[0] ), .A(to_acu0[43]), .B(n_38609), .Z
		(n_37082));
	notech_ao4 i_139573616(.A(n_58391), .B(n_39061), .C(n_58470), .D(n_39961
		), .Z(n_1587));
	notech_reg to_acu0_reg_44(.CP(n_61873), .D(n_37088), .CD(n_61312), .Q(to_acu0
		[44]));
	notech_mux2 i_44431(.S(\nbus_13539[0] ), .A(to_acu0[44]), .B(n_38610), .Z
		(n_37088));
	notech_reg to_acu0_reg_45(.CP(n_61873), .D(n_37094), .CD(n_61312), .Q(to_acu0
		[45]));
	notech_mux2 i_44439(.S(\nbus_13539[0] ), .A(to_acu0[45]), .B(n_38611), .Z
		(n_37094));
	notech_reg to_acu0_reg_46(.CP(n_61873), .D(n_37100), .CD(n_61312), .Q(to_acu0
		[46]));
	notech_mux2 i_44447(.S(n_55031), .A(to_acu0[46]), .B(n_38612), .Z(n_37100
		));
	notech_ao4 i_141273599(.A(n_58470), .B(n_39975), .C(n_2056), .D(n_161751607
		), .Z(n_1585));
	notech_reg to_acu0_reg_47(.CP(n_61873), .D(n_37106), .CD(n_61309), .Q(to_acu0
		[47]));
	notech_mux2 i_44455(.S(\nbus_13539[0] ), .A(to_acu0[47]), .B(n_38613), .Z
		(n_37106));
	notech_ao4 i_141373598(.A(n_58394), .B(n_39090), .C(n_58470), .D(n_39976
		), .Z(n_1584));
	notech_reg to_acu0_reg_48(.CP(n_61870), .D(n_37112), .CD(n_61309), .Q(to_acu0
		[48]));
	notech_mux2 i_44463(.S(\nbus_13539[0] ), .A(to_acu0[48]), .B(n_38614), .Z
		(n_37112));
	notech_ao4 i_141473597(.A(n_58394), .B(n_39092), .C(n_58470), .D(n_39977
		), .Z(n_1583));
	notech_reg to_acu0_reg_49(.CP(n_61870), .D(n_37118), .CD(n_61309), .Q(to_acu0
		[49]));
	notech_mux2 i_44471(.S(\nbus_13539[0] ), .A(to_acu0[49]), .B(n_38615), .Z
		(n_37118));
	notech_reg to_acu0_reg_50(.CP(n_61870), .D(n_37124), .CD(n_61309), .Q(to_acu0
		[50]));
	notech_mux2 i_44479(.S(\nbus_13539[0] ), .A(to_acu0[50]), .B(n_38616), .Z
		(n_37124));
	notech_reg to_acu0_reg_51(.CP(n_61870), .D(n_37130), .CD(n_61309), .Q(to_acu0
		[51]));
	notech_mux2 i_44487(.S(\nbus_13539[0] ), .A(to_acu0[51]), .B(n_38617), .Z
		(n_37130));
	notech_reg to_acu0_reg_52(.CP(n_61870), .D(n_37136), .CD(n_61309), .Q(to_acu0
		[52]));
	notech_mux2 i_44495(.S(n_55022), .A(to_acu0[52]), .B(n_38618), .Z(n_37136
		));
	notech_reg to_acu0_reg_53(.CP(n_61870), .D(n_37142), .CD(n_61309), .Q(to_acu0
		[53]));
	notech_mux2 i_44503(.S(n_55022), .A(to_acu0[53]), .B(n_38619), .Z(n_37142
		));
	notech_reg to_acu0_reg_54(.CP(n_61870), .D(n_37148), .CD(n_61309), .Q(to_acu0
		[54]));
	notech_mux2 i_44511(.S(n_55022), .A(to_acu0[54]), .B(n_38620), .Z(n_37148
		));
	notech_reg to_acu0_reg_55(.CP(n_61870), .D(n_37154), .CD(n_61309), .Q(to_acu0
		[55]));
	notech_mux2 i_44519(.S(n_55022), .A(to_acu0[55]), .B(n_38621), .Z(n_37154
		));
	notech_reg to_acu0_reg_56(.CP(n_61870), .D(n_37160), .CD(n_61309), .Q(to_acu0
		[56]));
	notech_mux2 i_44527(.S(n_55022), .A(to_acu0[56]), .B(n_38622), .Z(n_37160
		));
	notech_and4 i_143873573(.A(n_59686), .B(n_2126), .C(n_1574), .D(n_1563),
		 .Z(n_1577));
	notech_reg to_acu0_reg_57(.CP(n_61870), .D(n_37166), .CD(n_61309), .Q(to_acu0
		[57]));
	notech_mux2 i_44535(.S(n_55022), .A(to_acu0[57]), .B(n_38623), .Z(n_37166
		));
	notech_reg to_acu0_reg_58(.CP(n_61870), .D(n_37172), .CD(n_61309), .Q(to_acu0
		[58]));
	notech_mux2 i_44543(.S(n_55022), .A(to_acu0[58]), .B(n_38626), .Z(n_37172
		));
	notech_reg to_acu0_reg_59(.CP(n_61875), .D(n_37178), .CD(n_61309), .Q(to_acu0
		[59]));
	notech_mux2 i_44551(.S(n_55022), .A(to_acu0[59]), .B(n_38629), .Z(n_37178
		));
	notech_ao4 i_19474994(.A(n_2141), .B(n_39849), .C(n_38510), .D(n_39848),
		 .Z(n_1574));
	notech_reg to_acu0_reg_60(.CP(n_61875), .D(n_37184), .CD(n_61312), .Q(to_acu0
		[60]));
	notech_mux2 i_44559(.S(n_55017), .A(to_acu0[60]), .B(n_38632), .Z(n_37184
		));
	notech_reg to_acu0_reg_61(.CP(n_61875), .D(n_37191), .CD(n_61314), .Q(to_acu0
		[61]));
	notech_mux2 i_44567(.S(n_55017), .A(to_acu0[61]), .B(n_38635), .Z(n_37191
		));
	notech_and2 i_19174995(.A(n_40193), .B(n_59607), .Z(n_16150155));
	notech_reg to_acu0_reg_62(.CP(n_61873), .D(n_37197), .CD(n_61312), .Q(to_acu0
		[62]));
	notech_mux2 i_44575(.S(n_55017), .A(to_acu0[62]), .B(n_38636), .Z(n_37197
		));
	notech_ao4 i_144173570(.A(n_3247), .B(n_1480), .C(n_1479), .D(n_18050174
		), .Z(n_1572));
	notech_reg to_acu0_reg_63(.CP(n_61873), .D(n_37203), .CD(n_61312), .Q(to_acu0
		[63]));
	notech_mux2 i_44583(.S(n_55017), .A(to_acu0[63]), .B(n_38637), .Z(n_37203
		));
	notech_reg to_acu0_reg_64(.CP(n_61875), .D(n_37209), .CD(n_61312), .Q(to_acu0
		[64]));
	notech_mux2 i_44591(.S(n_55022), .A(to_acu0[64]), .B(n_38639), .Z(n_37209
		));
	notech_nand2 i_144373568(.A(n_2217), .B(n_2844), .Z(n_1570));
	notech_reg to_acu0_reg_65(.CP(n_61875), .D(n_37215), .CD(n_61314), .Q(to_acu0
		[65]));
	notech_mux2 i_44599(.S(n_55022), .A(to_acu0[65]), .B(n_38640), .Z(n_37215
		));
	notech_reg to_acu0_reg_66(.CP(n_61875), .D(n_37221), .CD(n_61314), .Q(to_acu0
		[66]));
	notech_mux2 i_44607(.S(n_55017), .A(to_acu0[66]), .B(n_38641), .Z(n_37221
		));
	notech_ao4 i_144573566(.A(pg_fault), .B(n_59607), .C(n_2833), .D(n_39848
		), .Z(n_1568));
	notech_reg to_acu0_reg_67(.CP(n_61875), .D(n_37227), .CD(n_61314), .Q(to_acu0
		[67]));
	notech_mux2 i_44615(.S(n_55017), .A(to_acu0[67]), .B(n_38642), .Z(n_37227
		));
	notech_or4 i_13674998(.A(n_58831), .B(pc_req), .C(pg_fault), .D(n_2138),
		 .Z(n_18050174));
	notech_reg to_acu0_reg_68(.CP(n_61875), .D(n_37233), .CD(n_61314), .Q(to_acu0
		[68]));
	notech_mux2 i_44623(.S(n_55022), .A(to_acu0[68]), .B(n_38341), .Z(n_37233
		));
	notech_and2 i_73618(.A(n_61314), .B(n_1411), .Z(\nbus_13559[0] ));
	notech_reg to_acu0_reg_69(.CP(n_61873), .D(n_37239), .CD(n_61312), .Q(to_acu0
		[69]));
	notech_mux2 i_44631(.S(n_55026), .A(to_acu0[69]), .B(n_38643), .Z(n_37239
		));
	notech_reg to_acu0_reg_70(.CP(n_61873), .D(n_37245), .CD(n_61312), .Q(to_acu0
		[70]));
	notech_mux2 i_44639(.S(n_55026), .A(to_acu0[70]), .B(n_38342), .Z(n_37245
		));
	notech_reg to_acu0_reg_71(.CP(n_61873), .D(n_37251), .CD(n_61312), .Q(to_acu0
		[71]));
	notech_mux2 i_44647(.S(n_55026), .A(to_acu0[71]), .B(n_38343), .Z(n_37251
		));
	notech_or2 i_122373788(.A(n_2056), .B(n_39849), .Z(n_1565));
	notech_reg to_acu0_reg_72(.CP(n_61873), .D(n_37257), .CD(n_61312), .Q(to_acu0
		[72]));
	notech_mux2 i_44655(.S(n_55026), .A(to_acu0[72]), .B(n_38344), .Z(n_37257
		));
	notech_reg to_acu0_reg_73(.CP(n_61873), .D(n_37263), .CD(n_61312), .Q(to_acu0
		[73]));
	notech_mux2 i_44663(.S(n_55026), .A(to_acu0[73]), .B(n_38345), .Z(n_37263
		));
	notech_or4 i_121773794(.A(n_56589), .B(pg_fault), .C(pc_req), .D(n_1476)
		, .Z(n_1563));
	notech_reg to_acu0_reg_74(.CP(n_61873), .D(n_37269), .CD(n_61312), .Q(to_acu0
		[74]));
	notech_mux2 i_44671(.S(n_55026), .A(to_acu0[74]), .B(n_38346), .Z(n_37269
		));
	notech_and3 i_2884(.A(n_39847), .B(n_1473), .C(n_2841), .Z(useq_ptr[1])
		);
	notech_reg to_acu0_reg_75(.CP(n_61873), .D(n_37275), .CD(n_61312), .Q(to_acu0
		[75]));
	notech_mux2 i_44679(.S(n_55026), .A(to_acu0[75]), .B(n_38347), .Z(n_37275
		));
	notech_reg to_acu0_reg_76(.CP(n_61873), .D(n_37281), .CD(n_61312), .Q(to_acu0
		[76]));
	notech_mux2 i_44687(.S(n_55026), .A(to_acu0[76]), .B(n_38348), .Z(n_37281
		));
	notech_reg to_acu0_reg_77(.CP(n_61873), .D(n_37287), .CD(n_61312), .Q(to_acu0
		[77]));
	notech_mux2 i_44695(.S(n_55022), .A(to_acu0[77]), .B(n_38349), .Z(n_37287
		));
	notech_reg to_acu0_reg_78(.CP(n_61873), .D(n_37293), .CD(n_61312), .Q(to_acu0
		[78]));
	notech_mux2 i_44703(.S(n_55022), .A(to_acu0[78]), .B(n_38350), .Z(n_37293
		));
	notech_reg to_acu0_reg_79(.CP(n_61873), .D(n_37299), .CD(n_61312), .Q(to_acu0
		[79]));
	notech_mux2 i_44711(.S(n_55022), .A(to_acu0[79]), .B(n_38351), .Z(n_37299
		));
	notech_reg to_acu0_reg_80(.CP(n_61840), .D(n_37305), .CD(n_61296), .Q(to_acu0
		[80]));
	notech_mux2 i_44719(.S(n_55022), .A(to_acu0[80]), .B(n_38352), .Z(n_37305
		));
	notech_reg to_acu0_reg_81(.CP(n_61840), .D(n_37311), .CD(n_61276), .Q(to_acu0
		[81]));
	notech_mux2 i_44727(.S(n_55026), .A(to_acu0[81]), .B(n_38353), .Z(n_37311
		));
	notech_nao3 i_26674743(.A(n_2847), .B(inst_deco1[113]), .C(n_1995), .Z(n_1556
		));
	notech_reg to_acu0_reg_82(.CP(n_61840), .D(n_37317), .CD(n_61279), .Q(to_acu0
		[82]));
	notech_mux2 i_44735(.S(n_55026), .A(to_acu0[82]), .B(n_38354), .Z(n_37317
		));
	notech_reg to_acu0_reg_83(.CP(n_61837), .D(n_37323), .CD(n_61276), .Q(to_acu0
		[83]));
	notech_mux2 i_44743(.S(n_55026), .A(to_acu0[83]), .B(n_38355), .Z(n_37323
		));
	notech_reg to_acu0_reg_84(.CP(n_61840), .D(n_37329), .CD(n_61276), .Q(to_acu0
		[84]));
	notech_mux2 i_44751(.S(n_55026), .A(to_acu0[84]), .B(n_38356), .Z(n_37329
		));
	notech_reg to_acu0_reg_85(.CP(n_61840), .D(n_37335), .CD(n_61276), .Q(to_acu0
		[85]));
	notech_mux2 i_44759(.S(n_54970), .A(to_acu0[85]), .B(n_38357), .Z(n_37335
		));
	notech_reg to_acu0_reg_86(.CP(n_61840), .D(n_37341), .CD(n_61279), .Q(to_acu0
		[86]));
	notech_mux2 i_44767(.S(n_54970), .A(to_acu0[86]), .B(n_38358), .Z(n_37341
		));
	notech_reg to_acu0_reg_87(.CP(n_61840), .D(n_37347), .CD(n_61279), .Q(to_acu0
		[87]));
	notech_mux2 i_44775(.S(n_54970), .A(to_acu0[87]), .B(n_38359), .Z(n_37347
		));
	notech_reg to_acu0_reg_88(.CP(n_61840), .D(n_37353), .CD(n_61279), .Q(to_acu0
		[88]));
	notech_mux2 i_44783(.S(n_54970), .A(to_acu0[88]), .B(n_38360), .Z(n_37353
		));
	notech_reg to_acu0_reg_89(.CP(n_61840), .D(n_37359), .CD(n_61279), .Q(to_acu0
		[89]));
	notech_mux2 i_44791(.S(n_54970), .A(to_acu0[89]), .B(n_38361), .Z(n_37359
		));
	notech_reg to_acu0_reg_90(.CP(n_61837), .D(n_37365), .CD(n_61279), .Q(to_acu0
		[90]));
	notech_mux2 i_44799(.S(n_54970), .A(to_acu0[90]), .B(n_38362), .Z(n_37365
		));
	notech_reg to_acu0_reg_91(.CP(n_61837), .D(n_37371), .CD(n_61276), .Q(to_acu0
		[91]));
	notech_mux2 i_44807(.S(n_54970), .A(to_acu0[91]), .B(n_38363), .Z(n_37371
		));
	notech_reg to_acu0_reg_92(.CP(n_61837), .D(n_37377), .CD(n_61276), .Q(to_acu0
		[92]));
	notech_mux2 i_44815(.S(n_54970), .A(to_acu0[92]), .B(n_38364), .Z(n_37377
		));
	notech_reg to_acu0_reg_93(.CP(n_61837), .D(n_37383), .CD(n_61276), .Q(to_acu0
		[93]));
	notech_mux2 i_44823(.S(n_54966), .A(to_acu0[93]), .B(n_38365), .Z(n_37383
		));
	notech_reg to_acu0_reg_94(.CP(n_61837), .D(n_37389), .CD(n_61276), .Q(to_acu0
		[94]));
	notech_mux2 i_44831(.S(n_54966), .A(to_acu0[94]), .B(n_38366), .Z(n_37389
		));
	notech_reg to_acu0_reg_95(.CP(n_61837), .D(n_37395), .CD(n_61276), .Q(to_acu0
		[95]));
	notech_mux2 i_44839(.S(n_54966), .A(to_acu0[95]), .B(n_38367), .Z(n_37395
		));
	notech_reg to_acu0_reg_96(.CP(n_61837), .D(n_37401), .CD(n_61276), .Q(to_acu0
		[96]));
	notech_mux2 i_44847(.S(n_54966), .A(to_acu0[96]), .B(n_38368), .Z(n_37401
		));
	notech_nao3 i_20774797(.A(n_2847), .B(inst_deco1[87]), .C(n_1995), .Z(n_1541
		));
	notech_reg to_acu0_reg_97(.CP(n_61837), .D(n_37407), .CD(n_61276), .Q(to_acu0
		[97]));
	notech_mux2 i_44855(.S(n_54966), .A(to_acu0[97]), .B(n_38369), .Z(n_37407
		));
	notech_reg to_acu0_reg_98(.CP(n_61837), .D(n_37413), .CD(n_61276), .Q(to_acu0
		[98]));
	notech_mux2 i_44863(.S(n_54966), .A(to_acu0[98]), .B(n_38370), .Z(n_37413
		));
	notech_reg to_acu0_reg_99(.CP(n_61837), .D(n_37419), .CD(n_61276), .Q(to_acu0
		[99]));
	notech_mux2 i_44871(.S(n_54966), .A(to_acu0[99]), .B(n_38371), .Z(n_37419
		));
	notech_nao3 i_19974803(.A(n_2847), .B(inst_deco1[85]), .C(n_1995), .Z(n_1538
		));
	notech_reg to_acu0_reg_100(.CP(n_61837), .D(n_37425), .CD(n_61276), .Q(to_acu0
		[100]));
	notech_mux2 i_44879(.S(n_54966), .A(to_acu0[100]), .B(n_38372), .Z(n_37425
		));
	notech_reg to_acu0_reg_101(.CP(n_61842), .D(n_37431), .CD(n_61276), .Q(to_acu0
		[101]));
	notech_mux2 i_44887(.S(n_54970), .A(to_acu0[101]), .B(n_38373), .Z(n_37431
		));
	notech_reg to_acu0_reg_102(.CP(n_61842), .D(n_37437), .CD(n_61281), .Q(to_acu0
		[102]));
	notech_mux2 i_44895(.S(n_54975), .A(to_acu0[102]), .B(n_38374), .Z(n_37437
		));
	notech_nao3 i_19674806(.A(n_2847), .B(inst_deco1[84]), .C(n_1995), .Z(n_1535
		));
	notech_reg to_acu0_reg_103(.CP(n_61842), .D(n_37443), .CD(n_61281), .Q(to_acu0
		[103]));
	notech_mux2 i_44903(.S(n_54975), .A(to_acu0[103]), .B(n_38375), .Z(n_37443
		));
	notech_reg to_acu0_reg_104(.CP(n_61842), .D(n_37449), .CD(n_61281), .Q(to_acu0
		[104]));
	notech_mux2 i_44911(.S(n_54975), .A(to_acu0[104]), .B(n_38376), .Z(n_37449
		));
	notech_reg to_acu0_reg_105(.CP(n_61842), .D(n_37455), .CD(n_61279), .Q(to_acu0
		[105]));
	notech_mux2 i_44919(.S(n_54975), .A(to_acu0[105]), .B(n_38377), .Z(n_37455
		));
	notech_nao3 i_19274809(.A(n_2847), .B(inst_deco1[83]), .C(n_1995), .Z(n_1532
		));
	notech_reg to_acu0_reg_106(.CP(n_61842), .D(n_37461), .CD(n_61281), .Q(to_acu0
		[106]));
	notech_mux2 i_44927(.S(n_54975), .A(to_acu0[106]), .B(n_38378), .Z(n_37461
		));
	notech_reg to_acu0_reg_107(.CP(n_61842), .D(n_37467), .CD(n_61281), .Q(to_acu0
		[107]));
	notech_mux2 i_44935(.S(n_54975), .A(to_acu0[107]), .B(n_38379), .Z(n_37467
		));
	notech_reg to_acu0_reg_108(.CP(n_61842), .D(n_37473), .CD(n_61281), .Q(to_acu0
		[108]));
	notech_mux2 i_44943(.S(n_54975), .A(to_acu0[108]), .B(n_38380), .Z(n_37473
		));
	notech_nao3 i_18874812(.A(n_2847), .B(inst_deco1[82]), .C(n_1995), .Z(n_1529
		));
	notech_reg to_acu0_reg_109(.CP(n_61842), .D(n_37479), .CD(n_61281), .Q(to_acu0
		[109]));
	notech_mux2 i_44951(.S(n_54975), .A(to_acu0[109]), .B(n_38381), .Z(n_37479
		));
	notech_reg to_acu0_reg_110(.CP(n_61842), .D(n_37485), .CD(n_61281), .Q(to_acu0
		[110]));
	notech_mux2 i_44959(.S(n_54970), .A(to_acu0[110]), .B(n_38382), .Z(n_37485
		));
	notech_reg to_acu0_reg_111(.CP(n_61842), .D(n_37491), .CD(n_61281), .Q(to_acu0
		[111]));
	notech_mux2 i_44967(.S(n_54970), .A(to_acu0[111]), .B(n_38383), .Z(n_37491
		));
	notech_reg to_acu0_reg_112(.CP(n_61840), .D(n_37497), .CD(n_61279), .Q(to_acu0
		[112]));
	notech_mux2 i_44975(.S(n_54970), .A(to_acu0[112]), .B(n_38644), .Z(n_37497
		));
	notech_reg to_acu0_reg_113(.CP(n_61840), .D(n_37503), .CD(n_61279), .Q(to_acu0
		[113]));
	notech_mux2 i_44983(.S(n_54970), .A(to_acu0[113]), .B(n_38384), .Z(n_37503
		));
	notech_reg to_acu0_reg_114(.CP(n_61840), .D(n_37509), .CD(n_61279), .Q(to_acu0
		[114]));
	notech_mux2 i_44991(.S(n_54975), .A(to_acu0[114]), .B(n_38385), .Z(n_37509
		));
	notech_reg to_acu0_reg_115(.CP(n_61840), .D(n_37515), .CD(n_61279), .Q(to_acu0
		[115]));
	notech_mux2 i_44999(.S(n_54975), .A(to_acu0[115]), .B(n_38386), .Z(n_37515
		));
	notech_reg to_acu0_reg_116(.CP(n_61840), .D(n_37521), .CD(n_61279), .Q(to_acu0
		[116]));
	notech_mux2 i_45007(.S(n_54970), .A(to_acu0[116]), .B(n_38387), .Z(n_37521
		));
	notech_reg to_acu0_reg_117(.CP(n_61840), .D(n_37527), .CD(n_61279), .Q(to_acu0
		[117]));
	notech_mux2 i_45015(.S(n_54970), .A(to_acu0[117]), .B(n_38645), .Z(n_37527
		));
	notech_reg to_acu0_reg_118(.CP(n_61842), .D(n_37533), .CD(n_61279), .Q(to_acu0
		[118]));
	notech_mux2 i_45023(.S(n_54957), .A(to_acu0[118]), .B(n_38388), .Z(n_37533
		));
	notech_reg to_acu0_reg_119(.CP(n_61840), .D(n_37539), .CD(n_61279), .Q(to_acu0
		[119]));
	notech_mux2 i_45031(.S(n_54957), .A(to_acu0[119]), .B(n_38646), .Z(n_37539
		));
	notech_reg to_acu0_reg_120(.CP(n_61840), .D(n_37545), .CD(n_61279), .Q(to_acu0
		[120]));
	notech_mux2 i_45039(.S(n_54957), .A(to_acu0[120]), .B(n_38389), .Z(n_37545
		));
	notech_reg to_acu0_reg_121(.CP(n_61840), .D(n_37551), .CD(n_61279), .Q(to_acu0
		[121]));
	notech_mux2 i_45047(.S(n_54957), .A(to_acu0[121]), .B(n_38390), .Z(n_37551
		));
	notech_reg to_acu0_reg_122(.CP(n_61837), .D(n_37557), .CD(n_61279), .Q(to_acu0
		[122]));
	notech_mux2 i_45055(.S(n_54961), .A(to_acu0[122]), .B(n_38391), .Z(n_37557
		));
	notech_reg to_acu0_reg_123(.CP(n_61832), .D(n_37563), .CD(n_61271), .Q(to_acu0
		[123]));
	notech_mux2 i_45063(.S(n_54961), .A(to_acu0[123]), .B(n_38648), .Z(n_37563
		));
	notech_reg to_acu0_reg_124(.CP(n_61832), .D(n_37569), .CD(n_61271), .Q(to_acu0
		[124]));
	notech_mux2 i_45071(.S(n_54961), .A(to_acu0[124]), .B(n_38650), .Z(n_37569
		));
	notech_reg to_acu0_reg_125(.CP(n_61832), .D(n_37575), .CD(n_61271), .Q(to_acu0
		[125]));
	notech_mux2 i_45079(.S(n_54961), .A(to_acu0[125]), .B(n_38392), .Z(n_37575
		));
	notech_reg to_acu0_reg_126(.CP(n_61832), .D(n_37581), .CD(n_61271), .Q(to_acu0
		[126]));
	notech_mux2 i_45087(.S(n_54957), .A(to_acu0[126]), .B(n_38651), .Z(n_37581
		));
	notech_reg to_acu0_reg_127(.CP(n_61832), .D(n_37587), .CD(n_61271), .Q(to_acu0
		[127]));
	notech_mux2 i_45095(.S(n_54957), .A(to_acu0[127]), .B(n_38652), .Z(n_37587
		));
	notech_reg to_acu0_reg_128(.CP(n_61835), .D(n_37593), .CD(n_61271), .Q(to_acu0
		[128]));
	notech_mux2 i_45103(.S(n_54957), .A(to_acu0[128]), .B(n_38654), .Z(n_37593
		));
	notech_reg to_acu0_reg_129(.CP(n_61835), .D(n_37599), .CD(n_61271), .Q(to_acu0
		[129]));
	notech_mux2 i_45111(.S(n_54957), .A(to_acu0[129]), .B(n_38393), .Z(n_37599
		));
	notech_reg to_acu0_reg_130(.CP(n_61832), .D(n_37605), .CD(n_61271), .Q(to_acu0
		[130]));
	notech_mux2 i_45119(.S(n_54957), .A(to_acu0[130]), .B(n_38655), .Z(n_37605
		));
	notech_reg to_acu0_reg_131(.CP(n_61832), .D(n_37611), .CD(n_61271), .Q(to_acu0
		[131]));
	notech_mux2 i_45127(.S(n_54957), .A(to_acu0[131]), .B(n_38657), .Z(n_37611
		));
	notech_reg to_acu0_reg_132(.CP(n_61832), .D(n_37617), .CD(n_61271), .Q(to_acu0
		[132]));
	notech_mux2 i_45135(.S(n_54957), .A(to_acu0[132]), .B(n_38658), .Z(n_37617
		));
	notech_reg to_acu0_reg_133(.CP(n_61832), .D(n_37623), .CD(n_61271), .Q(to_acu0
		[133]));
	notech_mux2 i_45143(.S(n_54957), .A(to_acu0[133]), .B(n_38660), .Z(n_37623
		));
	notech_reg to_acu0_reg_134(.CP(n_61832), .D(n_37629), .CD(n_61271), .Q(to_acu0
		[134]));
	notech_mux2 i_45151(.S(n_54961), .A(to_acu0[134]), .B(n_38662), .Z(n_37629
		));
	notech_reg to_acu0_reg_135(.CP(n_61832), .D(n_37635), .CD(n_61271), .Q(to_acu0
		[135]));
	notech_mux2 i_45159(.S(n_54966), .A(to_acu0[135]), .B(n_38663), .Z(n_37635
		));
	notech_reg to_acu0_reg_136(.CP(n_61832), .D(n_37641), .CD(n_61269), .Q(to_acu0
		[136]));
	notech_mux2 i_45167(.S(n_54966), .A(to_acu0[136]), .B(n_38665), .Z(n_37641
		));
	notech_reg to_acu0_reg_137(.CP(n_61830), .D(n_37647), .CD(n_61269), .Q(to_acu0
		[137]));
	notech_mux2 i_45175(.S(n_54961), .A(to_acu0[137]), .B(n_38394), .Z(n_37647
		));
	notech_reg to_acu0_reg_138(.CP(n_61832), .D(n_37653), .CD(n_61269), .Q(to_acu0
		[138]));
	notech_mux2 i_45183(.S(n_54966), .A(to_acu0[138]), .B(n_39854), .Z(n_37653
		));
	notech_reg to_acu0_reg_139(.CP(n_61832), .D(n_37659), .CD(n_61271), .Q(to_acu0
		[139]));
	notech_mux2 i_45191(.S(n_54966), .A(to_acu0[139]), .B(n_38667), .Z(n_37659
		));
	notech_reg to_acu0_reg_140(.CP(n_61832), .D(n_37665), .CD(n_61271), .Q(to_acu0
		[140]));
	notech_mux2 i_45199(.S(n_54966), .A(to_acu0[140]), .B(n_38670), .Z(n_37665
		));
	notech_reg to_acu0_reg_141(.CP(n_61832), .D(n_37671), .CD(n_61271), .Q(to_acu0
		[141]));
	notech_mux2 i_45207(.S(n_54966), .A(to_acu0[141]), .B(n_38673), .Z(n_37671
		));
	notech_reg to_acu0_reg_142(.CP(n_61832), .D(n_37677), .CD(n_61271), .Q(to_acu0
		[142]));
	notech_mux2 i_45215(.S(n_54966), .A(to_acu0[142]), .B(n_38675), .Z(n_37677
		));
	notech_reg to_acu0_reg_143(.CP(n_61832), .D(n_37683), .CD(n_61271), .Q(to_acu0
		[143]));
	notech_mux2 i_45223(.S(n_54961), .A(to_acu0[143]), .B(n_38677), .Z(n_37683
		));
	notech_reg to_acu0_reg_144(.CP(n_61835), .D(n_37689), .CD(n_61274), .Q(to_acu0
		[144]));
	notech_mux2 i_45231(.S(n_54961), .A(to_acu0[144]), .B(n_38679), .Z(n_37689
		));
	notech_reg to_acu0_reg_145(.CP(n_61835), .D(n_37695), .CD(n_61274), .Q(to_acu0
		[145]));
	notech_mux2 i_45239(.S(n_54961), .A(to_acu0[145]), .B(n_38682), .Z(n_37695
		));
	notech_reg to_acu0_reg_146(.CP(n_61835), .D(n_37701), .CD(n_61274), .Q(to_acu0
		[146]));
	notech_mux2 i_45247(.S(n_54961), .A(to_acu0[146]), .B(n_39855), .Z(n_37701
		));
	notech_reg to_acu0_reg_147(.CP(n_61835), .D(n_37707), .CD(n_61274), .Q(to_acu0
		[147]));
	notech_mux2 i_45255(.S(n_54961), .A(to_acu0[147]), .B(n_38685), .Z(n_37707
		));
	notech_and3 i_2940(.A(n_2124), .B(lenpc2[31]), .C(n_59607), .Z(n_44548)
		);
	notech_reg to_acu0_reg_148(.CP(n_61835), .D(n_37713), .CD(n_61274), .Q(to_acu0
		[148]));
	notech_mux2 i_45263(.S(n_54961), .A(to_acu0[148]), .B(n_38688), .Z(n_37713
		));
	notech_and3 i_2939(.A(n_2124), .B(lenpc2[30]), .C(n_59607), .Z(n_44542)
		);
	notech_reg to_acu0_reg_149(.CP(n_61837), .D(n_37719), .CD(n_61276), .Q(to_acu0
		[149]));
	notech_mux2 i_45271(.S(n_54961), .A(to_acu0[149]), .B(n_38691), .Z(n_37719
		));
	notech_and3 i_2938(.A(n_2124), .B(lenpc2[29]), .C(n_59607), .Z(n_44536)
		);
	notech_reg to_acu0_reg_150(.CP(n_61837), .D(n_37725), .CD(n_61276), .Q(to_acu0
		[150]));
	notech_mux2 i_45279(.S(n_54961), .A(to_acu0[150]), .B(n_38694), .Z(n_37725
		));
	notech_and3 i_2937(.A(n_2124), .B(lenpc2[28]), .C(n_59607), .Z(n_44530)
		);
	notech_reg to_acu0_reg_151(.CP(n_61837), .D(n_37731), .CD(n_61276), .Q(to_acu0
		[151]));
	notech_mux2 i_45287(.S(n_54975), .A(to_acu0[151]), .B(n_38697), .Z(n_37731
		));
	notech_and3 i_2936(.A(n_2124), .B(lenpc2[27]), .C(n_59607), .Z(n_44524)
		);
	notech_reg to_acu0_reg_152(.CP(n_61837), .D(n_37737), .CD(n_61274), .Q(to_acu0
		[152]));
	notech_mux2 i_45295(.S(n_54989), .A(to_acu0[152]), .B(n_38700), .Z(n_37737
		));
	notech_and3 i_2929(.A(n_59669), .B(lenpc2[20]), .C(n_59607), .Z(n_44482)
		);
	notech_reg to_acu0_reg_153(.CP(n_61837), .D(n_37743), .CD(n_61274), .Q(to_acu0
		[153]));
	notech_mux2 i_45303(.S(n_54989), .A(to_acu0[153]), .B(n_38703), .Z(n_37743
		));
	notech_and3 i_2928(.A(n_59669), .B(lenpc2[19]), .C(n_59607), .Z(n_44476)
		);
	notech_reg to_acu0_reg_154(.CP(n_61835), .D(n_37749), .CD(n_61274), .Q(to_acu0
		[154]));
	notech_mux2 i_45311(.S(n_54989), .A(to_acu0[154]), .B(n_38706), .Z(n_37749
		));
	notech_and3 i_2927(.A(n_59669), .B(lenpc2[18]), .C(n_59607), .Z(n_44470)
		);
	notech_reg to_acu0_reg_155(.CP(n_61835), .D(n_37755), .CD(n_61274), .Q(to_acu0
		[155]));
	notech_mux2 i_45319(.S(n_54989), .A(to_acu0[155]), .B(n_38709), .Z(n_37755
		));
	notech_and3 i_2926(.A(n_59669), .B(lenpc2[17]), .C(n_59607), .Z(n_44464)
		);
	notech_reg to_acu0_reg_156(.CP(n_61835), .D(n_37761), .CD(n_61274), .Q(to_acu0
		[156]));
	notech_mux2 i_45327(.S(n_54989), .A(to_acu0[156]), .B(n_38712), .Z(n_37761
		));
	notech_and3 i_2925(.A(n_59669), .B(lenpc2[16]), .C(n_59602), .Z(n_44458)
		);
	notech_reg to_acu0_reg_157(.CP(n_61835), .D(n_37767), .CD(n_61274), .Q(to_acu0
		[157]));
	notech_mux2 i_45335(.S(n_54989), .A(to_acu0[157]), .B(n_38715), .Z(n_37767
		));
	notech_and3 i_2924(.A(n_59669), .B(lenpc2[15]), .C(n_59602), .Z(n_44452)
		);
	notech_reg to_acu0_reg_158(.CP(n_61835), .D(n_37773), .CD(n_61274), .Q(to_acu0
		[158]));
	notech_mux2 i_45343(.S(n_54989), .A(to_acu0[158]), .B(n_38718), .Z(n_37773
		));
	notech_and3 i_2923(.A(n_59669), .B(lenpc2[14]), .C(n_59602), .Z(n_44446)
		);
	notech_reg to_acu0_reg_159(.CP(n_61835), .D(n_37779), .CD(n_61274), .Q(to_acu0
		[159]));
	notech_mux2 i_45351(.S(n_54989), .A(to_acu0[159]), .B(n_38721), .Z(n_37779
		));
	notech_and3 i_2922(.A(n_59669), .B(lenpc2[13]), .C(n_59602), .Z(n_44440)
		);
	notech_reg to_acu0_reg_160(.CP(n_61835), .D(n_37785), .CD(n_61274), .Q(to_acu0
		[160]));
	notech_mux2 i_45359(.S(n_54989), .A(to_acu0[160]), .B(n_38724), .Z(n_37785
		));
	notech_and3 i_2921(.A(n_59669), .B(lenpc2[12]), .C(n_59602), .Z(n_44434)
		);
	notech_reg to_acu0_reg_161(.CP(n_61835), .D(n_37791), .CD(n_61274), .Q(to_acu0
		[161]));
	notech_mux2 i_45367(.S(n_54989), .A(to_acu0[161]), .B(n_38727), .Z(n_37791
		));
	notech_and3 i_2920(.A(n_59669), .B(lenpc2[11]), .C(n_59602), .Z(n_44428)
		);
	notech_reg to_acu0_reg_162(.CP(n_61835), .D(n_37797), .CD(n_61274), .Q(to_acu0
		[162]));
	notech_mux2 i_45375(.S(n_54985), .A(to_acu0[162]), .B(n_38730), .Z(n_37797
		));
	notech_and3 i_2919(.A(n_59669), .B(lenpc2[10]), .C(n_59607), .Z(n_44422)
		);
	notech_reg to_acu0_reg_163(.CP(n_61835), .D(n_37803), .CD(n_61274), .Q(to_acu0
		[163]));
	notech_mux2 i_45383(.S(n_54989), .A(to_acu0[163]), .B(n_38733), .Z(n_37803
		));
	notech_and3 i_2918(.A(n_59669), .B(lenpc2[9]), .C(n_59607), .Z(n_44416)
		);
	notech_reg to_acu0_reg_164(.CP(n_61835), .D(n_37809), .CD(n_61274), .Q(to_acu0
		[164]));
	notech_mux2 i_45391(.S(n_54989), .A(to_acu0[164]), .B(n_38736), .Z(n_37809
		));
	notech_and3 i_2917(.A(n_59669), .B(lenpc2[8]), .C(n_59607), .Z(n_44410)
		);
	notech_reg to_acu0_reg_165(.CP(n_61852), .D(n_37815), .CD(n_61281), .Q(to_acu0
		[165]));
	notech_mux2 i_45399(.S(n_54989), .A(to_acu0[165]), .B(n_38739), .Z(n_37815
		));
	notech_and3 i_2916(.A(n_59669), .B(lenpc2[7]), .C(n_59602), .Z(n_44404)
		);
	notech_reg to_acu0_reg_166(.CP(n_61852), .D(n_37821), .CD(n_61291), .Q(to_acu0
		[166]));
	notech_mux2 i_45407(.S(n_54989), .A(to_acu0[166]), .B(n_38742), .Z(n_37821
		));
	notech_and3 i_2915(.A(n_59669), .B(lenpc2[6]), .C(n_59602), .Z(n_44398)
		);
	notech_reg to_acu0_reg_167(.CP(n_61852), .D(n_37827), .CD(n_61291), .Q(to_acu0
		[167]));
	notech_mux2 i_45415(.S(n_54989), .A(to_acu0[167]), .B(n_38745), .Z(n_37827
		));
	notech_and3 i_2914(.A(to_acu1[39]), .B(n_59669), .C(n_59602), .Z(n_43312
		));
	notech_reg to_acu0_reg_168(.CP(n_61852), .D(n_37833), .CD(n_61291), .Q(to_acu0
		[168]));
	notech_mux2 i_45423(.S(n_54994), .A(to_acu0[168]), .B(n_38748), .Z(n_37833
		));
	notech_and4 i_123373778(.A(n_5761), .B(n_1740), .C(n_2120), .D(\to_acu2_0[69] 
		), .Z(n_1490));
	notech_reg to_acu0_reg_169(.CP(n_61852), .D(n_37839), .CD(n_61291), .Q(to_acu0
		[169]));
	notech_mux2 i_45431(.S(n_54994), .A(to_acu0[169]), .B(n_39856), .Z(n_37839
		));
	notech_or2 i_123273779(.A(n_2798), .B(n_251191358), .Z(n_1489));
	notech_reg to_acu0_reg_170(.CP(n_61854), .D(n_37845), .CD(n_61291), .Q(to_acu0
		[170]));
	notech_mux2 i_45439(.S(n_54994), .A(to_acu0[170]), .B(n_38751), .Z(n_37845
		));
	notech_reg to_acu0_reg_171(.CP(n_61854), .D(n_37851), .CD(n_61291), .Q(to_acu0
		[171]));
	notech_mux2 i_45447(.S(n_54994), .A(to_acu0[171]), .B(n_38754), .Z(n_37851
		));
	notech_reg to_acu0_reg_172(.CP(n_61854), .D(n_37857), .CD(n_61293), .Q(to_acu0
		[172]));
	notech_mux2 i_45455(.S(n_54994), .A(to_acu0[172]), .B(n_38757), .Z(n_37857
		));
	notech_ao4 i_174989(.A(n_38425), .B(n_39570), .C(n_2958), .D(n_2798), .Z
		(n_1486));
	notech_reg to_acu0_reg_173(.CP(n_61852), .D(n_37863), .CD(n_61291), .Q(to_acu0
		[173]));
	notech_mux2 i_45463(.S(n_54998), .A(to_acu0[173]), .B(n_38760), .Z(n_37863
		));
	notech_nand2 i_122973782(.A(db67), .B(n_40106), .Z(n_1485));
	notech_reg to_acu0_reg_174(.CP(n_61854), .D(n_37869), .CD(n_61291), .Q(to_acu0
		[174]));
	notech_mux2 i_45471(.S(n_54998), .A(to_acu0[174]), .B(n_38763), .Z(n_37869
		));
	notech_nand2 i_122873783(.A(n_2120), .B(n_2125), .Z(n_1484));
	notech_reg to_acu0_reg_175(.CP(n_61852), .D(n_37875), .CD(n_61291), .Q(to_acu0
		[175]));
	notech_mux2 i_45479(.S(n_54994), .A(to_acu0[175]), .B(n_38766), .Z(n_37875
		));
	notech_and4 i_122773784(.A(n_2120), .B(n_1740), .C(n_2121), .D(n_2122), 
		.Z(n_1483));
	notech_reg to_acu0_reg_176(.CP(n_61852), .D(n_37881), .CD(n_61291), .Q(to_acu0
		[176]));
	notech_mux2 i_45487(.S(n_54994), .A(to_acu0[176]), .B(n_38769), .Z(n_37881
		));
	notech_reg to_acu0_reg_177(.CP(n_61852), .D(n_37887), .CD(n_61291), .Q(to_acu0
		[177]));
	notech_mux2 i_45495(.S(n_54994), .A(to_acu0[177]), .B(n_38772), .Z(n_37887
		));
	notech_ao4 i_122573786(.A(n_2834), .B(n_38661), .C(n_2833), .D(n_1570), 
		.Z(n_1481));
	notech_reg to_acu0_reg_178(.CP(n_61852), .D(n_37893), .CD(n_61291), .Q(to_acu0
		[178]));
	notech_mux2 i_45503(.S(n_54994), .A(to_acu0[178]), .B(n_38775), .Z(n_37893
		));
	notech_nor2 i_374987(.A(idx_deco[1]), .B(idx_deco[0]), .Z(n_1480));
	notech_reg to_acu0_reg_179(.CP(n_61852), .D(n_37899), .CD(n_61291), .Q(to_acu0
		[179]));
	notech_mux2 i_45511(.S(n_54994), .A(to_acu0[179]), .B(n_38778), .Z(n_37899
		));
	notech_and2 i_274988(.A(n_1994), .B(n_38329), .Z(n_1479));
	notech_reg to_acu0_reg_180(.CP(n_61852), .D(n_37905), .CD(n_61288), .Q(to_acu0
		[180]));
	notech_mux2 i_45519(.S(n_54994), .A(to_acu0[180]), .B(n_38781), .Z(n_37905
		));
	notech_reg to_acu0_reg_181(.CP(n_61852), .D(n_37911), .CD(n_61288), .Q(to_acu0
		[181]));
	notech_mux2 i_45527(.S(n_54994), .A(to_acu0[181]), .B(n_38784), .Z(n_37911
		));
	notech_reg to_acu0_reg_182(.CP(n_61852), .D(n_37917), .CD(n_61291), .Q(to_acu0
		[182]));
	notech_mux2 i_45535(.S(n_54994), .A(to_acu0[182]), .B(n_38787), .Z(n_37917
		));
	notech_ao3 i_474986(.A(n_2071), .B(n_39849), .C(ipg_fault), .Z(n_1476)
		);
	notech_reg to_acu0_reg_183(.CP(n_61852), .D(n_37923), .CD(n_61291), .Q(to_acu0
		[183]));
	notech_mux2 i_45543(.S(n_54994), .A(to_acu0[183]), .B(n_38790), .Z(n_37923
		));
	notech_and4 i_121673795(.A(n_17550169), .B(n_40176), .C(in128[0]), .D(\to_acu2_0[9] 
		), .Z(n_1475));
	notech_reg to_acu0_reg_184(.CP(n_61852), .D(n_37929), .CD(n_61291), .Q(to_acu0
		[184]));
	notech_mux2 i_45551(.S(n_54994), .A(to_acu0[184]), .B(n_38793), .Z(n_37929
		));
	notech_or4 i_121573796(.A(idx_deco[1]), .B(n_58470), .C(idx_deco[0]), .D
		(n_2138), .Z(n_1474));
	notech_reg to_acu0_reg_185(.CP(n_61852), .D(n_37935), .CD(n_61291), .Q(to_acu0
		[185]));
	notech_mux2 i_45559(.S(n_54955), .A(to_acu0[185]), .B(n_38796), .Z(n_37935
		));
	notech_or4 i_35674653(.A(i_ptr[1]), .B(i_ptr[0]), .C(i_ptr[3]), .D(i_ptr
		[2]), .Z(n_1473));
	notech_reg to_acu0_reg_186(.CP(n_61857), .D(n_37941), .CD(n_61291), .Q(to_acu0
		[186]));
	notech_mux2 i_45567(.S(n_54955), .A(to_acu0[186]), .B(n_38799), .Z(n_37941
		));
	notech_reg to_acu0_reg_187(.CP(n_61857), .D(n_37947), .CD(n_61293), .Q(to_acu0
		[187]));
	notech_mux2 i_45575(.S(n_54955), .A(to_acu0[187]), .B(n_38802), .Z(n_37947
		));
	notech_reg to_acu0_reg_188(.CP(n_61854), .D(n_37953), .CD(n_61293), .Q(to_acu0
		[188]));
	notech_mux2 i_45583(.S(n_54955), .A(to_acu0[188]), .B(n_38805), .Z(n_37953
		));
	notech_reg to_acu0_reg_189(.CP(n_61854), .D(n_37959), .CD(n_61293), .Q(to_acu0
		[189]));
	notech_mux2 i_45591(.S(n_54955), .A(to_acu0[189]), .B(n_38808), .Z(n_37959
		));
	notech_reg to_acu0_reg_190(.CP(n_61854), .D(n_37965), .CD(n_61293), .Q(to_acu0
		[190]));
	notech_mux2 i_45599(.S(n_54955), .A(to_acu0[190]), .B(n_38811), .Z(n_37965
		));
	notech_reg to_acu0_reg_191(.CP(n_61857), .D(n_37971), .CD(n_61293), .Q(to_acu0
		[191]));
	notech_mux2 i_45607(.S(n_54955), .A(to_acu0[191]), .B(n_38814), .Z(n_37971
		));
	notech_reg to_acu0_reg_192(.CP(n_61857), .D(n_37977), .CD(n_61296), .Q(to_acu0
		[192]));
	notech_mux2 i_45615(.S(n_54955), .A(to_acu0[192]), .B(n_38817), .Z(n_37977
		));
	notech_reg to_acu0_reg_193(.CP(n_61857), .D(n_37983), .CD(n_61296), .Q(to_acu0
		[193]));
	notech_mux2 i_45623(.S(n_54975), .A(to_acu0[193]), .B(n_38820), .Z(n_37983
		));
	notech_reg to_acu0_reg_194(.CP(n_61857), .D(n_37989), .CD(n_61296), .Q(to_acu0
		[194]));
	notech_mux2 i_45631(.S(n_54975), .A(to_acu0[194]), .B(n_38823), .Z(n_37989
		));
	notech_reg to_acu0_reg_195(.CP(n_61857), .D(n_37995), .CD(n_61293), .Q(to_acu0
		[195]));
	notech_mux2 i_45639(.S(n_54975), .A(to_acu0[195]), .B(n_38826), .Z(n_37995
		));
	notech_reg to_acu0_reg_196(.CP(n_61854), .D(n_38001), .CD(n_61296), .Q(to_acu0
		[196]));
	notech_mux2 i_45647(.S(n_54975), .A(to_acu0[196]), .B(n_38829), .Z(n_38001
		));
	notech_reg to_acu0_reg_197(.CP(n_61854), .D(n_38007), .CD(n_61293), .Q(to_acu0
		[197]));
	notech_mux2 i_45655(.S(n_54955), .A(to_acu0[197]), .B(n_38832), .Z(n_38007
		));
	notech_reg to_acu0_reg_198(.CP(n_61854), .D(n_38013), .CD(n_61293), .Q(to_acu0
		[198]));
	notech_mux2 i_45663(.S(n_54955), .A(to_acu0[198]), .B(n_38836), .Z(n_38013
		));
	notech_reg to_acu0_reg_199(.CP(n_61854), .D(n_38019), .CD(n_61293), .Q(to_acu0
		[199]));
	notech_mux2 i_45671(.S(n_54955), .A(to_acu0[199]), .B(n_38839), .Z(n_38019
		));
	notech_reg to_acu0_reg_200(.CP(n_61854), .D(n_38025), .CD(n_61293), .Q(to_acu0
		[200]));
	notech_mux2 i_45679(.S(n_54955), .A(to_acu0[200]), .B(n_38842), .Z(n_38025
		));
	notech_reg to_acu0_reg_201(.CP(n_61854), .D(n_38031), .CD(n_61293), .Q(to_acu0
		[201]));
	notech_mux2 i_45687(.S(n_54955), .A(to_acu0[201]), .B(n_38845), .Z(n_38031
		));
	notech_reg to_acu0_reg_202(.CP(n_61854), .D(n_38037), .CD(n_61293), .Q(to_acu0
		[202]));
	notech_mux2 i_45695(.S(n_54985), .A(to_acu0[202]), .B(n_38848), .Z(n_38037
		));
	notech_reg to_acu0_reg_203(.CP(n_61854), .D(n_38043), .CD(n_61293), .Q(to_acu0
		[203]));
	notech_mux2 i_45703(.S(n_54985), .A(to_acu0[203]), .B(n_38851), .Z(n_38043
		));
	notech_reg to_acu0_reg_204(.CP(n_61854), .D(n_38049), .CD(n_61293), .Q(to_acu0
		[204]));
	notech_mux2 i_45711(.S(n_54985), .A(to_acu0[204]), .B(n_38854), .Z(n_38049
		));
	notech_reg to_acu0_reg_205(.CP(n_61854), .D(n_38055), .CD(n_61293), .Q(to_acu0
		[205]));
	notech_mux2 i_45719(.S(n_54985), .A(to_acu0[205]), .B(n_38857), .Z(n_38055
		));
	notech_reg to_acu0_reg_206(.CP(n_61854), .D(n_38061), .CD(n_61293), .Q(to_acu0
		[206]));
	notech_mux2 i_45727(.S(n_54985), .A(to_acu0[206]), .B(n_38860), .Z(n_38061
		));
	notech_reg to_acu0_reg_207(.CP(n_61852), .D(n_38067), .CD(n_61293), .Q(to_acu0
		[207]));
	notech_mux2 i_45735(.S(n_54985), .A(to_acu0[207]), .B(n_38863), .Z(n_38067
		));
	notech_reg to_acu0_reg_208(.CP(n_61847), .D(n_38073), .CD(n_61286), .Q(to_acu0
		[208]));
	notech_mux2 i_45743(.S(n_54985), .A(to_acu0[208]), .B(n_38866), .Z(n_38073
		));
	notech_reg to_acu0_reg_209(.CP(n_61847), .D(n_38079), .CD(n_61286), .Q(to_acu0
		[209]));
	notech_mux2 i_45751(.S(n_54985), .A(to_acu0[209]), .B(n_38869), .Z(n_38079
		));
	notech_reg to_acu0_reg_210(.CP(n_61847), .D(n_38085), .CD(n_61286), .Q(to_acu0
		[210]));
	notech_mux2 i_45759(.S(n_54985), .A(to_acu0[210]), .B(n_39310), .Z(n_38085
		));
	notech_reg over_seg0_reg_5(.CP(n_61847), .D(n_38091), .CD(n_61286), .Q(\over_seg0[5] 
		));
	notech_mux2 i_45767(.S(n_54985), .A(\over_seg0[5] ), .B(n_38339), .Z(n_38091
		));
	notech_reg opz0_reg_0(.CP(n_61847), .D(n_38097), .CD(n_61286), .Q(opz0[0
		]));
	notech_mux2 i_45775(.S(n_54955), .A(opz0[0]), .B(n_39857), .Z(n_38097)
		);
	notech_reg opz0_reg_1(.CP(n_61847), .D(n_38103), .CD(n_61286), .Q(opz0[1
		]));
	notech_mux2 i_45783(.S(n_54955), .A(opz0[1]), .B(n_39858), .Z(n_38103)
		);
	notech_reg_set opz0_reg_2(.CP(n_61847), .D(n_38109), .SD(n_61286), .Q(opz0
		[2]));
	notech_mux2 i_45791(.S(n_54985), .A(opz0[2]), .B(n_277591622), .Z(n_38109
		));
	notech_reg lenpc_reg_0(.CP(n_61847), .D(n_38115), .CD(n_61286), .Q(lenpc
		[0]));
	notech_mux2 i_45799(.S(n_3146), .A(n_38333), .B(lenpc[0]), .Z(n_38115)
		);
	notech_reg lenpc_reg_1(.CP(n_61847), .D(n_38121), .CD(n_61286), .Q(lenpc
		[1]));
	notech_mux2 i_45807(.S(n_3146), .A(n_38334), .B(lenpc[1]), .Z(n_38121)
		);
	notech_reg lenpc_reg_2(.CP(n_61847), .D(n_38127), .CD(n_61286), .Q(lenpc
		[2]));
	notech_mux2 i_45815(.S(n_3146), .A(n_38335), .B(lenpc[2]), .Z(n_38127)
		);
	notech_reg lenpc_reg_3(.CP(n_61847), .D(n_38133), .CD(n_61286), .Q(lenpc
		[3]));
	notech_mux2 i_45823(.S(n_3146), .A(n_38336), .B(lenpc[3]), .Z(n_38133)
		);
	notech_reg lenpc_reg_4(.CP(n_61842), .D(n_38139), .CD(n_61281), .Q(lenpc
		[4]));
	notech_mux2 i_45831(.S(n_3146), .A(n_38337), .B(lenpc[4]), .Z(n_38139)
		);
	notech_reg lenpc_reg_5(.CP(n_61842), .D(n_38145), .CD(n_61281), .Q(lenpc
		[5]));
	notech_mux2 i_45839(.S(n_3146), .A(n_38338), .B(lenpc[5]), .Z(n_38145)
		);
	notech_reg lenpc_reg_6(.CP(n_61842), .D(n_38151), .CD(n_61281), .Q(lenpc
		[6]));
	notech_mux2 i_45847(.S(n_3146), .A(n_170893329), .B(lenpc[6]), .Z(n_38151
		));
	notech_reg lenpc_reg_7(.CP(n_61842), .D(n_38157), .CD(n_61281), .Q(lenpc
		[7]));
	notech_mux2 i_45855(.S(n_3146), .A(n_160793228), .B(lenpc[7]), .Z(n_38157
		));
	notech_reg lenpc_reg_8(.CP(n_61842), .D(n_38163), .CD(n_61281), .Q(lenpc
		[8]));
	notech_mux2 i_45863(.S(n_3146), .A(n_108392704), .B(lenpc[8]), .Z(n_38163
		));
	notech_reg lenpc_reg_9(.CP(n_61847), .D(n_38169), .CD(n_61286), .Q(lenpc
		[9]));
	notech_mux2 i_45871(.S(n_3146), .A(n_108492705), .B(lenpc[9]), .Z(n_38169
		));
	notech_reg lenpc_reg_10(.CP(n_61847), .D(n_38175), .CD(n_61286), .Q(lenpc
		[10]));
	notech_mux2 i_45879(.S(n_3146), .A(n_108592706), .B(lenpc[10]), .Z(n_38175
		));
	notech_reg lenpc_reg_11(.CP(n_61847), .D(n_38181), .CD(n_61281), .Q(lenpc
		[11]));
	notech_mux2 i_45887(.S(n_3146), .A(n_108692707), .B(lenpc[11]), .Z(n_38181
		));
	notech_reg lenpc_reg_12(.CP(n_61842), .D(n_38187), .CD(n_61281), .Q(lenpc
		[12]));
	notech_mux2 i_45895(.S(n_3146), .A(n_108792708), .B(lenpc[12]), .Z(n_38187
		));
	notech_reg lenpc_reg_13(.CP(n_61847), .D(n_38193), .CD(n_61281), .Q(lenpc
		[13]));
	notech_mux2 i_45903(.S(n_3146), .A(n_108892709), .B(lenpc[13]), .Z(n_38193
		));
	notech_reg lenpc_reg_14(.CP(n_61849), .D(n_38199), .CD(n_61288), .Q(lenpc
		[14]));
	notech_mux2 i_45911(.S(n_3146), .A(n_108992710), .B(lenpc[14]), .Z(n_38199
		));
	notech_reg lenpc_reg_15(.CP(n_61849), .D(n_38205), .CD(n_61288), .Q(lenpc
		[15]));
	notech_mux2 i_45919(.S(n_3146), .A(n_109092711), .B(lenpc[15]), .Z(n_38205
		));
	notech_reg lenpc_reg_16(.CP(n_61849), .D(n_38211), .CD(n_61288), .Q(lenpc
		[16]));
	notech_mux2 i_45927(.S(n_58455), .A(n_109192712), .B(lenpc[16]), .Z(n_38211
		));
	notech_reg lenpc_reg_17(.CP(n_61849), .D(n_38217), .CD(n_61288), .Q(lenpc
		[17]));
	notech_mux2 i_45935(.S(n_58455), .A(n_109292713), .B(lenpc[17]), .Z(n_38217
		));
	notech_reg lenpc_reg_18(.CP(n_61849), .D(n_38223), .CD(n_61288), .Q(lenpc
		[18]));
	notech_mux2 i_45943(.S(n_58455), .A(n_109392714), .B(lenpc[18]), .Z(n_38223
		));
	notech_reg lenpc_reg_19(.CP(n_61849), .D(n_38229), .CD(n_61288), .Q(lenpc
		[19]));
	notech_mux2 i_45951(.S(n_58455), .A(n_109492715), .B(lenpc[19]), .Z(n_38229
		));
	notech_reg lenpc_reg_20(.CP(n_61849), .D(n_38235), .CD(n_61288), .Q(lenpc
		[20]));
	notech_mux2 i_45959(.S(n_58455), .A(n_109592716), .B(lenpc[20]), .Z(n_38235
		));
	notech_reg lenpc_reg_21(.CP(n_61849), .D(n_38241), .CD(n_61288), .Q(lenpc
		[21]));
	notech_mux2 i_45967(.S(n_58455), .A(n_109692717), .B(lenpc[21]), .Z(n_38241
		));
	notech_reg lenpc_reg_22(.CP(n_61849), .D(n_38247), .CD(n_61288), .Q(lenpc
		[22]));
	notech_mux2 i_45975(.S(n_58455), .A(n_109792718), .B(lenpc[22]), .Z(n_38247
		));
	notech_reg lenpc_reg_23(.CP(n_61849), .D(n_38253), .CD(n_61288), .Q(lenpc
		[23]));
	notech_mux2 i_45983(.S(n_58455), .A(n_109892719), .B(lenpc[23]), .Z(n_38253
		));
	notech_reg lenpc_reg_24(.CP(n_61849), .D(n_38259), .CD(n_61288), .Q(lenpc
		[24]));
	notech_mux2 i_45991(.S(n_58455), .A(n_109992720), .B(lenpc[24]), .Z(n_38259
		));
	notech_reg lenpc_reg_25(.CP(n_61849), .D(n_38265), .CD(n_61286), .Q(lenpc
		[25]));
	notech_mux2 i_45999(.S(n_58455), .A(n_110092721), .B(lenpc[25]), .Z(n_38265
		));
	notech_nand3 i_26774742(.A(cpl[0]), .B(cpl[1]), .C(pg_fault), .Z(n_1418)
		);
	notech_reg lenpc_reg_26(.CP(n_61849), .D(n_38271), .CD(n_61286), .Q(lenpc
		[26]));
	notech_mux2 i_46007(.S(n_3146), .A(n_110192722), .B(lenpc[26]), .Z(n_38271
		));
	notech_reg lenpc_reg_27(.CP(n_61847), .D(n_38277), .CD(n_61286), .Q(lenpc
		[27]));
	notech_mux2 i_46015(.S(n_58455), .A(n_110292723), .B(lenpc[27]), .Z(n_38277
		));
	notech_reg lenpc_reg_28(.CP(n_61847), .D(n_38283), .CD(n_61286), .Q(lenpc
		[28]));
	notech_mux2 i_46023(.S(n_58455), .A(n_110392724), .B(lenpc[28]), .Z(n_38283
		));
	notech_reg lenpc_reg_29(.CP(n_61847), .D(n_38289), .CD(n_61286), .Q(lenpc
		[29]));
	notech_mux2 i_46031(.S(n_58455), .A(n_110492725), .B(lenpc[29]), .Z(n_38289
		));
	notech_reg lenpc_reg_30(.CP(n_61849), .D(n_38295), .CD(n_61288), .Q(lenpc
		[30]));
	notech_mux2 i_46039(.S(n_58455), .A(n_110592726), .B(lenpc[30]), .Z(n_38295
		));
	notech_reg lenpc_reg_31(.CP(n_61849), .D(n_38301), .CD(n_61288), .Q(lenpc
		[31]));
	notech_mux2 i_46047(.S(n_58455), .A(n_110692727), .B(lenpc[31]), .Z(n_38301
		));
	notech_reg reps0_reg_0(.CP(n_61849), .D(n_38307), .CD(n_61288), .Q(reps0
		[0]));
	notech_mux2 i_46055(.S(n_54985), .A(reps0[0]), .B(n_38519), .Z(n_38307)
		);
	notech_nao3 i_074990(.A(n_18050174), .B(n_1568), .C(n_1490), .Z(n_1411)
		);
	notech_reg reps0_reg_1(.CP(n_61849), .D(n_38313), .CD(n_61288), .Q(reps0
		[1]));
	notech_mux2 i_46063(.S(n_54985), .A(reps0[1]), .B(n_38331), .Z(n_38313)
		);
	notech_reg reps0_reg_2(.CP(n_61849), .D(n_38319), .CD(n_61288), .Q(reps0
		[2]));
	notech_mux2 i_46071(.S(n_54985), .A(reps0[2]), .B(n_38332), .Z(n_38319)
		);
	notech_inv i_51265(.A(n_168393304), .Z(n_38325));
	notech_inv i_51266(.A(n_168593306), .Z(n_38326));
	notech_inv i_51267(.A(n_134692967), .Z(n_38327));
	notech_inv i_51268(.A(n_9539), .Z(n_38328));
	notech_inv i_51269(.A(n_5408), .Z(n_38329));
	notech_inv i_51270(.A(n_1995), .Z(n_38330));
	notech_inv i_51271(.A(n_2797), .Z(n_38331));
	notech_inv i_51272(.A(n_2795), .Z(n_38332));
	notech_inv i_51273(.A(n_2793), .Z(n_38333));
	notech_inv i_51274(.A(n_2790), .Z(n_38334));
	notech_inv i_51275(.A(n_2787), .Z(n_38335));
	notech_inv i_51276(.A(n_2784), .Z(n_38336));
	notech_inv i_51277(.A(n_278191628), .Z(n_38337));
	notech_inv i_51278(.A(n_277891625), .Z(n_38338));
	notech_inv i_51279(.A(n_277391620), .Z(n_38339));
	notech_inv i_51280(.A(n_277191618), .Z(n_38340));
	notech_inv i_51281(.A(n_276991616), .Z(n_38341));
	notech_inv i_51282(.A(n_276791614), .Z(n_38342));
	notech_inv i_51283(.A(n_276591612), .Z(n_38343));
	notech_inv i_51284(.A(n_276391610), .Z(n_38344));
	notech_inv i_51285(.A(n_276191608), .Z(n_38345));
	notech_inv i_51286(.A(n_275991606), .Z(n_38346));
	notech_inv i_51287(.A(n_275791604), .Z(n_38347));
	notech_inv i_51288(.A(n_275591602), .Z(n_38348));
	notech_inv i_51289(.A(n_275391600), .Z(n_38349));
	notech_inv i_51290(.A(n_275191598), .Z(n_38350));
	notech_inv i_51291(.A(n_274991596), .Z(n_38351));
	notech_inv i_51292(.A(n_274791594), .Z(n_38352));
	notech_inv i_51293(.A(n_274591592), .Z(n_38353));
	notech_inv i_51294(.A(n_274391590), .Z(n_38354));
	notech_inv i_51295(.A(n_274191588), .Z(n_38355));
	notech_inv i_51296(.A(n_273991586), .Z(n_38356));
	notech_inv i_51297(.A(n_273791584), .Z(n_38357));
	notech_inv i_51298(.A(n_273591582), .Z(n_38358));
	notech_inv i_51299(.A(n_273391580), .Z(n_38359));
	notech_inv i_51300(.A(n_273191578), .Z(n_38360));
	notech_inv i_51301(.A(n_272991576), .Z(n_38361));
	notech_inv i_51302(.A(n_272791574), .Z(n_38362));
	notech_inv i_51303(.A(n_272591572), .Z(n_38363));
	notech_inv i_51304(.A(n_272391570), .Z(n_38364));
	notech_inv i_51305(.A(n_272191568), .Z(n_38365));
	notech_inv i_51306(.A(n_271991566), .Z(n_38366));
	notech_inv i_51307(.A(n_271791564), .Z(n_38367));
	notech_inv i_51308(.A(n_271591562), .Z(n_38368));
	notech_inv i_51309(.A(n_271391560), .Z(n_38369));
	notech_inv i_51310(.A(n_271191558), .Z(n_38370));
	notech_inv i_51311(.A(n_270991556), .Z(n_38371));
	notech_inv i_51312(.A(n_270791554), .Z(n_38372));
	notech_inv i_51313(.A(n_270591552), .Z(n_38373));
	notech_inv i_51314(.A(n_270391550), .Z(n_38374));
	notech_inv i_51315(.A(n_270191548), .Z(n_38375));
	notech_inv i_51316(.A(n_269991546), .Z(n_38376));
	notech_inv i_51317(.A(n_269791544), .Z(n_38377));
	notech_inv i_51318(.A(n_269591542), .Z(n_38378));
	notech_inv i_51319(.A(n_269391540), .Z(n_38379));
	notech_inv i_51320(.A(n_269191538), .Z(n_38380));
	notech_inv i_51321(.A(n_268991536), .Z(n_38381));
	notech_inv i_51322(.A(n_268791534), .Z(n_38382));
	notech_inv i_51323(.A(n_268591532), .Z(n_38383));
	notech_inv i_51324(.A(n_268391530), .Z(n_38384));
	notech_inv i_51325(.A(n_268191528), .Z(n_38385));
	notech_inv i_51326(.A(n_267991526), .Z(n_38386));
	notech_inv i_51327(.A(n_267791524), .Z(n_38387));
	notech_inv i_51328(.A(n_267591522), .Z(n_38388));
	notech_inv i_51329(.A(n_267391520), .Z(n_38389));
	notech_inv i_51330(.A(n_267191518), .Z(n_38390));
	notech_inv i_51331(.A(n_266991516), .Z(n_38391));
	notech_inv i_51332(.A(n_266791514), .Z(n_38392));
	notech_inv i_51333(.A(n_266591512), .Z(n_38393));
	notech_inv i_51334(.A(n_266391510), .Z(n_38394));
	notech_inv i_51335(.A(n_266191508), .Z(n_38395));
	notech_inv i_51336(.A(n_265291499), .Z(n_38396));
	notech_inv i_51337(.A(n_265091497), .Z(n_38397));
	notech_inv i_51338(.A(n_264891495), .Z(n_38398));
	notech_inv i_51339(.A(n_264691493), .Z(n_38399));
	notech_inv i_51340(.A(n_264491491), .Z(n_38400));
	notech_inv i_51341(.A(n_264291489), .Z(n_38401));
	notech_inv i_51342(.A(n_264091487), .Z(n_38402));
	notech_inv i_51343(.A(n_263891485), .Z(n_38403));
	notech_inv i_51344(.A(n_263691483), .Z(n_38404));
	notech_inv i_51345(.A(n_263491481), .Z(n_38405));
	notech_inv i_51346(.A(n_262791474), .Z(n_38406));
	notech_inv i_51347(.A(n_262191468), .Z(n_38407));
	notech_inv i_51348(.A(n_162793248), .Z(n_38408));
	notech_inv i_51349(.A(n_260691453), .Z(n_38409));
	notech_inv i_51350(.A(n_260491451), .Z(n_38410));
	notech_inv i_51351(.A(n_170793328), .Z(n_38411));
	notech_inv i_51352(.A(n_260291449), .Z(n_38412));
	notech_inv i_51353(.A(n_260091447), .Z(n_38413));
	notech_inv i_51354(.A(n_259891445), .Z(n_38414));
	notech_inv i_51355(.A(n_2217), .Z(n_38415));
	notech_inv i_51356(.A(n_259691443), .Z(n_38416));
	notech_inv i_51357(.A(n_2058), .Z(start));
	notech_inv i_51358(.A(n_259491441), .Z(n_38418));
	notech_inv i_51359(.A(n_259291439), .Z(n_38419));
	notech_inv i_51360(.A(n_259091437), .Z(n_38420));
	notech_inv i_51361(.A(term_f), .Z(n_38421));
	notech_inv i_51362(.A(n_258891435), .Z(n_38422));
	notech_inv i_51363(.A(n_258691433), .Z(n_38423));
	notech_inv i_51364(.A(n_258491431), .Z(n_38424));
	notech_inv i_51365(.A(\fpu_indrm[0] ), .Z(n_38425));
	notech_inv i_51366(.A(n_258291429), .Z(n_38426));
	notech_inv i_51367(.A(n_258091427), .Z(n_38427));
	notech_inv i_51368(.A(\fpu_indrm[2] ), .Z(n_38428));
	notech_inv i_51369(.A(n_257891425), .Z(n_38429));
	notech_inv i_51370(.A(n_257691423), .Z(n_38430));
	notech_inv i_51371(.A(\fpu_indrm[3] ), .Z(n_38431));
	notech_inv i_51372(.A(n_257491421), .Z(n_38432));
	notech_inv i_51373(.A(n_257291419), .Z(n_38433));
	notech_inv i_51374(.A(\fpu_indrm[4] ), .Z(n_38434));
	notech_inv i_51375(.A(n_257091417), .Z(n_38435));
	notech_inv i_51376(.A(n_256891415), .Z(n_38436));
	notech_inv i_51377(.A(n_256691413), .Z(n_38437));
	notech_inv i_51378(.A(n_256491411), .Z(n_38438));
	notech_inv i_51379(.A(n_256291409), .Z(n_38439));
	notech_inv i_51380(.A(n_256091407), .Z(n_38440));
	notech_inv i_51381(.A(n_255891405), .Z(n_38441));
	notech_inv i_51382(.A(n_255691403), .Z(n_38442));
	notech_inv i_51383(.A(n_255491401), .Z(n_38443));
	notech_inv i_51384(.A(n_255291399), .Z(n_38444));
	notech_inv i_51385(.A(n_255091397), .Z(n_38445));
	notech_inv i_51386(.A(n_254891395), .Z(n_38446));
	notech_inv i_51387(.A(n_254691393), .Z(n_38447));
	notech_inv i_51388(.A(n_254491391), .Z(n_38448));
	notech_inv i_51389(.A(n_254291389), .Z(n_38449));
	notech_inv i_51390(.A(n_254091387), .Z(n_38450));
	notech_inv i_51391(.A(n_253891385), .Z(n_38451));
	notech_inv i_51392(.A(n_253691383), .Z(n_38452));
	notech_inv i_51393(.A(n_253491381), .Z(n_38453));
	notech_inv i_51394(.A(n_253291379), .Z(n_38454));
	notech_inv i_51395(.A(n_253091377), .Z(n_38455));
	notech_inv i_51396(.A(\imm2[0] ), .Z(n_38456));
	notech_inv i_51397(.A(n_252891375), .Z(n_38457));
	notech_inv i_51398(.A(\imm2[1] ), .Z(n_38458));
	notech_inv i_51399(.A(n_252691373), .Z(n_38459));
	notech_inv i_51400(.A(\imm2[2] ), .Z(n_38460));
	notech_inv i_51401(.A(n_252491371), .Z(n_38461));
	notech_inv i_51402(.A(\imm2[3] ), .Z(n_38462));
	notech_inv i_51403(.A(n_252291369), .Z(n_38463));
	notech_inv i_51404(.A(\imm2[4] ), .Z(n_38464));
	notech_inv i_51405(.A(\imm2[5] ), .Z(n_38465));
	notech_inv i_51406(.A(\imm2[6] ), .Z(n_38466));
	notech_inv i_51407(.A(\imm2[7] ), .Z(n_38467));
	notech_inv i_51408(.A(\imm2[8] ), .Z(n_38468));
	notech_inv i_51409(.A(\imm2[9] ), .Z(n_38469));
	notech_inv i_51410(.A(\imm2[10] ), .Z(n_38470));
	notech_inv i_51411(.A(\imm2[11] ), .Z(n_38471));
	notech_inv i_51412(.A(\imm2[12] ), .Z(n_38472));
	notech_inv i_51413(.A(\imm2[13] ), .Z(n_38473));
	notech_inv i_51414(.A(\imm2[14] ), .Z(n_38474));
	notech_inv i_51415(.A(\imm2[15] ), .Z(n_38475));
	notech_inv i_51416(.A(\imm2[16] ), .Z(n_38476));
	notech_inv i_51417(.A(\imm2[17] ), .Z(n_38477));
	notech_inv i_51418(.A(\imm2[18] ), .Z(n_38478));
	notech_inv i_51419(.A(\imm2[19] ), .Z(n_38479));
	notech_inv i_51420(.A(\imm2[20] ), .Z(n_38480));
	notech_inv i_51421(.A(\imm2[21] ), .Z(n_38481));
	notech_inv i_51422(.A(\imm2[22] ), .Z(n_38482));
	notech_inv i_51423(.A(\imm2[23] ), .Z(n_38483));
	notech_inv i_51424(.A(\imm2[24] ), .Z(n_38484));
	notech_inv i_51425(.A(\imm2[25] ), .Z(n_38485));
	notech_inv i_51426(.A(\imm2[26] ), .Z(n_38486));
	notech_inv i_51427(.A(\imm2[27] ), .Z(n_38487));
	notech_inv i_51428(.A(\imm2[28] ), .Z(n_38488));
	notech_inv i_51429(.A(\imm2[29] ), .Z(n_38489));
	notech_inv i_51430(.A(\imm2[30] ), .Z(n_38490));
	notech_inv i_51431(.A(\imm2[31] ), .Z(n_38491));
	notech_inv i_51432(.A(\imm2[32] ), .Z(n_38492));
	notech_inv i_51433(.A(\imm2[33] ), .Z(n_38493));
	notech_inv i_51434(.A(\imm2[34] ), .Z(n_38494));
	notech_inv i_51435(.A(\imm2[35] ), .Z(n_38495));
	notech_inv i_51436(.A(\imm2[36] ), .Z(n_38496));
	notech_inv i_51437(.A(\imm2[37] ), .Z(n_38497));
	notech_inv i_51438(.A(\imm2[38] ), .Z(n_38498));
	notech_inv i_51439(.A(\imm2[39] ), .Z(n_38499));
	notech_inv i_51440(.A(\imm2[40] ), .Z(n_38500));
	notech_inv i_51441(.A(\imm2[41] ), .Z(n_38501));
	notech_inv i_51442(.A(\imm2[42] ), .Z(n_38502));
	notech_inv i_51443(.A(\imm2[43] ), .Z(n_38503));
	notech_inv i_51444(.A(\imm2[44] ), .Z(n_38504));
	notech_inv i_51445(.A(\imm2[45] ), .Z(n_38505));
	notech_inv i_51446(.A(\imm2[46] ), .Z(n_38506));
	notech_inv i_51447(.A(\imm2[47] ), .Z(n_38507));
	notech_inv i_51448(.A(n_2218), .Z(n_38508));
	notech_inv i_51449(.A(\imm1[0] ), .Z(n_38509));
	notech_inv i_51450(.A(n_2132), .Z(n_38510));
	notech_inv i_51451(.A(\imm1[1] ), .Z(n_38511));
	notech_inv i_51452(.A(\imm1[2] ), .Z(n_38512));
	notech_inv i_51453(.A(\imm1[3] ), .Z(n_38513));
	notech_inv i_51454(.A(\imm1[4] ), .Z(n_38514));
	notech_inv i_51455(.A(\imm1[5] ), .Z(n_38515));
	notech_inv i_51456(.A(n_261391460), .Z(n_38516));
	notech_inv i_51457(.A(n_3813), .Z(n_38517));
	notech_inv i_51458(.A(\imm1[6] ), .Z(n_38518));
	notech_inv i_51459(.A(n_3812), .Z(n_38519));
	notech_inv i_51460(.A(\imm1[7] ), .Z(n_38520));
	notech_inv i_51461(.A(n_3811), .Z(n_38521));
	notech_inv i_51462(.A(\imm1[8] ), .Z(n_38522));
	notech_inv i_51463(.A(n_3809), .Z(n_38523));
	notech_inv i_51464(.A(\imm1[9] ), .Z(n_38524));
	notech_inv i_51465(.A(n_3808), .Z(n_38525));
	notech_inv i_51466(.A(\imm1[10] ), .Z(n_38526));
	notech_inv i_51467(.A(n_3806), .Z(n_38527));
	notech_inv i_51468(.A(\imm1[11] ), .Z(n_38528));
	notech_inv i_51469(.A(n_3805), .Z(n_38529));
	notech_inv i_51470(.A(\imm1[12] ), .Z(n_38530));
	notech_inv i_51471(.A(n_3803), .Z(n_38531));
	notech_inv i_51472(.A(\imm1[13] ), .Z(n_38532));
	notech_inv i_51473(.A(n_3801), .Z(n_38533));
	notech_inv i_51474(.A(\imm1[14] ), .Z(n_38534));
	notech_inv i_51475(.A(n_3799), .Z(n_38535));
	notech_inv i_51476(.A(\imm1[15] ), .Z(n_38536));
	notech_inv i_51477(.A(n_3798), .Z(n_38537));
	notech_inv i_51478(.A(\imm1[16] ), .Z(n_38538));
	notech_inv i_51479(.A(n_3796), .Z(n_38539));
	notech_inv i_51480(.A(\imm1[17] ), .Z(n_38540));
	notech_inv i_51481(.A(n_3794), .Z(n_38541));
	notech_inv i_51482(.A(\imm1[18] ), .Z(n_38542));
	notech_inv i_51483(.A(n_3792), .Z(n_38543));
	notech_inv i_51484(.A(\imm1[19] ), .Z(n_38544));
	notech_inv i_51485(.A(n_3791), .Z(n_38545));
	notech_inv i_51486(.A(\imm1[20] ), .Z(n_38546));
	notech_inv i_51487(.A(n_3790), .Z(n_38547));
	notech_inv i_51488(.A(\imm1[21] ), .Z(n_38548));
	notech_inv i_51489(.A(n_3789), .Z(n_38549));
	notech_inv i_51490(.A(\imm1[22] ), .Z(n_38550));
	notech_inv i_51491(.A(n_3787), .Z(n_38551));
	notech_inv i_51492(.A(\imm1[23] ), .Z(n_38552));
	notech_inv i_51493(.A(n_3785), .Z(n_38553));
	notech_inv i_51494(.A(\imm1[24] ), .Z(n_38554));
	notech_inv i_51495(.A(n_3783), .Z(n_38555));
	notech_inv i_51496(.A(\imm1[25] ), .Z(n_38556));
	notech_inv i_51497(.A(n_3781), .Z(n_38557));
	notech_inv i_51498(.A(\imm1[26] ), .Z(n_38558));
	notech_inv i_51499(.A(n_3779), .Z(n_38559));
	notech_inv i_51500(.A(\imm1[27] ), .Z(n_38560));
	notech_inv i_51501(.A(n_3777), .Z(n_38561));
	notech_inv i_51502(.A(\imm1[28] ), .Z(n_38562));
	notech_inv i_51503(.A(n_3776), .Z(n_38563));
	notech_inv i_51504(.A(\imm1[29] ), .Z(n_38564));
	notech_inv i_51505(.A(n_3775), .Z(n_38565));
	notech_inv i_51506(.A(\imm1[30] ), .Z(n_38566));
	notech_inv i_51507(.A(n_3774), .Z(n_38567));
	notech_inv i_51508(.A(\imm1[31] ), .Z(n_38568));
	notech_inv i_51509(.A(n_3773), .Z(n_38569));
	notech_inv i_51510(.A(\imm1[32] ), .Z(n_38570));
	notech_inv i_51511(.A(n_3772), .Z(n_38571));
	notech_inv i_51512(.A(\imm1[33] ), .Z(n_38572));
	notech_inv i_51513(.A(n_3771), .Z(n_38573));
	notech_inv i_51514(.A(\imm1[34] ), .Z(n_38574));
	notech_inv i_51515(.A(n_3770), .Z(n_38575));
	notech_inv i_51516(.A(\imm1[35] ), .Z(n_38576));
	notech_inv i_51517(.A(n_3768), .Z(n_38577));
	notech_inv i_51518(.A(\imm1[36] ), .Z(n_38578));
	notech_inv i_51519(.A(n_46345), .Z(n_38579));
	notech_inv i_51520(.A(\imm1[37] ), .Z(n_38580));
	notech_inv i_51521(.A(n_3766), .Z(n_38581));
	notech_inv i_51522(.A(n_46351), .Z(n_38582));
	notech_inv i_51523(.A(\imm1[38] ), .Z(n_38583));
	notech_inv i_51524(.A(n_46357), .Z(n_38584));
	notech_inv i_51525(.A(\imm1[39] ), .Z(n_38585));
	notech_inv i_51526(.A(n_3764), .Z(n_38586));
	notech_inv i_51527(.A(n_46363), .Z(n_38587));
	notech_inv i_51528(.A(\imm1[40] ), .Z(n_38588));
	notech_inv i_51529(.A(n_3762), .Z(n_38589));
	notech_inv i_51530(.A(\imm1[41] ), .Z(n_38590));
	notech_inv i_51531(.A(n_3760), .Z(n_38591));
	notech_inv i_51532(.A(\imm1[42] ), .Z(n_38592));
	notech_inv i_51533(.A(n_3758), .Z(n_38593));
	notech_inv i_51534(.A(\imm1[43] ), .Z(n_38594));
	notech_inv i_51535(.A(n_46387), .Z(n_38595));
	notech_inv i_51536(.A(\imm1[44] ), .Z(n_38596));
	notech_inv i_51537(.A(n_3756), .Z(n_38597));
	notech_inv i_51538(.A(\imm1[45] ), .Z(n_38598));
	notech_inv i_51539(.A(n_3754), .Z(n_38599));
	notech_inv i_51540(.A(\imm1[46] ), .Z(n_38600));
	notech_inv i_51541(.A(n_3752), .Z(n_38601));
	notech_inv i_51542(.A(\imm1[47] ), .Z(n_38602));
	notech_inv i_51543(.A(n_3750), .Z(n_38603));
	notech_inv i_51544(.A(n_3748), .Z(n_38604));
	notech_inv i_51545(.A(trig_itf), .Z(n_38605));
	notech_inv i_51546(.A(intf), .Z(n_38606));
	notech_inv i_51547(.A(n_3746), .Z(n_38607));
	notech_inv i_51548(.A(n_3744), .Z(n_38608));
	notech_inv i_51549(.A(n_3742), .Z(n_38609));
	notech_inv i_51550(.A(n_3740), .Z(n_38610));
	notech_inv i_51551(.A(n_3738), .Z(n_38611));
	notech_inv i_51552(.A(n_3736), .Z(n_38612));
	notech_inv i_51553(.A(n_3734), .Z(n_38613));
	notech_inv i_51554(.A(n_3732), .Z(n_38614));
	notech_inv i_51555(.A(n_3730), .Z(n_38615));
	notech_inv i_51556(.A(n_3728), .Z(n_38616));
	notech_inv i_51557(.A(n_3726), .Z(n_38617));
	notech_inv i_51558(.A(n_3724), .Z(n_38618));
	notech_inv i_51559(.A(n_3722), .Z(n_38619));
	notech_inv i_51560(.A(n_3720), .Z(n_38620));
	notech_inv i_51561(.A(n_3718), .Z(n_38621));
	notech_inv i_51562(.A(n_3716), .Z(n_38622));
	notech_inv i_51563(.A(n_3714), .Z(n_38623));
	notech_inv i_51564(.A(ififo_rvect1[0]), .Z(n_38624));
	notech_inv i_51565(.A(ififo_rvect1[1]), .Z(n_38625));
	notech_inv i_51566(.A(n_3712), .Z(n_38626));
	notech_inv i_51567(.A(ififo_rvect1[2]), .Z(n_38627));
	notech_inv i_51568(.A(ififo_rvect1[3]), .Z(n_38628));
	notech_inv i_51569(.A(n_3710), .Z(n_38629));
	notech_inv i_51570(.A(ififo_rvect1[4]), .Z(n_38630));
	notech_inv i_51571(.A(ififo_rvect1[5]), .Z(n_38631));
	notech_inv i_51572(.A(n_3708), .Z(n_38632));
	notech_inv i_51573(.A(ififo_rvect1[6]), .Z(n_38633));
	notech_inv i_51574(.A(ififo_rvect1[7]), .Z(n_38634));
	notech_inv i_51575(.A(n_3706), .Z(n_38635));
	notech_inv i_51576(.A(n_3704), .Z(n_38636));
	notech_inv i_51577(.A(n_3702), .Z(n_38637));
	notech_inv i_51578(.A(int_excl[2]), .Z(n_38638));
	notech_inv i_51579(.A(n_3701), .Z(n_38639));
	notech_inv i_51580(.A(n_3700), .Z(n_38640));
	notech_inv i_51581(.A(n_3699), .Z(n_38641));
	notech_inv i_51582(.A(n_3698), .Z(n_38642));
	notech_inv i_51583(.A(n_3697), .Z(n_38643));
	notech_inv i_51584(.A(n_3696), .Z(n_38644));
	notech_inv i_51585(.A(n_3694), .Z(n_38645));
	notech_inv i_51586(.A(n_3692), .Z(n_38646));
	notech_inv i_51587(.A(n_44589), .Z(n_38647));
	notech_inv i_51588(.A(n_3691), .Z(n_38648));
	notech_inv i_51589(.A(n_49822), .Z(n_38649));
	notech_inv i_51590(.A(n_3690), .Z(n_38650));
	notech_inv i_51591(.A(n_3689), .Z(n_38651));
	notech_inv i_51592(.A(n_3688), .Z(n_38652));
	notech_inv i_51593(.A(i_ptr[2]), .Z(n_38653));
	notech_inv i_51594(.A(n_3686), .Z(n_38654));
	notech_inv i_51595(.A(n_3684), .Z(n_38655));
	notech_inv i_51596(.A(idx_deco[0]), .Z(n_38656));
	notech_inv i_51597(.A(n_3682), .Z(n_38657));
	notech_inv i_51598(.A(n_3680), .Z(n_38658));
	notech_inv i_51599(.A(fsm[0]), .Z(n_38659));
	notech_inv i_51600(.A(n_3678), .Z(n_38660));
	notech_inv i_51601(.A(fsm[1]), .Z(n_38661));
	notech_inv i_51602(.A(n_3676), .Z(n_38662));
	notech_inv i_51603(.A(n_3674), .Z(n_38663));
	notech_inv i_51604(.A(fsm[4]), .Z(n_38664));
	notech_inv i_51605(.A(n_3672), .Z(n_38665));
	notech_inv i_51606(.A(repz), .Z(n_38666));
	notech_inv i_51607(.A(n_3670), .Z(n_38667));
	notech_inv i_51608(.A(rep), .Z(n_38668));
	notech_inv i_51609(.A(reps2[0]), .Z(n_38669));
	notech_inv i_51610(.A(n_3668), .Z(n_38670));
	notech_inv i_51611(.A(reps2[1]), .Z(n_38671));
	notech_inv i_51612(.A(reps2[2]), .Z(n_38672));
	notech_inv i_51613(.A(n_3666), .Z(n_38673));
	notech_inv i_51614(.A(reps1[0]), .Z(n_38674));
	notech_inv i_51615(.A(n_3664), .Z(n_38675));
	notech_inv i_51616(.A(reps1[1]), .Z(n_38676));
	notech_inv i_51617(.A(n_3662), .Z(n_38677));
	notech_inv i_51618(.A(reps1[2]), .Z(n_38678));
	notech_inv i_51619(.A(n_3660), .Z(n_38679));
	notech_inv i_51620(.A(inst_deco2[0]), .Z(n_38680));
	notech_inv i_51621(.A(inst_deco2[1]), .Z(n_38681));
	notech_inv i_51622(.A(n_3658), .Z(n_38682));
	notech_inv i_51623(.A(inst_deco2[2]), .Z(n_38683));
	notech_inv i_51624(.A(inst_deco2[3]), .Z(n_38684));
	notech_inv i_51625(.A(n_3656), .Z(n_38685));
	notech_inv i_51626(.A(inst_deco2[4]), .Z(n_38686));
	notech_inv i_51627(.A(inst_deco2[5]), .Z(n_38687));
	notech_inv i_51628(.A(n_3654), .Z(n_38688));
	notech_inv i_51629(.A(inst_deco2[6]), .Z(n_38689));
	notech_inv i_51630(.A(inst_deco2[7]), .Z(n_38690));
	notech_inv i_51631(.A(n_3652), .Z(n_38691));
	notech_inv i_51632(.A(inst_deco2[8]), .Z(n_38692));
	notech_inv i_51633(.A(inst_deco2[9]), .Z(n_38693));
	notech_inv i_51634(.A(n_3650), .Z(n_38694));
	notech_inv i_51635(.A(inst_deco2[10]), .Z(n_38695));
	notech_inv i_51636(.A(inst_deco2[11]), .Z(n_38696));
	notech_inv i_51637(.A(n_3648), .Z(n_38697));
	notech_inv i_51638(.A(inst_deco2[12]), .Z(n_38698));
	notech_inv i_51639(.A(inst_deco2[13]), .Z(n_38699));
	notech_inv i_51640(.A(n_3646), .Z(n_38700));
	notech_inv i_51641(.A(inst_deco2[14]), .Z(n_38701));
	notech_inv i_51642(.A(inst_deco2[15]), .Z(n_38702));
	notech_inv i_51643(.A(n_3644), .Z(n_38703));
	notech_inv i_51644(.A(inst_deco2[16]), .Z(n_38704));
	notech_inv i_51645(.A(inst_deco2[17]), .Z(n_38705));
	notech_inv i_51646(.A(n_3642), .Z(n_38706));
	notech_inv i_51647(.A(inst_deco2[18]), .Z(n_38707));
	notech_inv i_51648(.A(inst_deco2[19]), .Z(n_38708));
	notech_inv i_51649(.A(n_3640), .Z(n_38709));
	notech_inv i_51650(.A(inst_deco2[20]), .Z(n_38710));
	notech_inv i_51651(.A(inst_deco2[21]), .Z(n_38711));
	notech_inv i_51652(.A(n_3638), .Z(n_38712));
	notech_inv i_51653(.A(inst_deco2[22]), .Z(n_38713));
	notech_inv i_51654(.A(inst_deco2[23]), .Z(n_38714));
	notech_inv i_51655(.A(n_3636), .Z(n_38715));
	notech_inv i_51656(.A(inst_deco2[24]), .Z(n_38716));
	notech_inv i_51657(.A(inst_deco2[25]), .Z(n_38717));
	notech_inv i_51658(.A(n_3634), .Z(n_38718));
	notech_inv i_51659(.A(inst_deco2[26]), .Z(n_38719));
	notech_inv i_51660(.A(inst_deco2[27]), .Z(n_38720));
	notech_inv i_51661(.A(n_3632), .Z(n_38721));
	notech_inv i_51662(.A(inst_deco2[28]), .Z(n_38722));
	notech_inv i_51663(.A(inst_deco2[29]), .Z(n_38723));
	notech_inv i_51664(.A(n_3630), .Z(n_38724));
	notech_inv i_51665(.A(inst_deco2[30]), .Z(n_38725));
	notech_inv i_51666(.A(inst_deco2[31]), .Z(n_38726));
	notech_inv i_51667(.A(n_3628), .Z(n_38727));
	notech_inv i_51668(.A(inst_deco2[32]), .Z(n_38728));
	notech_inv i_51669(.A(inst_deco2[33]), .Z(n_38729));
	notech_inv i_51670(.A(n_3626), .Z(n_38730));
	notech_inv i_51671(.A(inst_deco2[34]), .Z(n_38731));
	notech_inv i_51672(.A(inst_deco2[35]), .Z(n_38732));
	notech_inv i_51673(.A(n_3625), .Z(n_38733));
	notech_inv i_51674(.A(inst_deco2[36]), .Z(n_38734));
	notech_inv i_51675(.A(inst_deco2[37]), .Z(n_38735));
	notech_inv i_51676(.A(n_3624), .Z(n_38736));
	notech_inv i_51677(.A(inst_deco2[38]), .Z(n_38737));
	notech_inv i_51678(.A(inst_deco2[39]), .Z(n_38738));
	notech_inv i_51679(.A(n_3623), .Z(n_38739));
	notech_inv i_51680(.A(inst_deco2[40]), .Z(n_38740));
	notech_inv i_51681(.A(inst_deco2[41]), .Z(n_38741));
	notech_inv i_51682(.A(n_3622), .Z(n_38742));
	notech_inv i_51683(.A(inst_deco2[42]), .Z(n_38743));
	notech_inv i_51684(.A(inst_deco2[43]), .Z(n_38744));
	notech_inv i_51685(.A(n_3621), .Z(n_38745));
	notech_inv i_51686(.A(inst_deco2[44]), .Z(n_38746));
	notech_inv i_51687(.A(inst_deco2[45]), .Z(n_38747));
	notech_inv i_51688(.A(n_3620), .Z(n_38748));
	notech_inv i_51689(.A(inst_deco2[46]), .Z(n_38749));
	notech_inv i_51690(.A(inst_deco2[47]), .Z(n_38750));
	notech_inv i_51691(.A(n_3618), .Z(n_38751));
	notech_inv i_51692(.A(inst_deco2[48]), .Z(n_38752));
	notech_inv i_51693(.A(inst_deco2[49]), .Z(n_38753));
	notech_inv i_51694(.A(n_3616), .Z(n_38754));
	notech_inv i_51695(.A(inst_deco2[50]), .Z(n_38755));
	notech_inv i_51696(.A(inst_deco2[51]), .Z(n_38756));
	notech_inv i_51697(.A(n_3615), .Z(n_38757));
	notech_inv i_51698(.A(inst_deco2[52]), .Z(n_38758));
	notech_inv i_51699(.A(inst_deco2[53]), .Z(n_38759));
	notech_inv i_51700(.A(n_3614), .Z(n_38760));
	notech_inv i_51701(.A(inst_deco2[54]), .Z(n_38761));
	notech_inv i_51702(.A(inst_deco2[55]), .Z(n_38762));
	notech_inv i_51703(.A(n_3612), .Z(n_38763));
	notech_inv i_51704(.A(inst_deco2[56]), .Z(n_38764));
	notech_inv i_51705(.A(inst_deco2[57]), .Z(n_38765));
	notech_inv i_51706(.A(n_3611), .Z(n_38766));
	notech_inv i_51707(.A(inst_deco2[58]), .Z(n_38767));
	notech_inv i_51708(.A(inst_deco2[59]), .Z(n_38768));
	notech_inv i_51709(.A(n_3609), .Z(n_38769));
	notech_inv i_51710(.A(inst_deco2[60]), .Z(n_38770));
	notech_inv i_51711(.A(inst_deco2[61]), .Z(n_38771));
	notech_inv i_51712(.A(n_3607), .Z(n_38772));
	notech_inv i_51713(.A(inst_deco2[62]), .Z(n_38773));
	notech_inv i_51714(.A(inst_deco2[63]), .Z(n_38774));
	notech_inv i_51715(.A(n_3606), .Z(n_38775));
	notech_inv i_51716(.A(inst_deco2[64]), .Z(n_38776));
	notech_inv i_51717(.A(inst_deco2[65]), .Z(n_38777));
	notech_inv i_51718(.A(n_3604), .Z(n_38778));
	notech_inv i_51719(.A(inst_deco2[66]), .Z(n_38779));
	notech_inv i_51720(.A(inst_deco2[67]), .Z(n_38780));
	notech_inv i_51721(.A(n_3602), .Z(n_38781));
	notech_inv i_51722(.A(inst_deco2[68]), .Z(n_38782));
	notech_inv i_51723(.A(inst_deco2[69]), .Z(n_38783));
	notech_inv i_51724(.A(n_3600), .Z(n_38784));
	notech_inv i_51725(.A(inst_deco2[70]), .Z(n_38785));
	notech_inv i_51726(.A(inst_deco2[71]), .Z(n_38786));
	notech_inv i_51727(.A(n_3598), .Z(n_38787));
	notech_inv i_51728(.A(inst_deco2[72]), .Z(n_38788));
	notech_inv i_51729(.A(inst_deco2[73]), .Z(n_38789));
	notech_inv i_51730(.A(n_3596), .Z(n_38790));
	notech_inv i_51731(.A(inst_deco2[74]), .Z(n_38791));
	notech_inv i_51732(.A(inst_deco2[75]), .Z(n_38792));
	notech_inv i_51733(.A(n_3594), .Z(n_38793));
	notech_inv i_51734(.A(inst_deco2[76]), .Z(n_38794));
	notech_inv i_51735(.A(inst_deco2[77]), .Z(n_38795));
	notech_inv i_51736(.A(n_3592), .Z(n_38796));
	notech_inv i_51737(.A(inst_deco2[78]), .Z(n_38797));
	notech_inv i_51738(.A(inst_deco2[79]), .Z(n_38798));
	notech_inv i_51739(.A(n_3590), .Z(n_38799));
	notech_inv i_51740(.A(inst_deco2[80]), .Z(n_38800));
	notech_inv i_51741(.A(inst_deco2[81]), .Z(n_38801));
	notech_inv i_51742(.A(n_3588), .Z(n_38802));
	notech_inv i_51743(.A(inst_deco2[82]), .Z(n_38803));
	notech_inv i_51744(.A(inst_deco2[83]), .Z(n_38804));
	notech_inv i_51745(.A(n_3586), .Z(n_38805));
	notech_inv i_51746(.A(inst_deco2[84]), .Z(n_38806));
	notech_inv i_51747(.A(inst_deco2[85]), .Z(n_38807));
	notech_inv i_51748(.A(n_3584), .Z(n_38808));
	notech_inv i_51749(.A(inst_deco2[86]), .Z(n_38809));
	notech_inv i_51750(.A(inst_deco2[87]), .Z(n_38810));
	notech_inv i_51751(.A(n_3582), .Z(n_38811));
	notech_inv i_51752(.A(inst_deco2[88]), .Z(n_38812));
	notech_inv i_51753(.A(inst_deco2[89]), .Z(n_38813));
	notech_inv i_51754(.A(n_3580), .Z(n_38814));
	notech_inv i_51755(.A(inst_deco2[90]), .Z(n_38815));
	notech_inv i_51756(.A(inst_deco2[91]), .Z(n_38816));
	notech_inv i_51757(.A(n_3578), .Z(n_38817));
	notech_inv i_51758(.A(inst_deco2[92]), .Z(n_38818));
	notech_inv i_51759(.A(inst_deco2[93]), .Z(n_38819));
	notech_inv i_51760(.A(n_3576), .Z(n_38820));
	notech_inv i_51761(.A(inst_deco2[94]), .Z(n_38821));
	notech_inv i_51762(.A(inst_deco2[95]), .Z(n_38822));
	notech_inv i_51763(.A(n_3574), .Z(n_38823));
	notech_inv i_51764(.A(inst_deco2[96]), .Z(n_38824));
	notech_inv i_51765(.A(inst_deco2[97]), .Z(n_38825));
	notech_inv i_51766(.A(n_3572), .Z(n_38826));
	notech_inv i_51767(.A(inst_deco2[98]), .Z(n_38827));
	notech_inv i_51768(.A(inst_deco2[99]), .Z(n_38828));
	notech_inv i_51769(.A(n_3570), .Z(n_38829));
	notech_inv i_51770(.A(inst_deco2[100]), .Z(n_38830));
	notech_inv i_51771(.A(inst_deco2[101]), .Z(n_38831));
	notech_inv i_51772(.A(n_3569), .Z(n_38832));
	notech_inv i_51773(.A(inst_deco2[102]), .Z(n_38833));
	notech_inv i_51774(.A(n_42780), .Z(n_38834));
	notech_inv i_51775(.A(inst_deco2[103]), .Z(n_38835));
	notech_inv i_51776(.A(n_3568), .Z(n_38836));
	notech_inv i_51777(.A(inst_deco2[104]), .Z(n_38837));
	notech_inv i_51778(.A(inst_deco2[105]), .Z(n_38838));
	notech_inv i_51779(.A(n_3567), .Z(n_38839));
	notech_inv i_51780(.A(inst_deco2[106]), .Z(n_38840));
	notech_inv i_51781(.A(inst_deco2[107]), .Z(n_38841));
	notech_inv i_51782(.A(n_3566), .Z(n_38842));
	notech_inv i_51783(.A(inst_deco2[108]), .Z(n_38843));
	notech_inv i_51784(.A(inst_deco2[109]), .Z(n_38844));
	notech_inv i_51785(.A(n_3564), .Z(n_38845));
	notech_inv i_51786(.A(inst_deco2[110]), .Z(n_38846));
	notech_inv i_51787(.A(inst_deco2[111]), .Z(n_38847));
	notech_inv i_51788(.A(n_3563), .Z(n_38848));
	notech_inv i_51789(.A(inst_deco2[112]), .Z(n_38849));
	notech_inv i_51790(.A(inst_deco2[113]), .Z(n_38850));
	notech_inv i_51791(.A(n_3562), .Z(n_38851));
	notech_inv i_51792(.A(inst_deco2[114]), .Z(n_38852));
	notech_inv i_51793(.A(inst_deco2[115]), .Z(n_38853));
	notech_inv i_51794(.A(n_3560), .Z(n_38854));
	notech_inv i_51795(.A(inst_deco2[116]), .Z(n_38855));
	notech_inv i_51796(.A(inst_deco2[117]), .Z(n_38856));
	notech_inv i_51797(.A(n_3558), .Z(n_38857));
	notech_inv i_51798(.A(inst_deco2[118]), .Z(n_38858));
	notech_inv i_51799(.A(inst_deco2[119]), .Z(n_38859));
	notech_inv i_51800(.A(n_3556), .Z(n_38860));
	notech_inv i_51801(.A(inst_deco2[120]), .Z(n_38861));
	notech_inv i_51802(.A(inst_deco2[121]), .Z(n_38862));
	notech_inv i_51803(.A(n_3555), .Z(n_38863));
	notech_inv i_51804(.A(inst_deco2[122]), .Z(n_38864));
	notech_inv i_51805(.A(inst_deco2[123]), .Z(n_38865));
	notech_inv i_51806(.A(n_3553), .Z(n_38866));
	notech_inv i_51807(.A(inst_deco2[124]), .Z(n_38867));
	notech_inv i_51808(.A(inst_deco2[125]), .Z(n_38868));
	notech_inv i_51809(.A(n_3551), .Z(n_38869));
	notech_inv i_51810(.A(inst_deco2[126]), .Z(n_38870));
	notech_inv i_51811(.A(inst_deco2[127]), .Z(n_38871));
	notech_inv i_51812(.A(n_3550), .Z(n_38872));
	notech_inv i_51813(.A(inst_deco1[0]), .Z(n_38873));
	notech_inv i_51814(.A(n_3549), .Z(n_38874));
	notech_inv i_51815(.A(inst_deco1[1]), .Z(n_38875));
	notech_inv i_51816(.A(n_3548), .Z(n_38876));
	notech_inv i_51817(.A(inst_deco1[2]), .Z(n_38877));
	notech_inv i_51818(.A(n_3546), .Z(n_38878));
	notech_inv i_51819(.A(inst_deco1[3]), .Z(n_38879));
	notech_inv i_51820(.A(n_3544), .Z(n_38880));
	notech_inv i_51821(.A(n_3542), .Z(n_38881));
	notech_inv i_51822(.A(inst_deco1[5]), .Z(n_38882));
	notech_inv i_51823(.A(n_3540), .Z(n_38883));
	notech_inv i_51824(.A(inst_deco1[6]), .Z(n_38884));
	notech_inv i_51825(.A(n_3538), .Z(n_38885));
	notech_inv i_51826(.A(inst_deco1[7]), .Z(n_38886));
	notech_inv i_51827(.A(n_3536), .Z(n_38887));
	notech_inv i_51828(.A(inst_deco1[8]), .Z(n_38888));
	notech_inv i_51829(.A(n_3534), .Z(n_38889));
	notech_inv i_51830(.A(inst_deco1[9]), .Z(n_38890));
	notech_inv i_51831(.A(n_3532), .Z(n_38891));
	notech_inv i_51832(.A(inst_deco1[10]), .Z(n_38892));
	notech_inv i_51833(.A(n_3530), .Z(n_38893));
	notech_inv i_51834(.A(inst_deco1[11]), .Z(n_38894));
	notech_inv i_51835(.A(n_3528), .Z(n_38895));
	notech_inv i_51836(.A(inst_deco1[12]), .Z(n_38896));
	notech_inv i_51837(.A(n_3526), .Z(n_38897));
	notech_inv i_51838(.A(n_3524), .Z(n_38898));
	notech_inv i_51839(.A(inst_deco1[14]), .Z(n_38899));
	notech_inv i_51840(.A(n_3522), .Z(n_38900));
	notech_inv i_51841(.A(inst_deco1[15]), .Z(n_38901));
	notech_inv i_51842(.A(n_3520), .Z(n_38902));
	notech_inv i_51843(.A(inst_deco1[16]), .Z(n_38903));
	notech_inv i_51844(.A(n_3518), .Z(n_38904));
	notech_inv i_51845(.A(inst_deco1[17]), .Z(n_38905));
	notech_inv i_51846(.A(n_3516), .Z(n_38906));
	notech_inv i_51847(.A(inst_deco1[18]), .Z(n_38907));
	notech_inv i_51848(.A(n_3514), .Z(n_38908));
	notech_inv i_51849(.A(inst_deco1[19]), .Z(n_38909));
	notech_inv i_51850(.A(n_3512), .Z(n_38910));
	notech_inv i_51851(.A(inst_deco1[20]), .Z(n_38911));
	notech_inv i_51852(.A(n_3510), .Z(n_38912));
	notech_inv i_51853(.A(inst_deco1[21]), .Z(n_38913));
	notech_inv i_51854(.A(n_3509), .Z(n_38914));
	notech_inv i_51855(.A(inst_deco1[22]), .Z(n_38915));
	notech_inv i_51856(.A(n_3508), .Z(n_38916));
	notech_inv i_51857(.A(inst_deco1[23]), .Z(n_38917));
	notech_inv i_51858(.A(n_3507), .Z(n_38918));
	notech_inv i_51859(.A(inst_deco1[24]), .Z(n_38919));
	notech_inv i_51860(.A(n_3506), .Z(n_38920));
	notech_inv i_51861(.A(inst_deco1[25]), .Z(n_38921));
	notech_inv i_51862(.A(n_3505), .Z(n_38922));
	notech_inv i_51863(.A(inst_deco1[26]), .Z(n_38923));
	notech_inv i_51864(.A(n_3504), .Z(n_38924));
	notech_inv i_51865(.A(inst_deco1[27]), .Z(n_38925));
	notech_inv i_51866(.A(n_3503), .Z(n_38926));
	notech_inv i_51867(.A(inst_deco1[28]), .Z(n_38927));
	notech_inv i_51868(.A(n_3502), .Z(n_38928));
	notech_inv i_51869(.A(inst_deco1[29]), .Z(n_38929));
	notech_inv i_51870(.A(n_3501), .Z(n_38930));
	notech_inv i_51871(.A(inst_deco1[30]), .Z(n_38931));
	notech_inv i_51872(.A(n_3500), .Z(n_38932));
	notech_inv i_51873(.A(inst_deco1[31]), .Z(n_38933));
	notech_inv i_51874(.A(n_3499), .Z(n_38934));
	notech_inv i_51875(.A(inst_deco1[32]), .Z(n_38935));
	notech_inv i_51876(.A(n_3498), .Z(n_38936));
	notech_inv i_51877(.A(inst_deco1[33]), .Z(n_38937));
	notech_inv i_51878(.A(n_3497), .Z(n_38938));
	notech_inv i_51879(.A(inst_deco1[34]), .Z(n_38939));
	notech_inv i_51880(.A(n_3496), .Z(n_38940));
	notech_inv i_51881(.A(inst_deco1[35]), .Z(n_38941));
	notech_inv i_51882(.A(n_3495), .Z(n_38942));
	notech_inv i_51883(.A(inst_deco1[36]), .Z(n_38943));
	notech_inv i_51884(.A(n_3494), .Z(n_38944));
	notech_inv i_51885(.A(inst_deco1[37]), .Z(n_38945));
	notech_inv i_51886(.A(n_3493), .Z(n_38946));
	notech_inv i_51887(.A(inst_deco1[38]), .Z(n_38947));
	notech_inv i_51888(.A(n_3491), .Z(n_38948));
	notech_inv i_51889(.A(inst_deco1[39]), .Z(n_38949));
	notech_inv i_51890(.A(n_3489), .Z(n_38950));
	notech_inv i_51891(.A(inst_deco1[40]), .Z(n_38951));
	notech_inv i_51892(.A(n_3487), .Z(n_38952));
	notech_inv i_51893(.A(inst_deco1[41]), .Z(n_38953));
	notech_inv i_51894(.A(n_3486), .Z(n_38954));
	notech_inv i_51895(.A(inst_deco1[42]), .Z(n_38955));
	notech_inv i_51896(.A(n_3484), .Z(n_38956));
	notech_inv i_51897(.A(inst_deco1[43]), .Z(n_38957));
	notech_inv i_51898(.A(n_3482), .Z(n_38958));
	notech_inv i_51899(.A(inst_deco1[44]), .Z(n_38959));
	notech_inv i_51900(.A(n_3480), .Z(n_38960));
	notech_inv i_51901(.A(inst_deco1[45]), .Z(n_38961));
	notech_inv i_51902(.A(n_3478), .Z(n_38962));
	notech_inv i_51903(.A(inst_deco1[46]), .Z(n_38963));
	notech_inv i_51904(.A(n_3476), .Z(n_38964));
	notech_inv i_51905(.A(inst_deco1[47]), .Z(n_38965));
	notech_inv i_51906(.A(n_3474), .Z(n_38966));
	notech_inv i_51907(.A(inst_deco1[48]), .Z(n_38967));
	notech_inv i_51908(.A(n_3472), .Z(n_38968));
	notech_inv i_51909(.A(inst_deco1[49]), .Z(n_38969));
	notech_inv i_51910(.A(n_3470), .Z(n_38970));
	notech_inv i_51911(.A(inst_deco1[50]), .Z(n_38971));
	notech_inv i_51912(.A(n_3468), .Z(n_38972));
	notech_inv i_51913(.A(inst_deco1[51]), .Z(n_38973));
	notech_inv i_51914(.A(n_3466), .Z(n_38974));
	notech_inv i_51915(.A(inst_deco1[52]), .Z(n_38975));
	notech_inv i_51916(.A(n_3464), .Z(n_38976));
	notech_inv i_51917(.A(inst_deco1[53]), .Z(n_38977));
	notech_inv i_51918(.A(n_3462), .Z(n_38978));
	notech_inv i_51919(.A(inst_deco1[54]), .Z(n_38979));
	notech_inv i_51920(.A(n_3460), .Z(n_38980));
	notech_inv i_51921(.A(inst_deco1[55]), .Z(n_38981));
	notech_inv i_51922(.A(n_3458), .Z(n_38982));
	notech_inv i_51923(.A(inst_deco1[56]), .Z(n_38983));
	notech_inv i_51924(.A(n_3456), .Z(n_38984));
	notech_inv i_51925(.A(inst_deco1[57]), .Z(n_38985));
	notech_inv i_51926(.A(n_3454), .Z(n_38986));
	notech_inv i_51927(.A(inst_deco1[58]), .Z(n_38987));
	notech_inv i_51928(.A(n_3452), .Z(n_38988));
	notech_inv i_51929(.A(inst_deco1[59]), .Z(n_38989));
	notech_inv i_51930(.A(n_3450), .Z(n_38990));
	notech_inv i_51931(.A(inst_deco1[60]), .Z(n_38991));
	notech_inv i_51932(.A(n_3448), .Z(n_38992));
	notech_inv i_51933(.A(inst_deco1[61]), .Z(n_38993));
	notech_inv i_51934(.A(n_3446), .Z(n_38994));
	notech_inv i_51935(.A(inst_deco1[62]), .Z(n_38995));
	notech_inv i_51936(.A(n_3444), .Z(n_38996));
	notech_inv i_51937(.A(inst_deco1[63]), .Z(n_38997));
	notech_inv i_51938(.A(n_3442), .Z(n_38998));
	notech_inv i_51939(.A(inst_deco1[64]), .Z(n_38999));
	notech_inv i_51940(.A(n_3440), .Z(n_39000));
	notech_inv i_51941(.A(inst_deco1[65]), .Z(n_39001));
	notech_inv i_51942(.A(n_3438), .Z(n_39002));
	notech_inv i_51943(.A(inst_deco1[66]), .Z(n_39003));
	notech_inv i_51944(.A(n_3436), .Z(n_39004));
	notech_inv i_51945(.A(inst_deco1[67]), .Z(n_39005));
	notech_inv i_51946(.A(n_3434), .Z(n_39006));
	notech_inv i_51947(.A(inst_deco1[68]), .Z(n_39007));
	notech_inv i_51948(.A(n_3432), .Z(n_39008));
	notech_inv i_51949(.A(inst_deco1[69]), .Z(n_39009));
	notech_inv i_51950(.A(n_3430), .Z(n_39010));
	notech_inv i_51951(.A(inst_deco1[70]), .Z(n_39011));
	notech_inv i_51952(.A(n_3428), .Z(n_39012));
	notech_inv i_51953(.A(inst_deco1[71]), .Z(n_39013));
	notech_inv i_51954(.A(n_3426), .Z(n_39014));
	notech_inv i_51955(.A(inst_deco1[72]), .Z(n_39015));
	notech_inv i_51956(.A(n_3424), .Z(n_39016));
	notech_inv i_51957(.A(inst_deco1[73]), .Z(n_39017));
	notech_inv i_51958(.A(n_3422), .Z(n_39018));
	notech_inv i_51959(.A(inst_deco1[74]), .Z(n_39019));
	notech_inv i_51960(.A(n_3420), .Z(n_39020));
	notech_inv i_51961(.A(inst_deco1[75]), .Z(n_39021));
	notech_inv i_51962(.A(n_3418), .Z(n_39022));
	notech_inv i_51963(.A(inst_deco1[76]), .Z(n_39023));
	notech_inv i_51964(.A(n_3416), .Z(n_39024));
	notech_inv i_51965(.A(inst_deco1[77]), .Z(n_39025));
	notech_inv i_51966(.A(n_3414), .Z(n_39026));
	notech_inv i_51967(.A(inst_deco1[78]), .Z(n_39027));
	notech_inv i_51968(.A(n_3412), .Z(n_39028));
	notech_inv i_51969(.A(inst_deco1[79]), .Z(n_39029));
	notech_inv i_51970(.A(n_3410), .Z(n_39030));
	notech_inv i_51971(.A(n_3408), .Z(n_39031));
	notech_inv i_51972(.A(n_3406), .Z(n_39032));
	notech_inv i_51973(.A(n_3404), .Z(n_39033));
	notech_inv i_51974(.A(n_3402), .Z(n_39034));
	notech_inv i_51975(.A(n_3400), .Z(n_39035));
	notech_inv i_51976(.A(n_3398), .Z(n_39036));
	notech_inv i_51977(.A(n_3396), .Z(n_39037));
	notech_inv i_51978(.A(n_3394), .Z(n_39038));
	notech_inv i_51979(.A(inst_deco1[88]), .Z(n_39039));
	notech_inv i_51980(.A(n_3392), .Z(n_39040));
	notech_inv i_51981(.A(inst_deco1[89]), .Z(n_39041));
	notech_inv i_51982(.A(n_3390), .Z(n_39042));
	notech_inv i_51983(.A(inst_deco1[90]), .Z(n_39043));
	notech_inv i_51984(.A(n_3388), .Z(n_39044));
	notech_inv i_51985(.A(inst_deco1[91]), .Z(n_39045));
	notech_inv i_51986(.A(n_3386), .Z(n_39046));
	notech_inv i_51987(.A(inst_deco1[92]), .Z(n_39047));
	notech_inv i_51988(.A(n_3384), .Z(n_39048));
	notech_inv i_51989(.A(inst_deco1[93]), .Z(n_39049));
	notech_inv i_51990(.A(n_3382), .Z(n_39050));
	notech_inv i_51991(.A(inst_deco1[94]), .Z(n_39051));
	notech_inv i_51992(.A(n_3380), .Z(n_39052));
	notech_inv i_51993(.A(inst_deco1[95]), .Z(n_39053));
	notech_inv i_51994(.A(n_3378), .Z(n_39054));
	notech_inv i_51995(.A(inst_deco1[96]), .Z(n_39055));
	notech_inv i_51996(.A(n_3376), .Z(n_39056));
	notech_inv i_51997(.A(inst_deco1[97]), .Z(n_39057));
	notech_inv i_51998(.A(n_3374), .Z(n_39058));
	notech_inv i_51999(.A(inst_deco1[98]), .Z(n_39059));
	notech_inv i_52000(.A(n_3372), .Z(n_39060));
	notech_inv i_52001(.A(inst_deco1[99]), .Z(n_39061));
	notech_inv i_52002(.A(n_3370), .Z(n_39062));
	notech_inv i_52003(.A(inst_deco1[100]), .Z(n_39063));
	notech_inv i_52004(.A(n_3368), .Z(n_39064));
	notech_inv i_52005(.A(inst_deco1[101]), .Z(n_39065));
	notech_inv i_52006(.A(n_3366), .Z(n_39066));
	notech_inv i_52007(.A(inst_deco1[102]), .Z(n_39067));
	notech_inv i_52008(.A(n_3364), .Z(n_39068));
	notech_inv i_52009(.A(n_50550), .Z(n_39069));
	notech_inv i_52010(.A(inst_deco1[103]), .Z(n_39070));
	notech_inv i_52011(.A(n_3362), .Z(n_39071));
	notech_inv i_52012(.A(inst_deco1[104]), .Z(n_39072));
	notech_inv i_52013(.A(n_3360), .Z(n_39073));
	notech_inv i_52014(.A(inst_deco1[105]), .Z(n_39074));
	notech_inv i_52015(.A(n_3358), .Z(n_39075));
	notech_inv i_52016(.A(n_3356), .Z(n_39076));
	notech_inv i_52017(.A(inst_deco1[107]), .Z(n_39077));
	notech_inv i_52018(.A(n_3354), .Z(n_39078));
	notech_inv i_52019(.A(inst_deco1[108]), .Z(n_39079));
	notech_inv i_52020(.A(n_3352), .Z(n_39080));
	notech_inv i_52021(.A(inst_deco1[109]), .Z(n_39081));
	notech_inv i_52022(.A(n_3350), .Z(n_39082));
	notech_inv i_52023(.A(inst_deco1[110]), .Z(n_39083));
	notech_inv i_52024(.A(n_3348), .Z(n_39084));
	notech_inv i_52025(.A(inst_deco1[111]), .Z(n_39085));
	notech_inv i_52026(.A(n_3346), .Z(n_39086));
	notech_inv i_52027(.A(inst_deco1[112]), .Z(n_39087));
	notech_inv i_52028(.A(n_3344), .Z(n_39088));
	notech_inv i_52029(.A(n_3342), .Z(n_39089));
	notech_inv i_52030(.A(inst_deco1[114]), .Z(n_39090));
	notech_inv i_52031(.A(n_3340), .Z(n_39091));
	notech_inv i_52032(.A(inst_deco1[115]), .Z(n_39092));
	notech_inv i_52033(.A(n_3338), .Z(n_39093));
	notech_inv i_52034(.A(inst_deco1[116]), .Z(n_39094));
	notech_inv i_52035(.A(n_3336), .Z(n_39095));
	notech_inv i_52036(.A(inst_deco1[117]), .Z(n_39096));
	notech_inv i_52037(.A(n_3334), .Z(n_39097));
	notech_inv i_52038(.A(inst_deco1[118]), .Z(n_39098));
	notech_inv i_52039(.A(n_3332), .Z(n_39099));
	notech_inv i_52040(.A(inst_deco1[119]), .Z(n_39100));
	notech_inv i_52041(.A(n_3330), .Z(n_39101));
	notech_inv i_52042(.A(inst_deco1[120]), .Z(n_39102));
	notech_inv i_52043(.A(n_3328), .Z(n_39103));
	notech_inv i_52044(.A(inst_deco1[121]), .Z(n_39104));
	notech_inv i_52045(.A(n_3326), .Z(n_39105));
	notech_inv i_52046(.A(inst_deco1[122]), .Z(n_39106));
	notech_inv i_52047(.A(n_3324), .Z(n_39107));
	notech_inv i_52048(.A(inst_deco1[123]), .Z(n_39108));
	notech_inv i_52049(.A(n_3322), .Z(n_39109));
	notech_inv i_52050(.A(inst_deco1[124]), .Z(n_39110));
	notech_inv i_52051(.A(n_3320), .Z(n_39111));
	notech_inv i_52052(.A(inst_deco1[125]), .Z(n_39112));
	notech_inv i_52053(.A(n_3319), .Z(n_39113));
	notech_inv i_52054(.A(inst_deco1[126]), .Z(n_39114));
	notech_inv i_52055(.A(n_3318), .Z(n_39115));
	notech_inv i_52056(.A(inst_deco1[127]), .Z(n_39116));
	notech_inv i_52057(.A(n_41571), .Z(n_39117));
	notech_inv i_52058(.A(overgs), .Z(n_39118));
	notech_inv i_52059(.A(n_3316), .Z(n_39119));
	notech_inv i_52060(.A(\over_seg2[5] ), .Z(n_39120));
	notech_inv i_52061(.A(n_3315), .Z(n_39121));
	notech_inv i_52062(.A(\over_seg1[5] ), .Z(n_39122));
	notech_inv i_52063(.A(n_3314), .Z(n_39123));
	notech_inv i_52064(.A(to_acu2[0]), .Z(n_39124));
	notech_inv i_52065(.A(to_acu2[1]), .Z(n_39125));
	notech_inv i_52066(.A(n_3312), .Z(n_39126));
	notech_inv i_52067(.A(to_acu2[2]), .Z(n_39127));
	notech_inv i_52068(.A(to_acu2[3]), .Z(n_39128));
	notech_inv i_52069(.A(n_3311), .Z(n_39129));
	notech_inv i_52070(.A(to_acu2[4]), .Z(n_39130));
	notech_inv i_52071(.A(to_acu2[5]), .Z(n_39131));
	notech_inv i_52072(.A(n_3310), .Z(n_39132));
	notech_inv i_52073(.A(to_acu2[6]), .Z(n_39133));
	notech_inv i_52074(.A(to_acu2[7]), .Z(n_39134));
	notech_inv i_52075(.A(n_3309), .Z(n_39135));
	notech_inv i_52076(.A(to_acu2[8]), .Z(n_39136));
	notech_inv i_52077(.A(to_acu2[9]), .Z(n_39137));
	notech_inv i_52078(.A(n_3308), .Z(n_39138));
	notech_inv i_52079(.A(to_acu2[10]), .Z(n_39139));
	notech_inv i_52080(.A(to_acu2[11]), .Z(n_39140));
	notech_inv i_52081(.A(n_3306), .Z(n_39141));
	notech_inv i_52082(.A(to_acu2[12]), .Z(n_39142));
	notech_inv i_52083(.A(to_acu2[13]), .Z(n_39143));
	notech_inv i_52084(.A(n_3305), .Z(n_39144));
	notech_inv i_52085(.A(to_acu2[14]), .Z(n_39145));
	notech_inv i_52086(.A(to_acu2[15]), .Z(n_39146));
	notech_inv i_52087(.A(n_3303), .Z(n_39147));
	notech_inv i_52088(.A(to_acu2[16]), .Z(n_39148));
	notech_inv i_52089(.A(to_acu2[17]), .Z(n_39149));
	notech_inv i_52090(.A(n_3302), .Z(n_39150));
	notech_inv i_52091(.A(to_acu2[18]), .Z(n_39151));
	notech_inv i_52092(.A(to_acu2[19]), .Z(n_39152));
	notech_inv i_52093(.A(n_3301), .Z(n_39153));
	notech_inv i_52094(.A(to_acu2[20]), .Z(n_39154));
	notech_inv i_52095(.A(to_acu2[21]), .Z(n_39155));
	notech_inv i_52096(.A(n_3300), .Z(n_39156));
	notech_inv i_52097(.A(to_acu2[22]), .Z(n_39157));
	notech_inv i_52098(.A(to_acu2[23]), .Z(n_39158));
	notech_inv i_52099(.A(n_3299), .Z(n_39159));
	notech_inv i_52100(.A(to_acu2[24]), .Z(n_39160));
	notech_inv i_52101(.A(to_acu2[25]), .Z(n_39161));
	notech_inv i_52102(.A(n_3298), .Z(n_39162));
	notech_inv i_52103(.A(to_acu2[26]), .Z(n_39163));
	notech_inv i_52104(.A(to_acu2[27]), .Z(n_39164));
	notech_inv i_52105(.A(n_3297), .Z(n_39165));
	notech_inv i_52106(.A(to_acu2[28]), .Z(n_39166));
	notech_inv i_52107(.A(to_acu2[29]), .Z(n_39167));
	notech_inv i_52108(.A(n_3296), .Z(n_39168));
	notech_inv i_52109(.A(to_acu2[30]), .Z(n_39169));
	notech_inv i_52110(.A(to_acu2[31]), .Z(n_39170));
	notech_inv i_52111(.A(n_3295), .Z(n_39171));
	notech_inv i_52112(.A(to_acu2[32]), .Z(n_39172));
	notech_inv i_52113(.A(to_acu2[33]), .Z(n_39173));
	notech_inv i_52114(.A(n_3294), .Z(n_39174));
	notech_inv i_52115(.A(to_acu2[34]), .Z(n_39175));
	notech_inv i_52116(.A(to_acu2[35]), .Z(n_39176));
	notech_inv i_52117(.A(n_3293), .Z(n_39177));
	notech_inv i_52118(.A(to_acu2[36]), .Z(n_39178));
	notech_inv i_52119(.A(to_acu2[37]), .Z(n_39179));
	notech_inv i_52120(.A(n_3292), .Z(n_39180));
	notech_inv i_52121(.A(to_acu2[38]), .Z(n_39181));
	notech_inv i_52122(.A(n_3291), .Z(n_39182));
	notech_inv i_52123(.A(to_acu2[40]), .Z(n_39183));
	notech_inv i_52124(.A(to_acu2[41]), .Z(n_39184));
	notech_inv i_52125(.A(n_3290), .Z(n_39185));
	notech_inv i_52126(.A(to_acu2[42]), .Z(n_39186));
	notech_inv i_52127(.A(to_acu2[43]), .Z(n_39187));
	notech_inv i_52128(.A(n_3289), .Z(n_39188));
	notech_inv i_52129(.A(to_acu2[44]), .Z(n_39189));
	notech_inv i_52130(.A(to_acu2[45]), .Z(n_39190));
	notech_inv i_52131(.A(n_3288), .Z(n_39191));
	notech_inv i_52132(.A(to_acu2[46]), .Z(n_39192));
	notech_inv i_52133(.A(to_acu2[47]), .Z(n_39193));
	notech_inv i_52134(.A(n_3287), .Z(n_39194));
	notech_inv i_52135(.A(to_acu2[48]), .Z(n_39195));
	notech_inv i_52136(.A(to_acu2[49]), .Z(n_39196));
	notech_inv i_52137(.A(n_3286), .Z(n_39197));
	notech_inv i_52138(.A(to_acu2[50]), .Z(n_39198));
	notech_inv i_52139(.A(to_acu2[51]), .Z(n_39199));
	notech_inv i_52140(.A(n_3285), .Z(n_39200));
	notech_inv i_52141(.A(to_acu2[52]), .Z(n_39201));
	notech_inv i_52142(.A(to_acu2[53]), .Z(n_39202));
	notech_inv i_52143(.A(n_3284), .Z(n_39203));
	notech_inv i_52144(.A(to_acu2[54]), .Z(n_39204));
	notech_inv i_52145(.A(to_acu2[55]), .Z(n_39205));
	notech_inv i_52146(.A(n_3283), .Z(n_39206));
	notech_inv i_52147(.A(to_acu2[56]), .Z(n_39207));
	notech_inv i_52148(.A(to_acu2[57]), .Z(n_39208));
	notech_inv i_52149(.A(n_3282), .Z(n_39209));
	notech_inv i_52150(.A(to_acu2[58]), .Z(n_39210));
	notech_inv i_52151(.A(to_acu2[59]), .Z(n_39211));
	notech_inv i_52152(.A(n_3281), .Z(n_39212));
	notech_inv i_52153(.A(to_acu2[60]), .Z(n_39213));
	notech_inv i_52154(.A(to_acu2[61]), .Z(n_39214));
	notech_inv i_52155(.A(n_3280), .Z(n_39215));
	notech_inv i_52156(.A(to_acu2[62]), .Z(n_39216));
	notech_inv i_52157(.A(to_acu2[63]), .Z(n_39217));
	notech_inv i_52158(.A(n_3279), .Z(n_39218));
	notech_inv i_52159(.A(to_acu2[64]), .Z(n_39219));
	notech_inv i_52160(.A(to_acu2[65]), .Z(n_39220));
	notech_inv i_52161(.A(n_3278), .Z(n_39221));
	notech_inv i_52162(.A(to_acu2[66]), .Z(n_39222));
	notech_inv i_52163(.A(to_acu2[67]), .Z(n_39223));
	notech_inv i_52164(.A(n_3277), .Z(n_39224));
	notech_inv i_52165(.A(to_acu2[68]), .Z(n_39225));
	notech_inv i_52166(.A(to_acu2[69]), .Z(n_39226));
	notech_inv i_52167(.A(n_3276), .Z(n_39227));
	notech_inv i_52168(.A(to_acu2[70]), .Z(n_39228));
	notech_inv i_52169(.A(to_acu2[71]), .Z(n_39229));
	notech_inv i_52170(.A(n_3275), .Z(n_39230));
	notech_inv i_52171(.A(to_acu2[72]), .Z(n_39231));
	notech_inv i_52172(.A(to_acu2[73]), .Z(n_39232));
	notech_inv i_52173(.A(n_3274), .Z(n_39233));
	notech_inv i_52174(.A(to_acu2[74]), .Z(n_39234));
	notech_inv i_52175(.A(to_acu2[75]), .Z(n_39235));
	notech_inv i_52176(.A(n_3273), .Z(n_39236));
	notech_inv i_52177(.A(to_acu2[76]), .Z(n_39237));
	notech_inv i_52178(.A(to_acu2[77]), .Z(n_39238));
	notech_inv i_52179(.A(n_3272), .Z(n_39239));
	notech_inv i_52180(.A(to_acu2[78]), .Z(n_39240));
	notech_inv i_52181(.A(to_acu2[79]), .Z(n_39241));
	notech_inv i_52182(.A(n_3271), .Z(n_39242));
	notech_inv i_52183(.A(to_acu2[80]), .Z(n_39243));
	notech_inv i_52184(.A(to_acu2[81]), .Z(n_39244));
	notech_inv i_52185(.A(n_3270), .Z(n_39245));
	notech_inv i_52186(.A(to_acu2[82]), .Z(n_39246));
	notech_inv i_52187(.A(to_acu2[83]), .Z(n_39247));
	notech_inv i_52188(.A(n_3269), .Z(n_39248));
	notech_inv i_52189(.A(n_47603), .Z(n_39249));
	notech_inv i_52190(.A(to_acu2[84]), .Z(n_39250));
	notech_inv i_52191(.A(to_acu2[85]), .Z(n_39251));
	notech_inv i_52192(.A(n_3268), .Z(n_39252));
	notech_inv i_52193(.A(to_acu2[86]), .Z(n_39253));
	notech_inv i_52194(.A(to_acu2[87]), .Z(n_39254));
	notech_inv i_52195(.A(n_3267), .Z(n_39255));
	notech_inv i_52196(.A(to_acu2[88]), .Z(n_39256));
	notech_inv i_52197(.A(to_acu2[89]), .Z(n_39257));
	notech_inv i_52198(.A(n_3266), .Z(n_39258));
	notech_inv i_52199(.A(to_acu2[90]), .Z(n_39259));
	notech_inv i_52200(.A(to_acu2[91]), .Z(n_39260));
	notech_inv i_52201(.A(n_3265), .Z(n_39261));
	notech_inv i_52202(.A(to_acu2[92]), .Z(n_39262));
	notech_inv i_52203(.A(to_acu2[93]), .Z(n_39263));
	notech_inv i_52204(.A(n_3264), .Z(n_39264));
	notech_inv i_52205(.A(to_acu2[94]), .Z(n_39265));
	notech_inv i_52206(.A(to_acu2[95]), .Z(n_39266));
	notech_inv i_52207(.A(n_3263), .Z(n_39267));
	notech_inv i_52208(.A(to_acu2[96]), .Z(n_39268));
	notech_inv i_52209(.A(to_acu2[97]), .Z(n_39269));
	notech_inv i_52210(.A(n_3262), .Z(n_39270));
	notech_inv i_52211(.A(to_acu2[98]), .Z(n_39271));
	notech_inv i_52212(.A(to_acu2[99]), .Z(n_39272));
	notech_inv i_52213(.A(n_3261), .Z(n_39273));
	notech_inv i_52214(.A(to_acu2[100]), .Z(n_39274));
	notech_inv i_52215(.A(to_acu2[101]), .Z(n_39275));
	notech_inv i_52216(.A(n_3260), .Z(n_39276));
	notech_inv i_52217(.A(to_acu2[102]), .Z(n_39277));
	notech_inv i_52218(.A(to_acu2[103]), .Z(n_39278));
	notech_inv i_52219(.A(n_3259), .Z(n_39279));
	notech_inv i_52220(.A(to_acu2[104]), .Z(n_39280));
	notech_inv i_52221(.A(to_acu2[105]), .Z(n_39281));
	notech_inv i_52222(.A(n_3258), .Z(n_39282));
	notech_inv i_52223(.A(to_acu2[106]), .Z(n_39283));
	notech_inv i_52224(.A(to_acu2[107]), .Z(n_39284));
	notech_inv i_52225(.A(n_3257), .Z(n_39285));
	notech_inv i_52226(.A(to_acu2[108]), .Z(n_39286));
	notech_inv i_52227(.A(to_acu2[109]), .Z(n_39287));
	notech_inv i_52228(.A(n_3256), .Z(n_39288));
	notech_inv i_52229(.A(to_acu2[110]), .Z(n_39289));
	notech_inv i_52230(.A(to_acu2[111]), .Z(n_39290));
	notech_inv i_52231(.A(n_3255), .Z(n_39291));
	notech_inv i_52232(.A(to_acu2[112]), .Z(n_39292));
	notech_inv i_52233(.A(to_acu2[113]), .Z(n_39293));
	notech_inv i_52234(.A(n_3254), .Z(n_39294));
	notech_inv i_52235(.A(to_acu2[114]), .Z(n_39295));
	notech_inv i_52236(.A(to_acu2[115]), .Z(n_39296));
	notech_inv i_52237(.A(n_3253), .Z(n_39297));
	notech_inv i_52238(.A(to_acu2[116]), .Z(n_39298));
	notech_inv i_52239(.A(to_acu2[117]), .Z(n_39299));
	notech_inv i_52240(.A(n_3252), .Z(n_39300));
	notech_inv i_52241(.A(to_acu2[118]), .Z(n_39301));
	notech_inv i_52242(.A(to_acu2[119]), .Z(n_39302));
	notech_inv i_52243(.A(n_3251), .Z(n_39303));
	notech_inv i_52244(.A(to_acu2[120]), .Z(n_39304));
	notech_inv i_52245(.A(to_acu2[121]), .Z(n_39305));
	notech_inv i_52246(.A(to_acu2[122]), .Z(n_39306));
	notech_inv i_52247(.A(to_acu2[123]), .Z(n_39307));
	notech_inv i_52248(.A(to_acu2[124]), .Z(n_39308));
	notech_inv i_52249(.A(to_acu2[125]), .Z(n_39309));
	notech_inv i_52250(.A(n_3245), .Z(n_39310));
	notech_inv i_52251(.A(to_acu2[126]), .Z(n_39311));
	notech_inv i_52252(.A(to_acu2[127]), .Z(n_39312));
	notech_inv i_52253(.A(n_3243), .Z(n_39313));
	notech_inv i_52254(.A(to_acu2[128]), .Z(n_39314));
	notech_inv i_52255(.A(to_acu2[129]), .Z(n_39315));
	notech_inv i_52256(.A(n_3241), .Z(n_39316));
	notech_inv i_52257(.A(to_acu2[130]), .Z(n_39317));
	notech_inv i_52258(.A(to_acu2[131]), .Z(n_39318));
	notech_inv i_52259(.A(n_3240), .Z(n_39319));
	notech_inv i_52260(.A(to_acu2[132]), .Z(n_39320));
	notech_inv i_52261(.A(to_acu2[133]), .Z(n_39321));
	notech_inv i_52262(.A(n_3238), .Z(n_39322));
	notech_inv i_52263(.A(to_acu2[134]), .Z(n_39323));
	notech_inv i_52264(.A(to_acu2[135]), .Z(n_39324));
	notech_inv i_52265(.A(n_3236), .Z(n_39325));
	notech_inv i_52266(.A(to_acu2[136]), .Z(n_39326));
	notech_inv i_52267(.A(to_acu2[137]), .Z(n_39327));
	notech_inv i_52268(.A(to_acu2[138]), .Z(n_39328));
	notech_inv i_52269(.A(to_acu2[139]), .Z(n_39329));
	notech_inv i_52270(.A(to_acu2[140]), .Z(n_39330));
	notech_inv i_52271(.A(to_acu2[141]), .Z(n_39331));
	notech_inv i_52272(.A(to_acu2[142]), .Z(n_39332));
	notech_inv i_52273(.A(to_acu2[143]), .Z(n_39333));
	notech_inv i_52274(.A(to_acu2[144]), .Z(n_39334));
	notech_inv i_52275(.A(to_acu2[145]), .Z(n_39335));
	notech_inv i_52276(.A(to_acu2[146]), .Z(n_39336));
	notech_inv i_52277(.A(to_acu2[147]), .Z(n_39337));
	notech_inv i_52278(.A(to_acu2[148]), .Z(n_39338));
	notech_inv i_52279(.A(to_acu2[149]), .Z(n_39339));
	notech_inv i_52280(.A(to_acu2[150]), .Z(n_39340));
	notech_inv i_52281(.A(to_acu2[151]), .Z(n_39341));
	notech_inv i_52282(.A(to_acu2[152]), .Z(n_39342));
	notech_inv i_52283(.A(to_acu2[153]), .Z(n_39343));
	notech_inv i_52284(.A(to_acu2[154]), .Z(n_39344));
	notech_inv i_52285(.A(to_acu2[155]), .Z(n_39345));
	notech_inv i_52286(.A(to_acu2[156]), .Z(n_39346));
	notech_inv i_52287(.A(to_acu2[157]), .Z(n_39347));
	notech_inv i_52288(.A(to_acu2[158]), .Z(n_39348));
	notech_inv i_52289(.A(to_acu2[159]), .Z(n_39349));
	notech_inv i_52290(.A(to_acu2[160]), .Z(n_39350));
	notech_inv i_52291(.A(to_acu2[161]), .Z(n_39351));
	notech_inv i_52292(.A(to_acu2[162]), .Z(n_39352));
	notech_inv i_52293(.A(to_acu2[163]), .Z(n_39353));
	notech_inv i_52294(.A(to_acu2[164]), .Z(n_39354));
	notech_inv i_52295(.A(to_acu2[165]), .Z(n_39355));
	notech_inv i_52296(.A(to_acu2[166]), .Z(n_39356));
	notech_inv i_52297(.A(to_acu2[167]), .Z(n_39357));
	notech_inv i_52298(.A(n_3205), .Z(n_39358));
	notech_inv i_52299(.A(to_acu2[168]), .Z(n_39359));
	notech_inv i_52300(.A(to_acu2[169]), .Z(n_39360));
	notech_inv i_52301(.A(to_acu2[170]), .Z(n_39361));
	notech_inv i_52302(.A(n_3202), .Z(n_39362));
	notech_inv i_52303(.A(to_acu2[171]), .Z(n_39363));
	notech_inv i_52304(.A(to_acu2[172]), .Z(n_39364));
	notech_inv i_52305(.A(n_3200), .Z(n_39365));
	notech_inv i_52306(.A(to_acu2[173]), .Z(n_39366));
	notech_inv i_52307(.A(to_acu2[174]), .Z(n_39367));
	notech_inv i_52308(.A(n_3198), .Z(n_39368));
	notech_inv i_52309(.A(to_acu2[175]), .Z(n_39369));
	notech_inv i_52310(.A(to_acu2[176]), .Z(n_39370));
	notech_inv i_52311(.A(n_3197), .Z(n_39371));
	notech_inv i_52312(.A(to_acu2[177]), .Z(n_39372));
	notech_inv i_52313(.A(to_acu2[178]), .Z(n_39373));
	notech_inv i_52314(.A(n_3196), .Z(n_39374));
	notech_inv i_52315(.A(to_acu2[179]), .Z(n_39375));
	notech_inv i_52316(.A(to_acu2[180]), .Z(n_39376));
	notech_inv i_52317(.A(n_3195), .Z(n_39377));
	notech_inv i_52318(.A(to_acu2[181]), .Z(n_39378));
	notech_inv i_52319(.A(to_acu2[182]), .Z(n_39379));
	notech_inv i_52320(.A(n_3194), .Z(n_39380));
	notech_inv i_52321(.A(to_acu2[183]), .Z(n_39381));
	notech_inv i_52322(.A(to_acu2[184]), .Z(n_39382));
	notech_inv i_52323(.A(n_3193), .Z(n_39383));
	notech_inv i_52324(.A(to_acu2[185]), .Z(n_39384));
	notech_inv i_52325(.A(to_acu2[186]), .Z(n_39385));
	notech_inv i_52326(.A(n_3192), .Z(n_39386));
	notech_inv i_52327(.A(to_acu2[187]), .Z(n_39387));
	notech_inv i_52328(.A(to_acu2[188]), .Z(n_39388));
	notech_inv i_52329(.A(n_3191), .Z(n_39389));
	notech_inv i_52330(.A(to_acu2[189]), .Z(n_39390));
	notech_inv i_52331(.A(to_acu2[190]), .Z(n_39391));
	notech_inv i_52332(.A(n_3190), .Z(n_39392));
	notech_inv i_52333(.A(to_acu2[191]), .Z(n_39393));
	notech_inv i_52334(.A(to_acu2[192]), .Z(n_39394));
	notech_inv i_52335(.A(n_3189), .Z(n_39395));
	notech_inv i_52336(.A(to_acu2[193]), .Z(n_39396));
	notech_inv i_52337(.A(to_acu2[194]), .Z(n_39397));
	notech_inv i_52338(.A(n_3188), .Z(n_39398));
	notech_inv i_52339(.A(to_acu2[195]), .Z(n_39399));
	notech_inv i_52340(.A(to_acu2[196]), .Z(n_39400));
	notech_inv i_52341(.A(n_3187), .Z(n_39401));
	notech_inv i_52342(.A(to_acu2[197]), .Z(n_39402));
	notech_inv i_52343(.A(to_acu2[198]), .Z(n_39403));
	notech_inv i_52344(.A(n_3186), .Z(n_39404));
	notech_inv i_52345(.A(to_acu2[199]), .Z(n_39405));
	notech_inv i_52346(.A(to_acu2[200]), .Z(n_39406));
	notech_inv i_52347(.A(n_3185), .Z(n_39407));
	notech_inv i_52348(.A(to_acu2[201]), .Z(n_39408));
	notech_inv i_52349(.A(to_acu2[202]), .Z(n_39409));
	notech_inv i_52350(.A(n_3184), .Z(n_39410));
	notech_inv i_52351(.A(to_acu2[203]), .Z(n_39411));
	notech_inv i_52352(.A(to_acu2[204]), .Z(n_39412));
	notech_inv i_52353(.A(n_3183), .Z(n_39413));
	notech_inv i_52354(.A(to_acu2[205]), .Z(n_39414));
	notech_inv i_52355(.A(to_acu2[206]), .Z(n_39415));
	notech_inv i_52356(.A(n_3182), .Z(n_39416));
	notech_inv i_52357(.A(to_acu2[207]), .Z(n_39417));
	notech_inv i_52358(.A(to_acu2[208]), .Z(n_39418));
	notech_inv i_52359(.A(n_3181), .Z(n_39419));
	notech_inv i_52360(.A(to_acu2[209]), .Z(n_39420));
	notech_inv i_52361(.A(to_acu2[210]), .Z(n_39421));
	notech_inv i_52362(.A(n_3180), .Z(n_39422));
	notech_inv i_52363(.A(to_acu1[0]), .Z(n_39423));
	notech_inv i_52364(.A(n_3179), .Z(n_39424));
	notech_inv i_52365(.A(n_48404), .Z(n_39425));
	notech_inv i_52366(.A(to_acu1[1]), .Z(n_39426));
	notech_inv i_52367(.A(n_3178), .Z(n_39427));
	notech_inv i_52368(.A(to_acu1[2]), .Z(n_39428));
	notech_inv i_52369(.A(n_48416), .Z(n_39429));
	notech_inv i_52370(.A(to_acu1[3]), .Z(n_39430));
	notech_inv i_52371(.A(n_3177), .Z(n_39431));
	notech_inv i_52372(.A(to_acu1[4]), .Z(n_39432));
	notech_inv i_52373(.A(n_3176), .Z(n_39433));
	notech_inv i_52374(.A(n_48428), .Z(n_39434));
	notech_inv i_52375(.A(to_acu1[5]), .Z(n_39435));
	notech_inv i_52376(.A(n_48434), .Z(n_39436));
	notech_inv i_52377(.A(to_acu1[6]), .Z(n_39437));
	notech_inv i_52378(.A(n_3175), .Z(n_39438));
	notech_inv i_52379(.A(n_48440), .Z(n_39439));
	notech_inv i_52380(.A(to_acu1[7]), .Z(n_39440));
	notech_inv i_52381(.A(n_3174), .Z(n_39441));
	notech_inv i_52382(.A(to_acu1[8]), .Z(n_39442));
	notech_inv i_52383(.A(n_48452), .Z(n_39443));
	notech_inv i_52384(.A(to_acu1[9]), .Z(n_39444));
	notech_inv i_52385(.A(n_3173), .Z(n_39445));
	notech_inv i_52386(.A(n_48458), .Z(n_39446));
	notech_inv i_52387(.A(to_acu1[10]), .Z(n_39447));
	notech_inv i_52388(.A(n_48464), .Z(n_39448));
	notech_inv i_52389(.A(to_acu1[11]), .Z(n_39449));
	notech_inv i_52390(.A(n_3172), .Z(n_39450));
	notech_inv i_52391(.A(to_acu1[12]), .Z(n_39451));
	notech_inv i_52392(.A(n_3171), .Z(n_39452));
	notech_inv i_52393(.A(to_acu1[13]), .Z(n_39453));
	notech_inv i_52394(.A(n_3170), .Z(n_39454));
	notech_inv i_52395(.A(to_acu1[14]), .Z(n_39455));
	notech_inv i_52396(.A(n_3169), .Z(n_39456));
	notech_inv i_52397(.A(n_48488), .Z(n_39457));
	notech_inv i_52398(.A(to_acu1[15]), .Z(n_39458));
	notech_inv i_52399(.A(n_48494), .Z(n_39459));
	notech_inv i_52400(.A(to_acu1[16]), .Z(n_39460));
	notech_inv i_52401(.A(n_3168), .Z(n_39461));
	notech_inv i_52402(.A(n_48500), .Z(n_39462));
	notech_inv i_52403(.A(to_acu1[17]), .Z(n_39463));
	notech_inv i_52404(.A(n_48506), .Z(n_39464));
	notech_inv i_52405(.A(to_acu1[18]), .Z(n_39465));
	notech_inv i_52406(.A(n_3167), .Z(n_39466));
	notech_inv i_52407(.A(n_48512), .Z(n_39467));
	notech_inv i_52408(.A(to_acu1[19]), .Z(n_39468));
	notech_inv i_52409(.A(n_48518), .Z(n_39469));
	notech_inv i_52410(.A(to_acu1[20]), .Z(n_39470));
	notech_inv i_52411(.A(n_3166), .Z(n_39471));
	notech_inv i_52412(.A(n_48524), .Z(n_39472));
	notech_inv i_52413(.A(to_acu1[21]), .Z(n_39473));
	notech_inv i_52414(.A(n_3165), .Z(n_39474));
	notech_inv i_52415(.A(to_acu1[22]), .Z(n_39475));
	notech_inv i_52416(.A(n_3164), .Z(n_39476));
	notech_inv i_52417(.A(to_acu1[23]), .Z(n_39477));
	notech_inv i_52418(.A(n_3163), .Z(n_39478));
	notech_inv i_52419(.A(to_acu1[24]), .Z(n_39479));
	notech_inv i_52420(.A(n_3162), .Z(n_39480));
	notech_inv i_52421(.A(to_acu1[25]), .Z(n_39481));
	notech_inv i_52422(.A(n_3161), .Z(n_39482));
	notech_inv i_52423(.A(to_acu1[26]), .Z(n_39483));
	notech_inv i_52424(.A(n_3160), .Z(n_39484));
	notech_inv i_52425(.A(to_acu1[27]), .Z(n_39485));
	notech_inv i_52426(.A(n_3159), .Z(n_39486));
	notech_inv i_52427(.A(to_acu1[28]), .Z(n_39487));
	notech_inv i_52428(.A(n_48572), .Z(n_39488));
	notech_inv i_52429(.A(to_acu1[29]), .Z(n_39489));
	notech_inv i_52430(.A(n_3158), .Z(n_39490));
	notech_inv i_52431(.A(n_48578), .Z(n_39491));
	notech_inv i_52432(.A(to_acu1[30]), .Z(n_39492));
	notech_inv i_52433(.A(n_48584), .Z(n_39493));
	notech_inv i_52434(.A(to_acu1[31]), .Z(n_39494));
	notech_inv i_52435(.A(n_3157), .Z(n_39495));
	notech_inv i_52436(.A(n_48590), .Z(n_39496));
	notech_inv i_52437(.A(to_acu1[32]), .Z(n_39497));
	notech_inv i_52438(.A(n_48596), .Z(n_39498));
	notech_inv i_52439(.A(to_acu1[33]), .Z(n_39499));
	notech_inv i_52440(.A(n_3156), .Z(n_39500));
	notech_inv i_52441(.A(n_48602), .Z(n_39501));
	notech_inv i_52442(.A(to_acu1[34]), .Z(n_39502));
	notech_inv i_52443(.A(n_48608), .Z(n_39503));
	notech_inv i_52444(.A(to_acu1[35]), .Z(n_39504));
	notech_inv i_52445(.A(n_3155), .Z(n_39505));
	notech_inv i_52446(.A(n_48614), .Z(n_39506));
	notech_inv i_52447(.A(to_acu1[36]), .Z(n_39507));
	notech_inv i_52448(.A(n_48620), .Z(n_39508));
	notech_inv i_52449(.A(to_acu1[37]), .Z(n_39509));
	notech_inv i_52450(.A(n_3154), .Z(n_39510));
	notech_inv i_52451(.A(n_48626), .Z(n_39511));
	notech_inv i_52452(.A(to_acu1[38]), .Z(n_39512));
	notech_inv i_52453(.A(n_3153), .Z(n_39513));
	notech_inv i_52454(.A(n_48638), .Z(n_39514));
	notech_inv i_52455(.A(to_acu1[40]), .Z(n_39515));
	notech_inv i_52456(.A(n_3152), .Z(n_39516));
	notech_inv i_52457(.A(n_48644), .Z(n_39517));
	notech_inv i_52458(.A(to_acu1[41]), .Z(n_39518));
	notech_inv i_52459(.A(n_48650), .Z(n_39519));
	notech_inv i_52460(.A(to_acu1[42]), .Z(n_39520));
	notech_inv i_52461(.A(n_3151), .Z(n_39521));
	notech_inv i_52462(.A(n_48656), .Z(n_39522));
	notech_inv i_52463(.A(to_acu1[43]), .Z(n_39523));
	notech_inv i_52464(.A(n_48662), .Z(n_39524));
	notech_inv i_52465(.A(to_acu1[44]), .Z(n_39525));
	notech_inv i_52466(.A(n_3150), .Z(n_39526));
	notech_inv i_52467(.A(n_48668), .Z(n_39527));
	notech_inv i_52468(.A(to_acu1[45]), .Z(n_39528));
	notech_inv i_52469(.A(n_48674), .Z(n_39529));
	notech_inv i_52470(.A(to_acu1[46]), .Z(n_39530));
	notech_inv i_52471(.A(n_3149), .Z(n_39531));
	notech_inv i_52472(.A(n_48680), .Z(n_39532));
	notech_inv i_52473(.A(to_acu1[47]), .Z(n_39533));
	notech_inv i_52474(.A(n_48686), .Z(n_39534));
	notech_inv i_52475(.A(to_acu1[48]), .Z(n_39535));
	notech_inv i_52476(.A(n_3148), .Z(n_39536));
	notech_inv i_52477(.A(n_48692), .Z(n_39537));
	notech_inv i_52478(.A(to_acu1[49]), .Z(n_39538));
	notech_inv i_52479(.A(n_48698), .Z(n_39539));
	notech_inv i_52480(.A(to_acu1[50]), .Z(n_39540));
	notech_inv i_52481(.A(n_3147), .Z(n_39541));
	notech_inv i_52482(.A(n_48704), .Z(n_39542));
	notech_inv i_52483(.A(to_acu1[51]), .Z(n_39543));
	notech_inv i_52484(.A(n_48710), .Z(n_39544));
	notech_inv i_52485(.A(to_acu1[52]), .Z(n_39545));
	notech_inv i_52486(.A(n_48716), .Z(n_39546));
	notech_inv i_52487(.A(to_acu1[53]), .Z(n_39547));
	notech_inv i_52488(.A(n_48722), .Z(n_39548));
	notech_inv i_52489(.A(to_acu1[54]), .Z(n_39549));
	notech_inv i_52490(.A(n_48728), .Z(n_39550));
	notech_inv i_52491(.A(to_acu1[55]), .Z(n_39551));
	notech_inv i_52492(.A(n_48734), .Z(n_39552));
	notech_inv i_52493(.A(to_acu1[56]), .Z(n_39553));
	notech_inv i_52494(.A(n_48740), .Z(n_39554));
	notech_inv i_52495(.A(to_acu1[57]), .Z(n_39555));
	notech_inv i_52496(.A(n_48746), .Z(n_39556));
	notech_inv i_52497(.A(to_acu1[58]), .Z(n_39557));
	notech_inv i_52498(.A(n_48752), .Z(n_39558));
	notech_inv i_52499(.A(to_acu1[59]), .Z(n_39559));
	notech_inv i_52500(.A(n_48758), .Z(n_39560));
	notech_inv i_52501(.A(to_acu1[60]), .Z(n_39561));
	notech_inv i_52502(.A(n_48764), .Z(n_39562));
	notech_inv i_52503(.A(to_acu1[61]), .Z(n_39563));
	notech_inv i_52504(.A(n_48770), .Z(n_39564));
	notech_inv i_52505(.A(to_acu1[62]), .Z(n_39565));
	notech_inv i_52506(.A(n_48776), .Z(n_39566));
	notech_inv i_52507(.A(to_acu1[63]), .Z(n_39567));
	notech_inv i_52508(.A(to_acu1[64]), .Z(n_39568));
	notech_inv i_52509(.A(to_acu1[65]), .Z(n_39569));
	notech_inv i_52510(.A(n_2123), .Z(n_39570));
	notech_inv i_52511(.A(to_acu1[66]), .Z(n_39571));
	notech_inv i_52512(.A(to_acu1[67]), .Z(n_39572));
	notech_inv i_52513(.A(n_48806), .Z(n_39573));
	notech_inv i_52514(.A(to_acu1[68]), .Z(n_39574));
	notech_inv i_52515(.A(to_acu1[69]), .Z(n_39575));
	notech_inv i_52516(.A(to_acu1[70]), .Z(n_39576));
	notech_inv i_52517(.A(to_acu1[71]), .Z(n_39577));
	notech_inv i_52518(.A(to_acu1[72]), .Z(n_39578));
	notech_inv i_52519(.A(to_acu1[73]), .Z(n_39579));
	notech_inv i_52520(.A(to_acu1[74]), .Z(n_39580));
	notech_inv i_52521(.A(to_acu1[75]), .Z(n_39581));
	notech_inv i_52522(.A(to_acu1[76]), .Z(n_39582));
	notech_inv i_52523(.A(to_acu1[77]), .Z(n_39583));
	notech_inv i_52524(.A(to_acu1[78]), .Z(n_39584));
	notech_inv i_52525(.A(to_acu1[79]), .Z(n_39585));
	notech_inv i_52526(.A(to_acu1[80]), .Z(n_39586));
	notech_inv i_52527(.A(to_acu1[81]), .Z(n_39587));
	notech_inv i_52528(.A(n_48890), .Z(n_39588));
	notech_inv i_52529(.A(to_acu1[82]), .Z(n_39589));
	notech_inv i_52530(.A(n_48896), .Z(n_39590));
	notech_inv i_52531(.A(to_acu1[83]), .Z(n_39591));
	notech_inv i_52532(.A(to_acu1[84]), .Z(n_39592));
	notech_inv i_52533(.A(n_3116), .Z(n_39593));
	notech_inv i_52534(.A(to_acu1[85]), .Z(n_39594));
	notech_inv i_52535(.A(n_3115), .Z(n_39595));
	notech_inv i_52536(.A(to_acu1[86]), .Z(n_39596));
	notech_inv i_52537(.A(n_48920), .Z(n_39597));
	notech_inv i_52538(.A(to_acu1[87]), .Z(n_39598));
	notech_inv i_52539(.A(n_48926), .Z(n_39599));
	notech_inv i_52540(.A(to_acu1[88]), .Z(n_39600));
	notech_inv i_52541(.A(n_3114), .Z(n_39601));
	notech_inv i_52542(.A(n_48932), .Z(n_39602));
	notech_inv i_52543(.A(to_acu1[89]), .Z(n_39603));
	notech_inv i_52544(.A(to_acu1[90]), .Z(n_39604));
	notech_inv i_52545(.A(n_3113), .Z(n_39605));
	notech_inv i_52546(.A(to_acu1[91]), .Z(n_39606));
	notech_inv i_52547(.A(n_3112), .Z(n_39607));
	notech_inv i_52548(.A(to_acu1[92]), .Z(n_39608));
	notech_inv i_52549(.A(to_acu1[93]), .Z(n_39609));
	notech_inv i_52550(.A(n_3111), .Z(n_39610));
	notech_inv i_52551(.A(to_acu1[94]), .Z(n_39611));
	notech_inv i_52552(.A(n_3110), .Z(n_39612));
	notech_inv i_52553(.A(to_acu1[95]), .Z(n_39613));
	notech_inv i_52554(.A(to_acu1[96]), .Z(n_39614));
	notech_inv i_52555(.A(n_3109), .Z(n_39615));
	notech_inv i_52556(.A(to_acu1[97]), .Z(n_39616));
	notech_inv i_52557(.A(to_acu1[98]), .Z(n_39617));
	notech_inv i_52558(.A(to_acu1[99]), .Z(n_39618));
	notech_inv i_52559(.A(n_3105), .Z(n_39619));
	notech_inv i_52560(.A(to_acu1[100]), .Z(n_39620));
	notech_inv i_52561(.A(n_49004), .Z(n_39621));
	notech_inv i_52562(.A(to_acu1[101]), .Z(n_39622));
	notech_inv i_52563(.A(n_49010), .Z(n_39623));
	notech_inv i_52564(.A(to_acu1[102]), .Z(n_39624));
	notech_inv i_52565(.A(n_3104), .Z(n_39625));
	notech_inv i_52566(.A(n_49016), .Z(n_39626));
	notech_inv i_52567(.A(to_acu1[103]), .Z(n_39627));
	notech_inv i_52568(.A(n_49022), .Z(n_39628));
	notech_inv i_52569(.A(to_acu1[104]), .Z(n_39629));
	notech_inv i_52570(.A(n_49028), .Z(n_39630));
	notech_inv i_52571(.A(to_acu1[105]), .Z(n_39631));
	notech_inv i_52572(.A(n_3103), .Z(n_39632));
	notech_inv i_52573(.A(to_acu1[106]), .Z(n_39633));
	notech_inv i_52574(.A(n_49040), .Z(n_39634));
	notech_inv i_52575(.A(to_acu1[107]), .Z(n_39635));
	notech_inv i_52576(.A(n_3102), .Z(n_39636));
	notech_inv i_52577(.A(n_49046), .Z(n_39637));
	notech_inv i_52578(.A(to_acu1[108]), .Z(n_39638));
	notech_inv i_52579(.A(n_49052), .Z(n_39639));
	notech_inv i_52580(.A(to_acu1[109]), .Z(n_39640));
	notech_inv i_52581(.A(n_49058), .Z(n_39641));
	notech_inv i_52582(.A(to_acu1[110]), .Z(n_39642));
	notech_inv i_52583(.A(n_3101), .Z(n_39643));
	notech_inv i_52584(.A(n_49064), .Z(n_39644));
	notech_inv i_52585(.A(to_acu1[111]), .Z(n_39645));
	notech_inv i_52586(.A(to_acu1[112]), .Z(n_39646));
	notech_inv i_52587(.A(n_3100), .Z(n_39647));
	notech_inv i_52588(.A(n_49076), .Z(n_39648));
	notech_inv i_52589(.A(to_acu1[113]), .Z(n_39649));
	notech_inv i_52590(.A(n_49082), .Z(n_39650));
	notech_inv i_52591(.A(to_acu1[114]), .Z(n_39651));
	notech_inv i_52592(.A(n_49088), .Z(n_39652));
	notech_inv i_52593(.A(to_acu1[115]), .Z(n_39653));
	notech_inv i_52594(.A(n_3099), .Z(n_39654));
	notech_inv i_52595(.A(n_49094), .Z(n_39655));
	notech_inv i_52596(.A(to_acu1[116]), .Z(n_39656));
	notech_inv i_52597(.A(n_49100), .Z(n_39657));
	notech_inv i_52598(.A(to_acu1[117]), .Z(n_39658));
	notech_inv i_52599(.A(n_49106), .Z(n_39659));
	notech_inv i_52600(.A(to_acu1[118]), .Z(n_39660));
	notech_inv i_52601(.A(n_3098), .Z(n_39661));
	notech_inv i_52602(.A(n_49112), .Z(n_39662));
	notech_inv i_52603(.A(to_acu1[119]), .Z(n_39663));
	notech_inv i_52604(.A(n_49118), .Z(n_39664));
	notech_inv i_52605(.A(to_acu1[120]), .Z(n_39665));
	notech_inv i_52606(.A(n_49124), .Z(n_39666));
	notech_inv i_52607(.A(to_acu1[121]), .Z(n_39667));
	notech_inv i_52608(.A(n_49130), .Z(n_39668));
	notech_inv i_52609(.A(to_acu1[122]), .Z(n_39669));
	notech_inv i_52610(.A(to_acu1[123]), .Z(n_39670));
	notech_inv i_52611(.A(to_acu1[124]), .Z(n_39671));
	notech_inv i_52612(.A(to_acu1[125]), .Z(n_39672));
	notech_inv i_52613(.A(to_acu1[126]), .Z(n_39673));
	notech_inv i_52614(.A(to_acu1[127]), .Z(n_39674));
	notech_inv i_52615(.A(n_49166), .Z(n_39675));
	notech_inv i_52616(.A(to_acu1[128]), .Z(n_39676));
	notech_inv i_52617(.A(n_49172), .Z(n_39677));
	notech_inv i_52618(.A(to_acu1[129]), .Z(n_39678));
	notech_inv i_52619(.A(n_49178), .Z(n_39679));
	notech_inv i_52620(.A(to_acu1[130]), .Z(n_39680));
	notech_inv i_52621(.A(n_49184), .Z(n_39681));
	notech_inv i_52622(.A(to_acu1[131]), .Z(n_39682));
	notech_inv i_52623(.A(n_49190), .Z(n_39683));
	notech_inv i_52624(.A(to_acu1[132]), .Z(n_39684));
	notech_inv i_52625(.A(n_49196), .Z(n_39685));
	notech_inv i_52626(.A(to_acu1[133]), .Z(n_39686));
	notech_inv i_52627(.A(n_49202), .Z(n_39687));
	notech_inv i_52628(.A(to_acu1[134]), .Z(n_39688));
	notech_inv i_52629(.A(n_49208), .Z(n_39689));
	notech_inv i_52630(.A(to_acu1[135]), .Z(n_39690));
	notech_inv i_52631(.A(n_49214), .Z(n_39691));
	notech_inv i_52632(.A(to_acu1[136]), .Z(n_39692));
	notech_inv i_52633(.A(n_49220), .Z(n_39693));
	notech_inv i_52634(.A(to_acu1[137]), .Z(n_39694));
	notech_inv i_52635(.A(to_acu1[138]), .Z(n_39695));
	notech_inv i_52636(.A(n_49232), .Z(n_39696));
	notech_inv i_52637(.A(to_acu1[139]), .Z(n_39697));
	notech_inv i_52638(.A(n_49238), .Z(n_39698));
	notech_inv i_52639(.A(to_acu1[140]), .Z(n_39699));
	notech_inv i_52640(.A(n_49244), .Z(n_39700));
	notech_inv i_52641(.A(to_acu1[141]), .Z(n_39701));
	notech_inv i_52642(.A(n_49250), .Z(n_39702));
	notech_inv i_52643(.A(to_acu1[142]), .Z(n_39703));
	notech_inv i_52644(.A(n_49256), .Z(n_39704));
	notech_inv i_52645(.A(to_acu1[143]), .Z(n_39705));
	notech_inv i_52646(.A(n_49262), .Z(n_39706));
	notech_inv i_52647(.A(to_acu1[144]), .Z(n_39707));
	notech_inv i_52648(.A(n_49268), .Z(n_39708));
	notech_inv i_52649(.A(to_acu1[145]), .Z(n_39709));
	notech_inv i_52650(.A(to_acu1[146]), .Z(n_39710));
	notech_inv i_52651(.A(n_49280), .Z(n_39711));
	notech_inv i_52652(.A(to_acu1[147]), .Z(n_39712));
	notech_inv i_52653(.A(n_49286), .Z(n_39713));
	notech_inv i_52654(.A(to_acu1[148]), .Z(n_39714));
	notech_inv i_52655(.A(n_49292), .Z(n_39715));
	notech_inv i_52656(.A(to_acu1[149]), .Z(n_39716));
	notech_inv i_52657(.A(n_49298), .Z(n_39717));
	notech_inv i_52658(.A(to_acu1[150]), .Z(n_39718));
	notech_inv i_52659(.A(n_49304), .Z(n_39719));
	notech_inv i_52660(.A(to_acu1[151]), .Z(n_39720));
	notech_inv i_52661(.A(n_49310), .Z(n_39721));
	notech_inv i_52662(.A(to_acu1[152]), .Z(n_39722));
	notech_inv i_52663(.A(n_49316), .Z(n_39723));
	notech_inv i_52664(.A(to_acu1[153]), .Z(n_39724));
	notech_inv i_52665(.A(n_49322), .Z(n_39725));
	notech_inv i_52666(.A(to_acu1[154]), .Z(n_39726));
	notech_inv i_52667(.A(n_49328), .Z(n_39727));
	notech_inv i_52668(.A(to_acu1[155]), .Z(n_39728));
	notech_inv i_52669(.A(n_49334), .Z(n_39729));
	notech_inv i_52670(.A(to_acu1[156]), .Z(n_39730));
	notech_inv i_52671(.A(n_49340), .Z(n_39731));
	notech_inv i_52672(.A(to_acu1[157]), .Z(n_39732));
	notech_inv i_52673(.A(n_49346), .Z(n_39733));
	notech_inv i_52674(.A(to_acu1[158]), .Z(n_39734));
	notech_inv i_52675(.A(n_49352), .Z(n_39735));
	notech_inv i_52676(.A(to_acu1[159]), .Z(n_39736));
	notech_inv i_52677(.A(n_49358), .Z(n_39737));
	notech_inv i_52678(.A(to_acu1[160]), .Z(n_39738));
	notech_inv i_52679(.A(n_49364), .Z(n_39739));
	notech_inv i_52680(.A(to_acu1[161]), .Z(n_39740));
	notech_inv i_52681(.A(n_49370), .Z(n_39741));
	notech_inv i_52682(.A(to_acu1[162]), .Z(n_39742));
	notech_inv i_52683(.A(to_acu1[163]), .Z(n_39743));
	notech_inv i_52684(.A(to_acu1[164]), .Z(n_39744));
	notech_inv i_52685(.A(to_acu1[165]), .Z(n_39745));
	notech_inv i_52686(.A(to_acu1[166]), .Z(n_39746));
	notech_inv i_52687(.A(to_acu1[167]), .Z(n_39747));
	notech_inv i_52688(.A(to_acu1[168]), .Z(n_39748));
	notech_inv i_52689(.A(to_acu1[169]), .Z(n_39749));
	notech_inv i_52690(.A(n_49418), .Z(n_39750));
	notech_inv i_52691(.A(to_acu1[170]), .Z(n_39751));
	notech_inv i_52692(.A(n_49424), .Z(n_39752));
	notech_inv i_52693(.A(to_acu1[171]), .Z(n_39753));
	notech_inv i_52694(.A(to_acu1[172]), .Z(n_39754));
	notech_inv i_52695(.A(to_acu1[173]), .Z(n_39755));
	notech_inv i_52696(.A(n_49442), .Z(n_39756));
	notech_inv i_52697(.A(to_acu1[174]), .Z(n_39757));
	notech_inv i_52698(.A(to_acu1[175]), .Z(n_39758));
	notech_inv i_52699(.A(n_49454), .Z(n_39759));
	notech_inv i_52700(.A(to_acu1[176]), .Z(n_39760));
	notech_inv i_52701(.A(n_49460), .Z(n_39761));
	notech_inv i_52702(.A(to_acu1[177]), .Z(n_39762));
	notech_inv i_52703(.A(to_acu1[178]), .Z(n_39763));
	notech_inv i_52704(.A(n_49472), .Z(n_39764));
	notech_inv i_52705(.A(to_acu1[179]), .Z(n_39765));
	notech_inv i_52706(.A(n_49478), .Z(n_39766));
	notech_inv i_52707(.A(to_acu1[180]), .Z(n_39767));
	notech_inv i_52708(.A(n_49484), .Z(n_39768));
	notech_inv i_52709(.A(to_acu1[181]), .Z(n_39769));
	notech_inv i_52710(.A(n_49490), .Z(n_39770));
	notech_inv i_52711(.A(to_acu1[182]), .Z(n_39771));
	notech_inv i_52712(.A(n_49496), .Z(n_39772));
	notech_inv i_52713(.A(to_acu1[183]), .Z(n_39773));
	notech_inv i_52714(.A(n_49502), .Z(n_39774));
	notech_inv i_52715(.A(to_acu1[184]), .Z(n_39775));
	notech_inv i_52716(.A(n_49508), .Z(n_39776));
	notech_inv i_52717(.A(to_acu1[185]), .Z(n_39777));
	notech_inv i_52718(.A(n_49514), .Z(n_39778));
	notech_inv i_52719(.A(to_acu1[186]), .Z(n_39779));
	notech_inv i_52720(.A(n_49520), .Z(n_39780));
	notech_inv i_52721(.A(to_acu1[187]), .Z(n_39781));
	notech_inv i_52722(.A(n_49526), .Z(n_39782));
	notech_inv i_52723(.A(to_acu1[188]), .Z(n_39783));
	notech_inv i_52724(.A(n_49532), .Z(n_39784));
	notech_inv i_52725(.A(to_acu1[189]), .Z(n_39785));
	notech_inv i_52726(.A(n_49538), .Z(n_39786));
	notech_inv i_52727(.A(to_acu1[190]), .Z(n_39787));
	notech_inv i_52728(.A(n_49544), .Z(n_39788));
	notech_inv i_52729(.A(to_acu1[191]), .Z(n_39789));
	notech_inv i_52730(.A(n_49550), .Z(n_39790));
	notech_inv i_52731(.A(to_acu1[192]), .Z(n_39791));
	notech_inv i_52732(.A(n_49556), .Z(n_39792));
	notech_inv i_52733(.A(to_acu1[193]), .Z(n_39793));
	notech_inv i_52734(.A(n_49562), .Z(n_39794));
	notech_inv i_52735(.A(to_acu1[194]), .Z(n_39795));
	notech_inv i_52736(.A(n_49568), .Z(n_39796));
	notech_inv i_52737(.A(to_acu1[195]), .Z(n_39797));
	notech_inv i_52738(.A(n_49574), .Z(n_39798));
	notech_inv i_52739(.A(to_acu1[196]), .Z(n_39799));
	notech_inv i_52740(.A(to_acu1[197]), .Z(n_39800));
	notech_inv i_52741(.A(to_acu1[198]), .Z(n_39801));
	notech_inv i_52742(.A(to_acu1[199]), .Z(n_39802));
	notech_inv i_52743(.A(to_acu1[200]), .Z(n_39803));
	notech_inv i_52744(.A(n_49604), .Z(n_39804));
	notech_inv i_52745(.A(to_acu1[201]), .Z(n_39805));
	notech_inv i_52746(.A(to_acu1[202]), .Z(n_39806));
	notech_inv i_52747(.A(to_acu1[203]), .Z(n_39807));
	notech_inv i_52748(.A(n_49622), .Z(n_39808));
	notech_inv i_52749(.A(to_acu1[204]), .Z(n_39809));
	notech_inv i_52750(.A(n_49628), .Z(n_39810));
	notech_inv i_52751(.A(to_acu1[205]), .Z(n_39811));
	notech_inv i_52752(.A(n_49634), .Z(n_39812));
	notech_inv i_52753(.A(to_acu1[206]), .Z(n_39813));
	notech_inv i_52754(.A(to_acu1[207]), .Z(n_39814));
	notech_inv i_52755(.A(n_49646), .Z(n_39815));
	notech_inv i_52756(.A(to_acu1[208]), .Z(n_39816));
	notech_inv i_52757(.A(n_49652), .Z(n_39817));
	notech_inv i_52758(.A(to_acu1[209]), .Z(n_39818));
	notech_inv i_52759(.A(n_49658), .Z(n_39819));
	notech_inv i_52760(.A(to_acu1[210]), .Z(n_39820));
	notech_inv i_52761(.A(n_46767), .Z(n_39821));
	notech_inv i_52762(.A(opz2[0]), .Z(n_39822));
	notech_inv i_52763(.A(opz2[1]), .Z(n_39823));
	notech_inv i_52764(.A(opz1[0]), .Z(n_39824));
	notech_inv i_52765(.A(opz1[1]), .Z(n_39825));
	notech_inv i_52766(.A(n_2961), .Z(n_39826));
	notech_inv i_52767(.A(n_41904), .Z(n_39827));
	notech_inv i_52768(.A(lenpc2[0]), .Z(n_39828));
	notech_inv i_52769(.A(lenpc2[1]), .Z(n_39829));
	notech_inv i_52770(.A(lenpc2[2]), .Z(n_39830));
	notech_inv i_52771(.A(lenpc2[3]), .Z(n_39831));
	notech_inv i_52772(.A(lenpc2[4]), .Z(n_39832));
	notech_inv i_52773(.A(lenpc2[5]), .Z(n_39833));
	notech_inv i_52774(.A(n_2917), .Z(n_39834));
	notech_inv i_52775(.A(n_2890), .Z(n_39835));
	notech_inv i_52776(.A(lenpc1[0]), .Z(n_39836));
	notech_inv i_52777(.A(lenpc1[1]), .Z(n_39837));
	notech_inv i_52778(.A(n_2904), .Z(n_39838));
	notech_inv i_52779(.A(lenpc1[2]), .Z(n_39839));
	notech_inv i_52780(.A(lenpc1[3]), .Z(n_39840));
	notech_inv i_52781(.A(n_2155), .Z(n_39841));
	notech_inv i_52782(.A(lenpc1[4]), .Z(n_39842));
	notech_inv i_52783(.A(n_2900), .Z(n_39843));
	notech_inv i_52784(.A(lenpc1[5]), .Z(n_39844));
	notech_inv i_52785(.A(n_2893), .Z(n_39845));
	notech_inv i_52786(.A(n_2888), .Z(n_39846));
	notech_inv i_52787(.A(n_2138), .Z(n_39847));
	notech_inv i_52788(.A(n_2847), .Z(n_39848));
	notech_inv i_52789(.A(n_2844), .Z(n_39849));
	notech_inv i_52790(.A(n_2841), .Z(n_39850));
	notech_inv i_52791(.A(n_2837), .Z(n_39851));
	notech_inv i_52792(.A(n_2836), .Z(n_39852));
	notech_inv i_52793(.A(n_261791464), .Z(n_39853));
	notech_inv i_52794(.A(n_43906), .Z(n_39854));
	notech_inv i_52795(.A(n_43954), .Z(n_39855));
	notech_inv i_52796(.A(n_44092), .Z(n_39856));
	notech_inv i_52797(.A(n_42938), .Z(n_39857));
	notech_inv i_52798(.A(n_42944), .Z(n_39858));
	notech_inv i_52799(.A(imm_sz[1]), .Z(n_39859));
	notech_inv i_52800(.A(imm_sz[2]), .Z(n_39860));
	notech_inv i_52801(.A(displc[0]), .Z(n_39861));
	notech_inv i_52802(.A(udeco[0]), .Z(n_39862));
	notech_inv i_52803(.A(udeco[1]), .Z(n_39863));
	notech_inv i_52804(.A(udeco[2]), .Z(n_39864));
	notech_inv i_52805(.A(udeco[3]), .Z(n_39865));
	notech_inv i_52806(.A(udeco[4]), .Z(n_39866));
	notech_inv i_52807(.A(udeco[5]), .Z(n_39867));
	notech_inv i_52808(.A(udeco[6]), .Z(n_39868));
	notech_inv i_52809(.A(udeco[7]), .Z(n_39869));
	notech_inv i_52810(.A(udeco[8]), .Z(n_39870));
	notech_inv i_52811(.A(udeco[9]), .Z(n_39871));
	notech_inv i_52812(.A(udeco[10]), .Z(n_39872));
	notech_inv i_52813(.A(udeco[11]), .Z(n_39873));
	notech_inv i_52814(.A(udeco[12]), .Z(n_39874));
	notech_inv i_52815(.A(udeco[13]), .Z(n_39875));
	notech_inv i_52816(.A(udeco[14]), .Z(n_39876));
	notech_inv i_52817(.A(udeco[15]), .Z(n_39877));
	notech_inv i_52818(.A(udeco[16]), .Z(n_39878));
	notech_inv i_52819(.A(udeco[17]), .Z(n_39879));
	notech_inv i_52820(.A(udeco[18]), .Z(n_39880));
	notech_inv i_52821(.A(udeco[19]), .Z(n_39881));
	notech_inv i_52822(.A(udeco[20]), .Z(n_39882));
	notech_inv i_52823(.A(udeco[21]), .Z(n_39883));
	notech_inv i_52824(.A(udeco[22]), .Z(n_39884));
	notech_inv i_52825(.A(udeco[23]), .Z(n_39885));
	notech_inv i_52826(.A(udeco[24]), .Z(n_39886));
	notech_inv i_52827(.A(udeco[25]), .Z(n_39887));
	notech_inv i_52828(.A(udeco[26]), .Z(n_39888));
	notech_inv i_52829(.A(udeco[27]), .Z(n_39889));
	notech_inv i_52830(.A(udeco[28]), .Z(n_39890));
	notech_inv i_52831(.A(udeco[29]), .Z(n_39891));
	notech_inv i_52832(.A(udeco[30]), .Z(n_39892));
	notech_inv i_52833(.A(udeco[31]), .Z(n_39893));
	notech_inv i_52834(.A(udeco[32]), .Z(n_39894));
	notech_inv i_52835(.A(udeco[33]), .Z(n_39895));
	notech_inv i_52836(.A(udeco[34]), .Z(n_39896));
	notech_inv i_52837(.A(udeco[35]), .Z(n_39897));
	notech_inv i_52838(.A(udeco[36]), .Z(n_39898));
	notech_inv i_52839(.A(udeco[37]), .Z(n_39899));
	notech_inv i_52840(.A(udeco[38]), .Z(n_39900));
	notech_inv i_52841(.A(udeco[39]), .Z(n_39901));
	notech_inv i_52842(.A(udeco[40]), .Z(n_39902));
	notech_inv i_52843(.A(udeco[41]), .Z(n_39903));
	notech_inv i_52844(.A(udeco[42]), .Z(n_39904));
	notech_inv i_52845(.A(udeco[43]), .Z(n_39905));
	notech_inv i_52846(.A(udeco[44]), .Z(n_39906));
	notech_inv i_52847(.A(udeco[45]), .Z(n_39907));
	notech_inv i_52848(.A(udeco[46]), .Z(n_39908));
	notech_inv i_52849(.A(udeco[47]), .Z(n_39909));
	notech_inv i_52850(.A(udeco[48]), .Z(n_39910));
	notech_inv i_52851(.A(udeco[49]), .Z(n_39911));
	notech_inv i_52852(.A(udeco[50]), .Z(n_39912));
	notech_inv i_52853(.A(udeco[51]), .Z(n_39913));
	notech_inv i_52854(.A(udeco[52]), .Z(n_39914));
	notech_inv i_52855(.A(udeco[53]), .Z(n_39915));
	notech_inv i_52856(.A(udeco[54]), .Z(n_39916));
	notech_inv i_52857(.A(udeco[55]), .Z(n_39917));
	notech_inv i_52858(.A(udeco[56]), .Z(n_39918));
	notech_inv i_52859(.A(udeco[57]), .Z(n_39919));
	notech_inv i_52860(.A(udeco[58]), .Z(n_39920));
	notech_inv i_52861(.A(udeco[59]), .Z(n_39921));
	notech_inv i_52862(.A(udeco[60]), .Z(n_39922));
	notech_inv i_52863(.A(udeco[61]), .Z(n_39923));
	notech_inv i_52864(.A(udeco[62]), .Z(n_39924));
	notech_inv i_52865(.A(udeco[63]), .Z(n_39925));
	notech_inv i_52866(.A(udeco[64]), .Z(n_39926));
	notech_inv i_52867(.A(udeco[65]), .Z(n_39927));
	notech_inv i_52868(.A(udeco[66]), .Z(n_39928));
	notech_inv i_52869(.A(udeco[67]), .Z(n_39929));
	notech_inv i_52870(.A(udeco[68]), .Z(n_39930));
	notech_inv i_52871(.A(udeco[69]), .Z(n_39931));
	notech_inv i_52872(.A(udeco[70]), .Z(n_39932));
	notech_inv i_52873(.A(udeco[71]), .Z(n_39933));
	notech_inv i_52874(.A(udeco[72]), .Z(n_39934));
	notech_inv i_52875(.A(udeco[73]), .Z(n_39935));
	notech_inv i_52876(.A(udeco[74]), .Z(n_39936));
	notech_inv i_52877(.A(udeco[75]), .Z(n_39937));
	notech_inv i_52878(.A(udeco[76]), .Z(n_39938));
	notech_inv i_52879(.A(udeco[77]), .Z(n_39939));
	notech_inv i_52880(.A(udeco[78]), .Z(n_39940));
	notech_inv i_52881(.A(udeco[79]), .Z(n_39941));
	notech_inv i_52882(.A(udeco[80]), .Z(n_39942));
	notech_inv i_52883(.A(udeco[81]), .Z(n_39943));
	notech_inv i_52884(.A(udeco[82]), .Z(n_39944));
	notech_inv i_52885(.A(udeco[83]), .Z(n_39945));
	notech_inv i_52886(.A(udeco[84]), .Z(n_39946));
	notech_inv i_52887(.A(udeco[85]), .Z(n_39947));
	notech_inv i_52888(.A(udeco[86]), .Z(n_39948));
	notech_inv i_52889(.A(udeco[87]), .Z(n_39949));
	notech_inv i_52890(.A(udeco[88]), .Z(n_39950));
	notech_inv i_52891(.A(udeco[89]), .Z(n_39951));
	notech_inv i_52892(.A(udeco[90]), .Z(n_39952));
	notech_inv i_52893(.A(udeco[91]), .Z(n_39953));
	notech_inv i_52894(.A(udeco[92]), .Z(n_39954));
	notech_inv i_52895(.A(udeco[93]), .Z(n_39955));
	notech_inv i_52896(.A(udeco[94]), .Z(n_39956));
	notech_inv i_52897(.A(udeco[95]), .Z(n_39957));
	notech_inv i_52898(.A(udeco[96]), .Z(n_39958));
	notech_inv i_52899(.A(udeco[97]), .Z(n_39959));
	notech_inv i_52900(.A(udeco[98]), .Z(n_39960));
	notech_inv i_52901(.A(udeco[99]), .Z(n_39961));
	notech_inv i_52902(.A(udeco[100]), .Z(n_39962));
	notech_inv i_52903(.A(udeco[101]), .Z(n_39963));
	notech_inv i_52904(.A(udeco[102]), .Z(n_39964));
	notech_inv i_52905(.A(udeco[103]), .Z(n_39965));
	notech_inv i_52906(.A(udeco[104]), .Z(n_39966));
	notech_inv i_52907(.A(udeco[105]), .Z(n_39967));
	notech_inv i_52908(.A(udeco[106]), .Z(n_39968));
	notech_inv i_52909(.A(udeco[107]), .Z(n_39969));
	notech_inv i_52910(.A(udeco[108]), .Z(n_39970));
	notech_inv i_52911(.A(udeco[109]), .Z(n_39971));
	notech_inv i_52912(.A(udeco[110]), .Z(n_39972));
	notech_inv i_52913(.A(udeco[111]), .Z(n_39973));
	notech_inv i_52914(.A(udeco[112]), .Z(n_39974));
	notech_inv i_52915(.A(udeco[113]), .Z(n_39975));
	notech_inv i_52916(.A(udeco[114]), .Z(n_39976));
	notech_inv i_52917(.A(udeco[115]), .Z(n_39977));
	notech_inv i_52918(.A(udeco[116]), .Z(n_39978));
	notech_inv i_52919(.A(udeco[117]), .Z(n_39979));
	notech_inv i_52920(.A(udeco[118]), .Z(n_39980));
	notech_inv i_52921(.A(udeco[119]), .Z(n_39981));
	notech_inv i_52922(.A(udeco[120]), .Z(n_39982));
	notech_inv i_52923(.A(udeco[121]), .Z(n_39983));
	notech_inv i_52924(.A(udeco[122]), .Z(n_39984));
	notech_inv i_52925(.A(udeco[123]), .Z(n_39985));
	notech_inv i_52926(.A(udeco[124]), .Z(n_39986));
	notech_inv i_52927(.A(udeco[125]), .Z(n_39987));
	notech_inv i_52928(.A(udeco[126]), .Z(n_39988));
	notech_inv i_52929(.A(udeco[127]), .Z(n_39989));
	notech_inv i_52930(.A(valid_len[5]), .Z(n_39990));
	notech_inv i_52931(.A(in128[16]), .Z(n_39991));
	notech_inv i_52932(.A(in128[17]), .Z(n_39992));
	notech_inv i_52933(.A(in128[18]), .Z(n_39993));
	notech_inv i_52934(.A(in128[19]), .Z(n_39994));
	notech_inv i_52935(.A(in128[20]), .Z(n_39995));
	notech_inv i_52936(.A(in128[21]), .Z(n_39996));
	notech_inv i_52937(.A(in128[22]), .Z(n_39997));
	notech_inv i_52938(.A(in128[23]), .Z(n_39998));
	notech_inv i_52939(.A(in128[24]), .Z(n_39999));
	notech_inv i_52940(.A(in128[25]), .Z(n_40000));
	notech_inv i_52941(.A(in128[26]), .Z(n_40001));
	notech_inv i_52942(.A(in128[27]), .Z(n_40002));
	notech_inv i_52943(.A(in128[28]), .Z(n_40003));
	notech_inv i_52944(.A(in128[29]), .Z(n_40004));
	notech_inv i_52945(.A(in128[30]), .Z(n_40005));
	notech_inv i_52946(.A(in128[31]), .Z(n_40006));
	notech_inv i_52947(.A(in128[32]), .Z(n_40007));
	notech_inv i_52948(.A(in128[33]), .Z(n_40008));
	notech_inv i_52949(.A(in128[34]), .Z(n_40009));
	notech_inv i_52950(.A(in128[35]), .Z(n_40010));
	notech_inv i_52951(.A(in128[36]), .Z(n_40011));
	notech_inv i_52952(.A(in128[37]), .Z(n_40012));
	notech_inv i_52953(.A(in128[38]), .Z(n_40013));
	notech_inv i_52954(.A(in128[39]), .Z(n_40014));
	notech_inv i_52955(.A(in128[40]), .Z(n_40015));
	notech_inv i_52956(.A(in128[41]), .Z(n_40016));
	notech_inv i_52957(.A(in128[42]), .Z(n_40017));
	notech_inv i_52958(.A(in128[43]), .Z(n_40018));
	notech_inv i_52959(.A(in128[44]), .Z(n_40019));
	notech_inv i_52960(.A(in128[45]), .Z(n_40020));
	notech_inv i_52961(.A(in128[46]), .Z(n_40021));
	notech_inv i_52962(.A(in128[47]), .Z(n_40022));
	notech_inv i_52963(.A(in128[48]), .Z(n_40023));
	notech_inv i_52964(.A(in128[49]), .Z(n_40024));
	notech_inv i_52965(.A(in128[50]), .Z(n_40025));
	notech_inv i_52966(.A(in128[51]), .Z(n_40026));
	notech_inv i_52967(.A(in128[52]), .Z(n_40027));
	notech_inv i_52968(.A(in128[53]), .Z(n_40028));
	notech_inv i_52969(.A(in128[54]), .Z(n_40029));
	notech_inv i_52970(.A(in128[55]), .Z(n_40030));
	notech_inv i_52971(.A(in128[56]), .Z(n_40031));
	notech_inv i_52972(.A(in128[57]), .Z(n_40032));
	notech_inv i_52973(.A(in128[58]), .Z(n_40033));
	notech_inv i_52974(.A(in128[59]), .Z(n_40034));
	notech_inv i_52975(.A(in128[60]), .Z(n_40035));
	notech_inv i_52976(.A(in128[61]), .Z(n_40036));
	notech_inv i_52977(.A(in128[62]), .Z(n_40037));
	notech_inv i_52978(.A(in128[63]), .Z(n_40038));
	notech_inv i_52979(.A(in128[64]), .Z(n_40039));
	notech_inv i_52980(.A(in128[65]), .Z(n_40040));
	notech_inv i_52981(.A(in128[66]), .Z(n_40041));
	notech_inv i_52982(.A(in128[67]), .Z(n_40042));
	notech_inv i_52983(.A(in128[68]), .Z(n_40043));
	notech_inv i_52984(.A(in128[69]), .Z(n_40044));
	notech_inv i_52985(.A(in128[70]), .Z(n_40045));
	notech_inv i_52986(.A(in128[71]), .Z(n_40046));
	notech_inv i_52987(.A(in128[72]), .Z(n_40047));
	notech_inv i_52988(.A(in128[73]), .Z(n_40048));
	notech_inv i_52989(.A(in128[74]), .Z(n_40049));
	notech_inv i_52990(.A(in128[75]), .Z(n_40050));
	notech_inv i_52991(.A(in128[76]), .Z(n_40051));
	notech_inv i_52992(.A(in128[77]), .Z(n_40052));
	notech_inv i_52993(.A(in128[78]), .Z(n_40053));
	notech_inv i_52994(.A(in128[79]), .Z(n_40054));
	notech_inv i_52995(.A(in128[80]), .Z(n_40055));
	notech_inv i_52996(.A(in128[81]), .Z(n_40056));
	notech_inv i_52997(.A(in128[82]), .Z(n_40057));
	notech_inv i_52998(.A(in128[83]), .Z(n_40058));
	notech_inv i_52999(.A(in128[84]), .Z(n_40059));
	notech_inv i_53000(.A(in128[85]), .Z(n_40060));
	notech_inv i_53001(.A(in128[86]), .Z(n_40061));
	notech_inv i_53002(.A(in128[87]), .Z(n_40062));
	notech_inv i_53003(.A(in128[88]), .Z(n_40063));
	notech_inv i_53004(.A(in128[89]), .Z(n_40064));
	notech_inv i_53005(.A(in128[90]), .Z(n_40065));
	notech_inv i_53006(.A(in128[91]), .Z(n_40066));
	notech_inv i_53007(.A(in128[92]), .Z(n_40067));
	notech_inv i_53008(.A(in128[93]), .Z(n_40068));
	notech_inv i_53009(.A(in128[94]), .Z(n_40069));
	notech_inv i_53010(.A(in128[95]), .Z(n_40070));
	notech_inv i_53011(.A(in128[96]), .Z(n_40071));
	notech_inv i_53012(.A(in128[97]), .Z(n_40072));
	notech_inv i_53013(.A(in128[98]), .Z(n_40073));
	notech_inv i_53014(.A(in128[99]), .Z(n_40074));
	notech_inv i_53015(.A(in128[100]), .Z(n_40075));
	notech_inv i_53016(.A(in128[101]), .Z(n_40076));
	notech_inv i_53017(.A(in128[102]), .Z(n_40077));
	notech_inv i_53018(.A(in128[103]), .Z(n_40078));
	notech_inv i_53019(.A(in128[104]), .Z(n_40079));
	notech_inv i_53020(.A(in128[105]), .Z(n_40080));
	notech_inv i_53021(.A(in128[106]), .Z(n_40081));
	notech_inv i_53022(.A(in128[107]), .Z(n_40082));
	notech_inv i_53023(.A(in128[108]), .Z(n_40083));
	notech_inv i_53024(.A(in128[109]), .Z(n_40084));
	notech_inv i_53025(.A(in128[110]), .Z(n_40085));
	notech_inv i_53026(.A(in128[111]), .Z(n_40086));
	notech_inv i_53027(.A(in128[112]), .Z(n_40087));
	notech_inv i_53028(.A(in128[113]), .Z(n_40088));
	notech_inv i_53029(.A(in128[114]), .Z(n_40089));
	notech_inv i_53030(.A(in128[115]), .Z(n_40090));
	notech_inv i_53031(.A(in128[116]), .Z(n_40091));
	notech_inv i_53032(.A(in128[117]), .Z(n_40092));
	notech_inv i_53033(.A(in128[118]), .Z(n_40093));
	notech_inv i_53034(.A(in128[119]), .Z(n_40094));
	notech_inv i_53035(.A(in128[120]), .Z(n_40095));
	notech_inv i_53036(.A(in128[121]), .Z(n_40096));
	notech_inv i_53037(.A(in128[122]), .Z(n_40097));
	notech_inv i_53038(.A(in128[123]), .Z(n_40098));
	notech_inv i_53039(.A(in128[124]), .Z(n_40099));
	notech_inv i_53040(.A(in128[125]), .Z(n_40100));
	notech_inv i_53041(.A(in128[126]), .Z(n_40101));
	notech_inv i_53042(.A(in128[127]), .Z(n_40102));
	notech_inv i_53043(.A(pfx_sz[1]), .Z(n_40103));
	notech_inv i_53044(.A(opz[0]), .Z(n_40104));
	notech_inv i_53045(.A(opz[1]), .Z(n_40105));
	notech_inv i_53046(.A(n_1486), .Z(n_40106));
	notech_inv i_53047(.A(\to_acu2_0[67] ), .Z(n_40107));
	notech_inv i_53048(.A(\to_acu2_0[66] ), .Z(n_40108));
	notech_inv i_53049(.A(\to_acu2_0[65] ), .Z(n_40109));
	notech_inv i_53050(.A(\to_acu2_0[64] ), .Z(n_40110));
	notech_inv i_53051(.A(\to_acu2_0[63] ), .Z(n_40111));
	notech_inv i_53052(.A(\to_acu2_0[60] ), .Z(n_40112));
	notech_inv i_53053(.A(\to_acu2_0[49] ), .Z(n_40113));
	notech_inv i_53054(.A(\to_acu2_0[33] ), .Z(n_40114));
	notech_inv i_53055(.A(\to_acu2_0[32] ), .Z(n_40115));
	notech_inv i_53056(.A(\to_acu2_0[31] ), .Z(n_40116));
	notech_inv i_53057(.A(\to_acu2_0[30] ), .Z(n_40117));
	notech_inv i_53058(.A(\to_acu2_0[29] ), .Z(n_40118));
	notech_inv i_53059(.A(\to_acu2_0[6] ), .Z(n_40119));
	notech_inv i_53060(.A(\to_acu2_0[56] ), .Z(n_40120));
	notech_inv i_53061(.A(\to_acu2_0[50] ), .Z(n_40121));
	notech_inv i_53062(.A(\to_acu2_0[58] ), .Z(n_40122));
	notech_inv i_53063(.A(\to_acu2_0[57] ), .Z(n_40123));
	notech_inv i_53064(.A(\to_acu2_0[52] ), .Z(n_40124));
	notech_inv i_53065(.A(\to_acu2_0[51] ), .Z(n_40125));
	notech_inv i_53066(.A(\to_acu2_0[53] ), .Z(n_40126));
	notech_inv i_53067(.A(\to_acu2_0[55] ), .Z(n_40127));
	notech_inv i_53068(.A(\to_acu2_0[54] ), .Z(n_40128));
	notech_inv i_53069(.A(\to_acu2_0[59] ), .Z(n_40129));
	notech_inv i_53070(.A(\to_acu2_0[5] ), .Z(n_40130));
	notech_inv i_53071(.A(\to_acu2_0[48] ), .Z(n_40131));
	notech_inv i_53072(.A(\to_acu2_0[35] ), .Z(n_40132));
	notech_inv i_53073(.A(\to_acu2_0[34] ), .Z(n_40133));
	notech_inv i_53074(.A(\to_acu2_0[37] ), .Z(n_40134));
	notech_inv i_53075(.A(\to_acu2_0[36] ), .Z(n_40135));
	notech_inv i_53076(.A(\to_acu2_0[40] ), .Z(n_40136));
	notech_inv i_53077(.A(\to_acu2_0[38] ), .Z(n_40137));
	notech_inv i_53078(.A(\to_acu2_0[41] ), .Z(n_40138));
	notech_inv i_53079(.A(\to_acu2_0[43] ), .Z(n_40139));
	notech_inv i_53080(.A(\to_acu2_0[42] ), .Z(n_40140));
	notech_inv i_53081(.A(\to_acu2_0[44] ), .Z(n_40141));
	notech_inv i_53082(.A(\to_acu2_0[46] ), .Z(n_40142));
	notech_inv i_53083(.A(\to_acu2_0[45] ), .Z(n_40143));
	notech_inv i_53084(.A(\to_acu2_0[47] ), .Z(n_40144));
	notech_inv i_53085(.A(\to_acu2_0[61] ), .Z(n_40145));
	notech_inv i_53086(.A(\to_acu2_0[7] ), .Z(n_40146));
	notech_inv i_53087(.A(\to_acu2_0[2] ), .Z(n_40147));
	notech_inv i_53088(.A(\to_acu2_0[1] ), .Z(n_40148));
	notech_inv i_53089(.A(\to_acu2_0[15] ), .Z(n_40149));
	notech_inv i_53090(.A(\to_acu2_0[14] ), .Z(n_40150));
	notech_inv i_53091(.A(\to_acu2_0[13] ), .Z(n_40151));
	notech_inv i_53092(.A(\to_acu2_0[17] ), .Z(n_40152));
	notech_inv i_53093(.A(\to_acu2_0[18] ), .Z(n_40153));
	notech_inv i_53094(.A(\to_acu2_0[12] ), .Z(n_40154));
	notech_inv i_53095(.A(\to_acu2_0[20] ), .Z(n_40155));
	notech_inv i_53096(.A(\to_acu2_0[21] ), .Z(n_40156));
	notech_inv i_53097(.A(\to_acu2_0[23] ), .Z(n_40157));
	notech_inv i_53098(.A(\to_acu2_0[22] ), .Z(n_40158));
	notech_inv i_53099(.A(\to_acu2_0[27] ), .Z(n_40159));
	notech_inv i_53100(.A(\to_acu2_0[26] ), .Z(n_40160));
	notech_inv i_53101(.A(\to_acu2_0[24] ), .Z(n_40161));
	notech_inv i_53102(.A(\to_acu2_0[25] ), .Z(n_40162));
	notech_inv i_53103(.A(\to_acu2_0[28] ), .Z(n_40163));
	notech_inv i_53104(.A(\to_acu2_0[16] ), .Z(n_40164));
	notech_inv i_53105(.A(\to_acu2_0[62] ), .Z(n_40165));
	notech_inv i_53106(.A(\to_acu2_0[69] ), .Z(n_40166));
	notech_inv i_53107(.A(\to_acu2_0[8] ), .Z(n_40167));
	notech_inv i_53108(.A(\to_acu2_0[11] ), .Z(n_40168));
	notech_inv i_53109(.A(\to_acu2_0[10] ), .Z(n_40169));
	notech_inv i_53110(.A(\to_acu2_0[9] ), .Z(n_40170));
	notech_inv i_53111(.A(fpu), .Z(n_40171));
	notech_inv i_53112(.A(in128[15]), .Z(n_40172));
	notech_inv i_53113(.A(in128[14]), .Z(n_40173));
	notech_inv i_53114(.A(in128[8]), .Z(n_40174));
	notech_inv i_53115(.A(in128[2]), .Z(n_40175));
	notech_inv i_53116(.A(in128[1]), .Z(n_40176));
	notech_inv i_53117(.A(mod_dec), .Z(n_40177));
	notech_inv i_53118(.A(sib_dec), .Z(n_40178));
	notech_inv i_53119(.A(\to_acu2_0[80] ), .Z(n_40179));
	notech_inv i_53120(.A(\to_acu2_0[79] ), .Z(n_40180));
	notech_inv i_53121(.A(\to_acu2_0[78] ), .Z(n_40181));
	notech_inv i_53122(.A(\to_acu2_0[77] ), .Z(n_40182));
	notech_inv i_53123(.A(\to_acu2_0[76] ), .Z(n_40183));
	notech_inv i_53124(.A(\to_acu2_0[73] ), .Z(n_40184));
	notech_inv i_53125(.A(\to_acu2_0[72] ), .Z(n_40185));
	notech_inv i_53126(.A(\to_acu2_0[68] ), .Z(n_40186));
	notech_inv i_53127(.A(\to_acu2_0[19] ), .Z(n_40187));
	notech_inv i_53128(.A(\nbus_12535[5] ), .Z(n_40188));
	notech_inv i_53129(.A(\nbus_12535[4] ), .Z(n_40189));
	notech_inv i_53130(.A(\nbus_12535[3] ), .Z(n_40190));
	notech_inv i_53131(.A(\nbus_12535[2] ), .Z(n_40191));
	notech_inv i_53132(.A(\nbus_12535[1] ), .Z(n_40192));
	notech_inv i_53133(.A(pg_fault), .Z(n_40193));
	notech_inv i_53134(.A(\nbus_12535[0] ), .Z(n_40194));
	notech_inv i_53135(.A(pc_req), .Z(n_40195));
	notech_inv i_53136(.A(in128[9]), .Z(n_40196));
	notech_inv i_53137(.A(n_57713), .Z(n_40197));
	notech_inv i_53138(.A(in128[3]), .Z(n_40198));
	notech_inv i_53139(.A(in128[4]), .Z(n_40199));
	notech_inv i_53140(.A(in128[5]), .Z(n_40200));
	notech_inv i_53141(.A(in128[6]), .Z(n_40201));
	notech_inv i_53142(.A(in128[7]), .Z(n_40202));
	notech_inv i_53143(.A(\to_acu2_0[75] ), .Z(n_40203));
	notech_inv i_53144(.A(\to_acu2_0[70] ), .Z(n_40204));
	notech_inv i_53145(.A(\to_acu2_0[71] ), .Z(n_40205));
	notech_inv i_53146(.A(in128[13]), .Z(n_40206));
	notech_inv i_53147(.A(in128[12]), .Z(n_40207));
	notech_inv i_53148(.A(in128[11]), .Z(n_40208));
	notech_inv i_53149(.A(\to_acu2_0[4] ), .Z(n_40209));
	notech_inv i_53150(.A(twobyte), .Z(n_40210));
	notech_inv i_53151(.A(\to_acu2_0[74] ), .Z(n_40211));
	notech_inv i_53152(.A(\to_acu2_0[3] ), .Z(n_40212));
	notech_inv i_53153(.A(in128[0]), .Z(n_40213));
	notech_inv i_53154(.A(\to_acu2_0[0] ), .Z(n_40214));
	notech_inv i_53155(.A(int_main), .Z(n_40215));
	deco8 i_deco_1(.in8({in128[7], in128[6], in128[5], in128[4], in128[3], in128
		[2], in128[1], in128[0]}), .indic({\to_acu2_0[80] , \to_acu2_0[79] 
		, \to_acu2_0[78] , \to_acu2_0[77] , \to_acu2_0[76] , \to_acu2_0[75] 
		, \to_acu2_0[74] , \to_acu2_0[73] , \to_acu2_0[72] , \to_acu2_0[71] 
		, \to_acu2_0[70] , \to_acu2_0[69] , \to_acu2_0[68] , \to_acu2_0[67] 
		, \to_acu2_0[66] , \to_acu2_0[65] , \to_acu2_0[64] , \to_acu2_0[63] 
		, \to_acu2_0[62] , \to_acu2_0[61] , \to_acu2_0[60] , \to_acu2_0[59] 
		, \to_acu2_0[58] , \to_acu2_0[57] , \to_acu2_0[56] , \to_acu2_0[55] 
		, \to_acu2_0[54] , \to_acu2_0[53] , \to_acu2_0[52] , \to_acu2_0[51] 
		, \to_acu2_0[50] , \to_acu2_0[49] , \to_acu2_0[48] , \to_acu2_0[47] 
		, \to_acu2_0[46] , \to_acu2_0[45] , \to_acu2_0[44] , \to_acu2_0[43] 
		, \to_acu2_0[42] , \to_acu2_0[41] , \to_acu2_0[40] , 
		UNCONNECTED_000, \to_acu2_0[38] , \to_acu2_0[37] , \to_acu2_0[36] 
		, \to_acu2_0[35] , \to_acu2_0[34] , \to_acu2_0[33] , \to_acu2_0[32] 
		, \to_acu2_0[31] , \to_acu2_0[30] , \to_acu2_0[29] , \to_acu2_0[28] 
		, \to_acu2_0[27] , \to_acu2_0[26] , \to_acu2_0[25] , \to_acu2_0[24] 
		, \to_acu2_0[23] , \to_acu2_0[22] , \to_acu2_0[21] , \to_acu2_0[20] 
		, \to_acu2_0[19] , \to_acu2_0[18] , \to_acu2_0[17] , \to_acu2_0[16] 
		, \to_acu2_0[15] , \to_acu2_0[14] , \to_acu2_0[13] , \to_acu2_0[12] 
		, \to_acu2_0[11] , \to_acu2_0[10] , \to_acu2_0[9] , \to_acu2_0[8] 
		}));
	deco_rm i_deco_3(.in8({in128[15], in128[14], in128[13], in128[12], 
		UNCONNECTED_001, n_57712, in128[9], in128[8]}), .indic({\to_acu2_0[7] 
		, \to_acu2_0[6] , \to_acu2_0[5] , \to_acu2_0[4] , \to_acu2_0[3] 
		, \to_acu2_0[2] , \to_acu2_0[1] , \to_acu2_0[0] }));
	udecox i_udeco(.op({in128[7], in128[6], in128[5], in128[4], in128[3], in128
		[2], in128[1], in128[0]}), .modrm({in128[15], in128[14], in128[
		13], in128[12], in128[11], n_57713, in128[9], in128[8]}), .twobyte
		(twobyte), .cpl(cpl), .adz(adz), .opz(opz), .udeco(udeco), .fpu(fpu
		), .emul(cr0[2]), .ipg_fault(ipg_fault));
	AWDP_partition_1 i_65676(.O0({\nbus_12535[5] , \nbus_12535[4] , \nbus_12535[3] 
		, \nbus_12535[2] , \nbus_12535[1] , \nbus_12535[0] }), .mod_dec(mod_dec
		), .sib_dec(sib_dec), .displc(displc), .imm_sz(imm_sz), .pfx_sz(pfx_sz
		), .twobyte(twobyte), .fpu(fpu));
endmodule
module AWDP_ADD_0(O0, opd, I0);

	output [31:0] O0;
	input [31:0] opd;
	input [31:0] I0;

	wire \opd[2] ;
	wire \opd[3] ;
	wire \opd[4] ;
	wire \opd[5] ;
	wire \opd[6] ;
	wire \opd[7] ;
	wire \opd[8] ;
	wire \opd[9] ;
	wire \opd[10] ;
	wire \opd[11] ;
	wire \opd[12] ;
	wire \opd[13] ;
	wire \opd[14] ;
	wire \opd[15] ;
	wire \opd[16] ;
	wire \opd[17] ;
	wire \opd[18] ;
	wire \opd[19] ;
	wire \opd[20] ;
	wire \opd[21] ;
	wire \opd[22] ;
	wire \opd[23] ;
	wire \opd[24] ;
	wire \opd[25] ;
	wire \opd[26] ;
	wire \opd[27] ;
	wire \opd[28] ;
	wire \opd[29] ;
	wire \opd[30] ;
	wire \opd[31] ;


	assign O0[0] = opd[0];
	assign O0[1] = opd[1];
	assign \opd[2]  = opd[2];
	assign \opd[3]  = opd[3];
	assign \opd[4]  = opd[4];
	assign \opd[5]  = opd[5];
	assign \opd[6]  = opd[6];
	assign \opd[7]  = opd[7];
	assign \opd[8]  = opd[8];
	assign \opd[9]  = opd[9];
	assign \opd[10]  = opd[10];
	assign \opd[11]  = opd[11];
	assign \opd[12]  = opd[12];
	assign \opd[13]  = opd[13];
	assign \opd[14]  = opd[14];
	assign \opd[15]  = opd[15];
	assign \opd[16]  = opd[16];
	assign \opd[17]  = opd[17];
	assign \opd[18]  = opd[18];
	assign \opd[19]  = opd[19];
	assign \opd[20]  = opd[20];
	assign \opd[21]  = opd[21];
	assign \opd[22]  = opd[22];
	assign \opd[23]  = opd[23];
	assign \opd[24]  = opd[24];
	assign \opd[25]  = opd[25];
	assign \opd[26]  = opd[26];
	assign \opd[27]  = opd[27];
	assign \opd[28]  = opd[28];
	assign \opd[29]  = opd[29];
	assign \opd[30]  = opd[30];
	assign \opd[31]  = opd[31];

	notech_ha2 i_29(.A(\opd[31] ), .B(n_354), .Z(O0[31]));
	notech_ha2 i_28(.A(\opd[30] ), .B(n_352), .Z(O0[30]), .CO(n_354));
	notech_ha2 i_27(.A(\opd[29] ), .B(n_341), .Z(O0[29]), .CO(n_352));
	notech_fa2 i_26(.A(I0[28]), .B(n_339), .CI(\opd[28] ), .Z(O0[28]), .CO(n_341
		));
	notech_fa2 i_25(.A(I0[27]), .B(n_337), .CI(\opd[27] ), .Z(O0[27]), .CO(n_339
		));
	notech_fa2 i_24(.A(I0[26]), .B(n_335), .CI(\opd[26] ), .Z(O0[26]), .CO(n_337
		));
	notech_fa2 i_23(.A(I0[25]), .B(n_333), .CI(\opd[25] ), .Z(O0[25]), .CO(n_335
		));
	notech_fa2 i_22(.A(I0[24]), .B(n_331), .CI(\opd[24] ), .Z(O0[24]), .CO(n_333
		));
	notech_fa2 i_21(.A(I0[23]), .B(n_329), .CI(\opd[23] ), .Z(O0[23]), .CO(n_331
		));
	notech_fa2 i_20(.A(I0[22]), .B(n_327), .CI(\opd[22] ), .Z(O0[22]), .CO(n_329
		));
	notech_fa2 i_19(.A(I0[21]), .B(n_325), .CI(\opd[21] ), .Z(O0[21]), .CO(n_327
		));
	notech_fa2 i_18(.A(I0[20]), .B(n_323), .CI(\opd[20] ), .Z(O0[20]), .CO(n_325
		));
	notech_fa2 i_17(.A(I0[19]), .B(n_321), .CI(\opd[19] ), .Z(O0[19]), .CO(n_323
		));
	notech_fa2 i_16(.A(I0[18]), .B(n_319), .CI(\opd[18] ), .Z(O0[18]), .CO(n_321
		));
	notech_fa2 i_15(.A(I0[17]), .B(n_317), .CI(\opd[17] ), .Z(O0[17]), .CO(n_319
		));
	notech_fa2 i_14(.A(I0[16]), .B(n_315), .CI(\opd[16] ), .Z(O0[16]), .CO(n_317
		));
	notech_fa2 i_13(.A(I0[15]), .B(n_313), .CI(\opd[15] ), .Z(O0[15]), .CO(n_315
		));
	notech_fa2 i_12(.A(I0[14]), .B(n_311), .CI(\opd[14] ), .Z(O0[14]), .CO(n_313
		));
	notech_fa2 i_11(.A(I0[13]), .B(n_309), .CI(\opd[13] ), .Z(O0[13]), .CO(n_311
		));
	notech_fa2 i_10(.A(I0[12]), .B(n_307), .CI(\opd[12] ), .Z(O0[12]), .CO(n_309
		));
	notech_fa2 i_9(.A(I0[11]), .B(n_305), .CI(\opd[11] ), .Z(O0[11]), .CO(n_307
		));
	notech_fa2 i_8(.A(I0[10]), .B(n_303), .CI(\opd[10] ), .Z(O0[10]), .CO(n_305
		));
	notech_fa2 i_7(.A(I0[9]), .B(n_301), .CI(\opd[9] ), .Z(O0[9]), .CO(n_303
		));
	notech_fa2 i_6(.A(I0[8]), .B(n_299), .CI(\opd[8] ), .Z(O0[8]), .CO(n_301
		));
	notech_fa2 i_5(.A(I0[7]), .B(n_297), .CI(\opd[7] ), .Z(O0[7]), .CO(n_299
		));
	notech_fa2 i_4(.A(I0[6]), .B(n_295), .CI(\opd[6] ), .Z(O0[6]), .CO(n_297
		));
	notech_fa2 i_3(.A(I0[5]), .B(n_293), .CI(\opd[5] ), .Z(O0[5]), .CO(n_295
		));
	notech_fa2 i_2(.A(I0[4]), .B(n_291), .CI(\opd[4] ), .Z(O0[4]), .CO(n_293
		));
	notech_fa2 i_1(.A(I0[3]), .B(n_350), .CI(\opd[3] ), .Z(O0[3]), .CO(n_291
		));
	notech_ha2 i_0(.A(I0[2]), .B(\opd[2] ), .Z(O0[2]), .CO(n_350));
endmodule
module AWDP_ADD_100(O0, opb, I0);

	output [32:0] O0;
	input [31:0] opb;
	input [31:0] I0;




	notech_inv i_10767(.A(n_57116), .Z(n_57117));
	notech_inv i_10766(.A(I0[18]), .Z(n_57116));
	notech_fa2 i_31(.A(I0[18]), .B(n_354), .CI(opb[31]), .Z(O0[31]), .CO(O0[
		32]));
	notech_fa2 i_30(.A(I0[18]), .B(n_352), .CI(opb[30]), .Z(O0[30]), .CO(n_354
		));
	notech_fa2 i_29(.A(I0[18]), .B(n_350), .CI(opb[29]), .Z(O0[29]), .CO(n_352
		));
	notech_fa2 i_28(.A(I0[18]), .B(n_348), .CI(opb[28]), .Z(O0[28]), .CO(n_350
		));
	notech_fa2 i_27(.A(I0[18]), .B(n_346), .CI(opb[27]), .Z(O0[27]), .CO(n_348
		));
	notech_fa2 i_26(.A(I0[18]), .B(n_344), .CI(opb[26]), .Z(O0[26]), .CO(n_346
		));
	notech_fa2 i_25(.A(I0[18]), .B(n_342), .CI(opb[25]), .Z(O0[25]), .CO(n_344
		));
	notech_fa2 i_24(.A(I0[18]), .B(n_340), .CI(opb[24]), .Z(O0[24]), .CO(n_342
		));
	notech_fa2 i_23(.A(I0[18]), .B(n_338), .CI(opb[23]), .Z(O0[23]), .CO(n_340
		));
	notech_fa2 i_22(.A(I0[18]), .B(n_336), .CI(opb[22]), .Z(O0[22]), .CO(n_338
		));
	notech_fa2 i_21(.A(I0[18]), .B(n_334), .CI(opb[21]), .Z(O0[21]), .CO(n_336
		));
	notech_fa2 i_20(.A(I0[18]), .B(n_332), .CI(opb[20]), .Z(O0[20]), .CO(n_334
		));
	notech_fa2 i_19(.A(I0[18]), .B(n_330), .CI(opb[19]), .Z(O0[19]), .CO(n_332
		));
	notech_fa2 i_18(.A(I0[18]), .B(n_328), .CI(opb[18]), .Z(O0[18]), .CO(n_330
		));
	notech_fa2 i_17(.A(I0[18]), .B(n_326), .CI(opb[17]), .Z(O0[17]), .CO(n_328
		));
	notech_fa2 i_16(.A(n_57117), .B(n_324), .CI(opb[16]), .Z(O0[16]), .CO(n_326
		));
	notech_fa2 i_15(.A(n_57117), .B(n_322), .CI(opb[15]), .Z(O0[15]), .CO(n_324
		));
	notech_fa2 i_14(.A(n_57117), .B(n_320), .CI(opb[14]), .Z(O0[14]), .CO(n_322
		));
	notech_fa2 i_13(.A(n_57117), .B(n_318), .CI(opb[13]), .Z(O0[13]), .CO(n_320
		));
	notech_fa2 i_12(.A(n_57117), .B(n_316), .CI(opb[12]), .Z(O0[12]), .CO(n_318
		));
	notech_fa2 i_11(.A(n_57117), .B(n_314), .CI(opb[11]), .Z(O0[11]), .CO(n_316
		));
	notech_fa2 i_10(.A(n_57117), .B(n_312), .CI(opb[10]), .Z(O0[10]), .CO(n_314
		));
	notech_fa2 i_9(.A(n_57117), .B(n_310), .CI(opb[9]), .Z(O0[9]), .CO(n_312
		));
	notech_fa2 i_8(.A(n_57117), .B(n_308), .CI(opb[8]), .Z(O0[8]), .CO(n_310
		));
	notech_fa2 i_7(.A(n_57117), .B(n_306), .CI(opb[7]), .Z(O0[7]), .CO(n_308
		));
	notech_fa2 i_6(.A(n_57117), .B(n_304), .CI(opb[6]), .Z(O0[6]), .CO(n_306
		));
	notech_fa2 i_5(.A(n_57117), .B(n_302), .CI(opb[5]), .Z(O0[5]), .CO(n_304
		));
	notech_fa2 i_4(.A(n_57117), .B(n_300), .CI(opb[4]), .Z(O0[4]), .CO(n_302
		));
	notech_fa2 i_3(.A(n_57117), .B(n_298), .CI(opb[3]), .Z(O0[3]), .CO(n_300
		));
	notech_fa2 i_2(.A(n_57117), .B(n_296), .CI(opb[2]), .Z(O0[2]), .CO(n_298
		));
	notech_fa2 i_1(.A(I0[1]), .B(n_361), .CI(opb[1]), .Z(O0[1]), .CO(n_296)
		);
	notech_ha2 i_0(.A(opb[0]), .B(I0[0]), .Z(O0[0]), .CO(n_361));
endmodule
module AWDP_ADD_122(O0, opa, opd);
    output [32:0] O0;
    input [31:0] opa;
    input [31:0] opd;
    // Line 599
    wire [32:0] O0;
    // Line 599
    wire [32:0] N70;

    // Line 599
    assign O0 = N70;
    // Line 599
    assign N70 = opa + opd;
endmodule

module AWDP_ADD_13(O0, regs_7, opd);
    output [31:0] O0;
    input [31:0] regs_7;
    input [31:0] opd;
    // Line 348
    wire [31:0] O0;
    // Line 520
    wire [31:0] N82;

    // Line 348
    assign O0 = N82;
    // Line 520
    assign N82 = regs_7 + opd;
endmodule

module AWDP_ADD_136(O0, opa, I0);

	output [16:0] O0;
	input [15:0] opa;
	input [15:0] I0;




	notech_fa2 i_15(.A(I0[13]), .B(n_178), .CI(opa[15]), .Z(O0[15]), .CO(O0[
		16]));
	notech_fa2 i_14(.A(I0[13]), .B(n_176), .CI(opa[14]), .Z(O0[14]), .CO(n_178
		));
	notech_fa2 i_13(.A(I0[13]), .B(n_174), .CI(opa[13]), .Z(O0[13]), .CO(n_176
		));
	notech_fa2 i_12(.A(I0[13]), .B(n_172), .CI(opa[12]), .Z(O0[12]), .CO(n_174
		));
	notech_fa2 i_11(.A(I0[13]), .B(n_170), .CI(opa[11]), .Z(O0[11]), .CO(n_172
		));
	notech_fa2 i_10(.A(I0[13]), .B(n_168), .CI(opa[10]), .Z(O0[10]), .CO(n_170
		));
	notech_fa2 i_9(.A(I0[13]), .B(n_166), .CI(opa[9]), .Z(O0[9]), .CO(n_168)
		);
	notech_fa2 i_8(.A(I0[13]), .B(n_164), .CI(opa[8]), .Z(O0[8]), .CO(n_166)
		);
	notech_fa2 i_7(.A(I0[13]), .B(n_162), .CI(opa[7]), .Z(O0[7]), .CO(n_164)
		);
	notech_fa2 i_6(.A(I0[13]), .B(n_160), .CI(opa[6]), .Z(O0[6]), .CO(n_162)
		);
	notech_fa2 i_5(.A(I0[13]), .B(n_158), .CI(opa[5]), .Z(O0[5]), .CO(n_160)
		);
	notech_fa2 i_4(.A(I0[13]), .B(n_156), .CI(opa[4]), .Z(O0[4]), .CO(n_158)
		);
	notech_fa2 i_3(.A(I0[13]), .B(n_154), .CI(opa[3]), .Z(O0[3]), .CO(n_156)
		);
	notech_fa2 i_2(.A(I0[13]), .B(n_152), .CI(opa[2]), .Z(O0[2]), .CO(n_154)
		);
	notech_fa2 i_1(.A(I0[1]), .B(n_185), .CI(opa[1]), .Z(O0[1]), .CO(n_152)
		);
	notech_ha2 i_0(.A(opa[0]), .B(I0[0]), .Z(O0[0]), .CO(n_185));
endmodule
module AWDP_ADD_139(O0, opa, opd);
    output [16:0] O0;
    input [15:0] opa;
    input [15:0] opd;
    // Line 600
    wire [16:0] N109;
    // Line 600
    wire [16:0] O0;

    // Line 600
    assign N109 = opa + opd;
    // Line 600
    assign O0 = N109;
endmodule

module AWDP_ADD_14(O0, regs_4, calc_sz);
    output [31:0] O0;
    input [31:0] regs_4;
    input [2:0] calc_sz;
    // Line 348
    wire [31:0] O0;
    // Line 470
    wire [31:0] N121;

    // Line 348
    assign O0 = N121;
    // Line 470
    assign N121 = regs_4 + calc_sz;
endmodule

module AWDP_ADD_181(O0, idtr, I0);

	output [31:0] O0;
	input [31:0] idtr;
	input [18:0] I0;

	wire \idtr[3] ;
	wire \idtr[4] ;
	wire \idtr[5] ;
	wire \idtr[6] ;
	wire \idtr[7] ;
	wire \idtr[8] ;
	wire \idtr[9] ;
	wire \idtr[10] ;
	wire \idtr[11] ;
	wire \idtr[12] ;
	wire \idtr[13] ;
	wire \idtr[14] ;
	wire \idtr[15] ;
	wire \idtr[16] ;
	wire \idtr[17] ;
	wire \idtr[18] ;
	wire \idtr[19] ;
	wire \idtr[20] ;
	wire \idtr[21] ;
	wire \idtr[22] ;
	wire \idtr[23] ;
	wire \idtr[24] ;
	wire \idtr[25] ;
	wire \idtr[26] ;
	wire \idtr[27] ;
	wire \idtr[28] ;
	wire \idtr[29] ;
	wire \idtr[30] ;
	wire \idtr[31] ;


	assign O0[0] = idtr[0];
	assign O0[1] = idtr[1];
	assign O0[2] = idtr[2];
	assign \idtr[3]  = idtr[3];
	assign \idtr[4]  = idtr[4];
	assign \idtr[5]  = idtr[5];
	assign \idtr[6]  = idtr[6];
	assign \idtr[7]  = idtr[7];
	assign \idtr[8]  = idtr[8];
	assign \idtr[9]  = idtr[9];
	assign \idtr[10]  = idtr[10];
	assign \idtr[11]  = idtr[11];
	assign \idtr[12]  = idtr[12];
	assign \idtr[13]  = idtr[13];
	assign \idtr[14]  = idtr[14];
	assign \idtr[15]  = idtr[15];
	assign \idtr[16]  = idtr[16];
	assign \idtr[17]  = idtr[17];
	assign \idtr[18]  = idtr[18];
	assign \idtr[19]  = idtr[19];
	assign \idtr[20]  = idtr[20];
	assign \idtr[21]  = idtr[21];
	assign \idtr[22]  = idtr[22];
	assign \idtr[23]  = idtr[23];
	assign \idtr[24]  = idtr[24];
	assign \idtr[25]  = idtr[25];
	assign \idtr[26]  = idtr[26];
	assign \idtr[27]  = idtr[27];
	assign \idtr[28]  = idtr[28];
	assign \idtr[29]  = idtr[29];
	assign \idtr[30]  = idtr[30];
	assign \idtr[31]  = idtr[31];

	notech_ha2 i_28(.A(\idtr[31] ), .B(n_346), .Z(O0[31]));
	notech_ha2 i_27(.A(\idtr[30] ), .B(n_344), .Z(O0[30]), .CO(n_346));
	notech_ha2 i_26(.A(\idtr[29] ), .B(n_342), .Z(O0[29]), .CO(n_344));
	notech_ha2 i_25(.A(\idtr[28] ), .B(n_340), .Z(O0[28]), .CO(n_342));
	notech_ha2 i_24(.A(\idtr[27] ), .B(n_338), .Z(O0[27]), .CO(n_340));
	notech_ha2 i_23(.A(\idtr[26] ), .B(n_336), .Z(O0[26]), .CO(n_338));
	notech_ha2 i_22(.A(\idtr[25] ), .B(n_334), .Z(O0[25]), .CO(n_336));
	notech_ha2 i_21(.A(\idtr[24] ), .B(n_332), .Z(O0[24]), .CO(n_334));
	notech_ha2 i_20(.A(\idtr[23] ), .B(n_330), .Z(O0[23]), .CO(n_332));
	notech_ha2 i_19(.A(\idtr[22] ), .B(n_328), .Z(O0[22]), .CO(n_330));
	notech_ha2 i_18(.A(\idtr[21] ), .B(n_326), .Z(O0[21]), .CO(n_328));
	notech_ha2 i_17(.A(\idtr[20] ), .B(n_324), .Z(O0[20]), .CO(n_326));
	notech_ha2 i_16(.A(\idtr[19] ), .B(n_293), .Z(O0[19]), .CO(n_324));
	notech_fa2 i_15(.A(I0[18]), .B(n_291), .CI(\idtr[18] ), .Z(O0[18]), .CO(n_293
		));
	notech_fa2 i_14(.A(I0[17]), .B(n_289), .CI(\idtr[17] ), .Z(O0[17]), .CO(n_291
		));
	notech_fa2 i_13(.A(I0[16]), .B(n_287), .CI(\idtr[16] ), .Z(O0[16]), .CO(n_289
		));
	notech_fa2 i_12(.A(I0[15]), .B(n_285), .CI(\idtr[15] ), .Z(O0[15]), .CO(n_287
		));
	notech_fa2 i_11(.A(I0[14]), .B(n_283), .CI(\idtr[14] ), .Z(O0[14]), .CO(n_285
		));
	notech_fa2 i_10(.A(I0[13]), .B(n_281), .CI(\idtr[13] ), .Z(O0[13]), .CO(n_283
		));
	notech_fa2 i_9(.A(I0[12]), .B(n_279), .CI(\idtr[12] ), .Z(O0[12]), .CO(n_281
		));
	notech_fa2 i_8(.A(I0[11]), .B(n_277), .CI(\idtr[11] ), .Z(O0[11]), .CO(n_279
		));
	notech_fa2 i_7(.A(I0[10]), .B(n_275), .CI(\idtr[10] ), .Z(O0[10]), .CO(n_277
		));
	notech_fa2 i_6(.A(I0[9]), .B(n_273), .CI(\idtr[9] ), .Z(O0[9]), .CO(n_275
		));
	notech_fa2 i_5(.A(I0[8]), .B(n_271), .CI(\idtr[8] ), .Z(O0[8]), .CO(n_273
		));
	notech_fa2 i_4(.A(I0[7]), .B(n_269), .CI(\idtr[7] ), .Z(O0[7]), .CO(n_271
		));
	notech_fa2 i_3(.A(I0[6]), .B(n_267), .CI(\idtr[6] ), .Z(O0[6]), .CO(n_269
		));
	notech_fa2 i_2(.A(I0[5]), .B(n_265), .CI(\idtr[5] ), .Z(O0[5]), .CO(n_267
		));
	notech_fa2 i_1(.A(I0[4]), .B(n_322), .CI(\idtr[4] ), .Z(O0[4]), .CO(n_265
		));
	notech_ha2 i_0(.A(\idtr[3] ), .B(I0[3]), .Z(O0[3]), .CO(n_322));
endmodule
module AWDP_ADD_185(O0, opb, I0);

	output [31:0] O0;
	input [31:0] opb;
	input [31:0] I0;




	notech_ha2 i_31(.A(opb[31]), .B(n_400), .Z(O0[31]));
	notech_ha2 i_30(.A(opb[30]), .B(n_398), .Z(O0[30]), .CO(n_400));
	notech_ha2 i_29(.A(opb[29]), .B(n_396), .Z(O0[29]), .CO(n_398));
	notech_ha2 i_28(.A(opb[28]), .B(n_394), .Z(O0[28]), .CO(n_396));
	notech_ha2 i_27(.A(opb[27]), .B(n_392), .Z(O0[27]), .CO(n_394));
	notech_ha2 i_26(.A(opb[26]), .B(n_390), .Z(O0[26]), .CO(n_392));
	notech_ha2 i_25(.A(opb[25]), .B(n_388), .Z(O0[25]), .CO(n_390));
	notech_ha2 i_24(.A(opb[24]), .B(n_386), .Z(O0[24]), .CO(n_388));
	notech_ha2 i_23(.A(opb[23]), .B(n_384), .Z(O0[23]), .CO(n_386));
	notech_ha2 i_22(.A(opb[22]), .B(n_382), .Z(O0[22]), .CO(n_384));
	notech_ha2 i_21(.A(opb[21]), .B(n_380), .Z(O0[21]), .CO(n_382));
	notech_ha2 i_20(.A(opb[20]), .B(n_378), .Z(O0[20]), .CO(n_380));
	notech_ha2 i_19(.A(opb[19]), .B(n_376), .Z(O0[19]), .CO(n_378));
	notech_ha2 i_18(.A(opb[18]), .B(n_374), .Z(O0[18]), .CO(n_376));
	notech_ha2 i_17(.A(opb[17]), .B(n_372), .Z(O0[17]), .CO(n_374));
	notech_ha2 i_16(.A(opb[16]), .B(n_370), .Z(O0[16]), .CO(n_372));
	notech_ha2 i_15(.A(opb[15]), .B(n_368), .Z(O0[15]), .CO(n_370));
	notech_ha2 i_14(.A(opb[14]), .B(n_366), .Z(O0[14]), .CO(n_368));
	notech_ha2 i_13(.A(opb[13]), .B(n_364), .Z(O0[13]), .CO(n_366));
	notech_ha2 i_12(.A(opb[12]), .B(n_362), .Z(O0[12]), .CO(n_364));
	notech_ha2 i_11(.A(opb[11]), .B(n_360), .Z(O0[11]), .CO(n_362));
	notech_ha2 i_10(.A(opb[10]), .B(n_358), .Z(O0[10]), .CO(n_360));
	notech_ha2 i_9(.A(opb[9]), .B(n_356), .Z(O0[9]), .CO(n_358));
	notech_ha2 i_8(.A(opb[8]), .B(n_303), .Z(O0[8]), .CO(n_356));
	notech_fa2 i_7(.A(I0[7]), .B(n_301), .CI(opb[7]), .Z(O0[7]), .CO(n_303)
		);
	notech_fa2 i_6(.A(I0[6]), .B(n_299), .CI(opb[6]), .Z(O0[6]), .CO(n_301)
		);
	notech_fa2 i_5(.A(I0[5]), .B(n_297), .CI(opb[5]), .Z(O0[5]), .CO(n_299)
		);
	notech_fa2 i_4(.A(I0[4]), .B(n_295), .CI(opb[4]), .Z(O0[4]), .CO(n_297)
		);
	notech_fa2 i_3(.A(I0[3]), .B(n_293), .CI(opb[3]), .Z(O0[3]), .CO(n_295)
		);
	notech_fa2 i_2(.A(I0[2]), .B(n_291), .CI(opb[2]), .Z(O0[2]), .CO(n_293)
		);
	notech_fa2 i_1(.A(I0[1]), .B(n_354), .CI(opb[1]), .Z(O0[1]), .CO(n_291)
		);
	notech_ha2 i_0(.A(I0[0]), .B(opb[0]), .Z(O0[0]), .CO(n_354));
endmodule
module AWDP_ADD_194(O0, opa, opd);
    output [8:0] O0;
    input [7:0] opa;
    input [7:0] opd;
    // Line 601
    wire [8:0] N154;
    // Line 601
    wire [8:0] O0;

    // Line 601
    assign N154 = opa + opd;
    // Line 601
    assign O0 = N154;
endmodule

module AWDP_ADD_195(O0, opc, I0);
    output [31:0] O0;
    input [31:0] opc;
    input [31:0] I0;
    // Line 1006
    wire [31:0] N167;
    // Line 1006
    wire [31:0] O0;

    // Line 1006
    assign N167 = opc + I0;
    // Line 1006
    assign O0 = N167;
endmodule

module AWDP_ADD_198(O0, I0, add_len_pc);
    output [31:0] O0;
    input [31:0] I0;
    input [31:0] add_len_pc;
    // Line 879
    wire [31:0] N190;
    // Line 386
    wire [31:0] O0;

    // Line 879
    assign N190 = I0 + add_len_pc;
    // Line 386
    assign O0 = N190;
endmodule

module AWDP_ADD_207(O0, regs_6, opd);
    output [31:0] O0;
    input [31:0] regs_6;
    input [31:0] opd;
    // Line 348
    wire [31:0] O0;
    // Line 520
    wire [31:0] N199;

    // Line 348
    assign O0 = N199;
    // Line 520
    assign N199 = regs_6 + opd;
endmodule

module AWDP_ADD_22(O0, gdtr, I0);

	output [31:0] O0;
	input [31:0] gdtr;
	input [31:0] I0;

	wire \gdtr[1] ;
	wire \gdtr[2] ;
	wire \gdtr[3] ;
	wire \gdtr[4] ;
	wire \gdtr[5] ;
	wire \gdtr[6] ;
	wire \gdtr[7] ;
	wire \gdtr[8] ;
	wire \gdtr[9] ;
	wire \gdtr[10] ;
	wire \gdtr[11] ;
	wire \gdtr[12] ;
	wire \gdtr[13] ;
	wire \gdtr[14] ;
	wire \gdtr[15] ;
	wire \gdtr[16] ;
	wire \gdtr[17] ;
	wire \gdtr[18] ;
	wire \gdtr[19] ;
	wire \gdtr[20] ;
	wire \gdtr[21] ;
	wire \gdtr[22] ;
	wire \gdtr[23] ;
	wire \gdtr[24] ;
	wire \gdtr[25] ;
	wire \gdtr[26] ;
	wire \gdtr[27] ;
	wire \gdtr[28] ;
	wire \gdtr[29] ;
	wire \gdtr[30] ;
	wire \gdtr[31] ;


	assign O0[0] = gdtr[0];
	assign \gdtr[1]  = gdtr[1];
	assign \gdtr[2]  = gdtr[2];
	assign \gdtr[3]  = gdtr[3];
	assign \gdtr[4]  = gdtr[4];
	assign \gdtr[5]  = gdtr[5];
	assign \gdtr[6]  = gdtr[6];
	assign \gdtr[7]  = gdtr[7];
	assign \gdtr[8]  = gdtr[8];
	assign \gdtr[9]  = gdtr[9];
	assign \gdtr[10]  = gdtr[10];
	assign \gdtr[11]  = gdtr[11];
	assign \gdtr[12]  = gdtr[12];
	assign \gdtr[13]  = gdtr[13];
	assign \gdtr[14]  = gdtr[14];
	assign \gdtr[15]  = gdtr[15];
	assign \gdtr[16]  = gdtr[16];
	assign \gdtr[17]  = gdtr[17];
	assign \gdtr[18]  = gdtr[18];
	assign \gdtr[19]  = gdtr[19];
	assign \gdtr[20]  = gdtr[20];
	assign \gdtr[21]  = gdtr[21];
	assign \gdtr[22]  = gdtr[22];
	assign \gdtr[23]  = gdtr[23];
	assign \gdtr[24]  = gdtr[24];
	assign \gdtr[25]  = gdtr[25];
	assign \gdtr[26]  = gdtr[26];
	assign \gdtr[27]  = gdtr[27];
	assign \gdtr[28]  = gdtr[28];
	assign \gdtr[29]  = gdtr[29];
	assign \gdtr[30]  = gdtr[30];
	assign \gdtr[31]  = gdtr[31];

	notech_fa2 i_30(.A(I0[31]), .B(n_347), .CI(\gdtr[31] ), .Z(O0[31]));
	notech_fa2 i_29(.A(I0[30]), .B(n_345), .CI(\gdtr[30] ), .Z(O0[30]), .CO(n_347
		));
	notech_fa2 i_28(.A(I0[29]), .B(n_343), .CI(\gdtr[29] ), .Z(O0[29]), .CO(n_345
		));
	notech_fa2 i_27(.A(I0[28]), .B(n_341), .CI(\gdtr[28] ), .Z(O0[28]), .CO(n_343
		));
	notech_fa2 i_26(.A(I0[27]), .B(n_339), .CI(\gdtr[27] ), .Z(O0[27]), .CO(n_341
		));
	notech_fa2 i_25(.A(I0[26]), .B(n_337), .CI(\gdtr[26] ), .Z(O0[26]), .CO(n_339
		));
	notech_fa2 i_24(.A(I0[25]), .B(n_335), .CI(\gdtr[25] ), .Z(O0[25]), .CO(n_337
		));
	notech_fa2 i_23(.A(I0[24]), .B(n_333), .CI(\gdtr[24] ), .Z(O0[24]), .CO(n_335
		));
	notech_fa2 i_22(.A(I0[23]), .B(n_331), .CI(\gdtr[23] ), .Z(O0[23]), .CO(n_333
		));
	notech_fa2 i_21(.A(I0[22]), .B(n_329), .CI(\gdtr[22] ), .Z(O0[22]), .CO(n_331
		));
	notech_fa2 i_20(.A(I0[21]), .B(n_327), .CI(\gdtr[21] ), .Z(O0[21]), .CO(n_329
		));
	notech_fa2 i_19(.A(I0[20]), .B(n_325), .CI(\gdtr[20] ), .Z(O0[20]), .CO(n_327
		));
	notech_fa2 i_18(.A(I0[19]), .B(n_323), .CI(\gdtr[19] ), .Z(O0[19]), .CO(n_325
		));
	notech_fa2 i_17(.A(I0[18]), .B(n_321), .CI(\gdtr[18] ), .Z(O0[18]), .CO(n_323
		));
	notech_fa2 i_16(.A(I0[17]), .B(n_319), .CI(\gdtr[17] ), .Z(O0[17]), .CO(n_321
		));
	notech_fa2 i_15(.A(I0[16]), .B(n_317), .CI(\gdtr[16] ), .Z(O0[16]), .CO(n_319
		));
	notech_fa2 i_14(.A(I0[15]), .B(n_315), .CI(\gdtr[15] ), .Z(O0[15]), .CO(n_317
		));
	notech_fa2 i_13(.A(I0[14]), .B(n_313), .CI(\gdtr[14] ), .Z(O0[14]), .CO(n_315
		));
	notech_fa2 i_12(.A(I0[13]), .B(n_311), .CI(\gdtr[13] ), .Z(O0[13]), .CO(n_313
		));
	notech_fa2 i_11(.A(I0[12]), .B(n_309), .CI(\gdtr[12] ), .Z(O0[12]), .CO(n_311
		));
	notech_fa2 i_10(.A(I0[11]), .B(n_307), .CI(\gdtr[11] ), .Z(O0[11]), .CO(n_309
		));
	notech_fa2 i_9(.A(I0[10]), .B(n_305), .CI(\gdtr[10] ), .Z(O0[10]), .CO(n_307
		));
	notech_fa2 i_8(.A(I0[9]), .B(n_303), .CI(\gdtr[9] ), .Z(O0[9]), .CO(n_305
		));
	notech_fa2 i_7(.A(I0[8]), .B(n_301), .CI(\gdtr[8] ), .Z(O0[8]), .CO(n_303
		));
	notech_fa2 i_6(.A(I0[7]), .B(n_299), .CI(\gdtr[7] ), .Z(O0[7]), .CO(n_301
		));
	notech_fa2 i_5(.A(I0[6]), .B(n_297), .CI(\gdtr[6] ), .Z(O0[6]), .CO(n_299
		));
	notech_fa2 i_4(.A(I0[5]), .B(n_295), .CI(\gdtr[5] ), .Z(O0[5]), .CO(n_297
		));
	notech_fa2 i_3(.A(I0[4]), .B(n_293), .CI(\gdtr[4] ), .Z(O0[4]), .CO(n_295
		));
	notech_fa2 i_2(.A(I0[3]), .B(n_354), .CI(\gdtr[3] ), .Z(O0[3]), .CO(n_293
		));
	notech_ha2 i_1(.A(\gdtr[2] ), .B(\gdtr[1] ), .Z(O0[2]), .CO(n_354));
	notech_inv i_0(.A(\gdtr[1] ), .Z(O0[1]));
endmodule
module AWDP_ADD_238(O0, gdtr, I0);

	output [31:0] O0;
	input [31:0] gdtr;
	input [15:0] I0;

	wire \gdtr[1] ;
	wire \gdtr[2] ;
	wire \gdtr[3] ;
	wire \gdtr[4] ;
	wire \gdtr[5] ;
	wire \gdtr[6] ;
	wire \gdtr[7] ;
	wire \gdtr[8] ;
	wire \gdtr[9] ;
	wire \gdtr[10] ;
	wire \gdtr[11] ;
	wire \gdtr[12] ;
	wire \gdtr[13] ;
	wire \gdtr[14] ;
	wire \gdtr[15] ;
	wire \gdtr[16] ;
	wire \gdtr[17] ;
	wire \gdtr[18] ;
	wire \gdtr[19] ;
	wire \gdtr[20] ;
	wire \gdtr[21] ;
	wire \gdtr[22] ;
	wire \gdtr[23] ;
	wire \gdtr[24] ;
	wire \gdtr[25] ;
	wire \gdtr[26] ;
	wire \gdtr[27] ;
	wire \gdtr[28] ;
	wire \gdtr[29] ;
	wire \gdtr[30] ;
	wire \gdtr[31] ;


	assign O0[0] = gdtr[0];
	assign \gdtr[1]  = gdtr[1];
	assign \gdtr[2]  = gdtr[2];
	assign \gdtr[3]  = gdtr[3];
	assign \gdtr[4]  = gdtr[4];
	assign \gdtr[5]  = gdtr[5];
	assign \gdtr[6]  = gdtr[6];
	assign \gdtr[7]  = gdtr[7];
	assign \gdtr[8]  = gdtr[8];
	assign \gdtr[9]  = gdtr[9];
	assign \gdtr[10]  = gdtr[10];
	assign \gdtr[11]  = gdtr[11];
	assign \gdtr[12]  = gdtr[12];
	assign \gdtr[13]  = gdtr[13];
	assign \gdtr[14]  = gdtr[14];
	assign \gdtr[15]  = gdtr[15];
	assign \gdtr[16]  = gdtr[16];
	assign \gdtr[17]  = gdtr[17];
	assign \gdtr[18]  = gdtr[18];
	assign \gdtr[19]  = gdtr[19];
	assign \gdtr[20]  = gdtr[20];
	assign \gdtr[21]  = gdtr[21];
	assign \gdtr[22]  = gdtr[22];
	assign \gdtr[23]  = gdtr[23];
	assign \gdtr[24]  = gdtr[24];
	assign \gdtr[25]  = gdtr[25];
	assign \gdtr[26]  = gdtr[26];
	assign \gdtr[27]  = gdtr[27];
	assign \gdtr[28]  = gdtr[28];
	assign \gdtr[29]  = gdtr[29];
	assign \gdtr[30]  = gdtr[30];
	assign \gdtr[31]  = gdtr[31];

	notech_ha2 i_30(.A(\gdtr[31] ), .B(n_352), .Z(O0[31]));
	notech_ha2 i_29(.A(\gdtr[30] ), .B(n_350), .Z(O0[30]), .CO(n_352));
	notech_ha2 i_28(.A(\gdtr[29] ), .B(n_348), .Z(O0[29]), .CO(n_350));
	notech_ha2 i_27(.A(\gdtr[28] ), .B(n_346), .Z(O0[28]), .CO(n_348));
	notech_ha2 i_26(.A(\gdtr[27] ), .B(n_344), .Z(O0[27]), .CO(n_346));
	notech_ha2 i_25(.A(\gdtr[26] ), .B(n_342), .Z(O0[26]), .CO(n_344));
	notech_ha2 i_24(.A(\gdtr[25] ), .B(n_340), .Z(O0[25]), .CO(n_342));
	notech_ha2 i_23(.A(\gdtr[24] ), .B(n_338), .Z(O0[24]), .CO(n_340));
	notech_ha2 i_22(.A(\gdtr[23] ), .B(n_336), .Z(O0[23]), .CO(n_338));
	notech_ha2 i_21(.A(\gdtr[22] ), .B(n_334), .Z(O0[22]), .CO(n_336));
	notech_ha2 i_20(.A(\gdtr[21] ), .B(n_332), .Z(O0[21]), .CO(n_334));
	notech_ha2 i_19(.A(\gdtr[20] ), .B(n_330), .Z(O0[20]), .CO(n_332));
	notech_ha2 i_18(.A(\gdtr[19] ), .B(n_328), .Z(O0[19]), .CO(n_330));
	notech_ha2 i_17(.A(\gdtr[18] ), .B(n_326), .Z(O0[18]), .CO(n_328));
	notech_ha2 i_16(.A(\gdtr[17] ), .B(n_324), .Z(O0[17]), .CO(n_326));
	notech_ha2 i_15(.A(\gdtr[16] ), .B(n_285), .Z(O0[16]), .CO(n_324));
	notech_fa2 i_14(.A(I0[15]), .B(n_283), .CI(\gdtr[15] ), .Z(O0[15]), .CO(n_285
		));
	notech_fa2 i_13(.A(I0[14]), .B(n_281), .CI(\gdtr[14] ), .Z(O0[14]), .CO(n_283
		));
	notech_fa2 i_12(.A(I0[13]), .B(n_279), .CI(\gdtr[13] ), .Z(O0[13]), .CO(n_281
		));
	notech_fa2 i_11(.A(I0[12]), .B(n_277), .CI(\gdtr[12] ), .Z(O0[12]), .CO(n_279
		));
	notech_fa2 i_10(.A(I0[11]), .B(n_275), .CI(\gdtr[11] ), .Z(O0[11]), .CO(n_277
		));
	notech_fa2 i_9(.A(I0[10]), .B(n_273), .CI(\gdtr[10] ), .Z(O0[10]), .CO(n_275
		));
	notech_fa2 i_8(.A(I0[9]), .B(n_271), .CI(\gdtr[9] ), .Z(O0[9]), .CO(n_273
		));
	notech_fa2 i_7(.A(I0[8]), .B(n_269), .CI(\gdtr[8] ), .Z(O0[8]), .CO(n_271
		));
	notech_fa2 i_6(.A(I0[7]), .B(n_267), .CI(\gdtr[7] ), .Z(O0[7]), .CO(n_269
		));
	notech_fa2 i_5(.A(I0[6]), .B(n_265), .CI(\gdtr[6] ), .Z(O0[6]), .CO(n_267
		));
	notech_fa2 i_4(.A(I0[5]), .B(n_263), .CI(\gdtr[5] ), .Z(O0[5]), .CO(n_265
		));
	notech_fa2 i_3(.A(I0[4]), .B(n_261), .CI(\gdtr[4] ), .Z(O0[4]), .CO(n_263
		));
	notech_fa2 i_2(.A(I0[3]), .B(n_322), .CI(\gdtr[3] ), .Z(O0[3]), .CO(n_261
		));
	notech_ha2 i_1(.A(\gdtr[2] ), .B(\gdtr[1] ), .Z(O0[2]), .CO(n_322));
	notech_inv i_0(.A(\gdtr[1] ), .Z(O0[1]));
endmodule
module AWDP_ADD_239(O0, Daddrs);

	output [31:0] O0;
	input [31:0] Daddrs;

	wire \Daddrs[2] ;
	wire \Daddrs[3] ;
	wire \Daddrs[4] ;
	wire \Daddrs[5] ;
	wire \Daddrs[6] ;
	wire \Daddrs[7] ;
	wire \Daddrs[8] ;
	wire \Daddrs[9] ;
	wire \Daddrs[10] ;
	wire \Daddrs[11] ;
	wire \Daddrs[12] ;
	wire \Daddrs[13] ;
	wire \Daddrs[14] ;
	wire \Daddrs[15] ;
	wire \Daddrs[16] ;
	wire \Daddrs[17] ;
	wire \Daddrs[18] ;
	wire \Daddrs[19] ;
	wire \Daddrs[20] ;
	wire \Daddrs[21] ;
	wire \Daddrs[22] ;
	wire \Daddrs[23] ;
	wire \Daddrs[24] ;
	wire \Daddrs[25] ;
	wire \Daddrs[26] ;
	wire \Daddrs[27] ;
	wire \Daddrs[28] ;
	wire \Daddrs[29] ;
	wire \Daddrs[30] ;
	wire \Daddrs[31] ;


	assign O0[0] = Daddrs[0];
	assign O0[1] = Daddrs[1];
	assign \Daddrs[2]  = Daddrs[2];
	assign \Daddrs[3]  = Daddrs[3];
	assign \Daddrs[4]  = Daddrs[4];
	assign \Daddrs[5]  = Daddrs[5];
	assign \Daddrs[6]  = Daddrs[6];
	assign \Daddrs[7]  = Daddrs[7];
	assign \Daddrs[8]  = Daddrs[8];
	assign \Daddrs[9]  = Daddrs[9];
	assign \Daddrs[10]  = Daddrs[10];
	assign \Daddrs[11]  = Daddrs[11];
	assign \Daddrs[12]  = Daddrs[12];
	assign \Daddrs[13]  = Daddrs[13];
	assign \Daddrs[14]  = Daddrs[14];
	assign \Daddrs[15]  = Daddrs[15];
	assign \Daddrs[16]  = Daddrs[16];
	assign \Daddrs[17]  = Daddrs[17];
	assign \Daddrs[18]  = Daddrs[18];
	assign \Daddrs[19]  = Daddrs[19];
	assign \Daddrs[20]  = Daddrs[20];
	assign \Daddrs[21]  = Daddrs[21];
	assign \Daddrs[22]  = Daddrs[22];
	assign \Daddrs[23]  = Daddrs[23];
	assign \Daddrs[24]  = Daddrs[24];
	assign \Daddrs[25]  = Daddrs[25];
	assign \Daddrs[26]  = Daddrs[26];
	assign \Daddrs[27]  = Daddrs[27];
	assign \Daddrs[28]  = Daddrs[28];
	assign \Daddrs[29]  = Daddrs[29];
	assign \Daddrs[30]  = Daddrs[30];
	assign \Daddrs[31]  = Daddrs[31];

	notech_ha2 i_29(.A(\Daddrs[31] ), .B(n_308), .Z(O0[31]));
	notech_ha2 i_28(.A(\Daddrs[30] ), .B(n_306), .Z(O0[30]), .CO(n_308));
	notech_ha2 i_27(.A(\Daddrs[29] ), .B(n_304), .Z(O0[29]), .CO(n_306));
	notech_ha2 i_26(.A(\Daddrs[28] ), .B(n_302), .Z(O0[28]), .CO(n_304));
	notech_ha2 i_25(.A(\Daddrs[27] ), .B(n_300), .Z(O0[27]), .CO(n_302));
	notech_ha2 i_24(.A(\Daddrs[26] ), .B(n_298), .Z(O0[26]), .CO(n_300));
	notech_ha2 i_23(.A(\Daddrs[25] ), .B(n_296), .Z(O0[25]), .CO(n_298));
	notech_ha2 i_22(.A(\Daddrs[24] ), .B(n_294), .Z(O0[24]), .CO(n_296));
	notech_ha2 i_21(.A(\Daddrs[23] ), .B(n_292), .Z(O0[23]), .CO(n_294));
	notech_ha2 i_20(.A(\Daddrs[22] ), .B(n_290), .Z(O0[22]), .CO(n_292));
	notech_ha2 i_19(.A(\Daddrs[21] ), .B(n_288), .Z(O0[21]), .CO(n_290));
	notech_ha2 i_18(.A(\Daddrs[20] ), .B(n_286), .Z(O0[20]), .CO(n_288));
	notech_ha2 i_17(.A(\Daddrs[19] ), .B(n_284), .Z(O0[19]), .CO(n_286));
	notech_ha2 i_16(.A(\Daddrs[18] ), .B(n_282), .Z(O0[18]), .CO(n_284));
	notech_ha2 i_15(.A(\Daddrs[17] ), .B(n_280), .Z(O0[17]), .CO(n_282));
	notech_ha2 i_14(.A(\Daddrs[16] ), .B(n_278), .Z(O0[16]), .CO(n_280));
	notech_ha2 i_13(.A(\Daddrs[15] ), .B(n_276), .Z(O0[15]), .CO(n_278));
	notech_ha2 i_12(.A(\Daddrs[14] ), .B(n_274), .Z(O0[14]), .CO(n_276));
	notech_ha2 i_11(.A(\Daddrs[13] ), .B(n_272), .Z(O0[13]), .CO(n_274));
	notech_ha2 i_10(.A(\Daddrs[12] ), .B(n_270), .Z(O0[12]), .CO(n_272));
	notech_ha2 i_9(.A(\Daddrs[11] ), .B(n_268), .Z(O0[11]), .CO(n_270));
	notech_ha2 i_8(.A(\Daddrs[10] ), .B(n_266), .Z(O0[10]), .CO(n_268));
	notech_ha2 i_7(.A(\Daddrs[9] ), .B(n_264), .Z(O0[9]), .CO(n_266));
	notech_ha2 i_6(.A(\Daddrs[8] ), .B(n_262), .Z(O0[8]), .CO(n_264));
	notech_ha2 i_5(.A(\Daddrs[7] ), .B(n_260), .Z(O0[7]), .CO(n_262));
	notech_ha2 i_4(.A(\Daddrs[6] ), .B(n_258), .Z(O0[6]), .CO(n_260));
	notech_ha2 i_3(.A(\Daddrs[5] ), .B(n_256), .Z(O0[5]), .CO(n_258));
	notech_ha2 i_2(.A(\Daddrs[4] ), .B(n_254), .Z(O0[4]), .CO(n_256));
	notech_ha2 i_1(.A(\Daddrs[3] ), .B(\Daddrs[2] ), .Z(O0[3]), .CO(n_254)
		);
	notech_inv i_0(.A(\Daddrs[2] ), .Z(O0[2]));
endmodule
module AWDP_ADD_241(O0, opd, desc);
    output [31:0] O0;
    input [31:0] opd;
    input [31:0] desc;
    // Line 1144
    wire [31:0] O0;
    // Line 1146
    wire [31:0] N238;

    // Line 1144
    assign O0 = N238;
    // Line 1146
    assign N238 = desc + opd;
endmodule

module AWDP_ADD_25(add_len_pc16, regs_14, lenpc);
    output [15:0] add_len_pc16;
    input [15:0] regs_14;
    input [15:0] lenpc;
    // Line 156
    wire [15:0] add_len_pc16;
    // Line 154
    wire [15:0] N248;

    // Line 156
    assign add_len_pc16 = N248;
    // Line 154
    assign N248 = lenpc + regs_14;
endmodule

module AWDP_ADD_36(O0, opd);

	output [31:0] O0;
	input [31:0] opd;

	wire \opd[2] ;
	wire \opd[3] ;
	wire \opd[4] ;
	wire \opd[5] ;
	wire \opd[6] ;
	wire \opd[7] ;
	wire \opd[8] ;
	wire \opd[9] ;
	wire \opd[10] ;
	wire \opd[11] ;
	wire \opd[12] ;
	wire \opd[13] ;
	wire \opd[14] ;
	wire \opd[15] ;
	wire \opd[16] ;
	wire \opd[17] ;
	wire \opd[18] ;
	wire \opd[19] ;
	wire \opd[20] ;
	wire \opd[21] ;
	wire \opd[22] ;
	wire \opd[23] ;
	wire \opd[24] ;
	wire \opd[25] ;
	wire \opd[26] ;
	wire \opd[27] ;
	wire \opd[28] ;
	wire \opd[29] ;
	wire \opd[30] ;
	wire \opd[31] ;


	assign O0[0] = opd[0];
	assign O0[1] = opd[1];
	assign \opd[2]  = opd[2];
	assign \opd[3]  = opd[3];
	assign \opd[4]  = opd[4];
	assign \opd[5]  = opd[5];
	assign \opd[6]  = opd[6];
	assign \opd[7]  = opd[7];
	assign \opd[8]  = opd[8];
	assign \opd[9]  = opd[9];
	assign \opd[10]  = opd[10];
	assign \opd[11]  = opd[11];
	assign \opd[12]  = opd[12];
	assign \opd[13]  = opd[13];
	assign \opd[14]  = opd[14];
	assign \opd[15]  = opd[15];
	assign \opd[16]  = opd[16];
	assign \opd[17]  = opd[17];
	assign \opd[18]  = opd[18];
	assign \opd[19]  = opd[19];
	assign \opd[20]  = opd[20];
	assign \opd[21]  = opd[21];
	assign \opd[22]  = opd[22];
	assign \opd[23]  = opd[23];
	assign \opd[24]  = opd[24];
	assign \opd[25]  = opd[25];
	assign \opd[26]  = opd[26];
	assign \opd[27]  = opd[27];
	assign \opd[28]  = opd[28];
	assign \opd[29]  = opd[29];
	assign \opd[30]  = opd[30];
	assign \opd[31]  = opd[31];

	notech_ha2 i_29(.A(\opd[31] ), .B(n_308), .Z(O0[31]));
	notech_ha2 i_28(.A(\opd[30] ), .B(n_306), .Z(O0[30]), .CO(n_308));
	notech_ha2 i_27(.A(\opd[29] ), .B(n_304), .Z(O0[29]), .CO(n_306));
	notech_ha2 i_26(.A(\opd[28] ), .B(n_302), .Z(O0[28]), .CO(n_304));
	notech_ha2 i_25(.A(\opd[27] ), .B(n_300), .Z(O0[27]), .CO(n_302));
	notech_ha2 i_24(.A(\opd[26] ), .B(n_298), .Z(O0[26]), .CO(n_300));
	notech_ha2 i_23(.A(\opd[25] ), .B(n_296), .Z(O0[25]), .CO(n_298));
	notech_ha2 i_22(.A(\opd[24] ), .B(n_294), .Z(O0[24]), .CO(n_296));
	notech_ha2 i_21(.A(\opd[23] ), .B(n_292), .Z(O0[23]), .CO(n_294));
	notech_ha2 i_20(.A(\opd[22] ), .B(n_290), .Z(O0[22]), .CO(n_292));
	notech_ha2 i_19(.A(\opd[21] ), .B(n_288), .Z(O0[21]), .CO(n_290));
	notech_ha2 i_18(.A(\opd[20] ), .B(n_286), .Z(O0[20]), .CO(n_288));
	notech_ha2 i_17(.A(\opd[19] ), .B(n_284), .Z(O0[19]), .CO(n_286));
	notech_ha2 i_16(.A(\opd[18] ), .B(n_282), .Z(O0[18]), .CO(n_284));
	notech_ha2 i_15(.A(\opd[17] ), .B(n_280), .Z(O0[17]), .CO(n_282));
	notech_ha2 i_14(.A(\opd[16] ), .B(n_278), .Z(O0[16]), .CO(n_280));
	notech_ha2 i_13(.A(\opd[15] ), .B(n_276), .Z(O0[15]), .CO(n_278));
	notech_ha2 i_12(.A(\opd[14] ), .B(n_274), .Z(O0[14]), .CO(n_276));
	notech_ha2 i_11(.A(\opd[13] ), .B(n_272), .Z(O0[13]), .CO(n_274));
	notech_ha2 i_10(.A(\opd[12] ), .B(n_270), .Z(O0[12]), .CO(n_272));
	notech_ha2 i_9(.A(\opd[11] ), .B(n_268), .Z(O0[11]), .CO(n_270));
	notech_ha2 i_8(.A(\opd[10] ), .B(n_266), .Z(O0[10]), .CO(n_268));
	notech_ha2 i_7(.A(\opd[9] ), .B(n_264), .Z(O0[9]), .CO(n_266));
	notech_ha2 i_6(.A(\opd[8] ), .B(n_262), .Z(O0[8]), .CO(n_264));
	notech_ha2 i_5(.A(\opd[7] ), .B(n_260), .Z(O0[7]), .CO(n_262));
	notech_ha2 i_4(.A(\opd[6] ), .B(n_258), .Z(O0[6]), .CO(n_260));
	notech_ha2 i_3(.A(\opd[5] ), .B(n_256), .Z(O0[5]), .CO(n_258));
	notech_ha2 i_2(.A(\opd[4] ), .B(n_254), .Z(O0[4]), .CO(n_256));
	notech_ha2 i_1(.A(\opd[3] ), .B(\opd[2] ), .Z(O0[3]), .CO(n_254));
	notech_inv i_0(.A(\opd[2] ), .Z(O0[2]));
endmodule
module AWDP_ADD_40(O0, I0, I1);

	output [31:0] O0;
	input [31:0] I0;
	input [31:0] I1;

	wire \I0[4] ;
	wire \I0[5] ;
	wire \I0[6] ;
	wire \I0[7] ;
	wire \I0[8] ;
	wire \I0[9] ;
	wire \I0[10] ;
	wire \I0[11] ;
	wire \I0[12] ;
	wire \I0[13] ;
	wire \I0[14] ;
	wire \I0[15] ;


	assign O0[0] = I0[0];
	assign O0[1] = I0[1];
	assign O0[2] = I0[2];
	assign O0[3] = I0[3];
	assign \I0[4]  = I0[4];
	assign \I0[5]  = I0[5];
	assign \I0[6]  = I0[6];
	assign \I0[7]  = I0[7];
	assign \I0[8]  = I0[8];
	assign \I0[9]  = I0[9];
	assign \I0[10]  = I0[10];
	assign \I0[11]  = I0[11];
	assign \I0[12]  = I0[12];
	assign \I0[13]  = I0[13];
	assign \I0[14]  = I0[14];
	assign \I0[15]  = I0[15];

	notech_ha2 i_27(.A(I1[31]), .B(n_376), .Z(O0[31]));
	notech_ha2 i_26(.A(I1[30]), .B(n_374), .Z(O0[30]), .CO(n_376));
	notech_ha2 i_25(.A(I1[29]), .B(n_372), .Z(O0[29]), .CO(n_374));
	notech_ha2 i_24(.A(I1[28]), .B(n_370), .Z(O0[28]), .CO(n_372));
	notech_ha2 i_23(.A(I1[27]), .B(n_368), .Z(O0[27]), .CO(n_370));
	notech_ha2 i_22(.A(I1[26]), .B(n_366), .Z(O0[26]), .CO(n_368));
	notech_ha2 i_21(.A(I1[25]), .B(n_364), .Z(O0[25]), .CO(n_366));
	notech_ha2 i_20(.A(I1[24]), .B(n_362), .Z(O0[24]), .CO(n_364));
	notech_ha2 i_19(.A(I1[23]), .B(n_360), .Z(O0[23]), .CO(n_362));
	notech_ha2 i_18(.A(I1[22]), .B(n_358), .Z(O0[22]), .CO(n_360));
	notech_ha2 i_17(.A(I1[21]), .B(n_356), .Z(O0[21]), .CO(n_358));
	notech_ha2 i_16(.A(I1[20]), .B(n_354), .Z(O0[20]), .CO(n_356));
	notech_ha2 i_15(.A(I1[19]), .B(n_352), .Z(O0[19]), .CO(n_354));
	notech_ha2 i_14(.A(I1[18]), .B(n_350), .Z(O0[18]), .CO(n_352));
	notech_ha2 i_13(.A(I1[17]), .B(n_348), .Z(O0[17]), .CO(n_350));
	notech_ha2 i_12(.A(I1[16]), .B(n_311), .Z(O0[16]), .CO(n_348));
	notech_fa2 i_11(.A(\I0[15] ), .B(n_309), .CI(I1[15]), .Z(O0[15]), .CO(n_311
		));
	notech_fa2 i_10(.A(\I0[14] ), .B(n_307), .CI(I1[14]), .Z(O0[14]), .CO(n_309
		));
	notech_fa2 i_9(.A(\I0[13] ), .B(n_305), .CI(I1[13]), .Z(O0[13]), .CO(n_307
		));
	notech_fa2 i_8(.A(\I0[12] ), .B(n_303), .CI(I1[12]), .Z(O0[12]), .CO(n_305
		));
	notech_fa2 i_7(.A(\I0[11] ), .B(n_301), .CI(I1[11]), .Z(O0[11]), .CO(n_303
		));
	notech_fa2 i_6(.A(\I0[10] ), .B(n_299), .CI(I1[10]), .Z(O0[10]), .CO(n_301
		));
	notech_fa2 i_5(.A(\I0[9] ), .B(n_297), .CI(I1[9]), .Z(O0[9]), .CO(n_299)
		);
	notech_fa2 i_4(.A(\I0[8] ), .B(n_295), .CI(I1[8]), .Z(O0[8]), .CO(n_297)
		);
	notech_fa2 i_3(.A(\I0[7] ), .B(n_293), .CI(I1[7]), .Z(O0[7]), .CO(n_295)
		);
	notech_fa2 i_2(.A(\I0[6] ), .B(n_291), .CI(I1[6]), .Z(O0[6]), .CO(n_293)
		);
	notech_fa2 i_1(.A(\I0[5] ), .B(n_346), .CI(I1[5]), .Z(O0[5]), .CO(n_291)
		);
	notech_ha2 i_0(.A(\I0[4] ), .B(I1[4]), .Z(O0[4]), .CO(n_346));
endmodule
module AWDP_ADD_47(O0, opa, I0);

	output [32:0] O0;
	input [31:0] opa;
	input [31:0] I0;




	notech_inv i_10755(.A(n_57040), .Z(n_57045));
	notech_inv i_10751(.A(n_57040), .Z(n_57041));
	notech_inv i_10750(.A(I0[19]), .Z(n_57040));
	notech_fa2 i_31(.A(n_57045), .B(n_354), .CI(opa[31]), .Z(O0[31]), .CO(O0
		[32]));
	notech_fa2 i_30(.A(n_57045), .B(n_352), .CI(opa[30]), .Z(O0[30]), .CO(n_354
		));
	notech_fa2 i_29(.A(n_57045), .B(n_350), .CI(opa[29]), .Z(O0[29]), .CO(n_352
		));
	notech_fa2 i_28(.A(n_57045), .B(n_348), .CI(opa[28]), .Z(O0[28]), .CO(n_350
		));
	notech_fa2 i_27(.A(n_57045), .B(n_346), .CI(opa[27]), .Z(O0[27]), .CO(n_348
		));
	notech_fa2 i_26(.A(n_57045), .B(n_344), .CI(opa[26]), .Z(O0[26]), .CO(n_346
		));
	notech_fa2 i_25(.A(n_57045), .B(n_342), .CI(opa[25]), .Z(O0[25]), .CO(n_344
		));
	notech_fa2 i_24(.A(n_57045), .B(n_340), .CI(opa[24]), .Z(O0[24]), .CO(n_342
		));
	notech_fa2 i_23(.A(n_57045), .B(n_338), .CI(opa[23]), .Z(O0[23]), .CO(n_340
		));
	notech_fa2 i_22(.A(n_57045), .B(n_336), .CI(opa[22]), .Z(O0[22]), .CO(n_338
		));
	notech_fa2 i_21(.A(n_57045), .B(n_334), .CI(opa[21]), .Z(O0[21]), .CO(n_336
		));
	notech_fa2 i_20(.A(n_57045), .B(n_332), .CI(opa[20]), .Z(O0[20]), .CO(n_334
		));
	notech_fa2 i_19(.A(n_57045), .B(n_330), .CI(opa[19]), .Z(O0[19]), .CO(n_332
		));
	notech_fa2 i_18(.A(n_57045), .B(n_328), .CI(opa[18]), .Z(O0[18]), .CO(n_330
		));
	notech_fa2 i_17(.A(n_57045), .B(n_326), .CI(opa[17]), .Z(O0[17]), .CO(n_328
		));
	notech_fa2 i_16(.A(n_57041), .B(n_324), .CI(opa[16]), .Z(O0[16]), .CO(n_326
		));
	notech_fa2 i_15(.A(n_57041), .B(n_322), .CI(opa[15]), .Z(O0[15]), .CO(n_324
		));
	notech_fa2 i_14(.A(n_57041), .B(n_320), .CI(opa[14]), .Z(O0[14]), .CO(n_322
		));
	notech_fa2 i_13(.A(n_57041), .B(n_318), .CI(opa[13]), .Z(O0[13]), .CO(n_320
		));
	notech_fa2 i_12(.A(n_57041), .B(n_316), .CI(opa[12]), .Z(O0[12]), .CO(n_318
		));
	notech_fa2 i_11(.A(n_57041), .B(n_314), .CI(opa[11]), .Z(O0[11]), .CO(n_316
		));
	notech_fa2 i_10(.A(n_57041), .B(n_312), .CI(opa[10]), .Z(O0[10]), .CO(n_314
		));
	notech_fa2 i_9(.A(n_57041), .B(n_310), .CI(opa[9]), .Z(O0[9]), .CO(n_312
		));
	notech_fa2 i_8(.A(n_57045), .B(n_308), .CI(opa[8]), .Z(O0[8]), .CO(n_310
		));
	notech_fa2 i_7(.A(n_57045), .B(n_306), .CI(opa[7]), .Z(O0[7]), .CO(n_308
		));
	notech_fa2 i_6(.A(n_57045), .B(n_304), .CI(opa[6]), .Z(O0[6]), .CO(n_306
		));
	notech_fa2 i_5(.A(n_57045), .B(n_302), .CI(opa[5]), .Z(O0[5]), .CO(n_304
		));
	notech_fa2 i_4(.A(n_57041), .B(n_300), .CI(opa[4]), .Z(O0[4]), .CO(n_302
		));
	notech_fa2 i_3(.A(n_57041), .B(n_298), .CI(opa[3]), .Z(O0[3]), .CO(n_300
		));
	notech_fa2 i_2(.A(n_57045), .B(n_296), .CI(opa[2]), .Z(O0[2]), .CO(n_298
		));
	notech_fa2 i_1(.A(I0[1]), .B(n_361), .CI(opa[1]), .Z(O0[1]), .CO(n_296)
		);
	notech_ha2 i_0(.A(opa[0]), .B(I0[0]), .Z(O0[0]), .CO(n_361));
endmodule
module AWDP_ADD_6(O0, opd, I0);

	output [16:0] O0;
	input [15:0] opd;
	input [15:0] I0;




	notech_fa2 i_15(.A(I0[4]), .B(n_178), .CI(opd[15]), .Z(O0[15]), .CO(O0[
		16]));
	notech_fa2 i_14(.A(I0[4]), .B(n_176), .CI(opd[14]), .Z(O0[14]), .CO(n_178
		));
	notech_fa2 i_13(.A(I0[4]), .B(n_174), .CI(opd[13]), .Z(O0[13]), .CO(n_176
		));
	notech_fa2 i_12(.A(I0[4]), .B(n_172), .CI(opd[12]), .Z(O0[12]), .CO(n_174
		));
	notech_fa2 i_11(.A(I0[4]), .B(n_170), .CI(opd[11]), .Z(O0[11]), .CO(n_172
		));
	notech_fa2 i_10(.A(I0[4]), .B(n_168), .CI(opd[10]), .Z(O0[10]), .CO(n_170
		));
	notech_fa2 i_9(.A(I0[4]), .B(n_166), .CI(opd[9]), .Z(O0[9]), .CO(n_168)
		);
	notech_fa2 i_8(.A(I0[4]), .B(n_164), .CI(opd[8]), .Z(O0[8]), .CO(n_166)
		);
	notech_fa2 i_7(.A(I0[4]), .B(n_162), .CI(opd[7]), .Z(O0[7]), .CO(n_164)
		);
	notech_fa2 i_6(.A(I0[4]), .B(n_160), .CI(opd[6]), .Z(O0[6]), .CO(n_162)
		);
	notech_fa2 i_5(.A(I0[4]), .B(n_158), .CI(opd[5]), .Z(O0[5]), .CO(n_160)
		);
	notech_fa2 i_4(.A(I0[4]), .B(n_156), .CI(opd[4]), .Z(O0[4]), .CO(n_158)
		);
	notech_fa2 i_3(.A(I0[4]), .B(n_154), .CI(opd[3]), .Z(O0[3]), .CO(n_156)
		);
	notech_fa2 i_2(.A(I0[4]), .B(n_152), .CI(opd[2]), .Z(O0[2]), .CO(n_154)
		);
	notech_fa2 i_1(.A(I0[1]), .B(n_185), .CI(opd[1]), .Z(O0[1]), .CO(n_152)
		);
	notech_ha2 i_0(.A(opd[0]), .B(I0[0]), .Z(O0[0]), .CO(n_185));
endmodule
module AWDP_ADD_60(O0, opb, I0);

	output [16:0] O0;
	input [15:0] opb;
	input [15:0] I0;




	notech_fa2 i_15(.A(I0[15]), .B(n_178), .CI(opb[15]), .Z(O0[15]), .CO(O0[
		16]));
	notech_fa2 i_14(.A(I0[15]), .B(n_176), .CI(opb[14]), .Z(O0[14]), .CO(n_178
		));
	notech_fa2 i_13(.A(I0[15]), .B(n_174), .CI(opb[13]), .Z(O0[13]), .CO(n_176
		));
	notech_fa2 i_12(.A(I0[15]), .B(n_172), .CI(opb[12]), .Z(O0[12]), .CO(n_174
		));
	notech_fa2 i_11(.A(I0[15]), .B(n_170), .CI(opb[11]), .Z(O0[11]), .CO(n_172
		));
	notech_fa2 i_10(.A(I0[15]), .B(n_168), .CI(opb[10]), .Z(O0[10]), .CO(n_170
		));
	notech_fa2 i_9(.A(I0[15]), .B(n_166), .CI(opb[9]), .Z(O0[9]), .CO(n_168)
		);
	notech_fa2 i_8(.A(I0[15]), .B(n_164), .CI(opb[8]), .Z(O0[8]), .CO(n_166)
		);
	notech_fa2 i_7(.A(I0[15]), .B(n_162), .CI(opb[7]), .Z(O0[7]), .CO(n_164)
		);
	notech_fa2 i_6(.A(I0[15]), .B(n_160), .CI(opb[6]), .Z(O0[6]), .CO(n_162)
		);
	notech_fa2 i_5(.A(I0[15]), .B(n_158), .CI(opb[5]), .Z(O0[5]), .CO(n_160)
		);
	notech_fa2 i_4(.A(I0[15]), .B(n_156), .CI(opb[4]), .Z(O0[4]), .CO(n_158)
		);
	notech_fa2 i_3(.A(I0[15]), .B(n_154), .CI(opb[3]), .Z(O0[3]), .CO(n_156)
		);
	notech_fa2 i_2(.A(I0[15]), .B(n_152), .CI(opb[2]), .Z(O0[2]), .CO(n_154)
		);
	notech_fa2 i_1(.A(I0[1]), .B(n_185), .CI(opb[1]), .Z(O0[1]), .CO(n_152)
		);
	notech_ha2 i_0(.A(opb[0]), .B(I0[0]), .Z(O0[0]), .CO(n_185));
endmodule
module AWDP_ADD_69(O0, ldtr, I0);

	output [31:0] O0;
	input [31:0] ldtr;
	input [31:0] I0;

	wire \ldtr[1] ;
	wire \ldtr[2] ;
	wire \ldtr[3] ;
	wire \ldtr[4] ;
	wire \ldtr[5] ;
	wire \ldtr[6] ;
	wire \ldtr[7] ;
	wire \ldtr[8] ;
	wire \ldtr[9] ;
	wire \ldtr[10] ;
	wire \ldtr[11] ;
	wire \ldtr[12] ;
	wire \ldtr[13] ;
	wire \ldtr[14] ;
	wire \ldtr[15] ;
	wire \ldtr[16] ;
	wire \ldtr[17] ;
	wire \ldtr[18] ;
	wire \ldtr[19] ;
	wire \ldtr[20] ;
	wire \ldtr[21] ;
	wire \ldtr[22] ;
	wire \ldtr[23] ;
	wire \ldtr[24] ;
	wire \ldtr[25] ;
	wire \ldtr[26] ;
	wire \ldtr[27] ;
	wire \ldtr[28] ;
	wire \ldtr[29] ;
	wire \ldtr[30] ;
	wire \ldtr[31] ;


	assign O0[0] = ldtr[0];
	assign \ldtr[1]  = ldtr[1];
	assign \ldtr[2]  = ldtr[2];
	assign \ldtr[3]  = ldtr[3];
	assign \ldtr[4]  = ldtr[4];
	assign \ldtr[5]  = ldtr[5];
	assign \ldtr[6]  = ldtr[6];
	assign \ldtr[7]  = ldtr[7];
	assign \ldtr[8]  = ldtr[8];
	assign \ldtr[9]  = ldtr[9];
	assign \ldtr[10]  = ldtr[10];
	assign \ldtr[11]  = ldtr[11];
	assign \ldtr[12]  = ldtr[12];
	assign \ldtr[13]  = ldtr[13];
	assign \ldtr[14]  = ldtr[14];
	assign \ldtr[15]  = ldtr[15];
	assign \ldtr[16]  = ldtr[16];
	assign \ldtr[17]  = ldtr[17];
	assign \ldtr[18]  = ldtr[18];
	assign \ldtr[19]  = ldtr[19];
	assign \ldtr[20]  = ldtr[20];
	assign \ldtr[21]  = ldtr[21];
	assign \ldtr[22]  = ldtr[22];
	assign \ldtr[23]  = ldtr[23];
	assign \ldtr[24]  = ldtr[24];
	assign \ldtr[25]  = ldtr[25];
	assign \ldtr[26]  = ldtr[26];
	assign \ldtr[27]  = ldtr[27];
	assign \ldtr[28]  = ldtr[28];
	assign \ldtr[29]  = ldtr[29];
	assign \ldtr[30]  = ldtr[30];
	assign \ldtr[31]  = ldtr[31];

	notech_fa2 i_30(.A(I0[31]), .B(n_347), .CI(\ldtr[31] ), .Z(O0[31]));
	notech_fa2 i_29(.A(I0[30]), .B(n_345), .CI(\ldtr[30] ), .Z(O0[30]), .CO(n_347
		));
	notech_fa2 i_28(.A(I0[29]), .B(n_343), .CI(\ldtr[29] ), .Z(O0[29]), .CO(n_345
		));
	notech_fa2 i_27(.A(I0[28]), .B(n_341), .CI(\ldtr[28] ), .Z(O0[28]), .CO(n_343
		));
	notech_fa2 i_26(.A(I0[27]), .B(n_339), .CI(\ldtr[27] ), .Z(O0[27]), .CO(n_341
		));
	notech_fa2 i_25(.A(I0[26]), .B(n_337), .CI(\ldtr[26] ), .Z(O0[26]), .CO(n_339
		));
	notech_fa2 i_24(.A(I0[25]), .B(n_335), .CI(\ldtr[25] ), .Z(O0[25]), .CO(n_337
		));
	notech_fa2 i_23(.A(I0[24]), .B(n_333), .CI(\ldtr[24] ), .Z(O0[24]), .CO(n_335
		));
	notech_fa2 i_22(.A(I0[23]), .B(n_331), .CI(\ldtr[23] ), .Z(O0[23]), .CO(n_333
		));
	notech_fa2 i_21(.A(I0[22]), .B(n_329), .CI(\ldtr[22] ), .Z(O0[22]), .CO(n_331
		));
	notech_fa2 i_20(.A(I0[21]), .B(n_327), .CI(\ldtr[21] ), .Z(O0[21]), .CO(n_329
		));
	notech_fa2 i_19(.A(I0[20]), .B(n_325), .CI(\ldtr[20] ), .Z(O0[20]), .CO(n_327
		));
	notech_fa2 i_18(.A(I0[19]), .B(n_323), .CI(\ldtr[19] ), .Z(O0[19]), .CO(n_325
		));
	notech_fa2 i_17(.A(I0[18]), .B(n_321), .CI(\ldtr[18] ), .Z(O0[18]), .CO(n_323
		));
	notech_fa2 i_16(.A(I0[17]), .B(n_319), .CI(\ldtr[17] ), .Z(O0[17]), .CO(n_321
		));
	notech_fa2 i_15(.A(I0[16]), .B(n_317), .CI(\ldtr[16] ), .Z(O0[16]), .CO(n_319
		));
	notech_fa2 i_14(.A(I0[15]), .B(n_315), .CI(\ldtr[15] ), .Z(O0[15]), .CO(n_317
		));
	notech_fa2 i_13(.A(I0[14]), .B(n_313), .CI(\ldtr[14] ), .Z(O0[14]), .CO(n_315
		));
	notech_fa2 i_12(.A(I0[13]), .B(n_311), .CI(\ldtr[13] ), .Z(O0[13]), .CO(n_313
		));
	notech_fa2 i_11(.A(I0[12]), .B(n_309), .CI(\ldtr[12] ), .Z(O0[12]), .CO(n_311
		));
	notech_fa2 i_10(.A(I0[11]), .B(n_307), .CI(\ldtr[11] ), .Z(O0[11]), .CO(n_309
		));
	notech_fa2 i_9(.A(I0[10]), .B(n_305), .CI(\ldtr[10] ), .Z(O0[10]), .CO(n_307
		));
	notech_fa2 i_8(.A(I0[9]), .B(n_303), .CI(\ldtr[9] ), .Z(O0[9]), .CO(n_305
		));
	notech_fa2 i_7(.A(I0[8]), .B(n_301), .CI(\ldtr[8] ), .Z(O0[8]), .CO(n_303
		));
	notech_fa2 i_6(.A(I0[7]), .B(n_299), .CI(\ldtr[7] ), .Z(O0[7]), .CO(n_301
		));
	notech_fa2 i_5(.A(I0[6]), .B(n_297), .CI(\ldtr[6] ), .Z(O0[6]), .CO(n_299
		));
	notech_fa2 i_4(.A(I0[5]), .B(n_295), .CI(\ldtr[5] ), .Z(O0[5]), .CO(n_297
		));
	notech_fa2 i_3(.A(I0[4]), .B(n_293), .CI(\ldtr[4] ), .Z(O0[4]), .CO(n_295
		));
	notech_fa2 i_2(.A(I0[3]), .B(n_354), .CI(\ldtr[3] ), .Z(O0[3]), .CO(n_293
		));
	notech_ha2 i_1(.A(\ldtr[2] ), .B(\ldtr[1] ), .Z(O0[2]), .CO(n_354));
	notech_inv i_0(.A(\ldtr[1] ), .Z(O0[1]));
endmodule
module AWDP_ADD_8(O0, Daddrs);

	output [31:0] O0;
	input [31:0] Daddrs;

	wire \Daddrs[1] ;
	wire \Daddrs[2] ;
	wire \Daddrs[3] ;
	wire \Daddrs[4] ;
	wire \Daddrs[5] ;
	wire \Daddrs[6] ;
	wire \Daddrs[7] ;
	wire \Daddrs[8] ;
	wire \Daddrs[9] ;
	wire \Daddrs[10] ;
	wire \Daddrs[11] ;
	wire \Daddrs[12] ;
	wire \Daddrs[13] ;
	wire \Daddrs[14] ;
	wire \Daddrs[15] ;
	wire \Daddrs[16] ;
	wire \Daddrs[17] ;
	wire \Daddrs[18] ;
	wire \Daddrs[19] ;
	wire \Daddrs[20] ;
	wire \Daddrs[21] ;
	wire \Daddrs[22] ;
	wire \Daddrs[23] ;
	wire \Daddrs[24] ;
	wire \Daddrs[25] ;
	wire \Daddrs[26] ;
	wire \Daddrs[27] ;
	wire \Daddrs[28] ;
	wire \Daddrs[29] ;
	wire \Daddrs[30] ;
	wire \Daddrs[31] ;


	assign O0[0] = Daddrs[0];
	assign \Daddrs[1]  = Daddrs[1];
	assign \Daddrs[2]  = Daddrs[2];
	assign \Daddrs[3]  = Daddrs[3];
	assign \Daddrs[4]  = Daddrs[4];
	assign \Daddrs[5]  = Daddrs[5];
	assign \Daddrs[6]  = Daddrs[6];
	assign \Daddrs[7]  = Daddrs[7];
	assign \Daddrs[8]  = Daddrs[8];
	assign \Daddrs[9]  = Daddrs[9];
	assign \Daddrs[10]  = Daddrs[10];
	assign \Daddrs[11]  = Daddrs[11];
	assign \Daddrs[12]  = Daddrs[12];
	assign \Daddrs[13]  = Daddrs[13];
	assign \Daddrs[14]  = Daddrs[14];
	assign \Daddrs[15]  = Daddrs[15];
	assign \Daddrs[16]  = Daddrs[16];
	assign \Daddrs[17]  = Daddrs[17];
	assign \Daddrs[18]  = Daddrs[18];
	assign \Daddrs[19]  = Daddrs[19];
	assign \Daddrs[20]  = Daddrs[20];
	assign \Daddrs[21]  = Daddrs[21];
	assign \Daddrs[22]  = Daddrs[22];
	assign \Daddrs[23]  = Daddrs[23];
	assign \Daddrs[24]  = Daddrs[24];
	assign \Daddrs[25]  = Daddrs[25];
	assign \Daddrs[26]  = Daddrs[26];
	assign \Daddrs[27]  = Daddrs[27];
	assign \Daddrs[28]  = Daddrs[28];
	assign \Daddrs[29]  = Daddrs[29];
	assign \Daddrs[30]  = Daddrs[30];
	assign \Daddrs[31]  = Daddrs[31];

	notech_ha2 i_30(.A(\Daddrs[31] ), .B(n_312), .Z(O0[31]));
	notech_ha2 i_29(.A(\Daddrs[30] ), .B(n_310), .Z(O0[30]), .CO(n_312));
	notech_ha2 i_28(.A(\Daddrs[29] ), .B(n_308), .Z(O0[29]), .CO(n_310));
	notech_ha2 i_27(.A(\Daddrs[28] ), .B(n_306), .Z(O0[28]), .CO(n_308));
	notech_ha2 i_26(.A(\Daddrs[27] ), .B(n_304), .Z(O0[27]), .CO(n_306));
	notech_ha2 i_25(.A(\Daddrs[26] ), .B(n_302), .Z(O0[26]), .CO(n_304));
	notech_ha2 i_24(.A(\Daddrs[25] ), .B(n_300), .Z(O0[25]), .CO(n_302));
	notech_ha2 i_23(.A(\Daddrs[24] ), .B(n_298), .Z(O0[24]), .CO(n_300));
	notech_ha2 i_22(.A(\Daddrs[23] ), .B(n_296), .Z(O0[23]), .CO(n_298));
	notech_ha2 i_21(.A(\Daddrs[22] ), .B(n_294), .Z(O0[22]), .CO(n_296));
	notech_ha2 i_20(.A(\Daddrs[21] ), .B(n_292), .Z(O0[21]), .CO(n_294));
	notech_ha2 i_19(.A(\Daddrs[20] ), .B(n_290), .Z(O0[20]), .CO(n_292));
	notech_ha2 i_18(.A(\Daddrs[19] ), .B(n_288), .Z(O0[19]), .CO(n_290));
	notech_ha2 i_17(.A(\Daddrs[18] ), .B(n_286), .Z(O0[18]), .CO(n_288));
	notech_ha2 i_16(.A(\Daddrs[17] ), .B(n_284), .Z(O0[17]), .CO(n_286));
	notech_ha2 i_15(.A(\Daddrs[16] ), .B(n_282), .Z(O0[16]), .CO(n_284));
	notech_ha2 i_14(.A(\Daddrs[15] ), .B(n_280), .Z(O0[15]), .CO(n_282));
	notech_ha2 i_13(.A(\Daddrs[14] ), .B(n_278), .Z(O0[14]), .CO(n_280));
	notech_ha2 i_12(.A(\Daddrs[13] ), .B(n_276), .Z(O0[13]), .CO(n_278));
	notech_ha2 i_11(.A(\Daddrs[12] ), .B(n_274), .Z(O0[12]), .CO(n_276));
	notech_ha2 i_10(.A(\Daddrs[11] ), .B(n_272), .Z(O0[11]), .CO(n_274));
	notech_ha2 i_9(.A(\Daddrs[10] ), .B(n_270), .Z(O0[10]), .CO(n_272));
	notech_ha2 i_8(.A(\Daddrs[9] ), .B(n_268), .Z(O0[9]), .CO(n_270));
	notech_ha2 i_7(.A(\Daddrs[8] ), .B(n_266), .Z(O0[8]), .CO(n_268));
	notech_ha2 i_6(.A(\Daddrs[7] ), .B(n_264), .Z(O0[7]), .CO(n_266));
	notech_ha2 i_5(.A(\Daddrs[6] ), .B(n_262), .Z(O0[6]), .CO(n_264));
	notech_ha2 i_4(.A(\Daddrs[5] ), .B(n_260), .Z(O0[5]), .CO(n_262));
	notech_ha2 i_3(.A(\Daddrs[4] ), .B(n_258), .Z(O0[4]), .CO(n_260));
	notech_ha2 i_2(.A(\Daddrs[3] ), .B(n_256), .Z(O0[3]), .CO(n_258));
	notech_ha2 i_1(.A(\Daddrs[2] ), .B(\Daddrs[1] ), .Z(O0[2]), .CO(n_256)
		);
	notech_inv i_0(.A(\Daddrs[1] ), .Z(O0[1]));
endmodule
module AWDP_ADD_81(O0, opd, I0);

	output [32:0] O0;
	input [31:0] opd;
	input [31:0] I0;




	notech_inv i_10747(.A(n_57002), .Z(n_57007));
	notech_inv i_10743(.A(n_57002), .Z(n_57003));
	notech_inv i_10742(.A(I0[4]), .Z(n_57002));
	notech_fa2 i_31(.A(n_57007), .B(n_354), .CI(opd[31]), .Z(O0[31]), .CO(O0
		[32]));
	notech_fa2 i_30(.A(n_57007), .B(n_352), .CI(opd[30]), .Z(O0[30]), .CO(n_354
		));
	notech_fa2 i_29(.A(n_57007), .B(n_350), .CI(opd[29]), .Z(O0[29]), .CO(n_352
		));
	notech_fa2 i_28(.A(n_57007), .B(n_348), .CI(opd[28]), .Z(O0[28]), .CO(n_350
		));
	notech_fa2 i_27(.A(n_57007), .B(n_346), .CI(opd[27]), .Z(O0[27]), .CO(n_348
		));
	notech_fa2 i_26(.A(n_57007), .B(n_344), .CI(opd[26]), .Z(O0[26]), .CO(n_346
		));
	notech_fa2 i_25(.A(n_57007), .B(n_342), .CI(opd[25]), .Z(O0[25]), .CO(n_344
		));
	notech_fa2 i_24(.A(n_57007), .B(n_340), .CI(opd[24]), .Z(O0[24]), .CO(n_342
		));
	notech_fa2 i_23(.A(n_57007), .B(n_338), .CI(opd[23]), .Z(O0[23]), .CO(n_340
		));
	notech_fa2 i_22(.A(n_57007), .B(n_336), .CI(opd[22]), .Z(O0[22]), .CO(n_338
		));
	notech_fa2 i_21(.A(n_57007), .B(n_334), .CI(opd[21]), .Z(O0[21]), .CO(n_336
		));
	notech_fa2 i_20(.A(n_57007), .B(n_332), .CI(opd[20]), .Z(O0[20]), .CO(n_334
		));
	notech_fa2 i_19(.A(n_57007), .B(n_330), .CI(opd[19]), .Z(O0[19]), .CO(n_332
		));
	notech_fa2 i_18(.A(n_57007), .B(n_328), .CI(opd[18]), .Z(O0[18]), .CO(n_330
		));
	notech_fa2 i_17(.A(n_57007), .B(n_326), .CI(opd[17]), .Z(O0[17]), .CO(n_328
		));
	notech_fa2 i_16(.A(n_57003), .B(n_324), .CI(opd[16]), .Z(O0[16]), .CO(n_326
		));
	notech_fa2 i_15(.A(n_57003), .B(n_322), .CI(opd[15]), .Z(O0[15]), .CO(n_324
		));
	notech_fa2 i_14(.A(n_57003), .B(n_320), .CI(opd[14]), .Z(O0[14]), .CO(n_322
		));
	notech_fa2 i_13(.A(n_57003), .B(n_318), .CI(opd[13]), .Z(O0[13]), .CO(n_320
		));
	notech_fa2 i_12(.A(n_57003), .B(n_316), .CI(opd[12]), .Z(O0[12]), .CO(n_318
		));
	notech_fa2 i_11(.A(n_57003), .B(n_314), .CI(opd[11]), .Z(O0[11]), .CO(n_316
		));
	notech_fa2 i_10(.A(n_57003), .B(n_312), .CI(opd[10]), .Z(O0[10]), .CO(n_314
		));
	notech_fa2 i_9(.A(n_57003), .B(n_310), .CI(opd[9]), .Z(O0[9]), .CO(n_312
		));
	notech_fa2 i_8(.A(n_57007), .B(n_308), .CI(opd[8]), .Z(O0[8]), .CO(n_310
		));
	notech_fa2 i_7(.A(n_57007), .B(n_306), .CI(opd[7]), .Z(O0[7]), .CO(n_308
		));
	notech_fa2 i_6(.A(n_57007), .B(n_304), .CI(opd[6]), .Z(O0[6]), .CO(n_306
		));
	notech_fa2 i_5(.A(n_57007), .B(n_302), .CI(opd[5]), .Z(O0[5]), .CO(n_304
		));
	notech_fa2 i_4(.A(n_57003), .B(n_300), .CI(opd[4]), .Z(O0[4]), .CO(n_302
		));
	notech_fa2 i_3(.A(n_57003), .B(n_298), .CI(opd[3]), .Z(O0[3]), .CO(n_300
		));
	notech_fa2 i_2(.A(n_57007), .B(n_296), .CI(opd[2]), .Z(O0[2]), .CO(n_298
		));
	notech_fa2 i_1(.A(I0[1]), .B(n_361), .CI(opd[1]), .Z(O0[1]), .CO(n_296)
		);
	notech_ha2 i_0(.A(opd[0]), .B(I0[0]), .Z(O0[0]), .CO(n_361));
endmodule
module AWDP_ADD_97(add_len_pc32, regs_14, lenpc);
    output [31:0] add_len_pc32;
    input [31:0] regs_14;
    input [31:0] lenpc;
    // Line 155
    wire [31:0] N407;
    // Line 156
    wire [31:0] add_len_pc32;

    // Line 155
    assign N407 = lenpc + regs_14;
    // Line 156
    assign add_len_pc32 = N407;
endmodule

module AWDP_DEC_162(O0, cx);

	output [15:0] O0;
	input [15:0] cx;




	notech_ha2 i_16(.A(n_96), .B(n_126), .Z(O0[15]));
	notech_inv i_1(.A(cx[0]), .Z(O0[0]));
	notech_inv i_0(.A(cx[15]), .Z(n_96));
	notech_xor2 i_59682(.A(cx[14]), .B(n_124), .Z(n_42882));
	notech_inv i_59683(.A(n_42882), .Z(O0[14]));
	notech_or2 i_59681(.A(cx[14]), .B(n_124), .Z(n_126));
	notech_xor2 i_32(.A(cx[13]), .B(n_122), .Z(n_42909));
	notech_inv i_33(.A(n_42909), .Z(O0[13]));
	notech_or2 i_31(.A(cx[13]), .B(n_122), .Z(n_124));
	notech_xor2 i_30(.A(cx[12]), .B(n_120), .Z(n_42936));
	notech_inv i_3195048(.A(n_42936), .Z(O0[12]));
	notech_or2 i_29(.A(cx[12]), .B(n_120), .Z(n_122));
	notech_xor2 i_2995049(.A(cx[11]), .B(n_118), .Z(n_42963));
	notech_inv i_3095050(.A(n_42963), .Z(O0[11]));
	notech_or2 i_28(.A(cx[11]), .B(n_118), .Z(n_120));
	notech_xor2 i_2895051(.A(cx[10]), .B(n_116), .Z(n_42990));
	notech_inv i_2995052(.A(n_42990), .Z(O0[10]));
	notech_or2 i_27(.A(cx[10]), .B(n_116), .Z(n_118));
	notech_xor2 i_2795053(.A(cx[9]), .B(n_114), .Z(n_43017));
	notech_inv i_2895054(.A(n_43017), .Z(O0[9]));
	notech_or2 i_26(.A(cx[9]), .B(n_114), .Z(n_116));
	notech_xor2 i_2795055(.A(cx[8]), .B(n_112), .Z(n_43044));
	notech_inv i_2895056(.A(n_43044), .Z(O0[8]));
	notech_or2 i_2695057(.A(cx[8]), .B(n_112), .Z(n_114));
	notech_xor2 i_2795058(.A(cx[7]), .B(n_110), .Z(n_43071));
	notech_inv i_2895059(.A(n_43071), .Z(O0[7]));
	notech_or2 i_2695060(.A(cx[7]), .B(n_110), .Z(n_112));
	notech_xor2 i_2795061(.A(cx[6]), .B(n_108), .Z(n_43098));
	notech_inv i_2895062(.A(n_43098), .Z(O0[6]));
	notech_or2 i_2695063(.A(cx[6]), .B(n_108), .Z(n_110));
	notech_xor2 i_2795064(.A(cx[5]), .B(n_106), .Z(n_43125));
	notech_inv i_2895065(.A(n_43125), .Z(O0[5]));
	notech_or2 i_2695066(.A(cx[5]), .B(n_106), .Z(n_108));
	notech_xor2 i_2795067(.A(cx[4]), .B(n_104), .Z(n_43152));
	notech_inv i_2895068(.A(n_43152), .Z(O0[4]));
	notech_or2 i_2695069(.A(cx[4]), .B(n_104), .Z(n_106));
	notech_xor2 i_2795070(.A(cx[3]), .B(n_102), .Z(n_43179));
	notech_inv i_2895071(.A(n_43179), .Z(O0[3]));
	notech_or2 i_2695072(.A(cx[3]), .B(n_102), .Z(n_104));
	notech_xor2 i_2795073(.A(cx[2]), .B(n_100), .Z(n_43206));
	notech_inv i_2895074(.A(n_43206), .Z(O0[2]));
	notech_or2 i_2695075(.A(cx[2]), .B(n_100), .Z(n_102));
	notech_xor2 i_2795076(.A(cx[1]), .B(cx[0]), .Z(n_43234));
	notech_inv i_2895077(.A(n_43234), .Z(O0[1]));
	notech_or2 i_2695078(.A(cx[1]), .B(cx[0]), .Z(n_100));
endmodule
module AWDP_DEC_166(O0, ecx);

	output [31:0] O0;
	input [31:0] ecx;




	notech_ha2 i_32(.A(n_192), .B(n_254), .Z(O0[31]));
	notech_inv i_1(.A(ecx[0]), .Z(O0[0]));
	notech_inv i_0(.A(ecx[31]), .Z(n_192));
	notech_xor2 i_49(.A(ecx[30]), .B(n_252), .Z(n_43261));
	notech_inv i_50(.A(n_43261), .Z(O0[30]));
	notech_or2 i_48(.A(ecx[30]), .B(n_252), .Z(n_254));
	notech_xor2 i_4895079(.A(ecx[29]), .B(n_250), .Z(n_43288));
	notech_inv i_4995080(.A(n_43288), .Z(O0[29]));
	notech_or2 i_47(.A(ecx[29]), .B(n_250), .Z(n_252));
	notech_xor2 i_46(.A(ecx[28]), .B(n_248), .Z(n_43315));
	notech_inv i_4795081(.A(n_43315), .Z(O0[28]));
	notech_or2 i_45(.A(ecx[28]), .B(n_248), .Z(n_250));
	notech_xor2 i_4595082(.A(ecx[27]), .B(n_246), .Z(n_43342));
	notech_inv i_4695083(.A(n_43342), .Z(O0[27]));
	notech_or2 i_44(.A(ecx[27]), .B(n_246), .Z(n_248));
	notech_xor2 i_4495084(.A(ecx[26]), .B(n_244), .Z(n_43369));
	notech_inv i_4595085(.A(n_43369), .Z(O0[26]));
	notech_or2 i_43(.A(ecx[26]), .B(n_244), .Z(n_246));
	notech_xor2 i_4395086(.A(ecx[25]), .B(n_242), .Z(n_43396));
	notech_inv i_4495087(.A(n_43396), .Z(O0[25]));
	notech_or2 i_42(.A(ecx[25]), .B(n_242), .Z(n_244));
	notech_xor2 i_4295088(.A(ecx[24]), .B(n_240), .Z(n_43423));
	notech_inv i_4395089(.A(n_43423), .Z(O0[24]));
	notech_or2 i_41(.A(ecx[24]), .B(n_240), .Z(n_242));
	notech_xor2 i_4195090(.A(ecx[23]), .B(n_238), .Z(n_43450));
	notech_inv i_4295091(.A(n_43450), .Z(O0[23]));
	notech_or2 i_40(.A(ecx[23]), .B(n_238), .Z(n_240));
	notech_xor2 i_4095092(.A(ecx[22]), .B(n_236), .Z(n_43477));
	notech_inv i_4195093(.A(n_43477), .Z(O0[22]));
	notech_or2 i_39(.A(ecx[22]), .B(n_236), .Z(n_238));
	notech_xor2 i_3995094(.A(ecx[21]), .B(n_234), .Z(n_43504));
	notech_inv i_4095095(.A(n_43504), .Z(O0[21]));
	notech_or2 i_38(.A(ecx[21]), .B(n_234), .Z(n_236));
	notech_xor2 i_3895096(.A(ecx[20]), .B(n_232), .Z(n_43531));
	notech_inv i_3995097(.A(n_43531), .Z(O0[20]));
	notech_or2 i_37(.A(ecx[20]), .B(n_232), .Z(n_234));
	notech_xor2 i_3795098(.A(ecx[19]), .B(n_230), .Z(n_43558));
	notech_inv i_3895099(.A(n_43558), .Z(O0[19]));
	notech_or2 i_36(.A(ecx[19]), .B(n_230), .Z(n_232));
	notech_xor2 i_3695100(.A(ecx[18]), .B(n_228), .Z(n_43585));
	notech_inv i_3795101(.A(n_43585), .Z(O0[18]));
	notech_or2 i_35(.A(ecx[18]), .B(n_228), .Z(n_230));
	notech_xor2 i_3595102(.A(ecx[17]), .B(n_226), .Z(n_43612));
	notech_inv i_3695103(.A(n_43612), .Z(O0[17]));
	notech_or2 i_34(.A(ecx[17]), .B(n_226), .Z(n_228));
	notech_xor2 i_3495104(.A(ecx[16]), .B(n_224), .Z(n_43639));
	notech_inv i_3595105(.A(n_43639), .Z(O0[16]));
	notech_or2 i_33(.A(ecx[16]), .B(n_224), .Z(n_226));
	notech_xor2 i_3395106(.A(ecx[15]), .B(n_222), .Z(n_43666));
	notech_inv i_3495107(.A(n_43666), .Z(O0[15]));
	notech_or2 i_3295108(.A(ecx[15]), .B(n_222), .Z(n_224));
	notech_xor2 i_3295109(.A(ecx[14]), .B(n_220), .Z(n_43693));
	notech_inv i_3395110(.A(n_43693), .Z(O0[14]));
	notech_or2 i_31(.A(ecx[14]), .B(n_220), .Z(n_222));
	notech_xor2 i_3195111(.A(ecx[13]), .B(n_218), .Z(n_43720));
	notech_inv i_3295112(.A(n_43720), .Z(O0[13]));
	notech_or2 i_30(.A(ecx[13]), .B(n_218), .Z(n_220));
	notech_xor2 i_3095113(.A(ecx[12]), .B(n_216), .Z(n_43747));
	notech_inv i_3195114(.A(n_43747), .Z(O0[12]));
	notech_or2 i_29(.A(ecx[12]), .B(n_216), .Z(n_218));
	notech_xor2 i_2995115(.A(ecx[11]), .B(n_214), .Z(n_43774));
	notech_inv i_3095116(.A(n_43774), .Z(O0[11]));
	notech_or2 i_28(.A(ecx[11]), .B(n_214), .Z(n_216));
	notech_xor2 i_2895117(.A(ecx[10]), .B(n_212), .Z(n_43801));
	notech_inv i_2995118(.A(n_43801), .Z(O0[10]));
	notech_or2 i_27(.A(ecx[10]), .B(n_212), .Z(n_214));
	notech_xor2 i_2795119(.A(ecx[9]), .B(n_210), .Z(n_43828));
	notech_inv i_2895120(.A(n_43828), .Z(O0[9]));
	notech_or2 i_26(.A(ecx[9]), .B(n_210), .Z(n_212));
	notech_xor2 i_2795121(.A(ecx[8]), .B(n_208), .Z(n_43855));
	notech_inv i_2895122(.A(n_43855), .Z(O0[8]));
	notech_or2 i_2695123(.A(ecx[8]), .B(n_208), .Z(n_210));
	notech_xor2 i_2795124(.A(ecx[7]), .B(n_206), .Z(n_43882));
	notech_inv i_2895125(.A(n_43882), .Z(O0[7]));
	notech_or2 i_2695126(.A(ecx[7]), .B(n_206), .Z(n_208));
	notech_xor2 i_2795127(.A(ecx[6]), .B(n_204), .Z(n_43909));
	notech_inv i_2895128(.A(n_43909), .Z(O0[6]));
	notech_or2 i_2695129(.A(ecx[6]), .B(n_204), .Z(n_206));
	notech_xor2 i_2795130(.A(ecx[5]), .B(n_202), .Z(n_43936));
	notech_inv i_2895131(.A(n_43936), .Z(O0[5]));
	notech_or2 i_2695132(.A(ecx[5]), .B(n_202), .Z(n_204));
	notech_xor2 i_2795133(.A(ecx[4]), .B(n_200), .Z(n_43963));
	notech_inv i_2895134(.A(n_43963), .Z(O0[4]));
	notech_or2 i_2695135(.A(ecx[4]), .B(n_200), .Z(n_202));
	notech_xor2 i_2795136(.A(ecx[3]), .B(n_198), .Z(n_43990));
	notech_inv i_2895137(.A(n_43990), .Z(O0[3]));
	notech_or2 i_2695138(.A(ecx[3]), .B(n_198), .Z(n_200));
	notech_xor2 i_2795139(.A(ecx[2]), .B(n_196), .Z(n_44017));
	notech_inv i_2895140(.A(n_44017), .Z(O0[2]));
	notech_or2 i_2695141(.A(ecx[2]), .B(n_196), .Z(n_198));
	notech_xor2 i_2795142(.A(ecx[1]), .B(ecx[0]), .Z(n_44045));
	notech_inv i_2895143(.A(n_44045), .Z(O0[1]));
	notech_or2 i_2695144(.A(ecx[1]), .B(ecx[0]), .Z(n_196));
endmodule
module AWDP_DEC_2(O0, opc);

	output [31:0] O0;
	input [31:0] opc;




	notech_ha2 i_32(.A(n_192), .B(n_254), .Z(O0[31]));
	notech_inv i_1(.A(opc[0]), .Z(O0[0]));
	notech_inv i_0(.A(opc[31]), .Z(n_192));
	notech_xor2 i_49(.A(opc[30]), .B(n_252), .Z(n_44072));
	notech_inv i_50(.A(n_44072), .Z(O0[30]));
	notech_or2 i_48(.A(opc[30]), .B(n_252), .Z(n_254));
	notech_xor2 i_4895145(.A(opc[29]), .B(n_250), .Z(n_44099));
	notech_inv i_4995146(.A(n_44099), .Z(O0[29]));
	notech_or2 i_47(.A(opc[29]), .B(n_250), .Z(n_252));
	notech_xor2 i_46(.A(opc[28]), .B(n_248), .Z(n_44126));
	notech_inv i_4795147(.A(n_44126), .Z(O0[28]));
	notech_or2 i_45(.A(opc[28]), .B(n_248), .Z(n_250));
	notech_xor2 i_4595148(.A(opc[27]), .B(n_246), .Z(n_44153));
	notech_inv i_4695149(.A(n_44153), .Z(O0[27]));
	notech_or2 i_44(.A(opc[27]), .B(n_246), .Z(n_248));
	notech_xor2 i_4495150(.A(opc[26]), .B(n_244), .Z(n_44180));
	notech_inv i_4595151(.A(n_44180), .Z(O0[26]));
	notech_or2 i_43(.A(opc[26]), .B(n_244), .Z(n_246));
	notech_xor2 i_4395152(.A(opc[25]), .B(n_242), .Z(n_44207));
	notech_inv i_4495153(.A(n_44207), .Z(O0[25]));
	notech_or2 i_42(.A(opc[25]), .B(n_242), .Z(n_244));
	notech_xor2 i_4295154(.A(opc[24]), .B(n_240), .Z(n_44234));
	notech_inv i_4395155(.A(n_44234), .Z(O0[24]));
	notech_or2 i_41(.A(opc[24]), .B(n_240), .Z(n_242));
	notech_xor2 i_4195156(.A(opc[23]), .B(n_238), .Z(n_44261));
	notech_inv i_4295157(.A(n_44261), .Z(O0[23]));
	notech_or2 i_40(.A(opc[23]), .B(n_238), .Z(n_240));
	notech_xor2 i_4095158(.A(opc[22]), .B(n_236), .Z(n_44288));
	notech_inv i_4195159(.A(n_44288), .Z(O0[22]));
	notech_or2 i_39(.A(opc[22]), .B(n_236), .Z(n_238));
	notech_xor2 i_3995160(.A(opc[21]), .B(n_234), .Z(n_44315));
	notech_inv i_4095161(.A(n_44315), .Z(O0[21]));
	notech_or2 i_38(.A(opc[21]), .B(n_234), .Z(n_236));
	notech_xor2 i_3895162(.A(opc[20]), .B(n_232), .Z(n_44342));
	notech_inv i_3995163(.A(n_44342), .Z(O0[20]));
	notech_or2 i_37(.A(opc[20]), .B(n_232), .Z(n_234));
	notech_xor2 i_3795164(.A(opc[19]), .B(n_230), .Z(n_44369));
	notech_inv i_3895165(.A(n_44369), .Z(O0[19]));
	notech_or2 i_36(.A(opc[19]), .B(n_230), .Z(n_232));
	notech_xor2 i_3695166(.A(opc[18]), .B(n_228), .Z(n_44396));
	notech_inv i_3795167(.A(n_44396), .Z(O0[18]));
	notech_or2 i_35(.A(opc[18]), .B(n_228), .Z(n_230));
	notech_xor2 i_3595168(.A(opc[17]), .B(n_226), .Z(n_44423));
	notech_inv i_3695169(.A(n_44423), .Z(O0[17]));
	notech_or2 i_34(.A(opc[17]), .B(n_226), .Z(n_228));
	notech_xor2 i_3495170(.A(opc[16]), .B(n_224), .Z(n_44450));
	notech_inv i_3595171(.A(n_44450), .Z(O0[16]));
	notech_or2 i_33(.A(opc[16]), .B(n_224), .Z(n_226));
	notech_xor2 i_3395172(.A(opc[15]), .B(n_222), .Z(n_44477));
	notech_inv i_3495173(.A(n_44477), .Z(O0[15]));
	notech_or2 i_3295174(.A(opc[15]), .B(n_222), .Z(n_224));
	notech_xor2 i_3295175(.A(opc[14]), .B(n_220), .Z(n_44504));
	notech_inv i_3395176(.A(n_44504), .Z(O0[14]));
	notech_or2 i_31(.A(opc[14]), .B(n_220), .Z(n_222));
	notech_xor2 i_3195177(.A(opc[13]), .B(n_218), .Z(n_44531));
	notech_inv i_3295178(.A(n_44531), .Z(O0[13]));
	notech_or2 i_30(.A(opc[13]), .B(n_218), .Z(n_220));
	notech_xor2 i_3095179(.A(opc[12]), .B(n_216), .Z(n_44558));
	notech_inv i_3195180(.A(n_44558), .Z(O0[12]));
	notech_or2 i_29(.A(opc[12]), .B(n_216), .Z(n_218));
	notech_xor2 i_2995181(.A(opc[11]), .B(n_214), .Z(n_44585));
	notech_inv i_3095182(.A(n_44585), .Z(O0[11]));
	notech_or2 i_28(.A(opc[11]), .B(n_214), .Z(n_216));
	notech_xor2 i_2895183(.A(opc[10]), .B(n_212), .Z(n_44612));
	notech_inv i_2995184(.A(n_44612), .Z(O0[10]));
	notech_or2 i_27(.A(opc[10]), .B(n_212), .Z(n_214));
	notech_xor2 i_2795185(.A(opc[9]), .B(n_210), .Z(n_44639));
	notech_inv i_2895186(.A(n_44639), .Z(O0[9]));
	notech_or2 i_26(.A(opc[9]), .B(n_210), .Z(n_212));
	notech_xor2 i_2795187(.A(opc[8]), .B(n_208), .Z(n_44666));
	notech_inv i_2895188(.A(n_44666), .Z(O0[8]));
	notech_or2 i_2695189(.A(opc[8]), .B(n_208), .Z(n_210));
	notech_xor2 i_2795190(.A(opc[7]), .B(n_206), .Z(n_44693));
	notech_inv i_2895191(.A(n_44693), .Z(O0[7]));
	notech_or2 i_2695192(.A(opc[7]), .B(n_206), .Z(n_208));
	notech_xor2 i_2795193(.A(opc[6]), .B(n_204), .Z(n_44720));
	notech_inv i_2895194(.A(n_44720), .Z(O0[6]));
	notech_or2 i_2695195(.A(opc[6]), .B(n_204), .Z(n_206));
	notech_xor2 i_2795196(.A(opc[5]), .B(n_202), .Z(n_44747));
	notech_inv i_2895197(.A(n_44747), .Z(O0[5]));
	notech_or2 i_2695198(.A(opc[5]), .B(n_202), .Z(n_204));
	notech_xor2 i_2795199(.A(opc[4]), .B(n_200), .Z(n_44774));
	notech_inv i_2895200(.A(n_44774), .Z(O0[4]));
	notech_or2 i_2695201(.A(opc[4]), .B(n_200), .Z(n_202));
	notech_xor2 i_2795202(.A(opc[3]), .B(n_198), .Z(n_44801));
	notech_inv i_2895203(.A(n_44801), .Z(O0[3]));
	notech_or2 i_2695204(.A(opc[3]), .B(n_198), .Z(n_200));
	notech_xor2 i_2795205(.A(opc[2]), .B(n_196), .Z(n_44828));
	notech_inv i_2895206(.A(n_44828), .Z(O0[2]));
	notech_or2 i_2695207(.A(opc[2]), .B(n_196), .Z(n_198));
	notech_xor2 i_2795208(.A(opc[1]), .B(opc[0]), .Z(n_44856));
	notech_inv i_2895209(.A(n_44856), .Z(O0[1]));
	notech_or2 i_2695210(.A(opc[1]), .B(opc[0]), .Z(n_196));
endmodule
module AWDP_DEC_7(O0, opc);

	output [7:0] O0;
	input [7:0] opc;




	notech_ha2 i_8(.A(n_48), .B(n_62), .Z(O0[7]));
	notech_inv i_1(.A(opc[0]), .Z(O0[0]));
	notech_inv i_0(.A(opc[7]), .Z(n_48));
	notech_xor2 i_30(.A(opc[6]), .B(n_60), .Z(n_44883));
	notech_inv i_31(.A(n_44883), .Z(O0[6]));
	notech_or2 i_29(.A(opc[6]), .B(n_60), .Z(n_62));
	notech_xor2 i_27(.A(opc[5]), .B(n_58), .Z(n_44910));
	notech_inv i_28(.A(n_44910), .Z(O0[5]));
	notech_or2 i_26(.A(opc[5]), .B(n_58), .Z(n_60));
	notech_xor2 i_2795211(.A(opc[4]), .B(n_56), .Z(n_44937));
	notech_inv i_2895212(.A(n_44937), .Z(O0[4]));
	notech_or2 i_2695213(.A(opc[4]), .B(n_56), .Z(n_58));
	notech_xor2 i_2795214(.A(opc[3]), .B(n_54), .Z(n_44964));
	notech_inv i_2895215(.A(n_44964), .Z(O0[3]));
	notech_or2 i_2695216(.A(opc[3]), .B(n_54), .Z(n_56));
	notech_xor2 i_2795217(.A(opc[2]), .B(n_52), .Z(n_44991));
	notech_inv i_2895218(.A(n_44991), .Z(O0[2]));
	notech_or2 i_2695219(.A(opc[2]), .B(n_52), .Z(n_54));
	notech_xor2 i_2795220(.A(opc[1]), .B(opc[0]), .Z(n_45019));
	notech_inv i_2895221(.A(n_45019), .Z(O0[1]));
	notech_or2 i_2695222(.A(opc[1]), .B(opc[0]), .Z(n_52));
endmodule
module AWDP_EQ_125(O0, mul64);
    output [0:0] O0;
    input [63:32] mul64;
    // Line 131
    wire [0:0] O0;
    // Line 131
    wire [0:0] N551;

    // Line 131
    assign O0 = N551;
    // Line 131
    assign N551 = mul64 == 32'hffffffff;
endmodule

module AWDP_EQ_130(O0, mul64);
    output [0:0] O0;
    input [63:16] mul64;
    // Line 126
    wire [0:0] O0;
    // Line 126
    wire [0:0] N564;

    // Line 126
    assign O0 = N564;
    // Line 126
    assign N564 = mul64 == 48'h0;
endmodule

module AWDP_EQ_153(O0, mul64);
    output [0:0] O0;
    input [63:16] mul64;
    // Line 130
    wire [0:0] O0;
    // Line 130
    wire [0:0] N575;

    // Line 130
    assign O0 = N575;
    // Line 130
    assign N575 = mul64 == 48'hffffffff;
endmodule

module AWDP_EQ_218(O0, I0, I1);
    output [0:0] O0;
    input [63:0] I0;
    input [63:0] I1;
    // Line 790
    wire [0:0] N604;
    // Line 790
    wire [0:0] O0;

    // Line 790
    assign N604 = I0 == I1;
    // Line 790
    assign O0 = N604;
endmodule

module AWDP_EQ_58112339(O0, mul64);
    output [0:0] O0;
    input [63:8] mul64;
    // Line 129
    wire [0:0] N615;
    // Line 129
    wire [0:0] O0;

    // Line 129
    assign N615 = mul64 == 56'hffffffff;
    // Line 129
    assign O0 = N615;
endmodule

module AWDP_EQ_86(O0, mul64);
    output [0:0] O0;
    input [63:8] mul64;
    // Line 125
    wire [0:0] O0;
    // Line 125
    wire [0:0] N626;

    // Line 125
    assign O0 = N626;
    // Line 125
    assign N626 = mul64 == 56'h0;
endmodule

module AWDP_GE_12(O0, divr, divq);
    output [0:0] O0;
    input [63:0] divr;
    input [63:0] divq;
    // Line 1006
    wire [0:0] N639;
    // Line 1006
    wire [0:0] O0;

    // Line 1006
    assign N639 = divr >= divq;
    // Line 1006
    assign O0 = N639;
endmodule

module AWDP_INC_148(O0, I0);

	output [63:0] O0;
	input [63:0] I0;




	notech_ha2 i_63(.A(I0[63]), .B(n_636), .Z(O0[63]));
	notech_ha2 i_62(.A(I0[62]), .B(n_634), .Z(O0[62]), .CO(n_636));
	notech_ha2 i_61(.A(I0[61]), .B(n_632), .Z(O0[61]), .CO(n_634));
	notech_ha2 i_60(.A(I0[60]), .B(n_630), .Z(O0[60]), .CO(n_632));
	notech_ha2 i_59(.A(I0[59]), .B(n_628), .Z(O0[59]), .CO(n_630));
	notech_ha2 i_58(.A(I0[58]), .B(n_626), .Z(O0[58]), .CO(n_628));
	notech_ha2 i_57(.A(I0[57]), .B(n_624), .Z(O0[57]), .CO(n_626));
	notech_ha2 i_56(.A(I0[56]), .B(n_622), .Z(O0[56]), .CO(n_624));
	notech_ha2 i_55(.A(I0[55]), .B(n_620), .Z(O0[55]), .CO(n_622));
	notech_ha2 i_54(.A(I0[54]), .B(n_618), .Z(O0[54]), .CO(n_620));
	notech_ha2 i_53(.A(I0[53]), .B(n_616), .Z(O0[53]), .CO(n_618));
	notech_ha2 i_52(.A(I0[52]), .B(n_614), .Z(O0[52]), .CO(n_616));
	notech_ha2 i_51(.A(I0[51]), .B(n_612), .Z(O0[51]), .CO(n_614));
	notech_ha2 i_50(.A(I0[50]), .B(n_610), .Z(O0[50]), .CO(n_612));
	notech_ha2 i_49(.A(I0[49]), .B(n_608), .Z(O0[49]), .CO(n_610));
	notech_ha2 i_48(.A(I0[48]), .B(n_606), .Z(O0[48]), .CO(n_608));
	notech_ha2 i_47(.A(I0[47]), .B(n_604), .Z(O0[47]), .CO(n_606));
	notech_ha2 i_46(.A(I0[46]), .B(n_602), .Z(O0[46]), .CO(n_604));
	notech_ha2 i_45(.A(I0[45]), .B(n_600), .Z(O0[45]), .CO(n_602));
	notech_ha2 i_44(.A(I0[44]), .B(n_598), .Z(O0[44]), .CO(n_600));
	notech_ha2 i_43(.A(I0[43]), .B(n_596), .Z(O0[43]), .CO(n_598));
	notech_ha2 i_42(.A(I0[42]), .B(n_594), .Z(O0[42]), .CO(n_596));
	notech_ha2 i_41(.A(I0[41]), .B(n_592), .Z(O0[41]), .CO(n_594));
	notech_ha2 i_40(.A(I0[40]), .B(n_590), .Z(O0[40]), .CO(n_592));
	notech_ha2 i_39(.A(I0[39]), .B(n_588), .Z(O0[39]), .CO(n_590));
	notech_ha2 i_38(.A(I0[38]), .B(n_586), .Z(O0[38]), .CO(n_588));
	notech_ha2 i_37(.A(I0[37]), .B(n_584), .Z(O0[37]), .CO(n_586));
	notech_ha2 i_36(.A(I0[36]), .B(n_582), .Z(O0[36]), .CO(n_584));
	notech_ha2 i_35(.A(I0[35]), .B(n_580), .Z(O0[35]), .CO(n_582));
	notech_ha2 i_34(.A(I0[34]), .B(n_578), .Z(O0[34]), .CO(n_580));
	notech_ha2 i_33(.A(I0[33]), .B(n_576), .Z(O0[33]), .CO(n_578));
	notech_ha2 i_32(.A(I0[32]), .B(n_574), .Z(O0[32]), .CO(n_576));
	notech_ha2 i_31(.A(I0[31]), .B(n_572), .Z(O0[31]), .CO(n_574));
	notech_ha2 i_30(.A(I0[30]), .B(n_570), .Z(O0[30]), .CO(n_572));
	notech_ha2 i_29(.A(I0[29]), .B(n_568), .Z(O0[29]), .CO(n_570));
	notech_ha2 i_28(.A(I0[28]), .B(n_566), .Z(O0[28]), .CO(n_568));
	notech_ha2 i_27(.A(I0[27]), .B(n_564), .Z(O0[27]), .CO(n_566));
	notech_ha2 i_26(.A(I0[26]), .B(n_562), .Z(O0[26]), .CO(n_564));
	notech_ha2 i_25(.A(I0[25]), .B(n_560), .Z(O0[25]), .CO(n_562));
	notech_ha2 i_24(.A(I0[24]), .B(n_558), .Z(O0[24]), .CO(n_560));
	notech_ha2 i_23(.A(I0[23]), .B(n_556), .Z(O0[23]), .CO(n_558));
	notech_ha2 i_22(.A(I0[22]), .B(n_554), .Z(O0[22]), .CO(n_556));
	notech_ha2 i_21(.A(I0[21]), .B(n_552), .Z(O0[21]), .CO(n_554));
	notech_ha2 i_20(.A(I0[20]), .B(n_550), .Z(O0[20]), .CO(n_552));
	notech_ha2 i_19(.A(I0[19]), .B(n_548), .Z(O0[19]), .CO(n_550));
	notech_ha2 i_18(.A(I0[18]), .B(n_546), .Z(O0[18]), .CO(n_548));
	notech_ha2 i_17(.A(I0[17]), .B(n_544), .Z(O0[17]), .CO(n_546));
	notech_ha2 i_16(.A(I0[16]), .B(n_542), .Z(O0[16]), .CO(n_544));
	notech_ha2 i_15(.A(I0[15]), .B(n_540), .Z(O0[15]), .CO(n_542));
	notech_ha2 i_14(.A(I0[14]), .B(n_538), .Z(O0[14]), .CO(n_540));
	notech_ha2 i_13(.A(I0[13]), .B(n_536), .Z(O0[13]), .CO(n_538));
	notech_ha2 i_12(.A(I0[12]), .B(n_534), .Z(O0[12]), .CO(n_536));
	notech_ha2 i_11(.A(I0[11]), .B(n_532), .Z(O0[11]), .CO(n_534));
	notech_ha2 i_10(.A(I0[10]), .B(n_530), .Z(O0[10]), .CO(n_532));
	notech_ha2 i_9(.A(I0[9]), .B(n_528), .Z(O0[9]), .CO(n_530));
	notech_ha2 i_8(.A(I0[8]), .B(n_526), .Z(O0[8]), .CO(n_528));
	notech_ha2 i_7(.A(I0[7]), .B(n_524), .Z(O0[7]), .CO(n_526));
	notech_ha2 i_6(.A(I0[6]), .B(n_522), .Z(O0[6]), .CO(n_524));
	notech_ha2 i_5(.A(I0[5]), .B(n_520), .Z(O0[5]), .CO(n_522));
	notech_ha2 i_4(.A(I0[4]), .B(n_518), .Z(O0[4]), .CO(n_520));
	notech_ha2 i_3(.A(I0[3]), .B(n_516), .Z(O0[3]), .CO(n_518));
	notech_ha2 i_2(.A(I0[2]), .B(n_514), .Z(O0[2]), .CO(n_516));
	notech_ha2 i_1(.A(I0[1]), .B(I0[0]), .Z(O0[1]), .CO(n_514));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_INC_201(O0, tsc);

	output [63:0] O0;
	input [63:0] tsc;




	notech_ha2 i_63(.A(tsc[63]), .B(n_636), .Z(O0[63]));
	notech_ha2 i_62(.A(tsc[62]), .B(n_634), .Z(O0[62]), .CO(n_636));
	notech_ha2 i_61(.A(tsc[61]), .B(n_632), .Z(O0[61]), .CO(n_634));
	notech_ha2 i_60(.A(tsc[60]), .B(n_630), .Z(O0[60]), .CO(n_632));
	notech_ha2 i_59(.A(tsc[59]), .B(n_628), .Z(O0[59]), .CO(n_630));
	notech_ha2 i_58(.A(tsc[58]), .B(n_626), .Z(O0[58]), .CO(n_628));
	notech_ha2 i_57(.A(tsc[57]), .B(n_624), .Z(O0[57]), .CO(n_626));
	notech_ha2 i_56(.A(tsc[56]), .B(n_622), .Z(O0[56]), .CO(n_624));
	notech_ha2 i_55(.A(tsc[55]), .B(n_620), .Z(O0[55]), .CO(n_622));
	notech_ha2 i_54(.A(tsc[54]), .B(n_618), .Z(O0[54]), .CO(n_620));
	notech_ha2 i_53(.A(tsc[53]), .B(n_616), .Z(O0[53]), .CO(n_618));
	notech_ha2 i_52(.A(tsc[52]), .B(n_614), .Z(O0[52]), .CO(n_616));
	notech_ha2 i_51(.A(tsc[51]), .B(n_612), .Z(O0[51]), .CO(n_614));
	notech_ha2 i_50(.A(tsc[50]), .B(n_610), .Z(O0[50]), .CO(n_612));
	notech_ha2 i_49(.A(tsc[49]), .B(n_608), .Z(O0[49]), .CO(n_610));
	notech_ha2 i_48(.A(tsc[48]), .B(n_606), .Z(O0[48]), .CO(n_608));
	notech_ha2 i_47(.A(tsc[47]), .B(n_604), .Z(O0[47]), .CO(n_606));
	notech_ha2 i_46(.A(tsc[46]), .B(n_602), .Z(O0[46]), .CO(n_604));
	notech_ha2 i_45(.A(tsc[45]), .B(n_600), .Z(O0[45]), .CO(n_602));
	notech_ha2 i_44(.A(tsc[44]), .B(n_598), .Z(O0[44]), .CO(n_600));
	notech_ha2 i_43(.A(tsc[43]), .B(n_596), .Z(O0[43]), .CO(n_598));
	notech_ha2 i_42(.A(tsc[42]), .B(n_594), .Z(O0[42]), .CO(n_596));
	notech_ha2 i_41(.A(tsc[41]), .B(n_592), .Z(O0[41]), .CO(n_594));
	notech_ha2 i_40(.A(tsc[40]), .B(n_590), .Z(O0[40]), .CO(n_592));
	notech_ha2 i_39(.A(tsc[39]), .B(n_588), .Z(O0[39]), .CO(n_590));
	notech_ha2 i_38(.A(tsc[38]), .B(n_586), .Z(O0[38]), .CO(n_588));
	notech_ha2 i_37(.A(tsc[37]), .B(n_584), .Z(O0[37]), .CO(n_586));
	notech_ha2 i_36(.A(tsc[36]), .B(n_582), .Z(O0[36]), .CO(n_584));
	notech_ha2 i_35(.A(tsc[35]), .B(n_580), .Z(O0[35]), .CO(n_582));
	notech_ha2 i_34(.A(tsc[34]), .B(n_578), .Z(O0[34]), .CO(n_580));
	notech_ha2 i_33(.A(tsc[33]), .B(n_576), .Z(O0[33]), .CO(n_578));
	notech_ha2 i_32(.A(tsc[32]), .B(n_574), .Z(O0[32]), .CO(n_576));
	notech_ha2 i_31(.A(tsc[31]), .B(n_572), .Z(O0[31]), .CO(n_574));
	notech_ha2 i_30(.A(tsc[30]), .B(n_570), .Z(O0[30]), .CO(n_572));
	notech_ha2 i_29(.A(tsc[29]), .B(n_568), .Z(O0[29]), .CO(n_570));
	notech_ha2 i_28(.A(tsc[28]), .B(n_566), .Z(O0[28]), .CO(n_568));
	notech_ha2 i_27(.A(tsc[27]), .B(n_564), .Z(O0[27]), .CO(n_566));
	notech_ha2 i_26(.A(tsc[26]), .B(n_562), .Z(O0[26]), .CO(n_564));
	notech_ha2 i_25(.A(tsc[25]), .B(n_560), .Z(O0[25]), .CO(n_562));
	notech_ha2 i_24(.A(tsc[24]), .B(n_558), .Z(O0[24]), .CO(n_560));
	notech_ha2 i_23(.A(tsc[23]), .B(n_556), .Z(O0[23]), .CO(n_558));
	notech_ha2 i_22(.A(tsc[22]), .B(n_554), .Z(O0[22]), .CO(n_556));
	notech_ha2 i_21(.A(tsc[21]), .B(n_552), .Z(O0[21]), .CO(n_554));
	notech_ha2 i_20(.A(tsc[20]), .B(n_550), .Z(O0[20]), .CO(n_552));
	notech_ha2 i_19(.A(tsc[19]), .B(n_548), .Z(O0[19]), .CO(n_550));
	notech_ha2 i_18(.A(tsc[18]), .B(n_546), .Z(O0[18]), .CO(n_548));
	notech_ha2 i_17(.A(tsc[17]), .B(n_544), .Z(O0[17]), .CO(n_546));
	notech_ha2 i_16(.A(tsc[16]), .B(n_542), .Z(O0[16]), .CO(n_544));
	notech_ha2 i_15(.A(tsc[15]), .B(n_540), .Z(O0[15]), .CO(n_542));
	notech_ha2 i_14(.A(tsc[14]), .B(n_538), .Z(O0[14]), .CO(n_540));
	notech_ha2 i_13(.A(tsc[13]), .B(n_536), .Z(O0[13]), .CO(n_538));
	notech_ha2 i_12(.A(tsc[12]), .B(n_534), .Z(O0[12]), .CO(n_536));
	notech_ha2 i_11(.A(tsc[11]), .B(n_532), .Z(O0[11]), .CO(n_534));
	notech_ha2 i_10(.A(tsc[10]), .B(n_530), .Z(O0[10]), .CO(n_532));
	notech_ha2 i_9(.A(tsc[9]), .B(n_528), .Z(O0[9]), .CO(n_530));
	notech_ha2 i_8(.A(tsc[8]), .B(n_526), .Z(O0[8]), .CO(n_528));
	notech_ha2 i_7(.A(tsc[7]), .B(n_524), .Z(O0[7]), .CO(n_526));
	notech_ha2 i_6(.A(tsc[6]), .B(n_522), .Z(O0[6]), .CO(n_524));
	notech_ha2 i_5(.A(tsc[5]), .B(n_520), .Z(O0[5]), .CO(n_522));
	notech_ha2 i_4(.A(tsc[4]), .B(n_518), .Z(O0[4]), .CO(n_520));
	notech_ha2 i_3(.A(tsc[3]), .B(n_516), .Z(O0[3]), .CO(n_518));
	notech_ha2 i_2(.A(tsc[2]), .B(n_514), .Z(O0[2]), .CO(n_516));
	notech_ha2 i_1(.A(tsc[1]), .B(tsc[0]), .Z(O0[1]), .CO(n_514));
	notech_inv i_0(.A(tsc[0]), .Z(O0[0]));
endmodule
module AWDP_INC_235(O0, I0);

	output [31:0] O0;
	input [31:0] I0;




	notech_ha2 i_31(.A(I0[31]), .B(n_316), .Z(O0[31]));
	notech_ha2 i_30(.A(I0[30]), .B(n_314), .Z(O0[30]), .CO(n_316));
	notech_ha2 i_29(.A(I0[29]), .B(n_312), .Z(O0[29]), .CO(n_314));
	notech_ha2 i_28(.A(I0[28]), .B(n_310), .Z(O0[28]), .CO(n_312));
	notech_ha2 i_27(.A(I0[27]), .B(n_308), .Z(O0[27]), .CO(n_310));
	notech_ha2 i_26(.A(I0[26]), .B(n_306), .Z(O0[26]), .CO(n_308));
	notech_ha2 i_25(.A(I0[25]), .B(n_304), .Z(O0[25]), .CO(n_306));
	notech_ha2 i_24(.A(I0[24]), .B(n_302), .Z(O0[24]), .CO(n_304));
	notech_ha2 i_23(.A(I0[23]), .B(n_300), .Z(O0[23]), .CO(n_302));
	notech_ha2 i_22(.A(I0[22]), .B(n_298), .Z(O0[22]), .CO(n_300));
	notech_ha2 i_21(.A(I0[21]), .B(n_296), .Z(O0[21]), .CO(n_298));
	notech_ha2 i_20(.A(I0[20]), .B(n_294), .Z(O0[20]), .CO(n_296));
	notech_ha2 i_19(.A(I0[19]), .B(n_292), .Z(O0[19]), .CO(n_294));
	notech_ha2 i_18(.A(I0[18]), .B(n_290), .Z(O0[18]), .CO(n_292));
	notech_ha2 i_17(.A(I0[17]), .B(n_288), .Z(O0[17]), .CO(n_290));
	notech_ha2 i_16(.A(I0[16]), .B(n_286), .Z(O0[16]), .CO(n_288));
	notech_ha2 i_15(.A(I0[15]), .B(n_284), .Z(O0[15]), .CO(n_286));
	notech_ha2 i_14(.A(I0[14]), .B(n_282), .Z(O0[14]), .CO(n_284));
	notech_ha2 i_13(.A(I0[13]), .B(n_280), .Z(O0[13]), .CO(n_282));
	notech_ha2 i_12(.A(I0[12]), .B(n_278), .Z(O0[12]), .CO(n_280));
	notech_ha2 i_11(.A(I0[11]), .B(n_276), .Z(O0[11]), .CO(n_278));
	notech_ha2 i_10(.A(I0[10]), .B(n_274), .Z(O0[10]), .CO(n_276));
	notech_ha2 i_9(.A(I0[9]), .B(n_272), .Z(O0[9]), .CO(n_274));
	notech_ha2 i_8(.A(I0[8]), .B(n_270), .Z(O0[8]), .CO(n_272));
	notech_ha2 i_7(.A(I0[7]), .B(n_268), .Z(O0[7]), .CO(n_270));
	notech_ha2 i_6(.A(I0[6]), .B(n_266), .Z(O0[6]), .CO(n_268));
	notech_ha2 i_5(.A(I0[5]), .B(n_264), .Z(O0[5]), .CO(n_266));
	notech_ha2 i_4(.A(I0[4]), .B(n_262), .Z(O0[4]), .CO(n_264));
	notech_ha2 i_3(.A(I0[3]), .B(n_260), .Z(O0[3]), .CO(n_262));
	notech_ha2 i_2(.A(I0[2]), .B(n_258), .Z(O0[2]), .CO(n_260));
	notech_ha2 i_1(.A(I0[1]), .B(I0[0]), .Z(O0[1]), .CO(n_258));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_INC_26(O0, I0);

	output [31:0] O0;
	input [31:0] I0;




	notech_ha2 i_31(.A(I0[31]), .B(n_316), .Z(O0[31]));
	notech_ha2 i_30(.A(I0[30]), .B(n_314), .Z(O0[30]), .CO(n_316));
	notech_ha2 i_29(.A(I0[29]), .B(n_312), .Z(O0[29]), .CO(n_314));
	notech_ha2 i_28(.A(I0[28]), .B(n_310), .Z(O0[28]), .CO(n_312));
	notech_ha2 i_27(.A(I0[27]), .B(n_308), .Z(O0[27]), .CO(n_310));
	notech_ha2 i_26(.A(I0[26]), .B(n_306), .Z(O0[26]), .CO(n_308));
	notech_ha2 i_25(.A(I0[25]), .B(n_304), .Z(O0[25]), .CO(n_306));
	notech_ha2 i_24(.A(I0[24]), .B(n_302), .Z(O0[24]), .CO(n_304));
	notech_ha2 i_23(.A(I0[23]), .B(n_300), .Z(O0[23]), .CO(n_302));
	notech_ha2 i_22(.A(I0[22]), .B(n_298), .Z(O0[22]), .CO(n_300));
	notech_ha2 i_21(.A(I0[21]), .B(n_296), .Z(O0[21]), .CO(n_298));
	notech_ha2 i_20(.A(I0[20]), .B(n_294), .Z(O0[20]), .CO(n_296));
	notech_ha2 i_19(.A(I0[19]), .B(n_292), .Z(O0[19]), .CO(n_294));
	notech_ha2 i_18(.A(I0[18]), .B(n_290), .Z(O0[18]), .CO(n_292));
	notech_ha2 i_17(.A(I0[17]), .B(n_288), .Z(O0[17]), .CO(n_290));
	notech_ha2 i_16(.A(I0[16]), .B(n_286), .Z(O0[16]), .CO(n_288));
	notech_ha2 i_15(.A(I0[15]), .B(n_284), .Z(O0[15]), .CO(n_286));
	notech_ha2 i_14(.A(I0[14]), .B(n_282), .Z(O0[14]), .CO(n_284));
	notech_ha2 i_13(.A(I0[13]), .B(n_280), .Z(O0[13]), .CO(n_282));
	notech_ha2 i_12(.A(I0[12]), .B(n_278), .Z(O0[12]), .CO(n_280));
	notech_ha2 i_11(.A(I0[11]), .B(n_276), .Z(O0[11]), .CO(n_278));
	notech_ha2 i_10(.A(I0[10]), .B(n_274), .Z(O0[10]), .CO(n_276));
	notech_ha2 i_9(.A(I0[9]), .B(n_272), .Z(O0[9]), .CO(n_274));
	notech_ha2 i_8(.A(I0[8]), .B(n_270), .Z(O0[8]), .CO(n_272));
	notech_ha2 i_7(.A(I0[7]), .B(n_268), .Z(O0[7]), .CO(n_270));
	notech_ha2 i_6(.A(I0[6]), .B(n_266), .Z(O0[6]), .CO(n_268));
	notech_ha2 i_5(.A(I0[5]), .B(n_264), .Z(O0[5]), .CO(n_266));
	notech_ha2 i_4(.A(I0[4]), .B(n_262), .Z(O0[4]), .CO(n_264));
	notech_ha2 i_3(.A(I0[3]), .B(n_260), .Z(O0[3]), .CO(n_262));
	notech_ha2 i_2(.A(I0[2]), .B(n_258), .Z(O0[2]), .CO(n_260));
	notech_ha2 i_1(.A(I0[1]), .B(I0[0]), .Z(O0[1]), .CO(n_258));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_INC_77(O0, I0);

	output [15:0] O0;
	input [15:0] I0;




	notech_ha2 i_15(.A(I0[15]), .B(n_156), .Z(O0[15]));
	notech_ha2 i_14(.A(I0[14]), .B(n_154), .Z(O0[14]), .CO(n_156));
	notech_ha2 i_13(.A(I0[13]), .B(n_152), .Z(O0[13]), .CO(n_154));
	notech_ha2 i_12(.A(I0[12]), .B(n_150), .Z(O0[12]), .CO(n_152));
	notech_ha2 i_11(.A(I0[11]), .B(n_148), .Z(O0[11]), .CO(n_150));
	notech_ha2 i_10(.A(I0[10]), .B(n_146), .Z(O0[10]), .CO(n_148));
	notech_ha2 i_9(.A(I0[9]), .B(n_144), .Z(O0[9]), .CO(n_146));
	notech_ha2 i_8(.A(I0[8]), .B(n_142), .Z(O0[8]), .CO(n_144));
	notech_ha2 i_7(.A(I0[7]), .B(n_140), .Z(O0[7]), .CO(n_142));
	notech_ha2 i_6(.A(I0[6]), .B(n_138), .Z(O0[6]), .CO(n_140));
	notech_ha2 i_5(.A(I0[5]), .B(n_136), .Z(O0[5]), .CO(n_138));
	notech_ha2 i_4(.A(I0[4]), .B(n_134), .Z(O0[4]), .CO(n_136));
	notech_ha2 i_3(.A(I0[3]), .B(n_132), .Z(O0[3]), .CO(n_134));
	notech_ha2 i_2(.A(I0[2]), .B(n_130), .Z(O0[2]), .CO(n_132));
	notech_ha2 i_1(.A(I0[1]), .B(I0[0]), .Z(O0[1]), .CO(n_130));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_INC_78(O0, I0);

	output [31:0] O0;
	input [31:0] I0;




	notech_ha2 i_31(.A(I0[31]), .B(n_316), .Z(O0[31]));
	notech_ha2 i_30(.A(I0[30]), .B(n_314), .Z(O0[30]), .CO(n_316));
	notech_ha2 i_29(.A(I0[29]), .B(n_312), .Z(O0[29]), .CO(n_314));
	notech_ha2 i_28(.A(I0[28]), .B(n_310), .Z(O0[28]), .CO(n_312));
	notech_ha2 i_27(.A(I0[27]), .B(n_308), .Z(O0[27]), .CO(n_310));
	notech_ha2 i_26(.A(I0[26]), .B(n_306), .Z(O0[26]), .CO(n_308));
	notech_ha2 i_25(.A(I0[25]), .B(n_304), .Z(O0[25]), .CO(n_306));
	notech_ha2 i_24(.A(I0[24]), .B(n_302), .Z(O0[24]), .CO(n_304));
	notech_ha2 i_23(.A(I0[23]), .B(n_300), .Z(O0[23]), .CO(n_302));
	notech_ha2 i_22(.A(I0[22]), .B(n_298), .Z(O0[22]), .CO(n_300));
	notech_ha2 i_21(.A(I0[21]), .B(n_296), .Z(O0[21]), .CO(n_298));
	notech_ha2 i_20(.A(I0[20]), .B(n_294), .Z(O0[20]), .CO(n_296));
	notech_ha2 i_19(.A(I0[19]), .B(n_292), .Z(O0[19]), .CO(n_294));
	notech_ha2 i_18(.A(I0[18]), .B(n_290), .Z(O0[18]), .CO(n_292));
	notech_ha2 i_17(.A(I0[17]), .B(n_288), .Z(O0[17]), .CO(n_290));
	notech_ha2 i_16(.A(I0[16]), .B(n_286), .Z(O0[16]), .CO(n_288));
	notech_ha2 i_15(.A(I0[15]), .B(n_284), .Z(O0[15]), .CO(n_286));
	notech_ha2 i_14(.A(I0[14]), .B(n_282), .Z(O0[14]), .CO(n_284));
	notech_ha2 i_13(.A(I0[13]), .B(n_280), .Z(O0[13]), .CO(n_282));
	notech_ha2 i_12(.A(I0[12]), .B(n_278), .Z(O0[12]), .CO(n_280));
	notech_ha2 i_11(.A(I0[11]), .B(n_276), .Z(O0[11]), .CO(n_278));
	notech_ha2 i_10(.A(I0[10]), .B(n_274), .Z(O0[10]), .CO(n_276));
	notech_ha2 i_9(.A(I0[9]), .B(n_272), .Z(O0[9]), .CO(n_274));
	notech_ha2 i_8(.A(I0[8]), .B(n_270), .Z(O0[8]), .CO(n_272));
	notech_ha2 i_7(.A(I0[7]), .B(n_268), .Z(O0[7]), .CO(n_270));
	notech_ha2 i_6(.A(I0[6]), .B(n_266), .Z(O0[6]), .CO(n_268));
	notech_ha2 i_5(.A(I0[5]), .B(n_264), .Z(O0[5]), .CO(n_266));
	notech_ha2 i_4(.A(I0[4]), .B(n_262), .Z(O0[4]), .CO(n_264));
	notech_ha2 i_3(.A(I0[3]), .B(n_260), .Z(O0[3]), .CO(n_262));
	notech_ha2 i_2(.A(I0[2]), .B(n_258), .Z(O0[2]), .CO(n_260));
	notech_ha2 i_1(.A(I0[1]), .B(I0[0]), .Z(O0[1]), .CO(n_258));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_INC_99(O0, I0);

	output [63:0] O0;
	input [63:0] I0;




	notech_ha2 i_31(.A(I0[31]), .B(n_573), .Z(O0[31]), .CO(O0[32]));
	notech_ha2 i_30(.A(I0[30]), .B(n_571), .Z(O0[30]), .CO(n_573));
	notech_ha2 i_29(.A(I0[29]), .B(n_569), .Z(O0[29]), .CO(n_571));
	notech_ha2 i_28(.A(I0[28]), .B(n_567), .Z(O0[28]), .CO(n_569));
	notech_ha2 i_27(.A(I0[27]), .B(n_565), .Z(O0[27]), .CO(n_567));
	notech_ha2 i_26(.A(I0[26]), .B(n_563), .Z(O0[26]), .CO(n_565));
	notech_ha2 i_25(.A(I0[25]), .B(n_561), .Z(O0[25]), .CO(n_563));
	notech_ha2 i_24(.A(I0[24]), .B(n_559), .Z(O0[24]), .CO(n_561));
	notech_ha2 i_23(.A(I0[23]), .B(n_557), .Z(O0[23]), .CO(n_559));
	notech_ha2 i_22(.A(I0[22]), .B(n_555), .Z(O0[22]), .CO(n_557));
	notech_ha2 i_21(.A(I0[21]), .B(n_553), .Z(O0[21]), .CO(n_555));
	notech_ha2 i_20(.A(I0[20]), .B(n_551), .Z(O0[20]), .CO(n_553));
	notech_ha2 i_19(.A(I0[19]), .B(n_549), .Z(O0[19]), .CO(n_551));
	notech_ha2 i_18(.A(I0[18]), .B(n_547), .Z(O0[18]), .CO(n_549));
	notech_ha2 i_17(.A(I0[17]), .B(n_545), .Z(O0[17]), .CO(n_547));
	notech_ha2 i_16(.A(I0[16]), .B(n_543), .Z(O0[16]), .CO(n_545));
	notech_ha2 i_15(.A(I0[15]), .B(n_541), .Z(O0[15]), .CO(n_543));
	notech_ha2 i_14(.A(I0[14]), .B(n_539), .Z(O0[14]), .CO(n_541));
	notech_ha2 i_13(.A(I0[13]), .B(n_537), .Z(O0[13]), .CO(n_539));
	notech_ha2 i_12(.A(I0[12]), .B(n_535), .Z(O0[12]), .CO(n_537));
	notech_ha2 i_11(.A(I0[11]), .B(n_533), .Z(O0[11]), .CO(n_535));
	notech_ha2 i_10(.A(I0[10]), .B(n_531), .Z(O0[10]), .CO(n_533));
	notech_ha2 i_9(.A(I0[9]), .B(n_529), .Z(O0[9]), .CO(n_531));
	notech_ha2 i_8(.A(I0[8]), .B(n_527), .Z(O0[8]), .CO(n_529));
	notech_ha2 i_7(.A(I0[7]), .B(n_525), .Z(O0[7]), .CO(n_527));
	notech_ha2 i_6(.A(I0[6]), .B(n_523), .Z(O0[6]), .CO(n_525));
	notech_ha2 i_5(.A(I0[5]), .B(n_521), .Z(O0[5]), .CO(n_523));
	notech_ha2 i_4(.A(I0[4]), .B(n_519), .Z(O0[4]), .CO(n_521));
	notech_ha2 i_3(.A(I0[3]), .B(n_517), .Z(O0[3]), .CO(n_519));
	notech_ha2 i_2(.A(I0[2]), .B(n_515), .Z(O0[2]), .CO(n_517));
	notech_ha2 i_1(.A(I0[1]), .B(I0[0]), .Z(O0[1]), .CO(n_515));
	notech_inv i_0(.A(I0[0]), .Z(O0[0]));
endmodule
module AWDP_LE_209(O0, divq, I0);

	output [0:0] O0;
	input [63:0] divq;
	input [63:0] I0;




	notech_inv i_320(.A(n_710), .Z(O0[0]));
	notech_nand2 i_317(.A(n_703), .B(n_709), .Z(n_710));
	notech_inv i_506(.A(n_835), .Z(n_703));
	notech_or2 i_505(.A(n_834), .B(n_701), .Z(n_835));
	notech_and2 i_504(.A(n_702), .B(n_700), .Z(n_834));
	notech_inv i_315(.A(n_512), .Z(n_702));
	notech_inv i_314(.A(n_577), .Z(n_701));
	notech_inv i_503(.A(n_928), .Z(n_700));
	notech_nor2 i_502(.A(n_927), .B(n_866), .Z(n_928));
	notech_nor2 i_501(.A(n_699), .B(n_511), .Z(n_927));
	notech_inv i_500(.A(n_831), .Z(n_699));
	notech_or2 i_499(.A(n_830), .B(n_697), .Z(n_831));
	notech_and2 i_498(.A(n_698), .B(n_696), .Z(n_830));
	notech_inv i_311(.A(n_510), .Z(n_698));
	notech_inv i_310(.A(n_575), .Z(n_697));
	notech_inv i_497(.A(n_926), .Z(n_696));
	notech_nor2 i_496(.A(n_925), .B(n_865), .Z(n_926));
	notech_nor2 i_495(.A(n_695), .B(n_509), .Z(n_925));
	notech_inv i_494(.A(n_827), .Z(n_695));
	notech_or2 i_493(.A(n_826), .B(n_693), .Z(n_827));
	notech_and2 i_492(.A(n_694), .B(n_692), .Z(n_826));
	notech_inv i_307(.A(n_508), .Z(n_694));
	notech_inv i_306(.A(n_573), .Z(n_693));
	notech_inv i_491(.A(n_924), .Z(n_692));
	notech_nor2 i_490(.A(n_923), .B(n_864), .Z(n_924));
	notech_nor2 i_489(.A(n_691), .B(n_507), .Z(n_923));
	notech_inv i_488(.A(n_823), .Z(n_691));
	notech_or2 i_487(.A(n_822), .B(n_689), .Z(n_823));
	notech_and2 i_486(.A(n_690), .B(n_688), .Z(n_822));
	notech_inv i_303(.A(n_506), .Z(n_690));
	notech_inv i_302(.A(n_571), .Z(n_689));
	notech_inv i_485(.A(n_922), .Z(n_688));
	notech_nor2 i_484(.A(n_921), .B(n_863), .Z(n_922));
	notech_nor2 i_483(.A(n_687), .B(n_505), .Z(n_921));
	notech_inv i_482(.A(n_819), .Z(n_687));
	notech_or2 i_481(.A(n_818), .B(n_685), .Z(n_819));
	notech_and2 i_480(.A(n_686), .B(n_684), .Z(n_818));
	notech_inv i_299(.A(n_504), .Z(n_686));
	notech_inv i_298(.A(n_569), .Z(n_685));
	notech_inv i_479(.A(n_920), .Z(n_684));
	notech_nor2 i_478(.A(n_919), .B(n_862), .Z(n_920));
	notech_nor2 i_477(.A(n_683), .B(n_503), .Z(n_919));
	notech_inv i_476(.A(n_815), .Z(n_683));
	notech_or2 i_475(.A(n_814), .B(n_681), .Z(n_815));
	notech_and2 i_474(.A(n_682), .B(n_680), .Z(n_814));
	notech_inv i_295(.A(n_502), .Z(n_682));
	notech_inv i_294(.A(n_567), .Z(n_681));
	notech_inv i_473(.A(n_918), .Z(n_680));
	notech_nor2 i_472(.A(n_917), .B(n_861), .Z(n_918));
	notech_nor2 i_471(.A(n_679), .B(n_501), .Z(n_917));
	notech_inv i_470(.A(n_811), .Z(n_679));
	notech_or2 i_469(.A(n_810), .B(n_677), .Z(n_811));
	notech_and2 i_468(.A(n_678), .B(n_676), .Z(n_810));
	notech_inv i_291(.A(n_500), .Z(n_678));
	notech_inv i_290(.A(n_565), .Z(n_677));
	notech_inv i_467(.A(n_916), .Z(n_676));
	notech_nor2 i_466(.A(n_915), .B(n_860), .Z(n_916));
	notech_nor2 i_465(.A(n_675), .B(n_499), .Z(n_915));
	notech_inv i_464(.A(n_807), .Z(n_675));
	notech_or2 i_463(.A(n_806), .B(n_673), .Z(n_807));
	notech_and2 i_462(.A(n_674), .B(n_672), .Z(n_806));
	notech_inv i_287(.A(n_498), .Z(n_674));
	notech_inv i_286(.A(n_563), .Z(n_673));
	notech_inv i_461(.A(n_914), .Z(n_672));
	notech_nor2 i_460(.A(n_913), .B(n_859), .Z(n_914));
	notech_nor2 i_459(.A(n_671), .B(n_497), .Z(n_913));
	notech_inv i_458(.A(n_803), .Z(n_671));
	notech_or2 i_457(.A(n_802), .B(n_669), .Z(n_803));
	notech_and2 i_456(.A(n_670), .B(n_668), .Z(n_802));
	notech_inv i_283(.A(n_496), .Z(n_670));
	notech_inv i_282(.A(n_561), .Z(n_669));
	notech_inv i_455(.A(n_912), .Z(n_668));
	notech_nor2 i_454(.A(n_911), .B(n_858), .Z(n_912));
	notech_nor2 i_453(.A(n_667), .B(n_495), .Z(n_911));
	notech_inv i_452(.A(n_799), .Z(n_667));
	notech_or2 i_451(.A(n_798), .B(n_665), .Z(n_799));
	notech_and2 i_450(.A(n_666), .B(n_664), .Z(n_798));
	notech_inv i_279(.A(n_494), .Z(n_666));
	notech_inv i_278(.A(n_559), .Z(n_665));
	notech_inv i_449(.A(n_910), .Z(n_664));
	notech_nor2 i_448(.A(n_909), .B(n_857), .Z(n_910));
	notech_nor2 i_447(.A(n_663), .B(n_493), .Z(n_909));
	notech_inv i_446(.A(n_795), .Z(n_663));
	notech_or2 i_445(.A(n_794), .B(n_661), .Z(n_795));
	notech_and2 i_444(.A(n_662), .B(n_660), .Z(n_794));
	notech_inv i_275(.A(n_492), .Z(n_662));
	notech_inv i_274(.A(n_557), .Z(n_661));
	notech_inv i_443(.A(n_908), .Z(n_660));
	notech_nor2 i_442(.A(n_907), .B(n_856), .Z(n_908));
	notech_nor2 i_441(.A(n_659), .B(n_491), .Z(n_907));
	notech_inv i_440(.A(n_791), .Z(n_659));
	notech_or2 i_439(.A(n_790), .B(n_657), .Z(n_791));
	notech_and2 i_438(.A(n_658), .B(n_656), .Z(n_790));
	notech_inv i_271(.A(n_490), .Z(n_658));
	notech_inv i_270(.A(n_555), .Z(n_657));
	notech_inv i_437(.A(n_906), .Z(n_656));
	notech_nor2 i_436(.A(n_905), .B(n_855), .Z(n_906));
	notech_nor2 i_435(.A(n_655), .B(n_489), .Z(n_905));
	notech_inv i_434(.A(n_787), .Z(n_655));
	notech_or2 i_433(.A(n_786), .B(n_653), .Z(n_787));
	notech_and2 i_432(.A(n_654), .B(n_652), .Z(n_786));
	notech_inv i_267(.A(n_488), .Z(n_654));
	notech_inv i_266(.A(n_553), .Z(n_653));
	notech_inv i_431(.A(n_904), .Z(n_652));
	notech_nor2 i_430(.A(n_903), .B(n_854), .Z(n_904));
	notech_nor2 i_429(.A(n_651), .B(n_487), .Z(n_903));
	notech_inv i_428(.A(n_783), .Z(n_651));
	notech_or2 i_427(.A(n_782), .B(n_649), .Z(n_783));
	notech_and2 i_426(.A(n_650), .B(n_648), .Z(n_782));
	notech_inv i_263(.A(n_486), .Z(n_650));
	notech_inv i_262(.A(n_551), .Z(n_649));
	notech_inv i_425(.A(n_902), .Z(n_648));
	notech_nor2 i_424(.A(n_901), .B(n_853), .Z(n_902));
	notech_nor2 i_423(.A(n_647), .B(n_485), .Z(n_901));
	notech_inv i_422(.A(n_779), .Z(n_647));
	notech_or2 i_421(.A(n_778), .B(n_645), .Z(n_779));
	notech_and2 i_420(.A(n_646), .B(n_644), .Z(n_778));
	notech_inv i_259(.A(n_484), .Z(n_646));
	notech_inv i_258(.A(n_549), .Z(n_645));
	notech_inv i_419(.A(n_900), .Z(n_644));
	notech_nor2 i_418(.A(n_899), .B(n_852), .Z(n_900));
	notech_nor2 i_417(.A(n_643), .B(n_483), .Z(n_899));
	notech_inv i_416(.A(n_775), .Z(n_643));
	notech_or2 i_415(.A(n_774), .B(n_641), .Z(n_775));
	notech_and2 i_414(.A(n_642), .B(n_640), .Z(n_774));
	notech_inv i_255(.A(n_482), .Z(n_642));
	notech_inv i_254(.A(n_547), .Z(n_641));
	notech_inv i_413(.A(n_898), .Z(n_640));
	notech_nor2 i_412(.A(n_897), .B(n_851), .Z(n_898));
	notech_nor2 i_411(.A(n_639), .B(n_481), .Z(n_897));
	notech_inv i_410(.A(n_771), .Z(n_639));
	notech_or2 i_409(.A(n_770), .B(n_637), .Z(n_771));
	notech_and2 i_408(.A(n_638), .B(n_636), .Z(n_770));
	notech_inv i_251(.A(n_480), .Z(n_638));
	notech_inv i_250(.A(n_545), .Z(n_637));
	notech_inv i_407(.A(n_896), .Z(n_636));
	notech_nor2 i_406(.A(n_895), .B(n_850), .Z(n_896));
	notech_nor2 i_405(.A(n_635), .B(n_479), .Z(n_895));
	notech_inv i_404(.A(n_767), .Z(n_635));
	notech_or2 i_403(.A(n_766), .B(n_633), .Z(n_767));
	notech_and2 i_402(.A(n_634), .B(n_632), .Z(n_766));
	notech_inv i_247(.A(n_478), .Z(n_634));
	notech_inv i_246(.A(n_543), .Z(n_633));
	notech_inv i_401(.A(n_894), .Z(n_632));
	notech_nor2 i_400(.A(n_893), .B(n_849), .Z(n_894));
	notech_nor2 i_399(.A(n_631), .B(n_477), .Z(n_893));
	notech_inv i_398(.A(n_763), .Z(n_631));
	notech_or2 i_397(.A(n_762), .B(n_629), .Z(n_763));
	notech_and2 i_396(.A(n_630), .B(n_628), .Z(n_762));
	notech_inv i_243(.A(n_476), .Z(n_630));
	notech_inv i_242(.A(n_541), .Z(n_629));
	notech_inv i_395(.A(n_892), .Z(n_628));
	notech_nor2 i_394(.A(n_891), .B(n_848), .Z(n_892));
	notech_nor2 i_393(.A(n_627), .B(n_475), .Z(n_891));
	notech_inv i_392(.A(n_759), .Z(n_627));
	notech_or2 i_391(.A(n_758), .B(n_625), .Z(n_759));
	notech_and2 i_390(.A(n_626), .B(n_624), .Z(n_758));
	notech_inv i_239(.A(n_474), .Z(n_626));
	notech_inv i_238(.A(n_539), .Z(n_625));
	notech_inv i_389(.A(n_890), .Z(n_624));
	notech_nor2 i_388(.A(n_889), .B(n_847), .Z(n_890));
	notech_nor2 i_387(.A(n_623), .B(n_473), .Z(n_889));
	notech_inv i_386(.A(n_755), .Z(n_623));
	notech_or2 i_385(.A(n_754), .B(n_621), .Z(n_755));
	notech_and2 i_384(.A(n_622), .B(n_620), .Z(n_754));
	notech_inv i_235(.A(n_472), .Z(n_622));
	notech_inv i_234(.A(n_537), .Z(n_621));
	notech_inv i_383(.A(n_888), .Z(n_620));
	notech_nor2 i_382(.A(n_887), .B(n_846), .Z(n_888));
	notech_nor2 i_381(.A(n_619), .B(n_471), .Z(n_887));
	notech_inv i_380(.A(n_751), .Z(n_619));
	notech_or2 i_379(.A(n_750), .B(n_617), .Z(n_751));
	notech_and2 i_378(.A(n_618), .B(n_616), .Z(n_750));
	notech_inv i_231(.A(n_470), .Z(n_618));
	notech_inv i_230(.A(n_535), .Z(n_617));
	notech_inv i_377(.A(n_886), .Z(n_616));
	notech_nor2 i_376(.A(n_885), .B(n_845), .Z(n_886));
	notech_nor2 i_375(.A(n_615), .B(n_469), .Z(n_885));
	notech_inv i_374(.A(n_747), .Z(n_615));
	notech_or2 i_373(.A(n_746), .B(n_613), .Z(n_747));
	notech_and2 i_372(.A(n_614), .B(n_612), .Z(n_746));
	notech_inv i_227(.A(n_468), .Z(n_614));
	notech_inv i_226(.A(n_533), .Z(n_613));
	notech_inv i_371(.A(n_884), .Z(n_612));
	notech_nor2 i_370(.A(n_883), .B(n_844), .Z(n_884));
	notech_nor2 i_369(.A(n_611), .B(n_467), .Z(n_883));
	notech_inv i_368(.A(n_743), .Z(n_611));
	notech_or2 i_367(.A(n_742), .B(n_609), .Z(n_743));
	notech_and2 i_366(.A(n_610), .B(n_608), .Z(n_742));
	notech_inv i_223(.A(n_466), .Z(n_610));
	notech_inv i_222(.A(n_531), .Z(n_609));
	notech_inv i_365(.A(n_882), .Z(n_608));
	notech_nor2 i_364(.A(n_881), .B(n_843), .Z(n_882));
	notech_nor2 i_363(.A(n_607), .B(n_465), .Z(n_881));
	notech_inv i_362(.A(n_739), .Z(n_607));
	notech_or2 i_361(.A(n_738), .B(n_605), .Z(n_739));
	notech_and2 i_360(.A(n_606), .B(n_604), .Z(n_738));
	notech_inv i_219(.A(n_464), .Z(n_606));
	notech_inv i_218(.A(n_529), .Z(n_605));
	notech_inv i_359(.A(n_880), .Z(n_604));
	notech_nor2 i_358(.A(n_879), .B(n_842), .Z(n_880));
	notech_nor2 i_357(.A(n_603), .B(n_463), .Z(n_879));
	notech_inv i_356(.A(n_735), .Z(n_603));
	notech_or2 i_355(.A(n_734), .B(n_601), .Z(n_735));
	notech_and2 i_354(.A(n_602), .B(n_600), .Z(n_734));
	notech_inv i_215(.A(n_462), .Z(n_602));
	notech_inv i_214(.A(n_527), .Z(n_601));
	notech_inv i_353(.A(n_878), .Z(n_600));
	notech_nor2 i_352(.A(n_877), .B(n_841), .Z(n_878));
	notech_nor2 i_351(.A(n_599), .B(n_461), .Z(n_877));
	notech_inv i_350(.A(n_731), .Z(n_599));
	notech_or2 i_349(.A(n_730), .B(n_597), .Z(n_731));
	notech_and2 i_348(.A(n_598), .B(n_596), .Z(n_730));
	notech_inv i_211(.A(n_460), .Z(n_598));
	notech_inv i_210(.A(n_525), .Z(n_597));
	notech_inv i_347(.A(n_876), .Z(n_596));
	notech_nor2 i_346(.A(n_875), .B(n_840), .Z(n_876));
	notech_nor2 i_345(.A(n_595), .B(n_459), .Z(n_875));
	notech_inv i_344(.A(n_727), .Z(n_595));
	notech_or2 i_343(.A(n_726), .B(n_593), .Z(n_727));
	notech_and2 i_342(.A(n_594), .B(n_592), .Z(n_726));
	notech_inv i_207(.A(n_458), .Z(n_594));
	notech_inv i_206(.A(n_523), .Z(n_593));
	notech_inv i_341(.A(n_874), .Z(n_592));
	notech_nor2 i_340(.A(n_873), .B(n_839), .Z(n_874));
	notech_nor2 i_339(.A(n_591), .B(n_457), .Z(n_873));
	notech_inv i_338(.A(n_723), .Z(n_591));
	notech_or2 i_337(.A(n_722), .B(n_589), .Z(n_723));
	notech_and2 i_336(.A(n_590), .B(n_588), .Z(n_722));
	notech_inv i_203(.A(n_456), .Z(n_590));
	notech_inv i_202(.A(n_521), .Z(n_589));
	notech_inv i_335(.A(n_872), .Z(n_588));
	notech_nor2 i_334(.A(n_871), .B(n_838), .Z(n_872));
	notech_nor2 i_333(.A(n_587), .B(n_455), .Z(n_871));
	notech_inv i_332(.A(n_719), .Z(n_587));
	notech_or2 i_331(.A(n_718), .B(n_585), .Z(n_719));
	notech_and2 i_330(.A(n_586), .B(n_584), .Z(n_718));
	notech_inv i_199(.A(n_454), .Z(n_586));
	notech_inv i_198(.A(n_519), .Z(n_585));
	notech_inv i_329(.A(n_870), .Z(n_584));
	notech_nor2 i_328(.A(n_869), .B(n_837), .Z(n_870));
	notech_nor2 i_327(.A(n_583), .B(n_453), .Z(n_869));
	notech_inv i_326(.A(n_715), .Z(n_583));
	notech_or2 i_325(.A(n_714), .B(n_581), .Z(n_715));
	notech_and2 i_324(.A(n_582), .B(n_580), .Z(n_714));
	notech_inv i_195(.A(n_452), .Z(n_582));
	notech_inv i_194(.A(n_517), .Z(n_581));
	notech_inv i_323(.A(n_868), .Z(n_580));
	notech_nor2 i_322(.A(n_867), .B(n_836), .Z(n_868));
	notech_nor2 i_321(.A(n_451), .B(n_515), .Z(n_867));
	notech_inv i_191(.A(divq[63]), .Z(n_709));
	notech_nand2 i_190(.A(n_449), .B(divq[62]), .Z(n_577));
	notech_and2 i_189(.A(n_448), .B(divq[61]), .Z(n_866));
	notech_nand2 i_188(.A(n_447), .B(divq[60]), .Z(n_575));
	notech_and2 i_187(.A(n_446), .B(divq[59]), .Z(n_865));
	notech_nand2 i_186(.A(n_445), .B(divq[58]), .Z(n_573));
	notech_and2 i_185(.A(n_444), .B(divq[57]), .Z(n_864));
	notech_nand2 i_184(.A(n_443), .B(divq[56]), .Z(n_571));
	notech_and2 i_183(.A(n_442), .B(divq[55]), .Z(n_863));
	notech_nand2 i_182(.A(n_441), .B(divq[54]), .Z(n_569));
	notech_and2 i_181(.A(n_440), .B(divq[53]), .Z(n_862));
	notech_nand2 i_180(.A(n_439), .B(divq[52]), .Z(n_567));
	notech_and2 i_179(.A(n_438), .B(divq[51]), .Z(n_861));
	notech_nand2 i_178(.A(n_437), .B(divq[50]), .Z(n_565));
	notech_and2 i_177(.A(n_436), .B(divq[49]), .Z(n_860));
	notech_nand2 i_176(.A(n_435), .B(divq[48]), .Z(n_563));
	notech_and2 i_175(.A(n_434), .B(divq[47]), .Z(n_859));
	notech_nand2 i_174(.A(n_433), .B(divq[46]), .Z(n_561));
	notech_and2 i_173(.A(n_432), .B(divq[45]), .Z(n_858));
	notech_nand2 i_172(.A(n_431), .B(divq[44]), .Z(n_559));
	notech_and2 i_171(.A(n_430), .B(divq[43]), .Z(n_857));
	notech_nand2 i_170(.A(n_429), .B(divq[42]), .Z(n_557));
	notech_and2 i_169(.A(n_428), .B(divq[41]), .Z(n_856));
	notech_nand2 i_168(.A(n_427), .B(divq[40]), .Z(n_555));
	notech_and2 i_167(.A(n_426), .B(divq[39]), .Z(n_855));
	notech_nand2 i_166(.A(n_425), .B(divq[38]), .Z(n_553));
	notech_and2 i_165(.A(n_424), .B(divq[37]), .Z(n_854));
	notech_nand2 i_164(.A(n_423), .B(divq[36]), .Z(n_551));
	notech_and2 i_163(.A(n_422), .B(divq[35]), .Z(n_853));
	notech_nand2 i_162(.A(n_421), .B(divq[34]), .Z(n_549));
	notech_and2 i_161(.A(n_420), .B(divq[33]), .Z(n_852));
	notech_nand2 i_160(.A(n_419), .B(divq[32]), .Z(n_547));
	notech_and2 i_159(.A(n_418), .B(divq[31]), .Z(n_851));
	notech_nand2 i_158(.A(n_417), .B(divq[30]), .Z(n_545));
	notech_and2 i_157(.A(n_416), .B(divq[29]), .Z(n_850));
	notech_nand2 i_156(.A(n_415), .B(divq[28]), .Z(n_543));
	notech_and2 i_155(.A(n_414), .B(divq[27]), .Z(n_849));
	notech_nand2 i_154(.A(n_413), .B(divq[26]), .Z(n_541));
	notech_and2 i_153(.A(n_412), .B(divq[25]), .Z(n_848));
	notech_nand2 i_152(.A(n_411), .B(divq[24]), .Z(n_539));
	notech_and2 i_151(.A(n_410), .B(divq[23]), .Z(n_847));
	notech_nand2 i_150(.A(n_409), .B(divq[22]), .Z(n_537));
	notech_and2 i_149(.A(n_408), .B(divq[21]), .Z(n_846));
	notech_nand2 i_148(.A(n_407), .B(divq[20]), .Z(n_535));
	notech_and2 i_147(.A(n_406), .B(divq[19]), .Z(n_845));
	notech_nand2 i_146(.A(n_405), .B(divq[18]), .Z(n_533));
	notech_and2 i_145(.A(n_404), .B(divq[17]), .Z(n_844));
	notech_nand2 i_144(.A(n_403), .B(divq[16]), .Z(n_531));
	notech_and2 i_143(.A(n_402), .B(divq[15]), .Z(n_843));
	notech_nand2 i_142(.A(n_401), .B(divq[14]), .Z(n_529));
	notech_and2 i_141(.A(n_400), .B(divq[13]), .Z(n_842));
	notech_nand2 i_140(.A(n_399), .B(divq[12]), .Z(n_527));
	notech_and2 i_139(.A(n_398), .B(divq[11]), .Z(n_841));
	notech_nand2 i_138(.A(n_397), .B(divq[10]), .Z(n_525));
	notech_and2 i_137(.A(n_396), .B(divq[9]), .Z(n_840));
	notech_nand2 i_136(.A(n_395), .B(divq[8]), .Z(n_523));
	notech_and2 i_135(.A(n_394), .B(divq[7]), .Z(n_839));
	notech_nand2 i_134(.A(n_393), .B(divq[6]), .Z(n_521));
	notech_and2 i_133(.A(n_392), .B(divq[5]), .Z(n_838));
	notech_nand2 i_132(.A(n_391), .B(divq[4]), .Z(n_519));
	notech_and2 i_131(.A(n_390), .B(divq[3]), .Z(n_837));
	notech_nand2 i_130(.A(n_389), .B(divq[2]), .Z(n_517));
	notech_and2 i_129(.A(n_388), .B(divq[1]), .Z(n_836));
	notech_nand2 i_128(.A(n_387), .B(divq[0]), .Z(n_515));
	notech_nor2 i_125(.A(n_449), .B(divq[62]), .Z(n_512));
	notech_nor2 i_124(.A(n_448), .B(divq[61]), .Z(n_511));
	notech_nor2 i_123(.A(n_447), .B(divq[60]), .Z(n_510));
	notech_nor2 i_122(.A(n_446), .B(divq[59]), .Z(n_509));
	notech_nor2 i_121(.A(n_445), .B(divq[58]), .Z(n_508));
	notech_nor2 i_120(.A(n_444), .B(divq[57]), .Z(n_507));
	notech_nor2 i_119(.A(n_443), .B(divq[56]), .Z(n_506));
	notech_nor2 i_118(.A(n_442), .B(divq[55]), .Z(n_505));
	notech_nor2 i_117(.A(n_441), .B(divq[54]), .Z(n_504));
	notech_nor2 i_116(.A(n_440), .B(divq[53]), .Z(n_503));
	notech_nor2 i_115(.A(n_439), .B(divq[52]), .Z(n_502));
	notech_nor2 i_114(.A(n_438), .B(divq[51]), .Z(n_501));
	notech_nor2 i_113(.A(n_437), .B(divq[50]), .Z(n_500));
	notech_nor2 i_112(.A(n_436), .B(divq[49]), .Z(n_499));
	notech_nor2 i_111(.A(n_435), .B(divq[48]), .Z(n_498));
	notech_nor2 i_110(.A(n_434), .B(divq[47]), .Z(n_497));
	notech_nor2 i_109(.A(n_433), .B(divq[46]), .Z(n_496));
	notech_nor2 i_108(.A(n_432), .B(divq[45]), .Z(n_495));
	notech_nor2 i_107(.A(n_431), .B(divq[44]), .Z(n_494));
	notech_nor2 i_106(.A(n_430), .B(divq[43]), .Z(n_493));
	notech_nor2 i_105(.A(n_429), .B(divq[42]), .Z(n_492));
	notech_nor2 i_104(.A(n_428), .B(divq[41]), .Z(n_491));
	notech_nor2 i_103(.A(n_427), .B(divq[40]), .Z(n_490));
	notech_nor2 i_102(.A(n_426), .B(divq[39]), .Z(n_489));
	notech_nor2 i_101(.A(n_425), .B(divq[38]), .Z(n_488));
	notech_nor2 i_100(.A(n_424), .B(divq[37]), .Z(n_487));
	notech_nor2 i_99(.A(n_423), .B(divq[36]), .Z(n_486));
	notech_nor2 i_98(.A(n_422), .B(divq[35]), .Z(n_485));
	notech_nor2 i_97(.A(n_421), .B(divq[34]), .Z(n_484));
	notech_nor2 i_96(.A(n_420), .B(divq[33]), .Z(n_483));
	notech_nor2 i_95(.A(n_419), .B(divq[32]), .Z(n_482));
	notech_nor2 i_94(.A(n_418), .B(divq[31]), .Z(n_481));
	notech_nor2 i_93(.A(n_417), .B(divq[30]), .Z(n_480));
	notech_nor2 i_92(.A(n_416), .B(divq[29]), .Z(n_479));
	notech_nor2 i_91(.A(n_415), .B(divq[28]), .Z(n_478));
	notech_nor2 i_90(.A(n_414), .B(divq[27]), .Z(n_477));
	notech_nor2 i_89(.A(n_413), .B(divq[26]), .Z(n_476));
	notech_nor2 i_88(.A(n_412), .B(divq[25]), .Z(n_475));
	notech_nor2 i_87(.A(n_411), .B(divq[24]), .Z(n_474));
	notech_nor2 i_86(.A(n_410), .B(divq[23]), .Z(n_473));
	notech_nor2 i_85(.A(n_409), .B(divq[22]), .Z(n_472));
	notech_nor2 i_84(.A(n_408), .B(divq[21]), .Z(n_471));
	notech_nor2 i_83(.A(n_407), .B(divq[20]), .Z(n_470));
	notech_nor2 i_82(.A(n_406), .B(divq[19]), .Z(n_469));
	notech_nor2 i_81(.A(n_405), .B(divq[18]), .Z(n_468));
	notech_nor2 i_80(.A(n_404), .B(divq[17]), .Z(n_467));
	notech_nor2 i_79(.A(n_403), .B(divq[16]), .Z(n_466));
	notech_nor2 i_78(.A(n_402), .B(divq[15]), .Z(n_465));
	notech_nor2 i_77(.A(n_401), .B(divq[14]), .Z(n_464));
	notech_nor2 i_76(.A(n_400), .B(divq[13]), .Z(n_463));
	notech_nor2 i_75(.A(n_399), .B(divq[12]), .Z(n_462));
	notech_nor2 i_74(.A(n_398), .B(divq[11]), .Z(n_461));
	notech_nor2 i_73(.A(n_397), .B(divq[10]), .Z(n_460));
	notech_nor2 i_72(.A(n_396), .B(divq[9]), .Z(n_459));
	notech_nor2 i_71(.A(n_395), .B(divq[8]), .Z(n_458));
	notech_nor2 i_70(.A(n_394), .B(divq[7]), .Z(n_457));
	notech_nor2 i_69(.A(n_393), .B(divq[6]), .Z(n_456));
	notech_nor2 i_68(.A(n_392), .B(divq[5]), .Z(n_455));
	notech_nor2 i_67(.A(n_391), .B(divq[4]), .Z(n_454));
	notech_nor2 i_66(.A(n_390), .B(divq[3]), .Z(n_453));
	notech_nor2 i_65(.A(n_389), .B(divq[2]), .Z(n_452));
	notech_nor2 i_64(.A(n_388), .B(divq[1]), .Z(n_451));
	notech_inv i_62(.A(I0[62]), .Z(n_449));
	notech_inv i_61(.A(I0[61]), .Z(n_448));
	notech_inv i_60(.A(I0[60]), .Z(n_447));
	notech_inv i_59(.A(I0[59]), .Z(n_446));
	notech_inv i_58(.A(I0[58]), .Z(n_445));
	notech_inv i_57(.A(I0[57]), .Z(n_444));
	notech_inv i_56(.A(I0[56]), .Z(n_443));
	notech_inv i_55(.A(I0[55]), .Z(n_442));
	notech_inv i_54(.A(I0[54]), .Z(n_441));
	notech_inv i_53(.A(I0[53]), .Z(n_440));
	notech_inv i_52(.A(I0[52]), .Z(n_439));
	notech_inv i_51(.A(I0[51]), .Z(n_438));
	notech_inv i_50(.A(I0[50]), .Z(n_437));
	notech_inv i_49(.A(I0[49]), .Z(n_436));
	notech_inv i_48(.A(I0[48]), .Z(n_435));
	notech_inv i_47(.A(I0[47]), .Z(n_434));
	notech_inv i_46(.A(I0[46]), .Z(n_433));
	notech_inv i_45(.A(I0[45]), .Z(n_432));
	notech_inv i_44(.A(I0[44]), .Z(n_431));
	notech_inv i_43(.A(I0[43]), .Z(n_430));
	notech_inv i_42(.A(I0[42]), .Z(n_429));
	notech_inv i_41(.A(I0[41]), .Z(n_428));
	notech_inv i_40(.A(I0[40]), .Z(n_427));
	notech_inv i_39(.A(I0[39]), .Z(n_426));
	notech_inv i_38(.A(I0[38]), .Z(n_425));
	notech_inv i_37(.A(I0[37]), .Z(n_424));
	notech_inv i_36(.A(I0[36]), .Z(n_423));
	notech_inv i_35(.A(I0[35]), .Z(n_422));
	notech_inv i_34(.A(I0[34]), .Z(n_421));
	notech_inv i_33(.A(I0[33]), .Z(n_420));
	notech_inv i_32(.A(I0[32]), .Z(n_419));
	notech_inv i_31(.A(I0[31]), .Z(n_418));
	notech_inv i_30(.A(I0[30]), .Z(n_417));
	notech_inv i_29(.A(I0[29]), .Z(n_416));
	notech_inv i_28(.A(I0[28]), .Z(n_415));
	notech_inv i_27(.A(I0[27]), .Z(n_414));
	notech_inv i_26(.A(I0[26]), .Z(n_413));
	notech_inv i_25(.A(I0[25]), .Z(n_412));
	notech_inv i_24(.A(I0[24]), .Z(n_411));
	notech_inv i_23(.A(I0[23]), .Z(n_410));
	notech_inv i_22(.A(I0[22]), .Z(n_409));
	notech_inv i_21(.A(I0[21]), .Z(n_408));
	notech_inv i_20(.A(I0[20]), .Z(n_407));
	notech_inv i_19(.A(I0[19]), .Z(n_406));
	notech_inv i_18(.A(I0[18]), .Z(n_405));
	notech_inv i_17(.A(I0[17]), .Z(n_404));
	notech_inv i_16(.A(I0[16]), .Z(n_403));
	notech_inv i_15(.A(I0[15]), .Z(n_402));
	notech_inv i_14(.A(I0[14]), .Z(n_401));
	notech_inv i_13(.A(I0[13]), .Z(n_400));
	notech_inv i_12(.A(I0[12]), .Z(n_399));
	notech_inv i_11(.A(I0[11]), .Z(n_398));
	notech_inv i_10(.A(I0[10]), .Z(n_397));
	notech_inv i_9(.A(I0[9]), .Z(n_396));
	notech_inv i_8(.A(I0[8]), .Z(n_395));
	notech_inv i_7(.A(I0[7]), .Z(n_394));
	notech_inv i_6(.A(I0[6]), .Z(n_393));
	notech_inv i_5(.A(I0[5]), .Z(n_392));
	notech_inv i_4(.A(I0[4]), .Z(n_391));
	notech_inv i_3(.A(I0[3]), .Z(n_390));
	notech_inv i_2(.A(I0[2]), .Z(n_389));
	notech_inv i_1(.A(I0[1]), .Z(n_388));
	notech_inv i_0(.A(I0[0]), .Z(n_387));
endmodule
module AWDP_LSH_196(O0, opd);
    output [31:0] O0;
    input [5:0] opd;
    wire [31:0] O0;
    // Line 1006
    wire [31:0] N769;

    assign O0 = N769;
    // Line 1006
    assign N769 = 6'h1 << opd;
endmodule

module AWDP_LSH_43(O0, opb);
    output [31:0] O0;
    input [4:0] opb;
    // Line 348
    wire [31:0] O0;
    // Line 636
    wire [31:0] N785;

    // Line 348
    assign O0 = N785;
    // Line 636
    assign N785 = 5'h1 << opb;
endmodule

module AWDP_SUB_17(O0, regs_6, opd);
    output [31:0] O0;
    input [31:0] regs_6;
    input [31:0] opd;
    // Line 521
    wire [31:0] N800;
    // Line 348
    wire [31:0] O0;

    // Line 521
    assign N800 = regs_6 - opd;
    // Line 348
    assign O0 = N800;
endmodule

module AWDP_SUB_174(O0, divr, divq);
    output [63:0] O0;
    input [63:0] divr;
    input [63:0] divq;
    // Line 1006
    wire [63:0] N810;
    // Line 1006
    wire [63:0] O0;

    // Line 1006
    assign N810 = divr - divq;
    // Line 1006
    assign O0 = N810;
endmodule

module AWDP_SUB_200(O0, opd);

	output [31:0] O0;
	input [31:0] opd;

	wire \opd[2] ;
	wire \opd[3] ;
	wire \opd[4] ;
	wire \opd[5] ;
	wire \opd[6] ;
	wire \opd[7] ;
	wire \opd[8] ;
	wire \opd[9] ;
	wire \opd[10] ;
	wire \opd[11] ;
	wire \opd[12] ;
	wire \opd[13] ;
	wire \opd[14] ;
	wire \opd[15] ;
	wire \opd[16] ;
	wire \opd[17] ;
	wire \opd[18] ;
	wire \opd[19] ;
	wire \opd[20] ;
	wire \opd[21] ;
	wire \opd[22] ;
	wire \opd[23] ;
	wire \opd[24] ;
	wire \opd[25] ;
	wire \opd[26] ;
	wire \opd[27] ;
	wire \opd[28] ;
	wire \opd[29] ;
	wire \opd[30] ;
	wire \opd[31] ;


	assign O0[0] = opd[0];
	assign O0[1] = opd[1];
	assign \opd[2]  = opd[2];
	assign \opd[3]  = opd[3];
	assign \opd[4]  = opd[4];
	assign \opd[5]  = opd[5];
	assign \opd[6]  = opd[6];
	assign \opd[7]  = opd[7];
	assign \opd[8]  = opd[8];
	assign \opd[9]  = opd[9];
	assign \opd[10]  = opd[10];
	assign \opd[11]  = opd[11];
	assign \opd[12]  = opd[12];
	assign \opd[13]  = opd[13];
	assign \opd[14]  = opd[14];
	assign \opd[15]  = opd[15];
	assign \opd[16]  = opd[16];
	assign \opd[17]  = opd[17];
	assign \opd[18]  = opd[18];
	assign \opd[19]  = opd[19];
	assign \opd[20]  = opd[20];
	assign \opd[21]  = opd[21];
	assign \opd[22]  = opd[22];
	assign \opd[23]  = opd[23];
	assign \opd[24]  = opd[24];
	assign \opd[25]  = opd[25];
	assign \opd[26]  = opd[26];
	assign \opd[27]  = opd[27];
	assign \opd[28]  = opd[28];
	assign \opd[29]  = opd[29];
	assign \opd[30]  = opd[30];
	assign \opd[31]  = opd[31];

	notech_ha2 i_30(.A(n_192), .B(n_250), .Z(O0[31]));
	notech_inv i_1(.A(\opd[2] ), .Z(O0[2]));
	notech_inv i_0(.A(\opd[31] ), .Z(n_192));
	notech_xor2 i_47(.A(\opd[30] ), .B(n_248), .Z(n_45100));
	notech_inv i_48(.A(n_45100), .Z(O0[30]));
	notech_or2 i_46(.A(\opd[30] ), .B(n_248), .Z(n_250));
	notech_xor2 i_4695223(.A(\opd[29] ), .B(n_246), .Z(n_45127));
	notech_inv i_4795224(.A(n_45127), .Z(O0[29]));
	notech_or2 i_45(.A(\opd[29] ), .B(n_246), .Z(n_248));
	notech_xor2 i_44(.A(\opd[28] ), .B(n_244), .Z(n_45154));
	notech_inv i_4595225(.A(n_45154), .Z(O0[28]));
	notech_or2 i_43(.A(\opd[28] ), .B(n_244), .Z(n_246));
	notech_xor2 i_4395226(.A(\opd[27] ), .B(n_242), .Z(n_45181));
	notech_inv i_4495227(.A(n_45181), .Z(O0[27]));
	notech_or2 i_42(.A(\opd[27] ), .B(n_242), .Z(n_244));
	notech_xor2 i_4295228(.A(\opd[26] ), .B(n_240), .Z(n_45208));
	notech_inv i_4395229(.A(n_45208), .Z(O0[26]));
	notech_or2 i_41(.A(\opd[26] ), .B(n_240), .Z(n_242));
	notech_xor2 i_4195230(.A(\opd[25] ), .B(n_238), .Z(n_45235));
	notech_inv i_4295231(.A(n_45235), .Z(O0[25]));
	notech_or2 i_40(.A(\opd[25] ), .B(n_238), .Z(n_240));
	notech_xor2 i_4095232(.A(\opd[24] ), .B(n_236), .Z(n_45262));
	notech_inv i_4195233(.A(n_45262), .Z(O0[24]));
	notech_or2 i_39(.A(\opd[24] ), .B(n_236), .Z(n_238));
	notech_xor2 i_3995234(.A(\opd[23] ), .B(n_234), .Z(n_45289));
	notech_inv i_4095235(.A(n_45289), .Z(O0[23]));
	notech_or2 i_38(.A(\opd[23] ), .B(n_234), .Z(n_236));
	notech_xor2 i_3895236(.A(\opd[22] ), .B(n_232), .Z(n_45316));
	notech_inv i_3995237(.A(n_45316), .Z(O0[22]));
	notech_or2 i_37(.A(\opd[22] ), .B(n_232), .Z(n_234));
	notech_xor2 i_3795238(.A(\opd[21] ), .B(n_230), .Z(n_45343));
	notech_inv i_3895239(.A(n_45343), .Z(O0[21]));
	notech_or2 i_36(.A(\opd[21] ), .B(n_230), .Z(n_232));
	notech_xor2 i_3695240(.A(\opd[20] ), .B(n_228), .Z(n_45370));
	notech_inv i_3795241(.A(n_45370), .Z(O0[20]));
	notech_or2 i_35(.A(\opd[20] ), .B(n_228), .Z(n_230));
	notech_xor2 i_3595242(.A(\opd[19] ), .B(n_226), .Z(n_45397));
	notech_inv i_3695243(.A(n_45397), .Z(O0[19]));
	notech_or2 i_34(.A(\opd[19] ), .B(n_226), .Z(n_228));
	notech_xor2 i_3495244(.A(\opd[18] ), .B(n_224), .Z(n_45424));
	notech_inv i_3595245(.A(n_45424), .Z(O0[18]));
	notech_or2 i_33(.A(\opd[18] ), .B(n_224), .Z(n_226));
	notech_xor2 i_3395246(.A(\opd[17] ), .B(n_222), .Z(n_45451));
	notech_inv i_3495247(.A(n_45451), .Z(O0[17]));
	notech_or2 i_32(.A(\opd[17] ), .B(n_222), .Z(n_224));
	notech_xor2 i_3295248(.A(\opd[16] ), .B(n_220), .Z(n_45478));
	notech_inv i_3395249(.A(n_45478), .Z(O0[16]));
	notech_or2 i_31(.A(\opd[16] ), .B(n_220), .Z(n_222));
	notech_xor2 i_3195250(.A(\opd[15] ), .B(n_218), .Z(n_45505));
	notech_inv i_3295251(.A(n_45505), .Z(O0[15]));
	notech_or2 i_3095252(.A(\opd[15] ), .B(n_218), .Z(n_220));
	notech_xor2 i_3095253(.A(\opd[14] ), .B(n_216), .Z(n_45532));
	notech_inv i_3195254(.A(n_45532), .Z(O0[14]));
	notech_or2 i_29(.A(\opd[14] ), .B(n_216), .Z(n_218));
	notech_xor2 i_2995255(.A(\opd[13] ), .B(n_214), .Z(n_45559));
	notech_inv i_3095256(.A(n_45559), .Z(O0[13]));
	notech_or2 i_28(.A(\opd[13] ), .B(n_214), .Z(n_216));
	notech_xor2 i_2895257(.A(\opd[12] ), .B(n_212), .Z(n_45586));
	notech_inv i_2995258(.A(n_45586), .Z(O0[12]));
	notech_or2 i_27(.A(\opd[12] ), .B(n_212), .Z(n_214));
	notech_xor2 i_2795259(.A(\opd[11] ), .B(n_210), .Z(n_45613));
	notech_inv i_2895260(.A(n_45613), .Z(O0[11]));
	notech_or2 i_26(.A(\opd[11] ), .B(n_210), .Z(n_212));
	notech_xor2 i_2795261(.A(\opd[10] ), .B(n_208), .Z(n_45640));
	notech_inv i_2895262(.A(n_45640), .Z(O0[10]));
	notech_or2 i_2695263(.A(\opd[10] ), .B(n_208), .Z(n_210));
	notech_xor2 i_2795264(.A(\opd[9] ), .B(n_206), .Z(n_45667));
	notech_inv i_2895265(.A(n_45667), .Z(O0[9]));
	notech_or2 i_2695266(.A(\opd[9] ), .B(n_206), .Z(n_208));
	notech_xor2 i_2795267(.A(\opd[8] ), .B(n_204), .Z(n_45694));
	notech_inv i_2895268(.A(n_45694), .Z(O0[8]));
	notech_or2 i_2695269(.A(\opd[8] ), .B(n_204), .Z(n_206));
	notech_xor2 i_2795270(.A(\opd[7] ), .B(n_202), .Z(n_45721));
	notech_inv i_2895271(.A(n_45721), .Z(O0[7]));
	notech_or2 i_2695272(.A(\opd[7] ), .B(n_202), .Z(n_204));
	notech_xor2 i_2795273(.A(\opd[6] ), .B(n_200), .Z(n_45748));
	notech_inv i_2895274(.A(n_45748), .Z(O0[6]));
	notech_or2 i_2695275(.A(\opd[6] ), .B(n_200), .Z(n_202));
	notech_xor2 i_2795276(.A(\opd[5] ), .B(n_198), .Z(n_45775));
	notech_inv i_2895277(.A(n_45775), .Z(O0[5]));
	notech_or2 i_2695278(.A(\opd[5] ), .B(n_198), .Z(n_200));
	notech_xor2 i_2795279(.A(\opd[4] ), .B(n_196), .Z(n_45802));
	notech_inv i_2895280(.A(n_45802), .Z(O0[4]));
	notech_or2 i_2695281(.A(\opd[4] ), .B(n_196), .Z(n_198));
	notech_xor2 i_2795282(.A(\opd[3] ), .B(\opd[2] ), .Z(n_45830));
	notech_inv i_2895283(.A(n_45830), .Z(O0[3]));
	notech_or2 i_2695284(.A(\opd[3] ), .B(\opd[2] ), .Z(n_196));
endmodule
module AWDP_SUB_205(O0, opa, I0);

	output [16:0] O0;
	input [15:0] opa;
	input [15:0] I0;




	notech_inv i_10736(.A(I0[13]), .Z(n_56982));
	notech_inv i_32(.A(n_230), .Z(O0[16]));
	notech_fa2 i_31(.A(n_56982), .B(n_228), .CI(opa[15]), .Z(O0[15]), .CO(n_230
		));
	notech_fa2 i_30(.A(n_56982), .B(n_226), .CI(opa[14]), .Z(O0[14]), .CO(n_228
		));
	notech_fa2 i_29(.A(n_56982), .B(n_224), .CI(opa[13]), .Z(O0[13]), .CO(n_226
		));
	notech_fa2 i_28(.A(n_56982), .B(n_222), .CI(opa[12]), .Z(O0[12]), .CO(n_224
		));
	notech_fa2 i_27(.A(n_56982), .B(n_220), .CI(opa[11]), .Z(O0[11]), .CO(n_222
		));
	notech_fa2 i_26(.A(n_56982), .B(n_218), .CI(opa[10]), .Z(O0[10]), .CO(n_220
		));
	notech_fa2 i_25(.A(n_56982), .B(n_216), .CI(opa[9]), .Z(O0[9]), .CO(n_218
		));
	notech_fa2 i_24(.A(n_56982), .B(n_214), .CI(opa[8]), .Z(O0[8]), .CO(n_216
		));
	notech_fa2 i_23(.A(n_56982), .B(n_212), .CI(opa[7]), .Z(O0[7]), .CO(n_214
		));
	notech_fa2 i_22(.A(n_56982), .B(n_210), .CI(opa[6]), .Z(O0[6]), .CO(n_212
		));
	notech_fa2 i_21(.A(n_56982), .B(n_208), .CI(opa[5]), .Z(O0[5]), .CO(n_210
		));
	notech_fa2 i_20(.A(n_56982), .B(n_206), .CI(opa[4]), .Z(O0[4]), .CO(n_208
		));
	notech_fa2 i_19(.A(n_56982), .B(n_204), .CI(opa[3]), .Z(O0[3]), .CO(n_206
		));
	notech_fa2 i_18(.A(n_56982), .B(n_202), .CI(opa[2]), .Z(O0[2]), .CO(n_204
		));
	notech_fa2 i_17(.A(n_184), .B(n_200), .CI(opa[1]), .Z(O0[1]), .CO(n_202)
		);
	notech_inv i_1(.A(I0[1]), .Z(n_184));
	notech_inv i_0(.A(I0[0]), .Z(n_183));
	notech_xor2 i_49(.A(opa[0]), .B(n_183), .Z(n_45857));
	notech_inv i_50(.A(n_45857), .Z(O0[0]));
	notech_or2 i_48(.A(opa[0]), .B(n_183), .Z(n_200));
endmodule
module AWDP_SUB_233(O0, regs_4, calc_sz);
    output [31:0] O0;
    input [31:0] regs_4;
    input [2:0] calc_sz;
    // Line 456
    wire [31:0] N841;
    // Line 348
    wire [31:0] O0;

    // Line 456
    assign N841 = regs_4 - calc_sz;
    // Line 348
    assign O0 = N841;
endmodule

module AWDP_SUB_29(O0, regs_7, opd);
    output [31:0] O0;
    input [31:0] regs_7;
    input [31:0] opd;
    // Line 521
    wire [31:0] N860;
    // Line 348
    wire [31:0] O0;

    // Line 521
    assign N860 = regs_7 - opd;
    // Line 348
    assign O0 = N860;
endmodule

module AWDP_SUB_41(O0, opa, I0);

	output [32:0] O0;
	input [31:0] opa;
	input [31:0] I0;




	notech_inv i_10759(.A(n_57078), .Z(n_57079));
	notech_inv i_10758(.A(I0[19]), .Z(n_57078));
	notech_inv i_64(.A(n_454), .Z(O0[32]));
	notech_fa2 i_63(.A(n_57078), .B(n_452), .CI(opa[31]), .Z(O0[31]), .CO(n_454
		));
	notech_fa2 i_62(.A(n_57078), .B(n_450), .CI(opa[30]), .Z(O0[30]), .CO(n_452
		));
	notech_fa2 i_61(.A(n_57078), .B(n_448), .CI(opa[29]), .Z(O0[29]), .CO(n_450
		));
	notech_fa2 i_60(.A(n_57078), .B(n_446), .CI(opa[28]), .Z(O0[28]), .CO(n_448
		));
	notech_fa2 i_59(.A(n_57078), .B(n_444), .CI(opa[27]), .Z(O0[27]), .CO(n_446
		));
	notech_fa2 i_58(.A(n_57078), .B(n_442), .CI(opa[26]), .Z(O0[26]), .CO(n_444
		));
	notech_fa2 i_57(.A(n_57078), .B(n_440), .CI(opa[25]), .Z(O0[25]), .CO(n_442
		));
	notech_fa2 i_56(.A(n_57078), .B(n_438), .CI(opa[24]), .Z(O0[24]), .CO(n_440
		));
	notech_fa2 i_55(.A(n_57078), .B(n_436), .CI(opa[23]), .Z(O0[23]), .CO(n_438
		));
	notech_fa2 i_54(.A(n_57078), .B(n_434), .CI(opa[22]), .Z(O0[22]), .CO(n_436
		));
	notech_fa2 i_53(.A(n_57078), .B(n_432), .CI(opa[21]), .Z(O0[21]), .CO(n_434
		));
	notech_fa2 i_52(.A(n_57078), .B(n_430), .CI(opa[20]), .Z(O0[20]), .CO(n_432
		));
	notech_fa2 i_51(.A(n_57078), .B(n_428), .CI(opa[19]), .Z(O0[19]), .CO(n_430
		));
	notech_fa2 i_50(.A(n_57078), .B(n_426), .CI(opa[18]), .Z(O0[18]), .CO(n_428
		));
	notech_fa2 i_49(.A(n_57078), .B(n_424), .CI(opa[17]), .Z(O0[17]), .CO(n_426
		));
	notech_fa2 i_48(.A(n_361), .B(n_422), .CI(opa[16]), .Z(O0[16]), .CO(n_424
		));
	notech_fa2 i_47(.A(n_361), .B(n_420), .CI(opa[15]), .Z(O0[15]), .CO(n_422
		));
	notech_fa2 i_46(.A(n_361), .B(n_418), .CI(opa[14]), .Z(O0[14]), .CO(n_420
		));
	notech_fa2 i_45(.A(n_361), .B(n_416), .CI(opa[13]), .Z(O0[13]), .CO(n_418
		));
	notech_fa2 i_44(.A(n_361), .B(n_414), .CI(opa[12]), .Z(O0[12]), .CO(n_416
		));
	notech_fa2 i_43(.A(n_361), .B(n_412), .CI(opa[11]), .Z(O0[11]), .CO(n_414
		));
	notech_fa2 i_42(.A(n_361), .B(n_410), .CI(opa[10]), .Z(O0[10]), .CO(n_412
		));
	notech_fa2 i_41(.A(n_361), .B(n_408), .CI(opa[9]), .Z(O0[9]), .CO(n_410)
		);
	notech_fa2 i_40(.A(n_361), .B(n_406), .CI(opa[8]), .Z(O0[8]), .CO(n_408)
		);
	notech_fa2 i_39(.A(n_361), .B(n_404), .CI(opa[7]), .Z(O0[7]), .CO(n_406)
		);
	notech_fa2 i_38(.A(n_361), .B(n_402), .CI(opa[6]), .Z(O0[6]), .CO(n_404)
		);
	notech_fa2 i_37(.A(n_361), .B(n_400), .CI(opa[5]), .Z(O0[5]), .CO(n_402)
		);
	notech_fa2 i_36(.A(n_361), .B(n_398), .CI(opa[4]), .Z(O0[4]), .CO(n_400)
		);
	notech_fa2 i_35(.A(n_361), .B(n_396), .CI(opa[3]), .Z(O0[3]), .CO(n_398)
		);
	notech_fa2 i_34(.A(n_361), .B(n_394), .CI(opa[2]), .Z(O0[2]), .CO(n_396)
		);
	notech_fa2 i_33(.A(n_360), .B(n_392), .CI(opa[1]), .Z(O0[1]), .CO(n_394)
		);
	notech_inv i_2(.A(n_57079), .Z(n_361));
	notech_inv i_1(.A(I0[1]), .Z(n_360));
	notech_inv i_0(.A(I0[0]), .Z(n_359));
	notech_xor2 i_81(.A(opa[0]), .B(n_359), .Z(n_46694));
	notech_inv i_82(.A(n_46694), .Z(O0[0]));
	notech_or2 i_80(.A(opa[0]), .B(n_359), .Z(n_392));
endmodule
module AWMUX_16_1(I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14
		, I15, S, O0);

	input I0;
	input I1;
	input I2;
	input I3;
	input I4;
	input I5;
	input I6;
	input I7;
	input I8;
	input I9;
	input I10;
	input I11;
	input I12;
	input I13;
	input I14;
	input I15;
	input [3:0] S;
	output O0;




	notech_mux4 i_14(.S0(S[2]), .S1(S[3]), .A(n_23), .B(n_26), .C(n_29), .D(n_32
		), .Z(O0));
	notech_mux4 i_11(.S0(S[0]), .S1(S[1]), .A(I12), .B(n_14555), .C(I14), .D
		(n_14554), .Z(n_32));
	notech_mux4 i_8(.S0(S[0]), .S1(S[1]), .A(I8), .B(n_14557), .C(I10), .D(n_14556
		), .Z(n_29));
	notech_mux4 i_5(.S0(S[0]), .S1(S[1]), .A(I4), .B(n_14559), .C(I6), .D(n_14558
		), .Z(n_26));
	notech_mux4 i_2(.S0(S[0]), .S1(S[1]), .A(I0), .B(n_14561), .C(I2), .D(n_14560
		), .Z(n_23));
	notech_inv i_28(.A(I14), .Z(n_14554));
	notech_inv i_29(.A(I12), .Z(n_14555));
	notech_inv i_30(.A(I10), .Z(n_14556));
	notech_inv i_31(.A(I8), .Z(n_14557));
	notech_inv i_32(.A(I6), .Z(n_14558));
	notech_inv i_33(.A(I4), .Z(n_14559));
	notech_inv i_34(.A(I2), .Z(n_14560));
	notech_inv i_35(.A(I0), .Z(n_14561));
endmodule
module AWMUX_16_32_0(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_1(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_2(I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13,
		 I14, I15, S, O0);

	input [31:0] I0;
	input [31:0] I1;
	input [31:0] I2;
	input [31:0] I3;
	input [31:0] I4;
	input [31:0] I5;
	input [31:0] I6;
	input [31:0] I7;
	input [31:0] I8;
	input [31:0] I9;
	input [31:0] I10;
	input [31:0] I11;
	input [31:0] I12;
	input [31:0] I13;
	input [31:0] I14;
	input [31:0] I15;
	input [3:0] S;
	output [31:0] O0;




	notech_inv i_7660(.A(n_53072), .Z(n_53345));
	notech_inv i_7655(.A(n_53072), .Z(n_53340));
	notech_inv i_7650(.A(n_53061), .Z(n_53334));
	notech_inv i_7645(.A(n_53061), .Z(n_53329));
	notech_inv i_7418(.A(n_53094), .Z(n_53095));
	notech_inv i_7417(.A(n_14553), .Z(n_53094));
	notech_inv i_7415(.A(n_723), .Z(n_53091));
	notech_inv i_7413(.A(n_723), .Z(n_53089));
	notech_inv i_7410(.A(n_723), .Z(n_53086));
	notech_inv i_7408(.A(n_723), .Z(n_53084));
	notech_inv i_7398(.A(n_53072), .Z(n_53073));
	notech_inv i_7397(.A(n_548), .Z(n_53072));
	notech_inv i_7388(.A(n_53061), .Z(n_53062));
	notech_inv i_7387(.A(n_549), .Z(n_53061));
	notech_inv i_180(.A(S[3]), .Z(n_723));
	notech_inv i_179(.A(n_722), .Z(n_684));
	notech_inv i_178(.A(S[2]), .Z(n_722));
	notech_mux4 i_67(.S0(n_548), .S1(n_549), .A(I4[31]), .B(I5[31]), .C(I6[
		31]), .D(I7[31]), .Z(n_615));
	notech_mux4 i_66(.S0(n_548), .S1(n_549), .A(I4[30]), .B(I5[30]), .C(I6[
		30]), .D(I7[30]), .Z(n_614));
	notech_mux4 i_65(.S0(n_548), .S1(n_549), .A(I4[29]), .B(I5[29]), .C(I6[
		29]), .D(I7[29]), .Z(n_613));
	notech_mux4 i_64(.S0(n_548), .S1(n_549), .A(I4[28]), .B(I5[28]), .C(I6[
		28]), .D(I7[28]), .Z(n_612));
	notech_mux4 i_63(.S0(n_548), .S1(n_549), .A(I4[27]), .B(I5[27]), .C(I6[
		27]), .D(I7[27]), .Z(n_611));
	notech_mux4 i_62(.S0(n_548), .S1(n_549), .A(I4[26]), .B(I5[26]), .C(I6[
		26]), .D(I7[26]), .Z(n_610));
	notech_mux4 i_61(.S0(n_548), .S1(n_549), .A(I4[25]), .B(I5[25]), .C(I6[
		25]), .D(I7[25]), .Z(n_609));
	notech_mux4 i_60(.S0(n_548), .S1(n_549), .A(I4[24]), .B(I5[24]), .C(I6[
		24]), .D(I7[24]), .Z(n_608));
	notech_mux4 i_59(.S0(n_548), .S1(n_549), .A(I4[23]), .B(I5[23]), .C(I6[
		23]), .D(I7[23]), .Z(n_607));
	notech_mux4 i_58(.S0(n_548), .S1(n_549), .A(I4[22]), .B(I5[22]), .C(I6[
		22]), .D(I7[22]), .Z(n_606));
	notech_mux4 i_57(.S0(n_548), .S1(n_549), .A(I4[21]), .B(I5[21]), .C(I6[
		21]), .D(I7[21]), .Z(n_605));
	notech_mux4 i_56(.S0(n_548), .S1(n_549), .A(I4[20]), .B(I5[20]), .C(I6[
		20]), .D(I7[20]), .Z(n_604));
	notech_mux4 i_55(.S0(n_548), .S1(n_549), .A(I4[19]), .B(I5[19]), .C(I6[
		19]), .D(I7[19]), .Z(n_603));
	notech_mux4 i_54(.S0(n_548), .S1(n_549), .A(I4[18]), .B(I5[18]), .C(I6[
		18]), .D(I7[18]), .Z(n_602));
	notech_mux4 i_53(.S0(n_548), .S1(n_549), .A(I4[17]), .B(I5[17]), .C(I6[
		17]), .D(I7[17]), .Z(n_601));
	notech_mux4 i_52(.S0(n_548), .S1(n_549), .A(I4[16]), .B(I5[16]), .C(I6[
		16]), .D(I7[16]), .Z(n_600));
	notech_mux4 i_51(.S0(n_53073), .S1(n_53062), .A(I4[15]), .B(I5[15]), .C(I6
		[15]), .D(I7[15]), .Z(n_599));
	notech_mux4 i_50(.S0(n_53073), .S1(n_53062), .A(I4[14]), .B(I5[14]), .C(I6
		[14]), .D(I7[14]), .Z(n_598));
	notech_mux4 i_49(.S0(n_53073), .S1(n_53062), .A(I4[13]), .B(I5[13]), .C(I6
		[13]), .D(I7[13]), .Z(n_597));
	notech_mux4 i_48(.S0(n_53073), .S1(n_53062), .A(I4[12]), .B(I5[12]), .C(I6
		[12]), .D(I7[12]), .Z(n_596));
	notech_mux4 i_47(.S0(n_53073), .S1(n_53062), .A(I4[11]), .B(I5[11]), .C(I6
		[11]), .D(I7[11]), .Z(n_595));
	notech_mux4 i_46(.S0(n_53073), .S1(n_53062), .A(I4[10]), .B(I5[10]), .C(I6
		[10]), .D(I7[10]), .Z(n_594));
	notech_mux4 i_45(.S0(n_53073), .S1(n_53062), .A(I4[9]), .B(I5[9]), .C(I6
		[9]), .D(I7[9]), .Z(n_593));
	notech_mux4 i_44(.S0(n_53073), .S1(n_53062), .A(I4[8]), .B(I5[8]), .C(I6
		[8]), .D(I7[8]), .Z(n_592));
	notech_mux4 i_43(.S0(n_53073), .S1(n_53062), .A(I4[7]), .B(I5[7]), .C(I6
		[7]), .D(I7[7]), .Z(n_591));
	notech_mux4 i_42(.S0(n_53073), .S1(n_53062), .A(I4[6]), .B(I5[6]), .C(I6
		[6]), .D(I7[6]), .Z(n_590));
	notech_mux4 i_41(.S0(n_53073), .S1(n_53062), .A(I4[5]), .B(I5[5]), .C(I6
		[5]), .D(I7[5]), .Z(n_589));
	notech_mux4 i_40(.S0(n_53073), .S1(n_53062), .A(I4[4]), .B(I5[4]), .C(I6
		[4]), .D(I7[4]), .Z(n_588));
	notech_mux4 i_39(.S0(n_53073), .S1(n_53062), .A(I4[3]), .B(I5[3]), .C(I6
		[3]), .D(I7[3]), .Z(n_587));
	notech_mux4 i_38(.S0(n_53073), .S1(n_53062), .A(I4[2]), .B(I5[2]), .C(I6
		[2]), .D(I7[2]), .Z(n_586));
	notech_mux4 i_37(.S0(n_53073), .S1(n_53062), .A(I4[1]), .B(I5[1]), .C(I6
		[1]), .D(I7[1]), .Z(n_585));
	notech_mux4 i_36(.S0(n_53073), .S1(n_53062), .A(I4[0]), .B(I5[0]), .C(I6
		[0]), .D(I7[0]), .Z(n_584));
	notech_mux4 i_33(.S0(n_53340), .S1(n_53329), .A(I0[31]), .B(I1[31]), .C(I2
		[31]), .D(I3[31]), .Z(n_581));
	notech_mux4 i_32(.S0(n_53340), .S1(n_53329), .A(I0[30]), .B(I1[30]), .C(I2
		[30]), .D(I3[30]), .Z(n_580));
	notech_mux4 i_31(.S0(n_53340), .S1(n_53329), .A(I0[29]), .B(I1[29]), .C(I2
		[29]), .D(I3[29]), .Z(n_579));
	notech_mux4 i_30(.S0(n_53340), .S1(n_53329), .A(I0[28]), .B(I1[28]), .C(I2
		[28]), .D(I3[28]), .Z(n_578));
	notech_mux4 i_29(.S0(n_53340), .S1(n_53329), .A(I0[27]), .B(I1[27]), .C(I2
		[27]), .D(I3[27]), .Z(n_577));
	notech_mux4 i_28(.S0(n_53340), .S1(n_53329), .A(I0[26]), .B(I1[26]), .C(I2
		[26]), .D(I3[26]), .Z(n_576));
	notech_mux4 i_27(.S0(n_53340), .S1(n_53329), .A(I0[25]), .B(I1[25]), .C(I2
		[25]), .D(I3[25]), .Z(n_575));
	notech_mux4 i_26(.S0(n_53340), .S1(n_53329), .A(I0[24]), .B(I1[24]), .C(I2
		[24]), .D(I3[24]), .Z(n_574));
	notech_mux4 i_25(.S0(n_53340), .S1(n_53329), .A(I0[23]), .B(I1[23]), .C(I2
		[23]), .D(I3[23]), .Z(n_573));
	notech_mux4 i_24(.S0(n_53340), .S1(n_53329), .A(I0[22]), .B(I1[22]), .C(I2
		[22]), .D(I3[22]), .Z(n_572));
	notech_mux4 i_23(.S0(n_53340), .S1(n_53329), .A(I0[21]), .B(I1[21]), .C(I2
		[21]), .D(I3[21]), .Z(n_571));
	notech_mux4 i_22(.S0(n_53340), .S1(n_53329), .A(I0[20]), .B(I1[20]), .C(I2
		[20]), .D(I3[20]), .Z(n_570));
	notech_mux4 i_21(.S0(n_53340), .S1(n_53329), .A(I0[19]), .B(I1[19]), .C(I2
		[19]), .D(I3[19]), .Z(n_569));
	notech_mux4 i_20(.S0(n_53340), .S1(n_53329), .A(I0[18]), .B(I1[18]), .C(I2
		[18]), .D(I3[18]), .Z(n_568));
	notech_mux4 i_19(.S0(n_53340), .S1(n_53329), .A(I0[17]), .B(I1[17]), .C(I2
		[17]), .D(I3[17]), .Z(n_567));
	notech_mux4 i_18(.S0(n_53340), .S1(n_53329), .A(I0[16]), .B(I1[16]), .C(I2
		[16]), .D(I3[16]), .Z(n_566));
	notech_mux4 i_17(.S0(n_53345), .S1(n_53334), .A(I0[15]), .B(I1[15]), .C(I2
		[15]), .D(I3[15]), .Z(n_565));
	notech_mux4 i_16(.S0(n_53345), .S1(n_53334), .A(I0[14]), .B(I1[14]), .C(I2
		[14]), .D(I3[14]), .Z(n_564));
	notech_mux4 i_15(.S0(n_53345), .S1(n_53334), .A(I0[13]), .B(I1[13]), .C(I2
		[13]), .D(I3[13]), .Z(n_563));
	notech_mux4 i_14(.S0(n_53345), .S1(n_53334), .A(I0[12]), .B(I1[12]), .C(I2
		[12]), .D(I3[12]), .Z(n_562));
	notech_mux4 i_13(.S0(n_53345), .S1(n_53334), .A(I0[11]), .B(I1[11]), .C(I2
		[11]), .D(I3[11]), .Z(n_561));
	notech_mux4 i_12(.S0(n_53345), .S1(n_53334), .A(I0[10]), .B(I1[10]), .C(I2
		[10]), .D(I3[10]), .Z(n_560));
	notech_mux4 i_11(.S0(n_53345), .S1(n_53334), .A(I0[9]), .B(I1[9]), .C(I2
		[9]), .D(I3[9]), .Z(n_559));
	notech_mux4 i_10(.S0(n_53345), .S1(n_53334), .A(I0[8]), .B(I1[8]), .C(I2
		[8]), .D(I3[8]), .Z(n_558));
	notech_mux4 i_9(.S0(n_53345), .S1(n_53334), .A(I0[7]), .B(I1[7]), .C(I2[
		7]), .D(I3[7]), .Z(n_557));
	notech_mux4 i_8(.S0(n_53345), .S1(n_53334), .A(I0[6]), .B(I1[6]), .C(I2[
		6]), .D(I3[6]), .Z(n_556));
	notech_mux4 i_7(.S0(n_53345), .S1(n_53334), .A(I0[5]), .B(I1[5]), .C(I2[
		5]), .D(I3[5]), .Z(n_555));
	notech_mux4 i_6(.S0(n_53345), .S1(n_53334), .A(I0[4]), .B(I1[4]), .C(I2[
		4]), .D(I3[4]), .Z(n_554));
	notech_mux4 i_5(.S0(n_53345), .S1(n_53334), .A(I0[3]), .B(I1[3]), .C(I2[
		3]), .D(I3[3]), .Z(n_553));
	notech_mux4 i_4(.S0(n_53345), .S1(n_53334), .A(I0[2]), .B(I1[2]), .C(I2[
		2]), .D(I3[2]), .Z(n_552));
	notech_mux4 i_3(.S0(n_53345), .S1(n_53334), .A(I0[1]), .B(I1[1]), .C(I2[
		1]), .D(I3[1]), .Z(n_551));
	notech_mux4 i_2(.S0(n_53345), .S1(n_53334), .A(I0[0]), .B(I1[0]), .C(I2[
		0]), .D(I3[0]), .Z(n_550));
	notech_inv i_173(.A(n_719), .Z(n_549));
	notech_inv i_172(.A(S[1]), .Z(n_719));
	notech_inv i_171(.A(n_718), .Z(n_548));
	notech_inv i_170(.A(S[0]), .Z(n_718));
	notech_nand2 i_21804(.A(n_13791), .B(n_13794), .Z(O0[0]));
	notech_nao3 i_21796(.A(n_53094), .B(n_584), .C(n_53086), .Z(n_13794));
	notech_nao3 i_21793(.A(n_550), .B(n_14553), .C(n_53086), .Z(n_13791));
	notech_nand2 i_5094624(.A(n_13815), .B(n_13818), .Z(O0[1]));
	notech_nao3 i_4294625(.A(n_53094), .B(n_585), .C(n_53086), .Z(n_13818)
		);
	notech_nao3 i_3994626(.A(n_551), .B(n_53095), .C(n_53086), .Z(n_13815)
		);
	notech_nand2 i_5094628(.A(n_13839), .B(n_13842), .Z(O0[2]));
	notech_nao3 i_4294629(.A(n_53094), .B(n_586), .C(n_53086), .Z(n_13842)
		);
	notech_nao3 i_3994630(.A(n_552), .B(n_14553), .C(n_53086), .Z(n_13839)
		);
	notech_nand2 i_5094632(.A(n_13863), .B(n_13866), .Z(O0[3]));
	notech_nao3 i_4294633(.A(n_53094), .B(n_587), .C(n_53086), .Z(n_13866)
		);
	notech_nao3 i_3994634(.A(n_553), .B(n_53095), .C(n_53086), .Z(n_13863)
		);
	notech_nand2 i_5094636(.A(n_13887), .B(n_13890), .Z(O0[4]));
	notech_nao3 i_4294637(.A(n_53094), .B(n_588), .C(n_53086), .Z(n_13890)
		);
	notech_nao3 i_3994638(.A(n_554), .B(n_14553), .C(n_53086), .Z(n_13887)
		);
	notech_nand2 i_5094640(.A(n_13911), .B(n_13914), .Z(O0[5]));
	notech_nao3 i_4294641(.A(n_684), .B(n_589), .C(n_53086), .Z(n_13914));
	notech_nao3 i_3994642(.A(n_555), .B(n_53095), .C(n_53086), .Z(n_13911)
		);
	notech_nand2 i_5094644(.A(n_13935), .B(n_13938), .Z(O0[6]));
	notech_nao3 i_4294645(.A(n_53094), .B(n_590), .C(n_53086), .Z(n_13938)
		);
	notech_nao3 i_3994646(.A(n_556), .B(n_14553), .C(n_53086), .Z(n_13935)
		);
	notech_nand2 i_5094648(.A(n_13959), .B(n_13962), .Z(O0[7]));
	notech_nao3 i_4294649(.A(n_53094), .B(n_591), .C(n_53086), .Z(n_13962)
		);
	notech_nao3 i_3994650(.A(n_557), .B(n_53095), .C(n_53086), .Z(n_13959)
		);
	notech_nand2 i_5094652(.A(n_13983), .B(n_13986), .Z(O0[8]));
	notech_nao3 i_4294653(.A(n_53094), .B(n_592), .C(n_53084), .Z(n_13986)
		);
	notech_nao3 i_3994654(.A(n_558), .B(n_14553), .C(n_53084), .Z(n_13983)
		);
	notech_nand2 i_5094656(.A(n_14007), .B(n_14010), .Z(O0[9]));
	notech_nao3 i_4294657(.A(n_53094), .B(n_593), .C(n_53084), .Z(n_14010)
		);
	notech_nao3 i_3994658(.A(n_559), .B(n_53095), .C(n_53084), .Z(n_14007)
		);
	notech_nand2 i_5094660(.A(n_14031), .B(n_14034), .Z(O0[10]));
	notech_nao3 i_4294661(.A(n_53094), .B(n_594), .C(n_53084), .Z(n_14034)
		);
	notech_nao3 i_3994662(.A(n_560), .B(n_14553), .C(n_53084), .Z(n_14031)
		);
	notech_nand2 i_5094664(.A(n_14055), .B(n_14058), .Z(O0[11]));
	notech_nao3 i_4294665(.A(n_53094), .B(n_595), .C(n_53084), .Z(n_14058)
		);
	notech_nao3 i_3994666(.A(n_561), .B(n_53095), .C(n_53084), .Z(n_14055)
		);
	notech_nand2 i_5094668(.A(n_14079), .B(n_14082), .Z(O0[12]));
	notech_nao3 i_4294669(.A(n_53094), .B(n_596), .C(n_53084), .Z(n_14082)
		);
	notech_nao3 i_3994670(.A(n_562), .B(n_14553), .C(n_53084), .Z(n_14079)
		);
	notech_nand2 i_5094672(.A(n_14103), .B(n_14106), .Z(O0[13]));
	notech_nao3 i_4294673(.A(n_53094), .B(n_597), .C(n_53084), .Z(n_14106)
		);
	notech_nao3 i_3994674(.A(n_563), .B(n_53095), .C(n_53084), .Z(n_14103)
		);
	notech_nand2 i_5094676(.A(n_14127), .B(n_14130), .Z(O0[14]));
	notech_nao3 i_4294677(.A(n_53094), .B(n_598), .C(n_53084), .Z(n_14130)
		);
	notech_nao3 i_3994678(.A(n_564), .B(n_14553), .C(n_53084), .Z(n_14127)
		);
	notech_nand2 i_5094680(.A(n_14151), .B(n_14154), .Z(O0[15]));
	notech_nao3 i_4294681(.A(n_53094), .B(n_599), .C(n_53084), .Z(n_14154)
		);
	notech_nao3 i_3994682(.A(n_565), .B(n_53095), .C(n_53084), .Z(n_14151)
		);
	notech_nand2 i_5094684(.A(n_14175), .B(n_14178), .Z(O0[16]));
	notech_nao3 i_4294685(.A(n_684), .B(n_600), .C(n_53091), .Z(n_14178));
	notech_nao3 i_3994686(.A(n_566), .B(n_14553), .C(n_53091), .Z(n_14175)
		);
	notech_nand2 i_5094688(.A(n_14199), .B(n_14202), .Z(O0[17]));
	notech_nao3 i_4294689(.A(n_684), .B(n_601), .C(n_53091), .Z(n_14202));
	notech_nao3 i_3994690(.A(n_567), .B(n_53095), .C(n_53091), .Z(n_14199)
		);
	notech_nand2 i_5094692(.A(n_14223), .B(n_14226), .Z(O0[18]));
	notech_nao3 i_4294693(.A(n_684), .B(n_602), .C(n_53091), .Z(n_14226));
	notech_nao3 i_3994694(.A(n_568), .B(n_14553), .C(n_53091), .Z(n_14223)
		);
	notech_nand2 i_5094696(.A(n_14247), .B(n_14250), .Z(O0[19]));
	notech_nao3 i_4294697(.A(n_684), .B(n_603), .C(n_53091), .Z(n_14250));
	notech_nao3 i_3994698(.A(n_569), .B(n_53095), .C(n_53091), .Z(n_14247)
		);
	notech_nand2 i_5094700(.A(n_14271), .B(n_14274), .Z(O0[20]));
	notech_nao3 i_4294701(.A(n_684), .B(n_604), .C(n_53091), .Z(n_14274));
	notech_nao3 i_3994702(.A(n_570), .B(n_14553), .C(n_53091), .Z(n_14271)
		);
	notech_nand2 i_5094704(.A(n_14295), .B(n_14298), .Z(O0[21]));
	notech_nao3 i_4294705(.A(n_684), .B(n_605), .C(n_53091), .Z(n_14298));
	notech_nao3 i_3994706(.A(n_571), .B(n_14553), .C(n_53091), .Z(n_14295)
		);
	notech_nand2 i_5094708(.A(n_14319), .B(n_14322), .Z(O0[22]));
	notech_nao3 i_4294709(.A(n_684), .B(n_606), .C(n_53091), .Z(n_14322));
	notech_nao3 i_3994710(.A(n_572), .B(n_14553), .C(n_53091), .Z(n_14319)
		);
	notech_nand2 i_5094712(.A(n_14343), .B(n_14346), .Z(O0[23]));
	notech_nao3 i_4294713(.A(n_684), .B(n_607), .C(n_53091), .Z(n_14346));
	notech_nao3 i_3994714(.A(n_573), .B(n_53095), .C(n_53091), .Z(n_14343)
		);
	notech_nand2 i_5094716(.A(n_14367), .B(n_14370), .Z(O0[24]));
	notech_nao3 i_4294717(.A(n_684), .B(n_608), .C(n_53089), .Z(n_14370));
	notech_nao3 i_3994718(.A(n_574), .B(n_14553), .C(n_53089), .Z(n_14367)
		);
	notech_nand2 i_5094720(.A(n_14391), .B(n_14394), .Z(O0[25]));
	notech_nao3 i_4294721(.A(n_684), .B(n_609), .C(n_53089), .Z(n_14394));
	notech_nao3 i_3994722(.A(n_575), .B(n_53095), .C(n_53089), .Z(n_14391)
		);
	notech_nand2 i_5094724(.A(n_14415), .B(n_14418), .Z(O0[26]));
	notech_nao3 i_4294725(.A(n_684), .B(n_610), .C(n_53089), .Z(n_14418));
	notech_nao3 i_3994726(.A(n_576), .B(n_14553), .C(n_53089), .Z(n_14415)
		);
	notech_nand2 i_5094728(.A(n_14439), .B(n_14442), .Z(O0[27]));
	notech_nao3 i_4294729(.A(n_684), .B(n_611), .C(n_53089), .Z(n_14442));
	notech_nao3 i_3994730(.A(n_577), .B(n_53095), .C(n_53089), .Z(n_14439)
		);
	notech_nand2 i_5094732(.A(n_14463), .B(n_14466), .Z(O0[28]));
	notech_nao3 i_4294733(.A(n_684), .B(n_612), .C(n_53089), .Z(n_14466));
	notech_nao3 i_3994734(.A(n_578), .B(n_14553), .C(n_53089), .Z(n_14463)
		);
	notech_nand2 i_5094736(.A(n_14487), .B(n_14490), .Z(O0[29]));
	notech_nao3 i_4294737(.A(n_684), .B(n_613), .C(n_53089), .Z(n_14490));
	notech_nao3 i_3994738(.A(n_579), .B(n_53095), .C(n_53089), .Z(n_14487)
		);
	notech_nand2 i_5094740(.A(n_14511), .B(n_14514), .Z(O0[30]));
	notech_nao3 i_4294741(.A(n_684), .B(n_614), .C(n_53089), .Z(n_14514));
	notech_nao3 i_3994742(.A(n_580), .B(n_14553), .C(n_53089), .Z(n_14511)
		);
	notech_inv i_394743(.A(n_684), .Z(n_14553));
	notech_nand2 i_5094744(.A(n_14535), .B(n_14538), .Z(O0[31]));
	notech_nao3 i_4294745(.A(n_684), .B(n_615), .C(n_53089), .Z(n_14538));
	notech_nao3 i_3994746(.A(n_581), .B(n_53095), .C(n_53089), .Z(n_14535)
		);
endmodule
module AWMUX_16_32_3(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_4(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_5(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_6(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module AWMUX_16_32_7(I0 , I1 , I2 , I3 , I4 , I5 , I6 , I7 , I8 , I9 , I10 , I11 , I12 , I13 , I14 , I15 , S , O0);
input  [31:0] I0;
input  [31:0] I1;
input  [31:0] I2;
input  [31:0] I3;
input  [31:0] I4;
input  [31:0] I5;
input  [31:0] I6;
input  [31:0] I7;
input  [31:0] I8;
input  [31:0] I9;
input  [31:0] I10;
input  [31:0] I11;
input  [31:0] I12;
input  [31:0] I13;
input  [31:0] I14;
input  [31:0] I15;
input  [3:0] S;
output  [31:0] O0;
reg [31:0] O0;

always @(I0 or I1 or I2 or I3 or I4 or I5 or I6 or I7 or I8 or I9 or I10 or I11 or I12 or I13 or I14 or I15 or S or O0)
begin
	case(S)
	4'h0 : O0 = I0;
	4'h1 : O0 = I1;
	4'h2 : O0 = I2;
	4'h3 : O0 = I3;
	4'h4 : O0 = I4;
	4'h5 : O0 = I5;
	4'h6 : O0 = I6;
	4'h7 : O0 = I7;
	4'h8 : O0 = I8;
	4'h9 : O0 = I9;
	4'ha : O0 = I10;
	4'hb : O0 = I11;
	4'hc : O0 = I12;
	4'hd : O0 = I13;
	4'he : O0 = I14;
	default : O0 = I15;
	endcase
end
endmodule

module vliw(clk, rstn, instrc, ie, readio_data, io_add, writeio_data, writeio_req
		, readio_req, writeio_ack, readio_ack, read_reqs, read_ack, read_data
		, over_seg, cr3, cr2, icr2, cr1, cr0, write_reqs, write_ack, write_data
		, Daddr, write_sz, read_sz, cs, add_src, from_acu, to_acu, seg_src
		, pg_en, ready_vliw, valid_op, imm, lenpc, pc_out, pc_req, opz, reps
		, adz, flush_tlb, flush_Dtlb, terminate, start_up, pg_fault, ipg_fault
		, wr_fault, pt_fault, repbytecache);

	input clk;
	input rstn;
	input [127:0] instrc;
	output ie;
	input [31:0] readio_data;
	output [31:0] io_add;
	output [31:0] writeio_data;
	output writeio_req;
	output readio_req;
	input writeio_ack;
	input readio_ack;
	output read_reqs;
	input read_ack;
	input [31:0] read_data;
	input [5:0] over_seg;
	output [31:0] cr3;
	input [31:0] cr2;
	input [31:0] icr2;
	output [31:0] cr1;
	output [31:0] cr0;
	output write_reqs;
	input write_ack;
	output [31:0] write_data;
	output [31:0] Daddr;
	output [1:0] write_sz;
	output [1:0] read_sz;
	output [31:0] cs;
	input [31:0] add_src;
	input [7:0] from_acu;
	output [63:0] to_acu;
	input [2:0] seg_src;
	output pg_en;
	output ready_vliw;
	input valid_op;
	input [63:0] imm;
	input [31:0] lenpc;
	output [31:0] pc_out;
	output pc_req;
	input [2:0] opz;
	input [2:0] reps;
	input adz;
	output flush_tlb;
	output flush_Dtlb;
	output terminate;
	input start_up;
	input pg_fault;
	input ipg_fault;
	input wr_fault;
	input pt_fault;
	output repbytecache;

	wire [4:0] fsm;
	wire [31:0] opa;
	wire [31:0] opc;
	wire [31:0] nbus_11326;
	wire [31:0] nbus_11273;
	wire [31:0] opd;
	wire [31:0] gs;
	wire [2:0] mask8b;
	wire [4:0] vliw_pc;
	wire [31:0] sav_epc;
	wire [31:0] sav_esi;
	wire [31:0] sav_ecx;
	wire [31:0] cr2_reg;
	wire [31:0] nbus_14522;
	wire [31:0] temp_sp;
	wire [31:0] temp_ss;
	wire [31:0] errco;
	wire [31:0] Daddrgs;
	wire [31:0] sav_edi;
	wire [1:0] sav_cs;
	wire [4:0] fsmf;
	wire [31:0] sav_esp;
	wire [1:0] pipe_mul;
	wire [31:0] nbus_11348;
	wire [31:0] nbus_11313;
	wire [31:0] nbus_11304;
	wire [31:0] nbus_11279;
	wire [31:0] write_data_33;
	wire [31:0] write_data_32;
	wire [31:0] write_data_31;
	wire [31:0] write_data_30;
	wire [31:0] write_data_29;
	wire [31:0] write_data_28;
	wire [31:0] write_data_27;
	wire [31:0] write_data_26;
	wire [31:0] write_data_25;
	wire [31:0] Daddrs_8;
	wire [31:0] opc_14;
	wire [31:0] opc_10;
	wire [31:0] Daddrs_3;
	wire [31:0] Daddrs_1;
	wire [31:0] regs_4_2;
	wire [31:0] opa_0;
	wire [31:0] resa_arithbox;
	wire [63:0] divr_0;
	wire [16:0] nbus_144;
	wire [32:0] nbus_143;
	wire [16:0] nbus_142;
	wire [32:0] nbus_141;
	wire [16:0] nbus_140;
	wire [32:0] nbus_139;
	wire [16:0] nbus_138;
	wire [32:0] nbus_137;
	wire [8:0] nbus_136;
	wire [16:0] nbus_135;
	wire [32:0] nbus_134;
	wire [63:0] mul64;
	wire [31:0] add_len_pc32;
	wire [31:0] resb_shift4box;
	wire [31:0] resa_shift4box;
	wire [31:0] resb_shiftbox;
	wire [31:0] resa_shiftbox;
	wire [3:0] calc_sz;
	wire [63:0] tsc;
	wire [3:0] all_cnt;
	wire [31:0] regs_14;
	wire [31:0] regs_12;
	wire [31:0] regs_11;
	wire [31:0] regs_10;
	wire [31:0] regs_8;
	wire [31:0] regs_7;
	wire [31:0] regs_6;
	wire [31:0] regs_5;
	wire [31:0] regs_4;
	wire [31:0] regs_3;
	wire [31:0] regs_2;
	wire [31:0] opb;
	wire [63:0] divq;
	wire [63:0] divr;
	wire [31:0] ecx;
	wire [31:0] regs_0;
	wire [31:0] ldtr;
	wire [31:0] gdtr;
	wire [31:0] idtr;
	wire [31:0] desc;



	notech_inv i_16104(.A(n_62436), .Z(n_62437));
	notech_inv i_16103(.A(\opcode[1] ), .Z(n_62436));
	notech_inv i_16100(.A(n_62432), .Z(n_62433));
	notech_inv i_16099(.A(n_62423), .Z(n_62432));
	notech_inv i_16098(.A(n_62430), .Z(n_62431));
	notech_inv i_16097(.A(n_62415), .Z(n_62430));
	notech_inv i_16096(.A(n_62428), .Z(n_62429));
	notech_inv i_16095(.A(n_62411), .Z(n_62428));
	notech_inv i_16094(.A(n_62426), .Z(n_62427));
	notech_inv i_16093(.A(n_62409), .Z(n_62426));
	notech_inv i_16090(.A(n_62422), .Z(n_62423));
	notech_inv i_16089(.A(n_62427), .Z(n_62422));
	notech_inv i_16086(.A(n_62418), .Z(n_62419));
	notech_inv i_16085(.A(n_62403), .Z(n_62418));
	notech_inv i_16084(.A(n_62416), .Z(n_62417));
	notech_inv i_16083(.A(n_62401), .Z(n_62416));
	notech_inv i_16082(.A(n_62414), .Z(n_62415));
	notech_inv i_16081(.A(n_62417), .Z(n_62414));
	notech_inv i_16080(.A(n_62412), .Z(n_62413));
	notech_inv i_16079(.A(n_62399), .Z(n_62412));
	notech_inv i_16078(.A(n_62410), .Z(n_62411));
	notech_inv i_16077(.A(n_62413), .Z(n_62410));
	notech_inv i_16076(.A(n_62408), .Z(n_62409));
	notech_inv i_16075(.A(n_62429), .Z(n_62408));
	notech_inv i_16072(.A(n_62404), .Z(n_62405));
	notech_inv i_16071(.A(opcode_289113), .Z(n_62404));
	notech_inv i_16070(.A(n_62402), .Z(n_62403));
	notech_inv i_16069(.A(n_62405), .Z(n_62402));
	notech_inv i_16068(.A(n_62400), .Z(n_62401));
	notech_inv i_16067(.A(n_62419), .Z(n_62400));
	notech_inv i_16066(.A(n_62398), .Z(n_62399));
	notech_inv i_16065(.A(n_62431), .Z(n_62398));
	notech_inv i_16062(.A(n_62394), .Z(n_62395));
	notech_inv i_16061(.A(\opcode[0] ), .Z(n_62394));
	notech_inv i_16058(.A(n_62390), .Z(n_62391));
	notech_inv i_16057(.A(n_62377), .Z(n_62390));
	notech_inv i_16056(.A(n_62388), .Z(n_62389));
	notech_inv i_16055(.A(n_62365), .Z(n_62388));
	notech_inv i_16054(.A(n_62386), .Z(n_62387));
	notech_inv i_16053(.A(n_62355), .Z(n_62386));
	notech_inv i_16052(.A(n_62384), .Z(n_62385));
	notech_inv i_16051(.A(n_62347), .Z(n_62384));
	notech_inv i_16050(.A(n_62382), .Z(n_62383));
	notech_inv i_16049(.A(n_62341), .Z(n_62382));
	notech_inv i_16048(.A(n_62380), .Z(n_62381));
	notech_inv i_16047(.A(n_62337), .Z(n_62380));
	notech_inv i_16046(.A(n_62378), .Z(n_62379));
	notech_inv i_16045(.A(n_62335), .Z(n_62378));
	notech_inv i_16044(.A(n_62376), .Z(n_62377));
	notech_inv i_16043(.A(n_62379), .Z(n_62376));
	notech_inv i_16040(.A(n_62372), .Z(n_62373));
	notech_inv i_16039(.A(n_62317), .Z(n_62372));
	notech_inv i_16038(.A(n_62370), .Z(n_62371));
	notech_inv i_16037(.A(n_62311), .Z(n_62370));
	notech_inv i_16036(.A(n_62368), .Z(n_62369));
	notech_inv i_16035(.A(n_62307), .Z(n_62368));
	notech_inv i_16034(.A(n_62366), .Z(n_62367));
	notech_inv i_16033(.A(n_62305), .Z(n_62366));
	notech_inv i_16032(.A(n_62364), .Z(n_62365));
	notech_inv i_16031(.A(n_62367), .Z(n_62364));
	notech_inv i_16030(.A(n_62362), .Z(n_62363));
	notech_inv i_16029(.A(n_62297), .Z(n_62362));
	notech_inv i_16028(.A(n_62360), .Z(n_62361));
	notech_inv i_16027(.A(n_62291), .Z(n_62360));
	notech_inv i_16026(.A(n_62358), .Z(n_62359));
	notech_inv i_16025(.A(n_62287), .Z(n_62358));
	notech_inv i_16024(.A(n_62356), .Z(n_62357));
	notech_inv i_16023(.A(n_62285), .Z(n_62356));
	notech_inv i_16022(.A(n_62354), .Z(n_62355));
	notech_inv i_16021(.A(n_62357), .Z(n_62354));
	notech_inv i_16020(.A(n_62352), .Z(n_62353));
	notech_inv i_16019(.A(n_62279), .Z(n_62352));
	notech_inv i_16018(.A(n_62350), .Z(n_62351));
	notech_inv i_16017(.A(n_62275), .Z(n_62350));
	notech_inv i_16016(.A(n_62348), .Z(n_62349));
	notech_inv i_16015(.A(n_62273), .Z(n_62348));
	notech_inv i_16014(.A(n_62346), .Z(n_62347));
	notech_inv i_16013(.A(n_62349), .Z(n_62346));
	notech_inv i_16012(.A(n_62344), .Z(n_62345));
	notech_inv i_16011(.A(n_62269), .Z(n_62344));
	notech_inv i_16010(.A(n_62342), .Z(n_62343));
	notech_inv i_16009(.A(n_62267), .Z(n_62342));
	notech_inv i_16008(.A(n_62340), .Z(n_62341));
	notech_inv i_16007(.A(n_62343), .Z(n_62340));
	notech_inv i_16006(.A(n_62338), .Z(n_62339));
	notech_inv i_16005(.A(n_62265), .Z(n_62338));
	notech_inv i_16004(.A(n_62336), .Z(n_62337));
	notech_inv i_16003(.A(n_62339), .Z(n_62336));
	notech_inv i_16002(.A(n_62334), .Z(n_62335));
	notech_inv i_16001(.A(n_62381), .Z(n_62334));
	notech_inv i_15990(.A(n_62322), .Z(n_62323));
	notech_inv i_15989(.A(n_62239), .Z(n_62322));
	notech_inv i_15988(.A(n_62320), .Z(n_62321));
	notech_inv i_15987(.A(n_62235), .Z(n_62320));
	notech_inv i_15986(.A(n_62318), .Z(n_62319));
	notech_inv i_15985(.A(n_62233), .Z(n_62318));
	notech_inv i_15984(.A(n_62316), .Z(n_62317));
	notech_inv i_15983(.A(n_62319), .Z(n_62316));
	notech_inv i_15982(.A(n_62314), .Z(n_62315));
	notech_inv i_15981(.A(n_62229), .Z(n_62314));
	notech_inv i_15980(.A(n_62312), .Z(n_62313));
	notech_inv i_15979(.A(n_62227), .Z(n_62312));
	notech_inv i_15978(.A(n_62310), .Z(n_62311));
	notech_inv i_15977(.A(n_62313), .Z(n_62310));
	notech_inv i_15976(.A(n_62308), .Z(n_62309));
	notech_inv i_15975(.A(n_62225), .Z(n_62308));
	notech_inv i_15974(.A(n_62306), .Z(n_62307));
	notech_inv i_15973(.A(n_62309), .Z(n_62306));
	notech_inv i_15972(.A(n_62304), .Z(n_62305));
	notech_inv i_15971(.A(n_62369), .Z(n_62304));
	notech_inv i_15970(.A(n_62302), .Z(n_62303));
	notech_inv i_15969(.A(n_62219), .Z(n_62302));
	notech_inv i_15968(.A(n_62300), .Z(n_62301));
	notech_inv i_15967(.A(n_62215), .Z(n_62300));
	notech_inv i_15966(.A(n_62298), .Z(n_62299));
	notech_inv i_15965(.A(n_62213), .Z(n_62298));
	notech_inv i_15964(.A(n_62296), .Z(n_62297));
	notech_inv i_15963(.A(n_62299), .Z(n_62296));
	notech_inv i_15962(.A(n_62294), .Z(n_62295));
	notech_inv i_15961(.A(n_62209), .Z(n_62294));
	notech_inv i_15960(.A(n_62292), .Z(n_62293));
	notech_inv i_15959(.A(n_62207), .Z(n_62292));
	notech_inv i_15958(.A(n_62290), .Z(n_62291));
	notech_inv i_15957(.A(n_62293), .Z(n_62290));
	notech_inv i_15956(.A(n_62288), .Z(n_62289));
	notech_inv i_15955(.A(n_62205), .Z(n_62288));
	notech_inv i_15954(.A(n_62286), .Z(n_62287));
	notech_inv i_15953(.A(n_62289), .Z(n_62286));
	notech_inv i_15952(.A(n_62284), .Z(n_62285));
	notech_inv i_15951(.A(n_62359), .Z(n_62284));
	notech_inv i_15950(.A(n_62282), .Z(n_62283));
	notech_inv i_15949(.A(n_62201), .Z(n_62282));
	notech_inv i_15948(.A(n_62280), .Z(n_62281));
	notech_inv i_15947(.A(n_62199), .Z(n_62280));
	notech_inv i_15946(.A(n_62278), .Z(n_62279));
	notech_inv i_15945(.A(n_62281), .Z(n_62278));
	notech_inv i_15944(.A(n_62276), .Z(n_62277));
	notech_inv i_15943(.A(n_62197), .Z(n_62276));
	notech_inv i_15942(.A(n_62274), .Z(n_62275));
	notech_inv i_15941(.A(n_62277), .Z(n_62274));
	notech_inv i_15940(.A(n_62272), .Z(n_62273));
	notech_inv i_15939(.A(n_62351), .Z(n_62272));
	notech_inv i_15938(.A(n_62270), .Z(n_62271));
	notech_inv i_15937(.A(n_62195), .Z(n_62270));
	notech_inv i_15936(.A(n_62268), .Z(n_62269));
	notech_inv i_15935(.A(n_62271), .Z(n_62268));
	notech_inv i_15934(.A(n_62266), .Z(n_62267));
	notech_inv i_15933(.A(n_62345), .Z(n_62266));
	notech_inv i_15932(.A(n_62264), .Z(n_62265));
	notech_inv i_15931(.A(n_62383), .Z(n_62264));
	notech_inv i_15930(.A(n_62262), .Z(n_62263));
	notech_inv i_15929(.A(n_62189), .Z(n_62262));
	notech_inv i_15910(.A(n_62242), .Z(n_62243));
	notech_inv i_15909(.A(n_62171), .Z(n_62242));
	notech_inv i_15908(.A(n_62240), .Z(n_62241));
	notech_inv i_15907(.A(n_62169), .Z(n_62240));
	notech_inv i_15906(.A(n_62238), .Z(n_62239));
	notech_inv i_15905(.A(n_62241), .Z(n_62238));
	notech_inv i_15904(.A(n_62236), .Z(n_62237));
	notech_inv i_15903(.A(n_62167), .Z(n_62236));
	notech_inv i_15902(.A(n_62234), .Z(n_62235));
	notech_inv i_15901(.A(n_62237), .Z(n_62234));
	notech_inv i_15900(.A(n_62232), .Z(n_62233));
	notech_inv i_15899(.A(n_62321), .Z(n_62232));
	notech_inv i_15898(.A(n_62230), .Z(n_62231));
	notech_inv i_15897(.A(n_62165), .Z(n_62230));
	notech_inv i_15896(.A(n_62228), .Z(n_62229));
	notech_inv i_15895(.A(n_62231), .Z(n_62228));
	notech_inv i_15894(.A(n_62226), .Z(n_62227));
	notech_inv i_15893(.A(n_62315), .Z(n_62226));
	notech_inv i_15892(.A(n_62224), .Z(n_62225));
	notech_inv i_15891(.A(n_62371), .Z(n_62224));
	notech_inv i_15890(.A(n_62222), .Z(n_62223));
	notech_inv i_15889(.A(n_62161), .Z(n_62222));
	notech_inv i_15888(.A(n_62220), .Z(n_62221));
	notech_inv i_15887(.A(n_62159), .Z(n_62220));
	notech_inv i_15886(.A(n_62218), .Z(n_62219));
	notech_inv i_15885(.A(n_62221), .Z(n_62218));
	notech_inv i_15884(.A(n_62216), .Z(n_62217));
	notech_inv i_15883(.A(n_62157), .Z(n_62216));
	notech_inv i_15882(.A(n_62214), .Z(n_62215));
	notech_inv i_15881(.A(n_62217), .Z(n_62214));
	notech_inv i_15880(.A(n_62212), .Z(n_62213));
	notech_inv i_15879(.A(n_62301), .Z(n_62212));
	notech_inv i_15878(.A(n_62210), .Z(n_62211));
	notech_inv i_15877(.A(n_62155), .Z(n_62210));
	notech_inv i_15876(.A(n_62208), .Z(n_62209));
	notech_inv i_15875(.A(n_62211), .Z(n_62208));
	notech_inv i_15874(.A(n_62206), .Z(n_62207));
	notech_inv i_15873(.A(n_62295), .Z(n_62206));
	notech_inv i_15872(.A(n_62204), .Z(n_62205));
	notech_inv i_15871(.A(n_62361), .Z(n_62204));
	notech_inv i_15870(.A(n_62202), .Z(n_62203));
	notech_inv i_15869(.A(n_62153), .Z(n_62202));
	notech_inv i_15868(.A(n_62200), .Z(n_62201));
	notech_inv i_15867(.A(n_62203), .Z(n_62200));
	notech_inv i_15866(.A(n_62198), .Z(n_62199));
	notech_inv i_15865(.A(n_62283), .Z(n_62198));
	notech_inv i_15864(.A(n_62196), .Z(n_62197));
	notech_inv i_15863(.A(n_62353), .Z(n_62196));
	notech_inv i_15862(.A(n_62194), .Z(n_62195));
	notech_inv i_15861(.A(n_62385), .Z(n_62194));
	notech_inv i_15860(.A(n_62192), .Z(n_62193));
	notech_inv i_15859(.A(n_62147), .Z(n_62192));
	notech_inv i_15858(.A(n_62190), .Z(n_62191));
	notech_inv i_15857(.A(n_62119), .Z(n_62190));
	notech_inv i_15856(.A(n_62188), .Z(n_62189));
	notech_inv i_15855(.A(n_62191), .Z(n_62188));
	notech_inv i_15840(.A(n_62172), .Z(n_62173));
	notech_inv i_15839(.A(n_62077), .Z(n_62172));
	notech_inv i_15838(.A(n_62170), .Z(n_62171));
	notech_inv i_15837(.A(n_62173), .Z(n_62170));
	notech_inv i_15836(.A(n_62168), .Z(n_62169));
	notech_inv i_15835(.A(n_62243), .Z(n_62168));
	notech_inv i_15834(.A(n_62166), .Z(n_62167));
	notech_inv i_15833(.A(n_62323), .Z(n_62166));
	notech_inv i_15832(.A(n_62164), .Z(n_62165));
	notech_inv i_15831(.A(n_62373), .Z(n_62164));
	notech_inv i_15830(.A(n_62162), .Z(n_62163));
	notech_inv i_15829(.A(n_62061), .Z(n_62162));
	notech_inv i_15828(.A(n_62160), .Z(n_62161));
	notech_inv i_15827(.A(n_62163), .Z(n_62160));
	notech_inv i_15826(.A(n_62158), .Z(n_62159));
	notech_inv i_15825(.A(n_62223), .Z(n_62158));
	notech_inv i_15824(.A(n_62156), .Z(n_62157));
	notech_inv i_15823(.A(n_62303), .Z(n_62156));
	notech_inv i_15822(.A(n_62154), .Z(n_62155));
	notech_inv i_15821(.A(n_62363), .Z(n_62154));
	notech_inv i_15820(.A(n_62152), .Z(n_62153));
	notech_inv i_15819(.A(n_62387), .Z(n_62152));
	notech_inv i_15814(.A(n_62146), .Z(n_62147));
	notech_inv i_15813(.A(clk), .Z(n_62146));
	notech_inv i_15785(.A(n_62118), .Z(n_62119));
	notech_inv i_15784(.A(n_62193), .Z(n_62118));
	notech_inv i_15742(.A(n_62076), .Z(n_62077));
	notech_inv i_15741(.A(n_62263), .Z(n_62076));
	notech_inv i_15726(.A(n_62060), .Z(n_62061));
	notech_inv i_15725(.A(n_62389), .Z(n_62060));
	notech_inv i_14572(.A(n_61082), .Z(n_61216));
	notech_inv i_14571(.A(n_61082), .Z(n_61215));
	notech_inv i_14570(.A(n_61082), .Z(n_61214));
	notech_inv i_14569(.A(n_61082), .Z(n_61213));
	notech_inv i_14567(.A(n_61082), .Z(n_61211));
	notech_inv i_14566(.A(n_61082), .Z(n_61210));
	notech_inv i_14565(.A(n_61082), .Z(n_61209));
	notech_inv i_14564(.A(n_61082), .Z(n_61208));
	notech_inv i_14561(.A(n_61082), .Z(n_61205));
	notech_inv i_14560(.A(n_61082), .Z(n_61204));
	notech_inv i_14559(.A(n_61082), .Z(n_61203));
	notech_inv i_14558(.A(n_61082), .Z(n_61202));
	notech_inv i_14556(.A(n_61082), .Z(n_61200));
	notech_inv i_14555(.A(n_61082), .Z(n_61199));
	notech_inv i_14554(.A(n_61082), .Z(n_61198));
	notech_inv i_14553(.A(n_61082), .Z(n_61197));
	notech_inv i_14550(.A(n_61185), .Z(n_61194));
	notech_inv i_14549(.A(n_61185), .Z(n_61193));
	notech_inv i_14548(.A(n_61185), .Z(n_61192));
	notech_inv i_14547(.A(n_61185), .Z(n_61191));
	notech_inv i_14545(.A(n_61185), .Z(n_61189));
	notech_inv i_14544(.A(n_61185), .Z(n_61188));
	notech_inv i_14543(.A(n_61185), .Z(n_61187));
	notech_inv i_14542(.A(n_61185), .Z(n_61186));
	notech_inv i_14541(.A(n_61202), .Z(n_61185));
	notech_inv i_14539(.A(n_61185), .Z(n_61183));
	notech_inv i_14538(.A(n_61185), .Z(n_61182));
	notech_inv i_14537(.A(n_61185), .Z(n_61181));
	notech_inv i_14536(.A(n_61185), .Z(n_61180));
	notech_inv i_14534(.A(n_61185), .Z(n_61178));
	notech_inv i_14533(.A(n_61185), .Z(n_61177));
	notech_inv i_14532(.A(n_61185), .Z(n_61176));
	notech_inv i_14531(.A(n_61185), .Z(n_61175));
	notech_inv i_14527(.A(n_61162), .Z(n_61171));
	notech_inv i_14526(.A(n_61162), .Z(n_61170));
	notech_inv i_14525(.A(n_61162), .Z(n_61169));
	notech_inv i_14524(.A(n_61162), .Z(n_61168));
	notech_inv i_14522(.A(n_61162), .Z(n_61166));
	notech_inv i_14521(.A(n_61162), .Z(n_61165));
	notech_inv i_14520(.A(n_61162), .Z(n_61164));
	notech_inv i_14519(.A(n_61162), .Z(n_61163));
	notech_inv i_14518(.A(n_61208), .Z(n_61162));
	notech_inv i_14516(.A(n_61162), .Z(n_61160));
	notech_inv i_14515(.A(n_61162), .Z(n_61159));
	notech_inv i_14514(.A(n_61162), .Z(n_61158));
	notech_inv i_14513(.A(n_61162), .Z(n_61157));
	notech_inv i_14511(.A(n_61162), .Z(n_61155));
	notech_inv i_14510(.A(n_61162), .Z(n_61154));
	notech_inv i_14509(.A(n_61162), .Z(n_61153));
	notech_inv i_14508(.A(n_61162), .Z(n_61152));
	notech_inv i_14505(.A(n_61140), .Z(n_61149));
	notech_inv i_14504(.A(n_61140), .Z(n_61148));
	notech_inv i_14503(.A(n_61140), .Z(n_61147));
	notech_inv i_14502(.A(n_61140), .Z(n_61146));
	notech_inv i_14500(.A(n_61140), .Z(n_61144));
	notech_inv i_14499(.A(n_61140), .Z(n_61143));
	notech_inv i_14498(.A(n_61140), .Z(n_61142));
	notech_inv i_14497(.A(n_61140), .Z(n_61141));
	notech_inv i_14496(.A(n_61208), .Z(n_61140));
	notech_inv i_14494(.A(n_61140), .Z(n_61138));
	notech_inv i_14493(.A(n_61140), .Z(n_61137));
	notech_inv i_14492(.A(n_61140), .Z(n_61136));
	notech_inv i_14491(.A(n_61140), .Z(n_61135));
	notech_inv i_14489(.A(n_61140), .Z(n_61133));
	notech_inv i_14488(.A(n_61140), .Z(n_61132));
	notech_inv i_14487(.A(n_61140), .Z(n_61131));
	notech_inv i_14486(.A(n_61140), .Z(n_61130));
	notech_inv i_14482(.A(n_61117), .Z(n_61126));
	notech_inv i_14481(.A(n_61117), .Z(n_61125));
	notech_inv i_14480(.A(n_61117), .Z(n_61124));
	notech_inv i_14479(.A(n_61117), .Z(n_61123));
	notech_inv i_14477(.A(n_61117), .Z(n_61121));
	notech_inv i_14476(.A(n_61117), .Z(n_61120));
	notech_inv i_14475(.A(n_61117), .Z(n_61119));
	notech_inv i_14474(.A(n_61117), .Z(n_61118));
	notech_inv i_14473(.A(n_61202), .Z(n_61117));
	notech_inv i_14471(.A(n_61117), .Z(n_61115));
	notech_inv i_14470(.A(n_61117), .Z(n_61114));
	notech_inv i_14469(.A(n_61117), .Z(n_61113));
	notech_inv i_14468(.A(n_61117), .Z(n_61112));
	notech_inv i_14466(.A(n_61117), .Z(n_61110));
	notech_inv i_14465(.A(n_61117), .Z(n_61109));
	notech_inv i_14464(.A(n_61117), .Z(n_61108));
	notech_inv i_14463(.A(n_61117), .Z(n_61107));
	notech_inv i_14460(.A(n_61095), .Z(n_61104));
	notech_inv i_14459(.A(n_61095), .Z(n_61103));
	notech_inv i_14458(.A(n_61095), .Z(n_61102));
	notech_inv i_14457(.A(n_61095), .Z(n_61101));
	notech_inv i_14455(.A(n_61095), .Z(n_61099));
	notech_inv i_14454(.A(n_61095), .Z(n_61098));
	notech_inv i_14453(.A(n_61095), .Z(n_61097));
	notech_inv i_14452(.A(n_61095), .Z(n_61096));
	notech_inv i_14451(.A(n_61202), .Z(n_61095));
	notech_inv i_14449(.A(n_61095), .Z(n_61093));
	notech_inv i_14448(.A(n_61095), .Z(n_61092));
	notech_inv i_14447(.A(n_61095), .Z(n_61091));
	notech_inv i_14446(.A(n_61095), .Z(n_61090));
	notech_inv i_14444(.A(n_61095), .Z(n_61088));
	notech_inv i_14443(.A(n_61095), .Z(n_61087));
	notech_inv i_14442(.A(n_61095), .Z(n_61086));
	notech_inv i_14441(.A(n_61095), .Z(n_61085));
	notech_inv i_14438(.A(rstn), .Z(n_61082));
	notech_inv i_14152(.A(n_60760), .Z(n_60782));
	notech_inv i_14150(.A(n_60760), .Z(n_60780));
	notech_inv i_14149(.A(n_60760), .Z(n_60779));
	notech_inv i_14145(.A(n_60760), .Z(n_60775));
	notech_inv i_14143(.A(n_60760), .Z(n_60773));
	notech_inv i_14140(.A(n_60760), .Z(n_60770));
	notech_inv i_14138(.A(n_60760), .Z(n_60768));
	notech_inv i_14137(.A(n_60760), .Z(n_60767));
	notech_inv i_14132(.A(n_60760), .Z(n_60762));
	notech_inv i_14131(.A(n_60760), .Z(n_60761));
	notech_inv i_14130(.A(n_2580), .Z(n_60760));
	notech_inv i_14123(.A(n_60747), .Z(n_60752));
	notech_inv i_14119(.A(n_60747), .Z(n_60748));
	notech_inv i_14118(.A(fsm[3]), .Z(n_60747));
	notech_inv i_14111(.A(n_60734), .Z(n_60739));
	notech_inv i_14107(.A(n_60734), .Z(n_60735));
	notech_inv i_14106(.A(fsm[0]), .Z(n_60734));
	notech_inv i_14104(.A(n_60718), .Z(n_60731));
	notech_inv i_14102(.A(n_60718), .Z(n_60729));
	notech_inv i_14099(.A(n_60718), .Z(n_60726));
	notech_inv i_14097(.A(n_60718), .Z(n_60724));
	notech_inv i_14094(.A(n_60718), .Z(n_60721));
	notech_inv i_14092(.A(n_60718), .Z(n_60719));
	notech_inv i_14091(.A(n_244256260), .Z(n_60718));
	notech_inv i_13979(.A(n_60601), .Z(n_60602));
	notech_inv i_13978(.A(n_2647), .Z(n_60601));
	notech_inv i_13976(.A(n_60576), .Z(n_60598));
	notech_inv i_13974(.A(n_60576), .Z(n_60596));
	notech_inv i_13973(.A(n_60576), .Z(n_60595));
	notech_inv i_13969(.A(n_60576), .Z(n_60591));
	notech_inv i_13967(.A(n_60576), .Z(n_60589));
	notech_inv i_13964(.A(n_60576), .Z(n_60586));
	notech_inv i_13962(.A(n_60576), .Z(n_60584));
	notech_inv i_13961(.A(n_60576), .Z(n_60583));
	notech_inv i_13957(.A(n_60576), .Z(n_60579));
	notech_inv i_13955(.A(n_60576), .Z(n_60577));
	notech_inv i_13954(.A(pg_fault), .Z(n_60576));
	notech_inv i_13944(.A(n_60557), .Z(n_60563));
	notech_inv i_13939(.A(n_60557), .Z(n_60558));
	notech_inv i_13938(.A(n_28974), .Z(n_60557));
	notech_inv i_13931(.A(n_60548), .Z(n_60549));
	notech_inv i_13930(.A(instrc[123]), .Z(n_60548));
	notech_inv i_13923(.A(n_60535), .Z(n_60540));
	notech_inv i_13919(.A(n_60535), .Z(n_60536));
	notech_inv i_13918(.A(n_28975), .Z(n_60535));
	notech_inv i_13916(.A(n_60524), .Z(n_60532));
	notech_inv i_13914(.A(n_60524), .Z(n_60530));
	notech_inv i_13911(.A(n_60524), .Z(n_60527));
	notech_inv i_13909(.A(n_60524), .Z(n_60525));
	notech_inv i_13908(.A(instrc[122]), .Z(n_60524));
	notech_inv i_13901(.A(n_60515), .Z(n_60516));
	notech_inv i_13900(.A(instrc[121]), .Z(n_60515));
	notech_inv i_13898(.A(n_60502), .Z(n_60512));
	notech_inv i_13897(.A(n_60502), .Z(n_60511));
	notech_inv i_13893(.A(n_60502), .Z(n_60507));
	notech_inv i_13890(.A(n_60502), .Z(n_60504));
	notech_inv i_13889(.A(n_60502), .Z(n_60503));
	notech_inv i_13888(.A(n_28976), .Z(n_60502));
	notech_inv i_13881(.A(n_60489), .Z(n_60494));
	notech_inv i_13877(.A(n_60489), .Z(n_60490));
	notech_inv i_13876(.A(n_2550), .Z(n_60489));
	notech_inv i_13872(.A(n_60478), .Z(n_60484));
	notech_inv i_13867(.A(n_60478), .Z(n_60479));
	notech_inv i_13866(.A(n_165623643), .Z(n_60478));
	notech_inv i_13863(.A(n_60462), .Z(n_60474));
	notech_inv i_13862(.A(n_60462), .Z(n_60473));
	notech_inv i_13857(.A(n_60462), .Z(n_60468));
	notech_inv i_13852(.A(n_60462), .Z(n_60463));
	notech_inv i_13851(.A(n_56066), .Z(n_60462));
	notech_inv i_13842(.A(n_60451), .Z(n_60452));
	notech_inv i_13841(.A(n_301386333), .Z(n_60451));
	notech_inv i_13818(.A(n_60414), .Z(n_60424));
	notech_inv i_13817(.A(n_60414), .Z(n_60423));
	notech_inv i_13813(.A(n_60414), .Z(n_60419));
	notech_inv i_13809(.A(n_60414), .Z(n_60415));
	notech_inv i_13808(.A(ipg_fault), .Z(n_60414));
	notech_inv i_13635(.A(n_60123), .Z(n_60138));
	notech_inv i_13633(.A(n_60123), .Z(n_60136));
	notech_inv i_13626(.A(n_60123), .Z(n_60130));
	notech_inv i_13620(.A(n_60123), .Z(n_60125));
	notech_inv i_13619(.A(n_60123), .Z(cr0[0]));
	notech_inv i_13618(.A(\nbus_14527[0] ), .Z(n_60123));
	notech_inv i_13476(.A(n_59966), .Z(n_59967));
	notech_inv i_13475(.A(n_2572), .Z(n_59966));
	notech_inv i_13467(.A(n_59957), .Z(n_59958));
	notech_inv i_13466(.A(n_272788728), .Z(n_59957));
	notech_inv i_13458(.A(n_59948), .Z(n_59949));
	notech_inv i_13457(.A(n_300186321), .Z(n_59948));
	notech_inv i_13454(.A(n_59873), .Z(n_59945));
	notech_inv i_13453(.A(n_59873), .Z(n_59944));
	notech_inv i_13449(.A(n_59873), .Z(n_59940));
	notech_inv i_13444(.A(n_59873), .Z(n_59936));
	notech_inv i_13443(.A(n_59873), .Z(n_59935));
	notech_inv i_13438(.A(n_59873), .Z(n_59931));
	notech_inv i_13434(.A(n_59873), .Z(n_59927));
	notech_inv i_13433(.A(n_59873), .Z(n_59926));
	notech_inv i_13428(.A(n_59873), .Z(n_59922));
	notech_inv i_13424(.A(n_59873), .Z(n_59918));
	notech_inv i_13422(.A(n_59873), .Z(n_59917));
	notech_inv i_13418(.A(n_59873), .Z(n_59913));
	notech_inv i_13412(.A(n_59873), .Z(n_59908));
	notech_inv i_13411(.A(n_59873), .Z(n_59907));
	notech_inv i_13406(.A(n_59873), .Z(n_59903));
	notech_inv i_13402(.A(n_59893), .Z(n_59899));
	notech_inv i_13401(.A(n_59893), .Z(n_59898));
	notech_inv i_13397(.A(n_59893), .Z(n_59895));
	notech_inv i_13396(.A(n_59893), .Z(n_59894));
	notech_inv i_13395(.A(n_59907), .Z(n_59893));
	notech_inv i_13392(.A(n_59873), .Z(n_59890));
	notech_inv i_13390(.A(n_59873), .Z(n_59889));
	notech_inv i_13386(.A(n_59873), .Z(n_59885));
	notech_inv i_13381(.A(n_59875), .Z(n_59881));
	notech_inv i_13380(.A(n_59875), .Z(n_59880));
	notech_inv i_13376(.A(n_59875), .Z(n_59876));
	notech_inv i_13374(.A(n_59889), .Z(n_59875));
	notech_inv i_13372(.A(n_159623583), .Z(n_59873));
	notech_inv i_13364(.A(n_59864), .Z(n_59865));
	notech_inv i_13363(.A(n_59863), .Z(n_59864));
	notech_inv i_13362(.A(n_59898), .Z(n_59863));
	notech_inv i_13354(.A(n_59855), .Z(n_59856));
	notech_inv i_13353(.A(n_59854), .Z(n_59855));
	notech_inv i_13352(.A(n_59898), .Z(n_59854));
	notech_inv i_13344(.A(n_59846), .Z(n_59847));
	notech_inv i_13342(.A(n_59845), .Z(n_59846));
	notech_inv i_13341(.A(n_59898), .Z(n_59845));
	notech_inv i_13332(.A(n_59836), .Z(n_59837));
	notech_inv i_13331(.A(n_59835), .Z(n_59836));
	notech_inv i_13330(.A(n_59898), .Z(n_59835));
	notech_inv i_13322(.A(n_59827), .Z(n_59828));
	notech_inv i_13321(.A(n_59826), .Z(n_59827));
	notech_inv i_13320(.A(n_59898), .Z(n_59826));
	notech_inv i_13312(.A(n_59818), .Z(n_59819));
	notech_inv i_13310(.A(n_59817), .Z(n_59818));
	notech_inv i_13309(.A(n_59898), .Z(n_59817));
	notech_inv i_13300(.A(n_59808), .Z(n_59809));
	notech_inv i_13299(.A(n_59807), .Z(n_59808));
	notech_inv i_13298(.A(n_59898), .Z(n_59807));
	notech_inv i_13290(.A(n_59799), .Z(n_59800));
	notech_inv i_13289(.A(n_59789), .Z(n_59799));
	notech_inv i_13284(.A(n_59799), .Z(n_59795));
	notech_inv i_13280(.A(n_59799), .Z(n_59791));
	notech_inv i_13277(.A(n_59898), .Z(n_59789));
	notech_inv i_13268(.A(n_59779), .Z(n_59780));
	notech_inv i_13267(.A(n_273688719), .Z(n_59779));
	notech_inv i_13259(.A(n_59770), .Z(n_59771));
	notech_inv i_13258(.A(n_26629), .Z(n_59770));
	notech_inv i_13250(.A(n_59761), .Z(n_59762));
	notech_inv i_13249(.A(n_275288705), .Z(n_59761));
	notech_inv i_13241(.A(n_59752), .Z(n_59753));
	notech_inv i_13240(.A(\nbus_11276[1] ), .Z(n_59752));
	notech_inv i_13232(.A(n_59743), .Z(n_59744));
	notech_inv i_13231(.A(opa[7]), .Z(n_59743));
	notech_inv i_13223(.A(n_59734), .Z(n_59735));
	notech_inv i_13222(.A(opa[6]), .Z(n_59734));
	notech_inv i_13213(.A(n_59725), .Z(n_59726));
	notech_inv i_13212(.A(opa[4]), .Z(n_59725));
	notech_inv i_13204(.A(n_59716), .Z(n_59717));
	notech_inv i_13203(.A(opa[2]), .Z(n_59716));
	notech_inv i_13195(.A(n_59707), .Z(n_59708));
	notech_inv i_13194(.A(opa[1]), .Z(n_59707));
	notech_inv i_13185(.A(n_59698), .Z(n_59699));
	notech_inv i_13184(.A(opa[0]), .Z(n_59698));
	notech_inv i_12884(.A(n_59374), .Z(n_59380));
	notech_inv i_12878(.A(n_59374), .Z(n_59375));
	notech_inv i_12877(.A(n_28969), .Z(n_59374));
	notech_inv i_12874(.A(n_59363), .Z(n_59370));
	notech_inv i_12872(.A(n_59363), .Z(n_59369));
	notech_inv i_12867(.A(n_59363), .Z(n_59364));
	notech_inv i_12866(.A(n_2646), .Z(n_59363));
	notech_inv i_12858(.A(n_59354), .Z(n_59355));
	notech_inv i_12856(.A(n_274988708), .Z(n_59354));
	notech_inv i_12848(.A(n_59345), .Z(n_59346));
	notech_inv i_12847(.A(\nbus_11276[25] ), .Z(n_59345));
	notech_inv i_12839(.A(n_59336), .Z(n_59337));
	notech_inv i_12838(.A(\nbus_11276[26] ), .Z(n_59336));
	notech_inv i_12830(.A(n_59327), .Z(n_59328));
	notech_inv i_12829(.A(\nbus_11276[27] ), .Z(n_59327));
	notech_inv i_12821(.A(n_59318), .Z(n_59319));
	notech_inv i_12820(.A(\nbus_11276[23] ), .Z(n_59318));
	notech_inv i_12812(.A(n_59309), .Z(n_59310));
	notech_inv i_12811(.A(\nbus_11276[21] ), .Z(n_59309));
	notech_inv i_12800(.A(n_59298), .Z(n_59299));
	notech_inv i_12799(.A(instrc[115]), .Z(n_59298));
	notech_inv i_12791(.A(n_59289), .Z(n_59290));
	notech_inv i_12790(.A(instrc[112]), .Z(n_59289));
	notech_inv i_12782(.A(n_59276), .Z(n_59281));
	notech_inv i_12778(.A(n_59276), .Z(n_59277));
	notech_inv i_12776(.A(n_206288851), .Z(n_59276));
	notech_inv i_12774(.A(n_59267), .Z(n_59273));
	notech_inv i_12773(.A(n_59267), .Z(n_59272));
	notech_inv i_12768(.A(n_59267), .Z(n_59268));
	notech_inv i_12767(.A(instrc[114]), .Z(n_59267));
	notech_inv i_12765(.A(n_59258), .Z(n_59264));
	notech_inv i_12764(.A(n_59258), .Z(n_59263));
	notech_inv i_12759(.A(n_59258), .Z(n_59259));
	notech_inv i_12758(.A(instrc[113]), .Z(n_59258));
	notech_inv i_12750(.A(n_59249), .Z(n_59250));
	notech_inv i_12749(.A(n_273588720), .Z(n_59249));
	notech_inv i_12741(.A(n_59240), .Z(n_59241));
	notech_inv i_12740(.A(n_28567), .Z(n_59240));
	notech_inv i_12735(.A(n_60527), .Z(n_59235));
	notech_inv i_12730(.A(n_60527), .Z(n_59230));
	notech_inv i_12724(.A(n_59218), .Z(n_59224));
	notech_inv i_12716(.A(n_59218), .Z(n_59219));
	notech_inv i_12715(.A(n_56189), .Z(n_59218));
	notech_inv i_12707(.A(n_59209), .Z(n_59210));
	notech_inv i_12706(.A(n_272988726), .Z(n_59209));
	notech_inv i_12698(.A(n_59200), .Z(n_59201));
	notech_inv i_12697(.A(n_273188724), .Z(n_59200));
	notech_inv i_12694(.A(n_59171), .Z(n_59197));
	notech_inv i_12692(.A(n_59171), .Z(n_59195));
	notech_inv i_12690(.A(n_59171), .Z(n_59193));
	notech_inv i_12686(.A(n_59171), .Z(n_59190));
	notech_inv i_12684(.A(n_59171), .Z(n_59188));
	notech_inv i_12682(.A(n_59171), .Z(n_59186));
	notech_inv i_12678(.A(n_59171), .Z(n_59183));
	notech_inv i_12676(.A(n_59171), .Z(n_59181));
	notech_inv i_12674(.A(n_59171), .Z(n_59179));
	notech_inv i_12670(.A(n_59171), .Z(n_59176));
	notech_inv i_12668(.A(n_59171), .Z(n_59174));
	notech_inv i_12666(.A(n_59171), .Z(n_59172));
	notech_inv i_12665(.A(n_28984), .Z(n_59171));
	notech_inv i_12662(.A(n_59158), .Z(n_59168));
	notech_inv i_12661(.A(n_59158), .Z(n_59167));
	notech_inv i_12657(.A(n_59158), .Z(n_59163));
	notech_inv i_12652(.A(n_59158), .Z(n_59159));
	notech_inv i_12651(.A(n_123723224), .Z(n_59158));
	notech_inv i_12643(.A(n_59149), .Z(n_59150));
	notech_inv i_12642(.A(n_170914103), .Z(n_59149));
	notech_inv i_12634(.A(n_59140), .Z(n_59141));
	notech_inv i_12633(.A(tcmp), .Z(n_59140));
	notech_inv i_12630(.A(n_59121), .Z(n_59137));
	notech_inv i_12628(.A(n_59121), .Z(n_59135));
	notech_inv i_12627(.A(n_59121), .Z(n_59134));
	notech_inv i_12621(.A(n_59121), .Z(n_59129));
	notech_inv i_12613(.A(n_59121), .Z(n_59122));
	notech_inv i_12612(.A(n_55623), .Z(n_59121));
	notech_inv i_12604(.A(n_59112), .Z(n_59113));
	notech_inv i_12603(.A(opc[0]), .Z(n_59112));
	notech_inv i_12595(.A(n_59103), .Z(n_59104));
	notech_inv i_12594(.A(nbus_11326[29]), .Z(n_59103));
	notech_inv i_12586(.A(n_59094), .Z(n_59095));
	notech_inv i_12585(.A(nbus_11326[31]), .Z(n_59094));
	notech_inv i_12577(.A(n_59085), .Z(n_59086));
	notech_inv i_12576(.A(nbus_11326[24]), .Z(n_59085));
	notech_inv i_12568(.A(n_59076), .Z(n_59077));
	notech_inv i_12566(.A(nbus_11326[28]), .Z(n_59076));
	notech_inv i_12558(.A(n_59067), .Z(n_59068));
	notech_inv i_12557(.A(nbus_11326[26]), .Z(n_59067));
	notech_inv i_12549(.A(n_59058), .Z(n_59059));
	notech_inv i_12548(.A(nbus_11326[27]), .Z(n_59058));
	notech_inv i_12540(.A(n_59049), .Z(n_59050));
	notech_inv i_12539(.A(nbus_11326[30]), .Z(n_59049));
	notech_inv i_12531(.A(n_59040), .Z(n_59041));
	notech_inv i_12530(.A(nbus_11326[23]), .Z(n_59040));
	notech_inv i_12522(.A(n_59031), .Z(n_59032));
	notech_inv i_12521(.A(nbus_11326[22]), .Z(n_59031));
	notech_inv i_12513(.A(n_59022), .Z(n_59023));
	notech_inv i_12512(.A(nbus_11326[25]), .Z(n_59022));
	notech_inv i_12504(.A(n_59013), .Z(n_59014));
	notech_inv i_12502(.A(nbus_11326[19]), .Z(n_59013));
	notech_inv i_12494(.A(n_59004), .Z(n_59005));
	notech_inv i_12493(.A(nbus_11326[20]), .Z(n_59004));
	notech_inv i_12485(.A(n_58995), .Z(n_58996));
	notech_inv i_12484(.A(nbus_11326[21]), .Z(n_58995));
	notech_inv i_12476(.A(n_58986), .Z(n_58987));
	notech_inv i_12475(.A(nbus_11326[16]), .Z(n_58986));
	notech_inv i_12467(.A(n_58977), .Z(n_58978));
	notech_inv i_12466(.A(nbus_11326[17]), .Z(n_58977));
	notech_inv i_12458(.A(n_58968), .Z(n_58969));
	notech_inv i_12457(.A(nbus_11326[18]), .Z(n_58968));
	notech_inv i_12449(.A(n_58959), .Z(n_58960));
	notech_inv i_12448(.A(nbus_11273[0]), .Z(n_58959));
	notech_inv i_12439(.A(n_58950), .Z(n_58951));
	notech_inv i_12437(.A(nbus_11273[31]), .Z(n_58950));
	notech_inv i_12433(.A(n_58939), .Z(n_58945));
	notech_inv i_12427(.A(n_58939), .Z(n_58940));
	notech_inv i_12426(.A(n_273788718), .Z(n_58939));
	notech_inv i_12418(.A(n_58930), .Z(n_58931));
	notech_inv i_12417(.A(n_205588858), .Z(n_58930));
	notech_inv i_12409(.A(n_58921), .Z(n_58922));
	notech_inv i_12408(.A(n_55808), .Z(n_58921));
	notech_inv i_12400(.A(n_58912), .Z(n_58913));
	notech_inv i_12399(.A(n_2831), .Z(n_58912));
	notech_inv i_12391(.A(n_58903), .Z(n_58904));
	notech_inv i_12389(.A(n_2825), .Z(n_58903));
	notech_inv i_12381(.A(n_58894), .Z(n_58895));
	notech_inv i_12380(.A(n_2645), .Z(n_58894));
	notech_inv i_12372(.A(n_58885), .Z(n_58886));
	notech_inv i_12371(.A(n_55838), .Z(n_58885));
	notech_inv i_12150(.A(n_58655), .Z(n_58661));
	notech_inv i_12148(.A(n_58655), .Z(n_58660));
	notech_inv i_12144(.A(n_58655), .Z(n_58656));
	notech_inv i_12143(.A(n_274188716), .Z(n_58655));
	notech_inv i_12132(.A(n_58644), .Z(n_58645));
	notech_inv i_12131(.A(n_26390), .Z(n_58644));
	notech_inv i_12083(.A(n_58590), .Z(n_58591));
	notech_inv i_12082(.A(n_26498), .Z(n_58590));
	notech_inv i_12058(.A(n_27564), .Z(n_58566));
	notech_inv i_12040(.A(n_58547), .Z(n_58548));
	notech_inv i_12039(.A(n_27565), .Z(n_58547));
	notech_inv i_12024(.A(n_58531), .Z(n_58532));
	notech_inv i_12023(.A(n_57461), .Z(n_58531));
	notech_inv i_12015(.A(n_58522), .Z(n_58523));
	notech_inv i_12014(.A(n_358079925), .Z(n_58522));
	notech_inv i_12006(.A(n_58513), .Z(n_58514));
	notech_inv i_12004(.A(n_2193), .Z(n_58513));
	notech_inv i_11996(.A(n_58504), .Z(n_58505));
	notech_inv i_11995(.A(n_55943), .Z(n_58504));
	notech_inv i_11987(.A(n_58495), .Z(n_58496));
	notech_inv i_11986(.A(n_55131), .Z(n_58495));
	notech_inv i_11978(.A(n_58482), .Z(n_58487));
	notech_inv i_11974(.A(n_58482), .Z(n_58483));
	notech_inv i_11972(.A(n_55878), .Z(n_58482));
	notech_inv i_11004(.A(n_57437), .Z(n_57448));
	notech_inv i_10996(.A(n_57437), .Z(n_57438));
	notech_inv i_10995(.A(n_56099), .Z(n_57437));
	notech_inv i_10987(.A(n_57422), .Z(n_57424));
	notech_inv i_10986(.A(n_57413), .Z(n_57422));
	notech_inv i_10978(.A(n_57403), .Z(n_57404));
	notech_inv i_10977(.A(n_1844), .Z(n_57403));
	notech_inv i_10969(.A(n_57381), .Z(n_57383));
	notech_inv i_10968(.A(n_244656264), .Z(n_57381));
	notech_inv i_10966(.A(n_57366), .Z(n_57373));
	notech_inv i_10964(.A(n_57366), .Z(n_57371));
	notech_inv i_10960(.A(n_57366), .Z(n_57367));
	notech_inv i_10959(.A(n_193714331), .Z(n_57366));
	notech_inv i_10951(.A(n_57356), .Z(n_57358));
	notech_inv i_10950(.A(n_197114365), .Z(n_57356));
	notech_inv i_10945(.A(n_57337), .Z(n_57343));
	notech_inv i_10939(.A(n_57337), .Z(n_57338));
	notech_inv i_10938(.A(n_56179), .Z(n_57337));
	notech_inv i_10930(.A(n_57322), .Z(n_57326));
	notech_inv i_10929(.A(nbus_11273[7]), .Z(n_57322));
	notech_inv i_10921(.A(n_57311), .Z(n_57312));
	notech_inv i_10920(.A(n_2786), .Z(n_57311));
	notech_inv i_10910(.A(n_57297), .Z(n_57298));
	notech_inv i_10909(.A(n_2784), .Z(n_57297));
	notech_inv i_10798(.A(n_57176), .Z(n_57177));
	notech_inv i_10797(.A(n_2785), .Z(n_57176));
	notech_inv i_10789(.A(n_57167), .Z(n_57168));
	notech_inv i_10787(.A(n_2803), .Z(n_57167));
	notech_inv i_10783(.A(n_57154), .Z(n_57162));
	notech_inv i_10782(.A(n_57154), .Z(n_57161));
	notech_inv i_10777(.A(n_57154), .Z(n_57157));
	notech_inv i_10776(.A(n_57154), .Z(n_57156));
	notech_inv i_10775(.A(n_57154), .Z(n_57155));
	notech_inv i_10774(.A(instrc[106]), .Z(n_57154));
	notech_inv i_10724(.A(n_56971), .Z(n_56972));
	notech_inv i_10722(.A(n_2806), .Z(n_56971));
	notech_inv i_10714(.A(n_56962), .Z(n_56963));
	notech_inv i_10712(.A(n_2612), .Z(n_56962));
	notech_inv i_10702(.A(n_56951), .Z(n_56952));
	notech_inv i_10701(.A(n_2804), .Z(n_56951));
	notech_inv i_10693(.A(n_56942), .Z(n_56943));
	notech_inv i_10692(.A(\nbus_11276[31] ), .Z(n_56942));
	notech_inv i_10682(.A(n_56931), .Z(n_56932));
	notech_inv i_10680(.A(n_2810), .Z(n_56931));
	notech_inv i_10670(.A(n_56920), .Z(n_56921));
	notech_inv i_10669(.A(n_2808), .Z(n_56920));
	notech_inv i_10659(.A(n_56909), .Z(n_56910));
	notech_inv i_10658(.A(n_2807), .Z(n_56909));
	notech_inv i_10650(.A(n_56900), .Z(n_56901));
	notech_inv i_10648(.A(nbus_11273[30]), .Z(n_56900));
	notech_inv i_10640(.A(n_56891), .Z(n_56892));
	notech_inv i_10639(.A(nbus_11273[29]), .Z(n_56891));
	notech_inv i_10631(.A(n_56882), .Z(n_56883));
	notech_inv i_10630(.A(nbus_11273[28]), .Z(n_56882));
	notech_inv i_10622(.A(n_56873), .Z(n_56874));
	notech_inv i_10621(.A(nbus_11273[27]), .Z(n_56873));
	notech_inv i_10613(.A(n_56864), .Z(n_56865));
	notech_inv i_10612(.A(nbus_11273[26]), .Z(n_56864));
	notech_inv i_10604(.A(n_56855), .Z(n_56856));
	notech_inv i_10603(.A(nbus_11273[25]), .Z(n_56855));
	notech_inv i_10595(.A(n_56846), .Z(n_56847));
	notech_inv i_10594(.A(nbus_11273[24]), .Z(n_56846));
	notech_inv i_10586(.A(n_56837), .Z(n_56838));
	notech_inv i_10584(.A(nbus_11273[23]), .Z(n_56837));
	notech_inv i_10576(.A(n_56828), .Z(n_56829));
	notech_inv i_10575(.A(nbus_11273[22]), .Z(n_56828));
	notech_inv i_10567(.A(n_56819), .Z(n_56820));
	notech_inv i_10566(.A(nbus_11273[21]), .Z(n_56819));
	notech_inv i_10558(.A(n_56810), .Z(n_56811));
	notech_inv i_10557(.A(nbus_11273[20]), .Z(n_56810));
	notech_inv i_10549(.A(n_56801), .Z(n_56802));
	notech_inv i_10548(.A(nbus_11273[19]), .Z(n_56801));
	notech_inv i_10540(.A(n_56792), .Z(n_56793));
	notech_inv i_10539(.A(nbus_11273[18]), .Z(n_56792));
	notech_inv i_10531(.A(n_56783), .Z(n_56784));
	notech_inv i_10530(.A(nbus_11273[17]), .Z(n_56783));
	notech_inv i_10522(.A(n_56774), .Z(n_56775));
	notech_inv i_10520(.A(nbus_11273[16]), .Z(n_56774));
	notech_inv i_10512(.A(n_56765), .Z(n_56766));
	notech_inv i_10511(.A(nbus_11273[15]), .Z(n_56765));
	notech_inv i_10503(.A(n_56756), .Z(n_56757));
	notech_inv i_10502(.A(nbus_11273[14]), .Z(n_56756));
	notech_inv i_10494(.A(n_56747), .Z(n_56748));
	notech_inv i_10493(.A(nbus_11273[13]), .Z(n_56747));
	notech_inv i_10485(.A(n_56738), .Z(n_56739));
	notech_inv i_10484(.A(nbus_11273[12]), .Z(n_56738));
	notech_inv i_10476(.A(n_56729), .Z(n_56730));
	notech_inv i_10475(.A(nbus_11273[11]), .Z(n_56729));
	notech_inv i_10467(.A(n_56720), .Z(n_56721));
	notech_inv i_10466(.A(nbus_11273[10]), .Z(n_56720));
	notech_inv i_10458(.A(n_56711), .Z(n_56712));
	notech_inv i_10456(.A(nbus_11273[9]), .Z(n_56711));
	notech_inv i_10448(.A(n_56702), .Z(n_56703));
	notech_inv i_10447(.A(nbus_11273[8]), .Z(n_56702));
	notech_inv i_10439(.A(n_56693), .Z(n_56694));
	notech_inv i_10438(.A(nbus_11273[6]), .Z(n_56693));
	notech_inv i_10430(.A(n_56684), .Z(n_56685));
	notech_inv i_10429(.A(nbus_11273[5]), .Z(n_56684));
	notech_inv i_10421(.A(n_56675), .Z(n_56676));
	notech_inv i_10420(.A(nbus_11273[4]), .Z(n_56675));
	notech_inv i_10412(.A(n_56666), .Z(n_56667));
	notech_inv i_10411(.A(nbus_11273[3]), .Z(n_56666));
	notech_inv i_10403(.A(n_56657), .Z(n_56658));
	notech_inv i_10402(.A(nbus_11273[2]), .Z(n_56657));
	notech_inv i_10392(.A(n_56648), .Z(n_56649));
	notech_inv i_10390(.A(nbus_11273[1]), .Z(n_56648));
	notech_inv i_10382(.A(n_56639), .Z(n_56640));
	notech_inv i_10381(.A(n_55936), .Z(n_56639));
	notech_inv i_10373(.A(n_56626), .Z(n_56631));
	notech_inv i_10369(.A(n_56626), .Z(n_56627));
	notech_inv i_10368(.A(n_329546800), .Z(n_56626));
	notech_inv i_10360(.A(n_56617), .Z(n_56618));
	notech_inv i_10358(.A(n_55231), .Z(n_56617));
	notech_inv i_10350(.A(n_56608), .Z(n_56609));
	notech_inv i_10349(.A(n_287372184), .Z(n_56608));
	notech_inv i_10326(.A(n_56577), .Z(n_56583));
	notech_inv i_10321(.A(n_56577), .Z(n_56578));
	notech_inv i_10320(.A(n_57292), .Z(n_56577));
	notech_inv i_10317(.A(n_56568), .Z(n_56574));
	notech_inv i_10316(.A(n_56568), .Z(n_56573));
	notech_inv i_10312(.A(n_56568), .Z(n_56569));
	notech_inv i_10310(.A(n_56107), .Z(n_56568));
	notech_inv i_10302(.A(n_56559), .Z(n_56560));
	notech_inv i_10301(.A(n_56112), .Z(n_56559));
	notech_inv i_10293(.A(n_56546), .Z(n_56551));
	notech_inv i_10289(.A(n_56546), .Z(n_56547));
	notech_inv i_10288(.A(n_56104), .Z(n_56546));
	notech_inv i_10280(.A(n_56537), .Z(n_56538));
	notech_inv i_10278(.A(n_54520), .Z(n_56537));
	notech_inv i_10270(.A(n_56528), .Z(n_56529));
	notech_inv i_10269(.A(n_334662244), .Z(n_56528));
	notech_inv i_10261(.A(n_56519), .Z(n_56520));
	notech_inv i_10260(.A(n_341962313), .Z(n_56519));
	notech_inv i_10252(.A(n_56510), .Z(n_56511));
	notech_inv i_10251(.A(n_334762245), .Z(n_56510));
	notech_inv i_10243(.A(n_56497), .Z(n_56502));
	notech_inv i_10238(.A(n_56497), .Z(n_56498));
	notech_inv i_10237(.A(n_2044), .Z(n_56497));
	notech_inv i_10233(.A(n_56486), .Z(n_56492));
	notech_inv i_10227(.A(n_56486), .Z(n_56487));
	notech_inv i_10226(.A(instrc[117]), .Z(n_56486));
	notech_inv i_10218(.A(n_56477), .Z(n_56478));
	notech_inv i_10217(.A(instrc[118]), .Z(n_56477));
	notech_inv i_10209(.A(n_56468), .Z(n_56469));
	notech_inv i_10208(.A(instrc[119]), .Z(n_56468));
	notech_inv i_10205(.A(n_56457), .Z(n_56465));
	notech_inv i_10203(.A(n_56457), .Z(n_56463));
	notech_inv i_10200(.A(n_56457), .Z(n_56460));
	notech_inv i_10197(.A(n_56457), .Z(n_56458));
	notech_inv i_10196(.A(instrc[116]), .Z(n_56457));
	notech_inv i_10188(.A(n_56448), .Z(n_56449));
	notech_inv i_10187(.A(n_1976), .Z(n_56448));
	notech_inv i_10179(.A(n_56439), .Z(n_56440));
	notech_inv i_10178(.A(n_29010), .Z(n_56439));
	notech_inv i_10170(.A(n_56430), .Z(n_56431));
	notech_inv i_10169(.A(n_264436799), .Z(n_56430));
	notech_inv i_10164(.A(n_56419), .Z(n_56425));
	notech_inv i_10158(.A(n_56419), .Z(n_56420));
	notech_inv i_10157(.A(n_342162315), .Z(n_56419));
	notech_inv i_10154(.A(n_56403), .Z(n_56415));
	notech_inv i_10153(.A(n_56403), .Z(n_56414));
	notech_inv i_10147(.A(n_56403), .Z(n_56409));
	notech_inv i_10141(.A(n_56403), .Z(n_56404));
	notech_inv i_10140(.A(n_56180), .Z(n_56403));
	notech_inv i_10132(.A(n_56394), .Z(n_56395));
	notech_inv i_10131(.A(n_56183), .Z(n_56394));
	notech_inv i_10123(.A(n_56381), .Z(n_56386));
	notech_inv i_10118(.A(n_56381), .Z(n_56382));
	notech_inv i_10117(.A(n_54439), .Z(n_56381));
	notech_inv i_10113(.A(n_56362), .Z(n_56376));
	notech_inv i_10112(.A(n_56362), .Z(n_56375));
	notech_inv i_10105(.A(n_56362), .Z(n_56369));
	notech_inv i_10098(.A(n_56362), .Z(n_56363));
	notech_inv i_10097(.A(n_56064), .Z(n_56362));
	notech_inv i_10089(.A(n_56353), .Z(n_56354));
	notech_inv i_10088(.A(n_205088863), .Z(n_56353));
	notech_inv i_10080(.A(n_56344), .Z(n_56345));
	notech_inv i_10078(.A(n_2240), .Z(n_56344));
	notech_inv i_10070(.A(n_56335), .Z(n_56336));
	notech_inv i_10069(.A(n_334862246), .Z(n_56335));
	notech_inv i_10061(.A(n_56326), .Z(n_56327));
	notech_inv i_10060(.A(n_334962247), .Z(n_56326));
	notech_inv i_10050(.A(n_56315), .Z(n_56316));
	notech_inv i_10049(.A(\nbus_11332[0] ), .Z(n_56315));
	notech_inv i_10043(.A(n_56304), .Z(n_56310));
	notech_inv i_10037(.A(n_56304), .Z(n_56305));
	notech_inv i_10036(.A(n_56181), .Z(n_56304));
	notech_inv i_10028(.A(n_56295), .Z(n_56296));
	notech_inv i_10027(.A(n_56182), .Z(n_56295));
	notech_inv i_10023(.A(n_56284), .Z(n_56290));
	notech_inv i_10017(.A(n_56284), .Z(n_56285));
	notech_inv i_10016(.A(n_56185), .Z(n_56284));
	notech_inv i_10008(.A(n_56275), .Z(n_56276));
	notech_inv i_10007(.A(n_56186), .Z(n_56275));
	notech_inv i_10002(.A(n_56264), .Z(n_56270));
	notech_inv i_9996(.A(n_56264), .Z(n_56265));
	notech_inv i_9995(.A(n_56188), .Z(n_56264));
	notech_inv i_9987(.A(n_56254), .Z(n_56255));
	notech_inv i_9986(.A(n_2262), .Z(n_56254));
	notech_inv i_9978(.A(n_56245), .Z(n_56246));
	notech_inv i_9977(.A(n_2261), .Z(n_56245));
	notech_inv i_9972(.A(n_56234), .Z(n_56240));
	notech_inv i_9967(.A(n_56234), .Z(n_56235));
	notech_inv i_9965(.A(n_56175), .Z(n_56234));
	notech_inv i_9957(.A(n_56225), .Z(n_56226));
	notech_inv i_9956(.A(n_56178), .Z(n_56225));
	notech_inv i_9948(.A(n_56215), .Z(n_56216));
	notech_inv i_9947(.A(n_56057), .Z(n_56215));
	notech_inv i_9939(.A(n_56206), .Z(n_56207));
	notech_inv i_9938(.A(\nbus_11276[24] ), .Z(n_56206));
	notech_inv i_9936(.A(n_56195), .Z(n_56203));
	notech_inv i_9933(.A(n_56195), .Z(n_56201));
	notech_inv i_9929(.A(n_56195), .Z(n_56197));
	notech_inv i_9928(.A(n_56195), .Z(n_56196));
	notech_inv i_9927(.A(n_2197), .Z(n_56195));
	notech_inv i_9918(.A(n_56171), .Z(n_56177));
	notech_inv i_9913(.A(n_56171), .Z(n_56172));
	notech_inv i_9912(.A(n_204788866), .Z(n_56171));
	notech_inv i_9904(.A(n_56157), .Z(n_56163));
	notech_inv i_9899(.A(n_56157), .Z(n_56158));
	notech_inv i_9898(.A(n_274288715), .Z(n_56157));
	notech_inv i_9894(.A(n_56138), .Z(n_56151));
	notech_inv i_9888(.A(n_56138), .Z(n_56144));
	notech_inv i_9882(.A(n_56138), .Z(n_56139));
	notech_inv i_9881(.A(n_54446), .Z(n_56138));
	notech_inv i_9873(.A(n_56125), .Z(n_56130));
	notech_inv i_9868(.A(n_56125), .Z(n_56126));
	notech_inv i_9867(.A(n_54451), .Z(n_56125));
	notech_inv i_9864(.A(n_56106), .Z(n_56121));
	notech_inv i_9863(.A(n_56106), .Z(n_56120));
	notech_inv i_9857(.A(n_56106), .Z(n_56114));
	notech_inv i_9851(.A(n_56106), .Z(n_56108));
	notech_inv i_9850(.A(n_2189), .Z(n_56106));
	notech_inv i_9846(.A(n_56091), .Z(n_56097));
	notech_inv i_9840(.A(n_56091), .Z(n_56092));
	notech_inv i_9839(.A(n_54465), .Z(n_56091));
	notech_inv i_9834(.A(n_56073), .Z(n_56086));
	notech_inv i_9828(.A(n_56073), .Z(n_56081));
	notech_inv i_9823(.A(n_56073), .Z(n_56074));
	notech_inv i_9822(.A(n_274388714), .Z(n_56073));
	notech_inv i_9817(.A(n_56042), .Z(n_56068));
	notech_inv i_9811(.A(n_56042), .Z(n_56049));
	notech_inv i_9806(.A(n_56042), .Z(n_56043));
	notech_inv i_9804(.A(n_55868), .Z(n_56042));
	notech_inv i_9801(.A(n_56021), .Z(n_56035));
	notech_inv i_9800(.A(n_56021), .Z(n_56033));
	notech_inv i_9794(.A(n_56021), .Z(n_56023));
	notech_inv i_9793(.A(n_55869), .Z(n_56021));
	notech_inv i_9785(.A(n_56008), .Z(n_56013));
	notech_inv i_9780(.A(n_56008), .Z(n_56009));
	notech_inv i_9779(.A(n_55870), .Z(n_56008));
	notech_inv i_9775(.A(n_55991), .Z(n_55998));
	notech_inv i_9769(.A(n_55991), .Z(n_55992));
	notech_inv i_9768(.A(n_55871), .Z(n_55991));
	notech_inv i_9760(.A(n_55964), .Z(n_55972));
	notech_inv i_9755(.A(n_55964), .Z(n_55965));
	notech_inv i_9754(.A(n_55872), .Z(n_55964));
	notech_inv i_9746(.A(n_55946), .Z(n_55952));
	notech_inv i_9742(.A(n_55946), .Z(n_55947));
	notech_inv i_9740(.A(n_55873), .Z(n_55946));
	notech_inv i_9736(.A(n_55932), .Z(n_55940));
	notech_inv i_9730(.A(n_55932), .Z(n_55934));
	notech_inv i_9729(.A(n_2242), .Z(n_55932));
	notech_inv i_9721(.A(n_55918), .Z(n_55924));
	notech_inv i_9716(.A(n_55918), .Z(n_55919));
	notech_inv i_9715(.A(n_54535), .Z(n_55918));
	notech_inv i_9707(.A(n_55905), .Z(n_55910));
	notech_inv i_9703(.A(n_55905), .Z(n_55906));
	notech_inv i_9702(.A(n_55864), .Z(n_55905));
	notech_inv i_9697(.A(n_55887), .Z(n_55898));
	notech_inv i_9691(.A(n_55887), .Z(n_55893));
	notech_inv i_9686(.A(n_55887), .Z(n_55888));
	notech_inv i_9684(.A(n_55865), .Z(n_55887));
	notech_inv i_9676(.A(n_55863), .Z(n_55879));
	notech_inv i_9672(.A(n_55863), .Z(n_55866));
	notech_inv i_9671(.A(n_55867), .Z(n_55863));
	notech_inv i_9667(.A(n_55851), .Z(n_55859));
	notech_inv i_9666(.A(n_55851), .Z(n_55858));
	notech_inv i_9660(.A(n_55851), .Z(n_55852));
	notech_inv i_9659(.A(n_56062), .Z(n_55851));
	notech_inv i_9655(.A(n_55818), .Z(n_55837));
	notech_inv i_9649(.A(n_55818), .Z(n_55827));
	notech_inv i_9643(.A(n_55818), .Z(n_55820));
	notech_inv i_9642(.A(n_56065), .Z(n_55818));
	notech_inv i_9634(.A(n_55806), .Z(n_55807));
	notech_inv i_9633(.A(n_56063), .Z(n_55806));
	notech_inv i_9625(.A(n_55785), .Z(n_55798));
	notech_inv i_9620(.A(n_55785), .Z(n_55794));
	notech_inv i_9619(.A(n_54367), .Z(n_55785));
	notech_inv i_9511(.A(n_55666), .Z(n_55667));
	notech_inv i_9510(.A(n_56061), .Z(n_55666));
	notech_inv i_9502(.A(n_55655), .Z(n_55658));
	notech_inv i_9501(.A(n_56060), .Z(n_55655));
	notech_inv i_9493(.A(n_55646), .Z(n_55647));
	notech_inv i_9492(.A(\nbus_11276[22] ), .Z(n_55646));
	notech_inv i_9484(.A(n_55630), .Z(n_55631));
	notech_inv i_9482(.A(\nbus_11276[20] ), .Z(n_55630));
	notech_inv i_9474(.A(n_55618), .Z(n_55620));
	notech_inv i_9473(.A(\nbus_11276[19] ), .Z(n_55618));
	notech_inv i_9465(.A(n_55608), .Z(n_55609));
	notech_inv i_9464(.A(\nbus_11276[18] ), .Z(n_55608));
	notech_inv i_9456(.A(n_55599), .Z(n_55600));
	notech_inv i_9455(.A(\nbus_11276[17] ), .Z(n_55599));
	notech_inv i_9447(.A(n_55589), .Z(n_55590));
	notech_inv i_9446(.A(\nbus_11276[16] ), .Z(n_55589));
	notech_inv i_9438(.A(n_55577), .Z(n_55578));
	notech_inv i_9437(.A(\nbus_11276[15] ), .Z(n_55577));
	notech_inv i_9429(.A(n_55565), .Z(n_55566));
	notech_inv i_9428(.A(\nbus_11276[14] ), .Z(n_55565));
	notech_inv i_9420(.A(n_55551), .Z(n_55552));
	notech_inv i_9418(.A(\nbus_11276[13] ), .Z(n_55551));
	notech_inv i_9410(.A(n_55540), .Z(n_55542));
	notech_inv i_9409(.A(\nbus_11276[12] ), .Z(n_55540));
	notech_inv i_9401(.A(n_55521), .Z(n_55522));
	notech_inv i_9400(.A(n_2145), .Z(n_55521));
	notech_inv i_9390(.A(n_55507), .Z(n_55508));
	notech_inv i_9389(.A(n_26808), .Z(n_55507));
	notech_inv i_9378(.A(n_55491), .Z(n_55492));
	notech_inv i_9377(.A(n_2345), .Z(n_55491));
	notech_inv i_9373(.A(n_55477), .Z(n_55484));
	notech_inv i_9367(.A(n_55477), .Z(n_55478));
	notech_inv i_9366(.A(n_187871189), .Z(n_55477));
	notech_inv i_9358(.A(n_55468), .Z(n_55469));
	notech_inv i_9357(.A(\nbus_11276[11] ), .Z(n_55468));
	notech_inv i_9349(.A(n_55458), .Z(n_55460));
	notech_inv i_9348(.A(\eflags[10] ), .Z(n_55458));
	notech_inv i_9340(.A(n_55449), .Z(n_55450));
	notech_inv i_9338(.A(n_29091), .Z(n_55449));
	notech_inv i_9330(.A(n_55437), .Z(n_55438));
	notech_inv i_9329(.A(\nbus_11276[10] ), .Z(n_55437));
	notech_inv i_9321(.A(n_55423), .Z(n_55425));
	notech_inv i_9320(.A(\nbus_11276[9] ), .Z(n_55423));
	notech_inv i_9312(.A(n_55412), .Z(n_55413));
	notech_inv i_9311(.A(\nbus_11276[8] ), .Z(n_55412));
	notech_inv i_9302(.A(n_55399), .Z(n_55400));
	notech_inv i_9301(.A(\nbus_11276[7] ), .Z(n_55399));
	notech_inv i_9293(.A(n_55386), .Z(n_55387));
	notech_inv i_9292(.A(\nbus_11276[6] ), .Z(n_55386));
	notech_inv i_9284(.A(n_55374), .Z(n_55375));
	notech_inv i_9283(.A(\nbus_11276[5] ), .Z(n_55374));
	notech_inv i_9274(.A(n_55364), .Z(n_55365));
	notech_inv i_9272(.A(\nbus_11276[4] ), .Z(n_55364));
	notech_inv i_9264(.A(n_55352), .Z(n_55356));
	notech_inv i_9263(.A(\nbus_11276[0] ), .Z(n_55352));
	notech_inv i_9255(.A(n_55341), .Z(n_55342));
	notech_inv i_9254(.A(n_27561), .Z(n_55341));
	notech_inv i_9246(.A(n_55330), .Z(n_55331));
	notech_inv i_9245(.A(n_27562), .Z(n_55330));
	notech_inv i_9243(.A(n_55312), .Z(n_55326));
	notech_inv i_9242(.A(n_55312), .Z(n_55322));
	notech_inv i_9237(.A(n_55312), .Z(n_55315));
	notech_inv i_9236(.A(gs[2]), .Z(n_55312));
	notech_inv i_9228(.A(n_55298), .Z(n_55299));
	notech_inv i_9227(.A(n_27563), .Z(n_55298));
	notech_inv i_9219(.A(n_55288), .Z(n_55289));
	notech_inv i_9218(.A(\nbus_11276[2] ), .Z(n_55288));
	notech_inv i_9210(.A(n_55276), .Z(n_55277));
	notech_inv i_9208(.A(\nbus_11276[3] ), .Z(n_55276));
	notech_inv i_9200(.A(n_55260), .Z(n_55261));
	notech_inv i_9199(.A(\nbus_11276[28] ), .Z(n_55260));
	notech_inv i_9191(.A(n_55246), .Z(n_55249));
	notech_inv i_9190(.A(\nbus_11276[29] ), .Z(n_55246));
	notech_inv i_9182(.A(n_55233), .Z(n_55234));
	notech_inv i_9181(.A(\nbus_11276[30] ), .Z(n_55233));
	notech_inv i_9171(.A(n_55213), .Z(n_55214));
	notech_inv i_9170(.A(n_301086330), .Z(n_55213));
	notech_inv i_9162(.A(n_55203), .Z(n_55204));
	notech_inv i_9160(.A(n_55243), .Z(n_55203));
	notech_inv i_9150(.A(n_55191), .Z(n_55192));
	notech_inv i_9149(.A(n_2164), .Z(n_55191));
	notech_inv i_9139(.A(n_55180), .Z(n_55181));
	notech_inv i_9138(.A(n_2319), .Z(n_55180));
	notech_inv i_9127(.A(n_55169), .Z(n_55170));
	notech_inv i_9126(.A(n_2322), .Z(n_55169));
	notech_inv i_9118(.A(n_55160), .Z(n_55161));
	notech_inv i_9117(.A(n_2156), .Z(n_55160));
	notech_inv i_9109(.A(n_55148), .Z(n_55149));
	notech_inv i_9108(.A(n_1908), .Z(n_55148));
	notech_inv i_9098(.A(n_55134), .Z(n_55136));
	notech_inv i_9096(.A(n_2323), .Z(n_55134));
	notech_inv i_9086(.A(n_55121), .Z(n_55122));
	notech_inv i_9085(.A(n_54884), .Z(n_55121));
	notech_inv i_9076(.A(n_55110), .Z(n_55111));
	notech_inv i_9075(.A(n_54735), .Z(n_55110));
	notech_inv i_9067(.A(n_55101), .Z(n_55102));
	notech_inv i_9066(.A(n_55366), .Z(n_55101));
	notech_inv i_9058(.A(n_55090), .Z(n_55091));
	notech_inv i_9057(.A(n_55619), .Z(n_55090));
	notech_inv i_9046(.A(n_55074), .Z(n_55075));
	notech_inv i_9045(.A(n_2320), .Z(n_55074));
	notech_inv i_9019(.A(n_55039), .Z(n_55040));
	notech_inv i_9018(.A(n_26763), .Z(n_55039));
	notech_inv i_8926(.A(n_54939), .Z(n_54940));
	notech_inv i_8925(.A(n_2249), .Z(n_54939));
	notech_inv i_8915(.A(n_54925), .Z(n_54926));
	notech_inv i_8914(.A(n_2248), .Z(n_54925));
	notech_inv i_8904(.A(n_54907), .Z(n_54908));
	notech_inv i_8902(.A(n_2247), .Z(n_54907));
	notech_inv i_8892(.A(n_54885), .Z(n_54887));
	notech_inv i_8891(.A(n_2313), .Z(n_54885));
	notech_inv i_8873(.A(n_54861), .Z(n_54863));
	notech_inv i_8872(.A(n_2314), .Z(n_54861));
	notech_inv i_8861(.A(n_54846), .Z(n_54847));
	notech_inv i_8860(.A(n_231547139), .Z(n_54846));
	notech_inv i_8850(.A(n_54835), .Z(n_54836));
	notech_inv i_8849(.A(n_55009), .Z(n_54835));
	notech_inv i_8803(.A(n_54783), .Z(n_54785));
	notech_inv i_8802(.A(\nbus_11354[0] ), .Z(n_54783));
	notech_inv i_8794(.A(n_54768), .Z(n_54771));
	notech_inv i_8793(.A(n_55787), .Z(n_54768));
	notech_inv i_8788(.A(n_54753), .Z(n_54762));
	notech_inv i_8782(.A(n_54753), .Z(n_54754));
	notech_inv i_8781(.A(n_54901), .Z(n_54753));
	notech_inv i_8773(.A(n_54739), .Z(n_54742));
	notech_inv i_8772(.A(n_55788), .Z(n_54739));
	notech_inv i_8762(.A(n_54726), .Z(n_54727));
	notech_inv i_8761(.A(n_55793), .Z(n_54726));
	notech_inv i_8753(.A(n_54713), .Z(n_54714));
	notech_inv i_8752(.A(n_310388585), .Z(n_54713));
	notech_inv i_8743(.A(n_54700), .Z(n_54701));
	notech_inv i_8741(.A(n_26468), .Z(n_54700));
	notech_inv i_8730(.A(n_54684), .Z(n_54685));
	notech_inv i_8729(.A(n_310188587), .Z(n_54684));
	notech_inv i_8719(.A(n_54673), .Z(n_54674));
	notech_inv i_8718(.A(n_55848), .Z(n_54673));
	notech_inv i_8707(.A(n_54658), .Z(n_54659));
	notech_inv i_8706(.A(n_55849), .Z(n_54658));
	notech_inv i_8691(.A(n_54636), .Z(n_54642));
	notech_inv i_8686(.A(n_54636), .Z(n_54637));
	notech_inv i_8685(.A(n_54687), .Z(n_54636));
	notech_inv i_8585(.A(n_54518), .Z(n_54519));
	notech_inv i_8584(.A(n_312083095), .Z(n_54518));
	notech_inv i_8581(.A(n_54497), .Z(n_54514));
	notech_inv i_8579(.A(n_54497), .Z(n_54513));
	notech_inv i_8574(.A(n_54497), .Z(n_54504));
	notech_inv i_8568(.A(n_54497), .Z(n_54498));
	notech_inv i_8567(.A(n_316283137), .Z(n_54497));
	notech_inv i_8563(.A(n_54480), .Z(n_54492));
	notech_inv i_8562(.A(n_54480), .Z(n_54491));
	notech_inv i_8557(.A(n_54480), .Z(n_54486));
	notech_inv i_8551(.A(n_54480), .Z(n_54481));
	notech_inv i_8550(.A(n_316883143), .Z(n_54480));
	notech_inv i_8542(.A(n_54471), .Z(n_54472));
	notech_inv i_8541(.A(n_311483089), .Z(n_54471));
	notech_inv i_8533(.A(n_54448), .Z(n_54449));
	notech_inv i_8531(.A(n_311383088), .Z(n_54448));
	notech_inv i_8521(.A(n_54426), .Z(n_54427));
	notech_inv i_8520(.A(n_311683091), .Z(n_54426));
	notech_inv i_8510(.A(n_54415), .Z(n_54416));
	notech_inv i_8509(.A(n_311783092), .Z(n_54415));
	notech_inv i_8498(.A(n_54404), .Z(n_54405));
	notech_inv i_8497(.A(n_311583090), .Z(n_54404));
	notech_inv i_8495(.A(\nbus_11342[0] ), .Z(n_54401));
	notech_inv i_8493(.A(\nbus_11342[0] ), .Z(n_54399));
	notech_inv i_8489(.A(\nbus_11342[0] ), .Z(n_54396));
	notech_inv i_8487(.A(\nbus_11342[0] ), .Z(n_54394));
	notech_inv i_8481(.A(n_54377), .Z(n_54389));
	notech_inv i_8480(.A(n_54377), .Z(n_54388));
	notech_inv i_8475(.A(n_54377), .Z(n_54383));
	notech_inv i_8469(.A(n_54377), .Z(n_54378));
	notech_inv i_8468(.A(n_179381781), .Z(n_54377));
	notech_inv i_8465(.A(n_54363), .Z(n_54374));
	notech_inv i_8464(.A(n_54363), .Z(n_54373));
	notech_inv i_8460(.A(n_54363), .Z(n_54369));
	notech_inv i_8456(.A(n_54363), .Z(n_54365));
	notech_inv i_8455(.A(n_54363), .Z(n_54364));
	notech_inv i_8454(.A(n_230585627), .Z(n_54363));
	notech_inv i_8452(.A(\nbus_11277[0] ), .Z(n_54360));
	notech_inv i_8449(.A(\nbus_11277[0] ), .Z(n_54358));
	notech_inv i_8446(.A(\nbus_11277[0] ), .Z(n_54355));
	notech_inv i_8444(.A(\nbus_11277[0] ), .Z(n_54353));
	notech_inv i_8435(.A(n_54343), .Z(n_54344));
	notech_inv i_8433(.A(n_172881716), .Z(n_54343));
	notech_inv i_8425(.A(n_54334), .Z(n_54335));
	notech_inv i_8424(.A(n_119181179), .Z(n_54334));
	notech_inv i_8252(.A(n_54157), .Z(n_54158));
	notech_inv i_8251(.A(n_27163), .Z(n_54157));
	notech_inv i_8243(.A(n_54147), .Z(n_54148));
	notech_inv i_8241(.A(n_55142), .Z(n_54147));
	notech_inv i_8231(.A(n_54136), .Z(n_54137));
	notech_inv i_8230(.A(n_27035), .Z(n_54136));
	notech_inv i_8220(.A(n_54123), .Z(n_54128));
	notech_inv i_8214(.A(n_54123), .Z(n_54124));
	notech_inv i_8213(.A(n_1416), .Z(n_54123));
	notech_inv i_8203(.A(n_54111), .Z(n_54112));
	notech_inv i_8202(.A(n_27022), .Z(n_54111));
	notech_inv i_8192(.A(n_54100), .Z(n_54101));
	notech_inv i_8190(.A(n_27000), .Z(n_54100));
	notech_inv i_8182(.A(n_54091), .Z(n_54092));
	notech_inv i_8181(.A(n_56024), .Z(n_54091));
	notech_inv i_8171(.A(n_54079), .Z(n_54080));
	notech_inv i_8170(.A(n_55977), .Z(n_54079));
	notech_inv i_8160(.A(n_54065), .Z(n_54066));
	notech_inv i_8158(.A(n_262636781), .Z(n_54065));
	notech_inv i_8148(.A(n_54054), .Z(n_54055));
	notech_inv i_8147(.A(\nbus_11309[0] ), .Z(n_54054));
	notech_inv i_8139(.A(n_54045), .Z(n_54046));
	notech_inv i_8138(.A(n_54707), .Z(n_54045));
	notech_inv i_8128(.A(n_54034), .Z(n_54035));
	notech_inv i_8126(.A(\nbus_11331[0] ), .Z(n_54034));
	notech_inv i_8116(.A(n_54023), .Z(n_54024));
	notech_inv i_8115(.A(n_321788473), .Z(n_54023));
	notech_inv i_8107(.A(n_54014), .Z(n_54015));
	notech_inv i_8106(.A(n_232761396), .Z(n_54014));
	notech_inv i_8096(.A(n_54003), .Z(n_54004));
	notech_inv i_8094(.A(\nbus_11310[0] ), .Z(n_54003));
	notech_inv i_8084(.A(n_53992), .Z(n_53993));
	notech_inv i_8083(.A(n_262336778), .Z(n_53992));
	notech_inv i_8073(.A(n_53981), .Z(n_53982));
	notech_inv i_8072(.A(n_26881), .Z(n_53981));
	notech_inv i_8064(.A(n_53972), .Z(n_53973));
	notech_inv i_8062(.A(n_135360435), .Z(n_53972));
	notech_inv i_8054(.A(n_53963), .Z(n_53964));
	notech_inv i_8053(.A(n_170860790), .Z(n_53963));
	notech_inv i_8045(.A(n_53954), .Z(n_53955));
	notech_inv i_8044(.A(n_170960791), .Z(n_53954));
	notech_inv i_8036(.A(n_53945), .Z(n_53946));
	notech_inv i_8035(.A(n_171060792), .Z(n_53945));
	notech_inv i_8027(.A(n_53936), .Z(n_53937));
	notech_inv i_8026(.A(n_171160793), .Z(n_53936));
	notech_inv i_8015(.A(n_53925), .Z(n_53926));
	notech_inv i_8013(.A(n_26852), .Z(n_53925));
	notech_inv i_8003(.A(n_53914), .Z(n_53915));
	notech_inv i_8002(.A(n_26844), .Z(n_53914));
	notech_inv i_7994(.A(n_53905), .Z(n_53906));
	notech_inv i_7993(.A(n_176260844), .Z(n_53905));
	notech_inv i_7983(.A(n_53894), .Z(n_53895));
	notech_inv i_7981(.A(\nbus_11350[0] ), .Z(n_53894));
	notech_inv i_7971(.A(n_53883), .Z(n_53884));
	notech_inv i_7970(.A(\nbus_11351[0] ), .Z(n_53883));
	notech_inv i_7952(.A(n_53863), .Z(n_53864));
	notech_inv i_7951(.A(\nbus_11274[0] ), .Z(n_53863));
	notech_inv i_7940(.A(n_53852), .Z(n_53853));
	notech_inv i_7939(.A(n_301186331), .Z(n_53852));
	notech_inv i_7931(.A(n_53843), .Z(n_53844));
	notech_inv i_7930(.A(n_55901), .Z(n_53843));
	notech_inv i_7920(.A(n_53832), .Z(n_53833));
	notech_inv i_7919(.A(n_26800), .Z(n_53832));
	notech_inv i_7860(.A(n_53715), .Z(n_53716));
	notech_inv i_7859(.A(n_300886328), .Z(n_53715));
	notech_inv i_7849(.A(n_53704), .Z(n_53705));
	notech_inv i_7848(.A(n_300986329), .Z(n_53704));
	notech_inv i_7808(.A(n_53660), .Z(n_53661));
	notech_inv i_7807(.A(\nbus_11323[0] ), .Z(n_53660));
	notech_inv i_7796(.A(n_53649), .Z(n_53650));
	notech_inv i_7795(.A(n_237585695), .Z(n_53649));
	notech_inv i_7787(.A(n_53640), .Z(n_53641));
	notech_inv i_7786(.A(n_265085970), .Z(n_53640));
	notech_inv i_7776(.A(n_53629), .Z(n_53630));
	notech_inv i_7775(.A(n_335083325), .Z(n_53629));
	notech_inv i_7746(.A(n_53556), .Z(n_53557));
	notech_inv i_7745(.A(n_299986319), .Z(n_53556));
	notech_inv i_7665(.A(n_53350), .Z(n_53351));
	notech_inv i_7664(.A(n_27366), .Z(n_53350));
	notech_inv i_7634(.A(n_53317), .Z(n_53318));
	notech_inv i_7633(.A(n_152160603), .Z(n_53317));
	notech_inv i_7623(.A(n_53306), .Z(n_53307));
	notech_inv i_7622(.A(n_21051), .Z(n_53306));
	notech_inv i_7611(.A(n_53295), .Z(n_53296));
	notech_inv i_7610(.A(n_28442003), .Z(n_53295));
	notech_inv i_7600(.A(n_53284), .Z(n_53285));
	notech_inv i_7599(.A(n_27341992), .Z(n_53284));
	notech_inv i_7591(.A(n_53275), .Z(n_53276));
	notech_inv i_7590(.A(n_26595), .Z(n_53275));
	notech_inv i_7579(.A(n_53264), .Z(n_53265));
	notech_inv i_7578(.A(n_151760599), .Z(n_53264));
	notech_inv i_7570(.A(n_53255), .Z(n_53256));
	notech_inv i_7569(.A(n_151960601), .Z(n_53255));
	notech_inv i_7559(.A(n_53244), .Z(n_53245));
	notech_inv i_7558(.A(n_152060602), .Z(n_53244));
	notech_inv i_7547(.A(n_53233), .Z(n_53234));
	notech_inv i_7546(.A(n_56153), .Z(n_53233));
	notech_inv i_7436(.A(n_53112), .Z(n_53113));
	notech_inv i_7435(.A(n_151260594), .Z(n_53112));
	notech_inv i_7376(.A(n_53050), .Z(n_53051));
	notech_inv i_7375(.A(n_151060592), .Z(n_53050));
	notech_inv i_7264(.A(n_52929), .Z(n_52930));
	notech_inv i_7263(.A(n_56150), .Z(n_52929));
	notech_inv i_7155(.A(n_52810), .Z(n_52811));
	notech_inv i_7154(.A(n_150960591), .Z(n_52810));
	notech_inv i_7143(.A(n_52799), .Z(n_52800));
	notech_inv i_7142(.A(n_56147), .Z(n_52799));
	notech_inv i_7034(.A(n_52680), .Z(n_52681));
	notech_inv i_7033(.A(n_150660588), .Z(n_52680));
	notech_inv i_7022(.A(n_52669), .Z(n_52670));
	notech_inv i_7021(.A(n_150760589), .Z(n_52669));
	notech_inv i_7011(.A(n_52658), .Z(n_52659));
	notech_inv i_7010(.A(n_56160), .Z(n_52658));
	notech_inv i_6903(.A(n_52539), .Z(n_52540));
	notech_inv i_6901(.A(n_150460586), .Z(n_52539));
	notech_inv i_6891(.A(n_52528), .Z(n_52529));
	notech_inv i_6890(.A(\nbus_11327[0] ), .Z(n_52528));
	notech_inv i_6880(.A(n_52517), .Z(n_52518));
	notech_inv i_6879(.A(n_223485557), .Z(n_52517));
	notech_inv i_6877(.A(n_52511), .Z(n_52515));
	notech_inv i_6876(.A(n_52511), .Z(n_52514));
	notech_inv i_6875(.A(n_52511), .Z(n_52513));
	notech_inv i_6874(.A(n_52511), .Z(n_52512));
	notech_inv i_6873(.A(n_197285298), .Z(n_52511));
	notech_inv i_6872(.A(n_52506), .Z(n_52510));
	notech_inv i_6871(.A(n_52506), .Z(n_52509));
	notech_inv i_6869(.A(n_52506), .Z(n_52508));
	notech_inv i_6868(.A(n_52506), .Z(n_52507));
	notech_inv i_6867(.A(n_197285298), .Z(n_52506));
	notech_inv i_6866(.A(n_52501), .Z(n_52504));
	notech_inv i_6865(.A(n_52501), .Z(n_52503));
	notech_inv i_6864(.A(n_52501), .Z(n_52502));
	notech_inv i_6863(.A(n_197185297), .Z(n_52501));
	notech_inv i_6861(.A(n_52497), .Z(n_52500));
	notech_inv i_6860(.A(n_52497), .Z(n_52499));
	notech_inv i_6859(.A(n_52497), .Z(n_52498));
	notech_inv i_6858(.A(n_197185297), .Z(n_52497));
	notech_inv i_6857(.A(n_52491), .Z(n_52495));
	notech_inv i_6856(.A(n_52491), .Z(n_52494));
	notech_inv i_6855(.A(n_52491), .Z(n_52493));
	notech_inv i_6853(.A(n_52491), .Z(n_52492));
	notech_inv i_6852(.A(n_196985295), .Z(n_52491));
	notech_inv i_6851(.A(n_52486), .Z(n_52490));
	notech_inv i_6850(.A(n_52486), .Z(n_52489));
	notech_inv i_6849(.A(n_52486), .Z(n_52488));
	notech_inv i_6848(.A(n_52486), .Z(n_52487));
	notech_inv i_6847(.A(n_196985295), .Z(n_52486));
	notech_inv i_6845(.A(n_52481), .Z(n_52484));
	notech_inv i_6844(.A(n_52481), .Z(n_52483));
	notech_inv i_6843(.A(n_52481), .Z(n_52482));
	notech_inv i_6842(.A(n_196785293), .Z(n_52481));
	notech_inv i_6841(.A(n_52477), .Z(n_52480));
	notech_inv i_6840(.A(n_52477), .Z(n_52479));
	notech_inv i_6839(.A(n_52477), .Z(n_52478));
	notech_inv i_6837(.A(n_196785293), .Z(n_52477));
	notech_inv i_6836(.A(n_52471), .Z(n_52475));
	notech_inv i_6835(.A(n_52471), .Z(n_52474));
	notech_inv i_6834(.A(n_52471), .Z(n_52473));
	notech_inv i_6833(.A(n_52471), .Z(n_52472));
	notech_inv i_6832(.A(n_196385289), .Z(n_52471));
	notech_inv i_6831(.A(n_52466), .Z(n_52470));
	notech_inv i_6829(.A(n_52466), .Z(n_52469));
	notech_inv i_6828(.A(n_52466), .Z(n_52468));
	notech_inv i_6827(.A(n_52466), .Z(n_52467));
	notech_inv i_6826(.A(n_196385289), .Z(n_52466));
	notech_inv i_6825(.A(n_52461), .Z(n_52464));
	notech_inv i_6824(.A(n_52461), .Z(n_52463));
	notech_inv i_6823(.A(n_52461), .Z(n_52462));
	notech_inv i_6821(.A(n_196185287), .Z(n_52461));
	notech_inv i_6820(.A(n_52457), .Z(n_52460));
	notech_inv i_6819(.A(n_52457), .Z(n_52459));
	notech_inv i_6818(.A(n_52457), .Z(n_52458));
	notech_inv i_6817(.A(n_196185287), .Z(n_52457));
	notech_inv i_6816(.A(n_52451), .Z(n_52455));
	notech_inv i_6815(.A(n_52451), .Z(n_52454));
	notech_inv i_6813(.A(n_52451), .Z(n_52453));
	notech_inv i_6812(.A(n_52451), .Z(n_52452));
	notech_inv i_6811(.A(n_195585281), .Z(n_52451));
	notech_inv i_6810(.A(n_52446), .Z(n_52450));
	notech_inv i_6809(.A(n_52446), .Z(n_52449));
	notech_inv i_6808(.A(n_52446), .Z(n_52448));
	notech_inv i_6807(.A(n_52446), .Z(n_52447));
	notech_inv i_6805(.A(n_195585281), .Z(n_52446));
	notech_inv i_6804(.A(n_52440), .Z(n_52444));
	notech_inv i_6803(.A(n_52440), .Z(n_52443));
	notech_inv i_6802(.A(n_52440), .Z(n_52442));
	notech_inv i_6801(.A(n_52440), .Z(n_52441));
	notech_inv i_6800(.A(n_195685282), .Z(n_52440));
	notech_inv i_6799(.A(n_52435), .Z(n_52439));
	notech_inv i_6797(.A(n_52435), .Z(n_52438));
	notech_inv i_6796(.A(n_52435), .Z(n_52437));
	notech_inv i_6795(.A(n_52435), .Z(n_52436));
	notech_inv i_6794(.A(n_195685282), .Z(n_52435));
	notech_inv i_6793(.A(n_52429), .Z(n_52433));
	notech_inv i_6792(.A(n_52429), .Z(n_52432));
	notech_inv i_6791(.A(n_52429), .Z(n_52431));
	notech_inv i_6789(.A(n_52429), .Z(n_52430));
	notech_inv i_6788(.A(n_26623), .Z(n_52429));
	notech_inv i_6787(.A(n_52424), .Z(n_52428));
	notech_inv i_6786(.A(n_52424), .Z(n_52427));
	notech_inv i_6785(.A(n_52424), .Z(n_52426));
	notech_inv i_6784(.A(n_52424), .Z(n_52425));
	notech_inv i_6783(.A(n_26623), .Z(n_52424));
	notech_inv i_6781(.A(n_52418), .Z(n_52422));
	notech_inv i_6780(.A(n_52418), .Z(n_52421));
	notech_inv i_6779(.A(n_52418), .Z(n_52419));
	notech_inv i_6778(.A(n_93942658), .Z(n_52418));
	notech_inv i_6777(.A(n_52414), .Z(n_52417));
	notech_inv i_6776(.A(n_52414), .Z(n_52416));
	notech_inv i_6775(.A(n_52414), .Z(n_52415));
	notech_inv i_6773(.A(n_93942658), .Z(n_52414));
	notech_inv i_6772(.A(n_52408), .Z(n_52412));
	notech_inv i_6771(.A(n_52408), .Z(n_52411));
	notech_inv i_6770(.A(n_52408), .Z(n_52410));
	notech_inv i_6769(.A(n_52408), .Z(n_52409));
	notech_inv i_6768(.A(n_94242661), .Z(n_52408));
	notech_inv i_6767(.A(n_52403), .Z(n_52407));
	notech_inv i_6765(.A(n_52403), .Z(n_52406));
	notech_inv i_6764(.A(n_52403), .Z(n_52405));
	notech_inv i_6763(.A(n_52403), .Z(n_52404));
	notech_inv i_6762(.A(n_94242661), .Z(n_52403));
	notech_inv i_6761(.A(n_52398), .Z(n_52401));
	notech_inv i_6760(.A(n_52398), .Z(n_52400));
	notech_inv i_6759(.A(n_52398), .Z(n_52399));
	notech_inv i_6757(.A(n_94442663), .Z(n_52398));
	notech_inv i_6756(.A(n_52394), .Z(n_52397));
	notech_inv i_6755(.A(n_52394), .Z(n_52396));
	notech_inv i_6754(.A(n_52394), .Z(n_52395));
	notech_inv i_6753(.A(n_94442663), .Z(n_52394));
	notech_inv i_6752(.A(n_52388), .Z(n_52392));
	notech_inv i_6751(.A(n_52388), .Z(n_52391));
	notech_inv i_6749(.A(n_52388), .Z(n_52390));
	notech_inv i_6748(.A(n_52388), .Z(n_52389));
	notech_inv i_6747(.A(n_95042669), .Z(n_52388));
	notech_inv i_6746(.A(n_52383), .Z(n_52387));
	notech_inv i_6745(.A(n_52383), .Z(n_52386));
	notech_inv i_6744(.A(n_52383), .Z(n_52385));
	notech_inv i_6743(.A(n_52383), .Z(n_52384));
	notech_inv i_6741(.A(n_95042669), .Z(n_52383));
	notech_inv i_6740(.A(n_52378), .Z(n_52381));
	notech_inv i_6739(.A(n_52378), .Z(n_52380));
	notech_inv i_6738(.A(n_52378), .Z(n_52379));
	notech_inv i_6737(.A(n_95342672), .Z(n_52378));
	notech_inv i_6736(.A(n_52374), .Z(n_52377));
	notech_inv i_6735(.A(n_52374), .Z(n_52376));
	notech_inv i_6733(.A(n_52374), .Z(n_52375));
	notech_inv i_6732(.A(n_95342672), .Z(n_52374));
	notech_inv i_6731(.A(n_52368), .Z(n_52372));
	notech_inv i_6730(.A(n_52368), .Z(n_52371));
	notech_inv i_6729(.A(n_52368), .Z(n_52370));
	notech_inv i_6728(.A(n_52368), .Z(n_52369));
	notech_inv i_6727(.A(n_182885154), .Z(n_52368));
	notech_inv i_6725(.A(n_52363), .Z(n_52367));
	notech_inv i_6724(.A(n_52363), .Z(n_52366));
	notech_inv i_6723(.A(n_52363), .Z(n_52365));
	notech_inv i_6722(.A(n_52363), .Z(n_52364));
	notech_inv i_6721(.A(n_182885154), .Z(n_52363));
	notech_inv i_6720(.A(n_52249), .Z(n_52253));
	notech_inv i_6719(.A(n_52249), .Z(n_52252));
	notech_inv i_6717(.A(n_52249), .Z(n_52251));
	notech_inv i_6716(.A(n_52249), .Z(n_52250));
	notech_inv i_6715(.A(n_182985155), .Z(n_52249));
	notech_inv i_6714(.A(n_52244), .Z(n_52248));
	notech_inv i_6713(.A(n_52244), .Z(n_52247));
	notech_inv i_6712(.A(n_52244), .Z(n_52246));
	notech_inv i_6711(.A(n_52244), .Z(n_52245));
	notech_inv i_6709(.A(n_182985155), .Z(n_52244));
	notech_ao4 i_115641118(.A(n_310818885), .B(n_3214), .C(n_321588475), .D(n_310565422
		), .Z(n_317365490));
	notech_ao4 i_115241120(.A(n_131423301), .B(n_27584), .C(n_59190), .D(n_26651
		), .Z(n_317565492));
	notech_and4 i_115841116(.A(n_317565492), .B(n_317365490), .C(n_282465141
		), .D(n_282765144), .Z(n_317765494));
	notech_ao4 i_114941123(.A(n_55533), .B(\nbus_11276[18] ), .C(n_321388476
		), .D(n_29165), .Z(n_317865495));
	notech_ao4 i_114641125(.A(n_55131), .B(n_29230), .C(n_131123298), .D(nbus_11326
		[18]), .Z(n_318065497));
	notech_and4 i_115141121(.A(n_54860), .B(n_318065497), .C(n_317865495), .D
		(n_282165138), .Z(n_318265499));
	notech_and3 i_75860587(.A(n_56060), .B(n_2660), .C(n_1081), .Z(n_318365500
		));
	notech_and3 i_4539047(.A(n_56061), .B(n_318365500), .C(n_1079), .Z(n_318465501
		));
	notech_or2 i_86638258(.A(n_2177), .B(n_271888737), .Z(n_318565502));
	notech_or2 i_141537737(.A(n_55442), .B(n_271988736), .Z(n_319065507));
	notech_nao3 i_141737735(.A(opc_10[16]), .B(n_62417), .C(n_308618863), .Z
		(n_320165518));
	notech_or2 i_141637736(.A(n_55780), .B(n_272088735), .Z(n_320265519));
	notech_nand3 i_1721724(.A(n_330065604), .B(n_320265519), .C(n_319065507)
		, .Z(n_12863));
	notech_or2 i_144137713(.A(n_55519), .B(n_271888737), .Z(n_320365520));
	notech_or4 i_65260697(.A(instrc[115]), .B(instrc[112]), .C(n_274288715),
		 .D(n_2240), .Z(n_320465521));
	notech_or4 i_120555296(.A(n_56463), .B(n_264436799), .C(n_177764115), .D
		(instrc[119]), .Z(n_320565522));
	notech_or4 i_455290(.A(n_56463), .B(n_264436799), .C(n_178164119), .D(instrc
		[119]), .Z(n_320665523));
	notech_nand2 i_144037714(.A(sav_esp[14]), .B(n_60591), .Z(n_321565532)
		);
	notech_or4 i_144237712(.A(n_274288715), .B(n_56120), .C(n_2240), .D(n_272188734
		), .Z(n_321665533));
	notech_nand3 i_1521722(.A(n_331165615), .B(n_331065614), .C(n_320365520)
		, .Z(n_12851));
	notech_or2 i_151337642(.A(n_323365550), .B(n_2700), .Z(n_321965536));
	notech_or4 i_151537640(.A(n_56086), .B(n_56120), .C(n_55523), .D(n_2648)
		, .Z(n_322265539));
	notech_or2 i_151637639(.A(n_328565589), .B(nbus_11326[17]), .Z(n_322365540
		));
	notech_or2 i_151037645(.A(n_322965546), .B(n_28987), .Z(n_322665543));
	notech_or2 i_151137644(.A(n_323065547), .B(\nbus_11276[17] ), .Z(n_322765544
		));
	notech_nand2 i_1821917(.A(n_332065624), .B(n_321965536), .Z(n_12151));
	notech_or4 i_58963601(.A(instrc[115]), .B(instrc[112]), .C(n_56081), .D(n_56375
		), .Z(n_322865545));
	notech_and3 i_86939142(.A(n_2662), .B(n_101413408), .C(n_327765581), .Z(n_322965546
		));
	notech_and3 i_78739140(.A(n_56057), .B(n_328165585), .C(n_339065692), .Z
		(n_323065547));
	notech_ao4 i_78639139(.A(n_2658), .B(n_56029), .C(n_55325), .D(n_59926),
		 .Z(n_323165548));
	notech_nor2 i_153137624(.A(n_323365550), .B(n_271988736), .Z(n_323265549
		));
	notech_and3 i_86839141(.A(n_2663), .B(n_101213406), .C(n_327965583), .Z(n_323365550
		));
	notech_nand3 i_152637629(.A(n_1416), .B(tsc[48]), .C(n_59847), .Z(n_323465551
		));
	notech_or2 i_153437621(.A(n_328565589), .B(nbus_11326[16]), .Z(n_323665553
		));
	notech_or2 i_153037625(.A(n_323165548), .B(nbus_11273[16]), .Z(n_323765554
		));
	notech_ao3 i_153237623(.A(opc_10[16]), .B(opcode_289113), .C(n_328665590
		), .Z(n_324088257));
	notech_nor2 i_153337622(.A(n_272088735), .B(n_328765591), .Z(n_324165557
		));
	notech_or4 i_1721916(.A(n_324088257), .B(n_332765631), .C(n_324165557), 
		.D(n_323265549), .Z(n_12145));
	notech_or2 i_135060568(.A(n_2689), .B(n_142263760), .Z(n_324288256));
	notech_or2 i_123663595(.A(n_2689), .B(n_56025), .Z(n_324388255));
	notech_nand3 i_154537610(.A(n_1416), .B(tsc[46]), .C(n_59847), .Z(n_324488254
		));
	notech_nao3 i_155137604(.A(n_62409), .B(opc[14]), .C(n_324288256), .Z(n_324965560
		));
	notech_nao3 i_155237603(.A(opc_10[14]), .B(opcode_289113), .C(n_324388255
		), .Z(n_325088251));
	notech_or2 i_155037605(.A(n_2663), .B(n_271888737), .Z(n_325165561));
	notech_or4 i_155337602(.A(instrc[115]), .B(instrc[112]), .C(n_56081), .D
		(n_80913203), .Z(n_325265562));
	notech_nao3 i_1521914(.A(n_325265562), .B(n_333765641), .C(n_5990), .Z(n_12133
		));
	notech_or2 i_216436998(.A(n_321288477), .B(n_271988736), .Z(n_325388250)
		);
	notech_nand2 i_215937003(.A(sav_ecx[16]), .B(n_60591), .Z(n_325788247)
		);
	notech_nao3 i_216336999(.A(n_26549), .B(opc[16]), .C(n_316988520), .Z(n_325888246
		));
	notech_or2 i_216037002(.A(n_321388476), .B(n_29004), .Z(n_325988245));
	notech_nao3 i_216636996(.A(opc_10[16]), .B(n_62417), .C(n_321588475), .Z
		(n_326265566));
	notech_or2 i_216536997(.A(n_3214), .B(n_272088735), .Z(n_326365567));
	notech_nand3 i_1716666(.A(n_334765651), .B(n_326365567), .C(n_325388250)
		, .Z(n_11788));
	notech_nao3 i_224536917(.A(n_62409), .B(opc[14]), .C(n_336265664), .Z(n_327065574
		));
	notech_nao3 i_224636916(.A(opc_10[14]), .B(n_62417), .C(n_336065662), .Z
		(n_327165575));
	notech_or2 i_224436918(.A(n_350965798), .B(n_271888737), .Z(n_327265576)
		);
	notech_or4 i_224736915(.A(n_59264), .B(n_59272), .C(n_56120), .D(n_80913203
		), .Z(n_327365577));
	notech_nao3 i_1517241(.A(n_327365577), .B(n_335865660), .C(n_5990), .Z(n_15858
		));
	notech_and3 i_105460669(.A(n_339065692), .B(n_328165585), .C(n_327965583
		), .Z(n_327465578));
	notech_and2 i_94360680(.A(n_327765581), .B(n_2657), .Z(n_327565579));
	notech_and2 i_61960699(.A(n_322865545), .B(n_142563763), .Z(n_327665580)
		);
	notech_or2 i_74260694(.A(n_2658), .B(n_318365500), .Z(n_327765581));
	notech_or4 i_74360693(.A(n_2740), .B(n_1076), .C(n_60530), .D(n_318365500
		), .Z(n_327965583));
	notech_or4 i_9281(.A(n_2740), .B(n_1076), .C(n_56029), .D(n_60530), .Z(n_328165585
		));
	notech_or4 i_8439009(.A(n_56463), .B(n_56029), .C(n_1189), .D(n_60511), 
		.Z(n_328565589));
	notech_or2 i_7939014(.A(n_2689), .B(n_318465501), .Z(n_328665590));
	notech_or4 i_8139012(.A(instrc[115]), .B(instrc[112]), .C(n_56086), .D(n_55523
		), .Z(n_328765591));
	notech_ao4 i_86738257(.A(n_254834174), .B(\nbus_11276[14] ), .C(n_2331),
		 .D(n_29006), .Z(n_328865592));
	notech_ao4 i_87038256(.A(n_59847), .B(n_27533), .C(n_2333), .D(nbus_11273
		[14]), .Z(n_328965593));
	notech_nand3 i_64839081(.A(n_328965593), .B(n_328865592), .C(n_318565502
		), .Z(n_5990));
	notech_ao4 i_142037732(.A(n_55535), .B(\nbus_11276[16] ), .C(n_55536), .D
		(nbus_11273[16]), .Z(n_329165595));
	notech_ao4 i_142137731(.A(n_262536780), .B(n_27535), .C(n_55443), .D(n_29004
		), .Z(n_329265596));
	notech_ao4 i_142237730(.A(n_59190), .B(n_26701), .C(n_55135), .D(n_27582
		), .Z(n_329465598));
	notech_ao4 i_141837734(.A(n_55977), .B(n_28430), .C(n_262636781), .D(n_26955
		), .Z(n_329565599));
	notech_ao4 i_141937733(.A(nbus_11326[16]), .B(n_308518862), .C(n_56024),
		 .D(n_29243), .Z(n_329665600));
	notech_and3 i_142537727(.A(n_329665600), .B(n_329565599), .C(n_329465598
		), .Z(n_329865602));
	notech_and4 i_142737725(.A(n_329265596), .B(n_329165595), .C(n_320165518
		), .D(n_329865602), .Z(n_330065604));
	notech_ao4 i_144637708(.A(n_55520), .B(n_29006), .C(n_56024), .D(n_29244
		), .Z(n_330265606));
	notech_ao4 i_144737707(.A(n_55382), .B(nbus_11273[14]), .C(n_55381), .D(\nbus_11276[14] 
		), .Z(n_330365607));
	notech_ao4 i_144837706(.A(n_262536780), .B(n_27533), .C(n_55738), .D(n_27579
		), .Z(n_330565609));
	notech_ao4 i_144537709(.A(n_55977), .B(n_28428), .C(n_262636781), .D(n_26951
		), .Z(n_330665610));
	notech_and3 i_145137703(.A(n_330665610), .B(n_330565609), .C(n_321565532
		), .Z(n_330865612));
	notech_and4 i_145337701(.A(n_330365607), .B(n_330265606), .C(n_321665533
		), .D(n_330865612), .Z(n_331065614));
	notech_ao4 i_145437700(.A(n_320665523), .B(n_82713221), .C(n_320565522),
		 .D(n_82813222), .Z(n_331165615));
	notech_ao4 i_151737638(.A(n_322865545), .B(n_27583), .C(n_107626780), .D
		(n_28718), .Z(n_331365617));
	notech_and4 i_152037635(.A(n_331365617), .B(n_272488731), .C(n_322265539
		), .D(n_322365540), .Z(n_331665620));
	notech_ao4 i_152137634(.A(n_328665590), .B(n_63826342), .C(n_323165548),
		 .D(nbus_11273[17]), .Z(n_331865622));
	notech_and4 i_152437631(.A(n_331865622), .B(n_331665620), .C(n_322765544
		), .D(n_322665543), .Z(n_332065624));
	notech_ao4 i_153637619(.A(n_322865545), .B(n_27582), .C(n_59847), .D(n_27535
		), .Z(n_332265626));
	notech_and4 i_153837617(.A(n_55901), .B(n_332265626), .C(n_323465551), .D
		(n_323665553), .Z(n_332465628));
	notech_ao4 i_154037615(.A(n_323065547), .B(\nbus_11276[16] ), .C(n_322965546
		), .D(n_29004), .Z(n_332665630));
	notech_nand3 i_154137614(.A(n_332465628), .B(n_332665630), .C(n_323765554
		), .Z(n_332765631));
	notech_ao4 i_155637599(.A(n_327665580), .B(n_27579), .C(n_327565579), .D
		(nbus_11273[14]), .Z(n_333065634));
	notech_ao4 i_155537600(.A(n_327465578), .B(\nbus_11276[14] ), .C(n_2662)
		, .D(n_29006), .Z(n_333265636));
	notech_and4 i_155837597(.A(n_55901), .B(n_333265636), .C(n_333065634), .D
		(n_324488254), .Z(n_333465638));
	notech_and4 i_156137594(.A(n_324965560), .B(n_333465638), .C(n_325088251
		), .D(n_325165561), .Z(n_333765641));
	notech_ao4 i_216836994(.A(n_131423301), .B(n_27582), .C(n_170914103), .D
		(n_27535), .Z(n_333965643));
	notech_ao4 i_216736995(.A(n_55131), .B(n_29245), .C(n_1031), .D(n_60473)
		, .Z(n_334065644));
	notech_and4 i_217136991(.A(n_334065644), .B(n_333965643), .C(n_325788247
		), .D(n_325888246), .Z(n_334365647));
	notech_ao4 i_217336989(.A(n_55534), .B(nbus_11273[16]), .C(n_55533), .D(\nbus_11276[16] 
		), .Z(n_334565649));
	notech_and4 i_217536987(.A(n_334365647), .B(n_334565649), .C(n_325988245
		), .D(n_326265566), .Z(n_334765651));
	notech_ao4 i_225036912(.A(n_339065692), .B(nbus_11326[14]), .C(n_337665678
		), .D(n_27579), .Z(n_334965653));
	notech_ao4 i_224836914(.A(n_350865797), .B(n_29006), .C(n_107626780), .D
		(n_28709), .Z(n_335065654));
	notech_ao4 i_224936913(.A(n_26244), .B(nbus_11273[14]), .C(\nbus_11276[14] 
		), .D(n_26245), .Z(n_335165655));
	notech_and3 i_225236910(.A(n_335165655), .B(n_335065654), .C(n_334965653
		), .Z(n_335365657));
	notech_and4 i_225536907(.A(n_327065574), .B(n_335365657), .C(n_327165575
		), .D(n_327265576), .Z(n_335865660));
	notech_or4 i_125432977(.A(instrc[118]), .B(n_229364616), .C(n_351465803)
		, .D(instrc[119]), .Z(n_336065662));
	notech_and3 i_69632890(.A(n_354376379), .B(n_353688272), .C(n_343465724)
		, .Z(n_336165663));
	notech_or4 i_134232851(.A(instrc[118]), .B(n_229364616), .C(n_338065682)
		, .D(instrc[119]), .Z(n_336265664));
	notech_and4 i_15432725(.A(n_57419), .B(n_276588692), .C(n_2105), .D(n_55656
		), .Z(n_336365665));
	notech_and4 i_15532724(.A(n_2222), .B(n_349565784), .C(n_336165663), .D(n_339565697
		), .Z(n_336465666));
	notech_and4 i_15632723(.A(n_55684), .B(n_339065692), .C(n_55943), .D(n_350165790
		), .Z(n_336565667));
	notech_and2 i_15732722(.A(n_2157), .B(n_336765669), .Z(n_336665668));
	notech_or4 i_27032652(.A(n_275388704), .B(n_2835), .C(n_57444), .D(read_ack
		), .Z(n_336765669));
	notech_ao3 i_19132715(.A(n_2234), .B(n_349265781), .C(n_2203), .Z(n_337165673
		));
	notech_ao4 i_19232714(.A(n_26418), .B(n_54877), .C(n_2193), .D(n_2161), 
		.Z(n_337265674));
	notech_and4 i_19332713(.A(n_2168), .B(n_348965778), .C(n_57375), .D(n_26736
		), .Z(n_337365675));
	notech_and2 i_61833141(.A(n_351165800), .B(n_338465686), .Z(n_337665678)
		);
	notech_nand2 i_104733142(.A(n_55143), .B(n_213364467), .Z(n_337765679)
		);
	notech_nand2 i_104833143(.A(n_55142), .B(n_213464468), .Z(n_337865680)
		);
	notech_or4 i_45632491(.A(fsm[3]), .B(fsm[0]), .C(n_60775), .D(n_2236), .Z
		(n_337965681));
	notech_and2 i_46332484(.A(n_338165683), .B(n_351065799), .Z(n_338065682)
		);
	notech_and3 i_75749177(.A(n_56060), .B(n_213264466), .C(n_56032), .Z(n_338165683
		));
	notech_or4 i_59432401(.A(n_59263), .B(n_59272), .C(n_56120), .D(n_36952)
		, .Z(n_338465686));
	notech_and4 i_26432658(.A(n_2225), .B(n_26554), .C(n_275588702), .D(n_29376
		), .Z(n_338565687));
	notech_or4 i_54232998(.A(fsm[3]), .B(fsm[0]), .C(n_60775), .D(n_55843), 
		.Z(n_339065692));
	notech_nand2 i_26732655(.A(n_26496), .B(n_29376), .Z(n_339565697));
	notech_nand3 i_30932625(.A(n_1416), .B(tsc[15]), .C(n_59847), .Z(n_340065702
		));
	notech_or2 i_30732626(.A(n_356476400), .B(n_350965798), .Z(n_340365705)
		);
	notech_nand2 i_30332629(.A(opa[15]), .B(n_337765679), .Z(n_340665708));
	notech_or4 i_30032632(.A(n_60775), .B(n_60726), .C(n_55843), .D(nbus_11326
		[15]), .Z(n_340965711));
	notech_nand2 i_43132515(.A(sav_epc[28]), .B(n_60591), .Z(n_341265714));
	notech_or2 i_42732518(.A(n_55567), .B(nbus_11273[28]), .Z(n_342365717)
		);
	notech_or2 i_42432521(.A(n_55587), .B(n_57330), .Z(n_342765720));
	notech_nao3 i_42132524(.A(n_205688857), .B(n_6822), .C(n_205588858), .Z(n_343365723
		));
	notech_nand2 i_46032487(.A(n_26380), .B(n_29130), .Z(n_343465724));
	notech_nand2 i_25896(.A(opc_10[28]), .B(n_62417), .Z(n_343565725));
	notech_ao4 i_125883394(.A(n_55873), .B(n_29228), .C(n_55940), .D(n_27814
		), .Z(n_345465743));
	notech_ao4 i_125783395(.A(n_55998), .B(n_27981), .C(n_55872), .D(n_28015
		), .Z(n_345565744));
	notech_ao4 i_125531835(.A(n_56035), .B(n_27915), .C(n_55870), .D(n_27949
		), .Z(n_345765746));
	notech_ao4 i_125331836(.A(n_55867), .B(n_27846), .C(n_56068), .D(n_27881
		), .Z(n_345865747));
	notech_and4 i_126131834(.A(n_345865747), .B(n_345765746), .C(n_345565744
		), .D(n_345465743), .Z(n_346065749));
	notech_ao4 i_124931839(.A(n_55864), .B(n_27743), .C(n_55898), .D(n_27782
		), .Z(n_346165750));
	notech_ao4 i_124831840(.A(n_56097), .B(n_27711), .C(n_54535), .D(n_27398
		), .Z(n_346265751));
	notech_and2 i_125131838(.A(n_346265751), .B(n_346165750), .Z(n_346365752
		));
	notech_ao4 i_124631842(.A(n_56151), .B(n_27634), .C(n_54451), .D(n_27676
		), .Z(n_346465753));
	notech_ao4 i_124531843(.A(n_55878), .B(n_28047), .C(n_54439), .D(n_29229
		), .Z(n_346565754));
	notech_ao4 i_109831967(.A(n_2212), .B(nbus_11326[28]), .C(n_2211), .D(n_343565725
		), .Z(n_347065759));
	notech_ao4 i_109631969(.A(n_55811), .B(n_57306), .C(n_2345), .D(n_27551)
		, .Z(n_347265761));
	notech_and4 i_110031965(.A(n_347265761), .B(n_347065759), .C(n_342765720
		), .D(n_343365723), .Z(n_347465763));
	notech_ao4 i_109331972(.A(n_55597), .B(n_29219), .C(n_55568), .D(\nbus_11276[28] 
		), .Z(n_347565764));
	notech_ao4 i_109031974(.A(n_26435), .B(n_29246), .C(n_55842), .D(n_27596
		), .Z(n_347765766));
	notech_and4 i_109531970(.A(n_347765766), .B(n_347565764), .C(n_341265714
		), .D(n_342365717), .Z(n_347965768));
	notech_ao4 i_83532196(.A(n_177264110), .B(n_336065662), .C(n_177164109),
		 .D(n_336265664), .Z(n_348065769));
	notech_ao4 i_83332198(.A(n_337665678), .B(n_27581), .C(n_56035), .D(n_363688159
		), .Z(n_348265771));
	notech_and4 i_83832194(.A(n_348265771), .B(n_348065769), .C(n_340665708)
		, .D(n_340965711), .Z(n_348465773));
	notech_ao4 i_83032201(.A(n_350865797), .B(n_29087), .C(\nbus_11276[15] )
		, .D(n_26245), .Z(n_348565774));
	notech_and4 i_83232199(.A(n_363088165), .B(n_348565774), .C(n_340065702)
		, .D(n_340365705), .Z(n_348865777));
	notech_ao4 i_82032207(.A(n_2258), .B(n_55086), .C(n_205588858), .D(n_58945
		), .Z(n_348965778));
	notech_ao4 i_81832209(.A(n_337365675), .B(n_59926), .C(n_337265674), .D(n_275388704
		), .Z(n_349265781));
	notech_ao4 i_162832832(.A(n_60591), .B(n_337165673), .C(n_60473), .D(n_354676382
		), .Z(n_349465783));
	notech_mux2 i_79832228(.S(read_ack), .A(n_55641), .B(n_2821), .Z(n_349565784
		));
	notech_ao4 i_79032236(.A(n_335162249), .B(n_336465666), .C(n_336365665),
		 .D(n_60473), .Z(n_349865787));
	notech_ao4 i_79432232(.A(n_1907), .B(read_ack), .C(n_2193), .D(n_336665668
		), .Z(n_350065789));
	notech_and2 i_79532231(.A(n_350065789), .B(n_26608), .Z(n_350165790));
	notech_ao4 i_78932237(.A(n_2113), .B(n_614), .C(n_60591), .D(n_336565667
		), .Z(n_350465793));
	notech_nand2 i_79132235(.A(n_350465793), .B(n_349865787), .Z(n_350565794
		));
	notech_and4 i_125641019(.A(n_55901), .B(n_316965486), .C(n_307918856), .D
		(n_283065147), .Z(n_317265489));
	notech_nand3 i_620657(.A(n_131863656), .B(n_131763655), .C(n_132263660),
		 .Z(n_19815));
	notech_or4 i_620721(.A(n_130263640), .B(n_168864026), .C(n_132663664), .D
		(n_26369), .Z(n_19467));
	notech_or4 i_620817(.A(n_168864026), .B(n_129563633), .C(n_133363671), .D
		(n_26367), .Z(n_19119));
	notech_nand3 i_620945(.A(n_133963677), .B(n_133863676), .C(n_134363681),
		 .Z(n_9009));
	notech_or4 i_620977(.A(n_168864026), .B(n_128063618), .C(n_134863686), .D
		(n_26361), .Z(n_16729));
	notech_nand3 i_621041(.A(n_135463692), .B(n_135363691), .C(n_135863696),
		 .Z(n_13845));
	notech_nand3 i_621585(.A(n_136163699), .B(n_136063698), .C(n_136563703),
		 .Z(n_13145));
	notech_and4 i_621713(.A(n_137363711), .B(n_137263710), .C(n_137663714), 
		.D(n_137163709), .Z(n_12797));
	notech_and4 i_321710(.A(n_138563723), .B(n_138463722), .C(n_138363721), 
		.D(n_138863726), .Z(n_12779));
	notech_and4 i_821907(.A(n_139163729), .B(n_139363731), .C(n_139863736), 
		.D(n_123863576), .Z(n_12091));
	notech_nand2 i_621905(.A(n_140863746), .B(n_140463742), .Z(n_12079));
	notech_nand2 i_421903(.A(n_141863756), .B(n_141463752), .Z(n_12067));
	notech_and3 i_9863449(.A(n_55069), .B(n_2678), .C(n_2656), .Z(n_269939487
		));
	notech_and3 i_9963448(.A(n_55068), .B(n_2677), .C(n_2653), .Z(n_269839486
		));
	notech_and3 i_10063447(.A(n_326769066), .B(n_201467834), .C(n_54457), .Z
		(n_269739485));
	notech_ao3 i_10163446(.A(n_326669065), .B(n_54460), .C(n_201367833), .Z(n_269639484
		));
	notech_ao4 i_125441021(.A(n_328565589), .B(nbus_11326[18]), .C(n_323165548
		), .D(nbus_11273[18]), .Z(n_316965486));
	notech_and4 i_126141014(.A(n_316665483), .B(n_316465481), .C(n_283365150
		), .D(n_283665153), .Z(n_316865485));
	notech_ao4 i_125741018(.A(n_322965546), .B(n_29165), .C(n_322865545), .D
		(n_27584), .Z(n_316665483));
	notech_ao4 i_125941016(.A(n_310818885), .B(n_328765591), .C(n_310565422)
		, .D(n_328665590), .Z(n_316465481));
	notech_ao4 i_126241013(.A(n_27539), .B(n_59847), .C(n_107626780), .D(n_28719
		), .Z(n_316265479));
	notech_nand2 i_621169(.A(n_157363911), .B(n_156863906), .Z(n_13497));
	notech_and4 i_621553(.A(n_154363881), .B(n_158063918), .C(n_158363921), 
		.D(n_157963917), .Z(n_16380));
	notech_and4 i_821715(.A(n_159263930), .B(n_159163929), .C(n_159063928), 
		.D(n_159563933), .Z(n_12809));
	notech_and4 i_721714(.A(n_160463942), .B(n_160363941), .C(n_160263940), 
		.D(n_160763945), .Z(n_12803));
	notech_and4 i_521712(.A(n_161663954), .B(n_161563953), .C(n_161463952), 
		.D(n_161963957), .Z(n_12791));
	notech_and4 i_421711(.A(n_162863966), .B(n_162763965), .C(n_163163969), 
		.D(n_162663964), .Z(n_12785));
	notech_and4 i_221709(.A(n_164063978), .B(n_163963977), .C(n_163863976), 
		.D(n_164363981), .Z(n_12773));
	notech_nand3 i_621841(.A(n_164763985), .B(n_164663984), .C(n_165163989),
		 .Z(n_12431));
	notech_and4 i_1021909(.A(n_165263990), .B(n_165463992), .C(n_165963997),
		 .D(n_146663804), .Z(n_12103));
	notech_and4 i_921908(.A(n_166063998), .B(n_166264000), .C(n_166764005), 
		.D(n_145863796), .Z(n_12097));
	notech_nand2 i_3016679(.A(n_167764015), .B(n_167264010), .Z(n_11866));
	notech_nand2 i_917235(.A(n_168664024), .B(n_168264020), .Z(n_15822));
	notech_or2 i_207949248(.A(n_351565804), .B(n_351465803), .Z(n_350865797)
		);
	notech_or4 i_204549246(.A(n_212964463), .B(n_60530), .C(n_2739), .D(n_351465803
		), .Z(n_350965798));
	notech_nor2 i_128257938(.A(n_229564618), .B(n_26239), .Z(n_55097));
	notech_ao4 i_31949264(.A(n_2044), .B(n_54520), .C(n_56375), .D(n_26501),
		 .Z(n_351065799));
	notech_and2 i_147257937(.A(n_55142), .B(n_213764471), .Z(n_54948));
	notech_ao4 i_147157936(.A(n_212864462), .B(n_26303), .C(n_229564618), .D
		(n_26239), .Z(n_54949));
	notech_ao4 i_126341012(.A(n_323165548), .B(nbus_11273[19]), .C(n_323065547
		), .D(\nbus_11276[19] ), .Z(n_316065477));
	notech_and3 i_126941006(.A(n_315665473), .B(n_315865475), .C(n_284565162
		), .Z(n_315965476));
	notech_nand3 i_621297(.A(n_175064088), .B(n_174964087), .C(n_174864086),
		 .Z(n_20631));
	notech_nand2 i_817234(.A(n_176064098), .B(n_175664094), .Z(n_15816));
	notech_and4 i_617232(.A(n_176464102), .B(n_177064108), .C(n_170564043), 
		.D(n_176364101), .Z(n_15804));
	notech_ao4 i_127657868(.A(n_55854), .B(\nbus_11276[4] ), .C(n_1135), .D(n_29063
		), .Z(n_249134117));
	notech_or4 i_58849255(.A(n_59264), .B(n_59273), .C(n_56120), .D(n_56375)
		, .Z(n_351165800));
	notech_and3 i_61255357(.A(n_55135), .B(n_296165278), .C(n_280865125), .Z
		(n_55738));
	notech_or2 i_171145421(.A(n_55976), .B(n_26235), .Z(n_54749));
	notech_ao4 i_126641009(.A(n_322965546), .B(n_29167), .C(n_322865545), .D
		(n_27585), .Z(n_315865475));
	notech_or4 i_177745420(.A(n_1912), .B(n_243664753), .C(n_55976), .D(n_60530
		), .Z(n_54695));
	notech_ao4 i_83355353(.A(n_1970), .B(n_60473), .C(n_54935), .D(n_178164119
		), .Z(n_55520));
	notech_ao4 i_83455352(.A(n_54874), .B(n_56104), .C(n_260961637), .D(n_178164119
		), .Z(n_55519));
	notech_and4 i_98155343(.A(n_55790), .B(n_295965276), .C(n_54759), .D(n_189664231
		), .Z(n_55382));
	notech_and4 i_98255342(.A(n_55791), .B(n_55692), .C(n_54751), .D(n_193164266
		), .Z(n_55381));
	notech_ao4 i_126741008(.A(n_310718884), .B(n_328765591), .C(n_308065397)
		, .D(n_328665590), .Z(n_315665473));
	notech_and3 i_127341002(.A(n_315265469), .B(n_315465471), .C(n_284965166
		), .Z(n_315565472));
	notech_ao4 i_127041005(.A(n_27540), .B(n_59847), .C(n_107626780), .D(n_28720
		), .Z(n_315465471));
	notech_or4 i_9556(.A(n_1912), .B(n_243664753), .C(n_258664903), .D(n_60530
		), .Z(n_47687));
	notech_or4 i_158745423(.A(n_1912), .B(n_243664753), .C(n_60530), .D(n_26225
		), .Z(n_54852));
	notech_nor2 i_9558(.A(n_258664903), .B(n_26235), .Z(n_47685));
	notech_nand2 i_158645424(.A(n_55970), .B(n_54936), .Z(n_54853));
	notech_nand2 i_1621723(.A(n_194564280), .B(n_194064275), .Z(n_12857));
	notech_nand2 i_1321720(.A(n_195664291), .B(n_195164286), .Z(n_12839));
	notech_nand2 i_2521924(.A(n_196564300), .B(n_196164296), .Z(n_12193));
	notech_nand2 i_1621915(.A(n_197464309), .B(n_197064305), .Z(n_12139));
	notech_nand2 i_1421913(.A(n_198364318), .B(n_197964314), .Z(n_12127));
	notech_and4 i_1321912(.A(n_184064175), .B(n_198464319), .C(n_198664321),
		 .D(n_199164326), .Z(n_12121));
	notech_nand2 i_1221911(.A(n_200064335), .B(n_199664331), .Z(n_12115));
	notech_and4 i_1121910(.A(n_200164336), .B(n_200364338), .C(n_200864343),
		 .D(n_182264157), .Z(n_12109));
	notech_nand2 i_1417240(.A(n_201764352), .B(n_201364348), .Z(n_15852));
	notech_or4 i_1317239(.A(n_189974767), .B(n_179264130), .C(n_202464359), 
		.D(n_26311), .Z(n_15846));
	notech_or4 i_1217238(.A(n_239168196), .B(n_178264120), .C(n_203364368), 
		.D(n_26310), .Z(n_15840));
	notech_ao4 i_127141004(.A(n_323165548), .B(nbus_11273[20]), .C(n_323065547
		), .D(\nbus_11276[20] ), .Z(n_315265469));
	notech_ao4 i_127441001(.A(n_322965546), .B(n_29169), .C(n_322865545), .D
		(n_27586), .Z(n_315065467));
	notech_ao4 i_127541000(.A(n_310618883), .B(n_328765591), .C(n_315162155)
		, .D(n_328665590), .Z(n_314865465));
	notech_and4 i_143855363(.A(n_192664261), .B(n_192564260), .C(n_192164256
		), .D(n_192464259), .Z(n_57293));
	notech_and4 i_128140994(.A(n_55901), .B(n_314465461), .C(n_308018857), .D
		(n_285765174), .Z(n_314765464));
	notech_nand2 i_26826(.A(opc_10[5]), .B(opcode_289113), .Z(n_351265801)
		);
	notech_nand2 i_26827(.A(n_62409), .B(opc[5]), .Z(n_351365802));
	notech_ao4 i_32349263(.A(n_56502), .B(n_56551), .C(n_55859), .D(n_26501)
		, .Z(n_351465803));
	notech_and2 i_83049258(.A(n_55837), .B(n_55580), .Z(n_55523));
	notech_nor2 i_148449214(.A(n_212864462), .B(n_26303), .Z(n_351565804));
	notech_and2 i_78549250(.A(n_339065692), .B(n_213564469), .Z(n_351665805)
		);
	notech_and2 i_79049247(.A(n_350865797), .B(n_213364467), .Z(n_351765806)
		);
	notech_and2 i_79149245(.A(n_350965798), .B(n_213464468), .Z(n_351865807)
		);
	notech_nand3 i_100649235(.A(n_54642), .B(n_54762), .C(n_213564469), .Z(n_351965808
		));
	notech_ao4 i_101649233(.A(n_212864462), .B(n_26303), .C(n_229564618), .D
		(n_26248), .Z(n_352065809));
	notech_and2 i_101849231(.A(n_213764471), .B(n_355188244), .Z(n_352165810
		));
	notech_or2 i_123149224(.A(n_351565804), .B(n_351065799), .Z(n_55143));
	notech_or4 i_123249223(.A(n_212964463), .B(n_60530), .C(n_2739), .D(n_351065799
		), .Z(n_55142));
	notech_or4 i_33929(.A(n_59264), .B(n_59273), .C(n_56121), .D(n_55523), .Z
		(n_352265811));
	notech_or4 i_33915(.A(n_59264), .B(n_59273), .C(n_56120), .D(n_54367), .Z
		(n_352365812));
	notech_mux2 i_3011687(.S(n_60136), .A(regs_14[29]), .B(add_len_pc32[29])
		, .Z(n_352465813));
	notech_mux2 i_3111688(.S(n_60136), .A(regs_14[30]), .B(add_len_pc32[30])
		, .Z(n_352565814));
	notech_ao4 i_31749205(.A(n_56573), .B(n_2044), .C(n_55827), .D(n_26501),
		 .Z(n_56032));
	notech_and2 i_32149204(.A(n_56060), .B(n_213264466), .Z(n_352665815));
	notech_ao3 i_152549203(.A(n_59235), .B(n_26772), .C(n_212964463), .Z(n_54904
		));
	notech_or4 i_24249190(.A(instrc[118]), .B(n_56463), .C(n_56492), .D(instrc
		[119]), .Z(n_352765816));
	notech_or4 i_108749169(.A(instrc[118]), .B(n_229364616), .C(n_213864472)
		, .D(instrc[119]), .Z(n_352865817));
	notech_or4 i_141649162(.A(instrc[118]), .B(n_229364616), .C(instrc[119])
		, .D(n_213964473), .Z(n_352965818));
	notech_nand2 i_80439123(.A(n_322088470), .B(n_56057), .Z(n_353065819));
	notech_and3 i_89239125(.A(n_101413408), .B(n_54431), .C(n_323088460), .Z
		(n_353165820));
	notech_and2 i_80339122(.A(n_98113375), .B(n_97522962), .Z(n_353265821)
		);
	notech_and3 i_89139124(.A(n_101213406), .B(n_322988461), .C(n_54455), .Z
		(n_353365822));
	notech_or2 i_57755323(.A(n_56375), .B(n_55898), .Z(n_55772));
	notech_or2 i_31421(.A(n_55523), .B(n_55893), .Z(n_322631613));
	notech_nao3 i_31410(.A(n_56492), .B(n_268064997), .C(n_177364111), .Z(n_322931616
		));
	notech_nao3 i_4545332(.A(n_56492), .B(n_268064997), .C(n_242164740), .Z(n_302621913
		));
	notech_and3 i_79455354(.A(n_54852), .B(n_47687), .C(n_54695), .Z(n_55556
		));
	notech_ao3 i_79355355(.A(n_54853), .B(n_54749), .C(n_47685), .Z(n_55557)
		);
	notech_or2 i_63239105(.A(n_56375), .B(n_56049), .Z(n_353465823));
	notech_and3 i_102345413(.A(n_47687), .B(n_54695), .C(n_54852), .Z(n_55346
		));
	notech_ao3 i_102245412(.A(n_54749), .B(n_54853), .C(n_47685), .Z(n_55347
		));
	notech_and4 i_93945436(.A(n_267764994), .B(n_267664993), .C(n_267264989)
		, .D(n_267564992), .Z(n_57330));
	notech_ao4 i_37545426(.A(n_2044), .B(n_54520), .C(n_56375), .D(n_26512),
		 .Z(n_55974));
	notech_nand2 i_37945394(.A(n_56061), .B(n_243864755), .Z(n_55970));
	notech_ao4 i_37345395(.A(n_56573), .B(n_2044), .C(n_55827), .D(n_26512),
		 .Z(n_55976));
	notech_nand2 i_148845411(.A(n_268164998), .B(n_56260), .Z(n_54936));
	notech_mux2 i_2411681(.S(n_60136), .A(regs_14[23]), .B(add_len_pc32[23])
		, .Z(\add_len_pc[23] ));
	notech_mux2 i_2611683(.S(n_60136), .A(regs_14[25]), .B(add_len_pc32[25])
		, .Z(\add_len_pc[25] ));
	notech_or4 i_115145397(.A(n_1912), .B(n_243664753), .C(n_55974), .D(n_60530
		), .Z(n_55221));
	notech_or2 i_115245396(.A(n_55974), .B(n_26235), .Z(n_55220));
	notech_and4 i_93629160(.A(n_266364980), .B(n_266264979), .C(n_265864975)
		, .D(n_266164978), .Z(n_308821975));
	notech_and4 i_144845388(.A(n_269465011), .B(n_269365010), .C(n_268965006
		), .D(n_269265009), .Z(n_308421971));
	notech_nand2 i_2620645(.A(n_270665023), .B(n_270165018), .Z(n_20261));
	notech_nand2 i_2420643(.A(n_273165048), .B(n_272665043), .Z(n_20249));
	notech_or4 i_2921928(.A(n_313168930), .B(n_252064837), .C(n_273565052), 
		.D(n_26299), .Z(n_12217));
	notech_and4 i_2821927(.A(n_274465061), .B(n_274665063), .C(n_274365060),
		 .D(n_251364830), .Z(n_12211));
	notech_or4 i_2721926(.A(n_265975498), .B(n_250264819), .C(n_275165068), 
		.D(n_26298), .Z(n_12205));
	notech_or4 i_2621925(.A(n_173971058), .B(n_249464811), .C(n_275865075), 
		.D(n_26297), .Z(n_12199));
	notech_and4 i_2421923(.A(n_276665083), .B(n_276865085), .C(n_248864805),
		 .D(n_276565082), .Z(n_12187));
	notech_and4 i_2916678(.A(n_277565092), .B(n_277765094), .C(n_277465091),
		 .D(n_247864795), .Z(n_11860));
	notech_nand2 i_2816677(.A(n_278865105), .B(n_278365100), .Z(n_11854));
	notech_nand2 i_2716676(.A(n_279865115), .B(n_279365110), .Z(n_11848));
	notech_and4 i_2616675(.A(n_280465121), .B(n_280665123), .C(n_280365120),
		 .D(n_244564762), .Z(n_11842));
	notech_or2 i_3745340(.A(n_258764904), .B(n_55974), .Z(n_303421921));
	notech_ao4 i_127940996(.A(n_328565589), .B(nbus_11326[21]), .C(n_323165548
		), .D(nbus_11273[21]), .Z(n_314465461));
	notech_and4 i_145133114(.A(n_346565754), .B(n_346465753), .C(n_346065749
		), .D(n_346365752), .Z(n_57306));
	notech_and4 i_128640989(.A(n_314165458), .B(n_313965456), .C(n_286065177
		), .D(n_286365180), .Z(n_314365460));
	notech_and4 i_144645389(.A(n_271965036), .B(n_271865035), .C(n_271465031
		), .D(n_271765034), .Z(n_308521972));
	notech_and4 i_93429158(.A(n_264964966), .B(n_264864965), .C(n_264464961)
		, .D(n_264764964), .Z(n_308921976));
	notech_ao4 i_128240993(.A(n_322965546), .B(n_29172), .C(n_322865545), .D
		(n_27588), .Z(n_314165458));
	notech_and3 i_56942292(.A(n_320465521), .B(n_296165278), .C(n_280865125)
		, .Z(n_55780));
	notech_and3 i_91342287(.A(n_295965276), .B(n_55978), .C(n_296065277), .Z
		(n_55443));
	notech_and3 i_91542286(.A(n_295765274), .B(n_55979), .C(n_295865275), .Z
		(n_55442));
	notech_mux2 i_1911676(.S(n_60136), .A(regs_14[18]), .B(add_len_pc32[18])
		, .Z(\add_len_pc[18] ));
	notech_mux2 i_2011677(.S(n_60136), .A(regs_14[19]), .B(add_len_pc32[19])
		, .Z(\add_len_pc[19] ));
	notech_mux2 i_2311680(.S(n_60136), .A(regs_14[22]), .B(add_len_pc32[22])
		, .Z(\add_len_pc[22] ));
	notech_nand2 i_2320642(.A(n_307965396), .B(n_307465391), .Z(n_20243));
	notech_nand2 i_2020639(.A(n_310465421), .B(n_309965416), .Z(n_20225));
	notech_nand2 i_1920638(.A(n_312965446), .B(n_312465441), .Z(n_20219));
	notech_nand2 i_2321922(.A(n_313865455), .B(n_313465451), .Z(n_12181));
	notech_nand2 i_2221921(.A(n_314765464), .B(n_314365460), .Z(n_12175));
	notech_and4 i_2121920(.A(n_314865465), .B(n_315065467), .C(n_315565472),
		 .D(n_285465171), .Z(n_12169));
	notech_and4 i_2021919(.A(n_316065477), .B(n_316265479), .C(n_284065157),
		 .D(n_315965476), .Z(n_12163));
	notech_nand2 i_1921918(.A(n_317265489), .B(n_316865485), .Z(n_12157));
	notech_nand2 i_1916668(.A(n_318265499), .B(n_317765494), .Z(n_11800));
	notech_or4 i_114842241(.A(n_56463), .B(n_264436799), .C(n_281665133), .D
		(instrc[119]), .Z(n_308618863));
	notech_and4 i_144142263(.A(n_311765434), .B(n_311665433), .C(n_311265429
		), .D(n_311565432), .Z(n_310818885));
	notech_and4 i_92929153(.A(n_302165338), .B(n_302065337), .C(n_301665333)
		, .D(n_301965336), .Z(n_311318890));
	notech_and4 i_144242262(.A(n_309265409), .B(n_309165408), .C(n_308765404
		), .D(n_309065407), .Z(n_310718884));
	notech_and4 i_93029154(.A(n_303565352), .B(n_303465351), .C(n_303065347)
		, .D(n_303365350), .Z(n_311218889));
	notech_and4 i_144542259(.A(n_306765384), .B(n_306665383), .C(n_306265379
		), .D(n_306565382), .Z(n_310418881));
	notech_nand2 i_93329157(.A(n_305165368), .B(n_304465361), .Z(n_310918886
		));
	notech_ao4 i_128440991(.A(n_310518882), .B(n_328765591), .C(n_312662130)
		, .D(n_328665590), .Z(n_313965456));
	notech_and4 i_129040985(.A(n_55901), .B(n_313565452), .C(n_308218859), .D
		(n_286665183), .Z(n_313865455));
	notech_ao4 i_81939150(.A(n_316988520), .B(n_320888481), .C(n_54688), .D(n_60473
		), .Z(n_55533));
	notech_ao4 i_81839149(.A(n_316988520), .B(n_54938), .C(n_55325), .D(n_60473
		), .Z(n_55534));
	notech_or4 i_27361(.A(n_60752), .B(n_60739), .C(n_60775), .D(n_1970), .Z
		(n_2331));
	notech_or4 i_27355(.A(fsm[3]), .B(fsm[0]), .C(n_60775), .D(n_55001), .Z(n_2333
		));
	notech_or2 i_69433153(.A(n_2226), .B(n_2647), .Z(n_55656));
	notech_and3 i_129333144(.A(n_2180), .B(n_2192), .C(n_2325), .Z(n_55086)
		);
	notech_mux2 i_2911686(.S(n_60136), .A(regs_14[28]), .B(add_len_pc32[28])
		, .Z(\add_len_pc[28] ));
	notech_or4 i_66633109(.A(n_56117), .B(n_2572), .C(n_274988708), .D(n_59922
		), .Z(n_55684));
	notech_ao4 i_128840987(.A(n_328565589), .B(nbus_11326[22]), .C(n_323165548
		), .D(nbus_11273[22]), .Z(n_313565452));
	notech_and4 i_129540980(.A(n_313265449), .B(n_313065447), .C(n_286965186
		), .D(n_287265189), .Z(n_313465451));
	notech_ao4 i_129140984(.A(n_322965546), .B(n_29174), .C(n_322865545), .D
		(n_27589), .Z(n_313265449));
	notech_ao4 i_129340982(.A(n_310418881), .B(n_328765591), .C(n_305565372)
		, .D(n_328665590), .Z(n_313065447));
	notech_and4 i_187940413(.A(n_312765444), .B(n_312565442), .C(n_287565192
		), .D(n_287865195), .Z(n_312965446));
	notech_ao4 i_187540417(.A(n_55567), .B(nbus_11273[18]), .C(n_55568), .D(\nbus_11276[18] 
		), .Z(n_312765444));
	notech_nand2 i_59132974(.A(n_54967), .B(n_337965681), .Z(n_55758));
	notech_or4 i_142133152(.A(n_274588712), .B(n_2572), .C(n_272988726), .D(n_59922
		), .Z(n_54967));
	notech_nand2 i_2920648(.A(n_347965768), .B(n_347465763), .Z(n_20279));
	notech_nand2 i_1617242(.A(n_348865777), .B(n_348465773), .Z(n_15864));
	notech_or4 i_126951(.A(n_26232), .B(n_338565687), .C(n_26420), .D(n_350565794
		), .Z(n_14896));
	notech_nand2 i_54432899(.A(n_26498), .B(n_59847), .Z(n_2234));
	notech_or4 i_175232824(.A(n_275388704), .B(n_2835), .C(n_57445), .D(n_29130
		), .Z(n_2157));
	notech_or4 i_40633110(.A(n_274988708), .B(n_275288705), .C(n_2647), .D(n_59922
		), .Z(n_55943));
	notech_ao4 i_187740415(.A(n_2345), .B(n_27538), .C(n_55808), .D(n_29231)
		, .Z(n_312565442));
	notech_and4 i_188440408(.A(n_312265439), .B(n_312065437), .C(n_288165198
		), .D(n_288465201), .Z(n_312465441));
	notech_ao4 i_188040412(.A(n_59190), .B(n_26783), .C(n_26435), .D(n_29232
		), .Z(n_312265439));
	notech_ao4 i_188240410(.A(n_55811), .B(n_310818885), .C(n_2211), .D(n_310565422
		), .Z(n_312065437));
	notech_ao4 i_188540407(.A(n_54439), .B(n_29233), .C(n_56144), .D(n_27624
		), .Z(n_311765434));
	notech_ao4 i_188640406(.A(n_54451), .B(n_27661), .C(n_56097), .D(n_27701
		), .Z(n_311665433));
	notech_and2 i_189040402(.A(n_311465431), .B(n_311365430), .Z(n_311565432
		));
	notech_ao4 i_188840404(.A(n_55924), .B(n_27388), .C(n_55910), .D(n_27733
		), .Z(n_311465431));
	notech_ao4 i_188940403(.A(n_55898), .B(n_27769), .C(n_55940), .D(n_27804
		), .Z(n_311365430));
	notech_and4 i_189840394(.A(n_311065427), .B(n_310965426), .C(n_310765424
		), .D(n_310665423), .Z(n_311265429));
	notech_ao4 i_189240400(.A(n_55879), .B(n_27836), .C(n_56049), .D(n_27870
		), .Z(n_311065427));
	notech_ao4 i_189340399(.A(n_56035), .B(n_27905), .C(n_56013), .D(n_27938
		), .Z(n_310965426));
	notech_ao4 i_189540397(.A(n_55998), .B(n_27971), .C(n_55872), .D(n_28003
		), .Z(n_310765424));
	notech_ao4 i_189640396(.A(n_55873), .B(n_29234), .C(n_55878), .D(n_28037
		), .Z(n_310665423));
	notech_nand2 i_1842258(.A(opc_10[18]), .B(n_62401), .Z(n_310565422));
	notech_and4 i_190340389(.A(n_310265419), .B(n_310065417), .C(n_290365220
		), .D(n_290665223), .Z(n_310465421));
	notech_ao4 i_189940393(.A(n_55567), .B(nbus_11273[19]), .C(n_55568), .D(\nbus_11276[19] 
		), .Z(n_310265419));
	notech_ao4 i_190140391(.A(n_2345), .B(n_27539), .C(n_55808), .D(n_29235)
		, .Z(n_310065417));
	notech_and4 i_190840384(.A(n_309765414), .B(n_309565412), .C(n_290965226
		), .D(n_291265229), .Z(n_309965416));
	notech_ao4 i_190440388(.A(n_59190), .B(n_26784), .C(n_26435), .D(n_29236
		), .Z(n_309765414));
	notech_ao4 i_190640386(.A(n_55811), .B(n_310718884), .C(n_2211), .D(n_308065397
		), .Z(n_309565412));
	notech_ao4 i_190940383(.A(n_54439), .B(n_29237), .C(n_56144), .D(n_27625
		), .Z(n_309265409));
	notech_ao4 i_191040382(.A(n_56130), .B(n_27662), .C(n_56097), .D(n_27702
		), .Z(n_309165408));
	notech_and2 i_191440378(.A(n_308965406), .B(n_308865405), .Z(n_309065407
		));
	notech_ao4 i_191240380(.A(n_54535), .B(n_27389), .C(n_55910), .D(n_27734
		), .Z(n_308965406));
	notech_ao4 i_191340379(.A(n_55898), .B(n_27770), .C(n_55940), .D(n_27805
		), .Z(n_308865405));
	notech_and4 i_192240370(.A(n_308565402), .B(n_308465401), .C(n_308265399
		), .D(n_308165398), .Z(n_308765404));
	notech_ao4 i_191640376(.A(n_55867), .B(n_27837), .C(n_56068), .D(n_27871
		), .Z(n_308565402));
	notech_ao4 i_191740375(.A(n_56035), .B(n_27906), .C(n_56013), .D(n_27939
		), .Z(n_308465401));
	notech_ao4 i_191940373(.A(n_55998), .B(n_27972), .C(n_55972), .D(n_28006
		), .Z(n_308265399));
	notech_ao4 i_192040372(.A(n_55952), .B(n_29238), .C(n_55878), .D(n_28038
		), .Z(n_308165398));
	notech_nand2 i_1942257(.A(opc_10[19]), .B(opcode_289113), .Z(n_308065397
		));
	notech_and4 i_197540317(.A(n_307765394), .B(n_307565392), .C(n_293165248
		), .D(n_293465251), .Z(n_307965396));
	notech_ao4 i_197140321(.A(n_55567), .B(nbus_11273[22]), .C(n_55568), .D(\nbus_11276[22] 
		), .Z(n_307765394));
	notech_ao4 i_197340319(.A(n_2345), .B(n_27542), .C(n_55808), .D(n_29239)
		, .Z(n_307565392));
	notech_and4 i_198040312(.A(n_307265389), .B(n_307065387), .C(n_293765254
		), .D(n_294065257), .Z(n_307465391));
	notech_ao4 i_197640316(.A(n_59190), .B(n_26788), .C(n_26435), .D(n_29240
		), .Z(n_307265389));
	notech_ao4 i_197840314(.A(n_310418881), .B(n_55811), .C(n_305565372), .D
		(n_2211), .Z(n_307065387));
	notech_ao4 i_198140311(.A(n_55873), .B(n_29241), .C(n_55864), .D(n_27737
		), .Z(n_306765384));
	notech_ao4 i_198240310(.A(n_55867), .B(n_27840), .C(n_55872), .D(n_28009
		), .Z(n_306665383));
	notech_and2 i_198640306(.A(n_306465381), .B(n_306365380), .Z(n_306565382
		));
	notech_ao4 i_198440308(.A(n_55898), .B(n_27774), .C(n_55998), .D(n_27975
		), .Z(n_306465381));
	notech_ao4 i_198540307(.A(n_56151), .B(n_27628), .C(n_55870), .D(n_27943
		), .Z(n_306365380));
	notech_and4 i_199440298(.A(n_306065377), .B(n_305965376), .C(n_305765374
		), .D(n_305665373), .Z(n_306265379));
	notech_ao4 i_198840304(.A(n_54439), .B(n_29242), .C(n_56035), .D(n_27909
		), .Z(n_306065377));
	notech_ao4 i_198940303(.A(n_54451), .B(n_27669), .C(n_56068), .D(n_27874
		), .Z(n_305965376));
	notech_ao4 i_199140301(.A(n_56097), .B(n_27705), .C(n_55878), .D(n_28041
		), .Z(n_305765374));
	notech_ao4 i_199240300(.A(n_54535), .B(n_27392), .C(n_27808), .D(n_55940
		), .Z(n_305665373));
	notech_nand2 i_2342254(.A(opc_10[22]), .B(n_62401), .Z(n_305565372));
	notech_and4 i_201440278(.A(n_304965366), .B(n_304865365), .C(n_304665363
		), .D(n_304565362), .Z(n_305165368));
	notech_ao4 i_200840284(.A(n_2261), .B(n_29241), .C(n_56240), .D(n_27737)
		, .Z(n_304965366));
	notech_ao4 i_200940283(.A(n_27840), .B(n_197114365), .C(n_56178), .D(n_28009
		), .Z(n_304865365));
	notech_ao4 i_201140281(.A(n_57343), .B(n_27774), .C(n_56414), .D(n_27975
		), .Z(n_304665363));
	notech_ao4 i_201240280(.A(n_56310), .B(n_27628), .C(n_56182), .D(n_27943
		), .Z(n_304565362));
	notech_and4 i_202140271(.A(n_304265359), .B(n_304165358), .C(n_303965356
		), .D(n_303865355), .Z(n_304465361));
	notech_ao4 i_201540277(.A(n_56183), .B(n_29242), .C(n_60484), .D(n_27909
		), .Z(n_304265359));
	notech_ao4 i_201640276(.A(n_56290), .B(n_27669), .C(n_56186), .D(n_27874
		), .Z(n_304165358));
	notech_ao4 i_201840274(.A(n_56270), .B(n_27705), .C(n_59224), .D(n_28041
		), .Z(n_303965356));
	notech_ao4 i_201940273(.A(n_57373), .B(n_27392), .C(n_2262), .D(n_27808)
		, .Z(n_303865355));
	notech_ao4 i_205640236(.A(n_29238), .B(n_2261), .C(n_56240), .D(n_27734)
		, .Z(n_303565352));
	notech_ao4 i_205740235(.A(n_2262), .B(n_27805), .C(n_27837), .D(n_197114365
		), .Z(n_303465351));
	notech_and2 i_206140231(.A(n_303265349), .B(n_303165348), .Z(n_303365350
		));
	notech_ao4 i_205940233(.A(n_28006), .B(n_56178), .C(n_57343), .D(n_27770
		), .Z(n_303265349));
	notech_ao4 i_206040232(.A(n_56414), .B(n_27972), .C(n_56310), .D(n_27625
		), .Z(n_303165348));
	notech_and4 i_206940223(.A(n_302865345), .B(n_302765344), .C(n_302565342
		), .D(n_302465341), .Z(n_303065347));
	notech_ao4 i_206340229(.A(n_27939), .B(n_56182), .C(n_56183), .D(n_29237
		), .Z(n_302865345));
	notech_ao4 i_206440228(.A(n_60484), .B(n_27906), .C(n_56290), .D(n_27662
		), .Z(n_302765344));
	notech_ao4 i_206640226(.A(n_56186), .B(n_27871), .C(n_56270), .D(n_27702
		), .Z(n_302565342));
	notech_ao4 i_206740225(.A(n_59224), .B(n_28038), .C(n_57371), .D(n_27389
		), .Z(n_302465341));
	notech_ao4 i_207240220(.A(n_29234), .B(n_2261), .C(n_56240), .D(n_27733)
		, .Z(n_302165338));
	notech_ao4 i_207340219(.A(n_2262), .B(n_27804), .C(n_27836), .D(n_197114365
		), .Z(n_302065337));
	notech_and2 i_207740215(.A(n_301865335), .B(n_301765334), .Z(n_301965336
		));
	notech_ao4 i_207540217(.A(n_28003), .B(n_56178), .C(n_57343), .D(n_27769
		), .Z(n_301865335));
	notech_ao4 i_207640216(.A(n_56414), .B(n_27971), .C(n_56310), .D(n_27624
		), .Z(n_301765334));
	notech_and4 i_208540207(.A(n_301465331), .B(n_301365330), .C(n_301165328
		), .D(n_301065327), .Z(n_301665333));
	notech_ao4 i_207940213(.A(n_27938), .B(n_56182), .C(n_56183), .D(n_29233
		), .Z(n_301465331));
	notech_ao4 i_208040212(.A(n_60484), .B(n_27905), .C(n_56290), .D(n_27661
		), .Z(n_301365330));
	notech_ao4 i_208240210(.A(n_56186), .B(n_27870), .C(n_56270), .D(n_27701
		), .Z(n_301165328));
	notech_ao4 i_208340209(.A(n_59224), .B(n_28037), .C(n_57373), .D(n_27388
		), .Z(n_301065327));
	notech_or4 i_9923(.A(n_260688757), .B(n_2605), .C(n_205088863), .D(n_55998
		), .Z(n_296165278));
	notech_or2 i_74760692(.A(n_54935), .B(n_142063758), .Z(n_296065277));
	notech_or2 i_111360667(.A(n_54935), .B(n_280965126), .Z(n_295965276));
	notech_or2 i_74860691(.A(n_260961637), .B(n_142063758), .Z(n_295865275)
		);
	notech_or2 i_111660666(.A(n_260961637), .B(n_280965126), .Z(n_295765274)
		);
	notech_or2 i_95641312(.A(n_26618), .B(n_55587), .Z(n_294065257));
	notech_or2 i_96141309(.A(n_55842), .B(n_27589), .Z(n_293765254));
	notech_or2 i_96441306(.A(n_55597), .B(n_29174), .Z(n_293465251));
	notech_or2 i_96741303(.A(n_2212), .B(nbus_11326[22]), .Z(n_293165248));
	notech_or2 i_86841396(.A(n_55587), .B(n_311218889), .Z(n_291265229));
	notech_or2 i_87141393(.A(n_55842), .B(n_27585), .Z(n_290965226));
	notech_or2 i_87441390(.A(n_55597), .B(n_29167), .Z(n_290665223));
	notech_or2 i_87741387(.A(n_2212), .B(nbus_11326[19]), .Z(n_290365220));
	notech_or2 i_83741424(.A(n_55587), .B(n_311318890), .Z(n_288465201));
	notech_or2 i_84041421(.A(n_55842), .B(n_27584), .Z(n_288165198));
	notech_or2 i_84441418(.A(n_55597), .B(n_29165), .Z(n_287865195));
	notech_or2 i_84741415(.A(n_2212), .B(nbus_11326[18]), .Z(n_287565192));
	notech_or2 i_21942023(.A(n_26618), .B(n_323365550), .Z(n_287265189));
	notech_or2 i_22242020(.A(n_323065547), .B(\nbus_11276[22] ), .Z(n_286965186
		));
	notech_nand3 i_22542017(.A(n_1416), .B(tsc[54]), .C(n_59847), .Z(n_286665183
		));
	notech_or2 i_21042032(.A(n_311018887), .B(n_323365550), .Z(n_286365180)
		);
	notech_or2 i_21342029(.A(n_323065547), .B(\nbus_11276[21] ), .Z(n_286065177
		));
	notech_nand3 i_21642026(.A(n_1416), .B(tsc[53]), .C(n_59835), .Z(n_285765174
		));
	notech_or2 i_20142041(.A(n_311118888), .B(n_323365550), .Z(n_285465171)
		);
	notech_or2 i_20642036(.A(n_328565589), .B(nbus_11326[20]), .Z(n_284965166
		));
	notech_or2 i_19242050(.A(n_311218889), .B(n_323365550), .Z(n_284565162)
		);
	notech_or2 i_19742045(.A(n_328565589), .B(nbus_11326[19]), .Z(n_284065157
		));
	notech_or2 i_18342059(.A(n_311318890), .B(n_323365550), .Z(n_283665153)
		);
	notech_or2 i_18642056(.A(n_323065547), .B(\nbus_11276[18] ), .Z(n_283365150
		));
	notech_nand3 i_18942053(.A(n_1416), .B(tsc[50]), .C(n_59835), .Z(n_283065147
		));
	notech_or2 i_6842174(.A(n_311318890), .B(n_321288477), .Z(n_282765144)
		);
	notech_or4 i_7142171(.A(n_60591), .B(n_59835), .C(n_26629), .D(n_27538),
		 .Z(n_282465141));
	notech_or2 i_7442168(.A(n_55534), .B(nbus_11273[18]), .Z(n_282165138));
	notech_and2 i_99641274(.A(n_280965126), .B(n_142063758), .Z(n_281665133)
		);
	notech_ao4 i_52360711(.A(n_56574), .B(n_204988864), .C(n_2241), .D(n_26583
		), .Z(n_280965126));
	notech_or4 i_66160695(.A(n_56574), .B(n_205088863), .C(n_56163), .D(n_56120
		), .Z(n_280865125));
	notech_ao4 i_119444224(.A(n_55131), .B(n_29214), .C(n_131123298), .D(nbus_11326
		[25]), .Z(n_280665123));
	notech_ao4 i_119544223(.A(n_55533), .B(\nbus_11276[25] ), .C(n_170914103
		), .D(n_27548), .Z(n_280465121));
	notech_and4 i_120244216(.A(n_280165118), .B(n_279965116), .C(n_245164768
		), .D(n_244864765), .Z(n_280365120));
	notech_ao4 i_119844220(.A(n_59190), .B(n_26661), .C(n_242664743), .D(n_29215
		), .Z(n_280165118));
	notech_ao4 i_120044218(.A(n_268264999), .B(n_302421911), .C(n_308421971)
		, .D(n_302221909), .Z(n_279965116));
	notech_and4 i_120744211(.A(n_54860), .B(n_279665113), .C(n_279465111), .D
		(n_245664773), .Z(n_279865115));
	notech_ao4 i_120344215(.A(n_55131), .B(n_29216), .C(n_131123298), .D(nbus_11326
		[26]), .Z(n_279665113));
	notech_ao4 i_120544213(.A(n_55533), .B(\nbus_11276[26] ), .C(n_170914103
		), .D(n_27549), .Z(n_279465111));
	notech_and4 i_121244206(.A(n_279165108), .B(n_278965106), .C(n_246264779
		), .D(n_245964776), .Z(n_279365110));
	notech_ao4 i_120844210(.A(n_59188), .B(n_26664), .C(n_242664743), .D(n_29156
		), .Z(n_279165108));
	notech_ao4 i_121044208(.A(n_288561889), .B(n_302421911), .C(n_308321970)
		, .D(n_302221909), .Z(n_278965106));
	notech_and4 i_121744201(.A(n_54860), .B(n_278665103), .C(n_278465101), .D
		(n_246764784), .Z(n_278865105));
	notech_ao4 i_121344205(.A(n_55131), .B(n_29217), .C(n_131123298), .D(nbus_11326
		[27]), .Z(n_278665103));
	notech_ao4 i_121544203(.A(n_55533), .B(\nbus_11276[27] ), .C(n_170914103
		), .D(n_27550), .Z(n_278465101));
	notech_and4 i_122244196(.A(n_278165098), .B(n_277965096), .C(n_247364790
		), .D(n_247064787), .Z(n_278365100));
	notech_ao4 i_121844200(.A(n_59188), .B(n_26673), .C(n_242664743), .D(n_29154
		), .Z(n_278165098));
	notech_ao4 i_122044198(.A(n_286061878), .B(n_302421911), .C(n_308221969)
		, .D(n_302221909), .Z(n_277965096));
	notech_ao4 i_122344195(.A(n_55131), .B(n_29218), .C(n_131423301), .D(n_27596
		), .Z(n_277765094));
	notech_ao4 i_122444194(.A(n_55534), .B(nbus_11273[28]), .C(n_55533), .D(\nbus_11276[28] 
		), .Z(n_277565092));
	notech_and4 i_123144187(.A(n_277265089), .B(n_277065087), .C(n_248164798
		), .D(n_248464801), .Z(n_277465091));
	notech_ao4 i_122744191(.A(n_59188), .B(n_26674), .C(n_57330), .D(n_242764744
		), .Z(n_277265089));
	notech_ao4 i_122944189(.A(n_343565725), .B(n_302421911), .C(n_57306), .D
		(n_302221909), .Z(n_277065087));
	notech_ao4 i_129944120(.A(n_27545), .B(n_59835), .C(n_107626780), .D(n_28721
		), .Z(n_276865085));
	notech_ao4 i_130044119(.A(n_323165548), .B(nbus_11273[23]), .C(n_323065547
		), .D(\nbus_11276[23] ), .Z(n_276665083));
	notech_and3 i_130644113(.A(n_276265079), .B(n_276465081), .C(n_249364810
		), .Z(n_276565082));
	notech_ao4 i_130344116(.A(n_322965546), .B(n_29152), .C(n_27590), .D(n_322865545
		), .Z(n_276465081));
	notech_ao4 i_130444115(.A(n_308521972), .B(n_328765591), .C(n_270765024)
		, .D(n_328665590), .Z(n_276265079));
	notech_ao4 i_130844111(.A(n_328565589), .B(nbus_11326[25]), .C(n_243064747
		), .D(\nbus_11276[25] ), .Z(n_275965076));
	notech_nand3 i_131344106(.A(n_275565072), .B(n_275765074), .C(n_250164818
		), .Z(n_275865075));
	notech_ao4 i_131044109(.A(n_2657), .B(nbus_11273[25]), .C(n_242864745), 
		.D(n_29215), .Z(n_275765074));
	notech_ao4 i_131144108(.A(n_303921926), .B(n_55867), .C(n_268264999), .D
		(n_258464901), .Z(n_275565072));
	notech_ao4 i_131544104(.A(n_328565589), .B(nbus_11326[26]), .C(n_243064747
		), .D(\nbus_11276[26] ), .Z(n_275265069));
	notech_nand3 i_132044099(.A(n_274865065), .B(n_275065067), .C(n_250964826
		), .Z(n_275165068));
	notech_ao4 i_131744102(.A(n_2657), .B(nbus_11273[26]), .C(n_242864745), 
		.D(n_29156), .Z(n_275065067));
	notech_ao4 i_131844101(.A(n_304021927), .B(n_55879), .C(n_288561889), .D
		(n_258464901), .Z(n_274865065));
	notech_ao4 i_132144098(.A(n_1031), .B(n_59926), .C(n_107626780), .D(n_28722
		), .Z(n_274665063));
	notech_ao4 i_132244097(.A(n_323165548), .B(nbus_11273[27]), .C(n_323065547
		), .D(\nbus_11276[27] ), .Z(n_274465061));
	notech_and4 i_133044090(.A(n_274165058), .B(n_273965056), .C(n_251664833
		), .D(n_251964836), .Z(n_274365060));
	notech_ao4 i_132644094(.A(n_27550), .B(n_59835), .C(n_322865545), .D(n_27595
		), .Z(n_274165058));
	notech_ao4 i_132844092(.A(n_308221969), .B(n_328765591), .C(n_286061878)
		, .D(n_328665590), .Z(n_273965056));
	notech_ao4 i_133244088(.A(nbus_11326[28]), .B(n_328565589), .C(n_243064747
		), .D(\nbus_11276[28] ), .Z(n_273665053));
	notech_nand3 i_133744083(.A(n_273265049), .B(n_273465051), .C(n_252764844
		), .Z(n_273565052));
	notech_ao4 i_133444086(.A(n_2657), .B(nbus_11273[28]), .C(n_57330), .D(n_242964746
		), .Z(n_273465051));
	notech_ao4 i_133544085(.A(n_304221929), .B(n_55879), .C(n_343565725), .D
		(n_258464901), .Z(n_273265049));
	notech_and4 i_188843545(.A(n_272965046), .B(n_272765044), .C(n_253364850
		), .D(n_253064847), .Z(n_273165048));
	notech_ao4 i_188443549(.A(n_55567), .B(nbus_11273[23]), .C(n_55568), .D(\nbus_11276[23] 
		), .Z(n_272965046));
	notech_ao4 i_188643547(.A(n_2345), .B(n_27545), .C(n_55808), .D(n_29220)
		, .Z(n_272765044));
	notech_and4 i_189343540(.A(n_272465041), .B(n_272265039), .C(n_253664853
		), .D(n_253964856), .Z(n_272665043));
	notech_ao4 i_188943544(.A(n_59190), .B(n_26789), .C(n_26435), .D(n_29221
		), .Z(n_272465041));
	notech_ao4 i_189143542(.A(n_55811), .B(n_308521972), .C(n_2211), .D(n_270765024
		), .Z(n_272265039));
	notech_ao4 i_189443539(.A(n_54439), .B(n_29222), .C(n_56151), .D(n_27629
		), .Z(n_271965036));
	notech_ao4 i_189543538(.A(n_54451), .B(n_27670), .C(n_56097), .D(n_27706
		), .Z(n_271865035));
	notech_and2 i_189943534(.A(n_271665033), .B(n_271565032), .Z(n_271765034
		));
	notech_ao4 i_189743536(.A(n_54535), .B(n_27393), .C(n_55864), .D(n_27738
		), .Z(n_271665033));
	notech_ao4 i_189843535(.A(n_55898), .B(n_27777), .C(n_55940), .D(n_27809
		), .Z(n_271565032));
	notech_and4 i_190743526(.A(n_271265029), .B(n_271165028), .C(n_270965026
		), .D(n_270865025), .Z(n_271465031));
	notech_ao4 i_190143532(.A(n_55879), .B(n_27841), .C(n_56068), .D(n_27875
		), .Z(n_271265029));
	notech_ao4 i_190243531(.A(n_56035), .B(n_27910), .C(n_55870), .D(n_27944
		), .Z(n_271165028));
	notech_ao4 i_190443529(.A(n_55998), .B(n_27976), .C(n_55872), .D(n_28010
		), .Z(n_270965026));
	notech_ao4 i_190543528(.A(n_55873), .B(n_29223), .C(n_55878), .D(n_28042
		), .Z(n_270865025));
	notech_nand2 i_2545385(.A(opc_10[23]), .B(n_62401), .Z(n_270765024));
	notech_and4 i_191243521(.A(n_270465021), .B(n_270265019), .C(n_255864875
		), .D(n_256164878), .Z(n_270665023));
	notech_ao4 i_190843525(.A(n_55567), .B(nbus_11273[25]), .C(n_55568), .D(\nbus_11276[25] 
		), .Z(n_270465021));
	notech_ao4 i_191043523(.A(n_2345), .B(n_27548), .C(n_55808), .D(n_29224)
		, .Z(n_270265019));
	notech_and4 i_191743516(.A(n_269965016), .B(n_269765014), .C(n_256464881
		), .D(n_256764884), .Z(n_270165018));
	notech_ao4 i_191343520(.A(n_59190), .B(n_26791), .C(n_26435), .D(n_29225
		), .Z(n_269965016));
	notech_ao4 i_191543518(.A(n_55811), .B(n_308421971), .C(n_2211), .D(n_268264999
		), .Z(n_269765014));
	notech_ao4 i_191843515(.A(n_54439), .B(n_29226), .C(n_56151), .D(n_27631
		), .Z(n_269465011));
	notech_ao4 i_191943514(.A(n_54451), .B(n_27672), .C(n_56097), .D(n_27708
		), .Z(n_269365010));
	notech_and2 i_192343510(.A(n_269165008), .B(n_269065007), .Z(n_269265009
		));
	notech_ao4 i_192143512(.A(n_55924), .B(n_27395), .C(n_55864), .D(n_27740
		), .Z(n_269165008));
	notech_ao4 i_192243511(.A(n_55893), .B(n_27779), .C(n_55940), .D(n_27811
		), .Z(n_269065007));
	notech_and4 i_193143502(.A(n_268765004), .B(n_268665003), .C(n_268465001
		), .D(n_268365000), .Z(n_268965006));
	notech_ao4 i_192543508(.A(n_55879), .B(n_27843), .C(n_56068), .D(n_27878
		), .Z(n_268765004));
	notech_ao4 i_192643507(.A(n_56033), .B(n_27912), .C(n_55870), .D(n_27946
		), .Z(n_268665003));
	notech_ao4 i_192843505(.A(n_55998), .B(n_27978), .C(n_55872), .D(n_28012
		), .Z(n_268465001));
	notech_ao4 i_192943504(.A(n_55873), .B(n_29227), .C(n_55878), .D(n_28044
		), .Z(n_268365000));
	notech_nand2 i_2745384(.A(opc_10[25]), .B(opcode_289113), .Z(n_268264999
		));
	notech_ao4 i_201843415(.A(n_2263), .B(n_26236), .C(n_243664753), .D(n_26317
		), .Z(n_268164998));
	notech_ao3 i_201943414(.A(n_56463), .B(n_29010), .C(instrc[118]), .Z(n_268064997
		));
	notech_ao4 i_202843405(.A(n_2261), .B(n_29228), .C(n_56240), .D(n_27743)
		, .Z(n_267764994));
	notech_ao4 i_202943404(.A(n_2262), .B(n_27814), .C(n_197114365), .D(n_27846
		), .Z(n_267664993));
	notech_and2 i_203343400(.A(n_267464991), .B(n_267364990), .Z(n_267564992
		));
	notech_ao4 i_203143402(.A(n_56178), .B(n_28015), .C(n_57343), .D(n_27782
		), .Z(n_267464991));
	notech_ao4 i_203243401(.A(n_56414), .B(n_27981), .C(n_56310), .D(n_27634
		), .Z(n_267364990));
	notech_and4 i_204143392(.A(n_267064987), .B(n_266964986), .C(n_266764984
		), .D(n_266664983), .Z(n_267264989));
	notech_ao4 i_203543398(.A(n_56182), .B(n_27949), .C(n_56183), .D(n_29229
		), .Z(n_267064987));
	notech_ao4 i_203643397(.A(n_60484), .B(n_27915), .C(n_56290), .D(n_27676
		), .Z(n_266964986));
	notech_ao4 i_203843395(.A(n_56186), .B(n_27881), .C(n_56270), .D(n_27711
		), .Z(n_266764984));
	notech_ao4 i_203943394(.A(n_59224), .B(n_28047), .C(n_57373), .D(n_27398
		), .Z(n_266664983));
	notech_ao4 i_207643357(.A(n_2261), .B(n_29227), .C(n_56240), .D(n_27740)
		, .Z(n_266364980));
	notech_ao4 i_207743356(.A(n_2262), .B(n_27811), .C(n_197114365), .D(n_27843
		), .Z(n_266264979));
	notech_and2 i_208143352(.A(n_266064977), .B(n_265964976), .Z(n_266164978
		));
	notech_ao4 i_207943354(.A(n_56178), .B(n_28012), .C(n_57343), .D(n_27779
		), .Z(n_266064977));
	notech_ao4 i_208043353(.A(n_56414), .B(n_27978), .C(n_56310), .D(n_27631
		), .Z(n_265964976));
	notech_and4 i_208943344(.A(n_265664973), .B(n_265564972), .C(n_265364970
		), .D(n_265264969), .Z(n_265864975));
	notech_ao4 i_208343350(.A(n_56182), .B(n_27946), .C(n_56183), .D(n_29226
		), .Z(n_265664973));
	notech_ao4 i_208443349(.A(n_60484), .B(n_27912), .C(n_56290), .D(n_27672
		), .Z(n_265564972));
	notech_ao4 i_208643347(.A(n_56186), .B(n_27878), .C(n_56270), .D(n_27708
		), .Z(n_265364970));
	notech_ao4 i_208743346(.A(n_59224), .B(n_28044), .C(n_57373), .D(n_27395
		), .Z(n_265264969));
	notech_ao4 i_209243341(.A(n_2261), .B(n_29223), .C(n_56240), .D(n_27738)
		, .Z(n_264964966));
	notech_ao4 i_209343340(.A(n_2262), .B(n_27809), .C(n_197114365), .D(n_27841
		), .Z(n_264864965));
	notech_and2 i_209743336(.A(n_264664963), .B(n_264564962), .Z(n_264764964
		));
	notech_ao4 i_209543338(.A(n_56178), .B(n_28010), .C(n_57343), .D(n_27777
		), .Z(n_264664963));
	notech_ao4 i_209643337(.A(n_56415), .B(n_27976), .C(n_56310), .D(n_27629
		), .Z(n_264564962));
	notech_and4 i_210543328(.A(n_264264959), .B(n_264164958), .C(n_263964956
		), .D(n_263864955), .Z(n_264464961));
	notech_ao4 i_209943334(.A(n_56182), .B(n_27944), .C(n_56183), .D(n_29222
		), .Z(n_264264959));
	notech_ao4 i_210043333(.A(n_60484), .B(n_27910), .C(n_56290), .D(n_27670
		), .Z(n_264164958));
	notech_ao4 i_210243331(.A(n_56186), .B(n_27875), .C(n_56270), .D(n_27706
		), .Z(n_263964956));
	notech_ao4 i_210343330(.A(n_59224), .B(n_28042), .C(n_57371), .D(n_27393
		), .Z(n_263864955));
	notech_nand3 i_31400(.A(n_56492), .B(n_268064997), .C(n_62401), .Z(n_258764904
		));
	notech_ao4 i_5245325(.A(n_56502), .B(n_56112), .C(n_56063), .D(n_26512),
		 .Z(n_258664903));
	notech_or2 i_5345324(.A(n_2689), .B(n_242364742), .Z(n_258464901));
	notech_or2 i_90744490(.A(n_55587), .B(n_308821975), .Z(n_256764884));
	notech_or2 i_91144487(.A(n_55842), .B(n_27593), .Z(n_256464881));
	notech_or2 i_91444484(.A(n_55597), .B(n_29215), .Z(n_256164878));
	notech_or2 i_91744481(.A(n_2212), .B(nbus_11326[25]), .Z(n_255864875));
	notech_or2 i_87544518(.A(n_55587), .B(n_308921976), .Z(n_253964856));
	notech_or2 i_87844515(.A(n_55842), .B(n_27590), .Z(n_253664853));
	notech_or2 i_88144512(.A(n_55597), .B(n_29152), .Z(n_253364850));
	notech_or2 i_88444509(.A(n_2212), .B(nbus_11326[23]), .Z(n_253064847));
	notech_or2 i_27145107(.A(n_242864745), .B(n_29219), .Z(n_252764844));
	notech_and3 i_27645102(.A(n_54128), .B(tsc[60]), .C(n_59835), .Z(n_252064837
		));
	notech_or2 i_26145117(.A(n_308621973), .B(n_323365550), .Z(n_251964836)
		);
	notech_or2 i_26445114(.A(n_322965546), .B(n_29154), .Z(n_251664833));
	notech_or2 i_26745111(.A(n_328565589), .B(nbus_11326[27]), .Z(n_251364830
		));
	notech_or2 i_25345125(.A(n_308721974), .B(n_242964746), .Z(n_250964826)
		);
	notech_and3 i_25845120(.A(n_54128), .B(tsc[58]), .C(n_59835), .Z(n_250264819
		));
	notech_or2 i_24545133(.A(n_308821975), .B(n_242964746), .Z(n_250164818)
		);
	notech_and3 i_25045128(.A(n_54128), .B(tsc[57]), .C(n_59835), .Z(n_249464811
		));
	notech_or2 i_23545142(.A(n_308921976), .B(n_323365550), .Z(n_249364810)
		);
	notech_or2 i_24145137(.A(n_328565589), .B(nbus_11326[23]), .Z(n_248864805
		));
	notech_or2 i_15245225(.A(n_242664743), .B(n_29219), .Z(n_248464801));
	notech_or4 i_15545222(.A(n_60591), .B(n_59835), .C(n_26629), .D(n_27551)
		, .Z(n_248164798));
	notech_nao3 i_15845219(.A(n_26549), .B(opc[28]), .C(n_316988520), .Z(n_247864795
		));
	notech_or2 i_14145236(.A(n_308621973), .B(n_242764744), .Z(n_247364790)
		);
	notech_or4 i_14445233(.A(n_56376), .B(n_55924), .C(n_60591), .D(n_27595)
		, .Z(n_247064787));
	notech_or2 i_14745230(.A(n_55534), .B(nbus_11273[27]), .Z(n_246764784)
		);
	notech_or2 i_13045247(.A(n_308721974), .B(n_242764744), .Z(n_246264779)
		);
	notech_or4 i_13345244(.A(n_56375), .B(n_55924), .C(n_60591), .D(n_27594)
		, .Z(n_245964776));
	notech_or2 i_13645241(.A(n_55534), .B(nbus_11273[26]), .Z(n_245664773)
		);
	notech_or2 i_11945258(.A(n_308821975), .B(n_242764744), .Z(n_245164768)
		);
	notech_or4 i_12245255(.A(n_56375), .B(n_55924), .C(n_60591), .D(n_27593)
		, .Z(n_244864765));
	notech_or2 i_12545252(.A(n_55534), .B(nbus_11273[25]), .Z(n_244564762)
		);
	notech_nao3 i_24045381(.A(n_56463), .B(n_56492), .C(n_114626850), .Z(n_243964756
		));
	notech_or2 i_103044379(.A(n_55859), .B(n_26512), .Z(n_243864755));
	notech_ao4 i_102944380(.A(n_59380), .B(n_62401), .C(n_2264), .D(n_26236)
		, .Z(n_243664753));
	notech_and3 i_88663596(.A(n_54642), .B(n_54762), .C(n_328165585), .Z(n_243064747
		));
	notech_and2 i_102145415(.A(n_2661), .B(n_241764736), .Z(n_242964746));
	notech_and2 i_101945414(.A(n_2659), .B(n_241864737), .Z(n_242864745));
	notech_ao4 i_105945417(.A(n_215558439), .B(n_320888481), .C(n_26326), .D
		(n_54874), .Z(n_242764744));
	notech_and2 i_105845416(.A(n_55459), .B(n_55978), .Z(n_242664743));
	notech_and2 i_3345344(.A(n_2660), .B(n_120563543), .Z(n_242364742));
	notech_and4 i_2445349(.A(n_55976), .B(n_258664903), .C(n_56061), .D(n_243864755
		), .Z(n_242164740));
	notech_or2 i_81163598(.A(n_2658), .B(n_120563543), .Z(n_241864737));
	notech_or4 i_81263597(.A(n_2740), .B(n_1076), .C(n_120563543), .D(n_60530
		), .Z(n_241764736));
	notech_and4 i_210947155(.A(n_101523002), .B(n_241264731), .C(n_228964612
		), .D(n_228864611), .Z(n_241564734));
	notech_and4 i_210647158(.A(n_240964728), .B(n_228564608), .C(n_228664609
		), .D(n_228764610), .Z(n_241264731));
	notech_ao4 i_210347161(.A(n_107626780), .B(n_28712), .C(n_351165800), .D
		(n_27599), .Z(n_240964728));
	notech_and4 i_199647262(.A(n_240464723), .B(n_228064603), .C(n_227964602
		), .D(n_26207), .Z(n_240764726));
	notech_and4 i_199347265(.A(n_240164720), .B(n_227664599), .C(n_227764600
		), .D(n_227864601), .Z(n_240464723));
	notech_ao4 i_199047268(.A(n_56033), .B(n_102623013), .C(n_107626780), .D
		(n_28713), .Z(n_240164720));
	notech_and4 i_126947963(.A(n_239664715), .B(n_239564714), .C(n_239364712
		), .D(n_239264711), .Z(n_239864717));
	notech_ao4 i_126647966(.A(n_59188), .B(n_26683), .C(n_55534), .D(nbus_11273
		[31]), .Z(n_239664715));
	notech_ao4 i_126547967(.A(n_131423301), .B(n_27601), .C(n_170914103), .D
		(n_27554), .Z(n_239564714));
	notech_ao4 i_126447968(.A(n_242664743), .B(n_28996), .C(n_55533), .D(\nbus_11276[31] 
		), .Z(n_239364712));
	notech_ao4 i_126347969(.A(n_131123298), .B(nbus_11326[31]), .C(n_55131),
		 .D(n_29213), .Z(n_239264711));
	notech_and4 i_119848031(.A(n_238764706), .B(n_238664705), .C(n_238564704
		), .D(n_226064583), .Z(n_239064709));
	notech_ao4 i_119448035(.A(n_262936784), .B(n_55879), .C(n_242864745), .D
		(n_28977), .Z(n_238764706));
	notech_ao4 i_119348036(.A(n_242964746), .B(n_57329), .C(n_243064747), .D
		(\nbus_11276[29] ), .Z(n_238664705));
	notech_and3 i_119548034(.A(n_262736782), .B(n_225464577), .C(n_225964582
		), .Z(n_238564704));
	notech_nand3 i_117948050(.A(n_237964698), .B(n_224964572), .C(n_225064573
		), .Z(n_238164700));
	notech_and4 i_117748052(.A(n_55901), .B(n_237764696), .C(n_237564694), .D
		(n_224464567), .Z(n_237964698));
	notech_ao4 i_117448055(.A(n_322965546), .B(n_28997), .C(n_323065547), .D
		(\nbus_11276[30] ), .Z(n_237764696));
	notech_ao4 i_117548054(.A(n_323165548), .B(nbus_11273[30]), .C(n_322865545
		), .D(n_27599), .Z(n_237564694));
	notech_nand3 i_116148068(.A(n_237164690), .B(n_224164564), .C(n_224064563
		), .Z(n_237364692));
	notech_and4 i_115948070(.A(n_236864687), .B(n_236764686), .C(n_223864561
		), .D(n_223964562), .Z(n_237164690));
	notech_ao4 i_115648073(.A(n_2657), .B(nbus_11273[31]), .C(n_28996), .D(n_242864745
		), .Z(n_236864687));
	notech_ao4 i_115548074(.A(n_243064747), .B(\nbus_11276[31] ), .C(n_328565589
		), .D(nbus_11326[31]), .Z(n_236764686));
	notech_and4 i_114348086(.A(n_236364682), .B(n_236264681), .C(n_236064679
		), .D(n_235964678), .Z(n_236564684));
	notech_ao4 i_114048089(.A(n_55220), .B(nbus_11273[29]), .C(n_262936784),
		 .D(n_55893), .Z(n_236364682));
	notech_ao4 i_113948090(.A(n_55347), .B(n_28977), .C(n_55346), .D(n_57329
		), .Z(n_236264681));
	notech_ao4 i_113848091(.A(n_55221), .B(\nbus_11276[29] ), .C(n_303421921
		), .D(nbus_11326[29]), .Z(n_236064679));
	notech_and2 i_113748092(.A(n_55901), .B(n_262736782), .Z(n_235964678));
	notech_and4 i_112448104(.A(n_235364672), .B(n_235264671), .C(n_235164670
		), .D(n_221864546), .Z(n_235664675));
	notech_ao4 i_112048108(.A(n_55557), .B(n_28997), .C(n_55221), .D(\nbus_11276[30] 
		), .Z(n_235364672));
	notech_ao4 i_111948109(.A(n_1031), .B(n_59926), .C(n_303421921), .D(nbus_11326
		[30]), .Z(n_235264671));
	notech_ao4 i_112148107(.A(n_55220), .B(nbus_11273[30]), .C(n_55772), .D(n_27599
		), .Z(n_235164670));
	notech_and4 i_98848228(.A(n_234164660), .B(n_234064659), .C(n_220964538)
		, .D(n_234664665), .Z(n_234864667));
	notech_and3 i_98648230(.A(n_234464663), .B(n_234364662), .C(n_220864537)
		, .Z(n_234664665));
	notech_ao4 i_98048236(.A(n_55977), .B(n_28444), .C(n_262636781), .D(n_26985
		), .Z(n_234464663));
	notech_ao4 i_98348233(.A(n_55536), .B(nbus_11273[30]), .C(n_55135), .D(n_27599
		), .Z(n_234364662));
	notech_ao4 i_98248234(.A(n_262536780), .B(n_27553), .C(n_55535), .D(\nbus_11276[30] 
		), .Z(n_234164660));
	notech_ao4 i_98148235(.A(n_308518862), .B(nbus_11326[30]), .C(n_56024), 
		.D(n_29212), .Z(n_234064659));
	notech_and4 i_57148618(.A(n_233464653), .B(n_233264652), .C(n_224964572)
		, .D(n_219564525), .Z(n_233764656));
	notech_ao4 i_56748622(.A(n_26572), .B(\nbus_11276[30] ), .C(n_121623203)
		, .D(nbus_11326[30]), .Z(n_233464653));
	notech_ao4 i_56848621(.A(n_353465823), .B(n_27599), .C(n_353165820), .D(n_28997
		), .Z(n_233264652));
	notech_and4 i_68249178(.A(n_232864649), .B(n_218764518), .C(n_218864519)
		, .D(n_218564516), .Z(n_101523002));
	notech_ao4 i_44948729(.A(n_59835), .B(n_27553), .C(n_56057), .D(\nbus_11276[30] 
		), .Z(n_232864649));
	notech_nand3 i_41748761(.A(n_231864640), .B(n_231664639), .C(n_232364645
		), .Z(n_232464646));
	notech_and3 i_41648762(.A(n_232164643), .B(n_232064642), .C(n_218264513)
		, .Z(n_232364645));
	notech_ao4 i_41048768(.A(n_55568), .B(\nbus_11276[29] ), .C(n_2212), .D(nbus_11326
		[29]), .Z(n_232164643));
	notech_ao4 i_41348765(.A(n_55567), .B(nbus_11273[29]), .C(n_55842), .D(n_27597
		), .Z(n_232064642));
	notech_ao4 i_41248766(.A(n_55808), .B(n_29211), .C(n_2345), .D(n_27552),
		 .Z(n_231864640));
	notech_ao4 i_41148767(.A(n_55597), .B(n_28977), .C(n_55587), .D(n_57329)
		, .Z(n_231664639));
	notech_nand2 i_39148784(.A(n_231264635), .B(n_216864501), .Z(n_231364636
		));
	notech_and4 i_39048785(.A(n_231064633), .B(n_230964632), .C(n_230764630)
		, .D(n_230664629), .Z(n_231264635));
	notech_ao4 i_38748788(.A(n_59190), .B(n_26796), .C(n_55567), .D(nbus_11273
		[30]), .Z(n_231064633));
	notech_ao4 i_38648789(.A(n_55842), .B(n_27599), .C(n_55808), .D(n_29210)
		, .Z(n_230964632));
	notech_ao4 i_38548790(.A(n_2345), .B(n_27553), .C(n_55597), .D(n_28997),
		 .Z(n_230764630));
	notech_ao4 i_38448791(.A(n_55568), .B(\nbus_11276[30] ), .C(n_2212), .D(nbus_11326
		[30]), .Z(n_230664629));
	notech_nand2 i_33648837(.A(n_230264625), .B(n_215564489), .Z(n_230364626
		));
	notech_and4 i_33548838(.A(n_230064623), .B(n_229964622), .C(n_229764620)
		, .D(n_229664619), .Z(n_230264625));
	notech_ao4 i_33248841(.A(n_59190), .B(n_26797), .C(n_55567), .D(nbus_11273
		[31]), .Z(n_230064623));
	notech_ao4 i_33148842(.A(n_55842), .B(n_27601), .C(n_55808), .D(n_29209)
		, .Z(n_229964622));
	notech_ao4 i_33048843(.A(n_2345), .B(n_27554), .C(n_55597), .D(n_28996),
		 .Z(n_229764620));
	notech_ao4 i_32948844(.A(n_55568), .B(\nbus_11276[31] ), .C(n_2212), .D(nbus_11326
		[31]), .Z(n_229664619));
	notech_nand3 i_87749175(.A(n_56060), .B(n_213264466), .C(n_351465803), .Z
		(n_229564618));
	notech_ao4 i_16149003(.A(n_62427), .B(\opcode[1] ), .C(n_2263), .D(n_26237
		), .Z(n_229464617));
	notech_or2 i_15549007(.A(n_56492), .B(n_56463), .Z(n_229364616));
	notech_ao4 i_9349069(.A(n_28442003), .B(n_27331), .C(n_27341992), .D(n_27364
		), .Z(n_229164614));
	notech_nand3 i_3117257(.A(n_241564734), .B(n_229064613), .C(n_228264605)
		, .Z(n_15954));
	notech_or2 i_209947165(.A(n_351865807), .B(n_270988746), .Z(n_229064613)
		);
	notech_or2 i_209747167(.A(n_55143), .B(nbus_11273[30]), .Z(n_228964612)
		);
	notech_or2 i_209847166(.A(n_55142), .B(\nbus_11276[30] ), .Z(n_228864611
		));
	notech_nao3 i_210247162(.A(opc_10[30]), .B(opcode_289113), .C(n_352865817
		), .Z(n_228764610));
	notech_or4 i_210047164(.A(n_58661), .B(n_56120), .C(n_55523), .D(n_271188744
		), .Z(n_228664609));
	notech_or2 i_209547169(.A(n_351665805), .B(nbus_11326[30]), .Z(n_228564608
		));
	notech_or2 i_209647168(.A(n_351765806), .B(n_28997), .Z(n_228264605));
	notech_nand3 i_3217258(.A(n_240764726), .B(n_228164604), .C(n_227364596)
		, .Z(n_15960));
	notech_or2 i_198447273(.A(n_352165810), .B(n_271088745), .Z(n_228164604)
		);
	notech_or2 i_198247275(.A(n_55143), .B(nbus_11273[31]), .Z(n_228064603)
		);
	notech_or2 i_198347274(.A(n_55142), .B(\nbus_11276[31] ), .Z(n_227964602
		));
	notech_nao3 i_198947269(.A(opc_10[31]), .B(opcode_289113), .C(n_352965818
		), .Z(n_227864601));
	notech_or4 i_198547272(.A(n_58660), .B(n_56120), .C(n_55798), .D(n_271288743
		), .Z(n_227764600));
	notech_nand2 i_198047277(.A(n_351965808), .B(opc[31]), .Z(n_227664599)
		);
	notech_nand2 i_198147276(.A(n_352065809), .B(\regs_13_14[31] ), .Z(n_227364596
		));
	notech_or4 i_3216681(.A(n_227164594), .B(n_227264595), .C(n_226264585), 
		.D(n_26300), .Z(n_11878));
	notech_nor2 i_126147971(.A(n_302221909), .B(n_271288743), .Z(n_227264595
		));
	notech_ao3 i_126247970(.A(opc_10[31]), .B(n_62401), .C(n_302421911), .Z(n_227164594
		));
	notech_nor2 i_126047972(.A(n_242764744), .B(n_271088745), .Z(n_226264585
		));
	notech_nand3 i_3021929(.A(n_239064709), .B(n_225364576), .C(n_226164584)
		, .Z(n_12223));
	notech_nao3 i_119048039(.A(opc_10[29]), .B(n_62417), .C(n_258464901), .Z
		(n_226164584));
	notech_nand3 i_119148038(.A(n_54128), .B(tsc[61]), .C(n_59847), .Z(n_226064583
		));
	notech_or2 i_118848041(.A(n_2657), .B(nbus_11273[29]), .Z(n_225964582)
		);
	notech_or2 i_118348046(.A(n_328565589), .B(nbus_11326[29]), .Z(n_225464577
		));
	notech_or4 i_118948040(.A(n_56086), .B(n_56120), .C(n_54367), .D(n_270688747
		), .Z(n_225364576));
	notech_or4 i_3121930(.A(n_225164574), .B(n_238164700), .C(n_225264575), 
		.D(n_224364566), .Z(n_12229));
	notech_nor2 i_117048059(.A(n_328765591), .B(n_271188744), .Z(n_225264575
		));
	notech_ao3 i_117148058(.A(opc_10[30]), .B(n_62411), .C(n_328665590), .Z(n_225164574
		));
	notech_nand3 i_117248057(.A(n_54128), .B(tsc[62]), .C(n_59845), .Z(n_225064573
		));
	notech_nand2 i_165349161(.A(n_59926), .B(read_data[30]), .Z(n_224964572)
		);
	notech_or2 i_116448065(.A(n_328565589), .B(nbus_11326[30]), .Z(n_224464567
		));
	notech_nor2 i_116948060(.A(n_323365550), .B(n_270988746), .Z(n_224364566
		));
	notech_or4 i_3221931(.A(n_284968648), .B(n_297468773), .C(n_224264565), 
		.D(n_237364692), .Z(n_12235));
	notech_nor2 i_115048079(.A(n_242964746), .B(n_271088745), .Z(n_224264565
		));
	notech_or4 i_115148078(.A(n_56086), .B(n_56120), .C(n_54367), .D(n_271288743
		), .Z(n_224164564));
	notech_nao3 i_115248077(.A(opc_10[31]), .B(n_62399), .C(n_258464901), .Z
		(n_224064563));
	notech_nand3 i_115348076(.A(n_54128), .B(tsc[63]), .C(n_59845), .Z(n_223964562
		));
	notech_or4 i_115448075(.A(instrc[115]), .B(instrc[112]), .C(n_56086), .D
		(n_102623013), .Z(n_223864561));
	notech_nao3 i_3021865(.A(n_236564684), .B(n_222164549), .C(n_223164556),
		 .Z(n_12575));
	notech_ao3 i_113648093(.A(opc_10[29]), .B(n_62405), .C(n_302621913), .Z(n_223164556
		));
	notech_or4 i_113548094(.A(n_56081), .B(n_206288851), .C(n_54367), .D(n_270688747
		), .Z(n_222164549));
	notech_and4 i_3121866(.A(n_235664675), .B(n_101523002), .C(n_221964547),
		 .D(n_222064548), .Z(n_12581));
	notech_or2 i_111648112(.A(n_55556), .B(n_270988746), .Z(n_222064548));
	notech_or4 i_111748111(.A(n_56081), .B(n_206288851), .C(n_55523), .D(n_271188744
		), .Z(n_221964547));
	notech_nao3 i_111848110(.A(opc_10[30]), .B(n_62405), .C(n_322931616), .Z
		(n_221864546));
	notech_or4 i_3121738(.A(n_221064539), .B(n_221264540), .C(n_219864528), 
		.D(n_26301), .Z(n_12947));
	notech_nor2 i_97848238(.A(n_271188744), .B(n_110123088), .Z(n_221264540)
		);
	notech_nor2 i_97648240(.A(n_354688262), .B(n_28997), .Z(n_221064539));
	notech_nao3 i_97948237(.A(opc_10[30]), .B(n_62399), .C(n_110323090), .Z(n_220964538
		));
	notech_nand2 i_97548241(.A(sav_esp[30]), .B(n_60595), .Z(n_220864537));
	notech_nor2 i_97748239(.A(n_270988746), .B(n_354588263), .Z(n_219864528)
		);
	notech_or4 i_3120970(.A(n_219664526), .B(n_219764527), .C(n_218964520), 
		.D(n_26302), .Z(n_9159));
	notech_nor2 i_56548624(.A(n_271188744), .B(n_121523202), .Z(n_219764527)
		);
	notech_ao3 i_56648623(.A(opc_10[30]), .B(n_62399), .C(n_121723204), .Z(n_219664526
		));
	notech_or2 i_56348626(.A(n_353265821), .B(nbus_11273[30]), .Z(n_219564525
		));
	notech_nor2 i_56448625(.A(n_353365822), .B(n_270988746), .Z(n_218964520)
		);
	notech_or4 i_44748731(.A(n_60775), .B(n_60729), .C(n_54761), .D(n_28997)
		, .Z(n_218864519));
	notech_or2 i_44648732(.A(n_98113375), .B(nbus_11273[30]), .Z(n_218764518
		));
	notech_or2 i_44848730(.A(n_101213406), .B(n_270988746), .Z(n_218564516)
		);
	notech_or4 i_3020649(.A(n_218464515), .B(n_218364514), .C(n_232464646), 
		.D(n_217164504), .Z(n_20285));
	notech_ao3 i_40948769(.A(opc_10[29]), .B(n_62405), .C(n_2211), .Z(n_218464515
		));
	notech_and2 i_40848770(.A(n_352465813), .B(n_55819), .Z(n_218364514));
	notech_nand2 i_40648772(.A(sav_epc[29]), .B(n_60595), .Z(n_218264513));
	notech_nor2 i_40748771(.A(n_55811), .B(n_270688747), .Z(n_217164504));
	notech_or4 i_3120650(.A(n_216964502), .B(n_231364636), .C(n_217064503), 
		.D(n_215964492), .Z(n_20291));
	notech_nor2 i_38248793(.A(n_55811), .B(n_271188744), .Z(n_217064503));
	notech_ao3 i_38348792(.A(opc_10[30]), .B(n_62399), .C(n_2211), .Z(n_216964502
		));
	notech_nand2 i_38048795(.A(n_352565814), .B(n_55819), .Z(n_216864501));
	notech_nor2 i_38148794(.A(n_55587), .B(n_270988746), .Z(n_215964492));
	notech_or4 i_3220651(.A(n_215664490), .B(n_230364626), .C(n_215864491), 
		.D(n_214664480), .Z(n_20297));
	notech_nor2 i_32748846(.A(n_55811), .B(n_271288743), .Z(n_215864491));
	notech_ao3 i_32848845(.A(opc_10[31]), .B(n_62405), .C(n_2211), .Z(n_215664490
		));
	notech_nand2 i_32548848(.A(\add_len_pc[31] ), .B(n_55819), .Z(n_215564489
		));
	notech_nor2 i_32648847(.A(n_55587), .B(n_271088745), .Z(n_214664480));
	notech_mux2 i_3211689(.S(n_60136), .A(regs_14[31]), .B(add_len_pc32[31])
		, .Z(\add_len_pc[31] ));
	notech_nor2 i_22848936(.A(n_229564618), .B(n_26248), .Z(n_213964473));
	notech_and3 i_22748937(.A(n_56061), .B(n_338165683), .C(n_212664460), .Z
		(n_213864472));
	notech_nand2 i_80949232(.A(n_229564618), .B(n_54904), .Z(n_213764471));
	notech_or4 i_17148993(.A(n_114626850), .B(n_229364616), .C(n_60511), .D(n_351065799
		), .Z(n_213564469));
	notech_or4 i_74149252(.A(n_212964463), .B(n_60530), .C(n_2739), .D(n_338165683
		), .Z(n_213464468));
	notech_or2 i_74049253(.A(n_351565804), .B(n_338165683), .Z(n_213364467)
		);
	notech_or2 i_16548999(.A(n_56063), .B(n_26501), .Z(n_213264466));
	notech_ao4 i_83749174(.A(n_59380), .B(n_62413), .C(n_2264), .D(n_26237),
		 .Z(n_212964463));
	notech_and2 i_16049004(.A(n_60484), .B(n_26238), .Z(n_212864462));
	notech_or2 i_14049022(.A(n_55859), .B(n_26501), .Z(n_212664460));
	notech_nand3 i_3117833(.A(n_229164614), .B(n_212164455), .C(n_212464458)
		, .Z(write_data_26[30]));
	notech_nand3 i_9149071(.A(n_60530), .B(n_26772), .C(temp_sp[30]), .Z(n_212464458
		));
	notech_or2 i_9249070(.A(n_26595), .B(n_270988746), .Z(n_212164455));
	notech_and4 i_128850750(.A(n_211064445), .B(n_210964444), .C(n_211764451
		), .D(n_16825881), .Z(n_211964453));
	notech_and3 i_128650752(.A(n_211564449), .B(n_211464448), .C(n_211264447
		), .Z(n_211764451));
	notech_ao4 i_128050758(.A(n_295765274), .B(n_2699), .C(n_56024), .D(n_29208
		), .Z(n_211564449));
	notech_ao4 i_127950759(.A(n_55977), .B(n_28414), .C(n_262636781), .D(n_26923
		), .Z(n_211464448));
	notech_ao4 i_128350755(.A(n_59190), .B(n_26685), .C(n_262536780), .D(n_27519
		), .Z(n_211264447));
	notech_ao4 i_128250756(.A(n_208364418), .B(n_27561), .C(n_208164416), .D
		(\nbus_11276[0] ), .Z(n_211064445));
	notech_ao4 i_128150757(.A(n_208264417), .B(nbus_11273[0]), .C(n_295965276
		), .D(n_28986), .Z(n_210964444));
	notech_ao4 i_128950749(.A(n_43626149), .B(n_206764402), .C(n_206664401),
		 .D(n_46226175), .Z(n_210864443));
	notech_and4 i_68351324(.A(n_206064395), .B(n_205964394), .C(n_210364438)
		, .D(n_206364398), .Z(n_210664441));
	notech_and3 i_67951328(.A(n_210164436), .B(n_210064435), .C(n_205864393)
		, .Z(n_210364438));
	notech_ao4 i_67651331(.A(n_55808), .B(n_29207), .C(n_2345), .D(n_27524),
		 .Z(n_210164436));
	notech_ao4 i_67751330(.A(n_322788463), .B(n_55216), .C(n_55236), .D(n_29065
		), .Z(n_210064435));
	notech_ao4 i_68251325(.A(\nbus_11276[5] ), .B(n_2691), .C(n_2690), .D(n_27566
		), .Z(n_209964434));
	notech_ao4 i_68451323(.A(n_351365802), .B(n_55426267), .C(n_55687), .D(n_57321
		), .Z(n_209864433));
	notech_ao4 i_44851539(.A(n_58487), .B(n_28024), .C(n_55952), .D(n_29118)
		, .Z(n_209564430));
	notech_ao4 i_44751540(.A(n_55972), .B(n_27990), .C(n_55998), .D(n_27958)
		, .Z(n_209464429));
	notech_and2 i_45151536(.A(n_209264427), .B(n_209164426), .Z(n_209364428)
		);
	notech_ao4 i_44651541(.A(n_56013), .B(n_27924), .C(n_56033), .D(n_27891)
		, .Z(n_209264427));
	notech_ao4 i_44551542(.A(n_56049), .B(n_27855), .C(n_55867), .D(n_27823)
		, .Z(n_209164426));
	notech_and4 i_45351534(.A(n_208864423), .B(n_208764422), .C(n_208564420)
		, .D(n_208464419), .Z(n_209064425));
	notech_ao4 i_44451543(.A(n_55940), .B(n_27791), .C(n_55893), .D(n_27752)
		, .Z(n_208864423));
	notech_ao4 i_44351544(.A(n_55910), .B(n_27720), .C(n_55924), .D(n_27375)
		, .Z(n_208764422));
	notech_ao4 i_44251545(.A(n_56097), .B(n_27688), .C(n_56130), .D(n_27644)
		, .Z(n_208564420));
	notech_ao4 i_44151546(.A(n_56151), .B(n_27611), .C(n_56386), .D(n_29119)
		, .Z(n_208464419));
	notech_and3 i_61560700(.A(n_55135), .B(n_296165278), .C(n_320465521), .Z
		(n_208364418));
	notech_and2 i_85060689(.A(n_54759), .B(n_296065277), .Z(n_208264417));
	notech_and3 i_98060673(.A(n_55692), .B(n_295865275), .C(n_54751), .Z(n_208164416
		));
	notech_nand3 i_121708(.A(n_208064415), .B(n_211964453), .C(n_210864443),
		 .Z(n_12767));
	notech_or4 i_127650762(.A(n_56574), .B(n_205088863), .C(n_55998), .D(n_2688
		), .Z(n_208064415));
	notech_or4 i_120760576(.A(n_56463), .B(n_264436799), .C(n_280965126), .D
		(instrc[119]), .Z(n_206764402));
	notech_or4 i_119060577(.A(n_56463), .B(n_264436799), .C(n_142363761), .D
		(instrc[119]), .Z(n_206664401));
	notech_nand3 i_620625(.A(n_209964434), .B(n_209864433), .C(n_210664441),
		 .Z(n_20141));
	notech_nand2 i_67351334(.A(n_2692), .B(opa[5]), .Z(n_206364398));
	notech_nao3 i_67551332(.A(opc_10[5]), .B(n_62413), .C(n_54526258), .Z(n_206064395
		));
	notech_nand2 i_67051337(.A(\add_len_pc[5] ), .B(n_55819), .Z(n_205964394
		));
	notech_nand2 i_66751339(.A(sav_epc[5]), .B(n_60595), .Z(n_205864393));
	notech_mux2 i_611663(.S(n_60136), .A(n_561), .B(add_len_pc32[5]), .Z(\add_len_pc[5] 
		));
	notech_and4 i_142852031(.A(n_209564430), .B(n_209464429), .C(n_209064425
		), .D(n_209364428), .Z(n_57321));
	notech_nand2 i_123954107(.A(n_203264367), .B(n_178564123), .Z(n_203364368
		));
	notech_ao4 i_123854108(.A(n_29080), .B(n_350865797), .C(n_57347), .D(n_350965798
		), .Z(n_203264367));
	notech_and4 i_124554101(.A(n_202964364), .B(n_179164129), .C(n_202764362
		), .D(n_178864126), .Z(n_203164366));
	notech_ao4 i_124154105(.A(nbus_11273[11]), .B(n_26244), .C(n_337665678),
		 .D(n_27576), .Z(n_202964364));
	notech_ao4 i_124354103(.A(n_336065662), .B(n_171658004), .C(n_56033), .D
		(n_238768192), .Z(n_202764362));
	notech_nand2 i_124854098(.A(n_202364358), .B(n_179564133), .Z(n_202464359
		));
	notech_ao4 i_124754099(.A(n_350865797), .B(n_29084), .C(n_57346), .D(n_350965798
		), .Z(n_202364358));
	notech_and4 i_125454092(.A(n_202064355), .B(n_180164139), .C(n_201864353
		), .D(n_179864136), .Z(n_202264357));
	notech_ao4 i_125054096(.A(nbus_11273[12]), .B(n_26244), .C(n_337665678),
		 .D(n_27577), .Z(n_202064355));
	notech_ao4 i_125254094(.A(n_169057978), .B(n_336065662), .C(n_189074758)
		, .D(n_56033), .Z(n_201864353));
	notech_and4 i_125854088(.A(n_201464349), .B(n_26408), .C(n_180264140), .D
		(n_180564143), .Z(n_201764352));
	notech_ao4 i_125654090(.A(n_350865797), .B(n_29037), .C(n_57345), .D(n_350965798
		), .Z(n_201464349));
	notech_and4 i_126354083(.A(n_201164346), .B(n_181264149), .C(n_200964344
		), .D(n_180864146), .Z(n_201364348));
	notech_ao4 i_125954087(.A(nbus_11273[13]), .B(n_26244), .C(n_337665678),
		 .D(n_27578), .Z(n_201164346));
	notech_ao4 i_126154085(.A(n_336065662), .B(n_166457952), .C(n_56033), .D
		(n_187874746), .Z(n_200964344));
	notech_and4 i_134154007(.A(n_154070859), .B(n_55901), .C(n_200564340), .D
		(n_181764152), .Z(n_200864343));
	notech_ao4 i_133954009(.A(n_2662), .B(n_29077), .C(n_57348), .D(n_2663),
		 .Z(n_200564340));
	notech_ao4 i_134254006(.A(\nbus_11276[10] ), .B(n_177664114), .C(nbus_11273
		[10]), .D(n_26331), .Z(n_200364338));
	notech_ao4 i_134354005(.A(n_174258030), .B(n_324388255), .C(n_319431581)
		, .D(n_55867), .Z(n_200164336));
	notech_and4 i_134953999(.A(n_55901), .B(n_199764332), .C(n_182564160), .D
		(n_26247), .Z(n_200064335));
	notech_ao4 i_134754001(.A(n_2662), .B(n_29080), .C(n_57347), .D(n_2663),
		 .Z(n_199764332));
	notech_and4 i_135453994(.A(n_199464329), .B(n_183164166), .C(n_199264327
		), .D(n_182864163), .Z(n_199664331));
	notech_ao4 i_135053998(.A(n_327565579), .B(nbus_11273[11]), .C(n_327665580
		), .D(n_27576), .Z(n_199464329));
	notech_ao4 i_135253996(.A(n_171658004), .B(n_324388255), .C(n_238768192)
		, .D(n_55867), .Z(n_199264327));
	notech_and4 i_135853990(.A(n_198864323), .B(n_183264167), .C(n_183564170
		), .D(n_26409), .Z(n_199164326));
	notech_ao4 i_135653992(.A(n_57346), .B(n_2663), .C(\nbus_11276[12] ), .D
		(n_327465578), .Z(n_198864323));
	notech_ao4 i_135953989(.A(n_327565579), .B(nbus_11273[12]), .C(n_327665580
		), .D(n_27577), .Z(n_198664321));
	notech_ao4 i_136053988(.A(n_169057978), .B(n_324388255), .C(n_189074758)
		, .D(n_55867), .Z(n_198464319));
	notech_and4 i_136653982(.A(n_55901), .B(n_198064315), .C(n_26408), .D(n_184364178
		), .Z(n_198364318));
	notech_ao4 i_136453984(.A(n_2662), .B(n_29037), .C(n_57345), .D(n_2663),
		 .Z(n_198064315));
	notech_and4 i_137153977(.A(n_197764312), .B(n_184964184), .C(n_197564310
		), .D(n_184664181), .Z(n_197964314));
	notech_ao4 i_136753981(.A(nbus_11273[13]), .B(n_327565579), .C(n_27578),
		 .D(n_327665580), .Z(n_197764312));
	notech_ao4 i_136953979(.A(n_166457952), .B(n_324388255), .C(n_187874746)
		, .D(n_55867), .Z(n_197564310));
	notech_and4 i_137553973(.A(n_55876), .B(n_363088165), .C(n_197164306), .D
		(n_185264187), .Z(n_197464309));
	notech_ao4 i_137353975(.A(n_2662), .B(n_29087), .C(n_2663), .D(n_356476400
		), .Z(n_197164306));
	notech_and4 i_138053968(.A(n_196864303), .B(n_185864193), .C(n_196664301
		), .D(n_185564190), .Z(n_197064305));
	notech_ao4 i_137653972(.A(n_327565579), .B(nbus_11273[15]), .C(n_327665580
		), .D(n_27581), .Z(n_196864303));
	notech_ao4 i_137853970(.A(n_177164109), .B(n_324288256), .C(n_177264110)
		, .D(n_324388255), .Z(n_196664301));
	notech_and4 i_138453964(.A(n_55901), .B(n_196264297), .C(n_316831555), .D
		(n_186164196), .Z(n_196564300));
	notech_ao4 i_138253966(.A(n_328565589), .B(nbus_11326[24]), .C(n_323165548
		), .D(nbus_11273[24]), .Z(n_196264297));
	notech_and4 i_138953959(.A(n_195964294), .B(n_186764202), .C(n_195764292
		), .D(n_186464199), .Z(n_196164296));
	notech_ao4 i_138553963(.A(n_57334), .B(n_323365550), .C(n_29137), .D(n_322965546
		), .Z(n_195964294));
	notech_ao4 i_138753961(.A(n_322231609), .B(n_328765591), .C(n_251061538)
		, .D(n_328665590), .Z(n_195764292));
	notech_and4 i_148153876(.A(n_195464289), .B(n_195264287), .C(n_187064205
		), .D(n_187364208), .Z(n_195664291));
	notech_ao4 i_147553880(.A(n_55977), .B(n_28426), .C(n_56024), .D(n_29203
		), .Z(n_195464289));
	notech_ao4 i_147953878(.A(n_59190), .B(n_26697), .C(n_55738), .D(n_27577
		), .Z(n_195264287));
	notech_and4 i_148753870(.A(n_194964284), .B(n_194764282), .C(n_194664281
		), .D(n_187664211), .Z(n_195164286));
	notech_ao4 i_148253875(.A(n_57346), .B(n_55519), .C(n_55382), .D(nbus_11273
		[12]), .Z(n_194964284));
	notech_ao4 i_148453873(.A(n_55381), .B(\nbus_11276[12] ), .C(n_321931606
		), .D(n_320465521), .Z(n_194764282));
	notech_ao4 i_148553872(.A(n_169157979), .B(n_320565522), .C(n_169057978)
		, .D(n_320665523), .Z(n_194664281));
	notech_and4 i_150353854(.A(n_194364278), .B(n_194164276), .C(n_188364218
		), .D(n_188664221), .Z(n_194564280));
	notech_ao4 i_149953858(.A(n_55977), .B(n_28429), .C(n_56024), .D(n_29204
		), .Z(n_194364278));
	notech_nand2 i_110467190(.A(n_56310), .B(n_56178), .Z(n_127467094));
	notech_nand2 i_217804(.A(n_128667106), .B(n_128567105), .Z(write_data_26
		[1]));
	notech_nand2 i_1017812(.A(n_128867108), .B(n_128767107), .Z(write_data_26
		[9]));
	notech_ao4 i_111767177(.A(n_28442003), .B(n_27298), .C(n_56414), .D(n_26925
		), .Z(n_128567105));
	notech_ao4 i_111867176(.A(n_27341992), .B(n_27334), .C(n_26595), .D(n_57357
		), .Z(n_128667106));
	notech_ao4 i_117367121(.A(n_28442003), .B(n_27310), .C(n_56414), .D(n_26941
		), .Z(n_128767107));
	notech_ao4 i_117467120(.A(n_27341992), .B(n_27342), .C(n_57349), .D(n_26595
		), .Z(n_128867108));
	notech_ao4 i_8463463(.A(n_34533), .B(n_54507), .C(n_323688454), .D(n_59926
		), .Z(n_128967109));
	notech_nand3 i_22463335(.A(n_1416), .B(tsc[33]), .C(n_59845), .Z(n_129467114
		));
	notech_or2 i_21963340(.A(n_2665), .B(\nbus_11276[1] ), .Z(n_129967119)
		);
	notech_or4 i_23463326(.A(n_56081), .B(n_56120), .C(n_55837), .D(n_57324)
		, .Z(n_130367123));
	notech_or2 i_22963331(.A(n_2665), .B(\nbus_11276[2] ), .Z(n_130867128)
		);
	notech_or2 i_33363228(.A(n_54748), .B(n_29049), .Z(n_130967129));
	notech_or2 i_32863233(.A(n_54921), .B(nbus_11273[1]), .Z(n_131667136));
	notech_or2 i_34163220(.A(n_54748), .B(n_29050), .Z(n_131767137));
	notech_or2 i_33663225(.A(n_54921), .B(nbus_11273[2]), .Z(n_132467144));
	notech_or2 i_34963213(.A(n_54748), .B(n_29043), .Z(n_132567145));
	notech_nao3 i_37663189(.A(n_2420), .B(n_29091), .C(n_232761396), .Z(n_133667156
		));
	notech_or2 i_37363192(.A(n_55422), .B(n_322688464), .Z(n_133967159));
	notech_nao3 i_37063195(.A(opc_10[3]), .B(n_62413), .C(n_261136766), .Z(n_134267162
		));
	notech_or2 i_39763168(.A(n_54436), .B(n_29049), .Z(n_134367163));
	notech_nand2 i_39263173(.A(n_54665), .B(opa[1]), .Z(n_135067170));
	notech_or2 i_40563160(.A(n_54436), .B(n_29050), .Z(n_135167171));
	notech_nand2 i_40063165(.A(n_54665), .B(opa[2]), .Z(n_135867178));
	notech_or2 i_41263153(.A(n_54436), .B(n_29043), .Z(n_135967179));
	notech_or4 i_44463121(.A(n_59370), .B(n_2645), .C(n_59926), .D(nbus_11326
		[1]), .Z(n_136667186));
	notech_or2 i_44363122(.A(n_54435), .B(n_29049), .Z(n_136967189));
	notech_or2 i_43863127(.A(n_54565), .B(nbus_11273[1]), .Z(n_137467194));
	notech_or4 i_45363112(.A(n_59370), .B(n_2645), .C(n_59922), .D(nbus_11326
		[2]), .Z(n_137567195));
	notech_or2 i_45263113(.A(n_54435), .B(n_29050), .Z(n_137867198));
	notech_or2 i_44763118(.A(n_54565), .B(nbus_11273[2]), .Z(n_138367203));
	notech_or2 i_47863087(.A(n_356176397), .B(n_29049), .Z(n_138467204));
	notech_nand2 i_47363092(.A(n_54661), .B(opa[1]), .Z(n_139167211));
	notech_or2 i_48663079(.A(n_356176397), .B(n_29050), .Z(n_139267212));
	notech_nand2 i_48163084(.A(n_54661), .B(opa[2]), .Z(n_139967219));
	notech_or2 i_49363072(.A(n_356176397), .B(n_29043), .Z(n_140067220));
	notech_or2 i_53263033(.A(n_54450), .B(n_29050), .Z(n_140767227));
	notech_or2 i_52763038(.A(n_271668515), .B(nbus_11273[2]), .Z(n_141467234
		));
	notech_or2 i_53963026(.A(n_54450), .B(n_29043), .Z(n_141567235));
	notech_or2 i_54763018(.A(n_54450), .B(n_29063), .Z(n_142267242));
	notech_or2 i_54263023(.A(n_271668515), .B(nbus_11273[4]), .Z(n_142967249
		));
	notech_or2 i_56263003(.A(n_54450), .B(n_29068), .Z(n_143067250));
	notech_or2 i_55763008(.A(n_271668515), .B(nbus_11273[6]), .Z(n_143767257
		));
	notech_or2 i_57062995(.A(n_54468), .B(n_29049), .Z(n_143867258));
	notech_nand2 i_56563000(.A(n_2670), .B(opa[1]), .Z(n_144567265));
	notech_or2 i_57862987(.A(n_54468), .B(n_29050), .Z(n_144667266));
	notech_nand2 i_57362992(.A(n_2670), .B(opa[2]), .Z(n_145367273));
	notech_or2 i_58662980(.A(n_54468), .B(n_29043), .Z(n_145467274));
	notech_or4 i_62762941(.A(n_56201), .B(n_274288715), .C(n_55837), .D(n_57325
		), .Z(n_146167281));
	notech_or2 i_62262946(.A(n_54438), .B(n_29049), .Z(n_146867288));
	notech_or4 i_63662933(.A(n_56201), .B(n_274288715), .C(n_55837), .D(n_57324
		), .Z(n_146967289));
	notech_or2 i_63062938(.A(n_54438), .B(n_29050), .Z(n_147667296));
	notech_or2 i_64362926(.A(n_55972), .B(n_203567855), .Z(n_147767297));
	notech_ao4 i_143262160(.A(n_279739585), .B(n_353369305), .C(n_275539543)
		, .D(n_353269304), .Z(n_148767307));
	notech_ao4 i_143162161(.A(n_54469), .B(n_322688464), .C(n_54438), .D(n_29043
		), .Z(n_148867308));
	notech_ao4 i_142962163(.A(n_54656), .B(nbus_11273[3]), .C(n_54655), .D(\nbus_11276[3] 
		), .Z(n_149067310));
	notech_and3 i_143062162(.A(n_201667836), .B(n_149067310), .C(n_147767297
		), .Z(n_149267312));
	notech_ao4 i_142562167(.A(n_279739585), .B(n_353569307), .C(n_275539543)
		, .D(n_353469306), .Z(n_149367313));
	notech_ao4 i_142462168(.A(n_54655), .B(\nbus_11276[2] ), .C(n_54469), .D
		(n_322488466), .Z(n_149567315));
	notech_and3 i_142762165(.A(n_149367313), .B(n_149567315), .C(n_147667296
		), .Z(n_149667316));
	notech_ao4 i_142262170(.A(n_55756), .B(n_27563), .C(n_54656), .D(nbus_11273
		[2]), .Z(n_149767317));
	notech_ao4 i_141862174(.A(n_279739585), .B(n_353869309), .C(n_275539543)
		, .D(n_353769308), .Z(n_150067320));
	notech_ao4 i_141762175(.A(n_54655), .B(\nbus_11276[1] ), .C(n_54469), .D
		(n_57357), .Z(n_150267322));
	notech_and3 i_142062172(.A(n_150067320), .B(n_150267322), .C(n_146867288
		), .Z(n_150367323));
	notech_ao4 i_141562177(.A(n_55756), .B(n_27562), .C(n_54656), .D(nbus_11273
		[1]), .Z(n_150467324));
	notech_ao4 i_138362209(.A(n_269839486), .B(nbus_11273[3]), .C(n_353369305
		), .D(n_2684), .Z(n_150867328));
	notech_ao4 i_138162210(.A(n_56144), .B(n_203567855), .C(n_269939487), .D
		(\nbus_11276[3] ), .Z(n_150967329));
	notech_ao4 i_137962212(.A(n_54428), .B(n_322688464), .C(n_2685), .D(n_353269304
		), .Z(n_151167331));
	notech_and3 i_138062211(.A(n_201667836), .B(n_151167331), .C(n_145467274
		), .Z(n_151367333));
	notech_ao4 i_137562216(.A(n_56144), .B(n_212767947), .C(n_2671), .D(n_27563
		), .Z(n_151467334));
	notech_ao4 i_137462217(.A(n_2685), .B(n_353469306), .C(n_2669), .D(\nbus_11276[2] 
		), .Z(n_151667336));
	notech_ao4 i_137262219(.A(n_54428), .B(n_322488466), .C(n_2684), .D(n_353569307
		), .Z(n_151867338));
	notech_and3 i_137362218(.A(n_201867838), .B(n_151867338), .C(n_144667266
		), .Z(n_152067340));
	notech_ao4 i_136862223(.A(n_56144), .B(n_201967839), .C(n_2671), .D(n_27562
		), .Z(n_152167341));
	notech_ao4 i_136762224(.A(n_2685), .B(n_353769308), .C(n_2669), .D(\nbus_11276[1] 
		), .Z(n_152367343));
	notech_and3 i_137062221(.A(n_152167341), .B(n_152367343), .C(n_144567265
		), .Z(n_152467344));
	notech_ao4 i_136562226(.A(n_54428), .B(n_57357), .C(n_2684), .D(n_353869309
		), .Z(n_152567345));
	notech_ao4 i_136162230(.A(n_56013), .B(n_144377843), .C(n_27568), .D(n_271768516
		), .Z(n_152867348));
	notech_ao4 i_136062231(.A(n_316588524), .B(n_247534101), .C(\nbus_11276[6] 
		), .D(n_271568514), .Z(n_153067350));
	notech_ao4 i_135862233(.A(n_57352), .B(n_54456), .C(n_316488525), .D(n_154267362
		), .Z(n_153267352));
	notech_and4 i_135962232(.A(n_183578230), .B(n_183478229), .C(n_153267352
		), .D(n_143067250), .Z(n_153467354));
	notech_ao4 i_134762244(.A(n_56013), .B(n_139770716), .C(n_271768516), .D
		(n_27565), .Z(n_153567355));
	notech_ao4 i_134662245(.A(n_316288527), .B(n_247534101), .C(n_271568514)
		, .D(\nbus_11276[4] ), .Z(n_153767357));
	notech_ao4 i_134462247(.A(n_321188478), .B(n_54456), .C(n_316388526), .D
		(n_154267362), .Z(n_153967359));
	notech_and3 i_134562246(.A(n_137970698), .B(n_153967359), .C(n_142267242
		), .Z(n_154167361));
	notech_or2 i_134262249(.A(n_54071), .B(n_324669045), .Z(n_154267362));
	notech_ao4 i_134062251(.A(n_269639484), .B(nbus_11273[3]), .C(n_353369305
		), .D(n_154267362), .Z(n_154367363));
	notech_ao4 i_133962252(.A(n_56013), .B(n_203567855), .C(n_269739485), .D
		(\nbus_11276[3] ), .Z(n_154467364));
	notech_ao4 i_133762254(.A(n_54456), .B(n_322688464), .C(n_247534101), .D
		(n_353269304), .Z(n_154667366));
	notech_and3 i_133862253(.A(n_201667836), .B(n_154667366), .C(n_141567235
		), .Z(n_154867368));
	notech_ao4 i_133362258(.A(n_56013), .B(n_212767947), .C(n_271768516), .D
		(n_27563), .Z(n_154967369));
	notech_ao4 i_133262259(.A(n_247534101), .B(n_353469306), .C(n_271568514)
		, .D(\nbus_11276[2] ), .Z(n_155167371));
	notech_and3 i_133562256(.A(n_154967369), .B(n_155167371), .C(n_141467234
		), .Z(n_155267372));
	notech_ao4 i_133062261(.A(n_54456), .B(n_322488466), .C(n_353569307), .D
		(n_154267362), .Z(n_155367373));
	notech_ao4 i_129662293(.A(n_268739475), .B(\nbus_11276[3] ), .C(n_353369305
		), .D(n_356276398), .Z(n_155767377));
	notech_ao4 i_129562294(.A(n_56049), .B(n_203567855), .C(n_269539483), .D
		(nbus_11273[3]), .Z(n_155867378));
	notech_ao4 i_129362296(.A(n_356076396), .B(n_322688464), .C(n_356376399)
		, .D(n_353269304), .Z(n_156067380));
	notech_and3 i_129462295(.A(n_201667836), .B(n_156067380), .C(n_140067220
		), .Z(n_156267382));
	notech_ao4 i_128962300(.A(n_56049), .B(n_212767947), .C(n_55753), .D(n_27563
		), .Z(n_156367383));
	notech_ao4 i_128862301(.A(n_356376399), .B(n_353469306), .C(n_54631), .D
		(\nbus_11276[2] ), .Z(n_156567385));
	notech_ao4 i_128662303(.A(n_356076396), .B(n_322488466), .C(n_356276398)
		, .D(n_353569307), .Z(n_156767387));
	notech_and3 i_128762302(.A(n_201867838), .B(n_156767387), .C(n_139267212
		), .Z(n_156967389));
	notech_ao4 i_128262307(.A(n_56049), .B(n_201967839), .C(n_55753), .D(n_27562
		), .Z(n_157067390));
	notech_ao4 i_128162308(.A(n_356376399), .B(n_353769308), .C(n_54631), .D
		(\nbus_11276[1] ), .Z(n_157267392));
	notech_and3 i_128462305(.A(n_157067390), .B(n_157267392), .C(n_139167211
		), .Z(n_157367393));
	notech_ao4 i_127962310(.A(n_356076396), .B(n_57357), .C(n_356276398), .D
		(n_353869309), .Z(n_157467394));
	notech_ao4 i_125962330(.A(n_56386), .B(n_212767947), .C(n_26539), .D(n_27563
		), .Z(n_157767397));
	notech_ao4 i_125862331(.A(n_247234098), .B(n_353469306), .C(n_54563), .D
		(\nbus_11276[2] ), .Z(n_157967399));
	notech_ao4 i_125562334(.A(n_322488466), .B(n_54458), .C(n_247334099), .D
		(n_353569307), .Z(n_158167401));
	notech_and4 i_125762332(.A(n_201867838), .B(n_158167401), .C(n_137567195
		), .D(n_137867198), .Z(n_158467404));
	notech_ao4 i_125162338(.A(n_56386), .B(n_201967839), .C(n_26539), .D(n_27562
		), .Z(n_158567405));
	notech_ao4 i_125062339(.A(n_247234098), .B(n_353769308), .C(n_54563), .D
		(\nbus_11276[1] ), .Z(n_158767407));
	notech_ao4 i_124762342(.A(n_57357), .B(n_54458), .C(n_247334099), .D(n_353869309
		), .Z(n_158967409));
	notech_and4 i_124962340(.A(n_136667186), .B(n_201767837), .C(n_158967409
		), .D(n_136967189), .Z(n_159267412));
	notech_ao4 i_122162367(.A(nbus_11273[3]), .B(n_269339481), .C(n_353369305
		), .D(n_254734173), .Z(n_159467414));
	notech_ao4 i_122062368(.A(n_56130), .B(n_203567855), .C(n_269439482), .D
		(\nbus_11276[3] ), .Z(n_159567415));
	notech_ao4 i_121862370(.A(n_322688464), .B(n_54432), .C(n_254634172), .D
		(n_353269304), .Z(n_159767417));
	notech_and3 i_121962369(.A(n_201667836), .B(n_159767417), .C(n_135967179
		), .Z(n_159967419));
	notech_ao4 i_121462374(.A(n_56130), .B(n_212767947), .C(n_55757), .D(n_27563
		), .Z(n_160067420));
	notech_ao4 i_121362375(.A(n_254634172), .B(n_353469306), .C(n_54664), .D
		(\nbus_11276[2] ), .Z(n_160267422));
	notech_ao4 i_121162377(.A(n_322488466), .B(n_54432), .C(n_254734173), .D
		(n_353569307), .Z(n_160467424));
	notech_and3 i_121262376(.A(n_201867838), .B(n_160467424), .C(n_135167171
		), .Z(n_160667426));
	notech_ao4 i_120762381(.A(n_56130), .B(n_201967839), .C(n_55757), .D(n_27562
		), .Z(n_160767427));
	notech_ao4 i_120662382(.A(n_254634172), .B(n_353769308), .C(n_54664), .D
		(\nbus_11276[1] ), .Z(n_160967429));
	notech_and3 i_120962379(.A(n_160767427), .B(n_160967429), .C(n_135067170
		), .Z(n_161067430));
	notech_ao4 i_120462384(.A(n_57357), .B(n_54432), .C(n_254734173), .D(n_353869309
		), .Z(n_161167431));
	notech_ao4 i_118962398(.A(n_353369305), .B(n_260436759), .C(n_59193), .D
		(n_26742), .Z(n_161467434));
	notech_ao4 i_118762400(.A(n_55304), .B(\nbus_11276[3] ), .C(n_55316), .D
		(nbus_11273[3]), .Z(n_161667436));
	notech_and4 i_119162396(.A(n_161667436), .B(n_134267162), .C(n_161467434
		), .D(n_133967159), .Z(n_161867438));
	notech_ao4 i_118462403(.A(n_262336778), .B(n_29247), .C(n_55421), .D(n_29043
		), .Z(n_161967439));
	notech_ao4 i_118262405(.A(n_5577), .B(n_57323), .C(n_55951), .D(n_27564)
		, .Z(n_162167441));
	notech_and4 i_118662401(.A(n_176567585), .B(n_162167441), .C(n_161967439
		), .D(n_133667156), .Z(n_162367443));
	notech_nand3 i_116762420(.A(n_62433), .B(opc[3]), .C(n_26381), .Z(n_162467444
		));
	notech_ao4 i_116562422(.A(n_55910), .B(n_203567855), .C(n_273539523), .D
		(n_162467444), .Z(n_162567445));
	notech_ao4 i_116462423(.A(n_54921), .B(nbus_11273[3]), .C(n_248434110), 
		.D(n_353269304), .Z(n_162667446));
	notech_ao4 i_116262425(.A(n_322688464), .B(n_54740), .C(n_54920), .D(\nbus_11276[3] 
		), .Z(n_162867448));
	notech_and3 i_116362424(.A(n_201667836), .B(n_162867448), .C(n_132567145
		), .Z(n_163067450));
	notech_ao4 i_115862429(.A(n_55910), .B(n_212767947), .C(n_55730), .D(n_27563
		), .Z(n_163167451));
	notech_ao4 i_115762430(.A(n_248434110), .B(n_353469306), .C(n_54920), .D
		(\nbus_11276[2] ), .Z(n_163367453));
	notech_and3 i_116062427(.A(n_163167451), .B(n_163367453), .C(n_132467144
		), .Z(n_163467454));
	notech_ao4 i_115562432(.A(n_322488466), .B(n_54740), .C(n_248734113), .D
		(n_353569307), .Z(n_163567455));
	notech_ao4 i_115162436(.A(n_55910), .B(n_201967839), .C(n_55730), .D(n_27562
		), .Z(n_163867458));
	notech_ao4 i_115062437(.A(n_248434110), .B(n_353769308), .C(n_54920), .D
		(\nbus_11276[1] ), .Z(n_164067460));
	notech_and3 i_115362434(.A(n_163867458), .B(n_164067460), .C(n_131667136
		), .Z(n_164167461));
	notech_ao4 i_114862439(.A(n_57357), .B(n_54740), .C(n_248734113), .D(n_353869309
		), .Z(n_164267462));
	notech_ao4 i_105862526(.A(n_2666), .B(nbus_11273[2]), .C(n_2687), .D(n_27563
		), .Z(n_164567465));
	notech_ao4 i_105762527(.A(n_2697), .B(n_353569307), .C(n_54606), .D(n_353469306
		), .Z(n_164767467));
	notech_and3 i_106062524(.A(n_164567465), .B(n_164767467), .C(n_130867128
		), .Z(n_164867468));
	notech_ao4 i_105462530(.A(n_2667), .B(n_29050), .C(n_2668), .D(n_322488466
		), .Z(n_164967469));
	notech_ao4 i_105362531(.A(n_27521), .B(n_59845), .C(n_107626780), .D(n_28715
		), .Z(n_165167471));
	notech_ao4 i_105062534(.A(n_2666), .B(nbus_11273[1]), .C(n_2687), .D(n_27562
		), .Z(n_165367473));
	notech_ao4 i_104962535(.A(n_2697), .B(n_353869309), .C(n_54606), .D(n_353769308
		), .Z(n_165567475));
	notech_and3 i_105262532(.A(n_165367473), .B(n_165567475), .C(n_129967119
		), .Z(n_165667476));
	notech_ao4 i_104662538(.A(n_2667), .B(n_29049), .C(n_2668), .D(n_57357),
		 .Z(n_165767477));
	notech_ao4 i_104562539(.A(n_27520), .B(n_59845), .C(n_57325), .D(n_2686)
		, .Z(n_165967479));
	notech_and3 i_82559785(.A(n_56061), .B(n_212664460), .C(n_222068039), .Z
		(n_166367483));
	notech_nand3 i_82859782(.A(n_55976), .B(n_258664903), .C(n_55974), .Z(n_166467484
		));
	notech_and2 i_83059780(.A(n_324869047), .B(n_340469177), .Z(n_166567485)
		);
	notech_or2 i_86759749(.A(n_36952), .B(n_55893), .Z(n_166667486));
	notech_or2 i_87059746(.A(n_36952), .B(n_56013), .Z(n_166767487));
	notech_nand3 i_11360442(.A(n_1416), .B(tsc[1]), .C(n_59845), .Z(n_167167491
		));
	notech_or2 i_11060445(.A(n_271368512), .B(n_29049), .Z(n_167467494));
	notech_or4 i_10760448(.A(n_58661), .B(n_56120), .C(n_54089), .D(n_27562)
		, .Z(n_167767497));
	notech_nand3 i_12360432(.A(n_1416), .B(tsc[2]), .C(n_59845), .Z(n_168167501
		));
	notech_or2 i_12060435(.A(n_271368512), .B(n_29050), .Z(n_168467504));
	notech_or4 i_11760438(.A(n_58661), .B(n_56120), .C(n_54089), .D(n_27563)
		, .Z(n_168767507));
	notech_or2 i_13460421(.A(n_61624), .B(nbus_11326[3]), .Z(n_168867508));
	notech_nand3 i_13360422(.A(n_1416), .B(tsc[3]), .C(n_59845), .Z(n_169167511
		));
	notech_nao3 i_13060425(.A(n_26248), .B(\opa_12[3] ), .C(n_351565804), .Z
		(n_169467514));
	notech_or4 i_12760428(.A(n_58661), .B(n_56120), .C(n_55837), .D(n_57323)
		, .Z(n_169767517));
	notech_or2 i_14460411(.A(n_61624), .B(nbus_11326[4]), .Z(n_169867518));
	notech_nand3 i_14360412(.A(n_1416), .B(tsc[4]), .C(n_59845), .Z(n_170167521
		));
	notech_or2 i_14060415(.A(n_271368512), .B(n_29063), .Z(n_170467524));
	notech_or4 i_13760418(.A(n_58660), .B(n_56120), .C(n_54089), .D(n_27565)
		, .Z(n_170767527));
	notech_nand3 i_15360402(.A(n_1416), .B(tsc[6]), .C(n_59845), .Z(n_171167531
		));
	notech_or2 i_15060405(.A(n_271368512), .B(n_29068), .Z(n_171467534));
	notech_or4 i_14760408(.A(n_58660), .B(n_56121), .C(n_54089), .D(n_27568)
		, .Z(n_171767537));
	notech_or2 i_26560293(.A(n_55893), .B(n_203567855), .Z(n_171867538));
	notech_or4 i_28060278(.A(n_55859), .B(n_57300), .C(n_56081), .D(n_59281)
		, .Z(n_172767547));
	notech_or2 i_27560283(.A(n_54945), .B(\nbus_11276[8] ), .Z(n_173267552)
		);
	notech_or2 i_42160150(.A(n_55910), .B(n_55085), .Z(n_173367553));
	notech_ao3 i_43160140(.A(n_62429), .B(opc[1]), .C(n_320688483), .Z(n_174467564
		));
	notech_or2 i_42860143(.A(n_319088499), .B(nbus_11273[1]), .Z(n_174767567
		));
	notech_nand3 i_42360148(.A(n_59193), .B(n_59922), .C(read_data[1]), .Z(n_175167571
		));
	notech_ao3 i_44660128(.A(n_62429), .B(opc[2]), .C(n_320688483), .Z(n_175667576
		));
	notech_or2 i_44260131(.A(n_319088499), .B(nbus_11273[2]), .Z(n_175967579
		));
	notech_nand3 i_43660136(.A(n_59193), .B(n_59922), .C(read_data[2]), .Z(n_176367583
		));
	notech_or4 i_46360115(.A(n_317788512), .B(n_320988480), .C(n_28054), .D(n_60511
		), .Z(n_176467584));
	notech_nand3 i_11388(.A(n_59190), .B(n_59922), .C(read_data[3]), .Z(n_176567585
		));
	notech_or2 i_46260116(.A(n_55222), .B(n_29043), .Z(n_176867588));
	notech_or4 i_45760119(.A(n_56573), .B(n_205088863), .C(n_56097), .D(n_57323
		), .Z(n_177167591));
	notech_or4 i_46460114(.A(n_60595), .B(n_59922), .C(n_55854), .D(\nbus_11276[3] 
		), .Z(n_177867598));
	notech_or4 i_46560113(.A(n_1135), .B(n_60595), .C(n_59922), .D(n_29043),
		 .Z(n_177967599));
	notech_or2 i_52660055(.A(n_340969182), .B(n_27574), .Z(n_178467604));
	notech_nand2 i_52160058(.A(opa[9]), .B(n_238568190), .Z(n_178767607));
	notech_or4 i_55360029(.A(n_55827), .B(n_58487), .C(n_57325), .D(n_60591)
		, .Z(n_179667616));
	notech_or2 i_55060032(.A(n_55316), .B(nbus_11273[1]), .Z(n_179967619));
	notech_nao3 i_54760035(.A(n_2416), .B(n_29091), .C(n_232761396), .Z(n_180267622
		));
	notech_or4 i_58560001(.A(n_55827), .B(n_58487), .C(n_57324), .D(n_60591)
		, .Z(n_180767627));
	notech_or2 i_58260004(.A(n_55316), .B(nbus_11273[2]), .Z(n_181067630));
	notech_nao3 i_57960007(.A(n_2418), .B(n_29091), .C(n_232761396), .Z(n_181367633
		));
	notech_or4 i_74459859(.A(n_55859), .B(n_57300), .C(n_56081), .D(n_56201)
		, .Z(n_181467634));
	notech_or2 i_73759864(.A(n_341269185), .B(\nbus_11276[8] ), .Z(n_182167641
		));
	notech_nor2 i_75359852(.A(n_55085), .B(n_56013), .Z(n_182267642));
	notech_or4 i_74559858(.A(n_1976), .B(n_355988238), .C(n_353069302), .D(n_233368141
		), .Z(n_182767647));
	notech_nao3 i_74659857(.A(opc_10[9]), .B(n_62413), .C(n_328069079), .Z(n_182867648
		));
	notech_or2 i_76359844(.A(n_341669189), .B(nbus_11326[29]), .Z(n_182967649
		));
	notech_or2 i_75659849(.A(n_326669065), .B(nbus_11273[29]), .Z(n_183667656
		));
	notech_nor2 i_81259798(.A(n_98113375), .B(nbus_11273[9]), .Z(n_184167661
		));
	notech_mux2 i_166559015(.S(n_59922), .A(n_260636761), .B(n_27528), .Z(n_184867668
		));
	notech_ao4 i_166459016(.A(n_2177), .B(n_57349), .C(n_56034), .D(\nbus_11276[9] 
		), .Z(n_185067670));
	notech_nao3 i_43860597(.A(n_185067670), .B(n_184867668), .C(n_184167661)
		, .Z(n_185167671));
	notech_ao4 i_162359056(.A(n_326769066), .B(\nbus_11276[29] ), .C(n_262936784
		), .D(n_55870), .Z(n_185267672));
	notech_ao4 i_162259057(.A(n_28977), .B(n_26224), .C(n_57329), .D(n_327069069
		), .Z(n_185467674));
	notech_and3 i_162559054(.A(n_185267672), .B(n_185467674), .C(n_183667656
		), .Z(n_185567675));
	notech_ao4 i_162059059(.A(n_110923096), .B(n_341569188), .C(n_270688747)
		, .D(n_341769190), .Z(n_185667676));
	notech_ao4 i_161559064(.A(nbus_11273[9]), .B(n_222368042), .C(\nbus_11276[9] 
		), .D(n_222468043), .Z(n_186167681));
	notech_nand3 i_161759062(.A(n_182767647), .B(n_186167681), .C(n_182867648
		), .Z(n_186267682));
	notech_ao4 i_161359066(.A(n_57349), .B(n_54457), .C(n_54460), .D(n_29048
		), .Z(n_186367683));
	notech_ao4 i_160959070(.A(n_161957907), .B(n_328069079), .C(n_161857906)
		, .D(n_327969078), .Z(n_186667686));
	notech_ao4 i_160859071(.A(n_341469187), .B(n_27571), .C(nbus_11273[8]), 
		.D(n_341369186), .Z(n_186867688));
	notech_ao4 i_160659073(.A(n_57350), .B(n_54457), .C(n_29045), .D(n_54460
		), .Z(n_187067690));
	notech_and3 i_160759072(.A(n_181467634), .B(n_187067690), .C(n_26404), .Z
		(n_187267692));
	notech_ao4 i_142559239(.A(n_261136766), .B(n_353469306), .C(n_260436759)
		, .D(n_353569307), .Z(n_187367693));
	notech_ao4 i_142359241(.A(n_55304), .B(\nbus_11276[2] ), .C(n_262336778)
		, .D(n_29257), .Z(n_187567695));
	notech_and4 i_142759237(.A(n_187567695), .B(n_187367693), .C(n_181067630
		), .D(n_181367633), .Z(n_187767697));
	notech_ao4 i_142059244(.A(n_55422), .B(n_322488466), .C(n_55421), .D(n_29050
		), .Z(n_187867698));
	notech_ao4 i_141859246(.A(n_59190), .B(n_26741), .C(n_55951), .D(n_27563
		), .Z(n_188067700));
	notech_and4 i_142259242(.A(n_188067700), .B(n_187867698), .C(n_176367583
		), .D(n_180767627), .Z(n_188267702));
	notech_ao4 i_136159296(.A(n_261136766), .B(n_353769308), .C(n_260436759)
		, .D(n_353869309), .Z(n_188367703));
	notech_ao4 i_135959298(.A(n_55304), .B(\nbus_11276[1] ), .C(n_262336778)
		, .D(n_29256), .Z(n_188567705));
	notech_and4 i_136359294(.A(n_188567705), .B(n_188367703), .C(n_179967619
		), .D(n_180267622), .Z(n_188767707));
	notech_ao4 i_135659301(.A(n_55422), .B(n_57357), .C(n_55421), .D(n_29049
		), .Z(n_188867708));
	notech_ao4 i_135359303(.A(n_59190), .B(n_26740), .C(n_55951), .D(n_27562
		), .Z(n_189067710));
	notech_and4 i_135859299(.A(n_189067710), .B(n_188867708), .C(n_175167571
		), .D(n_179667616), .Z(n_189267712));
	notech_ao4 i_133459318(.A(n_317388516), .B(n_29048), .C(n_59190), .D(n_26724
		), .Z(n_189367713));
	notech_ao4 i_133259319(.A(n_332269121), .B(n_353069302), .C(n_317588514)
		, .D(n_57349), .Z(n_189467714));
	notech_ao4 i_132959321(.A(n_352969301), .B(n_332369122), .C(n_317088519)
		, .D(n_57299), .Z(n_189667716));
	notech_and4 i_133659316(.A(n_189667716), .B(n_189467714), .C(n_189367713
		), .D(n_178767607), .Z(n_189867718));
	notech_ao4 i_132559324(.A(n_238668191), .B(\nbus_11276[9] ), .C(n_27528)
		, .D(n_59167), .Z(n_189967719));
	notech_ao4 i_132359326(.A(n_321688474), .B(n_29255), .C(n_321788473), .D
		(n_29254), .Z(n_190167721));
	notech_and3 i_132459325(.A(n_116357451), .B(n_116257450), .C(n_190167721
		), .Z(n_190267722));
	notech_ao4 i_127059374(.A(n_318888501), .B(\nbus_11276[3] ), .C(n_59190)
		, .D(n_26719), .Z(n_190467724));
	notech_ao4 i_126959375(.A(n_321788473), .B(n_29253), .C(n_320688483), .D
		(n_353369305), .Z(n_190567725));
	notech_ao4 i_126759377(.A(n_319288497), .B(n_27564), .C(n_321688474), .D
		(n_29252), .Z(n_190767727));
	notech_and4 i_127259372(.A(n_177167591), .B(n_190767727), .C(n_190567725
		), .D(n_190467724), .Z(n_190967729));
	notech_ao4 i_126459380(.A(n_55238), .B(n_322688464), .C(n_319088499), .D
		(nbus_11273[3]), .Z(n_191067730));
	notech_and2 i_127459370(.A(n_177967599), .B(n_177867598), .Z(n_191367733
		));
	notech_ao4 i_127359371(.A(n_316688523), .B(nbus_11273[3]), .C(n_316788522
		), .D(n_322688464), .Z(n_191467734));
	notech_and4 i_126359381(.A(n_191467734), .B(n_191367733), .C(n_176467584
		), .D(n_176567585), .Z(n_191767737));
	notech_ao4 i_125959385(.A(n_59167), .B(n_27521), .C(n_59190), .D(n_26718
		), .Z(n_191967739));
	notech_ao4 i_125859386(.A(n_55688), .B(n_57324), .C(n_319288497), .D(n_27563
		), .Z(n_192067740));
	notech_ao4 i_125659388(.A(n_55222), .B(n_29050), .C(n_55238), .D(n_322488466
		), .Z(n_192267742));
	notech_and4 i_126159383(.A(n_192267742), .B(n_192067740), .C(n_191967739
		), .D(n_175967579), .Z(n_192467744));
	notech_ao4 i_125359391(.A(n_320188488), .B(n_353469306), .C(n_318888501)
		, .D(\nbus_11276[2] ), .Z(n_192567745));
	notech_ao4 i_125159393(.A(n_321688474), .B(n_29251), .C(n_321788473), .D
		(n_29250), .Z(n_192767747));
	notech_nand3 i_125259392(.A(n_120557493), .B(n_132857616), .C(n_192767747
		), .Z(n_192867748));
	notech_ao4 i_124859396(.A(n_59167), .B(n_27520), .C(n_59188), .D(n_26717
		), .Z(n_193067750));
	notech_ao4 i_124759397(.A(n_55688), .B(n_57325), .C(n_319288497), .D(n_27562
		), .Z(n_193167751));
	notech_ao4 i_124559399(.A(n_55222), .B(n_29049), .C(n_55238), .D(n_57357
		), .Z(n_193367753));
	notech_and4 i_125059394(.A(n_193367753), .B(n_193167751), .C(n_193067750
		), .D(n_174767567), .Z(n_193567755));
	notech_ao4 i_124259402(.A(n_320188488), .B(n_353769308), .C(n_318888501)
		, .D(\nbus_11276[1] ), .Z(n_193667756));
	notech_ao4 i_124059404(.A(n_321688474), .B(n_29249), .C(n_321788473), .D
		(n_29248), .Z(n_193867758));
	notech_nand3 i_124159403(.A(n_120457492), .B(n_132957617), .C(n_193867758
		), .Z(n_193967759));
	notech_ao4 i_123659407(.A(n_318031567), .B(n_352969301), .C(n_353069302)
		, .D(n_318231569), .Z(n_194267762));
	notech_ao4 i_123559408(.A(n_54944), .B(nbus_11273[9]), .C(n_54902), .D(n_29048
		), .Z(n_194367763));
	notech_ao4 i_123359410(.A(n_54872), .B(n_57349), .C(\nbus_11276[9] ), .D
		(n_54943), .Z(n_194567765));
	notech_and3 i_123459409(.A(n_194567765), .B(n_26240), .C(n_173367553), .Z
		(n_194767767));
	notech_ao4 i_106559568(.A(n_161857906), .B(n_333569134), .C(n_161957907)
		, .D(n_333669135), .Z(n_194867768));
	notech_ao4 i_106459569(.A(n_55725), .B(n_27571), .C(n_54946), .D(nbus_11273
		[8]), .Z(n_195067770));
	notech_ao4 i_106159572(.A(n_57350), .B(n_54852), .C(n_29045), .D(n_54853
		), .Z(n_195267772));
	notech_and4 i_106359570(.A(n_55901), .B(n_172767547), .C(n_195267772), .D
		(n_26404), .Z(n_195567775));
	notech_nao3 i_104759582(.A(n_56492), .B(n_268064997), .C(n_353369305), .Z
		(n_195767777));
	notech_ao4 i_104559584(.A(n_353269304), .B(n_259336748), .C(n_150774375)
		, .D(n_195767777), .Z(n_195867778));
	notech_ao4 i_104459585(.A(n_54923), .B(nbus_11273[3]), .C(n_54922), .D(\nbus_11276[3] 
		), .Z(n_195967779));
	notech_ao4 i_104259587(.A(n_322688464), .B(n_54695), .C(n_54749), .D(n_29043
		), .Z(n_196167781));
	notech_and3 i_104359586(.A(n_201667836), .B(n_196167781), .C(n_171867538
		), .Z(n_196367783));
	notech_ao4 i_93459685(.A(n_57320), .B(n_268368482), .C(n_316488525), .D(n_268468483
		), .Z(n_196467784));
	notech_ao4 i_93259687(.A(n_271268511), .B(nbus_11273[6]), .C(n_271168510
		), .D(\nbus_11276[6] ), .Z(n_196667786));
	notech_and4 i_93659683(.A(n_196667786), .B(n_196467784), .C(n_171467534)
		, .D(n_171767537), .Z(n_196867788));
	notech_ao4 i_92759690(.A(n_316588524), .B(n_54607), .C(n_57352), .D(n_271468513
		), .Z(n_196967789));
	notech_ao4 i_92659691(.A(n_27525), .B(n_59847), .C(n_61624), .D(nbus_11326
		[6]), .Z(n_197167791));
	notech_ao4 i_92359694(.A(n_319588494), .B(n_268368482), .C(n_316388526),
		 .D(n_268468483), .Z(n_197367793));
	notech_ao4 i_92159696(.A(n_271268511), .B(nbus_11273[4]), .C(n_271168510
		), .D(\nbus_11276[4] ), .Z(n_197567795));
	notech_and4 i_92559692(.A(n_197567795), .B(n_197367793), .C(n_170467524)
		, .D(n_170767527), .Z(n_197767797));
	notech_ao4 i_91859699(.A(n_316288527), .B(n_54607), .C(n_321188478), .D(n_271468513
		), .Z(n_197867798));
	notech_and2 i_91759700(.A(n_137377773), .B(n_169867518), .Z(n_198067800)
		);
	notech_or4 i_91659701(.A(instrc[118]), .B(n_229364616), .C(n_55097), .D(instrc
		[119]), .Z(n_198267802));
	notech_ao4 i_91359704(.A(n_263036785), .B(n_27564), .C(n_353369305), .D(n_198267802
		), .Z(n_198367803));
	notech_ao4 i_91159706(.A(n_322688464), .B(n_355188244), .C(n_54948), .D(\nbus_11276[3] 
		), .Z(n_198567805));
	notech_and4 i_91559702(.A(n_198567805), .B(n_169767517), .C(n_198367803)
		, .D(n_169467514), .Z(n_198767807));
	notech_ao4 i_90859709(.A(n_353269304), .B(n_54607), .C(nbus_11273[3]), .D
		(n_26204), .Z(n_198867808));
	notech_and4 i_91059707(.A(n_201667836), .B(n_198867808), .C(n_168867508)
		, .D(n_169167511), .Z(n_199167811));
	notech_ao4 i_90359713(.A(n_57324), .B(n_268368482), .C(n_353569307), .D(n_268468483
		), .Z(n_199267812));
	notech_ao4 i_90159715(.A(n_271268511), .B(nbus_11273[2]), .C(n_271168510
		), .D(\nbus_11276[2] ), .Z(n_199467814));
	notech_and4 i_90659711(.A(n_199467814), .B(n_199267812), .C(n_168467504)
		, .D(n_168767507), .Z(n_199667816));
	notech_ao4 i_89859718(.A(n_353469306), .B(n_54607), .C(n_322488466), .D(n_271468513
		), .Z(n_199767817));
	notech_ao4 i_89659720(.A(n_27521), .B(n_59847), .C(n_61624), .D(nbus_11326
		[2]), .Z(n_199967819));
	notech_and4 i_90059716(.A(n_55876), .B(n_199967819), .C(n_199767817), .D
		(n_168167501), .Z(n_200167821));
	notech_ao4 i_89359723(.A(n_57325), .B(n_268368482), .C(n_353869309), .D(n_268468483
		), .Z(n_200267822));
	notech_ao4 i_89159725(.A(n_271268511), .B(nbus_11273[1]), .C(n_271168510
		), .D(\nbus_11276[1] ), .Z(n_200467824));
	notech_and4 i_89559721(.A(n_200467824), .B(n_200267822), .C(n_167467494)
		, .D(n_167767497), .Z(n_200667826));
	notech_ao4 i_88859728(.A(n_353769308), .B(n_54607), .C(n_57357), .D(n_271468513
		), .Z(n_200767827));
	notech_ao4 i_88659730(.A(n_27520), .B(n_59847), .C(n_61624), .D(nbus_11326
		[1]), .Z(n_200967829));
	notech_and4 i_89059726(.A(n_55876), .B(n_200967829), .C(n_200767827), .D
		(n_167167491), .Z(n_201167831));
	notech_nor2 i_12720(.A(n_54525), .B(n_201567835), .Z(n_201367833));
	notech_or4 i_12719(.A(n_1913), .B(n_204067860), .C(n_201567835), .D(n_60530
		), .Z(n_201467834));
	notech_ao4 i_35857902(.A(n_56502), .B(n_56112), .C(n_56063), .D(n_26250)
		, .Z(n_201567835));
	notech_and3 i_43657900(.A(n_213967959), .B(n_214167961), .C(n_213267952)
		, .Z(n_201667836));
	notech_and2 i_67057891(.A(n_214567965), .B(n_214467964), .Z(n_201767837)
		);
	notech_and2 i_67157890(.A(n_214367963), .B(n_214267962), .Z(n_201867838)
		);
	notech_or2 i_68657887(.A(n_55827), .B(n_57325), .Z(n_201967839));
	notech_nand3 i_153457860(.A(n_273688719), .B(n_59922), .C(n_26606), .Z(n_202067840
		));
	notech_and2 i_34657943(.A(n_56058), .B(n_203767857), .Z(n_202167841));
	notech_and2 i_4457813(.A(nbus_11273[2]), .B(n_202467844), .Z(n_202267842
		));
	notech_and2 i_4557812(.A(n_251834144), .B(n_251934145), .Z(n_202367843)
		);
	notech_nand3 i_63357259(.A(calc_sz[0]), .B(n_2041), .C(\opa_12[2] ), .Z(n_202467844
		));
	notech_or4 i_66657229(.A(n_205588858), .B(n_59370), .C(n_56573), .D(n_59922
		), .Z(n_202567845));
	notech_ao4 i_151657931(.A(n_54089), .B(n_27564), .C(n_55827), .D(n_57323
		), .Z(n_203567855));
	notech_or2 i_89757018(.A(n_55827), .B(n_26250), .Z(n_203767857));
	notech_or2 i_89957016(.A(n_55859), .B(n_26250), .Z(n_203967859));
	notech_ao4 i_180457857(.A(n_59380), .B(n_62405), .C(n_2264), .D(n_26241)
		, .Z(n_204067860));
	notech_or2 i_92856989(.A(n_55580), .B(n_55870), .Z(n_204367863));
	notech_nao3 i_55157330(.A(opc_10[1]), .B(n_62405), .C(n_259336748), .Z(n_204767867
		));
	notech_nand2 i_54657335(.A(n_55729), .B(opd[1]), .Z(n_205267872));
	notech_nao3 i_55957322(.A(opc_10[2]), .B(n_62401), .C(n_259336748), .Z(n_205567875
		));
	notech_nand2 i_55457327(.A(n_55729), .B(opd[2]), .Z(n_206067880));
	notech_nand3 i_61557272(.A(n_273688719), .B(n_59922), .C(n_275888699), .Z
		(n_206167881));
	notech_or2 i_61457273(.A(n_55740), .B(n_27562), .Z(n_206467884));
	notech_or2 i_61157276(.A(n_55380), .B(\nbus_11276[1] ), .Z(n_206767887)
		);
	notech_or4 i_60757279(.A(n_2145), .B(n_1976), .C(n_120857496), .D(n_353869309
		), .Z(n_207067890));
	notech_nand3 i_63257260(.A(n_273688719), .B(n_59922), .C(read_data[2]), 
		.Z(n_207367893));
	notech_or4 i_62857263(.A(n_56201), .B(n_273588720), .C(n_55827), .D(n_57324
		), .Z(n_207667896));
	notech_or2 i_62457266(.A(n_249734123), .B(n_29050), .Z(n_207967899));
	notech_or4 i_61857269(.A(n_2145), .B(n_1976), .C(n_120857496), .D(n_353569307
		), .Z(n_208267902));
	notech_or4 i_63657256(.A(n_2145), .B(n_1976), .C(n_120857496), .D(n_353369305
		), .Z(n_209167911));
	notech_ao4 i_66457230(.A(n_26605), .B(n_26592), .C(n_55836), .D(n_26570)
		, .Z(n_209267912));
	notech_nand3 i_73257175(.A(opa[0]), .B(nbus_11273[2]), .C(opa[1]), .Z(n_209367913
		));
	notech_nand2 i_73357174(.A(n_55114), .B(opa[2]), .Z(n_209467914));
	notech_or4 i_75257158(.A(n_59370), .B(n_2645), .C(n_59927), .D(nbus_11326
		[3]), .Z(n_209567915));
	notech_or2 i_74657163(.A(n_54435), .B(n_29043), .Z(n_210267922));
	notech_or2 i_79757116(.A(n_271768516), .B(n_27562), .Z(n_210367923));
	notech_or4 i_79257121(.A(n_56201), .B(n_56081), .C(n_55827), .D(n_57325)
		, .Z(n_211067930));
	notech_or2 i_83057084(.A(n_271768516), .B(n_27570), .Z(n_211167931));
	notech_or4 i_82557089(.A(n_55837), .B(n_2675), .C(n_56201), .D(n_56081),
		 .Z(n_211867938));
	notech_or2 i_27530(.A(n_55837), .B(n_57324), .Z(n_212767947));
	notech_or4 i_86857047(.A(n_60775), .B(n_60729), .C(n_1135), .D(n_29043),
		 .Z(n_213267952));
	notech_ao4 i_171756241(.A(n_2263), .B(n_26241), .C(n_204067860), .D(n_26318
		), .Z(n_213667956));
	notech_ao4 i_169256265(.A(n_55810), .B(nbus_11273[3]), .C(n_56045), .D(\nbus_11276[3] 
		), .Z(n_213967959));
	notech_ao4 i_169156266(.A(n_27522), .B(n_59847), .C(n_55920), .D(n_322688464
		), .Z(n_214167961));
	notech_ao4 i_168956268(.A(n_55810), .B(nbus_11273[2]), .C(n_249234118), 
		.D(n_59927), .Z(n_214267962));
	notech_ao4 i_168856269(.A(n_55920), .B(n_322488466), .C(n_27521), .D(n_59847
		), .Z(n_214367963));
	notech_ao4 i_168756270(.A(n_55810), .B(nbus_11273[1]), .C(n_249334119), 
		.D(n_59927), .Z(n_214467964));
	notech_ao4 i_168656271(.A(n_55920), .B(n_57357), .C(n_27520), .D(n_59847
		), .Z(n_214567965));
	notech_ao4 i_167456283(.A(n_2679), .B(n_247534101), .C(n_2680), .D(n_154267362
		), .Z(n_214667966));
	notech_ao4 i_167356284(.A(n_57351), .B(n_54456), .C(n_28983), .D(n_54450
		), .Z(n_214867968));
	notech_ao4 i_167156286(.A(n_271668515), .B(nbus_11273[7]), .C(n_271568514
		), .D(\nbus_11276[7] ), .Z(n_215067970));
	notech_and4 i_167256285(.A(n_174064078), .B(n_173964077), .C(n_215067970
		), .D(n_211167931), .Z(n_215267972));
	notech_ao4 i_160356354(.A(n_247534101), .B(n_353769308), .C(n_353869309)
		, .D(n_154267362), .Z(n_215367973));
	notech_ao4 i_160256355(.A(n_54456), .B(n_57357), .C(n_54450), .D(n_29049
		), .Z(n_215567975));
	notech_and3 i_160556352(.A(n_211067930), .B(n_215367973), .C(n_215567975
		), .Z(n_215667976));
	notech_ao4 i_160056357(.A(nbus_11273[1]), .B(n_271668515), .C(n_271568514
		), .D(\nbus_11276[1] ), .Z(n_215767977));
	notech_ao4 i_152656428(.A(n_247334099), .B(n_353369305), .C(n_247234098)
		, .D(n_353269304), .Z(n_216067980));
	notech_ao4 i_152556429(.A(n_56386), .B(n_203567855), .C(n_322688464), .D
		(n_54458), .Z(n_216267982));
	notech_and3 i_152856426(.A(n_216067980), .B(n_216267982), .C(n_210267922
		), .Z(n_216367983));
	notech_ao4 i_152356431(.A(n_54565), .B(nbus_11273[3]), .C(n_54563), .D(\nbus_11276[3] 
		), .Z(n_216467984));
	notech_nand3 i_6857906(.A(n_55482), .B(n_209467914), .C(n_209367913), .Z
		(n_216967989));
	notech_xor2 i_127757867(.A(opa[3]), .B(opa[4]), .Z(n_217067990));
	notech_xor2 i_7857905(.A(n_217067990), .B(n_216967989), .Z(n_217167991)
		);
	notech_xor2 i_90957877(.A(nbus_11273[5]), .B(opa[7]), .Z(n_217267992));
	notech_xor2 i_128857865(.A(opa[6]), .B(n_217267992), .Z(n_217367993));
	notech_xor2 i_90257907(.A(n_217367993), .B(n_217167991), .Z(n_217467994)
		);
	notech_nor2 i_146156488(.A(n_55821), .B(n_26191), .Z(n_55562));
	notech_ao4 i_144356506(.A(n_56667), .B(n_248934115), .C(n_202067840), .D
		(n_27522), .Z(n_217667996));
	notech_ao4 i_144256507(.A(n_29043), .B(n_249834124), .C(n_249534121), .D
		(n_353269304), .Z(n_217867998));
	notech_and3 i_144556504(.A(n_209167911), .B(n_217667996), .C(n_217867998
		), .Z(n_217967999));
	notech_ao4 i_144056509(.A(n_55518), .B(n_322688464), .C(n_55380), .D(\nbus_11276[3] 
		), .Z(n_218068000));
	notech_ao4 i_143956510(.A(n_55740), .B(n_27564), .C(n_55685), .D(n_57323
		), .Z(n_218168001));
	notech_or4 i_143856511(.A(n_205588858), .B(n_59370), .C(n_59927), .D(n_56104
		), .Z(n_218368003));
	notech_ao4 i_143556514(.A(n_217467994), .B(n_202367843), .C(n_218368003)
		, .D(n_202267842), .Z(n_218468004));
	notech_ao4 i_143356516(.A(n_249634122), .B(nbus_11273[2]), .C(n_249534121
		), .D(n_353469306), .Z(n_218668006));
	notech_and4 i_143756512(.A(n_218668006), .B(n_218468004), .C(n_207967899
		), .D(n_208267902), .Z(n_218868008));
	notech_ao4 i_143056519(.A(n_55518), .B(n_322488466), .C(n_55380), .D(\nbus_11276[2] 
		), .Z(n_218968009));
	notech_ao4 i_142856521(.A(n_54822), .B(n_26892), .C(n_55740), .D(n_27563
		), .Z(n_219168011));
	notech_and4 i_143256517(.A(n_219168011), .B(n_218968009), .C(n_207367893
		), .D(n_207667896), .Z(n_219368013));
	notech_ao4 i_142556524(.A(n_248934115), .B(nbus_11273[1]), .C(n_202067840
		), .D(n_27520), .Z(n_219468014));
	notech_ao4 i_142356526(.A(n_249834124), .B(n_29049), .C(n_249534121), .D
		(n_353769308), .Z(n_219668016));
	notech_and4 i_142756522(.A(n_219668016), .B(n_219468014), .C(n_206767887
		), .D(n_207067890), .Z(n_219868018));
	notech_ao4 i_142056529(.A(n_55685), .B(n_57325), .C(n_55518), .D(n_57357
		), .Z(n_219968019));
	notech_and4 i_142256527(.A(n_219968019), .B(n_54822), .C(n_206167881), .D
		(n_206467884), .Z(n_220268022));
	notech_ao4 i_137856569(.A(n_55893), .B(n_212767947), .C(n_248634112), .D
		(n_353569307), .Z(n_220368023));
	notech_ao4 i_137756570(.A(n_54749), .B(n_29050), .C(n_54922), .D(\nbus_11276[2] 
		), .Z(n_220568025));
	notech_ao4 i_137356573(.A(n_54923), .B(nbus_11273[2]), .C(n_322488466), 
		.D(n_54695), .Z(n_220768027));
	notech_and4 i_137556571(.A(n_55901), .B(n_220768027), .C(n_201867838), .D
		(n_205567875), .Z(n_221068030));
	notech_ao4 i_136956577(.A(n_55893), .B(n_201967839), .C(n_248634112), .D
		(n_353869309), .Z(n_221168031));
	notech_ao4 i_136856578(.A(n_54922), .B(\nbus_11276[1] ), .C(n_54923), .D
		(nbus_11273[1]), .Z(n_221368033));
	notech_ao4 i_136556581(.A(n_57357), .B(n_54695), .C(n_54749), .D(n_29049
		), .Z(n_221568035));
	notech_and4 i_136756579(.A(n_55901), .B(n_221568035), .C(n_201767837), .D
		(n_204767867), .Z(n_221968038));
	notech_and3 i_180855332(.A(n_56060), .B(n_213264466), .C(n_351065799), .Z
		(n_222068039));
	notech_or4 i_2155277(.A(n_212964463), .B(n_352665815), .C(n_60530), .D(n_2739
		), .Z(n_222168040));
	notech_or2 i_2255276(.A(n_351565804), .B(n_352665815), .Z(n_222268041)
		);
	notech_ao3 i_194060629(.A(n_326669065), .B(n_54450), .C(n_201367833), .Z
		(n_222368042));
	notech_and3 i_194260628(.A(n_326769066), .B(n_201467834), .C(n_54456), .Z
		(n_222468043));
	notech_and3 i_119754148(.A(n_317788512), .B(n_319388496), .C(n_316888521
		), .Z(n_222568044));
	notech_nand3 i_6055245(.A(n_1416), .B(tsc[10]), .C(n_59845), .Z(n_222868047
		));
	notech_or2 i_5755248(.A(n_57348), .B(n_350965798), .Z(n_223168050));
	notech_nand3 i_4955251(.A(n_62429), .B(opc[10]), .C(n_54545), .Z(n_223468053
		));
	notech_nor2 i_23855067(.A(n_54853), .B(n_29080), .Z(n_223568054));
	notech_ao3 i_23355072(.A(n_62429), .B(opc[11]), .C(n_333569134), .Z(n_224268061
		));
	notech_nao3 i_42054885(.A(n_3363), .B(\eflags[10] ), .C(n_54707), .Z(n_224568064
		));
	notech_nand2 i_41754888(.A(sav_esi[8]), .B(n_60595), .Z(n_225368067));
	notech_or2 i_41454891(.A(n_57350), .B(n_340769180), .Z(n_225768070));
	notech_or4 i_41154894(.A(n_273588720), .B(n_2240), .C(n_57300), .D(n_56121
		), .Z(n_226068073));
	notech_nao3 i_43254873(.A(n_3367), .B(\eflags[10] ), .C(n_54707), .Z(n_226168074
		));
	notech_nand2 i_42754878(.A(sav_esi[10]), .B(n_60595), .Z(n_226868081));
	notech_nao3 i_45054857(.A(n_3369), .B(\eflags[10] ), .C(n_54707), .Z(n_227568088
		));
	notech_nand2 i_44654860(.A(sav_esi[11]), .B(n_60595), .Z(n_227868091));
	notech_or2 i_44354863(.A(n_57347), .B(n_340769180), .Z(n_228168094));
	notech_or4 i_44054866(.A(n_273588720), .B(n_56121), .C(n_2240), .D(n_322031607
		), .Z(n_228468097));
	notech_nao3 i_46254845(.A(n_3371), .B(\eflags[10] ), .C(n_54707), .Z(n_228768100
		));
	notech_nand2 i_45954848(.A(sav_esi[12]), .B(n_60589), .Z(n_229068103));
	notech_or2 i_45654851(.A(n_57346), .B(n_340769180), .Z(n_229368106));
	notech_or4 i_45354854(.A(n_273588720), .B(n_56121), .C(n_2240), .D(n_321931606
		), .Z(n_229668109));
	notech_nao3 i_47554833(.A(n_3373), .B(\eflags[10] ), .C(n_54707), .Z(n_229968112
		));
	notech_nand2 i_47154836(.A(sav_esi[13]), .B(n_60589), .Z(n_230268115));
	notech_or2 i_46854839(.A(n_57345), .B(n_340769180), .Z(n_230568118));
	notech_or4 i_46554842(.A(n_273588720), .B(n_56121), .C(n_2240), .D(n_321831605
		), .Z(n_230868121));
	notech_nao3 i_48754821(.A(n_3377), .B(\eflags[10] ), .C(n_54707), .Z(n_231568124
		));
	notech_nand2 i_48454824(.A(sav_esi[15]), .B(n_60589), .Z(n_231868127));
	notech_or2 i_48154827(.A(n_340869181), .B(n_29087), .Z(n_232168130));
	notech_or2 i_47854830(.A(n_340569178), .B(\nbus_11276[15] ), .Z(n_232468133
		));
	notech_or2 i_81454511(.A(n_54460), .B(n_29077), .Z(n_232568134));
	notech_or4 i_80854517(.A(n_1976), .B(n_355988238), .C(n_233368141), .D(n_174358031
		), .Z(n_233168139));
	notech_or2 i_80954516(.A(n_319431581), .B(n_55870), .Z(n_233268140));
	notech_and4 i_190060638(.A(n_56058), .B(n_201567835), .C(n_340469177), .D
		(n_203767857), .Z(n_233368141));
	notech_nor2 i_82254503(.A(n_54460), .B(n_29080), .Z(n_233468142));
	notech_ao3 i_81754508(.A(n_62429), .B(opc[11]), .C(n_327969078), .Z(n_234168149
		));
	notech_nor2 i_83054495(.A(n_54460), .B(n_29084), .Z(n_234268150));
	notech_ao3 i_82554500(.A(n_62411), .B(opc[12]), .C(n_327969078), .Z(n_235268157
		));
	notech_nor2 i_84054487(.A(n_54460), .B(n_29037), .Z(n_235368158));
	notech_ao3 i_83554492(.A(n_62429), .B(opc[13]), .C(n_327969078), .Z(n_236068165
		));
	notech_or2 i_85054479(.A(n_54460), .B(n_29087), .Z(n_236168166));
	notech_or4 i_84354484(.A(n_57293), .B(n_55858), .C(n_56201), .D(n_56086)
		, .Z(n_236868173));
	notech_nor2 i_86054471(.A(n_341669189), .B(nbus_11326[24]), .Z(n_236968174
		));
	notech_or4 i_85354476(.A(n_56201), .B(n_56086), .C(n_56375), .D(n_27592)
		, .Z(n_237668181));
	notech_or2 i_93654397(.A(n_254834174), .B(\nbus_11276[11] ), .Z(n_238168186
		));
	notech_nand3 i_84555324(.A(n_55222), .B(n_319188498), .C(n_317288517), .Z
		(n_238568190));
	notech_and2 i_84755325(.A(n_323731624), .B(n_317488515), .Z(n_238668191)
		);
	notech_or2 i_63955303(.A(n_322031607), .B(n_55858), .Z(n_238768192));
	notech_ao4 i_199453369(.A(n_2333), .B(nbus_11273[11]), .C(n_27530), .D(n_59847
		), .Z(n_238868193));
	notech_ao4 i_199353370(.A(n_2331), .B(n_29080), .C(n_57347), .D(n_2177),
		 .Z(n_239068195));
	notech_nand3 i_64555301(.A(n_238868193), .B(n_239068195), .C(n_238168186
		), .Z(n_239168196));
	notech_ao4 i_193053432(.A(n_322231609), .B(n_341769190), .C(n_251061538)
		, .D(n_341569188), .Z(n_239268197));
	notech_ao4 i_192953433(.A(n_57334), .B(n_327069069), .C(n_29137), .D(n_26224
		), .Z(n_239468199));
	notech_nand3 i_193253430(.A(n_237668181), .B(n_239268197), .C(n_239468199
		), .Z(n_239568200));
	notech_ao4 i_192753435(.A(n_326669065), .B(nbus_11273[24]), .C(n_326769066
		), .D(\nbus_11276[24] ), .Z(n_239668201));
	notech_ao4 i_192153439(.A(n_177164109), .B(n_327969078), .C(n_177264110)
		, .D(n_328069079), .Z(n_239968204));
	notech_ao4 i_192053440(.A(nbus_11273[15]), .B(n_341369186), .C(n_341469187
		), .D(n_27581), .Z(n_240168206));
	notech_and3 i_192353437(.A(n_236868173), .B(n_239968204), .C(n_240168206
		), .Z(n_240268207));
	notech_ao4 i_191853442(.A(n_356476400), .B(n_54457), .C(n_341269185), .D
		(\nbus_11276[15] ), .Z(n_240368208));
	notech_ao4 i_191453446(.A(n_166457952), .B(n_328069079), .C(n_187874746)
		, .D(n_55870), .Z(n_240668211));
	notech_ao4 i_191353447(.A(nbus_11273[13]), .B(n_341369186), .C(n_27578),
		 .D(n_341469187), .Z(n_240868213));
	notech_nao3 i_191653444(.A(n_240668211), .B(n_240868213), .C(n_236068165
		), .Z(n_240968214));
	notech_ao4 i_191153449(.A(n_57345), .B(n_54457), .C(n_341269185), .D(\nbus_11276[13] 
		), .Z(n_241068215));
	notech_ao4 i_190753453(.A(n_169057978), .B(n_328069079), .C(n_189074758)
		, .D(n_55870), .Z(n_241368218));
	notech_ao4 i_190653454(.A(nbus_11273[12]), .B(n_341369186), .C(n_341469187
		), .D(n_27577), .Z(n_241568220));
	notech_nao3 i_190953451(.A(n_241368218), .B(n_241568220), .C(n_235268157
		), .Z(n_242268221));
	notech_ao4 i_190453456(.A(n_57346), .B(n_54457), .C(n_341269185), .D(\nbus_11276[12] 
		), .Z(n_242368222));
	notech_ao4 i_190053460(.A(n_171658004), .B(n_328069079), .C(n_55870), .D
		(n_238768192), .Z(n_242668225));
	notech_ao4 i_189953461(.A(nbus_11273[11]), .B(n_341369186), .C(n_341469187
		), .D(n_27576), .Z(n_242868227));
	notech_nao3 i_190253458(.A(n_242668225), .B(n_242868227), .C(n_234168149
		), .Z(n_242968228));
	notech_ao4 i_189753463(.A(n_57347), .B(n_54457), .C(\nbus_11276[11] ), .D
		(n_341269185), .Z(n_243068229));
	notech_ao4 i_189253468(.A(n_222368042), .B(nbus_11273[10]), .C(n_174258030
		), .D(n_328069079), .Z(n_243568234));
	notech_and3 i_189453466(.A(n_233168139), .B(n_243568234), .C(n_233268140
		), .Z(n_243668235));
	notech_ao4 i_189053470(.A(n_57348), .B(n_54457), .C(n_222468043), .D(\nbus_11276[10] 
		), .Z(n_243768236));
	notech_ao4 i_162253736(.A(n_177164109), .B(n_332269121), .C(n_177264110)
		, .D(n_332369122), .Z(n_244068239));
	notech_ao4 i_162053738(.A(n_356476400), .B(n_340769180), .C(n_340669179)
		, .D(nbus_11273[15]), .Z(n_244268241));
	notech_and4 i_162453734(.A(n_244268241), .B(n_244068239), .C(n_232168130
		), .D(n_232468133), .Z(n_244468243));
	notech_ao4 i_161753741(.A(n_57293), .B(n_317088519), .C(n_340969182), .D
		(n_27581), .Z(n_244568244));
	notech_ao4 i_161553743(.A(n_321788473), .B(n_29263), .C(n_59167), .D(n_27534
		), .Z(n_244768246));
	notech_and4 i_161953739(.A(n_244768246), .B(n_244568244), .C(n_231568124
		), .D(n_231868127), .Z(n_244968248));
	notech_ao4 i_161253746(.A(n_166557953), .B(n_332269121), .C(n_166457952)
		, .D(n_332369122), .Z(n_245068249));
	notech_ao4 i_161053748(.A(n_340669179), .B(nbus_11273[13]), .C(n_340569178
		), .D(\nbus_11276[13] ), .Z(n_245268251));
	notech_and4 i_161453744(.A(n_245268251), .B(n_245068249), .C(n_230568118
		), .D(n_230868121), .Z(n_245468253));
	notech_ao4 i_160753751(.A(n_27578), .B(n_340969182), .C(n_29037), .D(n_340869181
		), .Z(n_245568254));
	notech_ao4 i_160553753(.A(n_321788473), .B(n_29262), .C(n_59167), .D(n_27532
		), .Z(n_245768256));
	notech_and4 i_160953749(.A(n_245768256), .B(n_245568254), .C(n_229968112
		), .D(n_230268115), .Z(n_245968258));
	notech_ao4 i_160253756(.A(n_169157979), .B(n_332269121), .C(n_169057978)
		, .D(n_332369122), .Z(n_246068259));
	notech_ao4 i_160053758(.A(nbus_11273[12]), .B(n_340669179), .C(n_340569178
		), .D(\nbus_11276[12] ), .Z(n_246268261));
	notech_and4 i_160453754(.A(n_246268261), .B(n_246068259), .C(n_229368106
		), .D(n_229668109), .Z(n_246468263));
	notech_ao4 i_159753761(.A(n_340969182), .B(n_27577), .C(n_340869181), .D
		(n_29084), .Z(n_246568264));
	notech_ao4 i_159553763(.A(n_321788473), .B(n_29261), .C(n_59167), .D(n_27531
		), .Z(n_246768266));
	notech_and4 i_159953759(.A(n_246768266), .B(n_246568264), .C(n_228768100
		), .D(n_229068103), .Z(n_246968268));
	notech_ao4 i_159253766(.A(n_171758005), .B(n_332269121), .C(n_171658004)
		, .D(n_332369122), .Z(n_247068269));
	notech_ao4 i_159053768(.A(n_340669179), .B(nbus_11273[11]), .C(n_340569178
		), .D(\nbus_11276[11] ), .Z(n_247268271));
	notech_and4 i_159453764(.A(n_247268271), .B(n_247068269), .C(n_228168094
		), .D(n_228468097), .Z(n_247468273));
	notech_ao4 i_158753771(.A(n_340969182), .B(n_27576), .C(n_340869181), .D
		(n_29080), .Z(n_247568274));
	notech_ao4 i_158553773(.A(n_321788473), .B(n_29260), .C(n_59167), .D(n_27530
		), .Z(n_247768276));
	notech_and4 i_158953769(.A(n_247768276), .B(n_247568274), .C(n_227568088
		), .D(n_227868091), .Z(n_247968278));
	notech_ao4 i_158253776(.A(n_174358031), .B(n_332269121), .C(n_174258030)
		, .D(n_332369122), .Z(n_248068279));
	notech_ao4 i_158153777(.A(nbus_11273[10]), .B(n_26194), .C(n_322131608),
		 .D(n_317088519), .Z(n_248168280));
	notech_ao4 i_157953779(.A(n_340969182), .B(n_27575), .C(\nbus_11276[10] 
		), .D(n_238668191), .Z(n_248368282));
	notech_and4 i_158453774(.A(n_248368282), .B(n_248168280), .C(n_248068279
		), .D(n_226868081), .Z(n_248568284));
	notech_ao4 i_157653782(.A(n_57348), .B(n_317588514), .C(n_59167), .D(n_27529
		), .Z(n_248668285));
	notech_ao4 i_157553783(.A(n_321788473), .B(n_29259), .C(n_317388516), .D
		(n_29077), .Z(n_248768286));
	notech_and3 i_157453784(.A(n_176558053), .B(n_176458052), .C(n_226168074
		), .Z(n_249068289));
	notech_ao4 i_157053788(.A(n_161857906), .B(n_332269121), .C(n_161957907)
		, .D(n_332369122), .Z(n_249268291));
	notech_ao4 i_156853790(.A(n_340669179), .B(nbus_11273[8]), .C(n_340569178
		), .D(\nbus_11276[8] ), .Z(n_249468293));
	notech_and4 i_157253786(.A(n_249468293), .B(n_226068073), .C(n_249268291
		), .D(n_225768070), .Z(n_249668295));
	notech_ao4 i_156553793(.A(n_340969182), .B(n_27571), .C(n_340869181), .D
		(n_29045), .Z(n_249768296));
	notech_ao4 i_156353795(.A(n_321788473), .B(n_29258), .C(n_59167), .D(n_27527
		), .Z(n_249968298));
	notech_and4 i_156753791(.A(n_249968298), .B(n_249768296), .C(n_224568064
		), .D(n_225368067), .Z(n_250168300));
	notech_ao4 i_140253946(.A(n_171658004), .B(n_333669135), .C(n_55898), .D
		(n_238768192), .Z(n_250268301));
	notech_ao4 i_140153947(.A(n_54946), .B(nbus_11273[11]), .C(n_55725), .D(n_27576
		), .Z(n_250468303));
	notech_nao3 i_140453944(.A(n_250268301), .B(n_250468303), .C(n_224268061
		), .Z(n_250568304));
	notech_ao4 i_139953949(.A(n_57347), .B(n_54852), .C(\nbus_11276[11] ), .D
		(n_54945), .Z(n_250668305));
	notech_ao4 i_123454112(.A(n_336065662), .B(n_174258030), .C(n_319431581)
		, .D(n_56035), .Z(n_250968308));
	notech_ao4 i_123254114(.A(n_54572), .B(\nbus_11276[10] ), .C(n_54573), .D
		(nbus_11273[10]), .Z(n_251168310));
	notech_and4 i_123654110(.A(n_251168310), .B(n_250968308), .C(n_223168050
		), .D(n_223468053), .Z(n_251368312));
	notech_ao4 i_122954117(.A(n_61624), .B(nbus_11326[10]), .C(n_350865797),
		 .D(n_29077), .Z(n_251468313));
	notech_and4 i_123154115(.A(n_154070859), .B(n_55876), .C(n_251468313), .D
		(n_222868047), .Z(n_251768316));
	notech_and4 i_53451460(.A(n_55846), .B(n_205188862), .C(n_55833), .D(n_1963
		), .Z(n_259068389));
	notech_nor2 i_56351431(.A(n_55811), .B(n_2648), .Z(n_259568394));
	notech_mux2 i_1811675(.S(n_60136), .A(regs_14[17]), .B(add_len_pc32[17])
		, .Z(\add_len_pc[17] ));
	notech_nand2 i_56251432(.A(sav_epc[17]), .B(n_60589), .Z(n_260468403));
	notech_and2 i_56451430(.A(\add_len_pc[17] ), .B(n_55819), .Z(n_260568404
		));
	notech_ao3 i_56551429(.A(opc_10[17]), .B(n_62405), .C(n_2211), .Z(n_260668405
		));
	notech_or4 i_1820637(.A(n_260668405), .B(n_260568404), .C(n_276768566), 
		.D(n_259568394), .Z(n_20213));
	notech_nor2 i_58451412(.A(n_57299), .B(n_55693), .Z(n_260768406));
	notech_and4 i_143252094(.A(n_270768506), .B(n_270668505), .C(n_270268501
		), .D(n_270568504), .Z(n_57299));
	notech_nand2 i_58351413(.A(sav_epc[9]), .B(n_60589), .Z(n_261268411));
	notech_nao3 i_58851408(.A(opc_10[9]), .B(n_62413), .C(n_354369313), .Z(n_261368412
		));
	notech_ao3 i_59051406(.A(n_62429), .B(opc[9]), .C(n_354469314), .Z(n_261468413
		));
	notech_or2 i_58751409(.A(n_354269312), .B(\nbus_11276[9] ), .Z(n_261768416
		));
	notech_nor2 i_58551411(.A(n_353969310), .B(n_27574), .Z(n_261868417));
	notech_or4 i_1020629(.A(n_261868417), .B(n_277668575), .C(n_260768406), 
		.D(n_26205), .Z(n_20165));
	notech_and4 i_142652033(.A(n_275768556), .B(n_275668555), .C(n_275268551
		), .D(n_275568554), .Z(n_57323));
	notech_mux2 i_411661(.S(n_60136), .A(n_559), .B(add_len_pc32[3]), .Z(\add_len_pc[3] 
		));
	notech_nand2 i_71651293(.A(sav_epc[3]), .B(n_60589), .Z(n_262368422));
	notech_nand2 i_71851291(.A(\add_len_pc[3] ), .B(n_55819), .Z(n_262468423
		));
	notech_nao3 i_72351286(.A(opc_10[3]), .B(n_62413), .C(n_54526258), .Z(n_262568424
		));
	notech_nand2 i_72151288(.A(n_2692), .B(opa[3]), .Z(n_262868427));
	notech_nand3 i_420623(.A(n_278168580), .B(n_278068579), .C(n_278868587),
		 .Z(n_20129));
	notech_and4 i_142552034(.A(n_274368542), .B(n_274268541), .C(n_273868537
		), .D(n_274168540), .Z(n_57324));
	notech_mux2 i_311660(.S(n_60136), .A(n_558), .B(add_len_pc32[2]), .Z(\add_len_pc[2] 
		));
	notech_nand2 i_73951270(.A(sav_epc[2]), .B(n_60589), .Z(n_263568434));
	notech_nand2 i_74151268(.A(\add_len_pc[2] ), .B(n_55819), .Z(n_263668435
		));
	notech_nao3 i_74651263(.A(opc_10[2]), .B(n_62419), .C(n_54526258), .Z(n_263768436
		));
	notech_nand2 i_74451265(.A(n_2692), .B(opa[2]), .Z(n_264068439));
	notech_nand3 i_320622(.A(n_279168590), .B(n_279068589), .C(n_279868597),
		 .Z(n_20123));
	notech_and4 i_142452035(.A(n_272968528), .B(n_272868527), .C(n_272468523
		), .D(n_272768526), .Z(n_57325));
	notech_mux2 i_211659(.S(n_60136), .A(n_557), .B(add_len_pc32[1]), .Z(\add_len_pc[1] 
		));
	notech_nand2 i_76251247(.A(sav_epc[1]), .B(n_60589), .Z(n_264768446));
	notech_nand2 i_76451245(.A(\add_len_pc[1] ), .B(n_55819), .Z(n_264868447
		));
	notech_nao3 i_76951240(.A(opc_10[1]), .B(n_62413), .C(n_54526258), .Z(n_264968448
		));
	notech_nand2 i_76751242(.A(n_2692), .B(opa[1]), .Z(n_265268451));
	notech_nand3 i_220621(.A(n_280168600), .B(n_280068599), .C(n_280868607),
		 .Z(n_20117));
	notech_mux2 i_111658(.S(n_60136), .A(n_556), .B(add_len_pc32[0]), .Z(\add_len_pc[0] 
		));
	notech_nand2 i_81551194(.A(sav_epc[0]), .B(n_60589), .Z(n_265968458));
	notech_nand2 i_81651193(.A(\add_len_pc[0] ), .B(n_55819), .Z(n_266068459
		));
	notech_or2 i_81851191(.A(n_2690), .B(n_27561), .Z(n_266168460));
	notech_ao3 i_82151188(.A(n_62429), .B(opc[0]), .C(n_55426267), .Z(n_266468463
		));
	notech_nao3 i_120620(.A(n_281968618), .B(n_281768616), .C(n_266468463), 
		.Z(n_20111));
	notech_nor2 i_101751008(.A(n_2648), .B(n_341769190), .Z(n_266768466));
	notech_or2 i_101151014(.A(n_341669189), .B(nbus_11326[17]), .Z(n_266868467
		));
	notech_or4 i_101651009(.A(n_56201), .B(n_56086), .C(n_56375), .D(n_27583
		), .Z(n_267368472));
	notech_ao3 i_101851007(.A(opc_10[17]), .B(n_62399), .C(n_341569188), .Z(n_267468473
		));
	notech_or4 i_1820829(.A(n_282468623), .B(n_282168620), .C(n_267468473), 
		.D(n_266768466), .Z(n_19191));
	notech_or4 i_103450991(.A(n_56201), .B(n_56086), .C(n_2688), .D(n_55837)
		, .Z(n_267568474));
	notech_or2 i_103150994(.A(n_271768516), .B(n_27561), .Z(n_268068479));
	notech_nao3 i_103250993(.A(n_62411), .B(opc[0]), .C(n_154267362), .Z(n_268168480
		));
	notech_nao3 i_103350992(.A(opc_10[0]), .B(n_62401), .C(n_247534101), .Z(n_268268481
		));
	notech_and4 i_120812(.A(n_41726130), .B(n_283168630), .C(n_267568474), .D
		(n_268268481), .Z(n_19089));
	notech_or4 i_196160552(.A(n_59263), .B(n_59272), .C(n_56121), .D(n_55837
		), .Z(n_268368482));
	notech_or4 i_196660551(.A(instrc[118]), .B(n_229364616), .C(n_166367483)
		, .D(instrc[119]), .Z(n_268468483));
	notech_nao3 i_150350553(.A(n_62411), .B(opc[0]), .C(n_268468483), .Z(n_269368492
		));
	notech_and4 i_117226(.A(n_2698), .B(n_284068639), .C(n_284368642), .D(n_269368492
		), .Z(n_15774));
	notech_ao4 i_12751846(.A(n_56144), .B(n_27615), .C(n_56386), .D(n_29264)
		, .Z(n_269668495));
	notech_ao4 i_12851845(.A(n_56097), .B(n_27692), .C(n_56130), .D(n_27650)
		, .Z(n_269768496));
	notech_ao4 i_12951844(.A(n_55910), .B(n_27724), .C(n_54535), .D(n_27379)
		, .Z(n_269968498));
	notech_ao4 i_13051843(.A(n_55940), .B(n_27795), .C(n_55898), .D(n_27756)
		, .Z(n_270068499));
	notech_and4 i_13951834(.A(n_270068499), .B(n_269968498), .C(n_269768496)
		, .D(n_269668495), .Z(n_270268501));
	notech_ao4 i_13151842(.A(n_56049), .B(n_27859), .C(n_55867), .D(n_27827)
		, .Z(n_270368502));
	notech_ao4 i_13251841(.A(n_55870), .B(n_27928), .C(n_56035), .D(n_27896)
		, .Z(n_270468503));
	notech_and2 i_13751836(.A(n_270468503), .B(n_270368502), .Z(n_270568504)
		);
	notech_ao4 i_13351840(.A(n_55972), .B(n_27994), .C(n_55998), .D(n_27962)
		, .Z(n_270668505));
	notech_ao4 i_13451839(.A(n_58487), .B(n_28028), .C(n_55952), .D(n_29265)
		, .Z(n_270768506));
	notech_and4 i_186660642(.A(n_55142), .B(n_222168040), .C(n_350965798), .D
		(n_56045), .Z(n_271168510));
	notech_and4 i_186460643(.A(n_55143), .B(n_350865797), .C(n_55810), .D(n_222268041
		), .Z(n_271268511));
	notech_ao4 i_183260644(.A(n_1135), .B(n_59927), .C(n_351565804), .D(n_56032
		), .Z(n_271368512));
	notech_and2 i_183160645(.A(n_55920), .B(n_355188244), .Z(n_271468513));
	notech_and3 i_182057948(.A(n_54457), .B(n_326769066), .C(n_201467834), .Z
		(n_271568514));
	notech_ao3 i_181957949(.A(n_54460), .B(n_326669065), .C(n_201367833), .Z
		(n_271668515));
	notech_and2 i_59557983(.A(n_326869067), .B(n_204367863), .Z(n_271768516)
		);
	notech_ao4 i_29551682(.A(n_56144), .B(n_27605), .C(n_56386), .D(n_27560)
		, .Z(n_271868517));
	notech_ao4 i_29651681(.A(n_56097), .B(n_27682), .C(n_56130), .D(n_27640)
		, .Z(n_271968518));
	notech_ao4 i_29751680(.A(n_55910), .B(n_27716), .C(n_54535), .D(n_27371)
		, .Z(n_272168520));
	notech_ao4 i_29851679(.A(n_55940), .B(n_27787), .C(n_55898), .D(n_27748)
		, .Z(n_272268521));
	notech_and4 i_30751670(.A(n_272268521), .B(n_272168520), .C(n_271968518)
		, .D(n_271868517), .Z(n_272468523));
	notech_ao4 i_29951678(.A(n_56049), .B(n_27851), .C(n_55867), .D(n_27819)
		, .Z(n_272568524));
	notech_ao4 i_30051677(.A(n_55870), .B(n_27920), .C(n_56035), .D(n_27886)
		, .Z(n_272668525));
	notech_and2 i_30551672(.A(n_272668525), .B(n_272568524), .Z(n_272768526)
		);
	notech_ao4 i_30151676(.A(n_55972), .B(n_27986), .C(n_55998), .D(n_27954)
		, .Z(n_272868527));
	notech_ao4 i_30251675(.A(n_58487), .B(n_28020), .C(n_55952), .D(n_29266)
		, .Z(n_272968528));
	notech_ao4 i_33351648(.A(n_56144), .B(n_27608), .C(n_54439), .D(n_29115)
		, .Z(n_273268531));
	notech_ao4 i_33451647(.A(n_56097), .B(n_27685), .C(n_56130), .D(n_27641)
		, .Z(n_273368532));
	notech_ao4 i_33551646(.A(n_55864), .B(n_27717), .C(n_54535), .D(n_27372)
		, .Z(n_273568534));
	notech_ao4 i_33651645(.A(n_55940), .B(n_27788), .C(n_55898), .D(n_27749)
		, .Z(n_273668535));
	notech_and4 i_34651636(.A(n_273668535), .B(n_273568534), .C(n_273368532)
		, .D(n_273268531), .Z(n_273868537));
	notech_ao4 i_33751644(.A(n_56049), .B(n_27852), .C(n_55867), .D(n_27820)
		, .Z(n_273968538));
	notech_ao4 i_33851643(.A(n_55870), .B(n_27921), .C(n_56035), .D(n_27887)
		, .Z(n_274068539));
	notech_and2 i_34351638(.A(n_274068539), .B(n_273968538), .Z(n_274168540)
		);
	notech_ao4 i_33951642(.A(n_55972), .B(n_27987), .C(n_55998), .D(n_27955)
		, .Z(n_274268541));
	notech_ao4 i_34051641(.A(n_58487), .B(n_28021), .C(n_55952), .D(n_29121)
		, .Z(n_274368542));
	notech_ao4 i_37151614(.A(n_56144), .B(n_27609), .C(n_54439), .D(n_29117)
		, .Z(n_274668545));
	notech_ao4 i_37251613(.A(n_56097), .B(n_27686), .C(n_54451), .D(n_27642)
		, .Z(n_274768546));
	notech_ao4 i_37351612(.A(n_55864), .B(n_27718), .C(n_54535), .D(n_27373)
		, .Z(n_274968548));
	notech_ao4 i_37451611(.A(n_55940), .B(n_27789), .C(n_55898), .D(n_27750)
		, .Z(n_275068549));
	notech_and4 i_38551602(.A(n_275068549), .B(n_274968548), .C(n_274768546)
		, .D(n_274668545), .Z(n_275268551));
	notech_ao4 i_37551610(.A(n_56068), .B(n_27853), .C(n_55867), .D(n_27821)
		, .Z(n_275368552));
	notech_ao4 i_37651609(.A(n_55870), .B(n_27922), .C(n_56035), .D(n_27888)
		, .Z(n_275468553));
	notech_and2 i_38251604(.A(n_275468553), .B(n_275368552), .Z(n_275568554)
		);
	notech_ao4 i_37751608(.A(n_55972), .B(n_27988), .C(n_55998), .D(n_27956)
		, .Z(n_275668555));
	notech_ao4 i_37851607(.A(n_55878), .B(n_28022), .C(n_55952), .D(n_29116)
		, .Z(n_275768556));
	notech_ao4 i_56751427(.A(n_55587), .B(n_2700), .C(n_55568), .D(\nbus_11276[17] 
		), .Z(n_276068559));
	notech_ao4 i_56851426(.A(n_2345), .B(n_27537), .C(n_55597), .D(n_28987),
		 .Z(n_276168560));
	notech_ao4 i_56951425(.A(n_55842), .B(n_27583), .C(n_55808), .D(n_29267)
		, .Z(n_276368562));
	notech_ao4 i_56651428(.A(n_55567), .B(nbus_11273[17]), .C(n_2212), .D(nbus_11326
		[17]), .Z(n_276468563));
	notech_and3 i_57351422(.A(n_276468563), .B(n_276368562), .C(n_260468403)
		, .Z(n_276668565));
	notech_nand3 i_57451421(.A(n_276168560), .B(n_276068559), .C(n_276668565
		), .Z(n_276768566));
	notech_ao4 i_59151405(.A(n_55808), .B(n_29268), .C(n_2345), .D(n_27528),
		 .Z(n_277068569));
	notech_ao4 i_59251404(.A(n_57349), .B(n_55264), .C(n_29048), .D(n_55263)
		, .Z(n_277268571));
	notech_and4 i_59751401(.A(n_261368412), .B(n_277268571), .C(n_277068569)
		, .D(n_261268411), .Z(n_277468573));
	notech_nao3 i_60051398(.A(n_277468573), .B(n_261768416), .C(n_261468413)
		, .Z(n_277668575));
	notech_ao4 i_59951399(.A(n_26435), .B(n_29269), .C(nbus_11273[9]), .D(n_26434
		), .Z(n_277768576));
	notech_ao4 i_73251277(.A(n_353369305), .B(n_55426267), .C(n_55687), .D(n_57323
		), .Z(n_278068579));
	notech_ao4 i_73051279(.A(n_2691), .B(n_55277), .C(n_2690), .D(n_27564), 
		.Z(n_278168580));
	notech_ao4 i_72551284(.A(n_322688464), .B(n_55216), .C(n_55236), .D(n_29043
		), .Z(n_278268581));
	notech_ao4 i_72451285(.A(n_55808), .B(n_29270), .C(n_2345), .D(n_27522),
		 .Z(n_278368582));
	notech_and3 i_72751282(.A(n_278368582), .B(n_278268581), .C(n_262368422)
		, .Z(n_278568584));
	notech_and4 i_73151278(.A(n_262568424), .B(n_262468423), .C(n_278568584)
		, .D(n_262868427), .Z(n_278868587));
	notech_ao4 i_75551254(.A(n_353569307), .B(n_55426267), .C(n_55687), .D(n_57324
		), .Z(n_279068589));
	notech_ao4 i_75351256(.A(n_2691), .B(n_55289), .C(n_2690), .D(n_55299), 
		.Z(n_279168590));
	notech_ao4 i_74851261(.A(n_322488466), .B(n_55216), .C(n_55236), .D(n_29050
		), .Z(n_279268591));
	notech_ao4 i_74751262(.A(n_55808), .B(n_29271), .C(n_2345), .D(n_27521),
		 .Z(n_279368592));
	notech_and3 i_75051259(.A(n_279368592), .B(n_279268591), .C(n_263568434)
		, .Z(n_279568594));
	notech_and4 i_75451255(.A(n_263768436), .B(n_263668435), .C(n_279568594)
		, .D(n_264068439), .Z(n_279868597));
	notech_ao4 i_77851231(.A(n_353869309), .B(n_55426267), .C(n_57325), .D(n_55687
		), .Z(n_280068599));
	notech_ao4 i_77651233(.A(n_2691), .B(n_59753), .C(n_2690), .D(n_55331), 
		.Z(n_280168600));
	notech_ao4 i_77151238(.A(n_57357), .B(n_55216), .C(n_55236), .D(n_29049)
		, .Z(n_280268601));
	notech_ao4 i_77051239(.A(n_55808), .B(n_29272), .C(n_2345), .D(n_27520),
		 .Z(n_280368602));
	notech_and3 i_77351236(.A(n_280368602), .B(n_280268601), .C(n_264768446)
		, .Z(n_280568604));
	notech_and4 i_77751232(.A(n_264968448), .B(n_264868447), .C(n_280568604)
		, .D(n_265268451), .Z(n_280868607));
	notech_ao4 i_82451185(.A(n_2699), .B(n_55216), .C(n_55236), .D(n_28986),
		 .Z(n_281068609));
	notech_ao4 i_82351186(.A(n_58922), .B(n_29273), .C(n_2345), .D(n_27519),
		 .Z(n_281168610));
	notech_and3 i_82651183(.A(n_281168610), .B(n_281068609), .C(n_265968458)
		, .Z(n_281368612));
	notech_ao4 i_82951180(.A(nbus_11273[0]), .B(n_26203), .C(n_2691), .D(\nbus_11276[0] 
		), .Z(n_281668615));
	notech_and4 i_83051179(.A(n_281668615), .B(n_266068459), .C(n_281368612)
		, .D(n_266168460), .Z(n_281768616));
	notech_ao4 i_83251177(.A(n_43626149), .B(n_54526258), .C(n_2688), .D(n_55687
		), .Z(n_281968618));
	notech_nand3 i_102251003(.A(n_43426147), .B(n_266868467), .C(n_267368472
		), .Z(n_282168620));
	notech_ao4 i_102051005(.A(n_326769066), .B(\nbus_11276[17] ), .C(n_326669065
		), .D(nbus_11273[17]), .Z(n_282268621));
	notech_ao4 i_102151004(.A(n_26224), .B(n_28987), .C(n_327069069), .D(n_2700
		), .Z(n_282368622));
	notech_nand2 i_102351002(.A(n_282368622), .B(n_282268621), .Z(n_282468623
		));
	notech_ao4 i_103650989(.A(n_271568514), .B(\nbus_11276[0] ), .C(n_271668515
		), .D(nbus_11273[0]), .Z(n_282768626));
	notech_ao4 i_103550990(.A(n_54450), .B(n_28986), .C(n_54456), .D(n_2699)
		, .Z(n_282868627));
	notech_and4 i_103950986(.A(n_282868627), .B(n_282768626), .C(n_268068479
		), .D(n_268168480), .Z(n_283168630));
	notech_ao4 i_150550551(.A(n_61624), .B(nbus_11326[0]), .C(n_107626780), 
		.D(n_28708), .Z(n_283468633));
	notech_ao4 i_150650550(.A(n_271368512), .B(n_28986), .C(n_271468513), .D
		(n_2699), .Z(n_283568634));
	notech_ao4 i_150750549(.A(n_271168510), .B(\nbus_11276[0] ), .C(n_271268511
		), .D(nbus_11273[0]), .Z(n_283768636));
	notech_ao4 i_150850548(.A(n_323631623), .B(n_59927), .C(n_263036785), .D
		(n_27561), .Z(n_283868637));
	notech_and4 i_151150545(.A(n_283868637), .B(n_283768636), .C(n_283568634
		), .D(n_283468633), .Z(n_284068639));
	notech_ao4 i_151450542(.A(n_43626149), .B(n_54607), .C(n_2688), .D(n_268368482
		), .Z(n_284368642));
	notech_nand3 i_63449254(.A(n_2203), .B(n_54520), .C(n_26887), .Z(n_284468643
		));
	notech_nor2 i_18248982(.A(n_55353), .B(n_26599), .Z(n_284768646));
	notech_nand2 i_4149207(.A(n_26229), .B(n_62413), .Z(n_56223));
	notech_and3 i_23148933(.A(n_55958), .B(n_55959), .C(n_55961), .Z(n_284868647
		));
	notech_nor2 i_42548753(.A(n_101213406), .B(n_271088745), .Z(n_284968648)
		);
	notech_or2 i_42348755(.A(n_98113375), .B(nbus_11273[31]), .Z(n_285268651
		));
	notech_or4 i_42448754(.A(n_60775), .B(n_60726), .C(n_54761), .D(n_28996)
		, .Z(n_285368652));
	notech_or4 i_43648742(.A(n_56201), .B(n_274288715), .C(n_56375), .D(n_27601
		), .Z(n_285868657));
	notech_nao3 i_43548743(.A(opc_10[31]), .B(n_62417), .C(n_306621953), .Z(n_285968658
		));
	notech_nor2 i_43448744(.A(n_271288743), .B(n_309921986), .Z(n_286068659)
		);
	notech_nor2 i_43348745(.A(n_55396), .B(n_271088745), .Z(n_286168660));
	notech_or4 i_3220683(.A(n_102723014), .B(n_286068659), .C(n_286168660), 
		.D(n_26208), .Z(n_19971));
	notech_or4 i_47848703(.A(n_204788866), .B(n_56163), .C(n_56375), .D(n_27601
		), .Z(n_286668665));
	notech_nao3 i_47748704(.A(opc_10[31]), .B(n_62413), .C(n_2694), .Z(n_286768666
		));
	notech_nor2 i_47648705(.A(n_2674), .B(n_271288743), .Z(n_286868667));
	notech_nor2 i_47548706(.A(n_271088745), .B(n_2655), .Z(n_286968668));
	notech_or4 i_3220747(.A(n_102723014), .B(n_286868667), .C(n_286968668), 
		.D(n_26209), .Z(n_19623));
	notech_or4 i_51348671(.A(n_56201), .B(n_56086), .C(n_56375), .D(n_27601)
		, .Z(n_287468673));
	notech_nao3 i_51248672(.A(opc_10[31]), .B(n_62413), .C(n_341569188), .Z(n_287568674
		));
	notech_nor2 i_51148673(.A(n_341769190), .B(n_271288743), .Z(n_287668675)
		);
	notech_nor2 i_51048674(.A(n_327069069), .B(n_271088745), .Z(n_287768676)
		);
	notech_or4 i_3220843(.A(n_102723014), .B(n_287668675), .C(n_287768676), 
		.D(n_26210), .Z(n_19275));
	notech_or2 i_52648658(.A(n_326669065), .B(nbus_11273[30]), .Z(n_288268681
		));
	notech_nao3 i_52948655(.A(opc_10[30]), .B(n_62417), .C(n_341569188), .Z(n_288368682
		));
	notech_or4 i_52848656(.A(n_56201), .B(n_56086), .C(n_55798), .D(n_271188744
		), .Z(n_288468683));
	notech_or2 i_52748657(.A(n_327069069), .B(n_270988746), .Z(n_288568684)
		);
	notech_and4 i_3120842(.A(n_300068799), .B(n_101523002), .C(n_288468683),
		 .D(n_288568684), .Z(n_19269));
	notech_or4 i_59948591(.A(n_59263), .B(n_59272), .C(n_56203), .D(n_102623013
		), .Z(n_289068689));
	notech_nao3 i_59848592(.A(opc_10[31]), .B(n_62413), .C(n_308418861), .Z(n_289168690
		));
	notech_nor2 i_59748593(.A(n_271288743), .B(n_309618873), .Z(n_289268691)
		);
	notech_nor2 i_59648594(.A(n_55404), .B(n_271088745), .Z(n_289368692));
	notech_or4 i_3221003(.A(n_102723014), .B(n_289268691), .C(n_289368692), 
		.D(n_26211), .Z(n_16885));
	notech_or2 i_61248578(.A(n_55064), .B(nbus_11273[30]), .Z(n_289868697)
		);
	notech_nao3 i_61548575(.A(opc_10[30]), .B(n_62413), .C(n_308418861), .Z(n_289968698
		));
	notech_or4 i_61448576(.A(n_56203), .B(n_58660), .C(n_55798), .D(n_271188744
		), .Z(n_290068699));
	notech_or2 i_61348577(.A(n_55404), .B(n_270988746), .Z(n_290168700));
	notech_and4 i_3121002(.A(n_301468813), .B(n_101523002), .C(n_290068699),
		 .D(n_290168700), .Z(n_16879));
	notech_or4 i_63048560(.A(n_56203), .B(n_58660), .C(n_55798), .D(n_270688747
		), .Z(n_290268701));
	notech_or2 i_62448566(.A(n_55424), .B(nbus_11326[29]), .Z(n_290368702)
		);
	notech_or2 i_62948561(.A(n_55064), .B(nbus_11273[29]), .Z(n_290868707)
		);
	notech_nao3 i_63148559(.A(opc_10[29]), .B(n_62413), .C(n_308418861), .Z(n_290968708
		));
	notech_nand3 i_3021001(.A(n_302268821), .B(n_290968708), .C(n_290268701)
		, .Z(n_16873));
	notech_or2 i_64748544(.A(n_123423221), .B(nbus_11326[31]), .Z(n_291268711
		));
	notech_nao3 i_64848543(.A(opc_10[31]), .B(n_62413), .C(n_123623223), .Z(n_291568714
		));
	notech_nor2 i_64548546(.A(n_271288743), .B(n_123223219), .Z(n_291668715)
		);
	notech_nor2 i_64448547(.A(n_271088745), .B(n_2702), .Z(n_291768716));
	notech_or4 i_3221067(.A(n_291668715), .B(n_291768716), .C(n_102723014), 
		.D(n_26212), .Z(n_14001));
	notech_or4 i_81848386(.A(n_56203), .B(n_273588720), .C(n_55798), .D(n_270688747
		), .Z(n_291868717));
	notech_nao3 i_81948385(.A(opc_10[29]), .B(n_62419), .C(n_302721914), .Z(n_292568724
		));
	notech_or2 i_82048384(.A(n_113313527), .B(nbus_11326[29]), .Z(n_292668725
		));
	notech_nand3 i_3021321(.A(n_303668835), .B(n_291868717), .C(n_292668725)
		, .Z(n_20775));
	notech_or2 i_89348318(.A(n_55219), .B(nbus_11273[31]), .Z(n_293168730)
		);
	notech_nao3 i_89648315(.A(opc_10[31]), .B(n_62417), .C(n_308718864), .Z(n_293268731
		));
	notech_nor2 i_89548316(.A(n_271288743), .B(n_309518872), .Z(n_293368732)
		);
	notech_nor2 i_89448317(.A(n_55554), .B(n_271088745), .Z(n_293468733));
	notech_or4 i_3221611(.A(n_102723014), .B(n_293368732), .C(n_293468733), 
		.D(n_26213), .Z(n_13301));
	notech_nand2 i_100048216(.A(sav_esp[29]), .B(n_60589), .Z(n_294368742)
		);
	notech_nao3 i_100448212(.A(opc_10[29]), .B(n_62419), .C(n_110323090), .Z
		(n_294468743));
	notech_or2 i_100248214(.A(n_354688262), .B(n_28977), .Z(n_294768746));
	notech_nand3 i_3021737(.A(n_305468853), .B(n_304568844), .C(n_294768746)
		, .Z(n_12941));
	notech_or2 i_109948129(.A(n_55220), .B(nbus_11273[31]), .Z(n_295268751)
		);
	notech_nao3 i_110248126(.A(opc_10[31]), .B(n_62403), .C(n_322931616), .Z
		(n_295368752));
	notech_nor2 i_110148127(.A(n_322631613), .B(n_271288743), .Z(n_295468753
		));
	notech_nor2 i_110048128(.A(n_271088745), .B(n_55556), .Z(n_295568754));
	notech_or4 i_3221867(.A(n_102723014), .B(n_295468753), .C(n_295568754), 
		.D(n_26214), .Z(n_12587));
	notech_nand3 i_164647600(.A(n_55159), .B(n_59847), .C(mul64[29]), .Z(n_295668755
		));
	notech_or4 i_165847589(.A(n_57445), .B(n_59826), .C(n_2792), .D(n_27552)
		, .Z(n_296768766));
	notech_nand3 i_1416823(.A(n_306568864), .B(n_306368862), .C(n_307368872)
		, .Z(n_9772));
	notech_ao4 i_18448980(.A(n_54530), .B(n_55961), .C(n_26326), .D(n_55841)
		, .Z(n_296868767));
	notech_ao4 i_42648752(.A(n_56057), .B(\nbus_11276[31] ), .C(n_59837), .D
		(n_27554), .Z(n_297268771));
	notech_nand3 i_42848750(.A(n_297268771), .B(n_285268651), .C(n_285368652
		), .Z(n_297468773));
	notech_or2 i_45449185(.A(n_284968648), .B(n_297468773), .Z(n_102723014)
		);
	notech_or2 i_45649184(.A(n_56375), .B(n_27601), .Z(n_102623013));
	notech_ao4 i_43748741(.A(n_55071), .B(\nbus_11276[31] ), .C(n_303521922)
		, .D(nbus_11326[31]), .Z(n_297568774));
	notech_ao4 i_43848740(.A(n_55070), .B(nbus_11273[31]), .C(n_55397), .D(n_28996
		), .Z(n_297668775));
	notech_and4 i_44148737(.A(n_297668775), .B(n_297568774), .C(n_285868657)
		, .D(n_285968658), .Z(n_297968778));
	notech_ao4 i_47948702(.A(n_55069), .B(\nbus_11276[31] ), .C(n_2672), .D(nbus_11326
		[31]), .Z(n_298268781));
	notech_ao4 i_48048701(.A(n_55068), .B(nbus_11273[31]), .C(n_28996), .D(n_26444
		), .Z(n_298368782));
	notech_and4 i_48348698(.A(n_298368782), .B(n_298268781), .C(n_286668665)
		, .D(n_286768666), .Z(n_298668785));
	notech_ao4 i_51448670(.A(n_326769066), .B(\nbus_11276[31] ), .C(n_341669189
		), .D(nbus_11326[31]), .Z(n_298968788));
	notech_ao4 i_51548669(.A(n_326669065), .B(nbus_11273[31]), .C(n_26224), 
		.D(n_28996), .Z(n_299068789));
	notech_and4 i_51848666(.A(n_299068789), .B(n_298968788), .C(n_287468673)
		, .D(n_287568674), .Z(n_299368792));
	notech_ao4 i_53148653(.A(n_326869067), .B(n_27599), .C(n_26224), .D(n_28997
		), .Z(n_299668795));
	notech_ao4 i_53048654(.A(n_326769066), .B(\nbus_11276[30] ), .C(n_341669189
		), .D(nbus_11326[30]), .Z(n_299768796));
	notech_and4 i_53748650(.A(n_299768796), .B(n_299668795), .C(n_288268681)
		, .D(n_288368682), .Z(n_300068799));
	notech_ao4 i_60048590(.A(n_55062), .B(\nbus_11276[31] ), .C(n_55424), .D
		(nbus_11326[31]), .Z(n_300368802));
	notech_ao4 i_60148589(.A(n_55064), .B(nbus_11273[31]), .C(n_55405), .D(n_28996
		), .Z(n_300468803));
	notech_and4 i_60448586(.A(n_300468803), .B(n_300368802), .C(n_289068689)
		, .D(n_289168690), .Z(n_300768806));
	notech_ao4 i_61748573(.A(n_55720), .B(n_27599), .C(n_55405), .D(n_28997)
		, .Z(n_301068809));
	notech_ao4 i_61648574(.A(n_55062), .B(\nbus_11276[30] ), .C(n_55424), .D
		(nbus_11326[30]), .Z(n_301168810));
	notech_and4 i_62048570(.A(n_301168810), .B(n_301068809), .C(n_289868697)
		, .D(n_289968698), .Z(n_301468813));
	notech_and2 i_63248558(.A(n_262736782), .B(n_290368702), .Z(n_301768816)
		);
	notech_ao4 i_63348557(.A(n_55404), .B(n_57329), .C(n_55062), .D(\nbus_11276[29] 
		), .Z(n_301968818));
	notech_ao4 i_63548556(.A(n_54439), .B(n_262936784), .C(n_55405), .D(n_28977
		), .Z(n_302068819));
	notech_and4 i_63848553(.A(n_302068819), .B(n_301968818), .C(n_301768816)
		, .D(n_290868707), .Z(n_302268821));
	notech_ao4 i_64948542(.A(n_55073), .B(nbus_11273[31]), .C(n_55072), .D(\nbus_11276[31] 
		), .Z(n_302468823));
	notech_ao4 i_65148540(.A(n_54451), .B(n_102623013), .C(n_28996), .D(n_26450
		), .Z(n_302668825));
	notech_and4 i_65348538(.A(n_302468823), .B(n_302668825), .C(n_291268711)
		, .D(n_291568714), .Z(n_302868827));
	notech_ao4 i_82348381(.A(n_55562), .B(nbus_11273[29]), .C(n_55952), .D(n_262936784
		), .Z(n_303168830));
	notech_ao4 i_82148383(.A(n_55269), .B(n_57329), .C(n_55447), .D(\nbus_11276[29] 
		), .Z(n_303268831));
	notech_ao4 i_82248382(.A(n_2193), .B(n_27552), .C(n_55267), .D(n_28977),
		 .Z(n_303368832));
	notech_and4 i_82648378(.A(n_303368832), .B(n_303268831), .C(n_303168830)
		, .D(n_292568724), .Z(n_303668835));
	notech_ao4 i_89848313(.A(n_55773), .B(n_27601), .C(n_55555), .D(n_28996)
		, .Z(n_303868837));
	notech_ao4 i_89748314(.A(n_55218), .B(\nbus_11276[31] ), .C(nbus_11326[
		31]), .D(n_308318860), .Z(n_303968838));
	notech_and4 i_90148310(.A(n_303968838), .B(n_303868837), .C(n_293168730)
		, .D(n_293268731), .Z(n_304268841));
	notech_ao4 i_101548202(.A(n_110123088), .B(n_270688747), .C(n_354588263)
		, .D(n_57329), .Z(n_304568844));
	notech_ao4 i_100748210(.A(n_308518862), .B(nbus_11326[29]), .C(n_56024),
		 .D(n_29274), .Z(n_304668845));
	notech_ao4 i_100848209(.A(n_262536780), .B(n_27552), .C(n_55535), .D(\nbus_11276[29] 
		), .Z(n_304768846));
	notech_ao4 i_100948208(.A(n_55536), .B(nbus_11273[29]), .C(n_55135), .D(n_27597
		), .Z(n_304968848));
	notech_ao4 i_100548211(.A(n_55977), .B(n_28443), .C(n_262636781), .D(n_26983
		), .Z(n_305068849));
	notech_and3 i_101248205(.A(n_305068849), .B(n_304968848), .C(n_294368742
		), .Z(n_305268851));
	notech_and4 i_101448203(.A(n_304768846), .B(n_304668845), .C(n_305268851
		), .D(n_294468743), .Z(n_305468853));
	notech_ao4 i_110448124(.A(n_55772), .B(n_27601), .C(n_55557), .D(n_28996
		), .Z(n_305668855));
	notech_ao4 i_110348125(.A(n_55221), .B(\nbus_11276[31] ), .C(n_303421921
		), .D(nbus_11326[31]), .Z(n_305768856));
	notech_and4 i_110748121(.A(n_305768856), .B(n_305668855), .C(n_295268751
		), .D(n_295368752), .Z(n_306068859));
	notech_ao4 i_166447583(.A(n_54735), .B(nbus_11326[29]), .C(n_2249), .D(n_29278
		), .Z(n_306368862));
	notech_and4 i_166547582(.A(n_2786), .B(n_2186), .C(n_295668755), .D(n_296768766
		), .Z(n_306568864));
	notech_ao4 i_166047587(.A(n_55009), .B(n_28064), .C(n_54884), .D(\nbus_11276[5] 
		), .Z(n_306768866));
	notech_ao4 i_166147586(.A(n_2314), .B(\nbus_11276[13] ), .C(n_231547139)
		, .D(nbus_11326[21]), .Z(n_306868867));
	notech_ao4 i_166247585(.A(n_2247), .B(n_29276), .C(n_2313), .D(n_28913),
		 .Z(n_307068869));
	notech_ao4 i_166347584(.A(n_329546800), .B(n_29277), .C(n_2248), .D(nbus_11348
		[13]), .Z(n_307168870));
	notech_and4 i_166947578(.A(n_307168870), .B(n_307068869), .C(n_306868867
		), .D(n_306768866), .Z(n_307368872));
	notech_and3 i_2245351(.A(n_55961), .B(n_55959), .C(n_55958), .Z(n_307568874
		));
	notech_nor2 i_73444657(.A(n_341669189), .B(nbus_11326[23]), .Z(n_307768876
		));
	notech_or2 i_72944662(.A(n_308921976), .B(n_327069069), .Z(n_308468883)
		);
	notech_nor2 i_74244649(.A(n_341669189), .B(nbus_11326[25]), .Z(n_308568884
		));
	notech_or4 i_73744654(.A(n_56203), .B(n_56086), .C(n_55798), .D(n_308421971
		), .Z(n_309268891));
	notech_nor2 i_75044641(.A(n_341669189), .B(nbus_11326[26]), .Z(n_309368892
		));
	notech_or4 i_74544646(.A(n_56203), .B(n_56086), .C(n_55798), .D(n_308321970
		), .Z(n_310068899));
	notech_nor2 i_75844633(.A(n_341669189), .B(nbus_11326[27]), .Z(n_310168900
		));
	notech_or4 i_75344638(.A(n_56203), .B(n_56086), .C(n_54367), .D(n_308221969
		), .Z(n_310868907));
	notech_nor2 i_76644625(.A(n_341669189), .B(nbus_11326[28]), .Z(n_310968908
		));
	notech_or2 i_76144630(.A(n_326769066), .B(\nbus_11276[28] ), .Z(n_311668915
		));
	notech_nor2 i_87044523(.A(n_56057), .B(\nbus_11276[28] ), .Z(n_312168920
		));
	notech_nao3 i_100544398(.A(n_54520), .B(n_59826), .C(n_55334), .Z(n_312268921
		));
	notech_ao4 i_188243551(.A(n_27551), .B(n_59826), .C(n_57330), .D(n_101213406
		), .Z(n_312868927));
	notech_ao4 i_188143552(.A(n_101413408), .B(n_29219), .C(n_98113375), .D(nbus_11273
		[28]), .Z(n_313068929));
	notech_nao3 i_44245375(.A(n_312868927), .B(n_313068929), .C(n_312168920)
		, .Z(n_313168930));
	notech_ao4 i_180043633(.A(n_57330), .B(n_327069069), .C(n_55870), .D(n_307421961
		), .Z(n_313268931));
	notech_ao4 i_179943634(.A(n_29219), .B(n_26224), .C(n_326669065), .D(nbus_11273
		[28]), .Z(n_313468933));
	notech_nand3 i_180243631(.A(n_313268931), .B(n_313468933), .C(n_311668915
		), .Z(n_313568934));
	notech_ao4 i_179743636(.A(n_343565725), .B(n_341569188), .C(n_57306), .D
		(n_341769190), .Z(n_313668935));
	notech_ao4 i_179343640(.A(n_286061878), .B(n_341569188), .C(n_303621923)
		, .D(n_55870), .Z(n_313968938));
	notech_ao4 i_179243641(.A(n_29154), .B(n_26224), .C(n_308621973), .D(n_327069069
		), .Z(n_314168940));
	notech_nand3 i_179543638(.A(n_313968938), .B(n_314168940), .C(n_310868907
		), .Z(n_314268941));
	notech_ao4 i_179043643(.A(n_326669065), .B(nbus_11273[27]), .C(n_326769066
		), .D(\nbus_11276[27] ), .Z(n_314368942));
	notech_ao4 i_178643647(.A(n_288561889), .B(n_341569188), .C(n_55870), .D
		(n_307621963), .Z(n_314668945));
	notech_ao4 i_178543648(.A(n_29156), .B(n_26224), .C(n_308721974), .D(n_327069069
		), .Z(n_314868947));
	notech_nand3 i_178843645(.A(n_314668945), .B(n_314868947), .C(n_310068899
		), .Z(n_314968948));
	notech_ao4 i_178343650(.A(n_326669065), .B(nbus_11273[26]), .C(n_326769066
		), .D(\nbus_11276[26] ), .Z(n_315068949));
	notech_ao4 i_177943654(.A(n_268264999), .B(n_341569188), .C(n_307521962)
		, .D(n_55870), .Z(n_315368952));
	notech_ao4 i_177843655(.A(n_29215), .B(n_26224), .C(n_308821975), .D(n_327069069
		), .Z(n_315568954));
	notech_nand3 i_178143652(.A(n_315368952), .B(n_315568954), .C(n_309268891
		), .Z(n_315668955));
	notech_ao4 i_177543657(.A(n_326669065), .B(nbus_11273[25]), .C(n_326769066
		), .D(\nbus_11276[25] ), .Z(n_315768956));
	notech_ao4 i_177143661(.A(n_308521972), .B(n_341769190), .C(n_270765024)
		, .D(n_341569188), .Z(n_316068959));
	notech_ao4 i_177043662(.A(n_29152), .B(n_26224), .C(n_27590), .D(n_326869067
		), .Z(n_316268961));
	notech_nand3 i_177343659(.A(n_316068959), .B(n_316268961), .C(n_308468883
		), .Z(n_316368962));
	notech_ao4 i_176843664(.A(n_326669065), .B(nbus_11273[23]), .C(n_326769066
		), .D(\nbus_11276[23] ), .Z(n_316468963));
	notech_and4 i_99541275(.A(n_56061), .B(n_293761941), .C(n_293161935), .D
		(n_55975), .Z(n_316768966));
	notech_nor2 i_69841559(.A(n_341669189), .B(nbus_11326[18]), .Z(n_316868967
		));
	notech_or2 i_69341564(.A(n_311318890), .B(n_327069069), .Z(n_317568974)
		);
	notech_nor2 i_70641551(.A(n_341669189), .B(nbus_11326[19]), .Z(n_317668975
		));
	notech_or2 i_70141556(.A(n_311218889), .B(n_327069069), .Z(n_318368982)
		);
	notech_nor2 i_71441543(.A(n_341669189), .B(nbus_11326[20]), .Z(n_318468983
		));
	notech_or2 i_70941548(.A(n_311118888), .B(n_327069069), .Z(n_319168990)
		);
	notech_nor2 i_72241535(.A(n_341669189), .B(nbus_11326[21]), .Z(n_319268991
		));
	notech_or2 i_71741540(.A(n_311018887), .B(n_327069069), .Z(n_319968998)
		);
	notech_or2 i_73041527(.A(n_341669189), .B(nbus_11326[22]), .Z(n_320068999
		));
	notech_or2 i_72541532(.A(n_26618), .B(n_327069069), .Z(n_320769006));
	notech_ao4 i_178740505(.A(n_310418881), .B(n_341769190), .C(n_305565372)
		, .D(n_341569188), .Z(n_321169010));
	notech_ao4 i_178640506(.A(n_29174), .B(n_26224), .C(n_326869067), .D(n_27589
		), .Z(n_321369012));
	notech_and3 i_178940503(.A(n_321169010), .B(n_321369012), .C(n_320769006
		), .Z(n_321469013));
	notech_ao4 i_178440508(.A(n_326669065), .B(nbus_11273[22]), .C(n_326769066
		), .D(\nbus_11276[22] ), .Z(n_321569014));
	notech_ao4 i_178040512(.A(n_310518882), .B(n_341769190), .C(n_312662130)
		, .D(n_341569188), .Z(n_321869017));
	notech_ao4 i_177940513(.A(n_29172), .B(n_26224), .C(n_326869067), .D(n_27588
		), .Z(n_322069019));
	notech_nand3 i_178240510(.A(n_321869017), .B(n_322069019), .C(n_319968998
		), .Z(n_322169020));
	notech_ao4 i_177740515(.A(n_326669065), .B(nbus_11273[21]), .C(n_326769066
		), .D(\nbus_11276[21] ), .Z(n_322269021));
	notech_ao4 i_177340519(.A(n_310618883), .B(n_341769190), .C(n_315162155)
		, .D(n_341569188), .Z(n_322569024));
	notech_ao4 i_177240520(.A(n_29169), .B(n_26224), .C(n_326869067), .D(n_27586
		), .Z(n_322769026));
	notech_nand3 i_177540517(.A(n_322569024), .B(n_322769026), .C(n_319168990
		), .Z(n_322869027));
	notech_ao4 i_177040522(.A(n_326669065), .B(nbus_11273[20]), .C(n_326769066
		), .D(\nbus_11276[20] ), .Z(n_322969028));
	notech_ao4 i_176640526(.A(n_310718884), .B(n_341769190), .C(n_308065397)
		, .D(n_341569188), .Z(n_323269031));
	notech_ao4 i_176540527(.A(n_29167), .B(n_26224), .C(n_326869067), .D(n_27585
		), .Z(n_323469033));
	notech_nand3 i_176840524(.A(n_323269031), .B(n_323469033), .C(n_318368982
		), .Z(n_323569034));
	notech_ao4 i_176340529(.A(n_326669065), .B(nbus_11273[19]), .C(n_326769066
		), .D(\nbus_11276[19] ), .Z(n_323669035));
	notech_ao4 i_175940533(.A(n_310818885), .B(n_341769190), .C(n_310565422)
		, .D(n_341569188), .Z(n_323969038));
	notech_ao4 i_175840534(.A(n_29165), .B(n_26224), .C(n_326869067), .D(n_27584
		), .Z(n_324169040));
	notech_nand3 i_176140531(.A(n_323969038), .B(n_324169040), .C(n_317568974
		), .Z(n_324269041));
	notech_ao4 i_175640536(.A(n_326669065), .B(nbus_11273[18]), .C(n_326769066
		), .D(\nbus_11276[18] ), .Z(n_324369042));
	notech_nao3 i_24557903(.A(n_56463), .B(instrc[119]), .C(n_355988238), .Z
		(n_324669045));
	notech_and3 i_4839044(.A(n_56061), .B(n_324869047), .C(n_203967859), .Z(n_324769046
		));
	notech_and3 i_90560581(.A(n_56058), .B(n_203767857), .C(n_201567835), .Z
		(n_324869047));
	notech_and2 i_36457927(.A(n_56061), .B(n_203967859), .Z(n_324969048));
	notech_or2 i_131257964(.A(n_54525), .B(n_340469177), .Z(n_326669065));
	notech_or4 i_131357963(.A(n_1913), .B(n_204067860), .C(n_340469177), .D(n_60530
		), .Z(n_326769066));
	notech_or2 i_62957984(.A(n_56375), .B(n_56009), .Z(n_326869067));
	notech_nand2 i_96239120(.A(n_54460), .B(n_340269175), .Z(n_326969068));
	notech_and2 i_96339121(.A(n_54457), .B(n_340369176), .Z(n_327069069));
	notech_or4 i_93338204(.A(n_56203), .B(n_56086), .C(n_56375), .D(n_27582)
		, .Z(n_327369072));
	notech_or2 i_93738202(.A(n_341669189), .B(nbus_11326[16]), .Z(n_327469073
		));
	notech_and2 i_93638203(.A(n_326969068), .B(\regs_13_14[16] ), .Z(n_327569074
		));
	notech_ao3 i_94138199(.A(opc_10[16]), .B(n_62419), .C(n_341569188), .Z(n_327669075
		));
	notech_nor2 i_94038200(.A(n_272088735), .B(n_341769190), .Z(n_327769076)
		);
	notech_nor2 i_93938201(.A(n_327069069), .B(n_271988736), .Z(n_327869077)
		);
	notech_or4 i_1720828(.A(n_324476083), .B(n_340976246), .C(n_327869077), 
		.D(n_342369196), .Z(n_19185));
	notech_or2 i_135260566(.A(n_324669045), .B(n_166567485), .Z(n_327969078)
		);
	notech_or2 i_132860572(.A(n_324669045), .B(n_324969048), .Z(n_328069079)
		);
	notech_nao3 i_95638185(.A(n_62411), .B(opc[14]), .C(n_327969078), .Z(n_328569084
		));
	notech_nao3 i_95738184(.A(opc_10[14]), .B(n_62399), .C(n_328069079), .Z(n_328669085
		));
	notech_nor2 i_95538186(.A(n_271888737), .B(n_54457), .Z(n_328769086));
	notech_nor2 i_95838183(.A(n_56009), .B(n_80913203), .Z(n_328869087));
	notech_or4 i_1520826(.A(n_5990), .B(n_328769086), .C(n_26233), .D(n_328869087
		), .Z(n_19173));
	notech_nor2 i_126037891(.A(n_354969318), .B(n_271988736), .Z(n_328969088
		));
	notech_ao3 i_126237889(.A(opc_10[16]), .B(n_62399), .C(n_113113525), .Z(n_329669095
		));
	notech_nor2 i_126137890(.A(n_354569315), .B(n_272088735), .Z(n_329769096
		));
	notech_or4 i_1721308(.A(n_329669095), .B(n_343669209), .C(n_329769096), 
		.D(n_328969088), .Z(n_20697));
	notech_nor2 i_129637855(.A(n_355488242), .B(n_2700), .Z(n_329869097));
	notech_ao3 i_129837853(.A(opc_10[17]), .B(n_62403), .C(n_353788271), .Z(n_330369102
		));
	notech_nor2 i_129437857(.A(n_271688739), .B(nbus_11273[17]), .Z(n_330869107
		));
	notech_or4 i_1821565(.A(n_330869107), .B(n_344769219), .C(n_329869097), 
		.D(n_26234), .Z(n_16452));
	notech_nor2 i_132037832(.A(n_355488242), .B(n_271988736), .Z(n_330969108
		));
	notech_nand2 i_131537837(.A(sav_esi[16]), .B(n_60591), .Z(n_331469113)
		);
	notech_or2 i_131937833(.A(n_55133), .B(nbus_11326[16]), .Z(n_331569114)
		);
	notech_or2 i_131637836(.A(n_355688241), .B(n_29004), .Z(n_331669115));
	notech_ao3 i_132237830(.A(opc_10[16]), .B(n_62413), .C(n_353788271), .Z(n_331969118
		));
	notech_nor2 i_132137831(.A(n_355788240), .B(n_272088735), .Z(n_332069119
		));
	notech_or4 i_1721564(.A(n_331969118), .B(n_345769229), .C(n_332069119), 
		.D(n_330969108), .Z(n_16446));
	notech_or2 i_134237810(.A(n_340769180), .B(n_271888737), .Z(n_332169120)
		);
	notech_or4 i_119155297(.A(n_56463), .B(instrc[119]), .C(n_2145), .D(n_222568044
		), .Z(n_332269121));
	notech_or4 i_355291(.A(n_56463), .B(n_2145), .C(n_55829), .D(instrc[119]
		), .Z(n_332369122));
	notech_or4 i_134337809(.A(n_273588720), .B(n_56121), .C(n_2240), .D(n_272188734
		), .Z(n_333269131));
	notech_and4 i_1521562(.A(n_333269131), .B(n_346669238), .C(n_346869240),
		 .D(n_332169120), .Z(n_16434));
	notech_nand3 i_135460565(.A(n_56492), .B(n_268064997), .C(n_166467484), 
		.Z(n_333569134));
	notech_nand3 i_137360563(.A(n_56492), .B(n_268064997), .C(n_55970), .Z(n_333669135
		));
	notech_or2 i_149137664(.A(n_54853), .B(n_29006), .Z(n_333769136));
	notech_or2 i_149437661(.A(n_55725), .B(n_27579), .Z(n_334069139));
	notech_ao3 i_149637659(.A(n_62411), .B(opc[14]), .C(n_333569134), .Z(n_334169140
		));
	notech_nao3 i_149737658(.A(opc_10[14]), .B(n_62403), .C(n_333669135), .Z
		(n_334269141));
	notech_nor2 i_149537660(.A(n_54852), .B(n_271888737), .Z(n_334369142));
	notech_nor2 i_149837657(.A(n_55898), .B(n_80913203), .Z(n_334469143));
	notech_or4 i_1521850(.A(n_334369142), .B(n_347569247), .C(n_5990), .D(n_334469143
		), .Z(n_12485));
	notech_and4 i_92039160(.A(n_339969172), .B(n_339869171), .C(n_339469167)
		, .D(n_339769170), .Z(n_57349));
	notech_nand2 i_183537322(.A(n_272388732), .B(opb[9]), .Z(n_334569144));
	notech_nand2 i_182937328(.A(add_src[9]), .B(n_26579), .Z(n_338269155));
	notech_or2 i_183037327(.A(n_57349), .B(n_2320), .Z(n_338369156));
	notech_nor2 i_183337324(.A(n_89513289), .B(n_27593), .Z(n_338669159));
	notech_nao3 i_183437323(.A(imm[41]), .B(n_26795), .C(n_2198), .Z(n_338769160
		));
	notech_and4 i_1016179(.A(n_338769160), .B(n_349169263), .C(n_349069262),
		 .D(n_334569144), .Z(n_14146));
	notech_ao4 i_19138902(.A(n_56240), .B(n_27724), .C(n_2261), .D(n_29265),
		 .Z(n_338869161));
	notech_ao4 i_19238901(.A(n_56178), .B(n_27994), .C(n_27827), .D(n_197114365
		), .Z(n_338969162));
	notech_ao4 i_19338900(.A(n_56414), .B(n_27962), .C(n_57343), .D(n_27756)
		, .Z(n_339169164));
	notech_ao4 i_19438899(.A(n_56182), .B(n_27928), .C(n_56310), .D(n_27615)
		, .Z(n_339269165));
	notech_and4 i_20338890(.A(n_339269165), .B(n_339169164), .C(n_338969162)
		, .D(n_338869161), .Z(n_339469167));
	notech_ao4 i_19538898(.A(n_60484), .B(n_27896), .C(n_56183), .D(n_29264)
		, .Z(n_339569168));
	notech_ao4 i_19638897(.A(n_56186), .B(n_27859), .C(n_56290), .D(n_27650)
		, .Z(n_339669169));
	notech_and2 i_20138892(.A(n_339669169), .B(n_339569168), .Z(n_339769170)
		);
	notech_ao4 i_19738896(.A(n_59224), .B(n_28028), .C(n_56270), .D(n_27692)
		, .Z(n_339869171));
	notech_ao4 i_19838895(.A(n_2262), .B(n_27795), .C(n_57371), .D(n_27379),
		 .Z(n_339969172));
	notech_or2 i_86260686(.A(n_324869047), .B(n_54525), .Z(n_340269175));
	notech_or4 i_86360685(.A(n_1913), .B(n_204067860), .C(n_324869047), .D(n_60532
		), .Z(n_340369176));
	notech_ao4 i_35257994(.A(n_56502), .B(n_54520), .C(n_56375), .D(n_26250)
		, .Z(n_340469177));
	notech_and3 i_105055340(.A(n_323731624), .B(n_317488515), .C(n_55791), .Z
		(n_340569178));
	notech_and4 i_104955341(.A(n_55222), .B(n_319188498), .C(n_317288517), .D
		(n_55790), .Z(n_340669179));
	notech_ao4 i_93355348(.A(n_54874), .B(n_56104), .C(n_55829), .D(n_320788482
		), .Z(n_340769180));
	notech_ao4 i_93255349(.A(n_1970), .B(n_60473), .C(n_317888511), .D(n_55829
		), .Z(n_340869181));
	notech_and2 i_57455361(.A(n_55688), .B(n_319988490), .Z(n_340969182));
	notech_and2 i_95060676(.A(n_340369176), .B(n_326769066), .Z(n_341269185)
		);
	notech_and2 i_94960677(.A(n_326669065), .B(n_340269175), .Z(n_341369186)
		);
	notech_and2 i_60160703(.A(n_326869067), .B(n_166767487), .Z(n_341469187)
		);
	notech_or2 i_27925(.A(n_324669045), .B(n_324769046), .Z(n_341569188));
	notech_or4 i_27931(.A(n_1976), .B(n_355988238), .C(n_340469177), .D(n_60511
		), .Z(n_341669189));
	notech_or2 i_27937(.A(n_56009), .B(n_54367), .Z(n_341769190));
	notech_ao4 i_94238198(.A(n_326769066), .B(\nbus_11276[16] ), .C(nbus_11273
		[16]), .D(n_326669065), .Z(n_341869191));
	notech_nand3 i_94438196(.A(n_327369072), .B(n_341869191), .C(n_327469073
		), .Z(n_342069193));
	notech_or4 i_94738193(.A(n_327569074), .B(n_342069193), .C(n_327669075),
		 .D(n_327769076), .Z(n_342369196));
	notech_ao4 i_95938182(.A(n_341269185), .B(\nbus_11276[14] ), .C(n_54460)
		, .D(n_29006), .Z(n_342569198));
	notech_ao4 i_96038181(.A(n_341469187), .B(n_27579), .C(n_341369186), .D(nbus_11273
		[14]), .Z(n_342669199));
	notech_and4 i_96538178(.A(n_342669199), .B(n_342569198), .C(n_328569084)
		, .D(n_328669085), .Z(n_342969202));
	notech_ao4 i_126537886(.A(n_55776), .B(n_27582), .C(n_2193), .D(n_27535)
		, .Z(n_343269205));
	notech_ao4 i_126337888(.A(n_55562), .B(nbus_11273[16]), .C(n_113313527),
		 .D(nbus_11326[16]), .Z(n_343369206));
	notech_ao4 i_126437887(.A(n_29004), .B(n_26571), .C(n_354669316), .D(\nbus_11276[16] 
		), .Z(n_343469207));
	notech_nand3 i_126737884(.A(n_343469207), .B(n_343369206), .C(n_343269205
		), .Z(n_343669209));
	notech_ao4 i_130637845(.A(n_271588740), .B(\nbus_11276[17] ), .C(n_355688241
		), .D(n_28987), .Z(n_343969212));
	notech_ao4 i_129937852(.A(n_321788473), .B(n_29280), .C(n_321688474), .D
		(n_29279), .Z(n_344069213));
	notech_ao4 i_130037851(.A(n_59186), .B(n_26726), .C(n_320088489), .D(n_27583
		), .Z(n_344169214));
	notech_and3 i_130237849(.A(n_344169214), .B(n_344069213), .C(n_355888239
		), .Z(n_344469216));
	notech_ao4 i_130437847(.A(n_55133), .B(nbus_11326[17]), .C(n_355788240),
		 .D(n_2648), .Z(n_344669218));
	notech_nao3 i_130537846(.A(n_344669218), .B(n_344469216), .C(n_330369102
		), .Z(n_344769219));
	notech_ao4 i_132437828(.A(n_320088489), .B(n_27582), .C(n_59163), .D(n_27535
		), .Z(n_345069222));
	notech_ao4 i_132337829(.A(n_321788473), .B(n_29282), .C(n_321688474), .D
		(n_29281), .Z(n_345169223));
	notech_and4 i_132737825(.A(n_345169223), .B(n_345069222), .C(n_331469113
		), .D(n_331569114), .Z(n_345469226));
	notech_ao4 i_132937823(.A(n_271688739), .B(nbus_11273[16]), .C(n_271588740
		), .D(\nbus_11276[16] ), .Z(n_345669228));
	notech_nand3 i_133037822(.A(n_345469226), .B(n_345669228), .C(n_331669115
		), .Z(n_345769229));
	notech_ao4 i_134637806(.A(n_321788473), .B(n_29284), .C(n_321688474), .D
		(n_29283), .Z(n_346069232));
	notech_ao4 i_134737805(.A(n_340569178), .B(\nbus_11276[14] ), .C(n_340869181
		), .D(n_29006), .Z(n_346169233));
	notech_ao4 i_134837804(.A(n_340969182), .B(n_27579), .C(n_340669179), .D
		(nbus_11273[14]), .Z(n_346369235));
	notech_ao4 i_134937803(.A(n_59186), .B(n_26725), .C(n_59163), .D(n_27533
		), .Z(n_346469236));
	notech_and4 i_135237800(.A(n_346469236), .B(n_346369235), .C(n_346169233
		), .D(n_346069232), .Z(n_346669238));
	notech_ao4 i_135437798(.A(n_82713221), .B(n_332369122), .C(n_82813222), 
		.D(n_332269121), .Z(n_346869240));
	notech_ao4 i_150037655(.A(n_54946), .B(nbus_11273[14]), .C(n_54945), .D(\nbus_11276[14] 
		), .Z(n_347069242));
	notech_and4 i_150237653(.A(n_55901), .B(n_347069242), .C(n_333769136), .D
		(n_334069139), .Z(n_347369245));
	notech_nao3 i_150437651(.A(n_347369245), .B(n_334269141), .C(n_334169140
		), .Z(n_347569247));
	notech_ao4 i_183937318(.A(n_55243), .B(n_27528), .C(n_2164), .D(nbus_11326
		[9]), .Z(n_347869250));
	notech_ao4 i_184037317(.A(n_55526), .B(n_28591), .C(n_55366), .D(n_28783
		), .Z(n_347969251));
	notech_ao4 i_183637321(.A(n_54884), .B(\nbus_11276[25] ), .C(n_54735), .D
		(nbus_11326[1]), .Z(n_348169253));
	notech_ao4 i_183737320(.A(n_2156), .B(n_28810), .C(n_2323), .D(n_27574),
		 .Z(n_348369255));
	notech_ao4 i_183837319(.A(n_2319), .B(n_29024), .C(n_2322), .D(nbus_11273
		[9]), .Z(n_348469256));
	notech_and4 i_184437313(.A(n_348469256), .B(n_348369255), .C(n_348169253
		), .D(n_338269155), .Z(n_348669258));
	notech_and4 i_184637311(.A(n_347969251), .B(n_347869250), .C(n_348669258
		), .D(n_36812763), .Z(n_348869260));
	notech_ao3 i_184937308(.A(n_348869260), .B(n_338369156), .C(n_338669159)
		, .Z(n_349069262));
	notech_ao4 i_184837309(.A(n_88913283), .B(n_28839), .C(n_88813282), .D(n_28410
		), .Z(n_349169263));
	notech_ao4 i_220433565(.A(n_57343), .B(n_27748), .C(n_59224), .D(n_28020
		), .Z(n_351069282));
	notech_ao4 i_220333566(.A(n_56270), .B(n_27682), .C(n_57371), .D(n_27371
		), .Z(n_351169283));
	notech_ao4 i_220133568(.A(n_56290), .B(n_27640), .C(n_56186), .D(n_27851
		), .Z(n_351369285));
	notech_ao4 i_220033569(.A(n_56183), .B(n_27560), .C(n_60484), .D(n_27886
		), .Z(n_351469286));
	notech_and4 i_220633563(.A(n_351469286), .B(n_351369285), .C(n_351169283
		), .D(n_351069282), .Z(n_351669288));
	notech_ao4 i_219733572(.A(n_56310), .B(n_27605), .C(n_56182), .D(n_27920
		), .Z(n_351769289));
	notech_ao4 i_219633573(.A(n_56178), .B(n_27986), .C(n_56414), .D(n_27954
		), .Z(n_351869290));
	notech_and2 i_219833571(.A(n_351869290), .B(n_351769289), .Z(n_351969291
		));
	notech_ao4 i_219433575(.A(n_2262), .B(n_27787), .C(n_197114365), .D(n_27819
		), .Z(n_352069292));
	notech_ao4 i_219333576(.A(n_2261), .B(n_29266), .C(n_56240), .D(n_27716)
		, .Z(n_352169293));
	notech_and2 i_88432884(.A(n_55961), .B(n_55959), .Z(n_352469296));
	notech_or2 i_54032440(.A(n_57374), .B(eval_flag), .Z(n_352569297));
	notech_or4 i_10468305(.A(n_1909), .B(n_28567), .C(n_60532), .D(n_26597),
		 .Z(n_28442003));
	notech_and4 i_10668304(.A(n_56186), .B(n_56310), .C(n_56414), .D(n_56178
		), .Z(n_27641995));
	notech_nand3 i_19268293(.A(n_56186), .B(n_56414), .C(n_127467094), .Z(n_27341992
		));
	notech_ao4 i_150153856(.A(n_59186), .B(n_26700), .C(n_57293), .D(n_320465521
		), .Z(n_194164276));
	notech_nand3 i_420655(.A(n_148867308), .B(n_148767307), .C(n_149267312),
		 .Z(n_19803));
	notech_and4 i_320654(.A(n_146967289), .B(n_201867838), .C(n_149767317), 
		.D(n_149667316), .Z(n_19797));
	notech_and4 i_220653(.A(n_146167281), .B(n_201767837), .C(n_150467324), 
		.D(n_150367323), .Z(n_19791));
	notech_nand3 i_420719(.A(n_150967329), .B(n_150867328), .C(n_151367333),
		 .Z(n_19455));
	notech_and4 i_320718(.A(n_151467334), .B(n_151667336), .C(n_145367273), 
		.D(n_152067340), .Z(n_19449));
	notech_and4 i_220717(.A(n_201767837), .B(n_152567345), .C(n_143867258), 
		.D(n_152467344), .Z(n_19443));
	notech_and4 i_720818(.A(n_152867348), .B(n_153067350), .C(n_153467354), 
		.D(n_143767257), .Z(n_19125));
	notech_and4 i_520816(.A(n_153567355), .B(n_153767357), .C(n_154167361), 
		.D(n_142967249), .Z(n_19113));
	notech_nand3 i_420815(.A(n_154467364), .B(n_154367363), .C(n_154867368),
		 .Z(n_19107));
	notech_and4 i_320814(.A(n_201867838), .B(n_155367373), .C(n_140767227), 
		.D(n_155267372), .Z(n_19101));
	notech_nand3 i_420943(.A(n_155867378), .B(n_155767377), .C(n_156267382),
		 .Z(n_8997));
	notech_and4 i_320942(.A(n_156367383), .B(n_156567385), .C(n_139967219), 
		.D(n_156967389), .Z(n_8991));
	notech_and4 i_220941(.A(n_201767837), .B(n_157467394), .C(n_138467204), 
		.D(n_157367393), .Z(n_8985));
	notech_and4 i_320974(.A(n_157767397), .B(n_157967399), .C(n_158467404), 
		.D(n_138367203), .Z(n_16711));
	notech_and4 i_220973(.A(n_158567405), .B(n_158767407), .C(n_159267412), 
		.D(n_137467194), .Z(n_16705));
	notech_nand3 i_421039(.A(n_159567415), .B(n_159467414), .C(n_159967419),
		 .Z(n_13833));
	notech_and4 i_321038(.A(n_160067420), .B(n_160267422), .C(n_135867178), 
		.D(n_160667426), .Z(n_13827));
	notech_and4 i_221037(.A(n_201767837), .B(n_161167431), .C(n_134367163), 
		.D(n_161067430), .Z(n_13821));
	notech_nand2 i_421167(.A(n_162367443), .B(n_161867438), .Z(n_13485));
	notech_nand3 i_421583(.A(n_162667446), .B(n_162567445), .C(n_163067450),
		 .Z(n_13133));
	notech_and4 i_321582(.A(n_201867838), .B(n_163567455), .C(n_131767137), 
		.D(n_163467454), .Z(n_13127));
	notech_and4 i_221581(.A(n_201767837), .B(n_164267462), .C(n_130967129), 
		.D(n_164167461), .Z(n_13121));
	notech_and4 i_321902(.A(n_164967469), .B(n_165167471), .C(n_130367123), 
		.D(n_164867468), .Z(n_12061));
	notech_and4 i_221901(.A(n_165767477), .B(n_165967479), .C(n_129467114), 
		.D(n_165667476), .Z(n_12055));
	notech_and4 i_6163486(.A(n_56061), .B(n_293761941), .C(n_55973), .D(n_293161935
		), .Z(n_273539523));
	notech_and4 i_150953848(.A(n_193864273), .B(n_193664271), .C(n_193564270
		), .D(n_188964224), .Z(n_194064275));
	notech_and3 i_10263445(.A(n_97522962), .B(n_355976395), .C(n_54431), .Z(n_269539483
		));
	notech_and3 i_10363444(.A(n_55072), .B(n_45384), .C(n_54454), .Z(n_269439482
		));
	notech_ao4 i_150453853(.A(n_55520), .B(n_29087), .C(n_356476400), .D(n_55519
		), .Z(n_193864273));
	notech_ao3 i_10463443(.A(n_55073), .B(n_54453), .C(n_45383), .Z(n_269339481
		));
	notech_and2 i_11163437(.A(n_54455), .B(n_128967109), .Z(n_268739475));
	notech_ao4 i_150653851(.A(n_55382), .B(nbus_11273[15]), .C(n_55381), .D(\nbus_11276[15] 
		), .Z(n_193664271));
	notech_ao4 i_150753850(.A(n_177164109), .B(n_320565522), .C(n_320665523)
		, .D(n_177264110), .Z(n_193564270));
	notech_and2 i_62560698(.A(n_55772), .B(n_166667486), .Z(n_55725));
	notech_ao3 i_147460658(.A(n_54749), .B(n_55220), .C(n_47685), .Z(n_54946
		));
	notech_and3 i_147560657(.A(n_47687), .B(n_54695), .C(n_55221), .Z(n_54945
		));
	notech_or2 i_209260615(.A(n_56006), .B(n_54528), .Z(n_54436));
	notech_or4 i_209760614(.A(n_997), .B(n_56006), .C(n_1909), .D(n_2202), .Z
		(n_54432));
	notech_and2 i_222453139(.A(n_295765274), .B(n_189564230), .Z(n_193164266
		));
	notech_or4 i_11859(.A(n_1909), .B(n_2202), .C(n_997), .D(n_263136786), .Z
		(n_45384));
	notech_nor2 i_11860(.A(n_54528), .B(n_263136786), .Z(n_45383));
	notech_ao4 i_223253131(.A(n_54439), .B(n_29205), .C(n_56151), .D(n_27621
		), .Z(n_192664261));
	notech_ao4 i_223353130(.A(n_54451), .B(n_27658), .C(n_56097), .D(n_27698
		), .Z(n_192564260));
	notech_and2 i_223753126(.A(n_192364258), .B(n_192264257), .Z(n_192464259
		));
	notech_ao4 i_223553128(.A(n_54535), .B(n_27385), .C(n_55864), .D(n_27730
		), .Z(n_192364258));
	notech_and4 i_3020841(.A(n_262736782), .B(n_185667676), .C(n_182967649),
		 .D(n_185567675), .Z(n_19263));
	notech_or4 i_1020821(.A(n_185167671), .B(n_182267642), .C(n_186267682), 
		.D(n_26202), .Z(n_19143));
	notech_and4 i_920820(.A(n_186667686), .B(n_186867688), .C(n_182167641), 
		.D(n_187267692), .Z(n_19137));
	notech_nand2 i_321166(.A(n_188267702), .B(n_187767697), .Z(n_13479));
	notech_nand2 i_221165(.A(n_189267712), .B(n_188767707), .Z(n_13473));
	notech_and4 i_1021557(.A(n_189967719), .B(n_189867718), .C(n_178467604),
		 .D(n_190267722), .Z(n_16404));
	notech_and4 i_421551(.A(n_191067730), .B(n_191767737), .C(n_190967729), 
		.D(n_176867588), .Z(n_16368));
	notech_or4 i_321550(.A(n_175667576), .B(n_192867748), .C(n_26195), .D(n_26197
		), .Z(n_16362));
	notech_or4 i_221549(.A(n_174467564), .B(n_193967759), .C(n_26192), .D(n_26193
		), .Z(n_16356));
	notech_nand3 i_1021589(.A(n_194367763), .B(n_194267762), .C(n_194767767)
		, .Z(n_13169));
	notech_and4 i_921844(.A(n_194867768), .B(n_195067770), .C(n_195567775), 
		.D(n_173267552), .Z(n_12449));
	notech_nand3 i_421839(.A(n_195967779), .B(n_195867778), .C(n_196367783),
		 .Z(n_12419));
	notech_and4 i_717233(.A(n_196967789), .B(n_197167791), .C(n_196867788), 
		.D(n_171167531), .Z(n_15810));
	notech_and4 i_517231(.A(n_197867798), .B(n_197767797), .C(n_170167521), 
		.D(n_198067800), .Z(n_15798));
	notech_nand2 i_417230(.A(n_199167811), .B(n_198767807), .Z(n_15792));
	notech_nand2 i_317229(.A(n_200167821), .B(n_199667816), .Z(n_15786));
	notech_nand2 i_217228(.A(n_201167831), .B(n_200667826), .Z(n_15780));
	notech_or4 i_39260599(.A(n_59263), .B(n_59272), .C(n_56121), .D(n_54089)
		, .Z(n_263036785));
	notech_ao4 i_122660575(.A(nbus_11273[9]), .B(n_54698), .C(n_1970), .D(n_29048
		), .Z(n_260636761));
	notech_ao4 i_223653127(.A(n_55898), .B(n_27764), .C(n_55940), .D(n_27801
		), .Z(n_192264257));
	notech_and4 i_224553118(.A(n_191964254), .B(n_191864253), .C(n_191664251
		), .D(n_191564250), .Z(n_192164256));
	notech_ao4 i_223953124(.A(n_55867), .B(n_27833), .C(n_56068), .D(n_27866
		), .Z(n_191964254));
	notech_ao4 i_224053123(.A(n_56035), .B(n_27902), .C(n_56009), .D(n_27934
		), .Z(n_191864253));
	notech_ao4 i_224253121(.A(n_55998), .B(n_27968), .C(n_55872), .D(n_28000
		), .Z(n_191664251));
	notech_ao4 i_224353120(.A(n_55873), .B(n_29206), .C(n_55878), .D(n_28034
		), .Z(n_191564250));
	notech_or2 i_73657976(.A(n_54505), .B(n_250234128), .Z(n_55614));
	notech_ao3 i_150657959(.A(n_54902), .B(n_55219), .C(n_46842), .Z(n_54921
		));
	notech_and3 i_150757958(.A(n_46844), .B(n_54872), .C(n_55218), .Z(n_54920
		));
	notech_or2 i_206357946(.A(n_54525), .B(n_324969048), .Z(n_54460));
	notech_or4 i_206757944(.A(n_1913), .B(n_204067860), .C(n_60532), .D(n_324969048
		), .Z(n_54457));
	notech_and4 i_251757940(.A(n_56061), .B(n_203967859), .C(n_201567835), .D
		(n_340469177), .Z(n_54071));
	notech_and4 i_251957939(.A(n_56060), .B(n_996), .C(n_56000), .D(n_55988)
		, .Z(n_54069));
	notech_or2 i_137657861(.A(n_55975), .B(n_294261946), .Z(n_248434110));
	notech_or2 i_11202(.A(n_55580), .B(n_55873), .Z(n_46041));
	notech_or4 i_28993(.A(n_56492), .B(instrc[118]), .C(n_2349), .D(n_56006)
		, .Z(n_254634172));
	notech_and2 i_198257930(.A(n_213667956), .B(n_56260), .Z(n_54525));
	notech_or2 i_202057926(.A(n_204067860), .B(n_56182), .Z(n_54494));
	notech_or4 i_206857925(.A(n_1913), .B(n_204067860), .C(n_202167841), .D(n_60532
		), .Z(n_54456));
	notech_or2 i_207557924(.A(n_54525), .B(n_202167841), .Z(n_54450));
	notech_and4 i_820819(.A(n_211867938), .B(n_214667966), .C(n_214867968), 
		.D(n_215267972), .Z(n_19131));
	notech_and4 i_220813(.A(n_201767837), .B(n_215767977), .C(n_210367923), 
		.D(n_215667976), .Z(n_19095));
	notech_and4 i_420975(.A(n_201667836), .B(n_216467984), .C(n_209567915), 
		.D(n_216367983), .Z(n_16717));
	notech_nand3 i_421295(.A(n_218168001), .B(n_218068000), .C(n_217967999),
		 .Z(n_20619));
	notech_nand2 i_321294(.A(n_219368013), .B(n_218868008), .Z(n_20613));
	notech_nand2 i_221293(.A(n_220268022), .B(n_219868018), .Z(n_20607));
	notech_and4 i_321838(.A(n_220368023), .B(n_220568025), .C(n_221068030), 
		.D(n_206067880), .Z(n_12413));
	notech_and4 i_221837(.A(n_221168031), .B(n_221368033), .C(n_221968038), 
		.D(n_205267872), .Z(n_12407));
	notech_ao4 i_73557880(.A(n_26591), .B(n_27019), .C(n_26189), .D(n_26231)
		, .Z(n_250334129));
	notech_and2 i_75157879(.A(n_55959), .B(n_55958), .Z(n_250234128));
	notech_and2 i_115757875(.A(n_55355), .B(n_202567845), .Z(n_249834124));
	notech_ao3 i_128157866(.A(n_55562), .B(n_26246), .C(n_209267912), .Z(n_248934115
		));
	notech_or2 i_190757852(.A(n_324669045), .B(n_202167841), .Z(n_247534101)
		);
	notech_or4 i_188355336(.A(instrc[118]), .B(n_229364616), .C(n_56469), .D
		(n_56032), .Z(n_54607));
	notech_nand2 i_195855335(.A(n_54607), .B(n_50635), .Z(n_54545));
	notech_and3 i_192555334(.A(n_55142), .B(n_222168040), .C(n_355188244), .Z
		(n_54572));
	notech_and3 i_192455333(.A(n_55143), .B(n_222268041), .C(n_355388243), .Z
		(n_54573));
	notech_or4 i_6602(.A(instrc[118]), .B(n_229364616), .C(n_56469), .D(n_222068039
		), .Z(n_50635));
	notech_or4 i_47355326(.A(fsm[3]), .B(fsm[0]), .C(n_60775), .D(n_249261520
		), .Z(n_55876));
	notech_or4 i_2520836(.A(n_252861556), .B(n_236968174), .C(n_239568200), 
		.D(n_26196), .Z(n_19233));
	notech_and4 i_1620827(.A(n_363088165), .B(n_240368208), .C(n_236168166),
		 .D(n_240268207), .Z(n_19179));
	notech_or4 i_1420825(.A(n_188774755), .B(n_235368158), .C(n_240968214), 
		.D(n_26198), .Z(n_19167));
	notech_or4 i_1320824(.A(n_189974767), .B(n_234268150), .C(n_242268221), 
		.D(n_26199), .Z(n_19161));
	notech_or4 i_1220823(.A(n_239168196), .B(n_233468142), .C(n_242968228), 
		.D(n_26200), .Z(n_19155));
	notech_and4 i_1120822(.A(n_154070859), .B(n_243768236), .C(n_232568134),
		 .D(n_243668235), .Z(n_19149));
	notech_nand2 i_1621563(.A(n_244968248), .B(n_244468243), .Z(n_16440));
	notech_nand2 i_1421561(.A(n_245968258), .B(n_245468253), .Z(n_16428));
	notech_nand2 i_1321560(.A(n_246968268), .B(n_246468263), .Z(n_16422));
	notech_nand2 i_1221559(.A(n_247968278), .B(n_247468273), .Z(n_16416));
	notech_and4 i_1121558(.A(n_248768286), .B(n_248668285), .C(n_248568284),
		 .D(n_249068289), .Z(n_16410));
	notech_nand2 i_921556(.A(n_250168300), .B(n_249668295), .Z(n_16398));
	notech_or4 i_1221847(.A(n_239168196), .B(n_223568054), .C(n_250568304), 
		.D(n_26201), .Z(n_12467));
	notech_nand2 i_1117237(.A(n_251768316), .B(n_251368312), .Z(n_15834));
	notech_or2 i_120054145(.A(n_54935), .B(n_177864116), .Z(n_189664231));
	notech_or2 i_119954146(.A(n_260961637), .B(n_177864116), .Z(n_189564230)
		);
	notech_nand2 i_26647(.A(opc_10[9]), .B(n_62413), .Z(n_352969301));
	notech_nand2 i_26648(.A(n_62411), .B(opc[9]), .Z(n_353069302));
	notech_mux2 i_1011667(.S(n_60136), .A(n_565), .B(add_len_pc32[9]), .Z(n_353169303
		));
	notech_nand2 i_26908(.A(opc_10[3]), .B(n_62403), .Z(n_353269304));
	notech_nand2 i_26909(.A(n_62429), .B(opc[3]), .Z(n_353369305));
	notech_nand2 i_26941(.A(opc_10[2]), .B(n_62403), .Z(n_353469306));
	notech_nand2 i_26942(.A(n_62411), .B(opc[2]), .Z(n_353569307));
	notech_nand2 i_26983(.A(opc_10[1]), .B(n_62401), .Z(n_353769308));
	notech_nand2 i_26984(.A(n_62411), .B(opc[1]), .Z(n_353869309));
	notech_and3 i_60952089(.A(n_2006), .B(n_55842), .C(n_55687), .Z(n_353969310
		));
	notech_nao3 i_97552075(.A(n_55236), .B(n_55567), .C(n_1897), .Z(n_354069311
		));
	notech_and3 i_97652074(.A(n_55216), .B(n_1898), .C(n_55568), .Z(n_354269312
		));
	notech_or4 i_26404(.A(n_56463), .B(n_2145), .C(n_55834), .D(n_29010), .Z
		(n_354369313));
	notech_or4 i_119251975(.A(n_56465), .B(n_2145), .C(n_259068389), .D(n_29010
		), .Z(n_354469314));
	notech_and2 i_54649259(.A(n_55685), .B(n_46041), .Z(n_354569315));
	notech_ao4 i_78949249(.A(n_55960), .B(n_54505), .C(n_54688), .D(n_2327),
		 .Z(n_354669316));
	notech_or4 i_87049242(.A(n_250334129), .B(n_284768646), .C(n_55831), .D(n_26206
		), .Z(n_354869317));
	notech_and3 i_87149241(.A(n_54722), .B(n_284468643), .C(n_55614), .Z(n_354969318
		));
	notech_or4 i_170049218(.A(n_212964463), .B(n_60532), .C(n_2739), .D(n_56032
		), .Z(n_355188244));
	notech_or2 i_170549217(.A(n_351565804), .B(n_56032), .Z(n_355388243));
	notech_or2 i_108449171(.A(n_2255), .B(n_284868647), .Z(n_113113525));
	notech_or4 i_140449163(.A(n_2145), .B(n_1976), .C(n_55960), .D(n_60511),
		 .Z(n_113313527));
	notech_or2 i_4445333(.A(n_2255), .B(n_307568874), .Z(n_302721914));
	notech_or4 i_141142238(.A(n_264436799), .B(n_231461383), .C(n_55973), .D
		(n_60511), .Z(n_308318860));
	notech_or2 i_54942250(.A(n_55523), .B(n_55864), .Z(n_309518872));
	notech_or2 i_108242242(.A(n_316768966), .B(n_294261946), .Z(n_308718864)
		);
	notech_and3 i_79642290(.A(n_46844), .B(n_54872), .C(n_54740), .Z(n_55554
		));
	notech_ao3 i_79542291(.A(n_54902), .B(n_54748), .C(n_46842), .Z(n_55555)
		);
	notech_ao4 i_90845403(.A(n_55960), .B(n_54505), .C(n_56057), .D(eval_flag
		), .Z(n_55447));
	notech_and3 i_110345404(.A(n_55527), .B(n_46073), .C(n_284468643), .Z(n_55269
		));
	notech_and3 i_110545405(.A(n_55528), .B(n_54760), .C(n_312268921), .Z(n_55267
		));
	notech_or2 i_82533096(.A(n_54530), .B(n_352469296), .Z(n_55528));
	notech_or2 i_82633168(.A(n_54505), .B(n_352469296), .Z(n_55527));
	notech_or4 i_2920840(.A(n_313168930), .B(n_310968908), .C(n_313568934), 
		.D(n_26215), .Z(n_19257));
	notech_or4 i_2820839(.A(n_264975488), .B(n_310168900), .C(n_314268941), 
		.D(n_26216), .Z(n_19251));
	notech_or4 i_2720838(.A(n_265975498), .B(n_309368892), .C(n_314968948), 
		.D(n_26217), .Z(n_19245));
	notech_or4 i_2620837(.A(n_173971058), .B(n_308568884), .C(n_315668955), 
		.D(n_26218), .Z(n_19239));
	notech_or4 i_2420835(.A(n_267675515), .B(n_307768876), .C(n_316368962), 
		.D(n_26219), .Z(n_19227));
	notech_or2 i_43445378(.A(n_56376), .B(n_27596), .Z(n_307421961));
	notech_or2 i_34254963(.A(n_55738), .B(n_27581), .Z(n_188964224));
	notech_and2 i_103533119(.A(n_2216), .B(n_352569297), .Z(n_55334));
	notech_or4 i_34554960(.A(n_59167), .B(n_26604), .C(n_26377), .D(n_27534)
		, .Z(n_188664221));
	notech_and4 i_2320834(.A(n_303675875), .B(n_321569014), .C(n_320068999),
		 .D(n_321469013), .Z(n_19221));
	notech_or4 i_2220833(.A(n_304775886), .B(n_319268991), .C(n_322169020), 
		.D(n_26220), .Z(n_19215));
	notech_or4 i_2120832(.A(n_320179591), .B(n_318468983), .C(n_322869027), 
		.D(n_26221), .Z(n_19209));
	notech_or4 i_2020831(.A(n_306575904), .B(n_317668975), .C(n_323569034), 
		.D(n_26222), .Z(n_19203));
	notech_or4 i_1920830(.A(n_320579595), .B(n_316868967), .C(n_324269041), 
		.D(n_26223), .Z(n_19197));
	notech_and3 i_91239138(.A(n_323731624), .B(n_317588514), .C(n_55979), .Z
		(n_355488242));
	notech_and4 i_91039137(.A(n_55222), .B(n_317388516), .C(n_55978), .D(n_319188498
		), .Z(n_355688241));
	notech_and3 i_56739134(.A(n_317088519), .B(n_55688), .C(n_319488495), .Z
		(n_355788240));
	notech_nand3 i_11572(.A(n_59186), .B(n_59927), .C(read_data[17]), .Z(n_355888239
		));
	notech_nand2 i_27917(.A(n_56492), .B(n_28967), .Z(n_355988238));
	notech_and4 i_91229141(.A(n_352169293), .B(n_352069292), .C(n_351669288)
		, .D(n_351969291), .Z(n_57357));
	notech_ao4 i_129433123(.A(n_54121), .B(n_27574), .C(n_55858), .D(n_57299
		), .Z(n_55085));
	notech_or2 i_34854957(.A(n_262636781), .B(n_26953), .Z(n_188364218));
	notech_ao4 i_83632883(.A(n_59370), .B(n_205588858), .C(n_57378), .D(eval_flag
		), .Z(n_2216));
	notech_or2 i_31654989(.A(n_55520), .B(n_29084), .Z(n_187664211));
	notech_or4 i_31954986(.A(n_59167), .B(n_26604), .C(n_26377), .D(n_27531)
		, .Z(n_187364208));
	notech_or2 i_32254983(.A(n_262636781), .B(n_26947), .Z(n_187064205));
	notech_or4 i_21755088(.A(n_56086), .B(n_56121), .C(n_56376), .D(n_27592)
		, .Z(n_186764202));
	notech_or2 i_22055085(.A(n_323065547), .B(\nbus_11276[24] ), .Z(n_186464199
		));
	notech_nand3 i_22355082(.A(n_1416), .B(tsc[56]), .C(n_59837), .Z(n_186164196
		));
	notech_or4 i_20855097(.A(n_57293), .B(n_55858), .C(n_56086), .D(n_56121)
		, .Z(n_185864193));
	notech_or2 i_21155094(.A(n_327465578), .B(\nbus_11276[15] ), .Z(n_185564190
		));
	notech_nand3 i_21455091(.A(n_1416), .B(tsc[47]), .C(n_59837), .Z(n_185264187
		));
	notech_nao3 i_19955106(.A(n_62411), .B(opc[13]), .C(n_324288256), .Z(n_184964184
		));
	notech_or2 i_20255103(.A(n_327465578), .B(\nbus_11276[13] ), .Z(n_184664181
		));
	notech_nand3 i_20555100(.A(n_1416), .B(tsc[45]), .C(n_59837), .Z(n_184364178
		));
	notech_nao3 i_19055115(.A(n_62433), .B(opc[12]), .C(n_324288256), .Z(n_184064175
		));
	notech_or2 i_19555110(.A(n_2662), .B(n_29084), .Z(n_183564170));
	notech_nand3 i_19655109(.A(n_1416), .B(tsc[44]), .C(n_59837), .Z(n_183264167
		));
	notech_nao3 i_18155124(.A(n_62411), .B(opc[11]), .C(n_324288256), .Z(n_183164166
		));
	notech_or2 i_18455121(.A(n_327465578), .B(\nbus_11276[11] ), .Z(n_182864163
		));
	notech_nand3 i_18755118(.A(n_1416), .B(tsc[43]), .C(n_59837), .Z(n_182564160
		));
	notech_nand3 i_17355132(.A(n_62433), .B(opc[10]), .C(n_177464112), .Z(n_182264157
		));
	notech_nand3 i_17855127(.A(n_54128), .B(tsc[42]), .C(n_59826), .Z(n_181764152
		));
	notech_nao3 i_8355222(.A(n_62429), .B(opc[13]), .C(n_336265664), .Z(n_181264149
		));
	notech_nand2 i_8655219(.A(n_337865680), .B(opb[13]), .Z(n_180864146));
	notech_or4 i_8955216(.A(n_60779), .B(n_60726), .C(n_55843), .D(nbus_11326
		[13]), .Z(n_180564143));
	notech_nand3 i_9055215(.A(n_54124), .B(tsc[13]), .C(n_59826), .Z(n_180264140
		));
	notech_nao3 i_7355232(.A(n_62433), .B(opc[12]), .C(n_336265664), .Z(n_180164139
		));
	notech_nand2 i_7655229(.A(n_337865680), .B(opb[12]), .Z(n_179864136));
	notech_or4 i_7955226(.A(n_60779), .B(n_60726), .C(n_55843), .D(nbus_11326
		[12]), .Z(n_179564133));
	notech_and3 i_8055225(.A(n_54124), .B(tsc[12]), .C(n_59826), .Z(n_179264130
		));
	notech_nao3 i_6355242(.A(n_62429), .B(opc[11]), .C(n_336265664), .Z(n_179164129
		));
	notech_nand2 i_6655239(.A(n_337865680), .B(opb[11]), .Z(n_178864126));
	notech_or4 i_6955236(.A(n_60779), .B(n_60729), .C(n_55843), .D(nbus_11326
		[11]), .Z(n_178564123));
	notech_and3 i_7055235(.A(n_54124), .B(tsc[11]), .C(n_59826), .Z(n_178264120
		));
	notech_ao4 i_52560710(.A(n_204988864), .B(n_56104), .C(n_2240), .D(n_26583
		), .Z(n_178164119));
	notech_and2 i_52760709(.A(n_55846), .B(n_142663764), .Z(n_177864116));
	notech_and4 i_119854147(.A(n_55846), .B(n_280965126), .C(n_55967), .D(n_142663764
		), .Z(n_177764115));
	notech_and4 i_195460623(.A(n_54642), .B(n_54762), .C(n_1082), .D(n_2661)
		, .Z(n_177664114));
	notech_nand3 i_192660635(.A(n_2657), .B(n_1083), .C(n_2659), .Z(n_177564113
		));
	notech_nand2 i_195960621(.A(n_54606), .B(n_141963757), .Z(n_177464112)
		);
	notech_and4 i_1355284(.A(n_56061), .B(n_243864755), .C(n_258664903), .D(n_55976
		), .Z(n_177364111));
	notech_nand2 i_5255310(.A(opc_10[15]), .B(n_62401), .Z(n_177264110));
	notech_nand2 i_1055314(.A(n_62433), .B(opc[15]), .Z(n_177164109));
	notech_and4 i_126356668(.A(n_176764105), .B(n_169964037), .C(n_170264040
		), .D(n_26339), .Z(n_177064108));
	notech_ao4 i_126156670(.A(n_27566), .B(n_263036785), .C(n_355188244), .D
		(n_322788463), .Z(n_176764105));
	notech_ao4 i_126556667(.A(n_54607), .B(n_351265801), .C(\nbus_11276[5] )
		, .D(n_54948), .Z(n_176464102));
	notech_and3 i_126856664(.A(n_170764045), .B(n_170664044), .C(n_170864046
		), .Z(n_176364101));
	notech_and4 i_127856658(.A(n_168964027), .B(n_175764095), .C(n_170964047
		), .D(n_171264050), .Z(n_176064098));
	notech_ao4 i_127256660(.A(n_27570), .B(n_351165800), .C(n_355188244), .D
		(n_57351), .Z(n_175764095));
	notech_and4 i_128556653(.A(n_175464092), .B(n_175264090), .C(n_171564053
		), .D(n_171864056), .Z(n_175664094));
	notech_ao4 i_127956657(.A(n_2679), .B(n_54607), .C(n_56035), .D(n_169464032
		), .Z(n_175464092));
	notech_ao4 i_128356655(.A(nbus_11273[7]), .B(n_169264030), .C(n_2680), .D
		(n_169164029), .Z(n_175264090));
	notech_ao4 i_145456495(.A(n_55740), .B(n_27566), .C(n_57321), .D(n_55685
		), .Z(n_175064088));
	notech_ao4 i_145556494(.A(n_55518), .B(n_322788463), .C(n_55380), .D(\nbus_11276[5] 
		), .Z(n_174964087));
	notech_and3 i_146056489(.A(n_174564083), .B(n_174764085), .C(n_172764065
		), .Z(n_174864086));
	notech_ao4 i_145756492(.A(n_249834124), .B(n_29065), .C(n_249534121), .D
		(n_351265801), .Z(n_174764085));
	notech_ao4 i_145856491(.A(n_248934115), .B(nbus_11273[5]), .C(n_202067840
		), .D(n_27524), .Z(n_174564083));
	notech_ao4 i_167956278(.A(n_316788522), .B(n_321188478), .C(n_249134117)
		, .D(n_60473), .Z(n_174464082));
	notech_ao4 i_169756260(.A(n_27524), .B(n_59826), .C(n_55920), .D(n_322788463
		), .Z(n_174364081));
	notech_ao4 i_169856259(.A(n_55810), .B(nbus_11273[5]), .C(n_56045), .D(\nbus_11276[5] 
		), .Z(n_174164079));
	notech_ao4 i_170356255(.A(n_27526), .B(n_59826), .C(n_57351), .D(n_55920
		), .Z(n_174064078));
	notech_ao4 i_170456254(.A(n_55810), .B(nbus_11273[7]), .C(n_247634102), 
		.D(n_59927), .Z(n_173964077));
	notech_or4 i_87857037(.A(n_60779), .B(n_60729), .C(n_1135), .D(n_29065),
		 .Z(n_173464072));
	notech_or4 i_65757237(.A(n_2145), .B(n_1976), .C(n_120857496), .D(n_351365802
		), .Z(n_172764065));
	notech_nand2 i_46057417(.A(opb[7]), .B(n_169364031), .Z(n_171864056));
	notech_nao3 i_46357414(.A(n_26248), .B(\opa_12[7] ), .C(n_351565804), .Z
		(n_171564053));
	notech_or4 i_46657411(.A(n_60779), .B(n_60729), .C(n_55843), .D(nbus_11326
		[7]), .Z(n_171264050));
	notech_nand3 i_46757410(.A(n_54124), .B(tsc[7]), .C(n_59826), .Z(n_170964047
		));
	notech_nand2 i_45057427(.A(opa[5]), .B(n_54949), .Z(n_170864046));
	notech_or4 i_44957428(.A(n_58660), .B(n_56121), .C(n_55837), .D(n_57321)
		, .Z(n_170764045));
	notech_or4 i_44857429(.A(n_351365802), .B(n_55097), .C(n_114626850), .D(n_229364616
		), .Z(n_170664044));
	notech_nao3 i_45357424(.A(n_26248), .B(\opa_12[5] ), .C(n_351565804), .Z
		(n_170564043));
	notech_nand3 i_45657421(.A(n_54124), .B(tsc[5]), .C(n_59826), .Z(n_170264040
		));
	notech_or2 i_45757420(.A(n_61624), .B(nbus_11326[5]), .Z(n_169964037));
	notech_or2 i_84157074(.A(n_316688523), .B(nbus_11273[4]), .Z(n_169564033
		));
	notech_ao4 i_138857935(.A(n_2675), .B(n_55837), .C(n_55580), .D(n_27570)
		, .Z(n_169464032));
	notech_nand3 i_4857809(.A(n_55142), .B(n_222168040), .C(n_350965798), .Z
		(n_169364031));
	notech_and3 i_4757810(.A(n_55143), .B(n_222268041), .C(n_350865797), .Z(n_169264030
		));
	notech_and2 i_4657811(.A(n_50635), .B(n_336065662), .Z(n_169164029));
	notech_and2 i_64257893(.A(n_174064078), .B(n_173964077), .Z(n_168964027)
		);
	notech_nand3 i_43757899(.A(n_173464072), .B(n_174164079), .C(n_174364081
		), .Z(n_168864026));
	notech_and4 i_94159679(.A(n_142963767), .B(n_168364021), .C(n_26404), .D
		(n_143263770), .Z(n_168664024));
	notech_ao4 i_93859681(.A(n_161857906), .B(n_336265664), .C(n_161957907),
		 .D(n_336065662), .Z(n_168364021));
	notech_and4 i_95459674(.A(n_143563773), .B(n_168064018), .C(n_167864016)
		, .D(n_143863776), .Z(n_168264020));
	notech_ao4 i_94459678(.A(n_27571), .B(n_337665678), .C(n_57350), .D(n_350965798
		), .Z(n_168064018));
	notech_ao4 i_94859676(.A(nbus_11273[8]), .B(n_26244), .C(n_350865797), .D
		(n_29045), .Z(n_167864016));
	notech_and4 i_101059619(.A(n_54860), .B(n_167564013), .C(n_167364011), .D
		(n_144363781), .Z(n_167764015));
	notech_ao4 i_100659623(.A(n_55131), .B(n_29190), .C(n_131423301), .D(n_27597
		), .Z(n_167564013));
	notech_ao4 i_100859621(.A(n_110923096), .B(n_302421911), .C(n_270688747)
		, .D(n_302221909), .Z(n_167364011));
	notech_and4 i_101559614(.A(n_167064008), .B(n_166864006), .C(n_144663784
		), .D(n_144963787), .Z(n_167264010));
	notech_ao4 i_101159618(.A(n_57329), .B(n_242764744), .C(n_55534), .D(nbus_11273
		[29]), .Z(n_167064008));
	notech_ao4 i_101359616(.A(n_170914103), .B(n_27552), .C(n_59186), .D(n_26676
		), .Z(n_166864006));
	notech_and4 i_102859601(.A(n_145063788), .B(n_145363791), .C(n_166464002
		), .D(n_26404), .Z(n_166764005));
	notech_ao4 i_102659603(.A(n_2662), .B(n_29045), .C(n_2663), .D(n_57350),
		 .Z(n_166464002));
	notech_ao4 i_102959600(.A(n_161957907), .B(n_324388255), .C(n_327665580)
		, .D(n_27571), .Z(n_166264000));
	notech_ao4 i_103059599(.A(n_327465578), .B(\nbus_11276[8] ), .C(n_161857906
		), .D(n_324288256), .Z(n_166063998));
	notech_and4 i_103659593(.A(n_53844), .B(n_165663994), .C(n_26240), .D(n_146163799
		), .Z(n_165963997));
	notech_ao4 i_103459595(.A(n_55085), .B(n_55867), .C(n_2662), .D(n_29048)
		, .Z(n_165663994));
	notech_ao4 i_103759592(.A(n_57349), .B(n_2663), .C(n_352969301), .D(n_324388255
		), .Z(n_165463992));
	notech_ao4 i_103859591(.A(n_177664114), .B(\nbus_11276[9] ), .C(n_353069302
		), .D(n_26330), .Z(n_165263990));
	notech_and3 i_105059579(.A(n_164963987), .B(n_146763805), .C(n_26339), .Z
		(n_165163989));
	notech_ao4 i_104959580(.A(n_54749), .B(n_29065), .C(n_54923), .D(nbus_11273
		[5]), .Z(n_164963987));
	notech_ao4 i_105559578(.A(n_54922), .B(\nbus_11276[5] ), .C(n_55898), .D
		(n_142163759), .Z(n_164763985));
	notech_ao4 i_105659577(.A(n_259336748), .B(n_351265801), .C(n_150774375)
		, .D(n_164563983), .Z(n_164663984));
	notech_nao3 i_105859575(.A(n_56492), .B(n_268064997), .C(n_351365802), .Z
		(n_164563983));
	notech_and3 i_107759557(.A(n_120457492), .B(n_132957617), .C(n_164263980
		), .Z(n_164363981));
	notech_ao4 i_107659558(.A(n_59186), .B(n_26686), .C(n_56024), .D(n_29191
		), .Z(n_164263980));
	notech_ao4 i_107859556(.A(n_55977), .B(n_28415), .C(n_208364418), .D(n_55331
		), .Z(n_164063978));
	notech_ao4 i_107959555(.A(n_57325), .B(n_280865125), .C(nbus_11273[1]), 
		.D(n_208264417), .Z(n_163963977));
	notech_and4 i_108759547(.A(n_163663974), .B(n_163463972), .C(n_163363971
		), .D(n_148263820), .Z(n_163863976));
	notech_ao4 i_108259552(.A(n_295965276), .B(n_29049), .C(n_57357), .D(n_295765274
		), .Z(n_163663974));
	notech_ao4 i_108459550(.A(n_262636781), .B(n_26925), .C(n_262536780), .D
		(n_27520), .Z(n_163463972));
	notech_ao4 i_108559549(.A(n_353869309), .B(n_206664401), .C(n_353769308)
		, .D(n_206764402), .Z(n_163363971));
	notech_and4 i_117059466(.A(n_191467734), .B(n_163063968), .C(n_177967599
		), .D(n_177867598), .Z(n_163163969));
	notech_ao4 i_116959467(.A(n_59186), .B(n_26688), .C(n_56024), .D(n_29194
		), .Z(n_163063968));
	notech_ao4 i_117159465(.A(n_55977), .B(n_28417), .C(n_208364418), .D(n_27564
		), .Z(n_162863966));
	notech_ao4 i_117259464(.A(n_57323), .B(n_280865125), .C(n_56667), .D(n_208264417
		), .Z(n_162763965));
	notech_and4 i_118259456(.A(n_162463962), .B(n_162263960), .C(n_162163959
		), .D(n_149563833), .Z(n_162663964));
	notech_ao4 i_117659461(.A(n_295965276), .B(n_29043), .C(n_322688464), .D
		(n_295765274), .Z(n_162463962));
	notech_ao4 i_117859459(.A(n_262636781), .B(n_26929), .C(n_262536780), .D
		(n_27522), .Z(n_162263960));
	notech_ao4 i_118059458(.A(n_353369305), .B(n_206664401), .C(n_353269304)
		, .D(n_206764402), .Z(n_162163959));
	notech_and3 i_118459454(.A(n_174464082), .B(n_161863956), .C(n_169564033
		), .Z(n_161963957));
	notech_ao4 i_118359455(.A(n_59186), .B(n_26689), .C(n_56024), .D(n_29195
		), .Z(n_161863956));
	notech_ao4 i_118559453(.A(n_55977), .B(n_28418), .C(n_208364418), .D(n_27565
		), .Z(n_161663954));
	notech_ao4 i_118659452(.A(n_319588494), .B(n_280865125), .C(nbus_11273[4
		]), .D(n_208264417), .Z(n_161563953));
	notech_and4 i_119659444(.A(n_161263950), .B(n_161063948), .C(n_160963947
		), .D(n_150863846), .Z(n_161463952));
	notech_ao4 i_119159449(.A(n_295965276), .B(n_29063), .C(n_321188478), .D
		(n_295765274), .Z(n_161263950));
	notech_ao4 i_119359447(.A(n_262636781), .B(n_26931), .C(n_262536780), .D
		(n_27523), .Z(n_161063948));
	notech_ao4 i_119459446(.A(n_316388526), .B(n_206664401), .C(n_316288527)
		, .D(n_206764402), .Z(n_160963947));
	notech_and3 i_119859442(.A(n_183678231), .B(n_160663944), .C(n_144577845
		), .Z(n_160763945));
	notech_ao4 i_119759443(.A(n_59186), .B(n_26691), .C(n_56024), .D(n_29198
		), .Z(n_160663944));
	notech_ao4 i_119959441(.A(n_55977), .B(n_28420), .C(n_208364418), .D(n_27568
		), .Z(n_160463942));
	notech_ao4 i_120059440(.A(n_57320), .B(n_280865125), .C(nbus_11273[6]), 
		.D(n_208264417), .Z(n_160363941));
	notech_and4 i_120959432(.A(n_160063938), .B(n_159863936), .C(n_159763935
		), .D(n_152163859), .Z(n_160263940));
	notech_ao4 i_120359437(.A(n_295965276), .B(n_29068), .C(n_57352), .D(n_295765274
		), .Z(n_160063938));
	notech_ao4 i_120559435(.A(n_262636781), .B(n_26935), .C(n_262536780), .D
		(n_27525), .Z(n_159863936));
	notech_ao4 i_120659434(.A(n_316488525), .B(n_206664401), .C(n_316588524)
		, .D(n_206764402), .Z(n_159763935));
	notech_and3 i_121159430(.A(n_158074448), .B(n_159463932), .C(n_150874376
		), .Z(n_159563933));
	notech_ao4 i_121059431(.A(n_59186), .B(n_26692), .C(n_56024), .D(n_29199
		), .Z(n_159463932));
	notech_ao4 i_121259429(.A(n_55977), .B(n_28421), .C(n_208364418), .D(n_27570
		), .Z(n_159263930));
	notech_ao4 i_121359428(.A(n_2675), .B(n_280865125), .C(nbus_11273[7]), .D
		(n_208264417), .Z(n_159163929));
	notech_and4 i_122259420(.A(n_158863926), .B(n_158663924), .C(n_158563923
		), .D(n_153463872), .Z(n_159063928));
	notech_ao4 i_121659425(.A(n_28983), .B(n_295965276), .C(n_57351), .D(n_295765274
		), .Z(n_158863926));
	notech_ao4 i_121859423(.A(n_262636781), .B(n_26937), .C(n_262536780), .D
		(n_27526), .Z(n_158663924));
	notech_ao4 i_122059422(.A(n_2680), .B(n_206664401), .C(n_2679), .D(n_206764402
		), .Z(n_158563923));
	notech_and3 i_128959356(.A(n_132757615), .B(n_132657614), .C(n_158263920
		), .Z(n_158363921));
	notech_ao4 i_128859357(.A(n_321688474), .B(n_29201), .C(n_321788473), .D
		(n_29200), .Z(n_158263920));
	notech_ao4 i_129059355(.A(n_318888501), .B(\nbus_11276[5] ), .C(n_319088499
		), .D(nbus_11273[5]), .Z(n_158063918));
	notech_and4 i_129959347(.A(n_157763915), .B(n_157563913), .C(n_157463912
		), .D(n_154663884), .Z(n_157963917));
	notech_ao4 i_129359352(.A(n_55238), .B(n_322788463), .C(n_55688), .D(n_57321
		), .Z(n_157763915));
	notech_ao4 i_129559350(.A(n_59167), .B(n_27524), .C(n_319288497), .D(n_27566
		), .Z(n_157563913));
	notech_ao4 i_129659349(.A(n_320688483), .B(n_351365802), .C(n_59186), .D
		(n_26721), .Z(n_157463912));
	notech_and4 i_144259222(.A(n_157163909), .B(n_155563893), .C(n_156963907
		), .D(n_154863886), .Z(n_157363911));
	notech_ao4 i_143859226(.A(n_59186), .B(n_26744), .C(n_55951), .D(n_27566
		), .Z(n_157163909));
	notech_ao4 i_144059224(.A(n_55422), .B(n_322788463), .C(n_55421), .D(n_29065
		), .Z(n_156963907));
	notech_and4 i_144759217(.A(n_156663904), .B(n_156463902), .C(n_155863896
		), .D(n_156163899), .Z(n_156863906));
	notech_ao4 i_144359221(.A(\nbus_11276[5] ), .B(n_55304), .C(n_262336778)
		, .D(n_29202), .Z(n_156663904));
	notech_ao4 i_144559219(.A(n_261136766), .B(n_351265801), .C(n_260436759)
		, .D(n_351365802), .Z(n_156463902));
	notech_nao3 i_60859983(.A(n_2424), .B(n_29091), .C(n_232761396), .Z(n_156163899
		));
	notech_or2 i_61259980(.A(n_55316), .B(nbus_11273[5]), .Z(n_155863896));
	notech_or4 i_61659977(.A(n_55837), .B(n_55878), .C(n_57321), .D(n_60589)
		, .Z(n_155563893));
	notech_nand3 i_48460095(.A(n_59188), .B(n_59927), .C(read_data[5]), .Z(n_154863886
		));
	notech_or2 i_48760092(.A(n_55222), .B(n_29065), .Z(n_154663884));
	notech_or4 i_49060089(.A(n_317788512), .B(n_320988480), .C(n_28056), .D(n_60511
		), .Z(n_154363881));
	notech_or2 i_39360177(.A(n_208164416), .B(\nbus_11276[7] ), .Z(n_153463872
		));
	notech_or2 i_37860190(.A(n_208164416), .B(\nbus_11276[6] ), .Z(n_152163859
		));
	notech_or2 i_36460203(.A(n_208164416), .B(\nbus_11276[4] ), .Z(n_150863846
		));
	notech_or2 i_34860216(.A(n_208164416), .B(n_55277), .Z(n_149563833));
	notech_or2 i_29460264(.A(n_208164416), .B(n_59753), .Z(n_148263820));
	notech_or2 i_27260286(.A(n_54695), .B(n_322788463), .Z(n_146763805));
	notech_nand2 i_25360305(.A(opa[9]), .B(n_177564113), .Z(n_146663804));
	notech_nand3 i_25860300(.A(n_54124), .B(tsc[41]), .C(n_59826), .Z(n_146163799
		));
	notech_or2 i_24360314(.A(n_327565579), .B(nbus_11273[8]), .Z(n_145863796
		));
	notech_or4 i_24960309(.A(instrc[115]), .B(instrc[112]), .C(n_157974447),
		 .D(n_56086), .Z(n_145363791));
	notech_nand3 i_25060308(.A(n_54124), .B(tsc[40]), .C(n_59826), .Z(n_145063788
		));
	notech_or2 i_22160334(.A(n_55533), .B(\nbus_11276[29] ), .Z(n_144963787)
		);
	notech_or2 i_22560331(.A(n_242664743), .B(n_28977), .Z(n_144663784));
	notech_nao3 i_22860328(.A(n_26549), .B(opc[29]), .C(n_316988520), .Z(n_144363781
		));
	notech_nand2 i_15760398(.A(opb[8]), .B(n_337865680), .Z(n_143863776));
	notech_or4 i_16060395(.A(instrc[115]), .B(instrc[112]), .C(n_157974447),
		 .D(n_58661), .Z(n_143563773));
	notech_or4 i_16360392(.A(n_60775), .B(n_60729), .C(n_55843), .D(nbus_11326
		[8]), .Z(n_143263770));
	notech_nand3 i_16460391(.A(n_54124), .B(tsc[8]), .C(n_59837), .Z(n_142963767
		));
	notech_or4 i_87259744(.A(n_260688757), .B(n_2605), .C(n_205088863), .D(n_26583
		), .Z(n_142663764));
	notech_or4 i_86859748(.A(instrc[115]), .B(instrc[112]), .C(n_56086), .D(n_36952
		), .Z(n_142563763));
	notech_and2 i_83959771(.A(n_55967), .B(n_142063758), .Z(n_142363761));
	notech_and2 i_82759783(.A(n_318365500), .B(n_56029), .Z(n_142263760));
	notech_ao4 i_151760612(.A(n_55837), .B(n_57321), .C(n_54089), .D(n_27566
		), .Z(n_142163759));
	notech_and3 i_76060586(.A(n_55846), .B(n_142663764), .C(n_178164119), .Z
		(n_142063758));
	notech_or2 i_9082(.A(n_2689), .B(n_54668), .Z(n_141963757));
	notech_and4 i_106462520(.A(n_53844), .B(n_121463552), .C(n_141563753), .D
		(n_201667836), .Z(n_141863756));
	notech_ao4 i_106262522(.A(n_107626780), .B(n_28716), .C(n_2687), .D(n_27564
		), .Z(n_141563753));
	notech_and4 i_106962515(.A(n_141263750), .B(n_141063748), .C(n_121763555
		), .D(n_122063558), .Z(n_141463752));
	notech_ao4 i_106562519(.A(n_2661), .B(n_322688464), .C(n_2659), .D(n_29043
		), .Z(n_141263750));
	notech_ao4 i_106762517(.A(n_120763545), .B(n_55277), .C(n_120663544), .D
		(n_140963747), .Z(n_141063748));
	notech_nao3 i_107062514(.A(n_62429), .B(opc[3]), .C(n_2689), .Z(n_140963747
		));
	notech_and4 i_108262502(.A(n_53844), .B(n_122363561), .C(n_140563743), .D
		(n_26339), .Z(n_140863746));
	notech_ao4 i_108062504(.A(n_107626780), .B(n_28717), .C(n_27566), .D(n_2687
		), .Z(n_140563743));
	notech_and4 i_108762497(.A(n_140263740), .B(n_140063738), .C(n_122663564
		), .D(n_122963567), .Z(n_140463742));
	notech_ao4 i_108362501(.A(n_2661), .B(n_322788463), .C(n_29065), .D(n_2659
		), .Z(n_140263740));
	notech_ao4 i_108562499(.A(\nbus_11276[5] ), .B(n_120763545), .C(n_120663544
		), .D(n_139963737), .Z(n_140063738));
	notech_nao3 i_108862496(.A(n_62433), .B(opc[5]), .C(n_2689), .Z(n_139963737
		));
	notech_and4 i_109262492(.A(n_139563733), .B(n_168964027), .C(n_123063568
		), .D(n_123363571), .Z(n_139863736));
	notech_ao4 i_109062494(.A(n_2679), .B(n_54606), .C(n_57351), .D(n_2661),
		 .Z(n_139563733));
	notech_ao4 i_109362491(.A(n_2659), .B(n_28983), .C(n_322865545), .D(n_27570
		), .Z(n_139363731));
	notech_ao4 i_109462490(.A(nbus_11273[7]), .B(n_121063548), .C(n_2680), .D
		(n_120963547), .Z(n_139163729));
	notech_and3 i_109962485(.A(n_120557493), .B(n_132857616), .C(n_138763725
		), .Z(n_138863726));
	notech_ao4 i_109862486(.A(n_57324), .B(n_280865125), .C(n_262536780), .D
		(n_27521), .Z(n_138763725));
	notech_ao4 i_110062484(.A(n_55977), .B(n_28416), .C(n_56024), .D(n_29188
		), .Z(n_138563723));
	notech_ao4 i_110162483(.A(n_295965276), .B(n_29050), .C(n_322488466), .D
		(n_295765274), .Z(n_138463722));
	notech_and4 i_110962475(.A(n_124863586), .B(n_138163719), .C(n_137963717
		), .D(n_137863716), .Z(n_138363721));
	notech_ao4 i_110462480(.A(n_353469306), .B(n_206764402), .C(n_208164416)
		, .D(n_55289), .Z(n_138163719));
	notech_ao4 i_110662478(.A(n_56658), .B(n_208264417), .C(n_208364418), .D
		(n_55299), .Z(n_137963717));
	notech_ao4 i_110762477(.A(n_26927), .B(n_262636781), .C(n_59188), .D(n_26687
		), .Z(n_137863716));
	notech_and3 i_111162473(.A(n_132757615), .B(n_132657614), .C(n_137563713
		), .Z(n_137663714));
	notech_ao4 i_111062474(.A(n_57321), .B(n_280865125), .C(n_27566), .D(n_208364418
		), .Z(n_137563713));
	notech_ao4 i_111262472(.A(n_262536780), .B(n_27524), .C(n_55977), .D(n_28419
		), .Z(n_137363711));
	notech_ao4 i_111362471(.A(n_56024), .B(n_29189), .C(n_295965276), .D(n_29065
		), .Z(n_137263710));
	notech_and4 i_112162463(.A(n_126163599), .B(n_136963707), .C(n_136763705
		), .D(n_136663704), .Z(n_137163709));
	notech_ao4 i_111662468(.A(\nbus_11276[5] ), .B(n_208164416), .C(nbus_11273
		[5]), .D(n_208264417), .Z(n_136963707));
	notech_ao4 i_111862466(.A(n_351265801), .B(n_206764402), .C(n_351365802)
		, .D(n_206664401), .Z(n_136763705));
	notech_ao4 i_111962465(.A(n_262636781), .B(n_26933), .C(n_59188), .D(n_26690
		), .Z(n_136663704));
	notech_and3 i_117762410(.A(n_136363701), .B(n_126663604), .C(n_26339), .Z
		(n_136563703));
	notech_ao4 i_117662411(.A(n_54740), .B(n_322788463), .C(n_54920), .D(\nbus_11276[5] 
		), .Z(n_136363701));
	notech_ao4 i_117862409(.A(n_54921), .B(nbus_11273[5]), .C(n_248434110), 
		.D(n_351265801), .Z(n_136163699));
	notech_ao4 i_117962408(.A(n_55864), .B(n_142163759), .C(n_273539523), .D
		(n_135963697), .Z(n_136063698));
	notech_nand3 i_118162406(.A(n_62429), .B(n_26381), .C(opc[5]), .Z(n_135963697
		));
	notech_and3 i_123362355(.A(n_135663694), .B(n_127363611), .C(n_26339), .Z
		(n_135863696));
	notech_ao4 i_123262356(.A(n_54432), .B(n_322788463), .C(n_254634172), .D
		(n_351265801), .Z(n_135663694));
	notech_ao4 i_123462354(.A(n_54451), .B(n_142163759), .C(n_269439482), .D
		(\nbus_11276[5] ), .Z(n_135463692));
	notech_ao4 i_123562353(.A(n_269339481), .B(nbus_11273[5]), .C(n_351365802
		), .D(n_254734173), .Z(n_135363691));
	notech_ao4 i_127162318(.A(n_54435), .B(n_29065), .C(n_54458), .D(n_322788463
		), .Z(n_134963687));
	notech_nand3 i_127662313(.A(n_128763625), .B(n_134563683), .C(n_134763685
		), .Z(n_134863686));
	notech_ao4 i_127362316(.A(n_54563), .B(\nbus_11276[5] ), .C(n_54565), .D
		(nbus_11273[5]), .Z(n_134763685));
	notech_ao4 i_127462315(.A(n_54439), .B(n_142163759), .C(n_351365802), .D
		(n_247334099), .Z(n_134563683));
	notech_and3 i_131062281(.A(n_134163679), .B(n_128863626), .C(n_26339), .Z
		(n_134363681));
	notech_ao4 i_130762282(.A(n_356076396), .B(n_322788463), .C(n_351265801)
		, .D(n_356376399), .Z(n_134163679));
	notech_ao4 i_131162280(.A(n_56068), .B(n_142163759), .C(n_269539483), .D
		(nbus_11273[5]), .Z(n_133963677));
	notech_ao4 i_131262279(.A(n_268739475), .B(n_55375), .C(n_351365802), .D
		(n_356276398), .Z(n_133863676));
	notech_ao4 i_135162240(.A(n_322788463), .B(n_54456), .C(n_351265801), .D
		(n_247534101), .Z(n_133463672));
	notech_nand3 i_135562236(.A(n_130063638), .B(n_133263670), .C(n_130163639
		), .Z(n_133363671));
	notech_ao4 i_135362238(.A(n_56009), .B(n_142163759), .C(n_55375), .D(n_269739485
		), .Z(n_133263670));
	notech_ao4 i_139462198(.A(n_54428), .B(n_322788463), .C(n_351265801), .D
		(n_2685), .Z(n_132763665));
	notech_nand3 i_139862194(.A(n_130763645), .B(n_132563663), .C(n_130863646
		), .Z(n_132663664));
	notech_ao4 i_139662196(.A(n_56151), .B(n_142163759), .C(n_55375), .D(n_269939487
		), .Z(n_132563663));
	notech_and3 i_144362149(.A(n_132063658), .B(n_130963647), .C(n_26339), .Z
		(n_132263660));
	notech_ao4 i_144262150(.A(n_54656), .B(nbus_11273[5]), .C(n_54655), .D(n_55375
		), .Z(n_132063658));
	notech_ao4 i_144462148(.A(n_322788463), .B(n_54469), .C(n_29065), .D(n_54438
		), .Z(n_131863656));
	notech_ao4 i_144562147(.A(n_279739585), .B(n_351365802), .C(n_275539543)
		, .D(n_351265801), .Z(n_131763655));
	notech_or2 i_65962911(.A(n_55872), .B(n_142163759), .Z(n_130963647));
	notech_or2 i_59862970(.A(n_269839486), .B(nbus_11273[5]), .Z(n_130863646
		));
	notech_or4 i_59762971(.A(n_264436799), .B(n_2664), .C(n_351365802), .D(n_2349
		), .Z(n_130763645));
	notech_nor2 i_60362965(.A(n_54468), .B(n_29065), .Z(n_130263640));
	notech_or2 i_54963016(.A(n_269639484), .B(nbus_11273[5]), .Z(n_130163639
		));
	notech_or4 i_54863017(.A(n_1976), .B(n_54071), .C(n_351365802), .D(n_355988238
		), .Z(n_130063638));
	notech_nor2 i_55463011(.A(n_54450), .B(n_29065), .Z(n_129563633));
	notech_or2 i_50863057(.A(n_356176397), .B(n_29065), .Z(n_128863626));
	notech_nao3 i_46563100(.A(opc_10[5]), .B(n_62401), .C(n_247234098), .Z(n_128763625
		));
	notech_ao3 i_47063095(.A(n_26826), .B(opc[5]), .C(n_2645), .Z(n_128063618
		));
	notech_or2 i_42763138(.A(n_54436), .B(n_29065), .Z(n_127363611));
	notech_or2 i_36763198(.A(n_54748), .B(n_29065), .Z(n_126663604));
	notech_or2 i_29363268(.A(n_322788463), .B(n_295765274), .Z(n_126163599)
		);
	notech_nao3 i_28063281(.A(n_62433), .B(opc[2]), .C(n_206664401), .Z(n_124863586
		));
	notech_or4 i_27363288(.A(n_2740), .B(n_1076), .C(n_60532), .D(n_56027), 
		.Z(n_123963577));
	notech_or2 i_26563295(.A(n_121163549), .B(\nbus_11276[7] ), .Z(n_123863576
		));
	notech_nand3 i_27163290(.A(n_54124), .B(tsc[39]), .C(n_59835), .Z(n_123363571
		));
	notech_or4 i_27263289(.A(instrc[115]), .B(instrc[112]), .C(n_56086), .D(n_169464032
		), .Z(n_123063568));
	notech_nand2 i_25663304(.A(n_120863546), .B(opa[5]), .Z(n_122963567));
	notech_nao3 i_25963301(.A(opc_10[5]), .B(n_62403), .C(n_54606), .Z(n_122663564
		));
	notech_or4 i_26263298(.A(n_56081), .B(n_56121), .C(n_55837), .D(n_57321)
		, .Z(n_122363561));
	notech_nand2 i_23863322(.A(n_120863546), .B(opa[3]), .Z(n_122063558));
	notech_nao3 i_24163319(.A(opc_10[3]), .B(n_62413), .C(n_54606), .Z(n_121763555
		));
	notech_or4 i_24463316(.A(n_55837), .B(n_57323), .C(n_56074), .D(n_56121)
		, .Z(n_121463552));
	notech_and4 i_19063361(.A(n_339065692), .B(n_328165585), .C(n_123963577)
		, .D(n_2663), .Z(n_121163549));
	notech_and3 i_18963362(.A(n_2657), .B(n_1083), .C(n_2662), .Z(n_121063548
		));
	notech_and2 i_18863363(.A(n_324388255), .B(n_141963757), .Z(n_120963547)
		);
	notech_nand2 i_10663442(.A(n_241864737), .B(n_2657), .Z(n_120863546));
	notech_and4 i_10763441(.A(n_54642), .B(n_54762), .C(n_328165585), .D(n_241764736
		), .Z(n_120763545));
	notech_and2 i_6563482(.A(n_56029), .B(n_120563543), .Z(n_120663544));
	notech_and4 i_3263515(.A(n_56060), .B(n_1081), .C(n_56061), .D(n_1079), 
		.Z(n_120563543));
	notech_and3 i_71432889(.A(n_346988339), .B(n_346888340), .C(n_347388335)
		, .Z(n_2223));
	notech_nand2 i_25641(.A(all_cnt[0]), .B(n_27556), .Z(n_2351));
	notech_nand3 i_176833045(.A(all_cnt[0]), .B(all_cnt[1]), .C(n_27557), .Z
		(n_54703));
	notech_nand3 i_129033046(.A(all_cnt[0]), .B(all_cnt[1]), .C(all_cnt[2]),
		 .Z(n_55089));
	notech_and2 i_104633047(.A(all_cnt[0]), .B(all_cnt[1]), .Z(n_55323));
	notech_nao3 i_18917(.A(n_26390), .B(n_26296), .C(n_206288851), .Z(n_38340
		));
	notech_or4 i_172133154(.A(n_28975), .B(n_244656264), .C(n_60511), .D(n_2586
		), .Z(n_54741));
	notech_or2 i_8218(.A(n_335262250), .B(n_29123), .Z(n_49023));
	notech_nand2 i_55070(.A(n_49023), .B(n_57470), .Z(\nbus_11355[0] ));
	notech_nand2 i_55071(.A(n_61176), .B(n_335562253), .Z(n_57470));
	notech_and4 i_54342(.A(n_341088366), .B(n_345388355), .C(n_346088348), .D
		(n_345088358), .Z(\nbus_11352[0] ));
	notech_or4 i_535677(.A(n_26380), .B(n_26629), .C(n_333188381), .D(n_331888394
		), .Z(n_328046808));
	notech_or4 i_235679(.A(n_2773), .B(n_2825), .C(n_260688757), .D(n_2605),
		 .Z(n_328246806));
	notech_nand2 i_114635763(.A(n_190488901), .B(n_57431), .Z(n_55226));
	notech_or4 i_124139103(.A(n_2145), .B(n_316888521), .C(n_319888491), .D(n_60507
		), .Z(n_55133));
	notech_nand2 i_1921182(.A(n_322562229), .B(n_322062224), .Z(n_13575));
	notech_nand2 i_2021183(.A(n_321562219), .B(n_321062214), .Z(n_13581));
	notech_nand2 i_2121184(.A(n_320562209), .B(n_320062204), .Z(n_13587));
	notech_nand2 i_2221185(.A(n_319562199), .B(n_319062194), .Z(n_13593));
	notech_nand2 i_2321186(.A(n_318562189), .B(n_318062184), .Z(n_13599));
	notech_nand2 i_2120640(.A(n_317562179), .B(n_317062174), .Z(n_20231));
	notech_nand2 i_2220641(.A(n_315062154), .B(n_314562149), .Z(n_20237));
	notech_and4 i_144442260(.A(n_313862142), .B(n_313762141), .C(n_313362137
		), .D(n_313662140), .Z(n_310518882));
	notech_and4 i_144342261(.A(n_316362167), .B(n_316262166), .C(n_315862162
		), .D(n_316162165), .Z(n_310618883));
	notech_and4 i_93229156(.A(n_312062124), .B(n_311962123), .C(n_311562119)
		, .D(n_311862122), .Z(n_311018887));
	notech_and4 i_93129155(.A(n_310662110), .B(n_310562109), .C(n_310162105)
		, .D(n_310462108), .Z(n_311118888));
	notech_mux2 i_2211679(.S(n_60136), .A(regs_14[21]), .B(add_len_pc32[21])
		, .Z(\add_len_pc[21] ));
	notech_mux2 i_2111678(.S(n_60136), .A(regs_14[20]), .B(add_len_pc32[20])
		, .Z(\add_len_pc[20] ));
	notech_ao4 i_37442270(.A(n_56573), .B(n_56502), .C(n_55837), .D(n_26513)
		, .Z(n_55975));
	notech_or4 i_156342278(.A(n_273888717), .B(n_294061944), .C(n_59235), .D
		(n_55969), .Z(n_54872));
	notech_or2 i_152842279(.A(n_55969), .B(n_293061934), .Z(n_54902));
	notech_nand2 i_2421187(.A(n_292961933), .B(n_292461928), .Z(n_13605));
	notech_nand2 i_2821191(.A(n_291961923), .B(n_291461918), .Z(n_13629));
	notech_nand2 i_2720646(.A(n_290961913), .B(n_290461908), .Z(n_20267));
	notech_nand2 i_2820647(.A(n_288461888), .B(n_287961883), .Z(n_20273));
	notech_and4 i_145045386(.A(n_2872), .B(n_2871), .C(n_2867), .D(n_2870), 
		.Z(n_308221969));
	notech_and4 i_144945387(.A(n_289761901), .B(n_289661900), .C(n_289261896
		), .D(n_289561899), .Z(n_308321970));
	notech_and4 i_93829162(.A(n_2857), .B(n_2856), .C(n_285261875), .D(n_2855
		), .Z(n_308621973));
	notech_and4 i_93729161(.A(n_284361868), .B(n_284261867), .C(n_283861866)
		, .D(n_2841), .Z(n_308721974));
	notech_mux2 i_2811685(.S(n_60136), .A(regs_14[27]), .B(add_len_pc32[27])
		, .Z(\add_len_pc[27] ));
	notech_mux2 i_2711684(.S(n_60138), .A(regs_14[26]), .B(add_len_pc32[26])
		, .Z(\add_len_pc[26] ));
	notech_or4 i_86745433(.A(n_1916), .B(n_148560567), .C(n_59235), .D(n_279961827
		), .Z(n_55487));
	notech_or2 i_86645435(.A(n_279961827), .B(n_54523), .Z(n_55488));
	notech_ao4 i_81542289(.A(n_55967), .B(n_54935), .C(n_55325), .D(n_60473)
		, .Z(n_55536));
	notech_and3 i_81642288(.A(n_54751), .B(n_55692), .C(n_56022), .Z(n_55535
		));
	notech_or4 i_123742240(.A(n_319888491), .B(n_264436799), .C(n_55967), .D
		(n_60507), .Z(n_308518862));
	notech_or2 i_58760592(.A(n_232761396), .B(n_29091), .Z(n_262336778));
	notech_or2 i_59060591(.A(n_232761396), .B(\eflags[10] ), .Z(n_262236777)
		);
	notech_or2 i_131949165(.A(n_323062234), .B(n_261361641), .Z(n_354988259)
		);
	notech_or4 i_124849167(.A(n_56465), .B(n_56469), .C(n_264436799), .D(n_261161639
		), .Z(n_110323090));
	notech_or4 i_39549187(.A(instrc[115]), .B(instrc[112]), .C(n_56163), .D(n_55088
		), .Z(n_110123088));
	notech_and4 i_106549226(.A(n_224461315), .B(n_55978), .C(n_225661327), .D
		(n_54710), .Z(n_354888260));
	notech_and3 i_106449227(.A(n_54774), .B(n_55584), .C(n_55979), .Z(n_354788261
		));
	notech_ao4 i_102749229(.A(n_54935), .B(n_261161639), .C(n_60473), .D(n_54761
		), .Z(n_354688262));
	notech_ao4 i_102649230(.A(n_261161639), .B(n_260961637), .C(n_26326), .D
		(n_54874), .Z(n_354588263));
	notech_ao4 i_93649238(.A(n_56040), .B(n_259561623), .C(n_54688), .D(n_60473
		), .Z(n_354488264));
	notech_and2 i_39749262(.A(n_5577), .B(n_45486), .Z(n_354388265));
	notech_and2 i_96645434(.A(n_55488), .B(n_54433), .Z(n_55397));
	notech_and2 i_96745432(.A(n_55487), .B(n_54445), .Z(n_55396));
	notech_or2 i_132345370(.A(n_151860600), .B(n_271761745), .Z(n_306621953)
		);
	notech_or2 i_27171(.A(n_54367), .B(n_55872), .Z(n_309921986));
	notech_or4 i_3645341(.A(n_1976), .B(n_264436799), .C(n_55999), .D(n_60507
		), .Z(n_303521922));
	notech_or4 i_66449257(.A(n_206288851), .B(n_205088863), .C(n_273588720),
		 .D(n_56551), .Z(n_354288266));
	notech_or2 i_29278(.A(n_323062234), .B(n_323262236), .Z(n_354188267));
	notech_or2 i_117739104(.A(n_323062234), .B(n_322962233), .Z(n_354088268)
		);
	notech_and4 i_93529159(.A(n_348988319), .B(n_348888320), .C(n_348488324)
		, .D(n_348788321), .Z(n_57334));
	notech_nand2 i_2555273(.A(read_data[24]), .B(n_59927), .Z(n_316831555)
		);
	notech_ao4 i_38042269(.A(n_56502), .B(n_56551), .C(n_55858), .D(n_26513)
		, .Z(n_55969));
	notech_or2 i_1255285(.A(n_55969), .B(n_294261946), .Z(n_318031567));
	notech_or2 i_855287(.A(n_55094), .B(n_294261946), .Z(n_318231569));
	notech_ao4 i_555289(.A(n_1970), .B(n_29077), .C(n_54698), .D(nbus_11273[
		10]), .Z(n_318431571));
	notech_and4 i_2521860(.A(n_238161449), .B(n_257261600), .C(n_257461602),
		 .D(n_257961607), .Z(n_12545));
	notech_and4 i_1121174(.A(n_256461592), .B(n_257161599), .C(n_239061458),
		 .D(n_256361591), .Z(n_13527));
	notech_nand2 i_1221175(.A(n_255861586), .B(n_255361581), .Z(n_13533));
	notech_nand2 i_1421177(.A(n_254861576), .B(n_254361571), .Z(n_13545));
	notech_nand2 i_2521188(.A(n_253861566), .B(n_253361561), .Z(n_13611));
	notech_and4 i_144755322(.A(n_252261550), .B(n_252161549), .C(n_251761545
		), .D(n_252061548), .Z(n_322231609));
	notech_or2 i_171342277(.A(n_55975), .B(n_293061934), .Z(n_54748));
	notech_nor2 i_10401(.A(n_293161935), .B(n_293061934), .Z(n_46842));
	notech_or4 i_172242276(.A(n_294061944), .B(n_55975), .C(n_59235), .D(n_273888717
		), .Z(n_54740));
	notech_or4 i_10399(.A(n_273888717), .B(n_294061944), .C(n_293161935), .D
		(n_59235), .Z(n_46844));
	notech_ao4 i_37642280(.A(n_56502), .B(n_54520), .C(n_56376), .D(n_26513)
		, .Z(n_55973));
	notech_or4 i_24962(.A(n_250861536), .B(n_250561533), .C(n_250161529), .D
		(n_249861526), .Z(n_321731604));
	notech_and3 i_128555331(.A(n_55975), .B(n_293161935), .C(n_55973), .Z(n_55094
		));
	notech_or2 i_154655337(.A(n_26616), .B(n_321731604), .Z(n_54886));
	notech_or4 i_115442271(.A(n_273888717), .B(n_294061944), .C(n_55973), .D
		(n_59235), .Z(n_55218));
	notech_and3 i_147755338(.A(n_54740), .B(n_46844), .C(n_55218), .Z(n_54943
		));
	notech_or2 i_115342273(.A(n_55973), .B(n_293061934), .Z(n_55219));
	notech_ao3 i_147655339(.A(n_54748), .B(n_55219), .C(n_46842), .Z(n_54944
		));
	notech_and2 i_30289(.A(n_55238), .B(n_318988500), .Z(n_323731624));
	notech_or2 i_57642268(.A(n_56376), .B(n_55864), .Z(n_55773));
	notech_and2 i_62455356(.A(n_55773), .B(n_237361441), .Z(n_55726));
	notech_or4 i_45260712(.A(n_56376), .B(n_206288851), .C(n_60591), .D(n_273588720
		), .Z(n_5538));
	notech_and3 i_77260583(.A(n_54851), .B(n_239561463), .C(n_225961330), .Z
		(n_261436769));
	notech_or4 i_46160594(.A(n_60591), .B(n_59835), .C(n_26604), .D(n_26377)
		, .Z(n_262536780));
	notech_nao3 i_46060595(.A(n_57458), .B(n_26377), .C(n_258636741), .Z(n_262636781
		));
	notech_and4 i_721170(.A(n_227661345), .B(n_236161429), .C(n_236461432), 
		.D(n_236061428), .Z(n_13503));
	notech_and4 i_821171(.A(n_228761356), .B(n_234961418), .C(n_235361421), 
		.D(n_234861417), .Z(n_13509));
	notech_and4 i_1021173(.A(n_233361402), .B(n_234061409), .C(n_230261371),
		 .D(n_233261401), .Z(n_13521));
	notech_and4 i_79882149(.A(n_351388295), .B(n_351088298), .C(n_351588293)
		, .D(n_351488294), .Z(n_57458));
	notech_nand3 i_171960555(.A(n_59188), .B(n_59927), .C(n_275788700), .Z(n_258636741
		));
	notech_nao3 i_11757(.A(n_26390), .B(n_55279), .C(n_59281), .Z(n_45486)
		);
	notech_nand3 i_11716(.A(n_59188), .B(n_59926), .C(read_data[29]), .Z(n_45527
		));
	notech_or2 i_176060646(.A(n_266361691), .B(n_56038), .Z(n_54710));
	notech_or2 i_170960647(.A(n_260961637), .B(n_55967), .Z(n_54751));
	notech_or2 i_169960648(.A(n_55967), .B(n_54935), .Z(n_54759));
	notech_or2 i_168160649(.A(n_56038), .B(n_259561623), .Z(n_54774));
	notech_or2 i_167360650(.A(n_56040), .B(n_259561623), .Z(n_54781));
	notech_or4 i_45160713(.A(n_59281), .B(n_55837), .C(n_273588720), .D(n_60591
		), .Z(n_5577));
	notech_ao4 i_80249243(.A(n_56040), .B(n_266361691), .C(n_55325), .D(n_60473
		), .Z(n_353988269));
	notech_or2 i_153860660(.A(n_56040), .B(n_266361691), .Z(n_54893));
	notech_or4 i_123960664(.A(n_56376), .B(n_56163), .C(n_56121), .D(n_60589
		), .Z(n_55135));
	notech_or2 i_76660690(.A(n_259561623), .B(n_261436769), .Z(n_55584));
	notech_ao4 i_38260715(.A(n_56059), .B(n_60589), .C(n_2250), .D(n_26583),
		 .Z(n_55967));
	notech_ao4 i_37260716(.A(n_275788700), .B(n_59167), .C(n_57420), .D(n_60473
		), .Z(n_55977));
	notech_ao4 i_32560720(.A(n_57419), .B(n_60473), .C(n_54890), .D(n_258636741
		), .Z(n_56024));
	notech_and2 i_31160721(.A(n_54900), .B(n_226961338), .Z(n_56038));
	notech_ao4 i_30960723(.A(n_56059), .B(n_60589), .C(n_2250), .D(n_26226),
		 .Z(n_56040));
	notech_nand2 i_101133063(.A(reps[2]), .B(n_344688362), .Z(n_57456));
	notech_and2 i_148960656(.A(n_231761386), .B(n_56260), .Z(n_54935));
	notech_or4 i_65860696(.A(n_2831), .B(n_2825), .C(n_275288705), .D(n_60473
		), .Z(n_55692));
	notech_or4 i_8239011(.A(n_56465), .B(n_56469), .C(n_2145), .D(n_323362237
		), .Z(n_353788271));
	notech_nao3 i_156682145(.A(n_349988309), .B(n_349488314), .C(n_275788700
		), .Z(n_353688272));
	notech_or4 i_132449209(.A(n_2145), .B(n_56040), .C(n_231461383), .D(n_60511
		), .Z(n_353488274));
	notech_or2 i_154260609(.A(n_57458), .B(n_57441), .Z(n_54890));
	notech_nand2 i_1821181(.A(n_224361314), .B(n_223861309), .Z(n_13569));
	notech_and2 i_138263575(.A(n_54880), .B(n_26551), .Z(n_55006));
	notech_ao4 i_35663562(.A(n_2044), .B(n_56112), .C(n_56063), .D(n_26312),
		 .Z(n_281539603));
	notech_or2 i_10999(.A(n_57378), .B(n_144960531), .Z(n_46244));
	notech_or4 i_15161(.A(n_60779), .B(n_60729), .C(n_55248), .D(n_60589), .Z
		(n_42082));
	notech_and2 i_112463577(.A(n_57420), .B(n_57419), .Z(n_55248));
	notech_nao3 i_11000(.A(n_163860720), .B(n_26487), .C(n_2007), .Z(n_46243
		));
	notech_and2 i_112563578(.A(n_26887), .B(n_145360535), .Z(n_55247));
	notech_or2 i_209663584(.A(n_54523), .B(n_55987), .Z(n_54433));
	notech_or4 i_208163586(.A(n_1916), .B(n_148560567), .C(n_55987), .D(n_59235
		), .Z(n_54445));
	notech_or4 i_153563592(.A(n_59168), .B(n_275388704), .C(n_273688719), .D
		(n_57456), .Z(n_54896));
	notech_and2 i_198563588(.A(n_181860893), .B(n_56260), .Z(n_54523));
	notech_or2 i_130963593(.A(n_54523), .B(n_55999), .Z(n_55070));
	notech_or4 i_130863594(.A(n_1916), .B(n_148560567), .C(n_55999), .D(n_59235
		), .Z(n_55071));
	notech_or2 i_63163599(.A(n_56376), .B(n_55872), .Z(n_55719));
	notech_ao4 i_36263602(.A(n_2044), .B(n_56551), .C(n_55859), .D(n_26312),
		 .Z(n_55987));
	notech_ao4 i_35063603(.A(n_2044), .B(n_54520), .C(n_56376), .D(n_26312),
		 .Z(n_55999));
	notech_ao4 i_34463604(.A(n_56573), .B(n_2044), .C(n_55837), .D(n_26312),
		 .Z(n_56005));
	notech_or4 i_830538(.A(instrc[125]), .B(n_28970), .C(instrc[124]), .D(instrc
		[127]), .Z(n_57292));
	notech_nand2 i_217932(.A(n_222461295), .B(n_222261294), .Z(write_data_27
		[1]));
	notech_and4 i_51634(.A(n_221361285), .B(n_221161284), .C(n_221661288), .D
		(n_221061283), .Z(\nbus_11330[0] ));
	notech_nand2 i_9063457(.A(n_60589), .B(fecx), .Z(n_270739495));
	notech_nao3 i_48861(.A(n_219961272), .B(n_270739495), .C(n_26598), .Z(\nbus_11305[0] 
		));
	notech_and4 i_49125(.A(n_216661239), .B(n_216561238), .C(n_217161244), .D
		(n_216461237), .Z(\nbus_11306[0] ));
	notech_and4 i_49382(.A(n_214161215), .B(n_214061214), .C(n_213961213), .D
		(n_215361227), .Z(\nbus_11307[0] ));
	notech_and4 i_49652(.A(n_212661200), .B(n_212561199), .C(n_208461158), .D
		(n_26474), .Z(\nbus_11308[0] ));
	notech_or2 i_51238(.A(n_353288276), .B(n_142560507), .Z(\nbus_11323[0] )
		);
	notech_or4 i_49905(.A(n_161160693), .B(n_206361137), .C(n_205861132), .D
		(n_26480), .Z(\nbus_11309[0] ));
	notech_or4 i_51987(.A(n_162460706), .B(n_204461118), .C(n_26484), .D(n_26483
		), .Z(\nbus_11331[0] ));
	notech_nao3 i_54736(.A(n_163460716), .B(n_55745), .C(n_163360715), .Z(\nbus_11353[1] 
		));
	notech_or4 i_50162(.A(n_165660738), .B(n_199361067), .C(n_26490), .D(n_26488
		), .Z(\nbus_11310[0] ));
	notech_and4 i_50415(.A(n_196461038), .B(n_196161035), .C(n_197661050), .D
		(n_197061044), .Z(\nbus_11311[0] ));
	notech_nand3 i_52241(.A(n_194761021), .B(n_195861032), .C(n_195161025), 
		.Z(\nbus_11332[0] ));
	notech_and4 i_47154(.A(n_169960781), .B(n_169860780), .C(n_192360997), .D
		(n_193961013), .Z(\nbus_11282[0] ));
	notech_and4 i_53605(.A(n_190560979), .B(n_189560969), .C(n_191360987), .D
		(n_172460806), .Z(\nbus_11349[0] ));
	notech_nand3 i_53858(.A(n_188360957), .B(n_187660950), .C(n_186960943), 
		.Z(\nbus_11350[0] ));
	notech_nao3 i_54111(.A(n_183760911), .B(n_186260936), .C(n_181160889), .Z
		(\nbus_11351[0] ));
	notech_or4 i_168035710(.A(n_59369), .B(n_2550), .C(n_274488713), .D(n_60473
		), .Z(n_54775));
	notech_and4 i_50597(.A(n_334588367), .B(n_334488368), .C(n_54775), .D(n_134360425
		), .Z(\nbus_11314[0] ));
	notech_or4 i_155363591(.A(n_274988708), .B(n_59369), .C(n_200761081), .D
		(n_2260), .Z(n_54880));
	notech_ao4 i_148365671(.A(n_134060422), .B(n_59168), .C(n_200861082), .D
		(n_60473), .Z(n_206841699));
	notech_and4 i_10046(.A(n_59188), .B(n_59837), .C(n_61176), .D(n_133260414
		), .Z(n_353288276));
	notech_or4 i_142068310(.A(n_60779), .B(n_60729), .C(n_60598), .D(n_55546
		), .Z(n_54968));
	notech_ao4 i_8563462(.A(n_221861290), .B(instrc[124]), .C(n_179160873), 
		.D(n_179960880), .Z(n_21051));
	notech_ao4 i_11263580(.A(n_341762311), .B(n_29122), .C(n_137760459), .D(n_26385
		), .Z(n_56153));
	notech_ao4 i_11563581(.A(n_341662310), .B(n_29022), .C(n_137160453), .D(n_26386
		), .Z(n_56150));
	notech_ao4 i_11863582(.A(n_29026), .B(n_26514), .C(n_136860450), .D(n_26387
		), .Z(n_56147));
	notech_ao4 i_10563583(.A(n_341862312), .B(n_29023), .C(n_136460446), .D(n_26388
		), .Z(n_56160));
	notech_nand2 i_2918599(.A(n_132660408), .B(n_132560407), .Z(write_data_32
		[28]));
	notech_nand2 i_1018452(.A(n_132460406), .B(n_132360405), .Z(write_data_31
		[9]));
	notech_nand2 i_1718331(.A(n_132260404), .B(n_132160403), .Z(write_data_30
		[16]));
	notech_nand2 i_1618202(.A(n_132060402), .B(n_131960401), .Z(write_data_29
		[15]));
	notech_nand2 i_118059(.A(n_131860400), .B(n_131760399), .Z(write_data_28
		[0]));
	notech_nand2 i_217676(.A(n_131660398), .B(n_131560397), .Z(write_data_25
		[1]));
	notech_or2 i_4282132(.A(n_352488284), .B(n_352388285), .Z(n_352588283)
		);
	notech_xor2 i_3882131(.A(cs[0]), .B(sav_cs[0]), .Z(n_352488284));
	notech_xor2 i_3782130(.A(cs[1]), .B(sav_cs[1]), .Z(n_352388285));
	notech_ao4 i_41182128(.A(n_351788291), .B(n_27557), .C(n_58661), .D(n_351988289
		), .Z(n_352188287));
	notech_or2 i_6782127(.A(n_351988289), .B(n_27557), .Z(n_352088288));
	notech_ao3 i_69882126(.A(instrc[112]), .B(n_27556), .C(all_cnt[0]), .Z(n_351988289
		));
	notech_and2 i_10382125(.A(n_351788291), .B(n_27557), .Z(n_351888290));
	notech_nand2 i_6482124(.A(n_351688292), .B(all_cnt[1]), .Z(n_351788291)
		);
	notech_nand2 i_6382123(.A(instrc[112]), .B(n_27555), .Z(n_351688292));
	notech_nand2 i_5282122(.A(instrc[115]), .B(n_27558), .Z(n_351588293));
	notech_nand3 i_44282121(.A(n_349488314), .B(n_352588283), .C(n_351188297
		), .Z(n_351488294));
	notech_or4 i_44382120(.A(all_cnt[1]), .B(all_cnt[2]), .C(n_351688292), .D
		(n_26395), .Z(n_351388295));
	notech_ao4 i_11282119(.A(n_352488284), .B(n_352388285), .C(n_349488314),
		 .D(n_26390), .Z(n_351288296));
	notech_or4 i_12282118(.A(n_350888300), .B(n_26390), .C(n_350988299), .D(n_350688302
		), .Z(n_351188297));
	notech_nao3 i_44082117(.A(n_349488314), .B(n_349988309), .C(n_352588283)
		, .Z(n_351088298));
	notech_ao3 i_43682116(.A(n_351788291), .B(n_27557), .C(n_59263), .Z(n_350988299
		));
	notech_ao3 i_43582115(.A(n_59263), .B(n_352088288), .C(n_59272), .Z(n_350888300
		));
	notech_nand3 i_11082114(.A(n_351688292), .B(all_cnt[2]), .C(all_cnt[1]),
		 .Z(n_350788301));
	notech_ao3 i_43782113(.A(n_59272), .B(n_350788301), .C(n_59264), .Z(n_350688302
		));
	notech_nand3 i_12982107(.A(n_352188287), .B(n_349888310), .C(n_349588313
		), .Z(n_350088308));
	notech_nand2 i_41482106(.A(n_351588293), .B(n_350088308), .Z(n_349988309
		));
	notech_or2 i_40982105(.A(n_59264), .B(n_352088288), .Z(n_349888310));
	notech_or2 i_41082102(.A(n_59273), .B(n_351888290), .Z(n_349588313));
	notech_or2 i_3482101(.A(instrc[115]), .B(n_27558), .Z(n_349488314));
	notech_or4 i_121931866(.A(n_275388704), .B(n_2835), .C(n_26612), .D(n_60598
		), .Z(n_349288316));
	notech_ao4 i_127231823(.A(n_27842), .B(n_197114365), .C(n_60484), .D(n_27911
		), .Z(n_348988319));
	notech_ao4 i_127331822(.A(n_57371), .B(n_27394), .C(n_59224), .D(n_28043
		), .Z(n_348888320));
	notech_and2 i_127731818(.A(n_348688322), .B(n_348588323), .Z(n_348788321
		));
	notech_ao4 i_127531820(.A(n_56240), .B(n_27739), .C(n_28011), .D(n_56178
		), .Z(n_348688322));
	notech_ao4 i_127631819(.A(n_27778), .B(n_57343), .C(n_56414), .D(n_27977
		), .Z(n_348588323));
	notech_and4 i_128531810(.A(n_348288326), .B(n_348188327), .C(n_347988329
		), .D(n_347888330), .Z(n_348488324));
	notech_ao4 i_127931816(.A(n_27630), .B(n_56310), .C(n_27945), .D(n_56182
		), .Z(n_348288326));
	notech_ao4 i_128031815(.A(n_56183), .B(n_29142), .C(n_56290), .D(n_27671
		), .Z(n_348188327));
	notech_ao4 i_128231813(.A(n_56186), .B(n_27877), .C(n_56270), .D(n_27707
		), .Z(n_347988329));
	notech_ao4 i_128331812(.A(n_2262), .B(n_27810), .C(n_2261), .D(n_29143),
		 .Z(n_347888330));
	notech_nand2 i_144931666(.A(n_2265), .B(n_29124), .Z(n_347788331));
	notech_or4 i_145831659(.A(fsm[2]), .B(n_60729), .C(n_2582), .D(n_2835), 
		.Z(n_347588333));
	notech_ao4 i_18826(.A(n_336162259), .B(n_60473), .C(n_346788341), .D(n_346688342
		), .Z(n_347488334));
	notech_and4 i_146131656(.A(n_57414), .B(n_57423), .C(n_57382), .D(n_55280
		), .Z(n_347388335));
	notech_ao4 i_146231655(.A(n_59369), .B(n_274688711), .C(n_274588712), .D
		(n_1844), .Z(n_346988339));
	notech_ao4 i_146331654(.A(n_56117), .B(n_2826), .C(n_273288723), .D(n_2221
		), .Z(n_346888340));
	notech_nao3 i_146631651(.A(n_57445), .B(n_26712), .C(n_177560857), .Z(n_346788341
		));
	notech_or4 i_146931649(.A(n_346288346), .B(n_346488344), .C(n_26629), .D
		(n_190388902), .Z(n_346688342));
	notech_nand3 i_147131647(.A(n_2822), .B(n_275788700), .C(n_57434), .Z(n_346488344
		));
	notech_or4 i_147331645(.A(n_26616), .B(n_321731604), .C(n_171560797), .D
		(n_26496), .Z(n_346288346));
	notech_and4 i_147831640(.A(n_54733), .B(n_54769), .C(n_54862), .D(n_345788351
		), .Z(n_346088348));
	notech_and4 i_147731641(.A(n_1958), .B(n_205988854), .C(n_340762305), .D
		(n_58922), .Z(n_345788351));
	notech_ao4 i_147931639(.A(n_2211), .B(n_166160743), .C(tcmp), .D(n_336462262
		), .Z(n_345388355));
	notech_ao3 i_148231636(.A(n_341288364), .B(n_341388363), .C(n_341188365)
		, .Z(n_345088358));
	notech_ao4 i_154131589(.A(first_rep), .B(n_338462282), .C(n_338362281), 
		.D(reps[0]), .Z(n_344688362));
	notech_nand3 i_72932288(.A(reps[0]), .B(reps[1]), .C(n_27146), .Z(n_342662320
		));
	notech_nand3 i_27016(.A(n_26606), .B(n_27558), .C(n_27555), .Z(n_342262316
		));
	notech_nao3 i_22460724(.A(n_28966), .B(n_29010), .C(n_264436799), .Z(n_342162315
		));
	notech_nand2 i_27027(.A(instrc[101]), .B(instrc[103]), .Z(n_342062314)
		);
	notech_or4 i_830550(.A(instrc[103]), .B(instrc[100]), .C(n_28971), .D(instrc
		[101]), .Z(n_341962313));
	notech_nand2 i_27062(.A(instrc[90]), .B(n_334962247), .Z(n_341862312));
	notech_nand2 i_27055(.A(n_57162), .B(n_334862246), .Z(n_341762311));
	notech_nand2 i_27044(.A(instrc[98]), .B(n_334762245), .Z(n_341662310));
	notech_or4 i_70232304(.A(n_54703), .B(n_137960461), .C(n_341762311), .D(n_29040
		), .Z(n_341562309));
	notech_or4 i_70132305(.A(n_341862312), .B(n_29017), .C(n_136660448), .D(n_55089
		), .Z(n_341462308));
	notech_or4 i_68232321(.A(n_336362261), .B(n_26629), .C(n_190388902), .D(n_2792
		), .Z(n_341388363));
	notech_or4 i_68132322(.A(tcmp), .B(n_221961291), .C(n_163260714), .D(n_336262260
		), .Z(n_341288364));
	notech_and4 i_68032323(.A(n_26712), .B(n_26629), .C(n_26776), .D(n_57456
		), .Z(n_341188365));
	notech_or4 i_68532318(.A(n_204788866), .B(tcmp), .C(n_2250), .D(n_273588720
		), .Z(n_341088366));
	notech_nand2 i_68632317(.A(fepc), .B(n_60598), .Z(n_340762305));
	notech_or4 i_10732772(.A(n_2792), .B(n_26629), .C(n_190388902), .D(n_335762255
		), .Z(n_340262300));
	notech_nao3 i_72632289(.A(reps[0]), .B(nZF), .C(reps[1]), .Z(n_338562283
		));
	notech_and3 i_12132758(.A(n_342662320), .B(n_338562283), .C(n_22579221),
		 .Z(n_338462282));
	notech_and2 i_12032759(.A(n_338562283), .B(n_22579221), .Z(n_338362281)
		);
	notech_nao3 i_70532301(.A(n_56414), .B(n_27557), .C(n_2262), .Z(n_338262280
		));
	notech_or4 i_70432302(.A(n_137360455), .B(n_27557), .C(n_341662310), .D(n_29016
		), .Z(n_338162279));
	notech_nand2 i_10632773(.A(n_338262280), .B(n_338162279), .Z(n_338062278
		));
	notech_nao3 i_70332303(.A(all_cnt[0]), .B(n_338062278), .C(all_cnt[1]), 
		.Z(n_337962277));
	notech_or4 i_70032306(.A(n_27557), .B(n_342062314), .C(instrc[100]), .D(n_28971
		), .Z(n_337862276));
	notech_or4 i_69932307(.A(n_221961291), .B(n_28970), .C(instrc[124]), .D(all_cnt
		[2]), .Z(n_337762275));
	notech_nand3 i_69832308(.A(n_56425), .B(n_27557), .C(n_2252), .Z(n_337662274
		));
	notech_or4 i_69732309(.A(n_162960711), .B(n_27557), .C(n_29026), .D(n_29030
		), .Z(n_337562273));
	notech_and2 i_10532774(.A(n_337762275), .B(n_337862276), .Z(n_337462272)
		);
	notech_and2 i_10332776(.A(n_337662274), .B(n_337562273), .Z(n_337262270)
		);
	notech_and3 i_10432775(.A(n_341562309), .B(n_341462308), .C(n_337962277)
		, .Z(n_337062268));
	notech_mux2 i_10232777(.S(all_cnt[1]), .A(n_337462272), .B(n_337262270),
		 .Z(n_336862266));
	notech_ao4 i_10032779(.A(n_337062268), .B(n_335062248), .C(n_342262316),
		 .D(n_336862266), .Z(n_336662264));
	notech_and4 i_10132778(.A(n_2212), .B(n_55811), .C(n_55568), .D(n_55587)
		, .Z(n_336462262));
	notech_ao4 i_9932780(.A(n_26625), .B(n_2594), .C(n_177560857), .D(n_336662264
		), .Z(n_336362261));
	notech_and2 i_9832781(.A(n_55567), .B(n_55597), .Z(n_336262260));
	notech_and2 i_19732709(.A(n_2223), .B(n_54741), .Z(n_336162259));
	notech_ao4 i_67332330(.A(n_274788710), .B(n_55878), .C(n_29130), .D(n_347588333
		), .Z(n_335762255));
	notech_nand3 i_10832771(.A(n_26498), .B(n_59835), .C(n_59188), .Z(n_335662254
		));
	notech_nand3 i_67232331(.A(n_340262300), .B(n_347488334), .C(n_335662254
		), .Z(n_335562253));
	notech_ao4 i_67132332(.A(n_2175), .B(n_347788331), .C(n_2113), .D(n_29187
		), .Z(n_335262250));
	notech_or4 i_107732868(.A(n_2793), .B(n_26629), .C(n_59835), .D(n_60598)
		, .Z(n_335162249));
	notech_nand2 i_98432877(.A(n_26606), .B(n_27558), .Z(n_335062248));
	notech_or4 i_830559(.A(instrc[88]), .B(instrc[89]), .C(n_29014), .D(instrc
		[91]), .Z(n_334962247));
	notech_or4 i_830547(.A(instrc[104]), .B(instrc[105]), .C(n_29008), .D(instrc
		[107]), .Z(n_334862246));
	notech_or4 i_830553(.A(n_29013), .B(instrc[97]), .C(instrc[96]), .D(instrc
		[99]), .Z(n_334762245));
	notech_or4 i_830556(.A(instrc[95]), .B(instrc[92]), .C(n_28972), .D(instrc
		[93]), .Z(n_334662244));
	notech_ao4 i_223933530(.A(n_1910), .B(n_212988815), .C(n_54764), .D(n_29130
		), .Z(n_334588367));
	notech_ao4 i_224033529(.A(n_332388389), .B(n_60474), .C(n_59168), .D(n_332288390
		), .Z(n_334488368));
	notech_and4 i_224333526(.A(n_54894), .B(n_57393), .C(n_305288635), .D(n_334088372
		), .Z(n_334388369));
	notech_and3 i_7235626(.A(n_57388), .B(n_54777), .C(n_328246806), .Z(n_334088372
		));
	notech_ao4 i_224533524(.A(n_272588730), .B(n_275288705), .C(n_2776), .D(n_27146
		), .Z(n_333588377));
	notech_or4 i_224833521(.A(n_2604), .B(n_2601), .C(n_26612), .D(n_2828), 
		.Z(n_333188381));
	notech_or4 i_119434555(.A(n_60540), .B(n_2588), .C(n_2777), .D(n_62403),
		 .Z(n_332888384));
	notech_or4 i_119134558(.A(n_331988393), .B(n_59224), .C(n_29040), .D(n_274788710
		), .Z(n_332488388));
	notech_and4 i_15735570(.A(n_332088392), .B(n_333588377), .C(n_334388369)
		, .D(n_332888384), .Z(n_332388389));
	notech_and2 i_14135571(.A(n_328046808), .B(n_332488388), .Z(n_332288390)
		);
	notech_or4 i_4935649(.A(n_60494), .B(n_1844), .C(n_60563), .D(\opcode[1] 
		), .Z(n_332188391));
	notech_and3 i_7335625(.A(n_57391), .B(n_57423), .C(n_332188391), .Z(n_332088392
		));
	notech_nao3 i_3235666(.A(n_26712), .B(n_273688719), .C(n_275088707), .Z(n_331988393
		));
	notech_and2 i_2935668(.A(n_55226), .B(n_54886), .Z(n_331888394));
	notech_and4 i_140137751(.A(n_331188397), .B(n_331088398), .C(n_327888425
		), .D(n_327988424), .Z(n_3314));
	notech_ao4 i_139837754(.A(n_55726), .B(n_27579), .C(n_54944), .D(nbus_11273
		[14]), .Z(n_331188397));
	notech_ao4 i_139737755(.A(n_54943), .B(\nbus_11276[14] ), .C(n_54902), .D
		(n_29006), .Z(n_331088398));
	notech_ao4 i_123337917(.A(n_354088268), .B(n_82713221), .C(n_354188267),
		 .D(n_82813222), .Z(n_330888400));
	notech_and4 i_123237918(.A(n_330088408), .B(n_327188432), .C(n_327088433
		), .D(n_330488404), .Z(n_330788401));
	notech_and3 i_122837922(.A(n_330288406), .B(n_330188407), .C(n_326788436
		), .Z(n_330488404));
	notech_ao4 i_122637924(.A(n_59188), .B(n_26756), .C(n_59168), .D(n_27533
		), .Z(n_330288406));
	notech_ao4 i_122537925(.A(n_262336778), .B(n_29186), .C(n_262236777), .D
		(n_29185), .Z(n_330188407));
	notech_ao4 i_122937921(.A(n_55308), .B(\nbus_11276[14] ), .C(n_55307), .D
		(nbus_11273[14]), .Z(n_330088408));
	notech_nand3 i_120937941(.A(n_329188417), .B(n_329062243), .C(n_329688412
		), .Z(n_329788411));
	notech_and3 i_120837942(.A(n_329488414), .B(n_329388415), .C(n_325688444
		), .Z(n_329688412));
	notech_ao4 i_120237948(.A(n_262336778), .B(n_29184), .C(n_262236777), .D
		(n_29183), .Z(n_329488414));
	notech_ao4 i_120537945(.A(n_5538), .B(n_27582), .C(n_59168), .D(n_27535)
		, .Z(n_329388415));
	notech_ao4 i_120437946(.A(n_323462238), .B(n_29004), .C(n_354488264), .D
		(\nbus_11276[16] ), .Z(n_329188417));
	notech_ao4 i_120337947(.A(n_353988269), .B(nbus_11273[16]), .C(n_353488274
		), .D(nbus_11326[16]), .Z(n_329062243));
	notech_or2 i_108549170(.A(n_323062234), .B(n_261261640), .Z(n_3288));
	notech_or4 i_1521594(.A(n_5990), .B(n_328088423), .C(n_26407), .D(n_328188422
		), .Z(n_13199));
	notech_nor2 i_139637756(.A(n_55864), .B(n_80913203), .Z(n_328188422));
	notech_nor2 i_139337759(.A(n_271888737), .B(n_54872), .Z(n_328088423));
	notech_nao3 i_139537757(.A(opc_10[14]), .B(n_62413), .C(n_318031567), .Z
		(n_327988424));
	notech_nao3 i_139437758(.A(n_62433), .B(opc[14]), .C(n_318231569), .Z(n_327888425
		));
	notech_nand3 i_1521178(.A(n_330888400), .B(n_330788401), .C(n_326288441)
		, .Z(n_13551));
	notech_or4 i_122237928(.A(n_273588720), .B(n_59281), .C(n_2240), .D(n_272188734
		), .Z(n_327188432));
	notech_nand2 i_122037930(.A(n_55728), .B(opd[14]), .Z(n_327088433));
	notech_or2 i_121937931(.A(n_55427), .B(n_29006), .Z(n_326788436));
	notech_and2 i_93539131(.A(n_55786), .B(n_322662230), .Z(n_55426));
	notech_or2 i_122137929(.A(n_55426), .B(n_271888737), .Z(n_326288441));
	notech_nand3 i_62239129(.A(n_5538), .B(n_323162235), .C(n_322862232), .Z
		(n_55728));
	notech_and2 i_93439130(.A(n_55789), .B(n_322762231), .Z(n_55427));
	notech_and4 i_106239132(.A(n_260561633), .B(n_259661624), .C(n_54781), .D
		(n_55791), .Z(n_55308));
	notech_and4 i_106339133(.A(n_259861626), .B(n_55790), .C(n_260261630), .D
		(n_54893), .Z(n_55307));
	notech_or4 i_1721180(.A(n_326088443), .B(n_329788411), .C(n_326188442), 
		.D(n_323562239), .Z(n_13563));
	notech_nor2 i_120037950(.A(n_323762241), .B(n_272088735), .Z(n_326188442
		));
	notech_ao3 i_120137949(.A(opc_10[16]), .B(n_62415), .C(n_3288), .Z(n_326088443
		));
	notech_nand2 i_119837952(.A(sav_edi[16]), .B(n_60598), .Z(n_325688444)
		);
	notech_and3 i_55149256(.A(n_354288266), .B(n_323162235), .C(n_322862232)
		, .Z(n_323762241));
	notech_and4 i_89049239(.A(n_260561633), .B(n_259661624), .C(n_322662230)
		, .D(n_55979), .Z(n_323662240));
	notech_nor2 i_119937951(.A(n_271988736), .B(n_323662240), .Z(n_323562239
		));
	notech_and4 i_88949240(.A(n_260261630), .B(n_259861626), .C(n_322762231)
		, .D(n_55978), .Z(n_323462238));
	notech_and3 i_4439048(.A(n_317788512), .B(n_319388496), .C(n_55829), .Z(n_323362237
		));
	notech_and4 i_4939043(.A(n_260461632), .B(n_56040), .C(n_55846), .D(n_260161629
		), .Z(n_323262236));
	notech_or4 i_11735(.A(n_59281), .B(n_205088863), .C(n_273588720), .D(n_56112
		), .Z(n_323162235));
	notech_nao3 i_24760602(.A(n_56492), .B(instrc[118]), .C(n_231461383), .Z
		(n_323062234));
	notech_ao4 i_53449260(.A(n_204988864), .B(n_56551), .C(n_2240), .D(n_26226
		), .Z(n_322962233));
	notech_or4 i_151949222(.A(n_59281), .B(n_56573), .C(n_205088863), .D(n_273588720
		), .Z(n_322862232));
	notech_or2 i_173849251(.A(n_322962233), .B(n_266361691), .Z(n_322762231)
		);
	notech_or2 i_167549244(.A(n_322962233), .B(n_259561623), .Z(n_322662230)
		);
	notech_and4 i_159840688(.A(n_322362227), .B(n_322162225), .C(n_294561949
		), .D(n_294861952), .Z(n_322562229));
	notech_ao4 i_159440692(.A(n_262336778), .B(n_29164), .C(n_353488274), .D
		(nbus_11326[18]), .Z(n_322362227));
	notech_ao4 i_159640690(.A(n_354488264), .B(\nbus_11276[18] ), .C(n_323462238
		), .D(n_29165), .Z(n_322162225));
	notech_and4 i_160340683(.A(n_321862222), .B(n_321662220), .C(n_295161955
		), .D(n_295461958), .Z(n_322062224));
	notech_ao4 i_159940687(.A(n_5538), .B(n_27584), .C(n_59188), .D(n_26759)
		, .Z(n_321862222));
	notech_ao4 i_160140685(.A(n_310818885), .B(n_323762241), .C(n_310565422)
		, .D(n_3288), .Z(n_321662220));
	notech_and4 i_160840678(.A(n_321362217), .B(n_321162215), .C(n_295761961
		), .D(n_296061964), .Z(n_321562219));
	notech_ao4 i_160440682(.A(n_262336778), .B(n_29166), .C(n_353488274), .D
		(nbus_11326[19]), .Z(n_321362217));
	notech_ao4 i_160640680(.A(n_354488264), .B(\nbus_11276[19] ), .C(n_323462238
		), .D(n_29167), .Z(n_321162215));
	notech_and4 i_161340673(.A(n_320862212), .B(n_320662210), .C(n_296361967
		), .D(n_296661970), .Z(n_321062214));
	notech_ao4 i_160940677(.A(n_5538), .B(n_27585), .C(n_59188), .D(n_26761)
		, .Z(n_320862212));
	notech_ao4 i_161140675(.A(n_310718884), .B(n_323762241), .C(n_308065397)
		, .D(n_3288), .Z(n_320662210));
	notech_and4 i_161840668(.A(n_320362207), .B(n_320162205), .C(n_296961973
		), .D(n_297261976), .Z(n_320562209));
	notech_ao4 i_161440672(.A(n_262336778), .B(n_29168), .C(n_353488274), .D
		(nbus_11326[20]), .Z(n_320362207));
	notech_ao4 i_161640670(.A(n_354488264), .B(\nbus_11276[20] ), .C(n_323462238
		), .D(n_29169), .Z(n_320162205));
	notech_and4 i_162340663(.A(n_319862202), .B(n_319662200), .C(n_297561979
		), .D(n_297861982), .Z(n_320062204));
	notech_ao4 i_161940667(.A(n_5538), .B(n_27586), .C(n_59188), .D(n_26762)
		, .Z(n_319862202));
	notech_ao4 i_162140665(.A(n_310618883), .B(n_323762241), .C(n_315162155)
		, .D(n_3288), .Z(n_319662200));
	notech_and4 i_162840658(.A(n_319362197), .B(n_319162195), .C(n_298161985
		), .D(n_298461988), .Z(n_319562199));
	notech_ao4 i_162440662(.A(n_262336778), .B(n_29170), .C(n_353488274), .D
		(nbus_11326[21]), .Z(n_319362197));
	notech_and3 i_44165256(.A(n_274788710), .B(n_59926), .C(n_57444), .Z(n_125170570
		));
	notech_ao3 i_86964831(.A(n_26390), .B(imm[16]), .C(n_56121), .Z(n_125270571
		));
	notech_ao4 i_29165401(.A(n_312283097), .B(n_125170570), .C(n_55484), .D(n_125270571
		), .Z(n_126170580));
	notech_nand3 i_41565678(.A(n_274788710), .B(n_59926), .C(n_26612), .Z(n_126470583
		));
	notech_ao4 i_116164541(.A(n_126470583), .B(n_27535), .C(n_207341704), .D
		(n_28627), .Z(n_126570584));
	notech_ao4 i_116064542(.A(n_311683091), .B(nbus_11273[16]), .C(nbus_11326
		[16]), .D(n_311783092), .Z(n_126770586));
	notech_ao3 i_116464539(.A(n_126570584), .B(n_126770586), .C(n_126170580)
		, .Z(n_126870587));
	notech_ao4 i_115864544(.A(n_311383088), .B(n_29287), .C(n_312083095), .D
		(n_28747), .Z(n_126970588));
	notech_ao4 i_115764545(.A(n_311583090), .B(n_29286), .C(n_311483089), .D
		(n_29285), .Z(n_127070589));
	notech_or2 i_42063145(.A(n_54436), .B(n_29063), .Z(n_127270591));
	notech_nand2 i_41563150(.A(opa[4]), .B(n_54665), .Z(n_127970598));
	notech_or2 i_43563130(.A(n_54436), .B(n_29068), .Z(n_128070599));
	notech_nand2 i_43063135(.A(n_54665), .B(opa[6]), .Z(n_128770606));
	notech_ao4 i_124362346(.A(n_144377843), .B(n_54451), .C(n_27568), .D(n_55757
		), .Z(n_128870607));
	notech_ao4 i_124262347(.A(n_316588524), .B(n_254634172), .C(\nbus_11276[6] 
		), .D(n_54664), .Z(n_129070609));
	notech_ao4 i_124062349(.A(n_57352), .B(n_54432), .C(n_316488525), .D(n_254734173
		), .Z(n_129270611));
	notech_and4 i_124162348(.A(n_183578230), .B(n_183478229), .C(n_129270611
		), .D(n_128070599), .Z(n_129470613));
	notech_ao4 i_122862360(.A(n_54451), .B(n_139770716), .C(n_55757), .D(n_27565
		), .Z(n_129570614));
	notech_ao4 i_122762361(.A(n_316288527), .B(n_254634172), .C(n_54664), .D
		(\nbus_11276[4] ), .Z(n_129770616));
	notech_ao4 i_122562363(.A(n_321188478), .B(n_54432), .C(n_316388526), .D
		(n_254734173), .Z(n_129970618));
	notech_and3 i_122662362(.A(n_137970698), .B(n_129970618), .C(n_127270591
		), .Z(n_130170620));
	notech_and4 i_82959781(.A(n_56060), .B(n_56001), .C(n_55995), .D(n_1021)
		, .Z(n_130270621));
	notech_or4 i_86959747(.A(n_59264), .B(n_59273), .C(n_56203), .D(n_36952)
		, .Z(n_130370622));
	notech_nor2 i_67159928(.A(n_161857906), .B(n_182471135), .Z(n_130470623)
		);
	notech_or4 i_66659933(.A(n_56290), .B(n_997), .C(n_55988), .D(n_57350), 
		.Z(n_131170630));
	notech_or4 i_70059899(.A(n_59264), .B(n_59273), .C(n_204788866), .D(n_55085
		), .Z(n_131270631));
	notech_or4 i_71059890(.A(n_59369), .B(n_59926), .C(n_2645), .D(nbus_11326
		[8]), .Z(n_131970638));
	notech_or4 i_70959891(.A(n_59264), .B(n_59273), .C(n_56203), .D(n_157974447
		), .Z(n_132270641));
	notech_or2 i_70459896(.A(n_183771148), .B(\nbus_11276[8] ), .Z(n_132770646
		));
	notech_nor2 i_72759874(.A(n_161857906), .B(n_184071151), .Z(n_132870647)
		);
	notech_or2 i_72259879(.A(n_177771096), .B(\nbus_11276[8] ), .Z(n_133570654
		));
	notech_or2 i_73459867(.A(n_56068), .B(n_55085), .Z(n_133670655));
	notech_or4 i_72859873(.A(n_355988238), .B(n_2349), .C(n_353069302), .D(n_54594
		), .Z(n_134170660));
	notech_nor2 i_72959872(.A(n_54547), .B(\nbus_11276[9] ), .Z(n_134270661)
		);
	notech_ao4 i_159959078(.A(n_352969301), .B(n_364788148), .C(n_54562), .D
		(nbus_11273[9]), .Z(n_134570664));
	notech_ao4 i_159759080(.A(n_54455), .B(n_57349), .C(n_54431), .D(n_29048
		), .Z(n_134770666));
	notech_nand3 i_159859079(.A(n_134770666), .B(n_26240), .C(n_133670655), 
		.Z(n_134970668));
	notech_ao4 i_159359084(.A(n_177971098), .B(nbus_11273[8]), .C(n_54431), 
		.D(n_29045), .Z(n_135070669));
	notech_ao4 i_159259085(.A(n_27571), .B(n_178071099), .C(n_54455), .D(n_57350
		), .Z(n_135270671));
	notech_nand3 i_159559082(.A(n_135070669), .B(n_135270671), .C(n_133570654
		), .Z(n_135370672));
	notech_ao4 i_159059087(.A(n_161957907), .B(n_364788148), .C(n_157974447)
		, .D(n_56068), .Z(n_135470673));
	notech_ao4 i_157859099(.A(n_161857906), .B(n_178871107), .C(n_161957907)
		, .D(n_178971108), .Z(n_135770676));
	notech_ao4 i_157759100(.A(n_183971150), .B(n_27571), .C(nbus_11273[8]), 
		.D(n_183871149), .Z(n_135970678));
	notech_ao4 i_157359103(.A(n_57350), .B(n_54441), .C(n_29045), .D(n_54459
		), .Z(n_136170680));
	notech_and4 i_157659101(.A(n_131970638), .B(n_132270641), .C(n_136170680
		), .D(n_26404), .Z(n_136470683));
	notech_nao3 i_157159105(.A(n_62423), .B(opc[9]), .C(n_142370742), .Z(n_136570684
		));
	notech_ao4 i_156959107(.A(n_352969301), .B(n_182571136), .C(n_263436789)
		, .D(n_136570684), .Z(n_136670685));
	notech_ao4 i_156859108(.A(n_57349), .B(n_54454), .C(n_29048), .D(n_54453
		), .Z(n_136770686));
	notech_ao4 i_156659110(.A(nbus_11273[9]), .B(n_141170730), .C(\nbus_11276[9] 
		), .D(n_141270731), .Z(n_136970688));
	notech_and3 i_156759109(.A(n_136970688), .B(n_26240), .C(n_131270631), .Z
		(n_137170690));
	notech_ao4 i_149259175(.A(n_54453), .B(n_29045), .C(n_161957907), .D(n_182571136
		), .Z(n_137270691));
	notech_ao4 i_149159176(.A(n_183471145), .B(\nbus_11276[8] ), .C(nbus_11273
		[8]), .D(n_26278), .Z(n_137470693));
	notech_nand3 i_149459173(.A(n_131170630), .B(n_137270691), .C(n_137470693
		), .Z(n_137570694));
	notech_ao4 i_148859178(.A(n_157974447), .B(n_54451), .C(n_27571), .D(n_183671147
		), .Z(n_137670695));
	notech_and2 i_67257889(.A(n_140270721), .B(n_140170720), .Z(n_137970698)
		);
	notech_or4 i_90057015(.A(n_1916), .B(n_1023), .C(n_252434150), .D(n_60532
		), .Z(n_138270701));
	notech_nor2 i_90157014(.A(n_54527), .B(n_252434150), .Z(n_138370702));
	notech_or4 i_92756990(.A(n_59264), .B(n_59273), .C(n_56203), .D(n_55580)
		, .Z(n_138470703));
	notech_or4 i_92956988(.A(n_59264), .B(n_59273), .C(n_204788866), .D(n_55580
		), .Z(n_138570704));
	notech_or4 i_74357166(.A(n_56290), .B(n_997), .C(n_56006), .D(n_57351), 
		.Z(n_138670705));
	notech_nao3 i_73857171(.A(opc[7]), .B(n_62401), .C(n_254734173), .Z(n_139370712
		));
	notech_or2 i_27507(.A(n_55837), .B(n_319588494), .Z(n_139770716));
	notech_ao4 i_169556262(.A(n_55810), .B(nbus_11273[4]), .C(n_249134117), 
		.D(n_59926), .Z(n_140170720));
	notech_ao4 i_169456263(.A(n_27523), .B(n_59835), .C(n_55920), .D(n_321188478
		), .Z(n_140270721));
	notech_ao4 i_151956435(.A(n_2679), .B(n_254634172), .C(n_54451), .D(n_251734143
		), .Z(n_140370722));
	notech_ao4 i_151856436(.A(nbus_11273[7]), .B(n_26307), .C(n_54664), .D(\nbus_11276[7] 
		), .Z(n_140570724));
	notech_ao4 i_151556438(.A(n_28983), .B(n_54436), .C(n_55757), .D(n_27570
		), .Z(n_140770726));
	notech_and4 i_151756437(.A(n_174064078), .B(n_173964077), .C(n_138670705
		), .D(n_140770726), .Z(n_140970728));
	notech_nor2 i_255292(.A(n_318931576), .B(n_26305), .Z(n_141070729));
	notech_ao3 i_192760634(.A(n_55073), .B(n_54436), .C(n_45383), .Z(n_141170730
		));
	notech_and3 i_193060633(.A(n_55072), .B(n_45384), .C(n_54432), .Z(n_141270731
		));
	notech_or4 i_120654140(.A(n_59264), .B(n_59273), .C(n_204788866), .D(n_36952
		), .Z(n_141570734));
	notech_or2 i_66554657(.A(n_54453), .B(n_29077), .Z(n_141670735));
	notech_and4 i_189660641(.A(n_56060), .B(n_56006), .C(n_996), .D(n_56000)
		, .Z(n_142370742));
	notech_nor2 i_67354649(.A(n_54453), .B(n_29080), .Z(n_142470743));
	notech_or4 i_66854654(.A(n_263436789), .B(n_28062), .C(n_60511), .D(n_55988
		), .Z(n_143170750));
	notech_nor2 i_68254641(.A(n_54453), .B(n_29084), .Z(n_143270751));
	notech_or4 i_67654646(.A(n_263436789), .B(n_28063), .C(n_60511), .D(n_55988
		), .Z(n_143970758));
	notech_nor2 i_69054633(.A(n_54453), .B(n_29037), .Z(n_144070759));
	notech_or4 i_68554638(.A(n_263436789), .B(n_28064), .C(n_60511), .D(n_55988
		), .Z(n_144770766));
	notech_or2 i_69854625(.A(n_54453), .B(n_29087), .Z(n_144870767));
	notech_or2 i_69354630(.A(n_183471145), .B(\nbus_11276[15] ), .Z(n_145570774
		));
	notech_or4 i_71454609(.A(n_59369), .B(n_2645), .C(n_59927), .D(nbus_11326
		[10]), .Z(n_145670775));
	notech_nao3 i_70954614(.A(opc_10[10]), .B(n_62415), .C(n_178971108), .Z(n_146370782
		));
	notech_ao3 i_72354600(.A(n_26826), .B(opc[11]), .C(n_2645), .Z(n_146470783
		));
	notech_nor2 i_72254601(.A(n_54459), .B(n_29080), .Z(n_146770786));
	notech_ao3 i_71754606(.A(n_62423), .B(opc[11]), .C(n_178871107), .Z(n_147270791
		));
	notech_ao3 i_73254591(.A(n_26826), .B(opc[12]), .C(n_2645), .Z(n_147370792
		));
	notech_nor2 i_73154592(.A(n_54459), .B(n_29084), .Z(n_147670795));
	notech_ao3 i_72654597(.A(n_62423), .B(opc[12]), .C(n_178871107), .Z(n_148170800
		));
	notech_ao3 i_74154582(.A(n_26826), .B(opc[13]), .C(n_2645), .Z(n_148270801
		));
	notech_nor2 i_74054583(.A(n_54459), .B(n_29037), .Z(n_148570804));
	notech_ao3 i_73554588(.A(n_62429), .B(opc[13]), .C(n_178871107), .Z(n_149070809
		));
	notech_or4 i_75054573(.A(n_59369), .B(n_2645), .C(n_59927), .D(nbus_11326
		[15]), .Z(n_149170810));
	notech_or2 i_74954574(.A(n_54459), .B(n_29087), .Z(n_149470813));
	notech_or4 i_74454579(.A(n_59264), .B(n_59273), .C(n_56203), .D(n_363688159
		), .Z(n_149970818));
	notech_nor2 i_77354550(.A(n_54431), .B(n_29080), .Z(n_150070819));
	notech_ao3 i_76854555(.A(n_62423), .B(opc[11]), .C(n_184071151), .Z(n_150770826
		));
	notech_nor2 i_78154542(.A(n_54431), .B(n_29084), .Z(n_150870827));
	notech_ao3 i_77654547(.A(n_62423), .B(opc[12]), .C(n_184071151), .Z(n_151570834
		));
	notech_nor2 i_78954534(.A(n_54431), .B(n_29037), .Z(n_151670835));
	notech_ao3 i_78454539(.A(n_62423), .B(opc[13]), .C(n_184071151), .Z(n_152370842
		));
	notech_or2 i_79954526(.A(n_54431), .B(n_29087), .Z(n_152470843));
	notech_or4 i_79254531(.A(n_204788866), .B(n_56074), .C(n_57293), .D(n_55859
		), .Z(n_153170850));
	notech_or2 i_91954412(.A(n_98113375), .B(nbus_11273[10]), .Z(n_153670855
		));
	notech_mux2 i_198353380(.S(n_59927), .A(n_318431571), .B(n_27529), .Z(n_153770856
		));
	notech_ao4 i_198253381(.A(n_2177), .B(n_57348), .C(n_56034), .D(\nbus_11276[10] 
		), .Z(n_153970858));
	notech_and3 i_43955305(.A(n_153770856), .B(n_153970858), .C(n_153670855)
		, .Z(n_154070859));
	notech_ao4 i_187853481(.A(n_177164109), .B(n_184071151), .C(n_177264110)
		, .D(n_364788148), .Z(n_154170860));
	notech_ao4 i_187753482(.A(n_177971098), .B(nbus_11273[15]), .C(n_178071099
		), .D(n_27581), .Z(n_154370862));
	notech_and3 i_188053479(.A(n_153170850), .B(n_154170860), .C(n_154370862
		), .Z(n_154470863));
	notech_ao4 i_187553484(.A(n_356476400), .B(n_54455), .C(n_177771096), .D
		(\nbus_11276[15] ), .Z(n_154570864));
	notech_ao4 i_187153488(.A(n_166457952), .B(n_364788148), .C(n_187874746)
		, .D(n_56068), .Z(n_154870867));
	notech_ao4 i_187053489(.A(nbus_11273[13]), .B(n_177971098), .C(n_178071099
		), .D(n_27578), .Z(n_155070869));
	notech_nao3 i_187353486(.A(n_154870867), .B(n_155070869), .C(n_152370842
		), .Z(n_155170870));
	notech_ao4 i_186853491(.A(n_57345), .B(n_54455), .C(n_177771096), .D(\nbus_11276[13] 
		), .Z(n_155270871));
	notech_ao4 i_186453495(.A(n_169057978), .B(n_364788148), .C(n_189074758)
		, .D(n_56068), .Z(n_155570874));
	notech_ao4 i_186353496(.A(nbus_11273[12]), .B(n_177971098), .C(n_178071099
		), .D(n_27577), .Z(n_155770876));
	notech_nao3 i_186653493(.A(n_155570874), .B(n_155770876), .C(n_151570834
		), .Z(n_155870877));
	notech_ao4 i_186153498(.A(n_57346), .B(n_54455), .C(n_177771096), .D(\nbus_11276[12] 
		), .Z(n_155970878));
	notech_ao4 i_185753502(.A(n_171658004), .B(n_364788148), .C(n_238768192)
		, .D(n_56068), .Z(n_156270881));
	notech_ao4 i_185653503(.A(n_177971098), .B(nbus_11273[11]), .C(n_178071099
		), .D(n_27576), .Z(n_156470883));
	notech_nao3 i_185953500(.A(n_156270881), .B(n_156470883), .C(n_150770826
		), .Z(n_156570884));
	notech_ao4 i_185453505(.A(n_57347), .B(n_54455), .C(\nbus_11276[11] ), .D
		(n_177771096), .Z(n_156670885));
	notech_ao4 i_183653523(.A(n_177164109), .B(n_178871107), .C(n_177264110)
		, .D(n_178971108), .Z(n_156970888));
	notech_ao4 i_183553524(.A(nbus_11273[15]), .B(n_183871149), .C(n_183971150
		), .D(n_27581), .Z(n_157170890));
	notech_ao4 i_183253527(.A(n_356476400), .B(n_54441), .C(n_183771148), .D
		(\nbus_11276[15] ), .Z(n_157370892));
	notech_and4 i_183453525(.A(n_363088165), .B(n_157370892), .C(n_149170810
		), .D(n_149470813), .Z(n_157670895));
	notech_ao4 i_182853531(.A(n_166457952), .B(n_178971108), .C(n_187874746)
		, .D(n_54439), .Z(n_157770896));
	notech_ao4 i_182753532(.A(nbus_11273[13]), .B(n_183871149), .C(n_27578),
		 .D(n_183971150), .Z(n_157970898));
	notech_ao4 i_182453535(.A(n_57345), .B(n_54441), .C(n_183771148), .D(\nbus_11276[13] 
		), .Z(n_158170900));
	notech_or4 i_182653533(.A(n_188774755), .B(n_148270801), .C(n_148570804)
		, .D(n_26261), .Z(n_158470903));
	notech_ao4 i_182053539(.A(n_169057978), .B(n_178971108), .C(n_189074758)
		, .D(n_54439), .Z(n_158570904));
	notech_ao4 i_181953540(.A(nbus_11273[12]), .B(n_183871149), .C(n_183971150
		), .D(n_27577), .Z(n_158770906));
	notech_ao4 i_181653543(.A(n_57346), .B(n_54441), .C(n_183771148), .D(\nbus_11276[12] 
		), .Z(n_158970908));
	notech_or4 i_181853541(.A(n_189974767), .B(n_147370792), .C(n_147670795)
		, .D(n_26264), .Z(n_159270911));
	notech_ao4 i_181253547(.A(n_171658004), .B(n_178971108), .C(n_238768192)
		, .D(n_54439), .Z(n_159370912));
	notech_ao4 i_181153548(.A(nbus_11273[11]), .B(n_183871149), .C(n_183971150
		), .D(n_27576), .Z(n_159570914));
	notech_ao4 i_180753551(.A(n_57347), .B(n_54441), .C(\nbus_11276[11] ), .D
		(n_183771148), .Z(n_159770916));
	notech_or4 i_181053549(.A(n_239168196), .B(n_146470783), .C(n_146770786)
		, .D(n_26268), .Z(n_160070919));
	notech_or4 i_180553553(.A(n_56492), .B(instrc[118]), .C(n_1976), .D(n_54595
		), .Z(n_160170920));
	notech_ao4 i_180253556(.A(n_54439), .B(n_319431581), .C(n_174358031), .D
		(n_160170920), .Z(n_160270921));
	notech_ao4 i_180153557(.A(\nbus_11276[10] ), .B(n_54564), .C(n_54566), .D
		(nbus_11273[10]), .Z(n_160470923));
	notech_ao4 i_179953559(.A(n_54459), .B(n_29077), .C(n_57348), .D(n_54441
		), .Z(n_160670925));
	notech_and3 i_180053558(.A(n_154070859), .B(n_160670925), .C(n_145670775
		), .Z(n_160870927));
	notech_ao4 i_178853570(.A(n_177264110), .B(n_182571136), .C(n_177164109)
		, .D(n_182471135), .Z(n_160970928));
	notech_ao4 i_178753571(.A(n_183671147), .B(n_27581), .C(nbus_11273[15]),
		 .D(n_26278), .Z(n_161170930));
	notech_and3 i_179053568(.A(n_160970928), .B(n_161170930), .C(n_145570774
		), .Z(n_161270931));
	notech_ao4 i_178553573(.A(n_356476400), .B(n_54454), .C(n_363688159), .D
		(n_54451), .Z(n_161370932));
	notech_ao4 i_178153577(.A(n_187874746), .B(n_54451), .C(n_182471135), .D
		(n_166557953), .Z(n_161670935));
	notech_ao4 i_178053578(.A(nbus_11273[13]), .B(n_26278), .C(n_183471145),
		 .D(\nbus_11276[13] ), .Z(n_161870937));
	notech_nand3 i_178353575(.A(n_144770766), .B(n_161670935), .C(n_161870937
		), .Z(n_161970938));
	notech_ao4 i_177853580(.A(n_57345), .B(n_54454), .C(n_183671147), .D(n_27578
		), .Z(n_162070939));
	notech_ao4 i_177453584(.A(n_189074758), .B(n_54451), .C(n_182471135), .D
		(n_169157979), .Z(n_162370942));
	notech_ao4 i_177353585(.A(nbus_11273[12]), .B(n_26278), .C(\nbus_11276[12] 
		), .D(n_183471145), .Z(n_162570944));
	notech_nand3 i_177653582(.A(n_143970758), .B(n_162370942), .C(n_162570944
		), .Z(n_162670945));
	notech_ao4 i_177153587(.A(n_57346), .B(n_54454), .C(n_183671147), .D(n_27577
		), .Z(n_162770946));
	notech_ao4 i_176753591(.A(n_238768192), .B(n_54451), .C(n_182471135), .D
		(n_171758005), .Z(n_163070949));
	notech_ao4 i_176653592(.A(nbus_11273[11]), .B(n_26278), .C(n_183471145),
		 .D(\nbus_11276[11] ), .Z(n_163270951));
	notech_nand3 i_176953589(.A(n_143170750), .B(n_163070949), .C(n_163270951
		), .Z(n_163370952));
	notech_ao4 i_176453594(.A(n_57347), .B(n_54454), .C(n_183671147), .D(n_27576
		), .Z(n_163470953));
	notech_or4 i_176253596(.A(n_56492), .B(instrc[118]), .C(n_2349), .D(n_142370742
		), .Z(n_163770956));
	notech_ao4 i_176053598(.A(n_54451), .B(n_319431581), .C(n_174358031), .D
		(n_163770956), .Z(n_163870957));
	notech_ao4 i_175953599(.A(n_141170730), .B(nbus_11273[10]), .C(n_174258030
		), .D(n_182571136), .Z(n_163970958));
	notech_ao4 i_175753601(.A(n_57348), .B(n_54454), .C(n_141270731), .D(\nbus_11276[10] 
		), .Z(n_164170960));
	notech_and3 i_175853600(.A(n_154070859), .B(n_164170960), .C(n_141670735
		), .Z(n_164370962));
	notech_or4 i_108350942(.A(n_56203), .B(n_58661), .C(n_2688), .D(n_55837)
		, .Z(n_164470963));
	notech_nao3 i_108150944(.A(n_62423), .B(opc[0]), .C(n_247334099), .Z(n_165170970
		));
	notech_nao3 i_108250943(.A(opc_10[0]), .B(n_62413), .C(n_247234098), .Z(n_165270971
		));
	notech_and4 i_120972(.A(n_41726130), .B(n_166670985), .C(n_164470963), .D
		(n_165270971), .Z(n_16699));
	notech_or4 i_110050925(.A(n_56177), .B(n_58661), .C(n_2688), .D(n_55820)
		, .Z(n_165370972));
	notech_or2 i_109750928(.A(n_55757), .B(n_27561), .Z(n_165870977));
	notech_nao3 i_109850927(.A(n_62433), .B(opc[0]), .C(n_254734173), .Z(n_165970978
		));
	notech_or4 i_109950926(.A(n_56006), .B(n_263436789), .C(n_28051), .D(n_60511
		), .Z(n_166070979));
	notech_and4 i_121036(.A(n_41726130), .B(n_167370992), .C(n_165370972), .D
		(n_166070979), .Z(n_13815));
	notech_ao4 i_108650939(.A(n_26539), .B(n_27561), .C(n_54563), .D(\nbus_11276[0] 
		), .Z(n_166170980));
	notech_ao4 i_108450941(.A(n_2699), .B(n_54458), .C(n_55903), .D(nbus_11326
		[0]), .Z(n_166270981));
	notech_ao4 i_108550940(.A(n_54565), .B(nbus_11273[0]), .C(n_54435), .D(n_28986
		), .Z(n_166370982));
	notech_and4 i_108950936(.A(n_166370982), .B(n_166270981), .C(n_166170980
		), .D(n_165170970), .Z(n_166670985));
	notech_ao4 i_110250923(.A(n_54664), .B(\nbus_11276[0] ), .C(n_26307), .D
		(nbus_11273[0]), .Z(n_166970988));
	notech_ao4 i_110150924(.A(n_54436), .B(n_28986), .C(n_2699), .D(n_54432)
		, .Z(n_167070989));
	notech_and4 i_110550920(.A(n_167070989), .B(n_166970988), .C(n_165870977
		), .D(n_165970978), .Z(n_167370992));
	notech_or2 i_65948532(.A(n_55073), .B(nbus_11273[30]), .Z(n_167870997)
		);
	notech_or2 i_66348528(.A(n_123423221), .B(nbus_11326[30]), .Z(n_167970998
		));
	notech_nand2 i_66048531(.A(n_2701), .B(\regs_13_14[30] ), .Z(n_168070999
		));
	notech_nao3 i_66548527(.A(opc_10[30]), .B(n_62411), .C(n_123623223), .Z(n_168171000
		));
	notech_or4 i_66248529(.A(n_56177), .B(n_58661), .C(n_54367), .D(n_271188744
		), .Z(n_168271001));
	notech_or2 i_66148530(.A(n_2702), .B(n_270988746), .Z(n_168371002));
	notech_nand3 i_3121066(.A(n_101523002), .B(n_168371002), .C(n_168971008)
		, .Z(n_13995));
	notech_ao4 i_66648526(.A(n_181471126), .B(n_27599), .C(n_55072), .D(\nbus_11276[30] 
		), .Z(n_168471003));
	notech_and3 i_66848524(.A(n_168471003), .B(n_167870997), .C(n_167970998)
		, .Z(n_168671005));
	notech_and4 i_67148521(.A(n_168070999), .B(n_168671005), .C(n_168171000)
		, .D(n_168271001), .Z(n_168971008));
	notech_nor2 i_61344777(.A(n_123423221), .B(nbus_11326[23]), .Z(n_169171010
		));
	notech_or2 i_60844782(.A(n_308921976), .B(n_2702), .Z(n_169871017));
	notech_nor2 i_62144769(.A(n_123423221), .B(nbus_11326[25]), .Z(n_169971018
		));
	notech_or4 i_61644774(.A(n_56177), .B(n_58661), .C(n_54367), .D(n_308421971
		), .Z(n_170671025));
	notech_nor2 i_62944761(.A(n_123423221), .B(nbus_11326[26]), .Z(n_170771026
		));
	notech_or4 i_62444766(.A(n_56177), .B(n_58661), .C(n_54367), .D(n_308321970
		), .Z(n_171471033));
	notech_nor2 i_63744753(.A(n_123423221), .B(nbus_11326[27]), .Z(n_171571034
		));
	notech_or4 i_63244758(.A(n_56177), .B(n_58661), .C(n_54367), .D(n_308221969
		), .Z(n_172271041));
	notech_nor2 i_64544745(.A(n_123423221), .B(nbus_11326[28]), .Z(n_172371042
		));
	notech_or2 i_64044750(.A(n_55072), .B(\nbus_11276[28] ), .Z(n_173071049)
		);
	notech_or4 i_82944562(.A(n_60773), .B(n_60726), .C(n_54761), .D(n_29215)
		, .Z(n_173571054));
	notech_ao4 i_185543578(.A(n_59835), .B(n_27548), .C(n_101213406), .D(n_308821975
		), .Z(n_173671055));
	notech_ao4 i_185443579(.A(n_98113375), .B(nbus_11273[25]), .C(n_56057), 
		.D(\nbus_11276[25] ), .Z(n_173871057));
	notech_nand3 i_44045377(.A(n_173671055), .B(n_173871057), .C(n_173571054
		), .Z(n_173971058));
	notech_ao4 i_169343738(.A(n_57330), .B(n_2702), .C(n_307421961), .D(n_56130
		), .Z(n_174071059));
	notech_ao4 i_169243739(.A(n_29219), .B(n_26450), .C(n_55073), .D(nbus_11273
		[28]), .Z(n_174271061));
	notech_nand3 i_169543736(.A(n_174071059), .B(n_174271061), .C(n_173071049
		), .Z(n_174371062));
	notech_ao4 i_169043741(.A(n_343565725), .B(n_123623223), .C(n_57306), .D
		(n_123223219), .Z(n_174471063));
	notech_ao4 i_168643745(.A(n_286061878), .B(n_123623223), .C(n_303621923)
		, .D(n_56126), .Z(n_174771066));
	notech_ao4 i_168543746(.A(n_29154), .B(n_26450), .C(n_308621973), .D(n_2702
		), .Z(n_174971068));
	notech_nand3 i_168843743(.A(n_174771066), .B(n_174971068), .C(n_172271041
		), .Z(n_175071069));
	notech_ao4 i_168343748(.A(n_55073), .B(nbus_11273[27]), .C(n_55072), .D(\nbus_11276[27] 
		), .Z(n_175171070));
	notech_ao4 i_167943752(.A(n_288561889), .B(n_123623223), .C(n_307621963)
		, .D(n_56126), .Z(n_175471073));
	notech_ao4 i_167843753(.A(n_29156), .B(n_26450), .C(n_308721974), .D(n_2702
		), .Z(n_175671075));
	notech_nand3 i_168143750(.A(n_175471073), .B(n_175671075), .C(n_171471033
		), .Z(n_175771076));
	notech_ao4 i_167643755(.A(n_55073), .B(nbus_11273[26]), .C(n_55072), .D(\nbus_11276[26] 
		), .Z(n_175871077));
	notech_ao4 i_167243759(.A(n_268264999), .B(n_123623223), .C(n_56126), .D
		(n_307521962), .Z(n_176171080));
	notech_ao4 i_167143760(.A(n_29215), .B(n_26450), .C(n_308821975), .D(n_2702
		), .Z(n_176371082));
	notech_nand3 i_167443757(.A(n_176171080), .B(n_176371082), .C(n_170671025
		), .Z(n_176471083));
	notech_ao4 i_166943762(.A(n_55073), .B(nbus_11273[25]), .C(n_55072), .D(\nbus_11276[25] 
		), .Z(n_176571084));
	notech_ao4 i_166543766(.A(n_308521972), .B(n_123223219), .C(n_270765024)
		, .D(n_123623223), .Z(n_176871087));
	notech_ao4 i_166443767(.A(n_29152), .B(n_26450), .C(n_27590), .D(n_181471126
		), .Z(n_177071089));
	notech_nand3 i_166743764(.A(n_176871087), .B(n_177071089), .C(n_169871017
		), .Z(n_177171090));
	notech_ao4 i_166243769(.A(nbus_11273[23]), .B(n_55073), .C(n_55072), .D(\nbus_11276[23] 
		), .Z(n_177271091));
	notech_and4 i_5439039(.A(n_323388457), .B(n_322288468), .C(n_56060), .D(n_238758633
		), .Z(n_177571094));
	notech_or2 i_65738455(.A(n_36952), .B(n_56068), .Z(n_177671095));
	notech_and2 i_106139128(.A(n_322088470), .B(n_322988461), .Z(n_177771096
		));
	notech_nor2 i_108938057(.A(n_177971098), .B(nbus_11273[14]), .Z(n_177871097
		));
	notech_and2 i_94839127(.A(n_323088460), .B(n_97522962), .Z(n_177971098)
		);
	notech_and2 i_60239126(.A(n_353465823), .B(n_177671095), .Z(n_178071099)
		);
	notech_nao3 i_109338053(.A(n_62427), .B(opc[14]), .C(n_184071151), .Z(n_178371102
		));
	notech_or2 i_109538051(.A(n_80913203), .B(n_56068), .Z(n_178471103));
	notech_or2 i_109238054(.A(n_271888737), .B(n_54455), .Z(n_178571104));
	notech_nor2 i_109138055(.A(n_54431), .B(n_29006), .Z(n_178671105));
	notech_nor2 i_108838058(.A(n_177771096), .B(\nbus_11276[14] ), .Z(n_178771106
		));
	notech_or4 i_1520954(.A(n_178671105), .B(n_184571156), .C(n_178771106), 
		.D(n_177871097), .Z(n_9063));
	notech_or4 i_135160567(.A(n_56492), .B(instrc[118]), .C(n_1976), .D(n_130270621
		), .Z(n_178871107));
	notech_or4 i_137260564(.A(n_56492), .B(instrc[118]), .C(n_1976), .D(n_55983
		), .Z(n_178971108));
	notech_or2 i_112538022(.A(n_183971150), .B(n_27579), .Z(n_179471113));
	notech_nao3 i_112738020(.A(n_62433), .B(opc[14]), .C(n_178871107), .Z(n_179571114
		));
	notech_nao3 i_112838019(.A(opc_10[14]), .B(n_62415), .C(n_178971108), .Z
		(n_179671115));
	notech_or2 i_112638021(.A(n_54441), .B(n_271888737), .Z(n_179971116));
	notech_or4 i_112938018(.A(n_59264), .B(n_59273), .C(n_56203), .D(n_80913203
		), .Z(n_180371117));
	notech_nao3 i_1520986(.A(n_180371117), .B(n_185471165), .C(n_5990), .Z(n_16783
		));
	notech_or2 i_114538002(.A(n_55072), .B(\nbus_11276[17] ), .Z(n_181171124
		));
	notech_or2 i_114638001(.A(n_2702), .B(n_2700), .Z(n_181371125));
	notech_nand3 i_1821053(.A(n_186171172), .B(n_43426147), .C(n_181371125),
		 .Z(n_13917));
	notech_or4 i_62755360(.A(n_59263), .B(n_59273), .C(n_56177), .D(n_56376)
		, .Z(n_181471126));
	notech_or4 i_115937988(.A(n_204788866), .B(n_58661), .C(n_56376), .D(n_27582
		), .Z(n_181971131));
	notech_nao3 i_116237985(.A(opc_10[16]), .B(n_62415), .C(n_123623223), .Z
		(n_182071132));
	notech_nor2 i_116137986(.A(n_123223219), .B(n_272088735), .Z(n_182171133
		));
	notech_nor2 i_116037987(.A(n_2702), .B(n_271988736), .Z(n_182371134));
	notech_or4 i_1721052(.A(n_82113215), .B(n_182171133), .C(n_182371134), .D
		(n_26279), .Z(n_13911));
	notech_or4 i_1555282(.A(n_56492), .B(instrc[118]), .C(n_2349), .D(n_141070729
		), .Z(n_182471135));
	notech_or4 i_133360570(.A(n_56492), .B(n_56478), .C(n_2349), .D(n_55988)
		, .Z(n_182571136));
	notech_nao3 i_117937971(.A(n_62427), .B(opc[14]), .C(n_182471135), .Z(n_183071141
		));
	notech_or4 i_118037970(.A(n_263436789), .B(n_28065), .C(n_60512), .D(n_55988
		), .Z(n_183171142));
	notech_nor2 i_117837972(.A(n_271888737), .B(n_54454), .Z(n_183271143));
	notech_nor2 i_118137969(.A(n_56126), .B(n_80913203), .Z(n_183371144));
	notech_or4 i_1521050(.A(n_5990), .B(n_183271143), .C(n_26280), .D(n_183371144
		), .Z(n_13899));
	notech_and2 i_94555346(.A(n_55497), .B(n_55072), .Z(n_183471145));
	notech_ao4 i_94455347(.A(n_26591), .B(n_29012), .C(n_318931576), .D(n_26305
		), .Z(n_183571146));
	notech_and2 i_59855359(.A(n_181471126), .B(n_141570734), .Z(n_183671147)
		);
	notech_and2 i_94760678(.A(n_55495), .B(n_55062), .Z(n_183771148));
	notech_and2 i_94660679(.A(n_55064), .B(n_55496), .Z(n_183871149));
	notech_and2 i_60360702(.A(n_55720), .B(n_130370622), .Z(n_183971150));
	notech_or4 i_28346(.A(n_56465), .B(n_355988238), .C(n_177571094), .D(n_29010
		), .Z(n_184071151));
	notech_ao4 i_109638050(.A(n_364788148), .B(n_82713221), .C(n_178071099),
		 .D(n_27579), .Z(n_184171152));
	notech_and3 i_109838048(.A(n_184171152), .B(n_178471103), .C(n_178371102
		), .Z(n_184371154));
	notech_nao3 i_110038046(.A(n_178571104), .B(n_184371154), .C(n_5990), .Z
		(n_184571156));
	notech_ao4 i_113138016(.A(n_183871149), .B(nbus_11273[14]), .C(n_183771148
		), .D(\nbus_11276[14] ), .Z(n_184871159));
	notech_ao4 i_113038017(.A(n_54459), .B(n_29006), .C(n_55903), .D(nbus_11326
		[14]), .Z(n_184971160));
	notech_and3 i_113338014(.A(n_184971160), .B(n_184871159), .C(n_179471113
		), .Z(n_185171162));
	notech_and4 i_113638011(.A(n_179571114), .B(n_185171162), .C(n_179671115
		), .D(n_179971116), .Z(n_185471165));
	notech_ao4 i_114738000(.A(n_123423221), .B(nbus_11326[17]), .C(n_123623223
		), .D(n_63826342), .Z(n_185671167));
	notech_ao4 i_114837999(.A(n_123223219), .B(n_2648), .C(n_181471126), .D(n_27583
		), .Z(n_185871169));
	notech_ao4 i_114937998(.A(n_55073), .B(nbus_11273[17]), .C(n_26450), .D(n_28987
		), .Z(n_185971170));
	notech_and4 i_115237995(.A(n_185971170), .B(n_185871169), .C(n_185671167
		), .D(n_181171124), .Z(n_186171172));
	notech_ao4 i_116437983(.A(n_26450), .B(n_29004), .C(n_55072), .D(\nbus_11276[16] 
		), .Z(n_186371174));
	notech_ao4 i_116337984(.A(n_55073), .B(nbus_11273[16]), .C(n_123423221),
		 .D(nbus_11326[16]), .Z(n_186471175));
	notech_and4 i_116837980(.A(n_181971131), .B(n_186471175), .C(n_186371174
		), .D(n_182071132), .Z(n_186771178));
	notech_ao4 i_118237968(.A(n_183471145), .B(\nbus_11276[14] ), .C(n_54453
		), .D(n_29006), .Z(n_187071181));
	notech_ao4 i_118337967(.A(n_183671147), .B(n_27579), .C(n_26278), .D(nbus_11273
		[14]), .Z(n_187171182));
	notech_and4 i_118637964(.A(n_187171182), .B(n_187071181), .C(n_183171142
		), .D(n_183071141), .Z(n_187471185));
	notech_nand3 i_6835630(.A(n_59188), .B(n_59926), .C(n_195371264), .Z(n_187771188
		));
	notech_or4 i_7435624(.A(n_49223), .B(n_26574), .C(n_26588), .D(n_187971190
		), .Z(n_187871189));
	notech_and2 i_4435654(.A(imm[7]), .B(n_26582), .Z(n_187971190));
	notech_and3 i_12535573(.A(n_199271303), .B(n_339372703), .C(n_199371304)
		, .Z(n_188071191));
	notech_ao4 i_12435574(.A(n_59926), .B(n_188871199), .C(n_2799), .D(nbus_11279
		[1]), .Z(n_188171192));
	notech_and2 i_12335575(.A(n_199271303), .B(n_354872858), .Z(n_188371194)
		);
	notech_and2 i_12235576(.A(n_199271303), .B(n_351972829), .Z(n_188471195)
		);
	notech_and2 i_12135577(.A(n_199271303), .B(n_349072800), .Z(n_188571196)
		);
	notech_and2 i_12035578(.A(n_199271303), .B(n_346172771), .Z(n_188671197)
		);
	notech_and2 i_11935579(.A(n_343272742), .B(n_199271303), .Z(n_188771198)
		);
	notech_and2 i_37735354(.A(n_54899), .B(n_339672706), .Z(n_188871199));
	notech_and2 i_11835580(.A(n_189071201), .B(n_339772707), .Z(n_188971200)
		);
	notech_or4 i_41035322(.A(n_60773), .B(n_60726), .C(n_2798), .D(nbus_11279
		[7]), .Z(n_189071201));
	notech_and2 i_41135321(.A(n_57398), .B(n_57397), .Z(n_189171202));
	notech_ao4 i_11735581(.A(n_2799), .B(nbus_11279[8]), .C(n_2390), .D(n_59917
		), .Z(n_189271203));
	notech_ao4 i_11635582(.A(n_2799), .B(nbus_11279[9]), .C(n_2390), .D(n_59917
		), .Z(n_189471205));
	notech_ao4 i_11535583(.A(n_2799), .B(nbus_11279[10]), .C(n_2390), .D(n_59913
		), .Z(n_189671207));
	notech_ao4 i_11435584(.A(n_2799), .B(nbus_11279[11]), .C(n_2390), .D(n_59913
		), .Z(n_189871209));
	notech_ao4 i_11335585(.A(n_2799), .B(nbus_11279[12]), .C(n_2390), .D(n_59913
		), .Z(n_190071211));
	notech_ao4 i_11235586(.A(n_2799), .B(nbus_11279[14]), .C(n_2390), .D(n_59917
		), .Z(n_190271213));
	notech_ao4 i_11135587(.A(n_2799), .B(nbus_11279[15]), .C(n_2390), .D(n_59917
		), .Z(n_190471215));
	notech_and4 i_11035588(.A(n_55231), .B(n_287372184), .C(n_287272183), .D
		(n_190771218), .Z(n_190671217));
	notech_or4 i_64435089(.A(n_60773), .B(n_60726), .C(n_2798), .D(nbus_11279
		[16]), .Z(n_190771218));
	notech_and4 i_10935589(.A(n_55231), .B(n_287372184), .C(n_287272183), .D
		(n_190971220), .Z(n_190871219));
	notech_or4 i_66635067(.A(n_60773), .B(n_60726), .C(n_2798), .D(nbus_11279
		[17]), .Z(n_190971220));
	notech_and4 i_10835590(.A(n_55231), .B(n_287372184), .C(n_287272183), .D
		(n_191171222), .Z(n_191071221));
	notech_or4 i_68835045(.A(n_60773), .B(n_60726), .C(n_2798), .D(nbus_11279
		[18]), .Z(n_191171222));
	notech_and4 i_10735591(.A(n_55231), .B(n_287372184), .C(n_287272183), .D
		(n_191371224), .Z(n_191271223));
	notech_or4 i_71135023(.A(n_60773), .B(n_60726), .C(n_2798), .D(nbus_11279
		[19]), .Z(n_191371224));
	notech_and4 i_10635592(.A(n_55231), .B(n_287372184), .C(n_287272183), .D
		(n_191571226), .Z(n_191471225));
	notech_or4 i_73535001(.A(n_60773), .B(n_60726), .C(n_2798), .D(nbus_11279
		[20]), .Z(n_191571226));
	notech_and4 i_10535593(.A(n_55231), .B(n_287372184), .C(n_287272183), .D
		(n_191771228), .Z(n_191671227));
	notech_or4 i_75734979(.A(n_60773), .B(n_60726), .C(n_2798), .D(nbus_11279
		[21]), .Z(n_191771228));
	notech_and4 i_10435594(.A(n_55231), .B(n_287372184), .C(n_287272183), .D
		(n_191971230), .Z(n_191871229));
	notech_or4 i_78034957(.A(n_60773), .B(n_60726), .C(n_2798), .D(nbus_11279
		[22]), .Z(n_191971230));
	notech_and4 i_10335595(.A(n_55231), .B(n_287372184), .C(n_287272183), .D
		(n_192171232), .Z(n_192071231));
	notech_or4 i_80334935(.A(n_60775), .B(n_60726), .C(n_2798), .D(nbus_11279
		[23]), .Z(n_192171232));
	notech_and4 i_10235596(.A(n_55231), .B(n_287372184), .C(n_287272183), .D
		(n_192371234), .Z(n_192271233));
	notech_or4 i_82734913(.A(n_60775), .B(n_60726), .C(n_2798), .D(nbus_11279
		[24]), .Z(n_192371234));
	notech_and4 i_10135597(.A(n_55231), .B(n_287372184), .C(n_287272183), .D
		(n_192571236), .Z(n_192471235));
	notech_or4 i_85134891(.A(n_60775), .B(n_60726), .C(n_2798), .D(nbus_11279
		[25]), .Z(n_192571236));
	notech_and4 i_10035598(.A(n_55231), .B(n_287372184), .C(n_287272183), .D
		(n_192771238), .Z(n_192671237));
	notech_or4 i_87434869(.A(n_60775), .B(n_60726), .C(n_2798), .D(nbus_11279
		[26]), .Z(n_192771238));
	notech_and4 i_9935599(.A(n_55231), .B(n_287372184), .C(n_287272183), .D(n_192971240
		), .Z(n_192871239));
	notech_or4 i_89634847(.A(n_60773), .B(n_60729), .C(n_2798), .D(nbus_11279
		[27]), .Z(n_192971240));
	notech_and4 i_9835600(.A(n_56618), .B(n_56609), .C(n_287272183), .D(n_193171242
		), .Z(n_193071241));
	notech_or4 i_91934825(.A(n_60773), .B(n_60731), .C(n_2798), .D(nbus_11279
		[28]), .Z(n_193171242));
	notech_and4 i_9735601(.A(n_56618), .B(n_56609), .C(n_287272183), .D(n_193371244
		), .Z(n_193271243));
	notech_or4 i_94134803(.A(n_60773), .B(n_60731), .C(n_2798), .D(nbus_11279
		[29]), .Z(n_193371244));
	notech_and4 i_9635602(.A(n_56618), .B(n_56609), .C(n_287272183), .D(n_193571246
		), .Z(n_193471245));
	notech_or4 i_96334781(.A(n_60773), .B(n_60731), .C(n_2798), .D(nbus_11279
		[30]), .Z(n_193571246));
	notech_and4 i_9535603(.A(n_56618), .B(n_56609), .C(n_287272183), .D(n_193771248
		), .Z(n_193671247));
	notech_or4 i_98534759(.A(n_60779), .B(n_60731), .C(n_2798), .D(nbus_11279
		[31]), .Z(n_193771248));
	notech_ao4 i_8735611(.A(CFOF_mul), .B(n_57387), .C(n_194471255), .D(n_280472115
		), .Z(n_193871249));
	notech_mux2 i_8835610(.S(n_57430), .A(nCF_shift4box), .B(nCF_shiftbox), 
		.Z(n_193971250));
	notech_and3 i_8935609(.A(n_279772108), .B(n_279672107), .C(n_194971260),
		 .Z(n_194071251));
	notech_and2 i_9035608(.A(n_286272173), .B(n_286172172), .Z(n_194171252)
		);
	notech_and4 i_9135607(.A(n_285772168), .B(n_285072161), .C(n_284272153),
		 .D(n_283572146), .Z(n_194271253));
	notech_ao4 i_6735631(.A(n_57412), .B(n_28123), .C(n_57399), .D(n_26281),
		 .Z(n_194471255));
	notech_or4 i_109334653(.A(n_274988708), .B(n_275488703), .C(n_2586), .D(n_28139
		), .Z(n_194971260));
	notech_ao3 i_8535613(.A(n_57409), .B(n_57410), .C(n_195271263), .Z(n_195171262
		));
	notech_ao4 i_117534574(.A(n_26294), .B(n_26293), .C(n_26605), .D(n_26594
		), .Z(n_195271263));
	notech_nand2 i_117834571(.A(n_328046808), .B(n_195471265), .Z(n_195371264
		));
	notech_or4 i_4835650(.A(n_276288695), .B(n_331988393), .C(n_26296), .D(n_28968
		), .Z(n_195471265));
	notech_and4 i_117934570(.A(n_57409), .B(n_57410), .C(n_57412), .D(n_57399
		), .Z(n_195571266));
	notech_and4 i_118034569(.A(n_57390), .B(n_281972130), .C(n_189171202), .D
		(n_280972120), .Z(n_195671267));
	notech_and3 i_118134568(.A(n_57371), .B(n_60484), .C(n_195971270), .Z(n_195771268
		));
	notech_and2 i_118234567(.A(n_197114365), .B(n_57343), .Z(n_195971270));
	notech_or4 i_118434565(.A(n_60782), .B(n_60731), .C(n_196171272), .D(n_60596
		), .Z(n_196071271));
	notech_ao4 i_8435614(.A(n_59370), .B(n_1911), .C(n_26292), .D(n_57415), 
		.Z(n_196171272));
	notech_nand3 i_18635541(.A(\opa_1[0] ), .B(n_26605), .C(n_26650), .Z(n_196671277
		));
	notech_nand3 i_17935548(.A(n_2771), .B(mul64[0]), .C(n_59835), .Z(n_197371284
		));
	notech_or2 i_17235555(.A(n_2804), .B(\nbus_11276[0] ), .Z(n_198071291)
		);
	notech_or4 i_16535562(.A(n_60782), .B(n_60731), .C(n_57390), .D(nbus_11273
		[8]), .Z(n_198771298));
	notech_or4 i_124935682(.A(fsm[3]), .B(fsm[0]), .C(n_60782), .D(n_188871199
		), .Z(n_199271303));
	notech_or4 i_18735540(.A(n_60782), .B(n_60731), .C(n_2798), .D(nbus_11279
		[0]), .Z(n_199371304));
	notech_nand3 i_21635511(.A(n_26650), .B(\opa_1[1] ), .C(n_26605), .Z(n_199671307
		));
	notech_nand3 i_20935518(.A(n_2771), .B(mul64[1]), .C(n_59835), .Z(n_200371314
		));
	notech_or2 i_20235525(.A(n_2804), .B(n_59753), .Z(n_201071321));
	notech_nand3 i_24635481(.A(n_26650), .B(\opa_1[2] ), .C(n_26605), .Z(n_202571336
		));
	notech_nand3 i_23935488(.A(n_2771), .B(mul64[2]), .C(n_59837), .Z(n_203271343
		));
	notech_or2 i_23235495(.A(n_2804), .B(n_55289), .Z(n_203971350));
	notech_nand3 i_27835450(.A(n_26650), .B(\opa_1[3] ), .C(n_26605), .Z(n_205671367
		));
	notech_nand3 i_27135457(.A(n_2771), .B(mul64[3]), .C(n_59837), .Z(n_206371374
		));
	notech_or2 i_26435464(.A(n_2804), .B(n_55277), .Z(n_207071381));
	notech_nand3 i_31035419(.A(n_26650), .B(\opa_1[4] ), .C(n_26605), .Z(n_208771398
		));
	notech_nand3 i_30335426(.A(n_2771), .B(mul64[4]), .C(n_59837), .Z(n_209471405
		));
	notech_or2 i_29635433(.A(n_2804), .B(\nbus_11276[4] ), .Z(n_210171412)
		);
	notech_nand3 i_34335388(.A(n_26650), .B(\opa_1[5] ), .C(n_26605), .Z(n_211871429
		));
	notech_nand3 i_33635395(.A(n_2771), .B(mul64[5]), .C(n_59837), .Z(n_212571436
		));
	notech_or2 i_32935402(.A(n_2804), .B(n_55375), .Z(n_213271443));
	notech_nand3 i_37435357(.A(n_26650), .B(\opa_1[6] ), .C(n_26605), .Z(n_214971460
		));
	notech_nand3 i_36735364(.A(n_2771), .B(mul64[6]), .C(n_59837), .Z(n_215671467
		));
	notech_nand2 i_36035371(.A(\nbus_14523[6] ), .B(n_26698), .Z(n_216371474
		));
	notech_nand2 i_39235339(.A(\nbus_14523[7] ), .B(n_26698), .Z(n_219471505
		));
	notech_nao3 i_42735306(.A(n_2613), .B(\nbus_14521[8] ), .C(n_2612), .Z(n_222571536
		));
	notech_nao3 i_45735276(.A(n_2613), .B(\nbus_14521[9] ), .C(n_2612), .Z(n_225471565
		));
	notech_nao3 i_48735246(.A(\nbus_14521[10] ), .B(n_2613), .C(n_2612), .Z(n_228371594
		));
	notech_nao3 i_51735216(.A(n_2613), .B(\nbus_14521[11] ), .C(n_2612), .Z(n_231271623
		));
	notech_nao3 i_54735186(.A(n_2613), .B(cr3[12]), .C(n_2612), .Z(n_234171652
		));
	notech_nao3 i_57735156(.A(n_2613), .B(cr3[14]), .C(n_2612), .Z(n_237071681
		));
	notech_nao3 i_60735126(.A(cr2_reg[15]), .B(n_26315), .C(n_2612), .Z(n_239971710
		));
	notech_or4 i_64335090(.A(n_58945), .B(n_2610), .C(n_59917), .D(n_27582),
		 .Z(n_241271723));
	notech_nand2 i_64235091(.A(resa_shiftbox[16]), .B(n_26288), .Z(n_241571726
		));
	notech_nao3 i_63935094(.A(n_2613), .B(cr3[16]), .C(n_2612), .Z(n_241871729
		));
	notech_or2 i_63635097(.A(n_2804), .B(\nbus_11276[16] ), .Z(n_242171732)
		);
	notech_nao3 i_63135102(.A(resa_shift4box[16]), .B(n_26856), .C(n_275988698
		), .Z(n_242671737));
	notech_nao3 i_62835105(.A(resa_arithbox[16]), .B(n_59837), .C(n_57413), 
		.Z(n_242971740));
	notech_or4 i_62535108(.A(n_2773), .B(n_2825), .C(n_59917), .D(nbus_11326
		[0]), .Z(n_243271743));
	notech_or2 i_66435069(.A(n_2784), .B(n_28987), .Z(n_243671747));
	notech_nao3 i_66135072(.A(cr2_reg[17]), .B(n_26315), .C(n_2612), .Z(n_243971750
		));
	notech_nao3 i_65835075(.A(nbus_134[17]), .B(n_59837), .C(n_57412), .Z(n_244271753
		));
	notech_nor2 i_65335080(.A(n_2808), .B(nbus_11326[17]), .Z(n_244771758)
		);
	notech_nao3 i_65035083(.A(resa_arithbox[17]), .B(n_59837), .C(n_57413), 
		.Z(n_245071761));
	notech_or4 i_64735086(.A(n_2773), .B(n_2825), .C(n_59917), .D(nbus_11326
		[1]), .Z(n_245371764));
	notech_or4 i_68735046(.A(n_58945), .B(n_2610), .C(n_59913), .D(n_27584),
		 .Z(n_245471765));
	notech_nand2 i_68635047(.A(resa_shiftbox[18]), .B(n_26288), .Z(n_245771768
		));
	notech_nao3 i_68335050(.A(n_2613), .B(cr3[18]), .C(n_2612), .Z(n_246071771
		));
	notech_or2 i_68035053(.A(n_2804), .B(\nbus_11276[18] ), .Z(n_246371774)
		);
	notech_nao3 i_67535058(.A(resa_shift4box[18]), .B(n_26856), .C(n_275988698
		), .Z(n_246871779));
	notech_nao3 i_67235061(.A(resa_arithbox[18]), .B(n_59837), .C(n_57413), 
		.Z(n_247171782));
	notech_or4 i_66935064(.A(n_2773), .B(n_2825), .C(n_59913), .D(nbus_11326
		[2]), .Z(n_247471785));
	notech_or4 i_71035024(.A(n_58945), .B(n_2610), .C(n_59913), .D(n_27585),
		 .Z(n_247571786));
	notech_nand2 i_70935025(.A(resa_shiftbox[19]), .B(n_26288), .Z(n_247871789
		));
	notech_nao3 i_70635028(.A(n_2613), .B(cr3[19]), .C(n_2612), .Z(n_248171792
		));
	notech_or2 i_70235031(.A(n_2804), .B(\nbus_11276[19] ), .Z(n_248471795)
		);
	notech_nao3 i_69735036(.A(resa_shift4box[19]), .B(n_26856), .C(n_275988698
		), .Z(n_248971800));
	notech_nao3 i_69435039(.A(resa_arithbox[19]), .B(n_59837), .C(n_57413), 
		.Z(n_249271803));
	notech_or4 i_69135042(.A(n_2773), .B(n_2825), .C(n_59913), .D(nbus_11326
		[3]), .Z(n_249571806));
	notech_or4 i_73435002(.A(n_58945), .B(n_2610), .C(n_59913), .D(n_27586),
		 .Z(n_249671807));
	notech_nand2 i_73335003(.A(resa_shiftbox[20]), .B(n_26288), .Z(n_249971810
		));
	notech_nao3 i_73035006(.A(n_2613), .B(cr3[20]), .C(n_2612), .Z(n_250271813
		));
	notech_or2 i_72735009(.A(n_2804), .B(\nbus_11276[20] ), .Z(n_250571816)
		);
	notech_nao3 i_72035014(.A(resa_shift4box[20]), .B(n_26856), .C(n_275988698
		), .Z(n_251071821));
	notech_nao3 i_71735017(.A(resa_arithbox[20]), .B(n_59845), .C(n_57413), 
		.Z(n_251371824));
	notech_or4 i_71435020(.A(n_2773), .B(n_2825), .C(n_59913), .D(nbus_11326
		[4]), .Z(n_251671827));
	notech_or4 i_75634980(.A(n_58945), .B(n_2610), .C(n_59913), .D(n_27588),
		 .Z(n_251771828));
	notech_nand2 i_75534981(.A(resa_shiftbox[21]), .B(n_26288), .Z(n_252071831
		));
	notech_nao3 i_75234984(.A(n_2613), .B(cr3[21]), .C(n_56963), .Z(n_252371834
		));
	notech_or2 i_74934987(.A(n_2804), .B(\nbus_11276[21] ), .Z(n_252671837)
		);
	notech_nao3 i_74434992(.A(resa_shift4box[21]), .B(n_26856), .C(n_275988698
		), .Z(n_253171842));
	notech_nao3 i_74134995(.A(resa_arithbox[21]), .B(n_59865), .C(n_57413), 
		.Z(n_253471845));
	notech_or4 i_73834998(.A(n_2773), .B(n_2825), .C(n_59913), .D(nbus_11326
		[5]), .Z(n_253771848));
	notech_or4 i_77934958(.A(n_58945), .B(n_2610), .C(n_59913), .D(n_27589),
		 .Z(n_253871849));
	notech_nand2 i_77834959(.A(resa_shiftbox[22]), .B(n_26288), .Z(n_254171852
		));
	notech_nao3 i_77534962(.A(n_2613), .B(cr3[22]), .C(n_56963), .Z(n_254471855
		));
	notech_or2 i_77134965(.A(n_2804), .B(\nbus_11276[22] ), .Z(n_254771858)
		);
	notech_nao3 i_76634970(.A(resa_shift4box[22]), .B(n_26856), .C(n_275988698
		), .Z(n_255271863));
	notech_nao3 i_76334973(.A(resa_arithbox[22]), .B(n_59865), .C(n_57413), 
		.Z(n_255571866));
	notech_or4 i_76034976(.A(n_2773), .B(n_2825), .C(n_59913), .D(nbus_11326
		[6]), .Z(n_255871869));
	notech_or2 i_80134937(.A(n_2784), .B(n_29152), .Z(n_256271873));
	notech_nao3 i_79834940(.A(cr2_reg[23]), .B(n_26315), .C(n_56963), .Z(n_256571876
		));
	notech_nao3 i_79534943(.A(nbus_134[23]), .B(n_59865), .C(n_57412), .Z(n_256871879
		));
	notech_or2 i_79034948(.A(n_2808), .B(nbus_11326[23]), .Z(n_257371884));
	notech_nao3 i_78734951(.A(resa_arithbox[23]), .B(n_59865), .C(n_57413), 
		.Z(n_257671887));
	notech_or4 i_78434954(.A(n_2773), .B(n_2825), .C(n_59913), .D(nbus_11326
		[7]), .Z(n_257971890));
	notech_or4 i_82634914(.A(n_58945), .B(n_2610), .C(n_59918), .D(n_27592),
		 .Z(n_258071891));
	notech_nand2 i_82534915(.A(resa_shiftbox[24]), .B(n_26288), .Z(n_258371894
		));
	notech_nao3 i_82134918(.A(n_2613), .B(cr3[24]), .C(n_56963), .Z(n_258671897
		));
	notech_or2 i_81834921(.A(n_2804), .B(\nbus_11276[24] ), .Z(n_258971900)
		);
	notech_nao3 i_81234926(.A(resa_shift4box[24]), .B(n_26856), .C(n_275988698
		), .Z(n_259471905));
	notech_nao3 i_80934929(.A(resa_arithbox[24]), .B(n_59865), .C(n_57413), 
		.Z(n_259771908));
	notech_or4 i_80634932(.A(n_2825), .B(n_2773), .C(n_59918), .D(nbus_11326
		[8]), .Z(n_260071911));
	notech_or4 i_85034892(.A(n_58945), .B(n_2610), .C(n_59918), .D(n_27593),
		 .Z(n_260171912));
	notech_nand2 i_84934893(.A(resa_shiftbox[25]), .B(n_26288), .Z(n_260471915
		));
	notech_nao3 i_84634896(.A(n_2613), .B(cr3[25]), .C(n_56963), .Z(n_260771918
		));
	notech_or2 i_84334899(.A(n_2804), .B(\nbus_11276[25] ), .Z(n_261071921)
		);
	notech_nao3 i_83734904(.A(resa_shift4box[25]), .B(n_26856), .C(n_275988698
		), .Z(n_261571926));
	notech_nao3 i_83434907(.A(resa_arithbox[25]), .B(n_59865), .C(n_57413), 
		.Z(n_261871929));
	notech_or4 i_83034910(.A(n_2773), .B(n_2825), .C(n_59918), .D(nbus_11326
		[9]), .Z(n_262171932));
	notech_or4 i_87334870(.A(n_58945), .B(n_2610), .C(n_59918), .D(n_27594),
		 .Z(n_262271933));
	notech_nand2 i_87134871(.A(resa_shiftbox[26]), .B(n_26288), .Z(n_262571936
		));
	notech_nao3 i_86834874(.A(n_2613), .B(cr3[26]), .C(n_56963), .Z(n_262871939
		));
	notech_or2 i_86534877(.A(n_2804), .B(\nbus_11276[26] ), .Z(n_263171942)
		);
	notech_nao3 i_86034882(.A(resa_shift4box[26]), .B(n_26856), .C(n_275988698
		), .Z(n_263671947));
	notech_nao3 i_85734885(.A(resa_arithbox[26]), .B(n_59865), .C(n_57413), 
		.Z(n_263971950));
	notech_or4 i_85434888(.A(n_2773), .B(n_2825), .C(n_59918), .D(nbus_11326
		[10]), .Z(n_264271953));
	notech_or4 i_89534848(.A(n_58945), .B(n_2610), .C(n_59918), .D(n_27595),
		 .Z(n_264371954));
	notech_nand2 i_89434849(.A(resa_shiftbox[27]), .B(n_26288), .Z(n_264671957
		));
	notech_nao3 i_89134852(.A(n_2613), .B(cr3[27]), .C(n_56963), .Z(n_264971960
		));
	notech_or2 i_88834855(.A(n_2804), .B(\nbus_11276[27] ), .Z(n_265271963)
		);
	notech_nao3 i_88334860(.A(resa_shift4box[27]), .B(n_26856), .C(n_275988698
		), .Z(n_265771968));
	notech_nao3 i_88034863(.A(resa_arithbox[27]), .B(n_59865), .C(n_57424), 
		.Z(n_266071971));
	notech_or4 i_87734866(.A(n_2773), .B(n_2825), .C(n_59918), .D(nbus_11326
		[11]), .Z(n_266371974));
	notech_or4 i_91734826(.A(n_58945), .B(n_2610), .C(n_59918), .D(n_27596),
		 .Z(n_266471975));
	notech_nand2 i_91634827(.A(resa_shiftbox[28]), .B(n_26288), .Z(n_266771978
		));
	notech_nao3 i_91334830(.A(n_2613), .B(cr3[28]), .C(n_56963), .Z(n_267071981
		));
	notech_or2 i_91034833(.A(n_56952), .B(\nbus_11276[28] ), .Z(n_267371984)
		);
	notech_nao3 i_90534838(.A(resa_shift4box[28]), .B(n_26856), .C(n_275988698
		), .Z(n_267871989));
	notech_nao3 i_90234841(.A(resa_arithbox[28]), .B(n_59865), .C(n_57424), 
		.Z(n_268171992));
	notech_or4 i_89934844(.A(n_2773), .B(n_58904), .C(n_59918), .D(nbus_11326
		[12]), .Z(n_268471995));
	notech_or4 i_94034804(.A(n_58945), .B(n_2610), .C(n_59918), .D(n_27597),
		 .Z(n_268571996));
	notech_nand2 i_93934805(.A(resa_shiftbox[29]), .B(n_26288), .Z(n_268871999
		));
	notech_nao3 i_93634808(.A(n_2613), .B(cr3[29]), .C(n_56963), .Z(n_269172002
		));
	notech_or2 i_93334811(.A(n_56952), .B(\nbus_11276[29] ), .Z(n_269472005)
		);
	notech_nao3 i_92834816(.A(resa_shift4box[29]), .B(n_26856), .C(n_275988698
		), .Z(n_269972010));
	notech_nao3 i_92534819(.A(resa_arithbox[29]), .B(n_59865), .C(n_57424), 
		.Z(n_270272013));
	notech_or4 i_92234822(.A(n_2773), .B(n_58904), .C(n_59917), .D(nbus_11326
		[13]), .Z(n_270572016));
	notech_or4 i_96234782(.A(n_58945), .B(n_2610), .C(n_59917), .D(n_27599),
		 .Z(n_270672017));
	notech_nand2 i_96134783(.A(resa_shiftbox[30]), .B(n_26288), .Z(n_270972020
		));
	notech_nao3 i_95834786(.A(n_2613), .B(cr3[30]), .C(n_56963), .Z(n_271272023
		));
	notech_or2 i_95534789(.A(n_56952), .B(\nbus_11276[30] ), .Z(n_271572026)
		);
	notech_nao3 i_95034794(.A(resa_shift4box[30]), .B(n_26856), .C(n_275988698
		), .Z(n_272072031));
	notech_nao3 i_94734797(.A(resa_arithbox[30]), .B(n_59854), .C(n_57424), 
		.Z(n_272372034));
	notech_or4 i_94434800(.A(n_2773), .B(n_58904), .C(n_59917), .D(nbus_11326
		[14]), .Z(n_272672037));
	notech_or4 i_98434760(.A(n_58945), .B(n_2610), .C(n_59917), .D(n_27601),
		 .Z(n_272772038));
	notech_nand2 i_98334761(.A(resa_shiftbox[31]), .B(n_26288), .Z(n_273072041
		));
	notech_nao3 i_98034764(.A(n_2613), .B(cr3[31]), .C(n_56963), .Z(n_273372044
		));
	notech_or2 i_97734767(.A(n_56952), .B(\nbus_11276[31] ), .Z(n_273672047)
		);
	notech_nao3 i_97234772(.A(resa_shift4box[31]), .B(n_26856), .C(n_275988698
		), .Z(n_274172052));
	notech_nao3 i_96934775(.A(resa_arithbox[31]), .B(n_59865), .C(n_57424), 
		.Z(n_274472055));
	notech_or4 i_96634778(.A(n_2773), .B(n_58904), .C(n_59917), .D(nbus_11326
		[15]), .Z(n_274772058));
	notech_nao3 i_108534661(.A(nCF_arithbox), .B(n_59854), .C(n_57424), .Z(n_275072061
		));
	notech_nao3 i_108234664(.A(n_57448), .B(nbus_144[16]), .C(n_312083095), 
		.Z(n_275372064));
	notech_nand2 i_107934667(.A(n_55569), .B(n_26289), .Z(n_275672067));
	notech_nand2 i_107634670(.A(n_193971250), .B(n_59918), .Z(n_275972070)
		);
	notech_nand3 i_109134655(.A(nbus_135[16]), .B(n_26605), .C(n_26294), .Z(n_279672107
		));
	notech_nand2 i_109234654(.A(nbus_140[16]), .B(n_26295), .Z(n_279772108)
		);
	notech_or4 i_117434575(.A(n_60780), .B(n_60731), .C(n_60596), .D(n_195171262
		), .Z(n_279872109));
	notech_or4 i_1235674(.A(n_59370), .B(n_60494), .C(n_106813462), .D(n_195771268
		), .Z(n_279972110));
	notech_nand2 i_118334566(.A(n_27146), .B(n_55154), .Z(n_280072111));
	notech_and2 i_34579(.A(n_187771188), .B(n_282272133), .Z(n_280172112));
	notech_or4 i_29524(.A(n_60780), .B(n_60731), .C(n_60596), .D(n_55324), .Z
		(n_280372114));
	notech_nand2 i_635676(.A(n_56112), .B(n_57448), .Z(n_280472115));
	notech_and3 i_223033539(.A(n_2788), .B(n_2787), .C(n_57392), .Z(n_280972120
		));
	notech_ao4 i_4035658(.A(n_273188724), .B(n_2610), .C(n_272588730), .D(n_58945
		), .Z(n_281572126));
	notech_and4 i_222533544(.A(n_281572126), .B(n_334088372), .C(n_57400), .D
		(n_279972110), .Z(n_281872129));
	notech_and4 i_222833541(.A(n_57418), .B(n_54914), .C(n_305088637), .D(n_281872129
		), .Z(n_281972130));
	notech_ao4 i_223733532(.A(n_190388902), .B(n_2190), .C(n_2798), .D(n_60474
		), .Z(n_282272133));
	notech_or4 i_213533634(.A(n_272788728), .B(n_260788756), .C(n_59918), .D
		(n_55245), .Z(n_282672137));
	notech_ao4 i_209833671(.A(n_193871249), .B(n_59918), .C(n_26292), .D(n_282672137
		), .Z(n_282772138));
	notech_ao4 i_212733642(.A(n_28086), .B(n_56667), .C(n_28084), .D(nbus_11273
		[1]), .Z(n_282972140));
	notech_ao4 i_212633643(.A(n_28088), .B(n_56685), .C(n_56658), .D(n_28085
		), .Z(n_283072141));
	notech_ao4 i_212433645(.A(nbus_11273[7]), .B(n_28090), .C(n_28087), .D(nbus_11273
		[4]), .Z(n_283272143));
	notech_ao4 i_212333646(.A(nbus_11273[9]), .B(n_28092), .C(nbus_11273[6])
		, .D(n_28089), .Z(n_283372144));
	notech_and4 i_212933640(.A(n_283372144), .B(n_283272143), .C(n_283072141
		), .D(n_282972140), .Z(n_283572146));
	notech_ao4 i_212033649(.A(nbus_11273[11]), .B(n_28094), .C(nbus_11273[8]
		), .D(n_28091), .Z(n_283672147));
	notech_ao4 i_211933650(.A(nbus_11273[12]), .B(n_28095), .C(n_28093), .D(nbus_11273
		[10]), .Z(n_283772148));
	notech_ao4 i_211733652(.A(nbus_11273[14]), .B(n_28097), .C(nbus_11273[15
		]), .D(n_28098), .Z(n_283972150));
	notech_ao4 i_211633653(.A(nbus_11273[16]), .B(n_28099), .C(nbus_11273[17
		]), .D(n_28100), .Z(n_284072151));
	notech_and4 i_212233647(.A(n_284072151), .B(n_283972150), .C(n_283772148
		), .D(n_283672147), .Z(n_284272153));
	notech_ao4 i_211233657(.A(nbus_11273[18]), .B(n_28101), .C(nbus_11273[19
		]), .D(n_28102), .Z(n_284472155));
	notech_ao4 i_211133658(.A(nbus_11273[20]), .B(n_28103), .C(nbus_11273[21
		]), .D(n_28104), .Z(n_284572156));
	notech_ao4 i_210933660(.A(nbus_11273[22]), .B(n_28105), .C(nbus_11273[23
		]), .D(n_28106), .Z(n_284772158));
	notech_ao4 i_210833661(.A(nbus_11273[24]), .B(n_28107), .C(nbus_11273[25
		]), .D(n_28108), .Z(n_284872159));
	notech_and4 i_211433655(.A(n_284872159), .B(n_284772158), .C(n_284572156
		), .D(n_284472155), .Z(n_285072161));
	notech_ao4 i_210533664(.A(nbus_11273[26]), .B(n_28109), .C(nbus_11273[27
		]), .D(n_28110), .Z(n_285172162));
	notech_ao4 i_210433665(.A(nbus_11273[28]), .B(n_28111), .C(nbus_11273[29
		]), .D(n_28112), .Z(n_285272163));
	notech_ao4 i_210233667(.A(nbus_11273[30]), .B(n_28113), .C(nbus_11273[31
		]), .D(n_28114), .Z(n_285472165));
	notech_ao4 i_210133668(.A(nbus_11273[13]), .B(n_28096), .C(n_28083), .D(nbus_11273
		[0]), .Z(n_285572166));
	notech_and4 i_210733662(.A(n_285572166), .B(n_285472165), .C(n_285272163
		), .D(n_285172162), .Z(n_285772168));
	notech_ao4 i_213233637(.A(n_57412), .B(n_28371), .C(n_57399), .D(n_26290
		), .Z(n_286172172));
	notech_ao4 i_213133638(.A(n_57409), .B(n_28340), .C(n_57410), .D(n_28302
		), .Z(n_286272173));
	notech_ao4 i_209633673(.A(n_305988628), .B(n_194171252), .C(n_305888629)
		, .D(n_194071251), .Z(n_286372174));
	notech_and4 i_210033669(.A(n_275672067), .B(n_286372174), .C(n_282772138
		), .D(n_275972070), .Z(n_286572176));
	notech_ao4 i_209333676(.A(n_304688641), .B(n_28412), .C(n_304588642), .D
		(n_28856), .Z(n_286672177));
	notech_ao4 i_209133678(.A(n_2778), .B(n_29288), .C(n_311983094), .D(n_28768
		), .Z(n_286872179));
	notech_and4 i_209533674(.A(n_286872179), .B(n_286672177), .C(n_275072061
		), .D(n_275372064), .Z(n_287072181));
	notech_and3 i_196933799(.A(n_55393), .B(n_55230), .C(n_55936), .Z(n_287272183
		));
	notech_or4 i_1835670(.A(n_59370), .B(n_272788728), .C(n_2588), .D(n_59917
		), .Z(n_287372184));
	notech_ao4 i_196333805(.A(n_56631), .B(n_29348), .C(n_193671247), .D(nbus_11273
		[31]), .Z(n_287672187));
	notech_ao4 i_196133807(.A(n_2838), .B(n_28252), .C(n_55936), .D(n_28114)
		, .Z(n_287872189));
	notech_and4 i_196533803(.A(n_287872189), .B(n_287672187), .C(n_274472055
		), .D(n_274772058), .Z(n_288072191));
	notech_ao4 i_195833810(.A(n_2810), .B(n_29347), .C(n_2808), .D(nbus_11326
		[31]), .Z(n_288172192));
	notech_ao4 i_195733811(.A(n_2807), .B(n_27198), .C(n_2834), .D(n_28339),
		 .Z(n_288372194));
	notech_and4 i_196633802(.A(n_288172192), .B(n_288372194), .C(n_288072191
		), .D(n_274172052), .Z(n_288572196));
	notech_ao4 i_195333815(.A(n_2805), .B(n_28370), .C(n_2806), .D(n_27369),
		 .Z(n_288672197));
	notech_ao4 i_195133817(.A(n_2803), .B(n_27229), .C(n_2833), .D(n_28301),
		 .Z(n_288872199));
	notech_and4 i_195533813(.A(n_288872199), .B(n_288672197), .C(n_273372044
		), .D(n_273672047), .Z(n_289072201));
	notech_ao4 i_194833820(.A(n_2784), .B(n_28996), .C(n_2785), .D(n_28173),
		 .Z(n_289172202));
	notech_and4 i_195033818(.A(n_2786), .B(n_289172202), .C(n_272772038), .D
		(n_273072041), .Z(n_289472205));
	notech_ao4 i_194333825(.A(n_329546800), .B(n_29346), .C(n_193471245), .D
		(nbus_11273[30]), .Z(n_289672207));
	notech_ao4 i_194133827(.A(n_2838), .B(n_28251), .C(n_55936), .D(n_28113)
		, .Z(n_289872209));
	notech_and4 i_194533823(.A(n_289872209), .B(n_272672037), .C(n_289672207
		), .D(n_272372034), .Z(n_290072211));
	notech_ao4 i_193833830(.A(n_2810), .B(n_29345), .C(n_2808), .D(nbus_11326
		[30]), .Z(n_290172212));
	notech_ao4 i_193733831(.A(n_2807), .B(n_27197), .C(n_2834), .D(n_28338),
		 .Z(n_290372214));
	notech_and4 i_194633822(.A(n_290172212), .B(n_290372214), .C(n_290072211
		), .D(n_272072031), .Z(n_290572216));
	notech_ao4 i_193333835(.A(n_2805), .B(n_28369), .C(n_2806), .D(n_27061),
		 .Z(n_290672217));
	notech_ao4 i_193133837(.A(n_2803), .B(n_27228), .C(n_2833), .D(n_28300),
		 .Z(n_290872219));
	notech_and4 i_193533833(.A(n_290872219), .B(n_290672217), .C(n_271272023
		), .D(n_271572026), .Z(n_291072221));
	notech_ao4 i_192833840(.A(n_2784), .B(n_28997), .C(n_2785), .D(n_28172),
		 .Z(n_291172222));
	notech_and4 i_193033838(.A(n_2786), .B(n_291172222), .C(n_270672017), .D
		(n_270972020), .Z(n_291472225));
	notech_ao4 i_192333845(.A(n_329546800), .B(n_29275), .C(n_193271243), .D
		(nbus_11273[29]), .Z(n_291672227));
	notech_ao4 i_192133847(.A(n_2838), .B(n_28250), .C(n_55936), .D(n_28112)
		, .Z(n_291872229));
	notech_and4 i_192533843(.A(n_291872229), .B(n_270572016), .C(n_291672227
		), .D(n_270272013), .Z(n_292072231));
	notech_ao4 i_191833850(.A(n_2808), .B(nbus_11326[29]), .C(n_2810), .D(n_29344
		), .Z(n_292172232));
	notech_ao4 i_191733851(.A(n_2807), .B(n_27196), .C(n_2834), .D(n_28337),
		 .Z(n_292372234));
	notech_and4 i_192633842(.A(n_292172232), .B(n_292372234), .C(n_292072231
		), .D(n_269972010), .Z(n_292572236));
	notech_ao4 i_191333855(.A(n_2805), .B(n_28368), .C(n_2806), .D(n_27060),
		 .Z(n_292672237));
	notech_ao4 i_191133857(.A(n_2803), .B(n_27227), .C(n_2833), .D(n_28299),
		 .Z(n_292872239));
	notech_and4 i_191533853(.A(n_292872239), .B(n_292672237), .C(n_269172002
		), .D(n_269472005), .Z(n_293072241));
	notech_ao4 i_190833860(.A(n_2784), .B(n_28977), .C(n_2785), .D(n_28171),
		 .Z(n_293172242));
	notech_and4 i_191033858(.A(n_2786), .B(n_293172242), .C(n_268571996), .D
		(n_268871999), .Z(n_293472245));
	notech_ao4 i_190333865(.A(n_329546800), .B(n_29343), .C(n_193071241), .D
		(nbus_11273[28]), .Z(n_293672247));
	notech_ao4 i_190133867(.A(n_2838), .B(n_28249), .C(n_55936), .D(n_28111)
		, .Z(n_293872249));
	notech_and4 i_190533863(.A(n_293872249), .B(n_268471995), .C(n_293672247
		), .D(n_268171992), .Z(n_294072251));
	notech_ao4 i_189833870(.A(n_2808), .B(nbus_11326[28]), .C(n_2810), .D(n_29342
		), .Z(n_294172252));
	notech_ao4 i_189733871(.A(n_2807), .B(n_27195), .C(n_2834), .D(n_28336),
		 .Z(n_294372254));
	notech_and4 i_190633862(.A(n_294172252), .B(n_294372254), .C(n_294072251
		), .D(n_267871989), .Z(n_294572256));
	notech_ao4 i_189333875(.A(n_2805), .B(n_28367), .C(n_2806), .D(n_27059),
		 .Z(n_294672257));
	notech_ao4 i_189133877(.A(n_2803), .B(n_27225), .C(n_2833), .D(n_28298),
		 .Z(n_294872259));
	notech_and4 i_189533873(.A(n_294872259), .B(n_294672257), .C(n_267071981
		), .D(n_267371984), .Z(n_295072261));
	notech_ao4 i_188833880(.A(n_2784), .B(n_29219), .C(n_2785), .D(n_28170),
		 .Z(n_295172262));
	notech_and4 i_189033878(.A(n_2786), .B(n_295172262), .C(n_266471975), .D
		(n_266771978), .Z(n_295472265));
	notech_ao4 i_188333885(.A(n_56631), .B(n_29341), .C(n_192871239), .D(nbus_11273
		[27]), .Z(n_295672267));
	notech_ao4 i_188133887(.A(n_2838), .B(n_28248), .C(n_55936), .D(n_28110)
		, .Z(n_295872269));
	notech_and4 i_188533883(.A(n_295872269), .B(n_266371974), .C(n_295672267
		), .D(n_266071971), .Z(n_296072271));
	notech_ao4 i_187833890(.A(n_2808), .B(nbus_11326[27]), .C(n_2810), .D(n_29340
		), .Z(n_296172272));
	notech_ao4 i_187733891(.A(n_2807), .B(n_27194), .C(n_2834), .D(n_28335),
		 .Z(n_296372274));
	notech_and4 i_188633882(.A(n_296172272), .B(n_296372274), .C(n_296072271
		), .D(n_265771968), .Z(n_296572276));
	notech_ao4 i_187333895(.A(n_2805), .B(n_28366), .C(n_2806), .D(n_27058),
		 .Z(n_296672277));
	notech_ao4 i_187133897(.A(n_2803), .B(n_27224), .C(n_2833), .D(n_28297),
		 .Z(n_296872279));
	notech_and4 i_187533893(.A(n_296872279), .B(n_296672277), .C(n_264971960
		), .D(n_265271963), .Z(n_297072281));
	notech_ao4 i_186733900(.A(n_2784), .B(n_29154), .C(n_2785), .D(n_28169),
		 .Z(n_297172282));
	notech_and4 i_187033898(.A(n_2786), .B(n_297172282), .C(n_264371954), .D
		(n_264671957), .Z(n_297472285));
	notech_ao4 i_186233905(.A(n_56631), .B(n_29339), .C(n_192671237), .D(nbus_11273
		[26]), .Z(n_297672287));
	notech_ao4 i_186033907(.A(n_2838), .B(n_28247), .C(n_55936), .D(n_28109)
		, .Z(n_297872289));
	notech_and4 i_186433903(.A(n_297872289), .B(n_264271953), .C(n_297672287
		), .D(n_263971950), .Z(n_298072291));
	notech_ao4 i_185733910(.A(n_2808), .B(nbus_11326[26]), .C(n_2810), .D(n_29338
		), .Z(n_298172292));
	notech_ao4 i_185633911(.A(n_2807), .B(n_27193), .C(n_2834), .D(n_28334),
		 .Z(n_298372294));
	notech_and4 i_186533902(.A(n_298172292), .B(n_298372294), .C(n_298072291
		), .D(n_263671947), .Z(n_298572296));
	notech_ao4 i_185233915(.A(n_2805), .B(n_28365), .C(n_2806), .D(n_27057),
		 .Z(n_298672297));
	notech_ao4 i_185033917(.A(n_2803), .B(n_27223), .C(n_2833), .D(n_28296),
		 .Z(n_298872299));
	notech_and4 i_185433913(.A(n_298872299), .B(n_298672297), .C(n_262871939
		), .D(n_263171942), .Z(n_299072301));
	notech_ao4 i_184733920(.A(n_2784), .B(n_29156), .C(n_2785), .D(n_28168),
		 .Z(n_299172302));
	notech_and4 i_184933918(.A(n_2786), .B(n_299172302), .C(n_262271933), .D
		(n_262571936), .Z(n_299472305));
	notech_ao4 i_184233925(.A(n_56631), .B(n_29337), .C(n_192471235), .D(nbus_11273
		[25]), .Z(n_299672307));
	notech_ao4 i_184033927(.A(n_2838), .B(n_28246), .C(n_55936), .D(n_28108)
		, .Z(n_299872309));
	notech_and4 i_184433923(.A(n_299872309), .B(n_262171932), .C(n_299672307
		), .D(n_261871929), .Z(n_300072311));
	notech_ao4 i_183733930(.A(n_2808), .B(nbus_11326[25]), .C(n_2810), .D(n_29336
		), .Z(n_300172312));
	notech_ao4 i_183633931(.A(n_2807), .B(n_27192), .C(n_2834), .D(n_28333),
		 .Z(n_300372314));
	notech_and4 i_184533922(.A(n_300172312), .B(n_300372314), .C(n_300072311
		), .D(n_261571926), .Z(n_300572316));
	notech_ao4 i_183233935(.A(n_2805), .B(n_28364), .C(n_2806), .D(n_27056),
		 .Z(n_300672317));
	notech_ao4 i_183033937(.A(n_2803), .B(n_27222), .C(n_2833), .D(n_28295),
		 .Z(n_300872319));
	notech_and4 i_183433933(.A(n_300872319), .B(n_300672317), .C(n_260771918
		), .D(n_261071921), .Z(n_301072321));
	notech_ao4 i_182733940(.A(n_2784), .B(n_29215), .C(n_2785), .D(n_28167),
		 .Z(n_301172322));
	notech_and4 i_182933938(.A(n_2786), .B(n_301172322), .C(n_260171912), .D
		(n_260471915), .Z(n_301472325));
	notech_ao4 i_182233945(.A(n_56631), .B(n_29335), .C(n_192271233), .D(nbus_11273
		[24]), .Z(n_301672327));
	notech_ao4 i_182033947(.A(n_2838), .B(n_28245), .C(n_55936), .D(n_28107)
		, .Z(n_301872329));
	notech_and4 i_182433943(.A(n_301872329), .B(n_260071911), .C(n_301672327
		), .D(n_259771908), .Z(n_302072331));
	notech_ao4 i_181733950(.A(n_2808), .B(nbus_11326[24]), .C(n_2810), .D(n_29334
		), .Z(n_302172332));
	notech_ao4 i_181533951(.A(n_2807), .B(n_27191), .C(n_2834), .D(n_28332),
		 .Z(n_302372334));
	notech_and4 i_182533942(.A(n_302172332), .B(n_302372334), .C(n_302072331
		), .D(n_259471905), .Z(n_302572336));
	notech_ao4 i_181133955(.A(n_2805), .B(n_28363), .C(n_2806), .D(n_27055),
		 .Z(n_302672337));
	notech_ao4 i_180933957(.A(n_2803), .B(n_27221), .C(n_2833), .D(n_28294),
		 .Z(n_302872339));
	notech_and4 i_181333953(.A(n_302872339), .B(n_302672337), .C(n_258671897
		), .D(n_258971900), .Z(n_303072341));
	notech_ao4 i_180633960(.A(n_2784), .B(n_29137), .C(n_2785), .D(n_28166),
		 .Z(n_303172342));
	notech_and4 i_180833958(.A(n_2786), .B(n_303172342), .C(n_258071891), .D
		(n_258371894), .Z(n_303472345));
	notech_ao4 i_180133965(.A(n_56631), .B(n_29333), .C(n_192071231), .D(nbus_11273
		[23]), .Z(n_303672347));
	notech_ao4 i_179933967(.A(n_2838), .B(n_28244), .C(n_55936), .D(n_28106)
		, .Z(n_303872349));
	notech_and4 i_180333963(.A(n_303872349), .B(n_257971890), .C(n_303672347
		), .D(n_257671887), .Z(n_304072351));
	notech_ao4 i_179633970(.A(n_29332), .B(n_2810), .C(n_280088689), .D(n_27590
		), .Z(n_304172352));
	notech_ao4 i_179533971(.A(n_2834), .B(n_28331), .C(n_2809), .D(n_28221),
		 .Z(n_304372354));
	notech_and3 i_179833968(.A(n_304172352), .B(n_304372354), .C(n_257371884
		), .Z(n_304472355));
	notech_ao4 i_179133975(.A(n_2806), .B(n_27054), .C(n_2807), .D(n_27190),
		 .Z(n_304672357));
	notech_ao4 i_178933977(.A(n_2833), .B(n_28293), .C(n_56952), .D(\nbus_11276[23] 
		), .Z(n_304872359));
	notech_and4 i_179333973(.A(n_304872359), .B(n_304672357), .C(n_256571876
		), .D(n_256871879), .Z(n_305072361));
	notech_ao4 i_178633980(.A(n_2785), .B(n_28165), .C(n_2802), .D(n_28203),
		 .Z(n_305172362));
	notech_ao4 i_178533981(.A(n_54899), .B(n_2597), .C(n_2783), .D(n_28196),
		 .Z(n_305372364));
	notech_and4 i_179433972(.A(n_305172362), .B(n_305372364), .C(n_305072361
		), .D(n_256271873), .Z(n_305572366));
	notech_ao4 i_178133985(.A(n_56631), .B(n_29331), .C(n_191871229), .D(nbus_11273
		[22]), .Z(n_305672367));
	notech_ao4 i_177933987(.A(n_2838), .B(n_28243), .C(n_55936), .D(n_28105)
		, .Z(n_305872369));
	notech_and4 i_178333983(.A(n_305872369), .B(n_255871869), .C(n_305672367
		), .D(n_255571866), .Z(n_306072371));
	notech_ao4 i_177633990(.A(n_2808), .B(nbus_11326[22]), .C(n_2810), .D(n_29330
		), .Z(n_306172372));
	notech_ao4 i_177533991(.A(n_2807), .B(n_27189), .C(n_2834), .D(n_28330),
		 .Z(n_306372374));
	notech_and4 i_178433982(.A(n_306172372), .B(n_306372374), .C(n_306072371
		), .D(n_255271863), .Z(n_306572376));
	notech_ao4 i_177133995(.A(n_2805), .B(n_28362), .C(n_2806), .D(n_27053),
		 .Z(n_306672377));
	notech_ao4 i_176933997(.A(n_2803), .B(n_27219), .C(n_2833), .D(n_28292),
		 .Z(n_306872379));
	notech_and4 i_177333993(.A(n_306872379), .B(n_306672377), .C(n_254471855
		), .D(n_254771858), .Z(n_307072381));
	notech_ao4 i_176634000(.A(n_2784), .B(n_29174), .C(n_2785), .D(n_28164),
		 .Z(n_307172382));
	notech_and4 i_176833998(.A(n_2786), .B(n_307172382), .C(n_253871849), .D
		(n_254171852), .Z(n_307472385));
	notech_ao4 i_176134005(.A(n_329546800), .B(n_29329), .C(n_191671227), .D
		(nbus_11273[21]), .Z(n_307672387));
	notech_ao4 i_175934007(.A(n_2838), .B(n_28242), .C(n_55936), .D(n_28104)
		, .Z(n_307872389));
	notech_and4 i_176334003(.A(n_307872389), .B(n_253771848), .C(n_307672387
		), .D(n_253471845), .Z(n_308072391));
	notech_ao4 i_175634010(.A(n_2808), .B(nbus_11326[21]), .C(n_2810), .D(n_29328
		), .Z(n_308172392));
	notech_ao4 i_175534011(.A(n_2807), .B(n_27188), .C(n_2834), .D(n_28329),
		 .Z(n_308372394));
	notech_and4 i_176434002(.A(n_308172392), .B(n_308372394), .C(n_308072391
		), .D(n_253171842), .Z(n_308572396));
	notech_ao4 i_175134015(.A(n_2805), .B(n_28361), .C(n_2806), .D(n_27052),
		 .Z(n_308672397));
	notech_ao4 i_174934017(.A(n_2803), .B(n_27218), .C(n_2833), .D(n_28289),
		 .Z(n_308872399));
	notech_and4 i_175334013(.A(n_308872399), .B(n_308672397), .C(n_252371834
		), .D(n_252671837), .Z(n_309072401));
	notech_ao4 i_174534020(.A(n_2784), .B(n_29172), .C(n_2785), .D(n_28163),
		 .Z(n_309172402));
	notech_and4 i_174834018(.A(n_2786), .B(n_309172402), .C(n_251771828), .D
		(n_252071831), .Z(n_309472405));
	notech_ao4 i_174034025(.A(n_329546800), .B(n_29327), .C(n_191471225), .D
		(nbus_11273[20]), .Z(n_309672407));
	notech_ao4 i_173834027(.A(n_2838), .B(n_28241), .C(n_55936), .D(n_28103)
		, .Z(n_309872409));
	notech_and4 i_174234023(.A(n_309872409), .B(n_251671827), .C(n_309672407
		), .D(n_251371824), .Z(n_310072411));
	notech_ao4 i_173534030(.A(n_2808), .B(nbus_11326[20]), .C(n_2810), .D(n_29326
		), .Z(n_310172412));
	notech_ao4 i_173434031(.A(n_2807), .B(n_27187), .C(n_2834), .D(n_28328),
		 .Z(n_310372414));
	notech_and4 i_174334022(.A(n_310172412), .B(n_310372414), .C(n_310072411
		), .D(n_251071821), .Z(n_310572416));
	notech_ao4 i_172934035(.A(n_2805), .B(n_28360), .C(n_2806), .D(n_27051),
		 .Z(n_310672417));
	notech_ao4 i_172734037(.A(n_2803), .B(n_27217), .C(n_2833), .D(n_28288),
		 .Z(n_310872419));
	notech_and4 i_173134033(.A(n_310872419), .B(n_310672417), .C(n_250271813
		), .D(n_250571816), .Z(n_311072421));
	notech_ao4 i_172434040(.A(n_2784), .B(n_29169), .C(n_2785), .D(n_28162),
		 .Z(n_311172422));
	notech_and4 i_172634038(.A(n_2786), .B(n_311172422), .C(n_249671807), .D
		(n_249971810), .Z(n_311472425));
	notech_ao4 i_171934045(.A(n_329546800), .B(n_29325), .C(n_191271223), .D
		(nbus_11273[19]), .Z(n_311672427));
	notech_ao4 i_171734047(.A(n_2838), .B(n_28240), .C(n_55936), .D(n_28102)
		, .Z(n_311872429));
	notech_and4 i_172134043(.A(n_311872429), .B(n_249571806), .C(n_311672427
		), .D(n_249271803), .Z(n_312072431));
	notech_ao4 i_171434050(.A(n_2808), .B(nbus_11326[19]), .C(n_2810), .D(n_29324
		), .Z(n_312172432));
	notech_ao4 i_171334051(.A(n_2807), .B(n_27186), .C(n_2834), .D(n_28327),
		 .Z(n_312372434));
	notech_and4 i_172234042(.A(n_312172432), .B(n_312372434), .C(n_312072431
		), .D(n_248971800), .Z(n_312572436));
	notech_ao4 i_170934055(.A(n_2805), .B(n_28359), .C(n_2806), .D(n_27050),
		 .Z(n_312672437));
	notech_ao4 i_170734057(.A(n_2803), .B(n_27216), .C(n_2833), .D(n_28287),
		 .Z(n_312872439));
	notech_and4 i_171134053(.A(n_312872439), .B(n_312672437), .C(n_248171792
		), .D(n_248471795), .Z(n_313072441));
	notech_ao4 i_170434060(.A(n_2784), .B(n_29167), .C(n_2785), .D(n_28161),
		 .Z(n_313172442));
	notech_and4 i_170634058(.A(n_2786), .B(n_313172442), .C(n_247571786), .D
		(n_247871789), .Z(n_313472445));
	notech_ao4 i_169934065(.A(n_329546800), .B(n_29323), .C(n_191071221), .D
		(nbus_11273[18]), .Z(n_313672447));
	notech_ao4 i_169734067(.A(n_2838), .B(n_28239), .C(n_55936), .D(n_28101)
		, .Z(n_313872449));
	notech_and4 i_170134063(.A(n_313872449), .B(n_247471785), .C(n_313672447
		), .D(n_247171782), .Z(n_314072451));
	notech_ao4 i_169434070(.A(n_2808), .B(nbus_11326[18]), .C(n_2810), .D(n_29322
		), .Z(n_314172452));
	notech_ao4 i_169334071(.A(n_2807), .B(n_27185), .C(n_2834), .D(n_28326),
		 .Z(n_314372454));
	notech_and4 i_170234062(.A(n_314172452), .B(n_314372454), .C(n_314072451
		), .D(n_246871779), .Z(n_314572456));
	notech_ao4 i_168934075(.A(n_2805), .B(n_28358), .C(n_2806), .D(n_27049),
		 .Z(n_314672457));
	notech_ao4 i_168734077(.A(n_2803), .B(n_27215), .C(n_2833), .D(n_28286),
		 .Z(n_314872459));
	notech_and4 i_169134073(.A(n_314872459), .B(n_314672457), .C(n_246071771
		), .D(n_246371774), .Z(n_315072461));
	notech_ao4 i_168434080(.A(n_2784), .B(n_29165), .C(n_2785), .D(n_28160),
		 .Z(n_315172462));
	notech_and4 i_168634078(.A(n_2786), .B(n_315172462), .C(n_245471765), .D
		(n_245771768), .Z(n_315472465));
	notech_ao4 i_167634085(.A(n_329546800), .B(n_29113), .C(n_190871219), .D
		(nbus_11273[17]), .Z(n_315672467));
	notech_ao4 i_167434087(.A(n_2838), .B(n_28238), .C(n_55936), .D(n_28100)
		, .Z(n_315872469));
	notech_and4 i_167934083(.A(n_315872469), .B(n_245371764), .C(n_315672467
		), .D(n_245071761), .Z(n_316072471));
	notech_ao4 i_167134090(.A(n_2810), .B(n_29321), .C(n_280088689), .D(n_27583
		), .Z(n_316172472));
	notech_ao4 i_167034091(.A(n_2834), .B(n_28325), .C(n_2809), .D(n_28220),
		 .Z(n_316372474));
	notech_ao3 i_167334088(.A(n_316172472), .B(n_316372474), .C(n_244771758)
		, .Z(n_316472475));
	notech_ao4 i_166534095(.A(n_2806), .B(n_27048), .C(n_2807), .D(n_27184),
		 .Z(n_316672477));
	notech_ao4 i_166334097(.A(n_2833), .B(n_28285), .C(n_56952), .D(\nbus_11276[17] 
		), .Z(n_316872479));
	notech_and4 i_166734093(.A(n_316872479), .B(n_316672477), .C(n_243971750
		), .D(n_244271753), .Z(n_317072481));
	notech_ao4 i_166034100(.A(n_2785), .B(n_28159), .C(n_2802), .D(n_28202),
		 .Z(n_317172482));
	notech_ao4 i_165934101(.A(n_2597), .B(n_54899), .C(n_2783), .D(n_28195),
		 .Z(n_317372484));
	notech_and4 i_166834092(.A(n_317172482), .B(n_317372484), .C(n_317072481
		), .D(n_243671747), .Z(n_317572486));
	notech_ao4 i_165534105(.A(n_329546800), .B(n_29320), .C(n_190671217), .D
		(nbus_11273[16]), .Z(n_317672487));
	notech_ao4 i_165334107(.A(n_28237), .B(n_2838), .C(n_55936), .D(n_28099)
		, .Z(n_317872489));
	notech_and4 i_165734103(.A(n_317872489), .B(n_243271743), .C(n_317672487
		), .D(n_242971740), .Z(n_318072491));
	notech_ao4 i_165034110(.A(n_2808), .B(nbus_11326[16]), .C(n_2810), .D(n_29319
		), .Z(n_318172492));
	notech_ao4 i_164934111(.A(n_2807), .B(n_27183), .C(n_2834), .D(n_28324),
		 .Z(n_318372494));
	notech_and4 i_165834102(.A(n_318172492), .B(n_318372494), .C(n_318072491
		), .D(n_242671737), .Z(n_318572496));
	notech_ao4 i_164534115(.A(n_2805), .B(n_28357), .C(n_2806), .D(n_28142),
		 .Z(n_318672497));
	notech_ao4 i_164334117(.A(n_2803), .B(n_27214), .C(n_2833), .D(n_28284),
		 .Z(n_318872499));
	notech_and4 i_164734113(.A(n_318872499), .B(n_318672497), .C(n_241871729
		), .D(n_242171732), .Z(n_319072501));
	notech_ao4 i_164034120(.A(n_2784), .B(n_29004), .C(n_2785), .D(n_28158),
		 .Z(n_319172502));
	notech_and4 i_164234118(.A(n_2786), .B(n_319172502), .C(n_241271723), .D
		(n_241571726), .Z(n_319472505));
	notech_ao4 i_163434125(.A(n_56640), .B(n_28098), .C(n_190471215), .D(nbus_11273
		[15]), .Z(n_319672507));
	notech_ao4 i_163334126(.A(n_55393), .B(nbus_11273[7]), .C(n_56618), .D(n_27570
		), .Z(n_319772508));
	notech_ao4 i_163134128(.A(n_2812), .B(nbus_11273[31]), .C(n_55230), .D(\nbus_11276[7] 
		), .Z(n_319972510));
	notech_ao4 i_163034129(.A(n_56952), .B(\nbus_11276[15] ), .C(n_2795), .D
		(n_28267), .Z(n_320072511));
	notech_and4 i_163734123(.A(n_320072511), .B(n_319972510), .C(n_319772508
		), .D(n_319672507), .Z(n_320272513));
	notech_ao4 i_162734132(.A(n_56932), .B(n_29318), .C(n_56921), .D(nbus_11326
		[15]), .Z(n_320372514));
	notech_ao4 i_162634133(.A(n_56910), .B(n_27181), .C(n_2809), .D(n_28219)
		, .Z(n_320472515));
	notech_ao4 i_162434135(.A(n_2820), .B(\nbus_11276[31] ), .C(n_56972), .D
		(n_27047), .Z(n_320672517));
	notech_and4 i_162934130(.A(n_320672517), .B(n_320472515), .C(n_320372514
		), .D(n_239971710), .Z(n_320872519));
	notech_ao4 i_162034139(.A(n_57177), .B(n_28157), .C(n_2802), .D(n_28200)
		, .Z(n_321072521));
	notech_ao4 i_161934140(.A(n_2783), .B(n_28194), .C(n_57298), .D(n_29087)
		, .Z(n_321172522));
	notech_ao4 i_161734142(.A(n_2794), .B(n_29317), .C(n_280088689), .D(n_27581
		), .Z(n_321372524));
	notech_ao4 i_161634143(.A(n_2818), .B(n_28283), .C(n_2819), .D(n_28386),
		 .Z(n_321472525));
	notech_and4 i_162234137(.A(n_321472525), .B(n_321372524), .C(n_321172522
		), .D(n_321072521), .Z(n_321672527));
	notech_ao4 i_161334146(.A(n_2815), .B(n_28323), .C(n_2817), .D(n_28138),
		 .Z(n_321772528));
	notech_ao4 i_161234147(.A(n_2814), .B(n_28236), .C(n_2816), .D(n_28356),
		 .Z(n_321872529));
	notech_ao4 i_160934149(.A(n_2811), .B(n_28402), .C(n_2813), .D(n_29316),
		 .Z(n_322072531));
	notech_and4 i_161534144(.A(n_2786), .B(n_322072531), .C(n_321872529), .D
		(n_321772528), .Z(n_322272533));
	notech_ao4 i_160534153(.A(n_56640), .B(n_28097), .C(n_190271213), .D(n_56757
		), .Z(n_322472535));
	notech_ao4 i_160434154(.A(n_55393), .B(nbus_11273[6]), .C(n_56618), .D(n_27568
		), .Z(n_322572536));
	notech_ao4 i_160234156(.A(nbus_11273[30]), .B(n_2812), .C(n_55230), .D(\nbus_11276[6] 
		), .Z(n_322772538));
	notech_ao4 i_160134157(.A(n_56952), .B(\nbus_11276[14] ), .C(n_2795), .D
		(n_28266), .Z(n_322872539));
	notech_and4 i_160734151(.A(n_322872539), .B(n_322772538), .C(n_322572536
		), .D(n_322472535), .Z(n_323072541));
	notech_ao4 i_159834160(.A(n_56921), .B(nbus_11326[14]), .C(n_56932), .D(n_29315
		), .Z(n_323172542));
	notech_ao4 i_159734161(.A(n_56910), .B(n_27180), .C(n_2809), .D(n_28218)
		, .Z(n_323272543));
	notech_ao4 i_159534163(.A(n_2803), .B(n_27213), .C(n_56972), .D(n_27046)
		, .Z(n_323472545));
	notech_and4 i_160034158(.A(n_323472545), .B(n_323272543), .C(n_323172542
		), .D(n_237071681), .Z(n_323672547));
	notech_ao4 i_159134167(.A(n_57298), .B(n_29006), .C(n_57177), .D(n_28156
		), .Z(n_323872549));
	notech_ao4 i_159034168(.A(n_280088689), .B(n_27579), .C(n_2783), .D(n_28193
		), .Z(n_323972550));
	notech_ao4 i_158834170(.A(n_2794), .B(n_29314), .C(n_2820), .D(\nbus_11276[30] 
		), .Z(n_324172552));
	notech_ao4 i_158734171(.A(n_2818), .B(n_28282), .C(n_2819), .D(n_28385),
		 .Z(n_324272553));
	notech_and4 i_159334165(.A(n_324272553), .B(n_324172552), .C(n_323972550
		), .D(n_323872549), .Z(n_324472555));
	notech_ao4 i_158434174(.A(n_2815), .B(n_28322), .C(n_2817), .D(n_28137),
		 .Z(n_324572556));
	notech_ao4 i_158334175(.A(n_2814), .B(n_28235), .C(n_2816), .D(n_28355),
		 .Z(n_324672557));
	notech_ao4 i_158134177(.A(n_2811), .B(n_28401), .C(n_2813), .D(n_29313),
		 .Z(n_324872559));
	notech_and4 i_158634172(.A(n_2786), .B(n_324872559), .C(n_324672557), .D
		(n_324572556), .Z(n_325072561));
	notech_ao4 i_157734181(.A(n_56640), .B(n_28095), .C(n_190071211), .D(nbus_11273
		[12]), .Z(n_325272563));
	notech_ao4 i_157634182(.A(n_55393), .B(nbus_11273[4]), .C(n_56618), .D(n_27565
		), .Z(n_325372564));
	notech_ao4 i_157434184(.A(n_2812), .B(nbus_11273[28]), .C(n_55230), .D(\nbus_11276[4] 
		), .Z(n_325572566));
	notech_ao4 i_157334185(.A(n_56932), .B(n_29312), .C(n_2795), .D(n_28265)
		, .Z(n_325672567));
	notech_and4 i_157934179(.A(n_325672567), .B(n_325572566), .C(n_325372564
		), .D(n_325272563), .Z(n_325872569));
	notech_ao4 i_157034188(.A(n_2809), .B(n_28217), .C(n_56921), .D(nbus_11326
		[12]), .Z(n_325972570));
	notech_ao4 i_156934189(.A(n_56972), .B(n_27044), .C(n_56910), .D(n_27178
		), .Z(n_326072571));
	notech_ao4 i_156734191(.A(n_57168), .B(n_27211), .C(n_56952), .D(\nbus_11276[12] 
		), .Z(n_326272573));
	notech_and4 i_157234186(.A(n_326272573), .B(n_326072571), .C(n_325972570
		), .D(n_234171652), .Z(n_326472575));
	notech_ao4 i_156334195(.A(n_57298), .B(n_29084), .C(n_57177), .D(n_28155
		), .Z(n_326672577));
	notech_ao4 i_156234196(.A(n_280088689), .B(n_27577), .C(n_2783), .D(n_28192
		), .Z(n_326772578));
	notech_ao4 i_156034198(.A(n_2794), .B(n_29311), .C(n_2820), .D(\nbus_11276[28] 
		), .Z(n_326972580));
	notech_ao4 i_155934199(.A(n_2818), .B(n_28280), .C(n_2819), .D(n_28384),
		 .Z(n_327072581));
	notech_and4 i_156534193(.A(n_327072581), .B(n_326972580), .C(n_326772578
		), .D(n_326672577), .Z(n_327272583));
	notech_ao4 i_155634202(.A(n_2815), .B(n_28320), .C(n_2817), .D(n_28136),
		 .Z(n_327372584));
	notech_ao4 i_155534203(.A(n_2814), .B(n_28234), .C(n_2816), .D(n_28353),
		 .Z(n_327472585));
	notech_ao4 i_155334205(.A(n_2811), .B(n_28399), .C(n_2813), .D(n_29310),
		 .Z(n_327672587));
	notech_and4 i_155834200(.A(n_2786), .B(n_327672587), .C(n_327472585), .D
		(n_327372584), .Z(n_327872589));
	notech_ao4 i_154934209(.A(n_56640), .B(n_28094), .C(n_189871209), .D(nbus_11273
		[11]), .Z(n_328072591));
	notech_ao4 i_154834210(.A(n_55393), .B(n_56667), .C(n_56618), .D(n_27564
		), .Z(n_328172592));
	notech_ao4 i_154634212(.A(n_2812), .B(nbus_11273[27]), .C(n_55230), .D(n_55277
		), .Z(n_328372594));
	notech_ao4 i_154534213(.A(n_56932), .B(n_29309), .C(n_2795), .D(n_28264)
		, .Z(n_328472595));
	notech_and4 i_155134207(.A(n_328472595), .B(n_328372594), .C(n_328172592
		), .D(n_328072591), .Z(n_328672597));
	notech_ao4 i_154234216(.A(n_2809), .B(n_28216), .C(n_56921), .D(nbus_11326
		[11]), .Z(n_328772598));
	notech_ao4 i_154134217(.A(n_56972), .B(n_27043), .C(n_56910), .D(n_27177
		), .Z(n_328872599));
	notech_ao4 i_153934219(.A(n_57168), .B(n_27210), .C(n_56952), .D(\nbus_11276[11] 
		), .Z(n_329172601));
	notech_and4 i_154434214(.A(n_329172601), .B(n_328872599), .C(n_328772598
		), .D(n_231271623), .Z(n_329372603));
	notech_ao4 i_153534223(.A(n_57298), .B(n_29080), .C(n_57177), .D(n_28154
		), .Z(n_329572605));
	notech_ao4 i_153434224(.A(n_280088689), .B(n_27576), .C(n_2783), .D(n_28191
		), .Z(n_329672606));
	notech_ao4 i_153134226(.A(n_2794), .B(n_29308), .C(n_2820), .D(\nbus_11276[27] 
		), .Z(n_329872608));
	notech_ao4 i_153034227(.A(n_2818), .B(n_28279), .C(n_2819), .D(n_28383),
		 .Z(n_329972609));
	notech_and4 i_153734221(.A(n_329972609), .B(n_329872608), .C(n_329672606
		), .D(n_329572605), .Z(n_330172611));
	notech_ao4 i_152734230(.A(n_2815), .B(n_28318), .C(n_2817), .D(n_28135),
		 .Z(n_330272612));
	notech_ao4 i_152634231(.A(n_2814), .B(n_28233), .C(n_2816), .D(n_28352),
		 .Z(n_330372613));
	notech_ao4 i_152434233(.A(n_2811), .B(n_28398), .C(n_2813), .D(n_29307),
		 .Z(n_330572615));
	notech_and4 i_152934228(.A(n_57312), .B(n_330572615), .C(n_330372613), .D
		(n_330272612), .Z(n_330772617));
	notech_ao4 i_152034237(.A(n_56640), .B(n_28093), .C(n_189671207), .D(nbus_11273
		[10]), .Z(n_330972619));
	notech_ao4 i_151934238(.A(n_55393), .B(n_56658), .C(n_56618), .D(n_55299
		), .Z(n_331072620));
	notech_ao4 i_151734240(.A(n_2812), .B(nbus_11273[26]), .C(n_55230), .D(n_55289
		), .Z(n_331272622));
	notech_ao4 i_151634241(.A(n_56932), .B(n_29306), .C(n_2795), .D(n_28263)
		, .Z(n_331372623));
	notech_and4 i_152234235(.A(n_331372623), .B(n_331272622), .C(n_331072620
		), .D(n_330972619), .Z(n_331572625));
	notech_ao4 i_151234244(.A(n_2809), .B(n_28215), .C(n_56921), .D(nbus_11326
		[10]), .Z(n_331672626));
	notech_ao4 i_151134245(.A(n_56972), .B(n_27042), .C(n_56910), .D(n_27176
		), .Z(n_331772627));
	notech_ao4 i_150934247(.A(n_57168), .B(n_27209), .C(n_56952), .D(\nbus_11276[10] 
		), .Z(n_331972629));
	notech_and4 i_151534242(.A(n_331972629), .B(n_331772627), .C(n_331672626
		), .D(n_228371594), .Z(n_332172631));
	notech_ao4 i_150534251(.A(n_57298), .B(n_29077), .C(n_57177), .D(n_28153
		), .Z(n_332372633));
	notech_ao4 i_150434252(.A(n_280088689), .B(n_27575), .C(n_2783), .D(n_28190
		), .Z(n_332472634));
	notech_ao4 i_150234254(.A(n_2794), .B(n_29305), .C(n_2820), .D(\nbus_11276[26] 
		), .Z(n_332672636));
	notech_ao4 i_150134255(.A(n_2818), .B(n_28278), .C(n_2819), .D(n_28382),
		 .Z(n_332772637));
	notech_and4 i_150734249(.A(n_332772637), .B(n_332672636), .C(n_332472634
		), .D(n_332372633), .Z(n_332972639));
	notech_ao4 i_149834258(.A(n_2815), .B(n_28317), .C(n_2817), .D(n_28134),
		 .Z(n_333072640));
	notech_ao4 i_149734259(.A(n_2814), .B(n_28232), .C(n_2816), .D(n_28351),
		 .Z(n_333172641));
	notech_ao4 i_149534261(.A(n_2811), .B(n_28397), .C(n_2813), .D(n_29304),
		 .Z(n_333372643));
	notech_and4 i_150034256(.A(n_57312), .B(n_333372643), .C(n_333172641), .D
		(n_333072640), .Z(n_333572645));
	notech_ao4 i_149134265(.A(n_56640), .B(n_28092), .C(n_189471205), .D(nbus_11273
		[9]), .Z(n_333772647));
	notech_ao4 i_149034266(.A(n_55393), .B(n_56649), .C(n_56618), .D(n_55331
		), .Z(n_333872648));
	notech_ao4 i_148834268(.A(n_2812), .B(nbus_11273[25]), .C(n_55230), .D(n_59753
		), .Z(n_334072650));
	notech_ao4 i_148734269(.A(n_56952), .B(\nbus_11276[9] ), .C(n_2795), .D(n_28262
		), .Z(n_334172651));
	notech_and4 i_149334263(.A(n_334172651), .B(n_334072650), .C(n_333872648
		), .D(n_333772647), .Z(n_334372653));
	notech_ao4 i_148434272(.A(n_56932), .B(n_29303), .C(n_56921), .D(nbus_11326
		[9]), .Z(n_334472654));
	notech_ao4 i_148334273(.A(n_56910), .B(n_27174), .C(n_2809), .D(n_28214)
		, .Z(n_334572655));
	notech_ao4 i_148134275(.A(n_57168), .B(n_27208), .C(n_56972), .D(n_27041
		), .Z(n_334772657));
	notech_and4 i_148634270(.A(n_334772657), .B(n_334572655), .C(n_334472654
		), .D(n_225471565), .Z(n_334972659));
	notech_ao4 i_147734279(.A(n_57298), .B(n_29048), .C(n_57177), .D(n_28152
		), .Z(n_335172661));
	notech_ao4 i_147634280(.A(n_280088689), .B(n_27574), .C(n_2783), .D(n_28189
		), .Z(n_335272662));
	notech_ao4 i_147434282(.A(n_2794), .B(n_29302), .C(n_2820), .D(\nbus_11276[25] 
		), .Z(n_335472664));
	notech_ao4 i_147334283(.A(n_2818), .B(n_28277), .C(n_2819), .D(n_28381),
		 .Z(n_335572665));
	notech_and4 i_147934277(.A(n_335572665), .B(n_335472664), .C(n_335272662
		), .D(n_335172661), .Z(n_335772667));
	notech_ao4 i_147034286(.A(n_2815), .B(n_28316), .C(n_2817), .D(n_28133),
		 .Z(n_335872668));
	notech_ao4 i_146934287(.A(n_2814), .B(n_28231), .C(n_2816), .D(n_28350),
		 .Z(n_335972669));
	notech_ao4 i_146734289(.A(n_2811), .B(n_28396), .C(n_2813), .D(n_29301),
		 .Z(n_336172671));
	notech_and4 i_147234284(.A(n_57312), .B(n_336172671), .C(n_335972669), .D
		(n_335872668), .Z(n_336372673));
	notech_ao4 i_146334293(.A(n_56640), .B(n_28091), .C(n_189271203), .D(nbus_11273
		[8]), .Z(n_336572675));
	notech_ao4 i_146234294(.A(n_56618), .B(n_27561), .C(n_55393), .D(nbus_11273
		[0]), .Z(n_336672676));
	notech_ao4 i_146034296(.A(n_2812), .B(nbus_11273[24]), .C(n_55230), .D(\nbus_11276[0] 
		), .Z(n_336872678));
	notech_ao4 i_145934297(.A(n_56932), .B(n_29300), .C(n_2795), .D(n_28261)
		, .Z(n_336972679));
	notech_and4 i_146534291(.A(n_336972679), .B(n_336872678), .C(n_336672676
		), .D(n_336572675), .Z(n_337172681));
	notech_ao4 i_145634300(.A(n_2809), .B(n_28213), .C(n_56921), .D(nbus_11326
		[8]), .Z(n_337272682));
	notech_ao4 i_145534301(.A(n_56972), .B(n_27040), .C(n_56910), .D(n_27173
		), .Z(n_337372683));
	notech_ao4 i_145334303(.A(n_57168), .B(n_27207), .C(n_56952), .D(\nbus_11276[8] 
		), .Z(n_337572685));
	notech_and4 i_145834298(.A(n_337572685), .B(n_337372683), .C(n_337272682
		), .D(n_222571536), .Z(n_337772687));
	notech_ao4 i_144934307(.A(n_57298), .B(n_29045), .C(n_57177), .D(n_28151
		), .Z(n_337972689));
	notech_ao4 i_144834308(.A(n_280088689), .B(n_27571), .C(n_2783), .D(n_28188
		), .Z(n_338072690));
	notech_ao4 i_144634310(.A(n_2794), .B(n_29299), .C(n_2820), .D(\nbus_11276[24] 
		), .Z(n_338272692));
	notech_ao4 i_144534311(.A(n_2818), .B(n_28276), .C(n_2819), .D(n_28380),
		 .Z(n_338372693));
	notech_and4 i_145134305(.A(n_338372693), .B(n_338272692), .C(n_338072690
		), .D(n_337972689), .Z(n_338572695));
	notech_ao4 i_144234314(.A(n_2815), .B(n_28315), .C(n_2817), .D(n_28132),
		 .Z(n_338672696));
	notech_ao4 i_144134315(.A(n_2814), .B(n_28230), .C(n_2816), .D(n_28349),
		 .Z(n_338772697));
	notech_ao4 i_143934317(.A(n_2811), .B(n_28395), .C(n_2813), .D(n_29298),
		 .Z(n_338972699));
	notech_and4 i_144434312(.A(n_57312), .B(n_338972699), .C(n_338772697), .D
		(n_338672696), .Z(n_339172701));
	notech_or4 i_77335688(.A(n_272788728), .B(n_260788756), .C(n_59917), .D(n_280472115
		), .Z(n_339372703));
	notech_or4 i_143834318(.A(n_57399), .B(n_59944), .C(n_280472115), .D(opa
		[7]), .Z(n_339472704));
	notech_and4 i_5335645(.A(n_272888727), .B(n_327246816), .C(n_57400), .D(n_281572126
		), .Z(n_339672706));
	notech_ao4 i_143734319(.A(n_339372703), .B(n_327446814), .C(n_339672706)
		, .D(n_59944), .Z(n_339772707));
	notech_ao4 i_143134325(.A(nbus_11273[7]), .B(n_188971200), .C(n_339472704
		), .D(n_26286), .Z(n_339872708));
	notech_or4 i_120035683(.A(n_57412), .B(n_56112), .C(n_59940), .D(n_26594
		), .Z(n_340072710));
	notech_ao4 i_143034326(.A(n_340072710), .B(n_28394), .C(n_56609), .D(\nbus_11276[15] 
		), .Z(n_340172711));
	notech_or4 i_119935684(.A(n_57412), .B(n_26594), .C(n_26605), .D(n_59940
		), .Z(n_340472714));
	notech_or4 i_119735685(.A(n_60752), .B(n_60739), .C(n_60782), .D(n_189171202
		), .Z(n_340572715));
	notech_ao4 i_142834328(.A(n_340572715), .B(n_27570), .C(n_340472714), .D
		(n_28122), .Z(n_340672716));
	notech_ao4 i_142734329(.A(n_55393), .B(nbus_11273[15]), .C(n_56640), .D(n_28090
		), .Z(n_340772717));
	notech_and4 i_143334323(.A(n_340772717), .B(n_340672716), .C(n_340172711
		), .D(n_339872708), .Z(n_340972719));
	notech_ao4 i_142434332(.A(n_56952), .B(\nbus_11276[7] ), .C(n_2795), .D(n_28260
		), .Z(n_341072720));
	notech_ao4 i_142334333(.A(n_56932), .B(n_29297), .C(n_56921), .D(nbus_11326
		[7]), .Z(n_341172721));
	notech_ao4 i_142134335(.A(n_56910), .B(n_27172), .C(n_2809), .D(n_28212)
		, .Z(n_341372723));
	notech_and4 i_142634330(.A(n_341372723), .B(n_341172721), .C(n_341072720
		), .D(n_219471505), .Z(n_341572725));
	notech_ao4 i_141734339(.A(n_2802), .B(n_27238), .C(n_57168), .D(n_27206)
		, .Z(n_341772727));
	notech_ao4 i_141634340(.A(n_57298), .B(n_28983), .C(n_57177), .D(n_28150
		), .Z(n_341872728));
	notech_ao4 i_141434342(.A(n_2820), .B(\nbus_11276[23] ), .C(n_2783), .D(n_28187
		), .Z(n_342072730));
	notech_ao4 i_141334343(.A(n_2819), .B(n_28379), .C(n_2794), .D(n_28569),
		 .Z(n_342172731));
	notech_and4 i_141934337(.A(n_342172731), .B(n_342072730), .C(n_341872728
		), .D(n_341772727), .Z(n_342372733));
	notech_ao4 i_141034346(.A(n_2817), .B(n_28131), .C(n_2818), .D(n_28275),
		 .Z(n_342472734));
	notech_ao4 i_140934347(.A(n_2816), .B(n_28348), .C(n_2815), .D(n_28310),
		 .Z(n_342572735));
	notech_ao4 i_140734349(.A(n_2813), .B(n_29296), .C(n_2814), .D(n_28229),
		 .Z(n_342772737));
	notech_and4 i_141234344(.A(n_57312), .B(n_342772737), .C(n_342572735), .D
		(n_342472734), .Z(n_342972739));
	notech_or4 i_140634350(.A(n_57399), .B(n_59940), .C(n_280472115), .D(opa
		[6]), .Z(n_343172741));
	notech_ao4 i_140534351(.A(n_2799), .B(nbus_11279[6]), .C(n_339372703), .D
		(n_327646812), .Z(n_343272742));
	notech_ao4 i_140134355(.A(nbus_11273[6]), .B(n_188771198), .C(n_343172741
		), .D(n_26285), .Z(n_343372743));
	notech_ao4 i_140034356(.A(n_340072710), .B(n_28393), .C(n_56609), .D(n_55566
		), .Z(n_343472744));
	notech_ao4 i_139834358(.A(n_340572715), .B(n_27568), .C(n_340472714), .D
		(n_28121), .Z(n_343672746));
	notech_ao4 i_139734359(.A(n_55393), .B(n_56757), .C(n_56640), .D(n_28089
		), .Z(n_343772747));
	notech_and4 i_140334353(.A(n_343772747), .B(n_343672746), .C(n_343472744
		), .D(n_343372743), .Z(n_343972749));
	notech_ao4 i_139434362(.A(n_56952), .B(\nbus_11276[6] ), .C(n_2795), .D(n_28259
		), .Z(n_344072750));
	notech_ao4 i_139334363(.A(n_56932), .B(n_29295), .C(n_56921), .D(nbus_11326
		[6]), .Z(n_344172751));
	notech_ao4 i_139134365(.A(n_56910), .B(n_27171), .C(n_28210), .D(n_2809)
		, .Z(n_344372753));
	notech_and4 i_139634360(.A(n_344372753), .B(n_344172751), .C(n_344072750
		), .D(n_216371474), .Z(n_344572755));
	notech_ao4 i_138734369(.A(n_2802), .B(n_27237), .C(n_57168), .D(n_27205)
		, .Z(n_344772757));
	notech_ao4 i_138634370(.A(n_57298), .B(n_29068), .C(n_57177), .D(n_28149
		), .Z(n_344872758));
	notech_ao4 i_138434372(.A(n_2820), .B(\nbus_11276[22] ), .C(n_2783), .D(n_28186
		), .Z(n_345072760));
	notech_and4 i_138934367(.A(n_345072760), .B(n_344872758), .C(n_344772757
		), .D(n_215671467), .Z(n_345272762));
	notech_ao4 i_138134375(.A(n_2818), .B(n_28274), .C(n_2819), .D(n_28378),
		 .Z(n_345372763));
	notech_ao4 i_138034376(.A(n_2815), .B(n_28309), .C(n_2817), .D(n_28130),
		 .Z(n_345472764));
	notech_ao4 i_137834378(.A(n_2814), .B(n_28228), .C(n_2816), .D(n_28347),
		 .Z(n_345672766));
	notech_and4 i_138334373(.A(n_345672766), .B(n_345472764), .C(n_345372763
		), .D(n_214971460), .Z(n_345872768));
	notech_or4 i_137734379(.A(n_57399), .B(n_59944), .C(n_280472115), .D(opa
		[5]), .Z(n_346072770));
	notech_ao4 i_137634380(.A(n_2799), .B(nbus_11279[5]), .C(n_339372703), .D
		(n_3290), .Z(n_346172771));
	notech_ao4 i_137234384(.A(n_56685), .B(n_188671197), .C(n_346072770), .D
		(n_26284), .Z(n_346272772));
	notech_ao4 i_137134385(.A(n_340072710), .B(n_28392), .C(n_56609), .D(\nbus_11276[13] 
		), .Z(n_346372773));
	notech_ao4 i_136934387(.A(n_27566), .B(n_340572715), .C(n_28120), .D(n_340472714
		), .Z(n_346572775));
	notech_ao4 i_136834388(.A(n_55393), .B(nbus_11273[13]), .C(n_56640), .D(n_28088
		), .Z(n_346672776));
	notech_and4 i_137434382(.A(n_346672776), .B(n_346572775), .C(n_346372773
		), .D(n_346272772), .Z(n_346872778));
	notech_ao4 i_136534391(.A(n_56932), .B(n_29294), .C(n_2795), .D(n_28258)
		, .Z(n_346972779));
	notech_ao4 i_136434392(.A(n_2809), .B(n_28209), .C(n_56921), .D(nbus_11326
		[5]), .Z(n_347072780));
	notech_ao4 i_136234394(.A(n_56972), .B(n_27039), .C(n_56910), .D(n_27170
		), .Z(n_347272782));
	notech_and4 i_136734389(.A(n_347272782), .B(n_347072780), .C(n_346972779
		), .D(n_213271443), .Z(n_347472784));
	notech_ao4 i_135834398(.A(n_2802), .B(n_27235), .C(n_57168), .D(n_27204)
		, .Z(n_347672786));
	notech_ao4 i_135734399(.A(n_57298), .B(n_29065), .C(n_57177), .D(n_28148
		), .Z(n_347772787));
	notech_ao4 i_135534401(.A(n_2820), .B(\nbus_11276[21] ), .C(n_2783), .D(n_28182
		), .Z(n_347972789));
	notech_and4 i_136034396(.A(n_347972789), .B(n_347772787), .C(n_347672786
		), .D(n_212571436), .Z(n_348172791));
	notech_ao4 i_135234404(.A(n_2818), .B(n_28273), .C(n_2819), .D(n_28377),
		 .Z(n_348272792));
	notech_ao4 i_135134405(.A(n_2815), .B(n_28308), .C(n_2817), .D(n_28129),
		 .Z(n_348372793));
	notech_ao4 i_134934407(.A(n_2814), .B(n_28227), .C(n_2816), .D(n_28346),
		 .Z(n_348572795));
	notech_and4 i_135434402(.A(n_348572795), .B(n_348372793), .C(n_348272792
		), .D(n_211871429), .Z(n_348772797));
	notech_or4 i_134734408(.A(n_57399), .B(n_59944), .C(n_280472115), .D(opa
		[4]), .Z(n_348972799));
	notech_ao4 i_134634409(.A(n_2799), .B(nbus_11279[4]), .C(n_339372703), .D
		(n_326046828), .Z(n_349072800));
	notech_ao4 i_134234413(.A(nbus_11273[4]), .B(n_188571196), .C(n_26283), 
		.D(n_348972799), .Z(n_349172801));
	notech_ao4 i_134134414(.A(n_340072710), .B(n_28391), .C(n_56609), .D(\nbus_11276[12] 
		), .Z(n_349272802));
	notech_ao4 i_133934416(.A(n_340572715), .B(n_27565), .C(n_340472714), .D
		(n_28119), .Z(n_349472804));
	notech_ao4 i_133834417(.A(n_55393), .B(nbus_11273[12]), .C(n_55936), .D(n_28087
		), .Z(n_349572805));
	notech_and4 i_134434411(.A(n_349572805), .B(n_349472804), .C(n_349272802
		), .D(n_349172801), .Z(n_349772807));
	notech_ao4 i_133534420(.A(n_56932), .B(n_29293), .C(n_2795), .D(n_28257)
		, .Z(n_349872808));
	notech_ao4 i_133434421(.A(n_2809), .B(n_28208), .C(n_56921), .D(nbus_11326
		[4]), .Z(n_349972809));
	notech_ao4 i_133234423(.A(n_56972), .B(n_27038), .C(n_56910), .D(n_27169
		), .Z(n_350172811));
	notech_and4 i_133734418(.A(n_350172811), .B(n_349972809), .C(n_349872808
		), .D(n_210171412), .Z(n_350372813));
	notech_ao4 i_132834427(.A(n_2802), .B(n_27234), .C(n_57168), .D(n_27203)
		, .Z(n_350572815));
	notech_ao4 i_132734428(.A(n_57298), .B(n_29063), .C(n_57177), .D(n_28147
		), .Z(n_350672816));
	notech_ao4 i_132534430(.A(n_2820), .B(\nbus_11276[20] ), .C(n_2783), .D(n_28179
		), .Z(n_350872818));
	notech_and4 i_133034425(.A(n_350872818), .B(n_350672816), .C(n_350572815
		), .D(n_209471405), .Z(n_351072820));
	notech_ao4 i_132234433(.A(n_2818), .B(n_28272), .C(n_2819), .D(n_28376),
		 .Z(n_351172821));
	notech_ao4 i_132134434(.A(n_2815), .B(n_28307), .C(n_2817), .D(n_28128),
		 .Z(n_351272822));
	notech_ao4 i_131934436(.A(n_2814), .B(n_28226), .C(n_2816), .D(n_28345),
		 .Z(n_351472824));
	notech_and4 i_132434431(.A(n_351472824), .B(n_351272822), .C(n_351172821
		), .D(n_208771398), .Z(n_351672826));
	notech_nand2 i_131834437(.A(n_55482), .B(n_56667), .Z(n_351872828));
	notech_ao4 i_131734438(.A(n_2799), .B(nbus_11279[3]), .C(n_55482), .D(n_339372703
		), .Z(n_351972829));
	notech_ao4 i_131334442(.A(n_56667), .B(n_188471195), .C(n_339372703), .D
		(n_351872828), .Z(n_352072830));
	notech_ao4 i_131234443(.A(n_340072710), .B(n_28390), .C(n_56609), .D(\nbus_11276[11] 
		), .Z(n_352172831));
	notech_ao4 i_131034445(.A(n_340572715), .B(n_27564), .C(n_340472714), .D
		(n_28118), .Z(n_352372833));
	notech_ao4 i_130934446(.A(n_55393), .B(nbus_11273[11]), .C(n_56640), .D(n_28086
		), .Z(n_352472834));
	notech_and4 i_131534440(.A(n_352472834), .B(n_352372833), .C(n_352172831
		), .D(n_352072830), .Z(n_352672836));
	notech_ao4 i_130634449(.A(n_56932), .B(n_29292), .C(n_2795), .D(n_28256)
		, .Z(n_352772837));
	notech_ao4 i_130534450(.A(n_2809), .B(n_28207), .C(n_56921), .D(nbus_11326
		[3]), .Z(n_352872838));
	notech_ao4 i_130334452(.A(n_56972), .B(n_27037), .C(n_56910), .D(n_27168
		), .Z(n_353072840));
	notech_and4 i_130834447(.A(n_353072840), .B(n_352872838), .C(n_352772837
		), .D(n_207071381), .Z(n_353272842));
	notech_ao4 i_129934456(.A(n_2802), .B(n_27233), .C(n_57168), .D(n_27202)
		, .Z(n_353472844));
	notech_ao4 i_129834457(.A(n_57298), .B(n_29043), .C(n_57177), .D(n_28146
		), .Z(n_353572845));
	notech_ao4 i_129634459(.A(n_2820), .B(\nbus_11276[19] ), .C(n_2783), .D(n_28178
		), .Z(n_353772847));
	notech_and4 i_130134454(.A(n_353772847), .B(n_353572845), .C(n_353472844
		), .D(n_206371374), .Z(n_353972849));
	notech_ao4 i_129334462(.A(n_2818), .B(n_28271), .C(n_2819), .D(n_28375),
		 .Z(n_354072850));
	notech_ao4 i_129234463(.A(n_2815), .B(n_28306), .C(n_2817), .D(n_28127),
		 .Z(n_354172851));
	notech_ao4 i_129034465(.A(n_2814), .B(n_28225), .C(n_2816), .D(n_28344),
		 .Z(n_354372853));
	notech_and4 i_129534460(.A(n_354372853), .B(n_354172851), .C(n_354072850
		), .D(n_205671367), .Z(n_354572855));
	notech_or4 i_128934466(.A(n_57399), .B(n_59944), .C(n_280472115), .D(opa
		[2]), .Z(n_354772857));
	notech_ao4 i_128834467(.A(n_2799), .B(nbus_11279[2]), .C(n_339372703), .D
		(n_326246826), .Z(n_354872858));
	notech_ao4 i_128434471(.A(n_56658), .B(n_188371194), .C(n_26282), .D(n_354772857
		), .Z(n_354972859));
	notech_ao4 i_128334472(.A(n_340072710), .B(n_28389), .C(n_56609), .D(\nbus_11276[10] 
		), .Z(n_355072860));
	notech_ao4 i_128134474(.A(n_340572715), .B(n_55299), .C(n_340472714), .D
		(n_28117), .Z(n_355288236));
	notech_ao4 i_128034475(.A(n_55393), .B(nbus_11273[10]), .C(n_56640), .D(n_28085
		), .Z(n_355372862));
	notech_and4 i_128634469(.A(n_355372862), .B(n_355288236), .C(n_355072860
		), .D(n_354972859), .Z(n_355588235));
	notech_ao4 i_127634478(.A(n_56932), .B(n_29291), .C(n_2795), .D(n_28255)
		, .Z(n_355672864));
	notech_ao4 i_127534479(.A(n_2809), .B(n_28206), .C(n_56921), .D(nbus_11326
		[2]), .Z(n_355772865));
	notech_ao4 i_127334481(.A(n_56972), .B(n_28141), .C(n_56910), .D(n_27167
		), .Z(n_355972867));
	notech_and4 i_127834476(.A(n_355972867), .B(n_355772865), .C(n_355672864
		), .D(n_203971350), .Z(n_356188234));
	notech_ao4 i_126934485(.A(n_2802), .B(n_27232), .C(n_57168), .D(n_27201)
		, .Z(n_356388232));
	notech_ao4 i_126834486(.A(n_57298), .B(n_29050), .C(n_57177), .D(n_28145
		), .Z(n_356488231));
	notech_ao4 i_126634488(.A(n_2820), .B(\nbus_11276[18] ), .C(n_2783), .D(n_28176
		), .Z(n_356688229));
	notech_and4 i_127134483(.A(n_356688229), .B(n_356488231), .C(n_356388232
		), .D(n_203271343), .Z(n_356888227));
	notech_ao4 i_126234491(.A(n_2818), .B(n_28270), .C(n_2819), .D(n_28374),
		 .Z(n_356988226));
	notech_ao4 i_126134492(.A(n_2815), .B(n_28305), .C(n_2817), .D(n_28126),
		 .Z(n_357088225));
	notech_ao4 i_125934494(.A(n_2814), .B(n_28224), .C(n_2816), .D(n_28343),
		 .Z(n_357288223));
	notech_and4 i_126434489(.A(n_357288223), .B(n_357088225), .C(n_356988226
		), .D(n_202571336), .Z(n_357488221));
	notech_ao4 i_125534498(.A(n_56609), .B(\nbus_11276[9] ), .C(n_188171192)
		, .D(n_56649), .Z(n_357688219));
	notech_ao4 i_125434499(.A(n_340472714), .B(n_28116), .C(n_340072710), .D
		(n_28388), .Z(n_357788218));
	notech_ao4 i_125234501(.A(n_339372703), .B(n_26309), .C(n_340572715), .D
		(n_55331), .Z(n_357988216));
	notech_ao4 i_125134502(.A(n_55393), .B(nbus_11273[9]), .C(n_56640), .D(n_28084
		), .Z(n_358088215));
	notech_and4 i_125734496(.A(n_358088215), .B(n_357988216), .C(n_357788218
		), .D(n_357688219), .Z(n_358288213));
	notech_ao4 i_124734505(.A(n_56921), .B(nbus_11326[1]), .C(n_2795), .D(n_28254
		), .Z(n_358388212));
	notech_ao4 i_124634506(.A(n_2809), .B(n_28205), .C(n_56932), .D(n_29290)
		, .Z(n_358488211));
	notech_ao4 i_124434508(.A(n_56972), .B(n_27036), .C(n_56910), .D(n_27166
		), .Z(n_358688209));
	notech_and4 i_125034503(.A(n_358688209), .B(n_358488211), .C(n_358388212
		), .D(n_201071321), .Z(n_358888207));
	notech_ao4 i_124034512(.A(n_2802), .B(n_27231), .C(n_57168), .D(n_27200)
		, .Z(n_359088205));
	notech_ao4 i_123934513(.A(n_57298), .B(n_29049), .C(n_57177), .D(n_28144
		), .Z(n_359188204));
	notech_ao4 i_123734515(.A(n_2820), .B(\nbus_11276[17] ), .C(n_2783), .D(n_28175
		), .Z(n_359388202));
	notech_and4 i_124234510(.A(n_359388202), .B(n_359188204), .C(n_359088205
		), .D(n_200371314), .Z(n_359588200));
	notech_ao4 i_123434518(.A(n_2818), .B(n_28269), .C(n_2819), .D(n_28373),
		 .Z(n_359688199));
	notech_ao4 i_123334519(.A(n_2815), .B(n_28304), .C(n_2817), .D(n_28125),
		 .Z(n_359788198));
	notech_ao4 i_123134521(.A(n_2814), .B(n_28223), .C(n_2816), .D(n_28342),
		 .Z(n_359988196));
	notech_and4 i_123634516(.A(n_359988196), .B(n_359788198), .C(n_359688199
		), .D(n_199671307), .Z(n_360188194));
	notech_ao4 i_122634526(.A(n_56609), .B(\nbus_11276[8] ), .C(nbus_11273[0
		]), .D(n_188071191), .Z(n_360488191));
	notech_ao4 i_122534527(.A(n_340472714), .B(n_28115), .C(n_340072710), .D
		(n_28387), .Z(n_360588190));
	notech_ao4 i_122334529(.A(n_56640), .B(n_28083), .C(n_340572715), .D(n_27561
		), .Z(n_360788188));
	notech_and4 i_122834524(.A(n_360788188), .B(n_360588190), .C(n_360488191
		), .D(n_198771298), .Z(n_360988186));
	notech_ao4 i_122034532(.A(n_56932), .B(n_29289), .C(n_2795), .D(n_28253)
		, .Z(n_361088185));
	notech_ao4 i_121934533(.A(n_2809), .B(n_28204), .C(n_56921), .D(nbus_11326
		[0]), .Z(n_361188184));
	notech_ao4 i_121734535(.A(n_56972), .B(n_28140), .C(n_56910), .D(n_27165
		), .Z(n_361388182));
	notech_and4 i_122234530(.A(n_361388182), .B(n_361188184), .C(n_361088185
		), .D(n_198071291), .Z(n_361588180));
	notech_ao4 i_121334539(.A(n_2802), .B(n_27230), .C(n_57168), .D(n_27199)
		, .Z(n_361788178));
	notech_ao4 i_121234540(.A(n_57298), .B(n_28986), .C(n_57177), .D(n_28143
		), .Z(n_361888177));
	notech_ao4 i_121034542(.A(n_2820), .B(\nbus_11276[16] ), .C(n_2783), .D(n_28174
		), .Z(n_362088175));
	notech_and4 i_121534537(.A(n_362088175), .B(n_361888177), .C(n_361788178
		), .D(n_197371284), .Z(n_362288173));
	notech_ao4 i_120734545(.A(n_2818), .B(n_28268), .C(n_2819), .D(n_28372),
		 .Z(n_362388172));
	notech_ao4 i_120634546(.A(n_2815), .B(n_28303), .C(n_2817), .D(n_28124),
		 .Z(n_362488171));
	notech_ao4 i_120434548(.A(n_2814), .B(n_28222), .C(n_2816), .D(n_28341),
		 .Z(n_362688169));
	notech_and4 i_120934543(.A(n_362688169), .B(n_362488171), .C(n_362388172
		), .D(n_196671277), .Z(n_362888167));
	notech_and4 i_64932892(.A(n_364588150), .B(n_363488161), .C(n_363388162)
		, .D(n_363588160), .Z(n_363088165));
	notech_or4 i_49132468(.A(n_60780), .B(n_60731), .C(n_1970), .D(n_29087),
		 .Z(n_363388162));
	notech_or2 i_49532467(.A(n_2177), .B(n_356476400), .Z(n_363488161));
	notech_or2 i_49632466(.A(n_2333), .B(nbus_11273[15]), .Z(n_363588160));
	notech_or2 i_27352(.A(n_57293), .B(n_55859), .Z(n_363688159));
	notech_or4 i_54932436(.A(n_60782), .B(n_60731), .C(n_57374), .D(n_26599)
		, .Z(n_363788158));
	notech_or4 i_55032435(.A(n_60782), .B(n_60731), .C(n_1900), .D(n_56112),
		 .Z(n_363888157));
	notech_ao4 i_122431861(.A(n_254834174), .B(\nbus_11276[15] ), .C(n_59854
		), .D(n_27534), .Z(n_364588150));
	notech_and4 i_52596(.A(n_280172112), .B(n_208741718), .C(n_55645), .D(n_54811
		), .Z(\nbus_11339[0] ));
	notech_nand2 i_104565718(.A(pipe_mul[1]), .B(n_26886), .Z(n_55324));
	notech_ao4 i_162640660(.A(n_354488264), .B(\nbus_11276[21] ), .C(n_323462238
		), .D(n_29172), .Z(n_319162195));
	notech_or2 i_26865706(.A(n_55484), .B(n_125270571), .Z(nbus_11313[16])
		);
	notech_and4 i_163340653(.A(n_318862192), .B(n_318662190), .C(n_298761991
		), .D(n_299061994), .Z(n_319062194));
	notech_nand3 i_21757(.A(n_2771), .B(n_26621), .C(n_26607), .Z(n_208741718
		));
	notech_ao4 i_162940657(.A(n_5538), .B(n_27588), .C(n_59188), .D(n_26764)
		, .Z(n_318862192));
	notech_nand3 i_1716218(.A(n_127070589), .B(n_126970588), .C(n_126870587)
		, .Z(n_21202));
	notech_nor2 i_30265681(.A(n_312283097), .B(n_125170570), .Z(n_207841709)
		);
	notech_ao4 i_76465676(.A(n_59865), .B(n_274788710), .C(n_207841709), .D(n_55878
		), .Z(n_207341704));
	notech_or4 i_163635711(.A(n_60782), .B(n_60731), .C(n_195571266), .D(n_60598
		), .Z(n_54811));
	notech_or4 i_70535740(.A(n_60782), .B(n_60729), .C(n_195671267), .D(n_60596
		), .Z(n_55645));
	notech_and4 i_721042(.A(n_128870607), .B(n_129070609), .C(n_129470613), 
		.D(n_128770606), .Z(n_13851));
	notech_and4 i_521040(.A(n_129570614), .B(n_129770616), .C(n_130170620), 
		.D(n_127970598), .Z(n_13839));
	notech_and4 i_189760640(.A(n_56060), .B(n_1021), .C(n_55995), .D(n_56001
		), .Z(n_54595));
	notech_ao3 i_193260632(.A(n_55064), .B(n_54435), .C(n_138370702), .Z(n_54566
		));
	notech_and3 i_193560631(.A(n_55062), .B(n_138270701), .C(n_54458), .Z(n_54564
		));
	notech_ao4 i_163140655(.A(n_310518882), .B(n_323762241), .C(n_312662130)
		, .D(n_3288), .Z(n_318662190));
	notech_and4 i_163840648(.A(n_318362187), .B(n_318162185), .C(n_299361997
		), .D(n_299662000), .Z(n_318562189));
	notech_ao4 i_163440652(.A(n_262336778), .B(n_29173), .C(n_353488274), .D
		(nbus_11326[22]), .Z(n_318362187));
	notech_or4 i_1020949(.A(n_26252), .B(n_134270661), .C(n_134970668), .D(n_26253
		), .Z(n_9033));
	notech_or4 i_920948(.A(n_145974327), .B(n_132870647), .C(n_135370672), .D
		(n_26254), .Z(n_9027));
	notech_and4 i_920980(.A(n_135770676), .B(n_135970678), .C(n_136470683), 
		.D(n_132770646), .Z(n_16747));
	notech_nand3 i_1021045(.A(n_136770686), .B(n_136670685), .C(n_137170690)
		, .Z(n_13869));
	notech_or4 i_921044(.A(n_145974327), .B(n_130470623), .C(n_137570694), .D
		(n_26255), .Z(n_13863));
	notech_or4 i_28343(.A(n_56465), .B(n_355988238), .C(n_29010), .D(n_26306
		), .Z(n_364788148));
	notech_and2 i_59257985(.A(n_181471126), .B(n_138570704), .Z(n_55757));
	notech_nao3 i_181357953(.A(n_55073), .B(n_54453), .C(n_45383), .Z(n_54665
		));
	notech_and3 i_181457952(.A(n_45384), .B(n_55072), .C(n_54454), .Z(n_54664
		));
	notech_or4 i_28992(.A(n_56492), .B(n_56478), .C(n_2349), .D(n_54069), .Z
		(n_254734173));
	notech_and4 i_251857932(.A(n_56061), .B(n_1022), .C(n_55995), .D(n_252434150
		), .Z(n_54070));
	notech_ao4 i_163640650(.A(n_354488264), .B(\nbus_11276[22] ), .C(n_323462238
		), .D(n_29174), .Z(n_318162185));
	notech_and4 i_164340643(.A(n_317862182), .B(n_317662180), .C(n_299962003
		), .D(n_300262006), .Z(n_318062184));
	notech_or4 i_206557921(.A(n_1916), .B(n_1023), .C(n_56001), .D(n_60532),
		 .Z(n_54458));
	notech_or2 i_209357920(.A(n_54527), .B(n_56001), .Z(n_54435));
	notech_and4 i_821043(.A(n_139370712), .B(n_140370722), .C(n_140570724), 
		.D(n_140970728), .Z(n_13857));
	notech_or4 i_191457850(.A(n_56487), .B(n_56478), .C(n_1976), .D(n_54070)
		, .Z(n_247334099));
	notech_or4 i_192057849(.A(n_56487), .B(n_56478), .C(n_56449), .D(n_56001
		), .Z(n_247234098));
	notech_and4 i_1620955(.A(n_363088165), .B(n_154570864), .C(n_152470843),
		 .D(n_154470863), .Z(n_9069));
	notech_or4 i_1420953(.A(n_188774755), .B(n_151670835), .C(n_155170870), 
		.D(n_26256), .Z(n_9057));
	notech_or4 i_1320952(.A(n_189974767), .B(n_150870827), .C(n_155870877), 
		.D(n_26257), .Z(n_9051));
	notech_or4 i_1220951(.A(n_239168196), .B(n_150070819), .C(n_156570884), 
		.D(n_26258), .Z(n_9045));
	notech_and4 i_1620987(.A(n_149970818), .B(n_156970888), .C(n_157170890),
		 .D(n_157670895), .Z(n_16789));
	notech_or4 i_1420985(.A(n_149070809), .B(n_158470903), .C(n_26259), .D(n_26260
		), .Z(n_16777));
	notech_or4 i_1320984(.A(n_148170800), .B(n_159270911), .C(n_26262), .D(n_26263
		), .Z(n_16771));
	notech_or4 i_1220983(.A(n_147270791), .B(n_160070919), .C(n_26265), .D(n_26266
		), .Z(n_16765));
	notech_and4 i_1120982(.A(n_160270921), .B(n_160470923), .C(n_146370782),
		 .D(n_160870927), .Z(n_16759));
	notech_and4 i_1621051(.A(n_363088165), .B(n_161370932), .C(n_144870767),
		 .D(n_161270931), .Z(n_13905));
	notech_or4 i_1421049(.A(n_188774755), .B(n_144070759), .C(n_161970938), 
		.D(n_26269), .Z(n_13893));
	notech_or4 i_1321048(.A(n_189974767), .B(n_143270751), .C(n_162670945), 
		.D(n_26270), .Z(n_13887));
	notech_or4 i_1221047(.A(n_239168196), .B(n_142470743), .C(n_163370952), 
		.D(n_26271), .Z(n_13881));
	notech_nand3 i_1121046(.A(n_163970958), .B(n_163870957), .C(n_164370962)
		, .Z(n_13875));
	notech_ao4 i_129555295(.A(n_54121), .B(n_27575), .C(n_322131608), .D(n_55859
		), .Z(n_319431581));
	notech_ao4 i_163940647(.A(n_5538), .B(n_27589), .C(n_59197), .D(n_26765)
		, .Z(n_317862182));
	notech_and3 i_181757950(.A(n_55062), .B(n_138270701), .C(n_54441), .Z(n_54563
		));
	notech_ao3 i_181557951(.A(n_55064), .B(n_54459), .C(n_138370702), .Z(n_54565
		));
	notech_nand2 i_59757982(.A(n_55720), .B(n_138470703), .Z(n_55752));
	notech_ao4 i_164140645(.A(n_310418881), .B(n_323762241), .C(n_305565372)
		, .D(n_3288), .Z(n_317662180));
	notech_and4 i_192740365(.A(n_317362177), .B(n_317162175), .C(n_300562009
		), .D(n_300862012), .Z(n_317562179));
	notech_or4 i_2921064(.A(n_313168930), .B(n_172371042), .C(n_174371062), 
		.D(n_26272), .Z(n_13983));
	notech_or4 i_2821063(.A(n_264975488), .B(n_171571034), .C(n_175071069), 
		.D(n_26273), .Z(n_13977));
	notech_or4 i_2721062(.A(n_265975498), .B(n_170771026), .C(n_175771076), 
		.D(n_26274), .Z(n_13971));
	notech_or4 i_2621061(.A(n_173971058), .B(n_169971018), .C(n_176471083), 
		.D(n_26275), .Z(n_13965));
	notech_or4 i_2421059(.A(n_267675515), .B(n_169171010), .C(n_177171090), 
		.D(n_26276), .Z(n_13953));
	notech_or2 i_43345379(.A(n_56376), .B(n_27593), .Z(n_307521962));
	notech_ao4 i_192340369(.A(n_55567), .B(nbus_11273[20]), .C(n_55568), .D(\nbus_11276[20] 
		), .Z(n_317362177));
	notech_nand2 i_46231(.A(n_300586325), .B(n_196071271), .Z(n_7432));
	notech_and4 i_52597(.A(n_55645), .B(n_208741718), .C(n_279872109), .D(n_280172112
		), .Z(\nbus_11339[8] ));
	notech_xor2 i_126535761(.A(opa[1]), .B(opa[0]), .Z(n_55114));
	notech_ao4 i_192540367(.A(n_55492), .B(n_27540), .C(n_58922), .D(n_29175
		), .Z(n_317162175));
	notech_ao3 i_78135712(.A(n_26652), .B(n_59865), .C(n_274988708), .Z(n_55569
		));
	notech_and4 i_151435708(.A(n_57380), .B(n_57423), .C(n_57424), .D(n_280072111
		), .Z(n_54914));
	notech_nand2 i_6435(.A(n_287072181), .B(n_286572176), .Z(n_7418));
	notech_nand3 i_3217418(.A(n_289472205), .B(n_289072201), .C(n_288572196)
		, .Z(n_17382));
	notech_nand3 i_3117417(.A(n_291472225), .B(n_291072221), .C(n_290572216)
		, .Z(n_17376));
	notech_nand3 i_3017416(.A(n_293472245), .B(n_293072241), .C(n_292572236)
		, .Z(n_17370));
	notech_nand3 i_2917415(.A(n_295472265), .B(n_295072261), .C(n_294572256)
		, .Z(n_17364));
	notech_nand3 i_2817414(.A(n_297472285), .B(n_297072281), .C(n_296572276)
		, .Z(n_17358));
	notech_nand3 i_2717413(.A(n_299472305), .B(n_299072301), .C(n_298572296)
		, .Z(n_17352));
	notech_nand3 i_2617412(.A(n_301472325), .B(n_301072321), .C(n_300572316)
		, .Z(n_17346));
	notech_nand3 i_2517411(.A(n_303472345), .B(n_303072341), .C(n_302572336)
		, .Z(n_17340));
	notech_nand3 i_2417410(.A(n_304072351), .B(n_305572366), .C(n_304472355)
		, .Z(n_17334));
	notech_nand3 i_2317409(.A(n_307472385), .B(n_307072381), .C(n_306572376)
		, .Z(n_17328));
	notech_nand3 i_2217408(.A(n_309472405), .B(n_309072401), .C(n_308572396)
		, .Z(n_17322));
	notech_nand3 i_2117407(.A(n_311472425), .B(n_311072421), .C(n_310572416)
		, .Z(n_17316));
	notech_nand3 i_2017406(.A(n_313472445), .B(n_313072441), .C(n_312572436)
		, .Z(n_17310));
	notech_nand3 i_1917405(.A(n_315472465), .B(n_315072461), .C(n_314572456)
		, .Z(n_17304));
	notech_nand3 i_1817404(.A(n_316072471), .B(n_317572486), .C(n_316472475)
		, .Z(n_17298));
	notech_nand3 i_1717403(.A(n_319472505), .B(n_319072501), .C(n_318572496)
		, .Z(n_17292));
	notech_and4 i_1617402(.A(n_322272533), .B(n_321672527), .C(n_320872519),
		 .D(n_320272513), .Z(n_17286));
	notech_and4 i_1517401(.A(n_325072561), .B(n_324472555), .C(n_323672547),
		 .D(n_323072541), .Z(n_17280));
	notech_and4 i_1317399(.A(n_327872589), .B(n_327272583), .C(n_326472575),
		 .D(n_325872569), .Z(n_17268));
	notech_and4 i_1217398(.A(n_330772617), .B(n_330172611), .C(n_329372603),
		 .D(n_328672597), .Z(n_17262));
	notech_and4 i_1117397(.A(n_333572645), .B(n_332972639), .C(n_332172631),
		 .D(n_331572625), .Z(n_17256));
	notech_and4 i_1017396(.A(n_336372673), .B(n_335772667), .C(n_334972659),
		 .D(n_334372653), .Z(n_17250));
	notech_and4 i_917395(.A(n_339172701), .B(n_338572695), .C(n_337772687), 
		.D(n_337172681), .Z(n_17244));
	notech_and4 i_817394(.A(n_342972739), .B(n_342372733), .C(n_341572725), 
		.D(n_340972719), .Z(n_17238));
	notech_and4 i_717393(.A(n_345872768), .B(n_345272762), .C(n_344572755), 
		.D(n_343972749), .Z(n_17232));
	notech_and4 i_617392(.A(n_348772797), .B(n_348172791), .C(n_347472784), 
		.D(n_346872778), .Z(n_17226));
	notech_and4 i_517391(.A(n_351672826), .B(n_351072820), .C(n_350372813), 
		.D(n_349772807), .Z(n_17220));
	notech_and4 i_417390(.A(n_354572855), .B(n_353972849), .C(n_353272842), 
		.D(n_352672836), .Z(n_17214));
	notech_and4 i_317389(.A(n_357488221), .B(n_356888227), .C(n_356188234), 
		.D(n_355588235), .Z(n_17208));
	notech_and4 i_217388(.A(n_360188194), .B(n_359588200), .C(n_358888207), 
		.D(n_358288213), .Z(n_17202));
	notech_and4 i_117387(.A(n_362888167), .B(n_362288173), .C(n_361588180), 
		.D(n_360988186), .Z(n_17196));
	notech_or4 i_2735669(.A(n_2550), .B(n_1844), .C(n_60563), .D(n_59380), .Z
		(n_327246816));
	notech_and4 i_31533120(.A(n_56057), .B(n_55920), .C(n_363888157), .D(n_363788158
		), .Z(n_56034));
	notech_and2 i_2467(.A(n_56376), .B(n_36952), .Z(n_54121));
	notech_and4 i_193240360(.A(n_316862172), .B(n_316662170), .C(n_301162015
		), .D(n_301462018), .Z(n_317062174));
	notech_ao4 i_192840364(.A(n_59197), .B(n_26786), .C(n_26435), .D(n_29176
		), .Z(n_316862172));
	notech_ao4 i_193040362(.A(n_55811), .B(n_310618883), .C(n_2211), .D(n_315162155
		), .Z(n_316662170));
	notech_ao4 i_193340359(.A(n_54439), .B(n_29177), .C(n_56151), .D(n_27626
		), .Z(n_316362167));
	notech_ao4 i_193440358(.A(n_56126), .B(n_27666), .C(n_56097), .D(n_27703
		), .Z(n_316262166));
	notech_and2 i_193840354(.A(n_316062164), .B(n_315962163), .Z(n_316162165
		));
	notech_ao4 i_193640356(.A(n_54535), .B(n_27390), .C(n_55864), .D(n_27735
		), .Z(n_316062164));
	notech_ao4 i_193740355(.A(n_55898), .B(n_27772), .C(n_55940), .D(n_27806
		), .Z(n_315962163));
	notech_and4 i_194640346(.A(n_315662160), .B(n_315562159), .C(n_315362157
		), .D(n_315262156), .Z(n_315862162));
	notech_ao4 i_194040352(.A(n_55879), .B(n_27838), .C(n_56068), .D(n_27872
		), .Z(n_315662160));
	notech_ao4 i_194140351(.A(n_56035), .B(n_27907), .C(n_56009), .D(n_27940
		), .Z(n_315562159));
	notech_ao4 i_194340349(.A(n_55998), .B(n_27973), .C(n_55872), .D(n_28007
		), .Z(n_315362157));
	notech_ao4 i_194440348(.A(n_55873), .B(n_29178), .C(n_55878), .D(n_28039
		), .Z(n_315262156));
	notech_nand2 i_2142256(.A(opc_10[20]), .B(n_62399), .Z(n_315162155));
	notech_and4 i_195140341(.A(n_314862152), .B(n_314662150), .C(n_303362037
		), .D(n_303662040), .Z(n_315062154));
	notech_ao4 i_194740345(.A(n_55567), .B(nbus_11273[21]), .C(n_55568), .D(\nbus_11276[21] 
		), .Z(n_314862152));
	notech_ao4 i_194940343(.A(n_55492), .B(n_27541), .C(n_58922), .D(n_29179
		), .Z(n_314662150));
	notech_and4 i_195640336(.A(n_314362147), .B(n_314162145), .C(n_303962043
		), .D(n_304262046), .Z(n_314562149));
	notech_ao4 i_195240340(.A(n_59195), .B(n_26787), .C(n_26435), .D(n_29180
		), .Z(n_314362147));
	notech_ao4 i_195440338(.A(n_55811), .B(n_310518882), .C(n_2211), .D(n_312662130
		), .Z(n_314162145));
	notech_ao4 i_195740335(.A(n_54439), .B(n_29181), .C(n_56151), .D(n_27627
		), .Z(n_313862142));
	notech_ao4 i_195840334(.A(n_56126), .B(n_27667), .C(n_56097), .D(n_27704
		), .Z(n_313762141));
	notech_and2 i_196240330(.A(n_313562139), .B(n_313462138), .Z(n_313662140
		));
	notech_ao4 i_196040332(.A(n_54535), .B(n_27391), .C(n_55864), .D(n_27736
		), .Z(n_313562139));
	notech_ao4 i_196140331(.A(n_55898), .B(n_27773), .C(n_55940), .D(n_27807
		), .Z(n_313462138));
	notech_and4 i_197040322(.A(n_313162135), .B(n_313062134), .C(n_312862132
		), .D(n_312762131), .Z(n_313362137));
	notech_ao4 i_196440328(.A(n_55866), .B(n_27839), .C(n_56068), .D(n_27873
		), .Z(n_313162135));
	notech_ao4 i_196540327(.A(n_56035), .B(n_27908), .C(n_56009), .D(n_27942
		), .Z(n_313062134));
	notech_ao4 i_196740325(.A(n_55998), .B(n_27974), .C(n_55872), .D(n_28008
		), .Z(n_312862132));
	notech_ao4 i_196840324(.A(n_55873), .B(n_29182), .C(n_55878), .D(n_28040
		), .Z(n_312762131));
	notech_nand2 i_2242255(.A(opc_10[21]), .B(n_62399), .Z(n_312662130));
	notech_or2 i_158242272(.A(n_294061944), .B(n_56240), .Z(n_312462128));
	notech_ao4 i_200440288(.A(n_2263), .B(n_26381), .C(n_294061944), .D(n_26314
		), .Z(n_312362127));
	notech_ao4 i_202440268(.A(n_29182), .B(n_2261), .C(n_56240), .D(n_27736)
		, .Z(n_312062124));
	notech_ao4 i_202540267(.A(n_2262), .B(n_27807), .C(n_27839), .D(n_197114365
		), .Z(n_311962123));
	notech_and2 i_202940263(.A(n_311762121), .B(n_311662120), .Z(n_311862122
		));
	notech_ao4 i_202740265(.A(n_28008), .B(n_56178), .C(n_57343), .D(n_27773
		), .Z(n_311762121));
	notech_ao4 i_202840264(.A(n_56414), .B(n_27974), .C(n_56310), .D(n_27627
		), .Z(n_311662120));
	notech_and4 i_203740255(.A(n_311362117), .B(n_311262116), .C(n_311062114
		), .D(n_310962113), .Z(n_311562119));
	notech_ao4 i_203140261(.A(n_27942), .B(n_56182), .C(n_56183), .D(n_29181
		), .Z(n_311362117));
	notech_ao4 i_203240260(.A(n_60484), .B(n_27908), .C(n_56290), .D(n_27667
		), .Z(n_311262116));
	notech_ao4 i_203440258(.A(n_56186), .B(n_27873), .C(n_56270), .D(n_27704
		), .Z(n_311062114));
	notech_ao4 i_203540257(.A(n_59224), .B(n_28040), .C(n_57373), .D(n_27391
		), .Z(n_310962113));
	notech_ao4 i_204040252(.A(n_29178), .B(n_2261), .C(n_56240), .D(n_27735)
		, .Z(n_310662110));
	notech_ao4 i_204140251(.A(n_2262), .B(n_27806), .C(n_27838), .D(n_197114365
		), .Z(n_310562109));
	notech_and2 i_204540247(.A(n_310362107), .B(n_310262106), .Z(n_310462108
		));
	notech_ao4 i_204340249(.A(n_28007), .B(n_56178), .C(n_57343), .D(n_27772
		), .Z(n_310362107));
	notech_ao4 i_204440248(.A(n_56414), .B(n_27973), .C(n_56310), .D(n_27626
		), .Z(n_310262106));
	notech_and4 i_205340239(.A(n_309962103), .B(n_309862102), .C(n_309662100
		), .D(n_309562099), .Z(n_310162105));
	notech_ao4 i_204740245(.A(n_27940), .B(n_56182), .C(n_56183), .D(n_29177
		), .Z(n_309962103));
	notech_ao4 i_204840244(.A(n_60484), .B(n_27907), .C(n_56290), .D(n_27666
		), .Z(n_309862102));
	notech_ao4 i_205040242(.A(n_56186), .B(n_27872), .C(n_56270), .D(n_27703
		), .Z(n_309662100));
	notech_ao4 i_205140241(.A(n_59224), .B(n_28039), .C(n_57373), .D(n_27390
		), .Z(n_309562099));
	notech_or4 i_30894(.A(n_56465), .B(n_264436799), .C(n_56469), .D(n_60512
		), .Z(n_306062064));
	notech_or2 i_92741340(.A(n_55587), .B(n_311018887), .Z(n_304262046));
	notech_or2 i_93041337(.A(n_55842), .B(n_27588), .Z(n_303962043));
	notech_or2 i_93341334(.A(n_55597), .B(n_29172), .Z(n_303662040));
	notech_or2 i_93641331(.A(n_2212), .B(nbus_11326[21]), .Z(n_303362037));
	notech_or2 i_89641368(.A(n_55587), .B(n_311118888), .Z(n_301462018));
	notech_or2 i_89941365(.A(n_55842), .B(n_27586), .Z(n_301162015));
	notech_or2 i_90241362(.A(n_55597), .B(n_29169), .Z(n_300862012));
	notech_or2 i_90641359(.A(n_2212), .B(nbus_11326[20]), .Z(n_300562009));
	notech_nand2 i_55341696(.A(n_26415), .B(n_310918886), .Z(n_300262006));
	notech_nand3 i_55641693(.A(n_59197), .B(n_59944), .C(read_data[22]), .Z(n_299962003
		));
	notech_or2 i_55941690(.A(n_353988269), .B(nbus_11273[22]), .Z(n_299662000
		));
	notech_nao3 i_56241687(.A(n_2458), .B(n_29091), .C(n_232761396), .Z(n_299361997
		));
	notech_or2 i_54041708(.A(n_311018887), .B(n_323662240), .Z(n_299061994)
		);
	notech_nand3 i_54341705(.A(n_59197), .B(n_59944), .C(read_data[21]), .Z(n_298761991
		));
	notech_or2 i_54641702(.A(n_353988269), .B(nbus_11273[21]), .Z(n_298461988
		));
	notech_nao3 i_55041699(.A(n_2456), .B(n_29091), .C(n_232761396), .Z(n_298161985
		));
	notech_or2 i_52841720(.A(n_311118888), .B(n_323662240), .Z(n_297861982)
		);
	notech_nand3 i_53141717(.A(n_59197), .B(n_59940), .C(read_data[20]), .Z(n_297561979
		));
	notech_or2 i_53441714(.A(n_353988269), .B(nbus_11273[20]), .Z(n_297261976
		));
	notech_nao3 i_53741711(.A(n_2454), .B(n_29091), .C(n_232761396), .Z(n_296961973
		));
	notech_or2 i_51641732(.A(n_311218889), .B(n_323662240), .Z(n_296661970)
		);
	notech_nand3 i_51941729(.A(n_59195), .B(n_59940), .C(read_data[19]), .Z(n_296361967
		));
	notech_or2 i_52241726(.A(n_353988269), .B(nbus_11273[19]), .Z(n_296061964
		));
	notech_nao3 i_52541723(.A(n_2452), .B(n_29091), .C(n_232761396), .Z(n_295761961
		));
	notech_or2 i_50441744(.A(n_311318890), .B(n_323662240), .Z(n_295461958)
		);
	notech_nand3 i_50741741(.A(n_59195), .B(n_59940), .C(read_data[18]), .Z(n_295161955
		));
	notech_or2 i_51041738(.A(n_353988269), .B(nbus_11273[18]), .Z(n_294861952
		));
	notech_nao3 i_51341735(.A(n_2450), .B(n_29091), .C(n_232761396), .Z(n_294561949
		));
	notech_nao3 i_23842253(.A(n_56465), .B(n_29010), .C(n_264436799), .Z(n_294261946
		));
	notech_ao4 i_84342244(.A(n_59380), .B(n_62415), .C(n_2264), .D(n_26381),
		 .Z(n_294061944));
	notech_or2 i_99941271(.A(n_55859), .B(n_26513), .Z(n_293761941));
	notech_ao4 i_37842252(.A(n_2044), .B(n_56112), .C(n_56063), .D(n_26513),
		 .Z(n_293161935));
	notech_and2 i_149042275(.A(n_312362127), .B(n_56260), .Z(n_293061934));
	notech_and4 i_161543816(.A(n_292761931), .B(n_292561929), .C(n_272061748
		), .D(n_272361751), .Z(n_292961933));
	notech_ao4 i_161143820(.A(n_262336778), .B(n_29151), .C(n_353488274), .D
		(nbus_11326[23]), .Z(n_292761931));
	notech_ao4 i_161343818(.A(n_354488264), .B(\nbus_11276[23] ), .C(n_323462238
		), .D(n_29152), .Z(n_292561929));
	notech_and4 i_162043811(.A(n_292261926), .B(n_292061924), .C(n_272661754
		), .D(n_272961757), .Z(n_292461928));
	notech_ao4 i_161643815(.A(n_5538), .B(n_27590), .C(n_59195), .D(n_26766)
		, .Z(n_292261926));
	notech_ao4 i_161843813(.A(n_308521972), .B(n_323762241), .C(n_270765024)
		, .D(n_3288), .Z(n_292061924));
	notech_and4 i_164543786(.A(n_291761921), .B(n_291561919), .C(n_273261760
		), .D(n_273561763), .Z(n_291961923));
	notech_ao4 i_164143790(.A(n_262336778), .B(n_29153), .C(n_353488274), .D
		(nbus_11326[27]), .Z(n_291761921));
	notech_ao4 i_164343788(.A(n_354488264), .B(\nbus_11276[27] ), .C(n_29154
		), .D(n_354888260), .Z(n_291561919));
	notech_and4 i_165043781(.A(n_291261916), .B(n_291061914), .C(n_273861766
		), .D(n_274161769), .Z(n_291461918));
	notech_ao4 i_164643785(.A(n_5538), .B(n_27595), .C(n_59195), .D(n_26770)
		, .Z(n_291261916));
	notech_ao4 i_164843783(.A(n_354388265), .B(n_308221969), .C(n_286061878)
		, .D(n_354988259), .Z(n_291061914));
	notech_and4 i_193643497(.A(n_290761911), .B(n_290561909), .C(n_274461772
		), .D(n_274761775), .Z(n_290961913));
	notech_ao4 i_193243501(.A(n_55567), .B(nbus_11273[26]), .C(n_55568), .D(\nbus_11276[26] 
		), .Z(n_290761911));
	notech_ao4 i_193443499(.A(n_55492), .B(n_27549), .C(n_58922), .D(n_29155
		), .Z(n_290561909));
	notech_and4 i_194143492(.A(n_290261906), .B(n_290061904), .C(n_275061778
		), .D(n_275361781), .Z(n_290461908));
	notech_ao4 i_193743496(.A(n_59195), .B(n_26793), .C(n_26435), .D(n_29157
		), .Z(n_290261906));
	notech_ao4 i_193943494(.A(n_55811), .B(n_308321970), .C(n_2211), .D(n_288561889
		), .Z(n_290061904));
	notech_ao4 i_194243491(.A(n_54439), .B(n_29158), .C(n_56151), .D(n_27632
		), .Z(n_289761901));
	notech_ao4 i_194343490(.A(n_56126), .B(n_27673), .C(n_56097), .D(n_27709
		), .Z(n_289661900));
	notech_and2 i_194743486(.A(n_289461898), .B(n_289361897), .Z(n_289561899
		));
	notech_ao4 i_194543488(.A(n_54535), .B(n_27396), .C(n_55864), .D(n_27741
		), .Z(n_289461898));
	notech_ao4 i_194643487(.A(n_55898), .B(n_27780), .C(n_55940), .D(n_27812
		), .Z(n_289361897));
	notech_and4 i_195543478(.A(n_289061894), .B(n_288961893), .C(n_288761891
		), .D(n_288661890), .Z(n_289261896));
	notech_ao4 i_194943484(.A(n_55866), .B(n_27844), .C(n_56068), .D(n_27879
		), .Z(n_289061894));
	notech_ao4 i_195043483(.A(n_56035), .B(n_27913), .C(n_56009), .D(n_27947
		), .Z(n_288961893));
	notech_ao4 i_195243481(.A(n_55998), .B(n_27979), .C(n_55872), .D(n_28013
		), .Z(n_288761891));
	notech_ao4 i_195343480(.A(n_55873), .B(n_29159), .C(n_55878), .D(n_28045
		), .Z(n_288661890));
	notech_nand2 i_2845383(.A(opc_10[26]), .B(n_62399), .Z(n_288561889));
	notech_and4 i_196043473(.A(n_288261886), .B(n_288061884), .C(n_277261800
		), .D(n_277561803), .Z(n_288461888));
	notech_ao4 i_195643477(.A(n_55567), .B(nbus_11273[27]), .C(n_55568), .D(\nbus_11276[27] 
		), .Z(n_288261886));
	notech_ao4 i_195843475(.A(n_55492), .B(n_27550), .C(n_58922), .D(n_29160
		), .Z(n_288061884));
	notech_and4 i_196543468(.A(n_2877), .B(n_2875), .C(n_277861806), .D(n_278161809
		), .Z(n_287961883));
	notech_ao4 i_196143472(.A(n_59195), .B(n_26794), .C(n_26435), .D(n_29161
		), .Z(n_2877));
	notech_ao4 i_196343470(.A(n_55811), .B(n_308221969), .C(n_2211), .D(n_286061878
		), .Z(n_2875));
	notech_ao4 i_196643467(.A(n_55873), .B(n_29162), .C(n_55864), .D(n_27742
		), .Z(n_2872));
	notech_ao4 i_196743466(.A(n_55866), .B(n_27845), .C(n_55872), .D(n_28014
		), .Z(n_2871));
	notech_and2 i_197143462(.A(n_2869), .B(n_2868), .Z(n_2870));
	notech_ao4 i_196943464(.A(n_55898), .B(n_27781), .C(n_55998), .D(n_27980
		), .Z(n_2869));
	notech_ao4 i_197043463(.A(n_56151), .B(n_27633), .C(n_56009), .D(n_27948
		), .Z(n_2868));
	notech_and4 i_197943454(.A(n_286561881), .B(n_2864), .C(n_286261879), .D
		(n_2861), .Z(n_2867));
	notech_ao4 i_197343460(.A(n_56386), .B(n_29163), .C(n_56035), .D(n_27914
		), .Z(n_286561881));
	notech_ao4 i_197443459(.A(n_56126), .B(n_27674), .C(n_56068), .D(n_27880
		), .Z(n_2864));
	notech_ao4 i_197643457(.A(n_56097), .B(n_27710), .C(n_55878), .D(n_28046
		), .Z(n_286261879));
	notech_ao4 i_197743456(.A(n_54535), .B(n_27397), .C(n_55940), .D(n_27813
		), .Z(n_2861));
	notech_nand2 i_2945382(.A(opc_10[27]), .B(n_62399), .Z(n_286061878));
	notech_ao4 i_204443389(.A(n_2261), .B(n_29162), .C(n_56240), .D(n_27742)
		, .Z(n_2857));
	notech_ao4 i_204543388(.A(n_2262), .B(n_27813), .C(n_27845), .D(n_197114365
		), .Z(n_2856));
	notech_and2 i_204943384(.A(n_2854), .B(n_285361876), .Z(n_2855));
	notech_ao4 i_204743386(.A(n_56178), .B(n_28014), .C(n_57343), .D(n_27781
		), .Z(n_2854));
	notech_ao4 i_204843385(.A(n_56415), .B(n_27980), .C(n_56310), .D(n_27633
		), .Z(n_285361876));
	notech_and4 i_205743376(.A(n_2850), .B(n_284961873), .C(n_284761871), .D
		(n_284661870), .Z(n_285261875));
	notech_ao4 i_205143382(.A(n_56182), .B(n_27948), .C(n_56183), .D(n_29163
		), .Z(n_2850));
	notech_ao4 i_205243381(.A(n_60484), .B(n_27914), .C(n_56290), .D(n_27674
		), .Z(n_284961873));
	notech_ao4 i_205443379(.A(n_56186), .B(n_27880), .C(n_56270), .D(n_27710
		), .Z(n_284761871));
	notech_ao4 i_205543378(.A(n_59224), .B(n_28046), .C(n_57373), .D(n_27397
		), .Z(n_284661870));
	notech_ao4 i_206043373(.A(n_29159), .B(n_2261), .C(n_56240), .D(n_27741)
		, .Z(n_284361868));
	notech_ao4 i_206143372(.A(n_2262), .B(n_27812), .C(n_27844), .D(n_197114365
		), .Z(n_284261867));
	notech_and2 i_206543368(.A(n_2840), .B(n_2839), .Z(n_2841));
	notech_ao4 i_206343370(.A(n_28013), .B(n_56178), .C(n_57343), .D(n_27780
		), .Z(n_2840));
	notech_ao4 i_206443369(.A(n_56415), .B(n_27979), .C(n_56310), .D(n_27632
		), .Z(n_2839));
	notech_and4 i_207343360(.A(n_283661864), .B(n_283561863), .C(n_283361861
		), .D(n_283261860), .Z(n_283861866));
	notech_ao4 i_206743366(.A(n_27947), .B(n_56182), .C(n_56183), .D(n_29158
		), .Z(n_283661864));
	notech_ao4 i_206843365(.A(n_60484), .B(n_27913), .C(n_56290), .D(n_27673
		), .Z(n_283561863));
	notech_ao4 i_207043363(.A(n_56186), .B(n_27879), .C(n_56270), .D(n_27709
		), .Z(n_283361861));
	notech_ao4 i_207143362(.A(n_59224), .B(n_28045), .C(n_57373), .D(n_27396
		), .Z(n_283261860));
	notech_and3 i_5445323(.A(n_55658), .B(n_135960441), .C(n_56005), .Z(n_279961827
		));
	notech_or2 i_96944434(.A(n_55587), .B(n_308621973), .Z(n_278161809));
	notech_or2 i_97244431(.A(n_55842), .B(n_27595), .Z(n_277861806));
	notech_or2 i_97544428(.A(n_55597), .B(n_29154), .Z(n_277561803));
	notech_or2 i_97844425(.A(n_2212), .B(nbus_11326[27]), .Z(n_277261800));
	notech_or2 i_93644462(.A(n_55587), .B(n_308721974), .Z(n_275361781));
	notech_or2 i_94044459(.A(n_55842), .B(n_27594), .Z(n_275061778));
	notech_or2 i_94344456(.A(n_55597), .B(n_29156), .Z(n_274761775));
	notech_or2 i_94644453(.A(n_2212), .B(nbus_11326[26]), .Z(n_274461772));
	notech_or2 i_58444806(.A(n_354788261), .B(n_308621973), .Z(n_274161769)
		);
	notech_nand3 i_58744803(.A(n_59197), .B(n_59940), .C(read_data[27]), .Z(n_273861766
		));
	notech_or2 i_59044800(.A(n_353988269), .B(nbus_11273[27]), .Z(n_273561763
		));
	notech_nao3 i_59344797(.A(n_2468), .B(n_29091), .C(n_232761396), .Z(n_273261760
		));
	notech_or2 i_54844842(.A(n_308921976), .B(n_323662240), .Z(n_272961757)
		);
	notech_nand3 i_55144839(.A(n_59197), .B(n_59940), .C(read_data[23]), .Z(n_272661754
		));
	notech_or2 i_55444836(.A(n_353988269), .B(nbus_11273[23]), .Z(n_272361751
		));
	notech_nao3 i_55744833(.A(n_2460), .B(n_29091), .C(n_232761396), .Z(n_272061748
		));
	notech_and3 i_100344400(.A(n_56061), .B(n_279961827), .C(n_136060442), .Z
		(n_271761745));
	notech_and4 i_96348253(.A(n_270361731), .B(n_270261730), .C(n_265961687)
		, .D(n_270861736), .Z(n_271061738));
	notech_and3 i_96148255(.A(n_270661734), .B(n_270561733), .C(n_265861686)
		, .Z(n_270861736));
	notech_ao4 i_95348261(.A(n_55977), .B(n_28445), .C(n_262636781), .D(n_26987
		), .Z(n_270661734));
	notech_ao4 i_95848258(.A(n_55536), .B(n_58951), .C(n_55135), .D(n_27601)
		, .Z(n_270561733));
	notech_ao4 i_95548259(.A(n_262536780), .B(n_27554), .C(n_55535), .D(n_56943
		), .Z(n_270361731));
	notech_ao4 i_95448260(.A(n_308518862), .B(nbus_11326[31]), .C(n_56024), 
		.D(n_29150), .Z(n_270261730));
	notech_and4 i_75948437(.A(n_269861726), .B(n_269261720), .C(n_264361671)
		, .D(n_269661724), .Z(n_270061728));
	notech_ao4 i_75548440(.A(n_354888260), .B(n_28977), .C(n_353988269), .D(nbus_11273
		[29]), .Z(n_269861726));
	notech_and3 i_75348442(.A(n_269461722), .B(n_269361721), .C(n_264261670)
		, .Z(n_269661724));
	notech_ao4 i_75048445(.A(n_59168), .B(n_27552), .C(n_262236777), .D(n_29148
		), .Z(n_269461722));
	notech_ao4 i_75148444(.A(n_5538), .B(n_27597), .C(n_262336778), .D(n_29149
		), .Z(n_269361721));
	notech_ao4 i_75648439(.A(n_353488274), .B(nbus_11326[29]), .C(n_354488264
		), .D(\nbus_11276[29] ), .Z(n_269261720));
	notech_nao3 i_73348460(.A(n_268761715), .B(n_268661714), .C(n_263561663)
		, .Z(n_268961717));
	notech_ao4 i_73148462(.A(n_353488274), .B(nbus_11326[30]), .C(n_354488264
		), .D(\nbus_11276[30] ), .Z(n_268761715));
	notech_and4 i_73048463(.A(n_268361711), .B(n_268261710), .C(n_263161659)
		, .D(n_263261660), .Z(n_268661714));
	notech_ao4 i_72648467(.A(n_262336778), .B(n_29147), .C(n_262236777), .D(n_29146
		), .Z(n_268361711));
	notech_ao4 i_72748466(.A(n_5538), .B(n_27599), .C(n_27553), .D(n_59168),
		 .Z(n_268261710));
	notech_and4 i_71148482(.A(n_267761705), .B(n_267261700), .C(n_262461652)
		, .D(n_262361651), .Z(n_268061708));
	notech_and4 i_70748486(.A(n_267461702), .B(n_267361701), .C(n_261961647)
		, .D(n_262061648), .Z(n_267761705));
	notech_ao4 i_70348490(.A(n_262336778), .B(n_29145), .C(n_262236777), .D(n_29144
		), .Z(n_267461702));
	notech_ao4 i_70448489(.A(n_5538), .B(n_27601), .C(n_27554), .D(n_59168),
		 .Z(n_267361701));
	notech_ao4 i_70848485(.A(n_354488264), .B(n_56943), .C(n_353988269), .D(n_58951
		), .Z(n_267261700));
	notech_and2 i_53549179(.A(n_55846), .B(n_260161629), .Z(n_266461692));
	notech_and2 i_197760620(.A(n_231961388), .B(n_56260), .Z(n_266361691));
	notech_or4 i_3221739(.A(n_266061688), .B(n_266161689), .C(n_264961677), 
		.D(n_26437), .Z(n_12953));
	notech_nor2 i_95148263(.A(n_110123088), .B(n_271288743), .Z(n_266161689)
		);
	notech_nor2 i_94948265(.A(n_354688262), .B(n_28996), .Z(n_266061688));
	notech_nao3 i_95248262(.A(opc_10[31]), .B(n_62399), .C(n_110323090), .Z(n_265961687
		));
	notech_nand2 i_94848266(.A(sav_esp[31]), .B(n_60598), .Z(n_265861686));
	notech_nor2 i_95048264(.A(n_354588263), .B(n_271088745), .Z(n_264961677)
		);
	notech_nand3 i_3021193(.A(n_264861676), .B(n_270061728), .C(n_263861666)
		, .Z(n_13641));
	notech_nao3 i_74948446(.A(opc_10[29]), .B(n_62415), .C(n_354988259), .Z(n_264861676
		));
	notech_or2 i_74548450(.A(n_354788261), .B(n_57329), .Z(n_264361671));
	notech_nand2 i_74248453(.A(sav_edi[29]), .B(n_60598), .Z(n_264261670));
	notech_or2 i_74748448(.A(n_354388265), .B(n_270688747), .Z(n_263861666)
		);
	notech_or4 i_3121194(.A(n_263661664), .B(n_268961717), .C(n_263761665), 
		.D(n_262661654), .Z(n_13647));
	notech_nor2 i_72048473(.A(n_323462238), .B(n_28997), .Z(n_263761665));
	notech_nor2 i_72448469(.A(n_323762241), .B(n_271188744), .Z(n_263661664)
		);
	notech_ao3 i_72548468(.A(opc_10[30]), .B(n_62399), .C(n_3288), .Z(n_263561663
		));
	notech_or2 i_71948474(.A(n_353988269), .B(n_56901), .Z(n_263261660));
	notech_nand2 i_71848475(.A(sav_edi[30]), .B(n_60598), .Z(n_263161659));
	notech_nor2 i_72348470(.A(n_270988746), .B(n_323662240), .Z(n_262661654)
		);
	notech_nand3 i_3221195(.A(n_268061708), .B(n_262561653), .C(n_261461642)
		, .Z(n_13653));
	notech_or2 i_70148492(.A(n_354388265), .B(n_271288743), .Z(n_262561653)
		);
	notech_nao3 i_70248491(.A(opc_10[31]), .B(n_62415), .C(n_354988259), .Z(n_262461652
		));
	notech_or2 i_69948494(.A(n_353488274), .B(nbus_11326[31]), .Z(n_262361651
		));
	notech_or2 i_69848495(.A(n_354888260), .B(n_28996), .Z(n_262061648));
	notech_nand2 i_69548498(.A(sav_edi[31]), .B(n_60598), .Z(n_261961647));
	notech_or2 i_70048493(.A(n_354788261), .B(n_271088745), .Z(n_261461642)
		);
	notech_and3 i_27848888(.A(n_54900), .B(n_261436769), .C(n_226961338), .Z
		(n_261361641));
	notech_and4 i_23248932(.A(n_55846), .B(n_260161629), .C(n_260461632), .D
		(n_322962233), .Z(n_261261640));
	notech_and4 i_246349168(.A(n_54851), .B(n_54900), .C(n_54876), .D(n_26442
		), .Z(n_261161639));
	notech_nao3 i_152360558(.A(n_60532), .B(n_26772), .C(n_226061331), .Z(n_260961637
		));
	notech_ao4 i_21248952(.A(n_56163), .B(n_56121), .C(n_26443), .D(n_54151)
		, .Z(n_260661634));
	notech_or2 i_11730(.A(n_259561623), .B(n_266461692), .Z(n_260561633));
	notech_ao4 i_53349208(.A(n_56574), .B(n_204988864), .C(n_2241), .D(n_26226
		), .Z(n_260461632));
	notech_or2 i_11732(.A(n_266461692), .B(n_266361691), .Z(n_260261630));
	notech_or4 i_18948975(.A(n_260688757), .B(n_2605), .C(n_205088863), .D(n_26226
		), .Z(n_260161629));
	notech_or2 i_173249216(.A(n_266361691), .B(n_260461632), .Z(n_259861626)
		);
	notech_or2 i_176949215(.A(n_260461632), .B(n_259561623), .Z(n_259661624)
		);
	notech_or2 i_201260550(.A(n_225761328), .B(n_59224), .Z(n_259561623));
	notech_nand2 i_85351163(.A(n_259161619), .B(n_259061618), .Z(n_259261620
		));
	notech_ao4 i_84751165(.A(n_55397), .B(n_28987), .C(n_55396), .D(n_2700),
		 .Z(n_259161619));
	notech_ao4 i_84651166(.A(n_55071), .B(\nbus_11276[17] ), .C(n_55070), .D
		(nbus_11273[17]), .Z(n_259061618));
	notech_nand3 i_85051164(.A(n_43426147), .B(n_258161609), .C(n_258661614)
		, .Z(n_258961617));
	notech_or4 i_1820669(.A(n_259261620), .B(n_258961617), .C(n_258761615), 
		.D(n_258061608), .Z(n_19887));
	notech_ao3 i_84351168(.A(opc_10[17]), .B(n_62399), .C(n_306621953), .Z(n_258761615
		));
	notech_or4 i_84151170(.A(n_56201), .B(n_56163), .C(n_56376), .D(n_27583)
		, .Z(n_258661614));
	notech_or2 i_83451175(.A(n_303521922), .B(nbus_11326[17]), .Z(n_258161609
		));
	notech_nor2 i_84251169(.A(n_2648), .B(n_309921986), .Z(n_258061608));
	notech_and4 i_143053918(.A(n_53844), .B(n_257661604), .C(n_237661444), .D
		(n_26375), .Z(n_257961607));
	notech_ao4 i_142853920(.A(n_55220), .B(nbus_11273[24]), .C(n_55221), .D(\nbus_11276[24] 
		), .Z(n_257661604));
	notech_ao4 i_143253917(.A(n_55557), .B(n_29137), .C(n_55556), .D(n_57334
		), .Z(n_257461602));
	notech_ao4 i_143753916(.A(n_322631613), .B(n_322231609), .C(n_251061538)
		, .D(n_322931616), .Z(n_257261600));
	notech_and4 i_169753661(.A(n_256961597), .B(n_256761595), .C(n_238461452
		), .D(n_238761455), .Z(n_257161599));
	notech_ao4 i_169353665(.A(n_53993), .B(n_29138), .C(n_224461315), .D(n_29077
		), .Z(n_256961597));
	notech_ao4 i_169553663(.A(n_236961437), .B(\nbus_11276[10] ), .C(n_236861436
		), .D(nbus_11273[10]), .Z(n_256761595));
	notech_ao4 i_169853660(.A(n_59168), .B(n_27529), .C(n_59197), .D(n_26750
		), .Z(n_256461592));
	notech_and3 i_170253656(.A(n_239461462), .B(n_239361461), .C(n_256261590
		), .Z(n_256361591));
	notech_ao4 i_170053658(.A(n_174358031), .B(n_236661434), .C(n_318431571)
		, .D(n_60474), .Z(n_256261590));
	notech_and4 i_171053648(.A(n_255661584), .B(n_255461582), .C(n_239861466
		), .D(n_240161469), .Z(n_255861586));
	notech_ao4 i_170653652(.A(n_53993), .B(n_29139), .C(n_55427), .D(n_29080
		), .Z(n_255661584));
	notech_ao4 i_170853650(.A(n_55308), .B(\nbus_11276[11] ), .C(n_55307), .D
		(nbus_11273[11]), .Z(n_255461582));
	notech_and4 i_171553643(.A(n_255161579), .B(n_240761475), .C(n_254961577
		), .D(n_240461472), .Z(n_255361581));
	notech_ao4 i_171153647(.A(n_59168), .B(n_27530), .C(n_59197), .D(n_26752
		), .Z(n_255161579));
	notech_ao4 i_171353645(.A(n_171758005), .B(n_354188267), .C(n_171658004)
		, .D(n_354088268), .Z(n_254961577));
	notech_and4 i_173053628(.A(n_254661574), .B(n_254461572), .C(n_241061478
		), .D(n_241361481), .Z(n_254861576));
	notech_ao4 i_172653632(.A(n_53993), .B(n_29140), .C(n_55427), .D(n_29037
		), .Z(n_254661574));
	notech_ao4 i_172853630(.A(n_55308), .B(\nbus_11276[13] ), .C(n_55307), .D
		(nbus_11273[13]), .Z(n_254461572));
	notech_and4 i_173553623(.A(n_254161569), .B(n_241961487), .C(n_253961567
		), .D(n_241661484), .Z(n_254361571));
	notech_ao4 i_173153627(.A(n_59167), .B(n_27532), .C(n_59197), .D(n_26754
		), .Z(n_254161569));
	notech_ao4 i_173353625(.A(n_166557953), .B(n_354188267), .C(n_166457952)
		, .D(n_354088268), .Z(n_253961567));
	notech_and4 i_175053608(.A(n_253661564), .B(n_253461562), .C(n_242261490
		), .D(n_242561493), .Z(n_253861566));
	notech_ao4 i_174653612(.A(n_53993), .B(n_29141), .C(n_353488274), .D(nbus_11326
		[24]), .Z(n_253661564));
	notech_ao4 i_174853610(.A(n_354488264), .B(\nbus_11276[24] ), .C(n_57334
		), .D(n_323662240), .Z(n_253461562));
	notech_and4 i_175553603(.A(n_253161559), .B(n_252961557), .C(n_243861496
		), .D(n_244561499), .Z(n_253361561));
	notech_ao4 i_175153607(.A(n_27546), .B(n_59168), .C(n_5538), .D(n_27592)
		, .Z(n_253161559));
	notech_ao4 i_175353605(.A(n_322231609), .B(n_323762241), .C(n_251061538)
		, .D(n_3288), .Z(n_252961557));
	notech_nao3 i_68155298(.A(n_252561553), .B(n_252761555), .C(n_246761503)
		, .Z(n_252861556));
	notech_ao4 i_203053333(.A(n_27546), .B(n_59865), .C(n_98113375), .D(nbus_11273
		[24]), .Z(n_252761555));
	notech_ao4 i_203153332(.A(n_101213406), .B(n_57334), .C(n_101413408), .D
		(n_29137), .Z(n_252561553));
	notech_ao4 i_215953204(.A(n_56382), .B(n_29142), .C(n_56151), .D(n_27630
		), .Z(n_252261550));
	notech_ao4 i_216053203(.A(n_56126), .B(n_27671), .C(n_27707), .D(n_56097
		), .Z(n_252161549));
	notech_and2 i_216453199(.A(n_251961547), .B(n_251861546), .Z(n_252061548
		));
	notech_ao4 i_216253201(.A(n_54535), .B(n_27394), .C(n_55864), .D(n_27739
		), .Z(n_251961547));
	notech_ao4 i_216353200(.A(n_55898), .B(n_27778), .C(n_55879), .D(n_27842
		), .Z(n_251861546));
	notech_and4 i_217253191(.A(n_251561543), .B(n_251461542), .C(n_251261540
		), .D(n_251161539), .Z(n_251761545));
	notech_ao4 i_216653197(.A(n_56068), .B(n_27877), .C(n_56035), .D(n_27911
		), .Z(n_251561543));
	notech_ao4 i_216753196(.A(n_56009), .B(n_27945), .C(n_55998), .D(n_27977
		), .Z(n_251461542));
	notech_ao4 i_216953194(.A(n_55872), .B(n_28011), .C(n_55873), .D(n_29143
		), .Z(n_251261540));
	notech_ao4 i_217053193(.A(n_55878), .B(n_28043), .C(n_55940), .D(n_27810
		), .Z(n_251161539));
	notech_nand2 i_2655312(.A(opc_10[24]), .B(n_62431), .Z(n_251061538));
	notech_or4 i_220953154(.A(fsmf[4]), .B(fsmf[2]), .C(fsmf[3]), .D(n_51741
		), .Z(n_250861536));
	notech_or4 i_221253151(.A(fsmf[0]), .B(fsmf[1]), .C(instrc[6]), .D(instrc
		[4]), .Z(n_250561533));
	notech_or4 i_221653147(.A(instrc[7]), .B(instrc[5]), .C(instrc[1]), .D(instrc
		[3]), .Z(n_250161529));
	notech_or4 i_221953144(.A(instrc[2]), .B(n_28499), .C(n_26226), .D(n_29009
		), .Z(n_249861526));
	notech_nao3 i_31679(.A(n_57433), .B(n_26243), .C(n_2647), .Z(n_249261520
		));
	notech_nor2 i_98954350(.A(n_56057), .B(\nbus_11276[24] ), .Z(n_246761503
		));
	notech_nand2 i_64954673(.A(sav_edi[24]), .B(n_60598), .Z(n_244561499));
	notech_or2 i_65254670(.A(n_323462238), .B(n_29137), .Z(n_243861496));
	notech_or2 i_65554667(.A(n_353988269), .B(nbus_11273[24]), .Z(n_242561493
		));
	notech_nao3 i_65854664(.A(n_2462), .B(n_29091), .C(n_232761396), .Z(n_242261490
		));
	notech_or4 i_61754697(.A(n_273588720), .B(n_59281), .C(n_2240), .D(n_321831605
		), .Z(n_241961487));
	notech_nand2 i_62054694(.A(opd[13]), .B(n_55728), .Z(n_241661484));
	notech_or2 i_62354691(.A(n_57345), .B(n_55426), .Z(n_241361481));
	notech_nao3 i_62854688(.A(n_2440), .B(n_29091), .C(n_54015), .Z(n_241061478
		));
	notech_or4 i_59054721(.A(n_273588720), .B(n_59281), .C(n_2240), .D(n_322031607
		), .Z(n_240761475));
	notech_nand2 i_59354718(.A(n_55728), .B(opd[11]), .Z(n_240461472));
	notech_or2 i_59654715(.A(n_57347), .B(n_55426), .Z(n_240161469));
	notech_nao3 i_60154712(.A(n_2436), .B(n_29091), .C(n_54015), .Z(n_239861466
		));
	notech_ao4 i_31060722(.A(n_56061), .B(n_60598), .C(n_26226), .D(n_56053)
		, .Z(n_239561463));
	notech_or4 i_57554735(.A(n_55859), .B(n_55878), .C(n_322131608), .D(n_60598
		), .Z(n_239461462));
	notech_or4 i_57354736(.A(n_323062234), .B(n_239561463), .C(n_28061), .D(n_60512
		), .Z(n_239361461));
	notech_or2 i_58154730(.A(n_236761435), .B(n_27575), .Z(n_239061458));
	notech_or2 i_58454727(.A(n_57348), .B(n_237061438), .Z(n_238761455));
	notech_nao3 i_58754724(.A(n_2434), .B(n_55450), .C(n_54015), .Z(n_238461452
		));
	notech_or4 i_26555040(.A(n_56074), .B(n_206288851), .C(n_56376), .D(n_27592
		), .Z(n_238161449));
	notech_or2 i_27055035(.A(n_303421921), .B(nbus_11326[24]), .Z(n_237661444
		));
	notech_or2 i_120354142(.A(n_36952), .B(n_55864), .Z(n_237361441));
	notech_ao4 i_121960665(.A(n_54874), .B(n_56551), .C(n_239561463), .D(n_259561623
		), .Z(n_237061438));
	notech_and4 i_151260651(.A(n_54781), .B(n_55422), .C(n_56022), .D(n_232461393
		), .Z(n_236961437));
	notech_and3 i_150260655(.A(n_54710), .B(n_225661327), .C(n_353988269), .Z
		(n_236861436));
	notech_and3 i_151160652(.A(n_5538), .B(n_5577), .C(n_231161380), .Z(n_236761435
		));
	notech_and2 i_140060659(.A(n_261136766), .B(n_225361324), .Z(n_236661434
		));
	notech_and4 i_144959215(.A(n_144577845), .B(n_183678231), .C(n_130277702
		), .D(n_236361431), .Z(n_236461432));
	notech_ao4 i_144859216(.A(n_57352), .B(n_259661624), .C(n_259861626), .D
		(n_29068), .Z(n_236361431));
	notech_ao4 i_145059214(.A(n_59197), .B(n_26746), .C(n_53993), .D(n_29133
		), .Z(n_236161429));
	notech_and4 i_145759207(.A(n_235861426), .B(n_235661424), .C(n_227961348
		), .D(n_228261351), .Z(n_236061428));
	notech_ao4 i_145359211(.A(\nbus_11276[6] ), .B(n_224861319), .C(nbus_11273
		[6]), .D(n_224761318), .Z(n_235861426));
	notech_ao4 i_145559209(.A(n_27568), .B(n_224561316), .C(n_235561423), .D
		(n_323062234), .Z(n_235661424));
	notech_nao3 i_145859206(.A(opc_10[6]), .B(n_62399), .C(n_260461632), .Z(n_235561423
		));
	notech_and4 i_146059204(.A(n_150874376), .B(n_158074448), .C(n_137474242
		), .D(n_235261420), .Z(n_235361421));
	notech_ao4 i_145959205(.A(n_57351), .B(n_259661624), .C(n_28983), .D(n_259861626
		), .Z(n_235261420));
	notech_ao4 i_146159203(.A(n_59197), .B(n_26747), .C(n_53993), .D(n_29134
		), .Z(n_234961418));
	notech_and4 i_146859196(.A(n_234661415), .B(n_234261411), .C(n_229061359
		), .D(n_229361362), .Z(n_234861417));
	notech_ao4 i_146459200(.A(n_224861319), .B(\nbus_11276[7] ), .C(n_224761318
		), .D(nbus_11273[7]), .Z(n_234661415));
	notech_ao4 i_146659198(.A(n_224561316), .B(n_27570), .C(n_323062234), .D
		(n_234161410), .Z(n_234261411));
	notech_nao3 i_147159193(.A(opc_10[7]), .B(n_62431), .C(n_260461632), .Z(n_234161410
		));
	notech_and4 i_147859188(.A(n_233861407), .B(n_233661405), .C(n_229661365
		), .D(n_229961368), .Z(n_234061409));
	notech_ao4 i_147259192(.A(n_59197), .B(n_26749), .C(n_57349), .D(n_237061438
		), .Z(n_233861407));
	notech_ao4 i_147659190(.A(nbus_11273[9]), .B(n_236861436), .C(n_27574), 
		.D(n_236761435), .Z(n_233661405));
	notech_ao4 i_147959187(.A(n_53993), .B(n_29136), .C(n_262236777), .D(n_29135
		), .Z(n_233361402));
	notech_and3 i_148359183(.A(n_230661375), .B(n_230561374), .C(n_233161400
		), .Z(n_233261401));
	notech_ao4 i_148159185(.A(n_29048), .B(n_224461315), .C(n_260636761), .D
		(n_60474), .Z(n_233161400));
	notech_or4 i_166360610(.A(n_60782), .B(n_60729), .C(n_225161322), .D(n_60598
		), .Z(n_232761396));
	notech_and3 i_169258990(.A(n_230961378), .B(n_230861377), .C(n_231061379
		), .Z(n_232461393));
	notech_ao4 i_170258981(.A(n_2263), .B(n_26379), .C(n_225761328), .D(n_26321
		), .Z(n_231961388));
	notech_and2 i_31260601(.A(n_54851), .B(n_225961330), .Z(n_231861387));
	notech_ao4 i_170658977(.A(n_2263), .B(n_26382), .C(n_226061331), .D(n_26597
		), .Z(n_231761386));
	notech_nand2 i_29071(.A(n_56465), .B(n_29010), .Z(n_231461383));
	notech_or4 i_84659765(.A(n_206288851), .B(n_56063), .C(n_273588720), .D(n_60598
		), .Z(n_231161380));
	notech_or4 i_84559766(.A(calc_sz[3]), .B(calc_sz[2]), .C(n_260688757), .D
		(n_54874), .Z(n_231061379));
	notech_or2 i_84459767(.A(n_259561623), .B(n_231861387), .Z(n_230961378)
		);
	notech_or4 i_84359768(.A(n_57374), .B(n_60598), .C(n_59940), .D(n_26599)
		, .Z(n_230861377));
	notech_or4 i_64959947(.A(n_55859), .B(n_57299), .C(n_55878), .D(n_60595)
		, .Z(n_230661375));
	notech_or4 i_64859948(.A(n_239561463), .B(n_323062234), .C(n_28060), .D(n_60512
		), .Z(n_230561374));
	notech_or2 i_65559942(.A(n_236961437), .B(\nbus_11276[9] ), .Z(n_230261371
		));
	notech_nao3 i_65959939(.A(n_62427), .B(opc[9]), .C(n_236661434), .Z(n_229961368
		));
	notech_nand3 i_66359936(.A(n_59197), .B(n_59940), .C(read_data[9]), .Z(n_229661365
		));
	notech_nand3 i_63659959(.A(n_224661317), .B(opc[7]), .C(n_62401), .Z(n_229361362
		));
	notech_nao3 i_63959956(.A(n_2428), .B(n_55450), .C(n_54015), .Z(n_229061359
		));
	notech_or4 i_64259953(.A(n_58487), .B(n_2675), .C(n_56574), .D(n_205088863
		), .Z(n_228761356));
	notech_nand3 i_62359971(.A(n_62427), .B(opc[6]), .C(n_224661317), .Z(n_228261351
		));
	notech_nao3 i_62759968(.A(n_2426), .B(n_55450), .C(n_54015), .Z(n_227961348
		));
	notech_or4 i_63059965(.A(n_56574), .B(n_205088863), .C(n_58483), .D(n_57320
		), .Z(n_227661345));
	notech_nao3 i_88359733(.A(n_59197), .B(n_58483), .C(n_55820), .Z(n_226961338
		));
	notech_ao4 i_84260582(.A(n_59380), .B(n_62431), .C(n_2264), .D(n_26382),
		 .Z(n_226061331));
	notech_nao3 i_86159753(.A(n_59197), .B(n_58483), .C(n_56063), .Z(n_225961330
		));
	notech_ao4 i_179960554(.A(n_59380), .B(n_62431), .C(n_2264), .D(n_26379)
		, .Z(n_225761328));
	notech_or2 i_85759757(.A(n_266361691), .B(n_231861387), .Z(n_225661327)
		);
	notech_and3 i_3760518(.A(n_54851), .B(n_225961330), .C(n_56040), .Z(n_225461325
		));
	notech_or2 i_84859763(.A(n_323062234), .B(n_225461325), .Z(n_225361324)
		);
	notech_ao4 i_83759773(.A(n_1901), .B(n_273288723), .C(n_272688729), .D(n_274988708
		), .Z(n_225161322));
	notech_and3 i_6160494(.A(n_55846), .B(n_260161629), .C(n_56040), .Z(n_225061321
		));
	notech_or2 i_64759949(.A(n_323062234), .B(n_225061321), .Z(n_224961320)
		);
	notech_and3 i_139660561(.A(n_322662230), .B(n_260561633), .C(n_54781), .Z
		(n_224861319));
	notech_and3 i_139760560(.A(n_322762231), .B(n_260261630), .C(n_54893), .Z
		(n_224761318));
	notech_nand2 i_139960559(.A(n_354088268), .B(n_224961320), .Z(n_224661317
		));
	notech_and3 i_6060495(.A(n_5538), .B(n_323162235), .C(n_354288266), .Z(n_224561316
		));
	notech_or2 i_175560585(.A(n_266361691), .B(n_239561463), .Z(n_224461315)
		);
	notech_and4 i_119762391(.A(n_355888239), .B(n_224161312), .C(n_223961310
		), .D(n_149560577), .Z(n_224361314));
	notech_ao4 i_119262395(.A(n_353488274), .B(nbus_11326[17]), .C(n_63826342
		), .D(n_3288), .Z(n_224161312));
	notech_ao4 i_119462393(.A(n_2700), .B(n_323662240), .C(n_323462238), .D(n_28987
		), .Z(n_223961310));
	notech_and4 i_120262386(.A(n_223661307), .B(n_223461305), .C(n_149860580
		), .D(n_150160583), .Z(n_223861309));
	notech_ao4 i_119862390(.A(n_262236777), .B(n_29132), .C(n_53993), .D(n_29131
		), .Z(n_223661307));
	notech_ao4 i_120062388(.A(n_2648), .B(n_323762241), .C(n_59197), .D(n_26758
		), .Z(n_223461305));
	notech_ao4 i_147462118(.A(n_29020), .B(n_29023), .C(instrc[90]), .D(n_26545
		), .Z(n_223361304));
	notech_ao4 i_149662096(.A(n_56425), .B(n_26925), .C(n_151760599), .D(n_28052
		), .Z(n_222461295));
	notech_ao4 i_149762095(.A(n_151960601), .B(n_27298), .C(n_152060602), .D
		(n_27334), .Z(n_222261294));
	notech_nand2 i_5363494(.A(instrc[125]), .B(instrc[127]), .Z(n_221961291)
		);
	notech_nao3 i_1263535(.A(instrc[127]), .B(instrc[126]), .C(instrc[125]),
		 .Z(n_221861290));
	notech_and4 i_150862084(.A(n_54860), .B(n_153760619), .C(n_152260604), .D
		(n_216961242), .Z(n_221661288));
	notech_ao4 i_150962083(.A(n_191060984), .B(n_2739), .C(n_148060562), .D(n_352765816
		), .Z(n_221361285));
	notech_ao4 i_151062082(.A(n_60484), .B(n_185560929), .C(n_56023), .D(n_148160563
		), .Z(n_221161284));
	notech_and4 i_151962073(.A(n_153060612), .B(n_220861281), .C(n_220461277
		), .D(n_26463), .Z(n_221061283));
	notech_ao4 i_151362079(.A(n_147960561), .B(n_138360465), .C(n_187860952)
		, .D(n_213361207), .Z(n_220861281));
	notech_ao4 i_152062072(.A(n_352765816), .B(n_182360897), .C(n_148160563)
		, .D(n_138360465), .Z(n_220661279));
	notech_or4 i_152162071(.A(n_351565804), .B(instrc[124]), .C(instrc[126])
		, .D(n_60563), .Z(n_220561278));
	notech_and4 i_151862074(.A(n_153260614), .B(n_153160613), .C(n_153360615
		), .D(n_153460616), .Z(n_220461277));
	notech_and4 i_71163558(.A(n_153760619), .B(n_154160623), .C(n_219661269)
		, .D(n_54860), .Z(n_219961272));
	notech_ao4 i_152962063(.A(n_207461148), .B(n_138760469), .C(n_138660468)
		, .D(n_219061263), .Z(n_219661269));
	notech_mux2 i_154862045(.S(n_54535), .A(n_141760499), .B(n_139160473), .Z
		(n_219561268));
	notech_nand2 i_863539(.A(n_139560477), .B(n_320888481), .Z(n_219361266)
		);
	notech_or4 i_155262041(.A(instrc[125]), .B(n_29032), .C(instrc[126]), .D
		(instrc[127]), .Z(n_219061263));
	notech_or4 i_153662057(.A(n_154860630), .B(n_154760629), .C(n_26467), .D
		(n_154560627), .Z(n_218561258));
	notech_and2 i_154662047(.A(n_29013), .B(n_29016), .Z(n_217461247));
	notech_or4 i_4063507(.A(n_275388704), .B(n_177660858), .C(n_26629), .D(n_59168
		), .Z(n_217361246));
	notech_and4 i_155662038(.A(n_54860), .B(n_153760619), .C(n_155360635), .D
		(n_216961242), .Z(n_217161244));
	notech_ao4 i_7963468(.A(n_2204), .B(n_2180), .C(n_60474), .D(n_216861241
		), .Z(n_216961242));
	notech_or2 i_156862026(.A(n_55843), .B(nZF), .Z(n_216861241));
	notech_ao4 i_155762037(.A(n_191060984), .B(n_2740), .C(n_2689), .D(n_148060562
		), .Z(n_216661239));
	notech_ao4 i_155862036(.A(n_185560929), .B(n_197114365), .C(n_148160563)
		, .D(n_55879), .Z(n_216561238));
	notech_and4 i_156762027(.A(n_216261235), .B(n_216061234), .C(n_215861232
		), .D(n_215561229), .Z(n_216461237));
	notech_ao4 i_156162033(.A(n_147960561), .B(n_139960481), .C(n_199961073)
		, .D(n_191760991), .Z(n_216261235));
	notech_ao4 i_156262032(.A(n_192861002), .B(n_197861052), .C(n_213661210)
		, .D(n_137960461), .Z(n_216061234));
	notech_ao4 i_156462030(.A(n_213261206), .B(n_137360455), .C(n_139860480)
		, .D(n_26227), .Z(n_215861232));
	notech_ao4 i_156962025(.A(n_2689), .B(n_182360897), .C(n_148160563), .D(n_139960481
		), .Z(n_215761231));
	notech_or4 i_157062024(.A(n_2658), .B(instrc[124]), .C(instrc[126]), .D(n_60563
		), .Z(n_215661230));
	notech_ao4 i_156562029(.A(n_212861202), .B(n_193161005), .C(n_213361207)
		, .D(n_203561109), .Z(n_215561229));
	notech_and3 i_157462020(.A(n_54860), .B(n_153760619), .C(n_215261226), .Z
		(n_215361227));
	notech_ao4 i_157362021(.A(n_184760921), .B(n_258764904), .C(n_1912), .D(n_191060984
		), .Z(n_215261226));
	notech_or4 i_158862006(.A(opa[7]), .B(opa[5]), .C(opa[2]), .D(n_214961223
		), .Z(n_215061224));
	notech_or4 i_158562009(.A(opa[3]), .B(n_59726), .C(opa[1]), .D(nbus_11273
		[0]), .Z(n_214961223));
	notech_or4 i_159162003(.A(n_249261520), .B(n_56067), .C(n_60595), .D(n_59940
		), .Z(n_214461218));
	notech_ao4 i_157562019(.A(n_148060562), .B(n_243964756), .C(n_57343), .D
		(n_185560929), .Z(n_214161215));
	notech_ao4 i_157662018(.A(n_148160563), .B(n_55898), .C(n_147960561), .D
		(n_140560487), .Z(n_214061214));
	notech_and4 i_158462010(.A(n_157660658), .B(n_213761211), .C(n_213461208
		), .D(n_213161205), .Z(n_213961213));
	notech_ao4 i_157962015(.A(n_197861052), .B(n_188660960), .C(n_213661210)
		, .D(n_189660970), .Z(n_213761211));
	notech_or2 i_15363398(.A(n_57162), .B(n_199761071), .Z(n_213661210));
	notech_ao4 i_158162013(.A(n_213361207), .B(n_190160975), .C(n_190260976)
		, .D(n_213261206), .Z(n_213461208));
	notech_nand2 i_11763433(.A(n_29014), .B(n_29017), .Z(n_213361207));
	notech_nand3 i_15763394(.A(n_26531), .B(n_29016), .C(n_29013), .Z(n_213261206
		));
	notech_ao4 i_158262012(.A(n_140460486), .B(n_26512), .C(n_188460958), .D
		(n_212861202), .Z(n_213161205));
	notech_ao4 i_159362001(.A(n_243964756), .B(n_182360897), .C(n_148160563)
		, .D(n_140560487), .Z(n_213061204));
	notech_or4 i_159462000(.A(n_29032), .B(instrc[126]), .C(n_60563), .D(n_26235
		), .Z(n_212961203));
	notech_nao3 i_159561999(.A(n_29029), .B(instrc[101]), .C(n_180560886), .Z
		(n_212861202));
	notech_ao4 i_159661998(.A(n_275288705), .B(n_2005), .C(n_55248), .D(n_60474
		), .Z(n_212661200));
	notech_ao4 i_159761997(.A(n_335162249), .B(n_353688272), .C(n_59197), .D
		(n_26684), .Z(n_212561199));
	notech_or4 i_160461990(.A(temp_sp[1]), .B(temp_sp[0]), .C(temp_sp[2]), .D
		(temp_sp[3]), .Z(n_212061194));
	notech_or4 i_160761987(.A(temp_sp[4]), .B(temp_sp[6]), .C(temp_sp[5]), .D
		(temp_sp[7]), .Z(n_211761191));
	notech_or4 i_161561979(.A(temp_sp[8]), .B(n_211061184), .C(temp_sp[9]), 
		.D(n_211161185), .Z(n_211461188));
	notech_nand2 i_161061984(.A(n_26943), .B(n_26945), .Z(n_211161185));
	notech_or4 i_161461980(.A(temp_sp[12]), .B(temp_sp[13]), .C(temp_sp[15])
		, .D(temp_sp[14]), .Z(n_211061184));
	notech_or4 i_163161963(.A(n_210561179), .B(n_210261176), .C(n_209861172)
		, .D(n_209561169), .Z(n_210761181));
	notech_or4 i_161961975(.A(temp_sp[18]), .B(temp_sp[19]), .C(temp_sp[17])
		, .D(temp_sp[16]), .Z(n_210561179));
	notech_or4 i_162261972(.A(temp_sp[20]), .B(temp_sp[21]), .C(temp_sp[22])
		, .D(temp_sp[23]), .Z(n_210261176));
	notech_or4 i_162661968(.A(temp_sp[25]), .B(temp_sp[26]), .C(temp_sp[27])
		, .D(temp_sp[24]), .Z(n_209861172));
	notech_or4 i_162961965(.A(temp_sp[29]), .B(temp_sp[28]), .C(temp_sp[31])
		, .D(temp_sp[30]), .Z(n_209561169));
	notech_ao4 i_160061994(.A(n_140960491), .B(n_207461148), .C(n_140860490)
		, .D(n_207361147), .Z(n_208461158));
	notech_ao4 i_163861956(.A(n_56583), .B(n_141860500), .C(n_55998), .D(n_141760499
		), .Z(n_208361157));
	notech_and4 i_6663481(.A(n_55667), .B(n_56058), .C(n_55658), .D(n_56059)
		, .Z(n_208061154));
	notech_nand2 i_563542(.A(n_260961637), .B(n_142460506), .Z(n_207661150)
		);
	notech_or2 i_763540(.A(tcmp), .B(n_60595), .Z(n_207461148));
	notech_or4 i_663541(.A(n_2193), .B(n_26496), .C(n_4737261), .D(n_349288316
		), .Z(n_207361147));
	notech_ao4 i_164461950(.A(n_142860510), .B(n_342262316), .C(n_335062248)
		, .D(n_142760509), .Z(n_207261146));
	notech_ao4 i_12463427(.A(n_334862246), .B(n_54703), .C(n_334962247), .D(n_55089
		), .Z(n_207161145));
	notech_and4 i_164961945(.A(n_206861142), .B(n_206661140), .C(n_160660688
		), .D(n_160960691), .Z(n_207061144));
	notech_ao4 i_164561949(.A(n_148060562), .B(n_294261946), .C(n_56240), .D
		(n_185560929), .Z(n_206861142));
	notech_ao4 i_164761947(.A(n_147960561), .B(n_144560527), .C(n_199861072)
		, .D(n_178060862), .Z(n_206661140));
	notech_nao3 i_165061944(.A(n_206261136), .B(n_144660528), .C(n_161060692
		), .Z(n_206361137));
	notech_ao4 i_165661938(.A(n_182360897), .B(n_294261946), .C(n_148160563)
		, .D(n_144560527), .Z(n_206261136));
	notech_or4 i_165461940(.A(n_161360695), .B(n_161260694), .C(n_161560697)
		, .D(n_26481), .Z(n_205861132));
	notech_and4 i_166861926(.A(n_54707), .B(n_205061124), .C(n_204861122), .D
		(n_162160703), .Z(n_205261126));
	notech_ao4 i_166461930(.A(n_59195), .B(n_26630), .C(n_56270), .D(n_185560929
		), .Z(n_205061124));
	notech_ao4 i_166661928(.A(n_135060432), .B(n_199961073), .C(n_197861052)
		, .D(n_162960711), .Z(n_204861122));
	notech_ao4 i_166961925(.A(n_320988480), .B(n_185960933), .C(n_353788271)
		, .D(n_166160743), .Z(n_204561119));
	notech_or4 i_167361921(.A(n_162860710), .B(n_162760709), .C(n_162660708)
		, .D(n_162560707), .Z(n_204461118));
	notech_and4 i_167961915(.A(n_317088519), .B(n_55688), .C(n_163060712), .D
		(n_319988490), .Z(n_204061114));
	notech_nao3 i_168361911(.A(n_184460918), .B(instrc[89]), .C(instrc[88]),
		 .Z(n_203561109));
	notech_or4 i_21441(.A(n_164260724), .B(n_164160723), .C(n_164460726), .D
		(n_164360725), .Z(n_203261106));
	notech_and2 i_170461890(.A(instrc[92]), .B(instrc[95]), .Z(n_202261096)
		);
	notech_ao4 i_170661888(.A(n_2261), .B(n_26524), .C(n_2255), .D(n_26523),
		 .Z(n_202061094));
	notech_or2 i_168761907(.A(n_163560717), .B(n_60596), .Z(n_201661090));
	notech_ao4 i_168861906(.A(n_57378), .B(n_144960531), .C(n_1900), .D(n_55247
		), .Z(n_201561089));
	notech_or2 i_169061904(.A(n_54530), .B(n_60563), .Z(n_201361087));
	notech_nao3 i_1363534(.A(n_26390), .B(\opcode[3] ), .C(n_56197), .Z(n_200961083
		));
	notech_ao4 i_104263576(.A(n_144960531), .B(n_57374), .C(n_200661080), .D
		(n_26887), .Z(n_200861082));
	notech_or4 i_6063487(.A(tcmp), .B(n_221961291), .C(n_29032), .D(n_28970)
		, .Z(n_200761081));
	notech_or4 i_169461900(.A(n_273288723), .B(n_275288705), .C(n_2258), .D(reps
		[2]), .Z(n_200661080));
	notech_and4 i_171661878(.A(n_54015), .B(n_200361077), .C(n_200161075), .D
		(n_200061074), .Z(n_200561079));
	notech_ao4 i_171161883(.A(n_59193), .B(n_26630), .C(n_134960431), .D(n_58483
		), .Z(n_200361077));
	notech_ao4 i_171361881(.A(n_59224), .B(n_185560929), .C(n_1912), .D(n_183460908
		), .Z(n_200161075));
	notech_ao4 i_171461880(.A(n_199961073), .B(n_179160873), .C(n_189660970)
		, .D(n_199861072), .Z(n_200061074));
	notech_nao3 i_11963432(.A(instrc[125]), .B(n_29028), .C(n_176360845), .Z
		(n_199961073));
	notech_nand2 i_14563406(.A(n_57162), .B(n_26489), .Z(n_199861072));
	notech_nand2 i_7163476(.A(n_177960861), .B(n_29040), .Z(n_199761071));
	notech_ao4 i_171761877(.A(n_184060914), .B(n_190160975), .C(n_3288), .D(n_166160743
		), .Z(n_199461068));
	notech_or4 i_172161873(.A(n_165760739), .B(n_166060742), .C(n_165860740)
		, .D(n_165960741), .Z(n_199361067));
	notech_and4 i_172461870(.A(n_260561633), .B(n_259661624), .C(n_322662230
		), .D(n_54781), .Z(n_199161065));
	notech_nand2 i_83163552(.A(instrc[125]), .B(n_29028), .Z(n_198661060));
	notech_and2 i_6863479(.A(n_29016), .B(n_26531), .Z(n_198461058));
	notech_and2 i_6963478(.A(n_29029), .B(n_26528), .Z(n_198161055));
	notech_and2 i_11463435(.A(instrc[101]), .B(instrc[102]), .Z(n_198061054)
		);
	notech_nand3 i_12163430(.A(n_183060904), .B(n_29030), .C(instrc[93]), .Z
		(n_197861052));
	notech_and4 i_173661858(.A(n_166660748), .B(n_197461048), .C(n_197261046
		), .D(n_166960751), .Z(n_197661050));
	notech_ao4 i_173261862(.A(n_263436789), .B(n_148060562), .C(n_56290), .D
		(n_185560929), .Z(n_197461048));
	notech_ao4 i_173461860(.A(n_147960561), .B(n_145860540), .C(n_187860952)
		, .D(n_189960973), .Z(n_197261046));
	notech_ao4 i_148664231(.A(n_55763), .B(n_29130), .C(n_2822), .D(n_353776373
		), .Z(n_125874126));
	notech_nor2 i_12663425(.A(n_54523), .B(n_281539603), .Z(n_126074128));
	notech_or4 i_13463417(.A(n_1916), .B(n_148560567), .C(n_281539603), .D(n_59235
		), .Z(n_126174129));
	notech_and4 i_67662894(.A(n_55667), .B(n_136060442), .C(n_55999), .D(n_281539603
		), .Z(n_126274130));
	notech_or2 i_67962891(.A(n_55580), .B(n_55872), .Z(n_126374131));
	notech_or2 i_50163064(.A(n_356176397), .B(n_29063), .Z(n_126474132));
	notech_nand2 i_49663069(.A(opa[4]), .B(n_54661), .Z(n_127174139));
	notech_or2 i_51663049(.A(n_356176397), .B(n_29068), .Z(n_127274140));
	notech_nand2 i_51163054(.A(n_54661), .B(n_59735), .Z(n_127974147));
	notech_or2 i_52463041(.A(n_356176397), .B(n_28983), .Z(n_128074148));
	notech_nand2 i_51963046(.A(n_54661), .B(opa[7]), .Z(n_128774155));
	notech_or2 i_59662972(.A(n_54468), .B(n_29063), .Z(n_128874156));
	notech_nand2 i_59062977(.A(opa[4]), .B(n_2670), .Z(n_129574163));
	notech_or2 i_61162957(.A(n_54468), .B(n_29068), .Z(n_129674164));
	notech_nand2 i_60662962(.A(n_2670), .B(opa[6]), .Z(n_130374171));
	notech_or2 i_61962949(.A(n_54468), .B(n_28983), .Z(n_130474172));
	notech_nand2 i_61462954(.A(n_2670), .B(opa[7]), .Z(n_131174179));
	notech_or4 i_67562895(.A(n_56197), .B(n_56163), .C(n_55820), .D(n_2675),
		 .Z(n_131274180));
	notech_or2 i_67062900(.A(n_54438), .B(n_28983), .Z(n_131974187));
	notech_ao4 i_145862134(.A(n_279739585), .B(n_2680), .C(n_275539543), .D(n_2679
		), .Z(n_132574193));
	notech_ao4 i_145762135(.A(\nbus_11276[7] ), .B(n_54655), .C(n_57351), .D
		(n_54469), .Z(n_132774195));
	notech_ao4 i_145562137(.A(n_55756), .B(n_27570), .C(n_54656), .D(nbus_11273
		[7]), .Z(n_132974197));
	notech_and4 i_145662136(.A(n_174064078), .B(n_173964077), .C(n_131274180
		), .D(n_132974197), .Z(n_133174199));
	notech_ao4 i_141162181(.A(n_56151), .B(n_251734143), .C(n_27570), .D(n_2671
		), .Z(n_133274200));
	notech_ao4 i_141062182(.A(n_2685), .B(n_2679), .C(n_2669), .D(\nbus_11276[7] 
		), .Z(n_133474202));
	notech_ao4 i_140862184(.A(n_54428), .B(n_57351), .C(n_2680), .D(n_2684),
		 .Z(n_133674204));
	notech_and4 i_140962183(.A(n_174064078), .B(n_173964077), .C(n_133674204
		), .D(n_130474172), .Z(n_133874206));
	notech_ao4 i_140462188(.A(n_144377843), .B(n_56151), .C(n_2671), .D(n_27568
		), .Z(n_133974207));
	notech_ao4 i_140362189(.A(n_2685), .B(n_316588524), .C(\nbus_11276[6] ),
		 .D(n_2669), .Z(n_134174209));
	notech_ao4 i_140162191(.A(n_54428), .B(n_57352), .C(n_2684), .D(n_316488525
		), .Z(n_134374211));
	notech_and4 i_140262190(.A(n_183578230), .B(n_183478229), .C(n_134374211
		), .D(n_129674164), .Z(n_134574213));
	notech_ao4 i_139062202(.A(n_139770716), .B(n_56151), .C(n_2671), .D(n_27565
		), .Z(n_134674214));
	notech_ao4 i_138962203(.A(n_2685), .B(n_316288527), .C(n_2669), .D(\nbus_11276[4] 
		), .Z(n_134874216));
	notech_ao4 i_138762205(.A(n_54428), .B(n_321188478), .C(n_2684), .D(n_316388526
		), .Z(n_135074218));
	notech_and3 i_138862204(.A(n_137970698), .B(n_135074218), .C(n_128874156
		), .Z(n_135274220));
	notech_ao4 i_132662265(.A(n_56049), .B(n_251734143), .C(n_55753), .D(n_27570
		), .Z(n_135374221));
	notech_ao4 i_132562266(.A(n_2679), .B(n_356376399), .C(n_54631), .D(\nbus_11276[7] 
		), .Z(n_135574223));
	notech_ao4 i_132362268(.A(n_57351), .B(n_356076396), .C(n_2680), .D(n_356276398
		), .Z(n_135774225));
	notech_and4 i_132462267(.A(n_174064078), .B(n_173964077), .C(n_135774225
		), .D(n_128074148), .Z(n_135974227));
	notech_ao4 i_131962272(.A(n_144377843), .B(n_56043), .C(n_55753), .D(n_27568
		), .Z(n_136074228));
	notech_ao4 i_131862273(.A(n_316588524), .B(n_356376399), .C(\nbus_11276[6] 
		), .D(n_54631), .Z(n_136274230));
	notech_ao4 i_131662275(.A(n_57352), .B(n_356076396), .C(n_316488525), .D
		(n_356276398), .Z(n_136474232));
	notech_and4 i_131762274(.A(n_183578230), .B(n_183478229), .C(n_136474232
		), .D(n_127274140), .Z(n_136674234));
	notech_ao4 i_130362286(.A(n_139770716), .B(n_56043), .C(n_55753), .D(n_27565
		), .Z(n_136774235));
	notech_ao4 i_130262287(.A(n_316288527), .B(n_356376399), .C(n_54631), .D
		(\nbus_11276[4] ), .Z(n_136974237));
	notech_ao4 i_130062289(.A(n_321188478), .B(n_356076396), .C(n_316388526)
		, .D(n_356276398), .Z(n_137174239));
	notech_and3 i_130162288(.A(n_137970698), .B(n_137174239), .C(n_126474132
		), .Z(n_137374241));
	notech_nand3 i_64659950(.A(n_59193), .B(n_59940), .C(read_data[7]), .Z(n_137474242
		));
	notech_and2 i_83159779(.A(n_2673), .B(n_2651), .Z(n_137574243));
	notech_or2 i_87159745(.A(n_36952), .B(n_56151), .Z(n_137674244));
	notech_or4 i_51260067(.A(n_182758113), .B(n_56270), .C(n_317788512), .D(n_57351
		), .Z(n_138174249));
	notech_or2 i_50960070(.A(n_319288497), .B(n_27570), .Z(n_138474252));
	notech_or2 i_50660073(.A(n_318888501), .B(\nbus_11276[7] ), .Z(n_138774255
		));
	notech_nand3 i_60559986(.A(n_59193), .B(n_59940), .C(read_data[4]), .Z(n_139074258
		));
	notech_or4 i_59959989(.A(n_55820), .B(n_58483), .C(n_319588494), .D(n_60596
		), .Z(n_139374261));
	notech_or2 i_59659992(.A(n_55316), .B(nbus_11273[4]), .Z(n_139674264));
	notech_nao3 i_59359995(.A(n_2422), .B(n_55450), .C(n_54015), .Z(n_139974267
		));
	notech_or4 i_77459836(.A(n_55859), .B(n_57300), .C(n_204788866), .D(n_56163
		), .Z(n_140074268));
	notech_or2 i_76859841(.A(n_339176228), .B(\nbus_11276[8] ), .Z(n_140774275
		));
	notech_nor2 i_78159829(.A(n_55085), .B(n_56151), .Z(n_140874276));
	notech_or4 i_77559835(.A(n_2349), .B(n_264436799), .C(n_353069302), .D(n_177074638
		), .Z(n_141374281));
	notech_nao3 i_77659834(.A(opc_10[9]), .B(n_62401), .C(n_327576114), .Z(n_141474282
		));
	notech_or2 i_78959821(.A(n_2672), .B(nbus_11326[29]), .Z(n_141574283));
	notech_or2 i_78459826(.A(n_55068), .B(nbus_11273[29]), .Z(n_142274290)
		);
	notech_or4 i_79759813(.A(n_163674504), .B(n_161857906), .C(n_56449), .D(n_264436799
		), .Z(n_142374291));
	notech_or2 i_79259818(.A(n_57350), .B(n_54445), .Z(n_143074298));
	notech_or4 i_80059810(.A(n_60782), .B(n_60729), .C(n_1970), .D(n_29045),
		 .Z(n_143574303));
	notech_or2 i_82459786(.A(n_303521922), .B(nbus_11326[29]), .Z(n_143674304
		));
	notech_or2 i_81959791(.A(n_55070), .B(nbus_11273[29]), .Z(n_144374311)
		);
	notech_ao4 i_167259008(.A(n_55071), .B(\nbus_11276[29] ), .C(n_55872), .D
		(n_262936784), .Z(n_144474312));
	notech_ao4 i_167159009(.A(n_55397), .B(n_28977), .C(n_55396), .D(n_57329
		), .Z(n_144674314));
	notech_and3 i_167559006(.A(n_144474312), .B(n_144674314), .C(n_144374311
		), .Z(n_144774315));
	notech_ao4 i_166959011(.A(n_110923096), .B(n_306621953), .C(n_270688747)
		, .D(n_309921986), .Z(n_144874316));
	notech_ao4 i_165159028(.A(n_161957907), .B(n_325776096), .C(n_157974447)
		, .D(n_55872), .Z(n_145174319));
	notech_ao4 i_165059029(.A(nbus_11273[8]), .B(n_339576232), .C(n_54433), 
		.D(n_29045), .Z(n_145374321));
	notech_nand3 i_165359026(.A(n_145174319), .B(n_145374321), .C(n_143074298
		), .Z(n_145474322));
	notech_ao4 i_164859031(.A(n_339676233), .B(n_27571), .C(n_339476231), .D
		(\nbus_11276[8] ), .Z(n_145574323));
	notech_ao4 i_165559024(.A(n_2177), .B(n_57350), .C(n_27527), .D(n_59865)
		, .Z(n_145674324));
	notech_ao4 i_165459025(.A(n_254834174), .B(\nbus_11276[8] ), .C(n_2333),
		 .D(n_56703), .Z(n_145874326));
	notech_nand3 i_64460590(.A(n_145674324), .B(n_145874326), .C(n_143574303
		), .Z(n_145974327));
	notech_ao4 i_164459035(.A(n_55069), .B(\nbus_11276[29] ), .C(n_56151), .D
		(n_262936784), .Z(n_146274330));
	notech_ao4 i_164359036(.A(n_28977), .B(n_26444), .C(n_57329), .D(n_2655)
		, .Z(n_146474332));
	notech_and3 i_164659033(.A(n_146274330), .B(n_146474332), .C(n_142274290
		), .Z(n_146574333));
	notech_ao4 i_164159038(.A(n_110923096), .B(n_2694), .C(n_270688747), .D(n_2674
		), .Z(n_146674334));
	notech_ao4 i_163659043(.A(nbus_11273[9]), .B(n_164274510), .C(\nbus_11276[9] 
		), .D(n_164374511), .Z(n_147174339));
	notech_nand3 i_163859041(.A(n_141374281), .B(n_147174339), .C(n_141474282
		), .Z(n_147274340));
	notech_ao4 i_163459045(.A(n_57349), .B(n_2656), .C(n_2653), .D(n_29048),
		 .Z(n_147374341));
	notech_ao4 i_163059049(.A(n_161957907), .B(n_327576114), .C(n_161857906)
		, .D(n_327476113), .Z(n_147674344));
	notech_ao4 i_162959050(.A(n_339376230), .B(n_27571), .C(n_56703), .D(n_339276229
		), .Z(n_147874346));
	notech_ao4 i_162759052(.A(n_2656), .B(n_57350), .C(n_2653), .D(n_29045),
		 .Z(n_148074348));
	notech_and3 i_162859051(.A(n_140074268), .B(n_148074348), .C(n_26404), .Z
		(n_148274350));
	notech_ao4 i_143559229(.A(n_316288527), .B(n_261136766), .C(n_260436759)
		, .D(n_316388526), .Z(n_148474352));
	notech_ao4 i_143359231(.A(n_55304), .B(\nbus_11276[4] ), .C(n_53993), .D
		(n_29351), .Z(n_148674354));
	notech_and4 i_143759227(.A(n_148674354), .B(n_148474352), .C(n_139674264
		), .D(n_139974267), .Z(n_148874356));
	notech_ao4 i_143059234(.A(n_55422), .B(n_321188478), .C(n_55421), .D(n_29063
		), .Z(n_148974357));
	notech_ao4 i_142859236(.A(n_59193), .B(n_26743), .C(n_55951), .D(n_27565
		), .Z(n_149174359));
	notech_and4 i_143259232(.A(n_149174359), .B(n_139374261), .C(n_148974357
		), .D(n_139074258), .Z(n_149374361));
	notech_ao4 i_132059329(.A(n_320188488), .B(n_2679), .C(n_59193), .D(n_26723
		), .Z(n_149474362));
	notech_ao4 i_131859331(.A(n_320688483), .B(n_2680), .C(n_319088499), .D(nbus_11273
		[7]), .Z(n_149674364));
	notech_and4 i_132259327(.A(n_149674364), .B(n_149474362), .C(n_138474252
		), .D(n_138774255), .Z(n_149874366));
	notech_ao4 i_131559334(.A(n_28983), .B(n_55222), .C(n_55688), .D(n_2675)
		, .Z(n_149974367));
	notech_ao4 i_131359336(.A(n_321688474), .B(n_29350), .C(n_321788473), .D
		(n_29349), .Z(n_150174369));
	notech_and4 i_131459335(.A(n_150874376), .B(n_158074448), .C(n_150174369
		), .D(n_137474242), .Z(n_150274370));
	notech_and2 i_4957808(.A(n_35657), .B(n_55546), .Z(n_150574373));
	notech_and2 i_4157816(.A(n_249634122), .B(n_186374731), .Z(n_150674374)
		);
	notech_and4 i_83157083(.A(n_55667), .B(n_243864755), .C(n_258664903), .D
		(n_55974), .Z(n_150774375));
	notech_or2 i_85557060(.A(n_316688523), .B(nbus_11273[7]), .Z(n_150874376
		));
	notech_or4 i_90557011(.A(n_60752), .B(n_60739), .C(n_60782), .D(n_55546)
		, .Z(n_151174379));
	notech_or2 i_92556992(.A(n_55580), .B(n_55893), .Z(n_151274380));
	notech_nao3 i_56857314(.A(opc_10[4]), .B(n_62401), .C(n_259336748), .Z(n_151374381
		));
	notech_nand2 i_56257319(.A(n_55729), .B(opd[4]), .Z(n_152074388));
	notech_nao3 i_57757306(.A(opc_10[6]), .B(n_62431), .C(n_259336748), .Z(n_152374391
		));
	notech_nand2 i_57157311(.A(opd[6]), .B(n_55729), .Z(n_152874396));
	notech_nao3 i_58557298(.A(opc_10[7]), .B(n_62431), .C(n_259336748), .Z(n_152974397
		));
	notech_nand2 i_58057303(.A(opd[7]), .B(n_55729), .Z(n_153674404));
	notech_or4 i_60457282(.A(n_56240), .B(n_294061944), .C(n_55975), .D(n_57351
		), .Z(n_153774405));
	notech_or4 i_59957287(.A(n_274288715), .B(n_206288851), .C(n_55820), .D(n_2675
		), .Z(n_154474412));
	notech_or4 i_65257242(.A(n_56197), .B(n_273588720), .C(n_55820), .D(n_319588494
		), .Z(n_154974417));
	notech_nand2 i_64757247(.A(nAF), .B(n_208474952), .Z(n_155474422));
	notech_nand3 i_70257203(.A(n_273688719), .B(n_59940), .C(read_data[7]), 
		.Z(n_155774425));
	notech_or2 i_69757206(.A(n_55518), .B(n_57351), .Z(n_156074428));
	notech_nao3 i_69457209(.A(n_35829), .B(opa[15]), .C(n_252034146), .Z(n_156374431
		));
	notech_or4 i_68957212(.A(n_55522), .B(n_56449), .C(n_55961), .D(n_2679),
		 .Z(n_156674434));
	notech_nor2 i_21599(.A(n_217467994), .B(n_150574373), .Z(n_156774435));
	notech_or4 i_78957124(.A(n_59370), .B(n_2645), .C(n_59945), .D(nbus_11326
		[7]), .Z(n_156874436));
	notech_nand2 i_78857125(.A(n_55752), .B(opd[7]), .Z(n_157174439));
	notech_or4 i_78357130(.A(n_59259), .B(n_59273), .C(n_56197), .D(n_251734143
		), .Z(n_157674444));
	notech_or2 i_27449(.A(n_55859), .B(n_57300), .Z(n_157974447));
	notech_ao4 i_168556272(.A(n_57351), .B(n_316788522), .C(n_247634102), .D
		(n_60474), .Z(n_158074448));
	notech_ao4 i_159656361(.A(n_247334099), .B(n_2680), .C(n_247234098), .D(n_2679
		), .Z(n_158174449));
	notech_ao4 i_159556362(.A(n_54458), .B(n_57351), .C(n_54435), .D(n_28983
		), .Z(n_158374451));
	notech_ao4 i_159256365(.A(n_54565), .B(nbus_11273[7]), .C(n_54563), .D(\nbus_11276[7] 
		), .Z(n_158574453));
	notech_and4 i_159456363(.A(n_168964027), .B(n_158574453), .C(n_156874436
		), .D(n_157174439), .Z(n_158874456));
	notech_ao4 i_148256469(.A(n_249434120), .B(n_2680), .C(n_57326), .D(n_150674374
		), .Z(n_158974457));
	notech_ao4 i_148056471(.A(n_55873), .B(n_251734143), .C(n_249734123), .D
		(n_28983), .Z(n_159174459));
	notech_and4 i_148456467(.A(n_159174459), .B(n_156674434), .C(n_158974457
		), .D(n_156374431), .Z(n_159374461));
	notech_ao4 i_147756474(.A(n_55380), .B(\nbus_11276[7] ), .C(n_251934145)
		, .D(n_58951), .Z(n_159474462));
	notech_ao4 i_147556476(.A(n_54822), .B(n_26894), .C(n_55740), .D(n_27570
		), .Z(n_159674464));
	notech_and4 i_147956472(.A(n_159674464), .B(n_159474462), .C(n_155774425
		), .D(n_156074428), .Z(n_159874466));
	notech_ao4 i_145156498(.A(n_316288527), .B(n_249534121), .C(n_316388526)
		, .D(n_249434120), .Z(n_159974467));
	notech_ao4 i_145056499(.A(n_55355), .B(n_29063), .C(n_55270), .D(nbus_11273
		[4]), .Z(n_160174469));
	notech_and3 i_145356496(.A(n_159974467), .B(n_160174469), .C(n_155474422
		), .Z(n_160274470));
	notech_ao4 i_144756502(.A(n_55518), .B(n_321188478), .C(n_55380), .D(\nbus_11276[4] 
		), .Z(n_160374471));
	notech_ao4 i_144656503(.A(n_2193), .B(n_27523), .C(n_55740), .D(n_27565)
		, .Z(n_160574473));
	notech_ao4 i_141656533(.A(n_2680), .B(n_248734113), .C(n_248434110), .D(n_2679
		), .Z(n_160774475));
	notech_ao4 i_141556534(.A(n_54921), .B(n_57326), .C(n_54920), .D(n_55400
		), .Z(n_160974477));
	notech_ao4 i_141356536(.A(n_54748), .B(n_28983), .C(n_55730), .D(n_27570
		), .Z(n_161174479));
	notech_and4 i_141456535(.A(n_174064078), .B(n_173964077), .C(n_153774405
		), .D(n_161174479), .Z(n_161374481));
	notech_ao4 i_140256547(.A(n_55888), .B(n_251734143), .C(n_2680), .D(n_248634112
		), .Z(n_161474482));
	notech_ao4 i_140156548(.A(n_54749), .B(n_28983), .C(n_54922), .D(n_55400
		), .Z(n_161674484));
	notech_ao4 i_139956550(.A(n_54923), .B(n_57326), .C(n_54695), .D(n_57351
		), .Z(n_161874486));
	notech_and4 i_140056549(.A(n_174064078), .B(n_173964077), .C(n_161874486
		), .D(n_152974397), .Z(n_162074488));
	notech_ao4 i_139556554(.A(n_55888), .B(n_144377843), .C(n_248634112), .D
		(n_316488525), .Z(n_162174489));
	notech_ao4 i_139456555(.A(n_54749), .B(n_29068), .C(n_54922), .D(\nbus_11276[6] 
		), .Z(n_162374491));
	notech_ao4 i_139156558(.A(n_54923), .B(nbus_11273[6]), .C(n_54695), .D(n_57352
		), .Z(n_162574493));
	notech_and4 i_139356556(.A(n_53844), .B(n_162574493), .C(n_144277842), .D
		(n_152374391), .Z(n_162874496));
	notech_ao4 i_138556562(.A(n_55888), .B(n_139770716), .C(n_248634112), .D
		(n_316388526), .Z(n_162974497));
	notech_ao4 i_138456563(.A(n_54749), .B(n_29063), .C(n_54922), .D(\nbus_11276[4] 
		), .Z(n_163174499));
	notech_ao4 i_138256565(.A(n_54923), .B(nbus_11273[4]), .C(n_54695), .D(n_321188478
		), .Z(n_163374501));
	notech_and3 i_138356564(.A(n_137970698), .B(n_163374501), .C(n_151374381
		), .Z(n_163574503));
	notech_and4 i_155293(.A(n_55658), .B(n_56005), .C(n_55999), .D(n_135960441
		), .Z(n_163674504));
	notech_ao3 i_2955270(.A(n_54711), .B(n_29011), .C(n_163974507), .Z(n_163774505
		));
	notech_ao4 i_3055269(.A(n_55353), .B(n_56551), .C(n_55958), .D(n_54530),
		 .Z(n_163874506));
	notech_ao4 i_52254786(.A(n_55836), .B(n_26327), .C(n_56104), .D(n_35829)
		, .Z(n_163974507));
	notech_and3 i_194560627(.A(n_55068), .B(n_2677), .C(n_54468), .Z(n_164274510
		));
	notech_and3 i_194760626(.A(n_55069), .B(n_2678), .C(n_54428), .Z(n_164374511
		));
	notech_or2 i_120454141(.A(n_55872), .B(n_36952), .Z(n_165074518));
	notech_nand3 i_9955206(.A(n_54124), .B(tsc[24]), .C(n_59865), .Z(n_165174519
		));
	notech_or2 i_9855207(.A(n_351665805), .B(nbus_11326[24]), .Z(n_165474522
		));
	notech_or4 i_9355212(.A(n_58661), .B(n_56121), .C(n_56376), .D(n_27592),
		 .Z(n_165974527));
	notech_or2 i_25455051(.A(n_54853), .B(n_29037), .Z(n_166274530));
	notech_nao3 i_24955056(.A(n_62427), .B(opc[13]), .C(n_333569134), .Z(n_166774535
		));
	notech_or2 i_29655009(.A(n_262636781), .B(n_26943), .Z(n_167074538));
	notech_or4 i_29355012(.A(n_59168), .B(n_26604), .C(n_26377), .D(n_27529)
		, .Z(n_167374541));
	notech_or2 i_29055015(.A(n_55520), .B(n_29077), .Z(n_167674544));
	notech_nor2 i_39254913(.A(n_54872), .B(n_57345), .Z(n_168174549));
	notech_or4 i_38754918(.A(n_274288715), .B(n_206288851), .C(n_321831605),
		 .D(n_55859), .Z(n_168874556));
	notech_nand2 i_52154787(.A(nOF), .B(n_26580), .Z(n_169174559));
	notech_or2 i_51854790(.A(n_55727), .B(n_27576), .Z(n_169474562));
	notech_or4 i_51554793(.A(n_55252), .B(n_260988754), .C(n_260888755), .D(n_252034146
		), .Z(n_169774565));
	notech_nao3 i_53554773(.A(n_62433), .B(opc[13]), .C(n_248534111), .Z(n_171174579
		));
	notech_nao3 i_57254737(.A(n_2430), .B(n_55450), .C(n_54015), .Z(n_171474582
		));
	notech_or2 i_56954740(.A(n_55426), .B(n_57350), .Z(n_171774585));
	notech_nand2 i_56654743(.A(n_55728), .B(opd[8]), .Z(n_172074588));
	notech_or4 i_56354746(.A(n_206288851), .B(n_57300), .C(n_59250), .D(n_2240
		), .Z(n_172374591));
	notech_nao3 i_61454700(.A(n_2438), .B(n_55450), .C(n_54015), .Z(n_172674594
		));
	notech_or2 i_61054703(.A(n_57346), .B(n_55426), .Z(n_172974597));
	notech_nand2 i_60754706(.A(n_55728), .B(opd[12]), .Z(n_173274600));
	notech_or4 i_60454709(.A(n_59250), .B(n_206288851), .C(n_2240), .D(n_321931606
		), .Z(n_173574603));
	notech_nao3 i_64354676(.A(n_2444), .B(n_55450), .C(n_232761396), .Z(n_173874606
		));
	notech_or2 i_63854679(.A(n_356476400), .B(n_55426), .Z(n_174174609));
	notech_nand2 i_63454682(.A(n_55728), .B(opd[15]), .Z(n_174474612));
	notech_or4 i_63154685(.A(n_59250), .B(n_206288851), .C(n_2240), .D(n_57293
		), .Z(n_174774615));
	notech_nor2 i_75854565(.A(n_55424), .B(nbus_11326[24]), .Z(n_174874616)
		);
	notech_or4 i_75354570(.A(n_56197), .B(n_58660), .C(n_56376), .D(n_27592)
		, .Z(n_175574623));
	notech_or2 i_76554558(.A(n_54431), .B(n_29077), .Z(n_175674624));
	notech_or2 i_86754464(.A(n_2653), .B(n_29077), .Z(n_176374631));
	notech_and4 i_190160637(.A(n_56058), .B(n_2673), .C(n_1188), .D(n_1071),
		 .Z(n_177074638));
	notech_nor2 i_87554456(.A(n_2653), .B(n_29080), .Z(n_177174639));
	notech_ao3 i_87054461(.A(n_62427), .B(opc[11]), .C(n_327476113), .Z(n_177874646
		));
	notech_nor2 i_88354448(.A(n_2653), .B(n_29084), .Z(n_177974647));
	notech_ao3 i_87854453(.A(n_62409), .B(opc[12]), .C(n_327476113), .Z(n_178674654
		));
	notech_nor2 i_89154440(.A(n_2653), .B(n_29037), .Z(n_178774655));
	notech_ao3 i_88654445(.A(n_62433), .B(opc[13]), .C(n_327476113), .Z(n_179474662
		));
	notech_or2 i_89954432(.A(n_2653), .B(n_29087), .Z(n_179574663));
	notech_or4 i_89454437(.A(n_57293), .B(n_55859), .C(n_204788866), .D(n_274288715
		), .Z(n_180274670));
	notech_nor2 i_90754424(.A(n_2672), .B(nbus_11326[24]), .Z(n_180374671)
		);
	notech_or4 i_90254429(.A(n_204788866), .B(n_274288715), .C(n_56376), .D(n_27592
		), .Z(n_181074678));
	notech_nor2 i_93154400(.A(n_57347), .B(n_54445), .Z(n_181174679));
	notech_or4 i_92654405(.A(n_322031607), .B(n_55859), .C(n_56197), .D(n_274288715
		), .Z(n_181874686));
	notech_nor2 i_94854387(.A(n_57346), .B(n_54445), .Z(n_181974687));
	notech_or4 i_94154392(.A(n_56197), .B(n_274288715), .C(n_321931606), .D(n_55852
		), .Z(n_182674694));
	notech_or2 i_95154384(.A(n_254834174), .B(\nbus_11276[12] ), .Z(n_183174699
		));
	notech_nor2 i_96354374(.A(n_57345), .B(n_54445), .Z(n_183274700));
	notech_or4 i_95854379(.A(n_56196), .B(n_274288715), .C(n_321831605), .D(n_55852
		), .Z(n_183974707));
	notech_or2 i_96654371(.A(n_254834174), .B(\nbus_11276[13] ), .Z(n_184474712
		));
	notech_or4 i_97654361(.A(n_57293), .B(n_55852), .C(n_56196), .D(n_274288715
		), .Z(n_184574713));
	notech_or2 i_97154366(.A(n_339476231), .B(\nbus_11276[15] ), .Z(n_185274720
		));
	notech_nor2 i_98654353(.A(n_303521922), .B(nbus_11326[24]), .Z(n_185374721
		));
	notech_or4 i_97954358(.A(n_56196), .B(n_274288715), .C(n_56376), .D(n_27592
		), .Z(n_186074728));
	notech_or2 i_2855271(.A(opbs), .B(opas), .Z(n_186174729));
	notech_nand2 i_2755272(.A(opbs), .B(opas), .Z(n_186274730));
	notech_or2 i_21417(.A(n_252034146), .B(n_56104), .Z(n_186374731));
	notech_ao4 i_202753336(.A(n_322231609), .B(n_309921986), .C(n_251061538)
		, .D(n_306621953), .Z(n_186474732));
	notech_ao4 i_202653337(.A(n_57334), .B(n_55396), .C(n_29137), .D(n_55397
		), .Z(n_186674734));
	notech_nand3 i_202953334(.A(n_186074728), .B(n_186474732), .C(n_186674734
		), .Z(n_186774735));
	notech_ao4 i_202453339(.A(nbus_11273[24]), .B(n_55070), .C(n_55071), .D(\nbus_11276[24] 
		), .Z(n_186874736));
	notech_ao4 i_202053343(.A(n_177264110), .B(n_325776096), .C(n_177164109)
		, .D(n_325676095), .Z(n_187174739));
	notech_ao4 i_201953344(.A(n_339676233), .B(n_27581), .C(nbus_11273[15]),
		 .D(n_339576232), .Z(n_187374741));
	notech_and3 i_202253341(.A(n_187174739), .B(n_187374741), .C(n_185274720
		), .Z(n_187474742));
	notech_ao4 i_201753346(.A(n_356476400), .B(n_54445), .C(n_54433), .D(n_29087
		), .Z(n_187574743));
	notech_or2 i_64055302(.A(n_321831605), .B(n_55858), .Z(n_187874746));
	notech_ao4 i_201053353(.A(n_166457952), .B(n_325776096), .C(n_166557953)
		, .D(n_325676095), .Z(n_187974747));
	notech_ao4 i_200953354(.A(nbus_11273[13]), .B(n_339576232), .C(n_339476231
		), .D(\nbus_11276[13] ), .Z(n_188174749));
	notech_nand3 i_201253351(.A(n_183974707), .B(n_187974747), .C(n_188174749
		), .Z(n_188274750));
	notech_ao4 i_200753356(.A(n_54433), .B(n_29037), .C(n_27578), .D(n_339676233
		), .Z(n_188374751));
	notech_ao4 i_201453349(.A(n_2333), .B(nbus_11273[13]), .C(n_27532), .D(n_59865
		), .Z(n_188474752));
	notech_ao4 i_201353350(.A(n_2331), .B(n_29037), .C(n_57345), .D(n_2177),
		 .Z(n_188674754));
	notech_nand3 i_64755299(.A(n_188474752), .B(n_188674754), .C(n_184474712
		), .Z(n_188774755));
	notech_or2 i_63655304(.A(n_321931606), .B(n_55852), .Z(n_189074758));
	notech_ao4 i_200053363(.A(n_169057978), .B(n_325776096), .C(n_169157979)
		, .D(n_325676095), .Z(n_189174759));
	notech_ao4 i_199953364(.A(nbus_11273[12]), .B(n_339576232), .C(\nbus_11276[12] 
		), .D(n_339476231), .Z(n_189374761));
	notech_nand3 i_200253361(.A(n_182674694), .B(n_189174759), .C(n_189374761
		), .Z(n_189474762));
	notech_ao4 i_199753366(.A(n_54433), .B(n_29084), .C(n_339676233), .D(n_27577
		), .Z(n_189574763));
	notech_ao4 i_200453359(.A(nbus_11273[12]), .B(n_2333), .C(n_27531), .D(n_59863
		), .Z(n_189674764));
	notech_ao4 i_200353360(.A(n_2331), .B(n_29084), .C(n_57346), .D(n_2177),
		 .Z(n_189874766));
	notech_nand3 i_64655300(.A(n_189674764), .B(n_189874766), .C(n_183174699
		), .Z(n_189974767));
	notech_ao4 i_199053373(.A(n_171658004), .B(n_325776096), .C(n_171758005)
		, .D(n_325676095), .Z(n_190274770));
	notech_ao4 i_198953374(.A(n_56730), .B(n_339576232), .C(n_339476231), .D
		(\nbus_11276[11] ), .Z(n_190474772));
	notech_nand3 i_199253371(.A(n_181874686), .B(n_190274770), .C(n_190474772
		), .Z(n_190574773));
	notech_ao4 i_198753376(.A(n_54433), .B(n_29080), .C(n_339676233), .D(n_27576
		), .Z(n_190674774));
	notech_ao4 i_197353390(.A(n_322231609), .B(n_2674), .C(n_251061538), .D(n_2694
		), .Z(n_190974777));
	notech_ao4 i_197253391(.A(n_57334), .B(n_2655), .C(n_29137), .D(n_26444)
		, .Z(n_191174779));
	notech_nand3 i_197553388(.A(n_181074678), .B(n_190974777), .C(n_191174779
		), .Z(n_191274780));
	notech_ao4 i_197053393(.A(n_55068), .B(nbus_11273[24]), .C(n_55069), .D(\nbus_11276[24] 
		), .Z(n_191374781));
	notech_ao4 i_196653397(.A(n_177164109), .B(n_327476113), .C(n_177264110)
		, .D(n_327576114), .Z(n_191674784));
	notech_ao4 i_196553398(.A(nbus_11273[15]), .B(n_339276229), .C(n_339376230
		), .D(n_27581), .Z(n_191874786));
	notech_and3 i_196853395(.A(n_180274670), .B(n_191674784), .C(n_191874786
		), .Z(n_191974787));
	notech_ao4 i_196353400(.A(n_356476400), .B(n_2656), .C(n_339176228), .D(\nbus_11276[15] 
		), .Z(n_192074788));
	notech_ao4 i_195953404(.A(n_166457952), .B(n_327576114), .C(n_56151), .D
		(n_187874746), .Z(n_192374791));
	notech_ao4 i_195753405(.A(nbus_11273[13]), .B(n_339276229), .C(n_27578),
		 .D(n_339376230), .Z(n_192574793));
	notech_nao3 i_196153402(.A(n_192374791), .B(n_192574793), .C(n_179474662
		), .Z(n_192674794));
	notech_ao4 i_195553407(.A(n_57345), .B(n_2656), .C(n_339176228), .D(\nbus_11276[13] 
		), .Z(n_192774795));
	notech_ao4 i_195153411(.A(n_169057978), .B(n_327576114), .C(n_56151), .D
		(n_189074758), .Z(n_193074798));
	notech_ao4 i_195053412(.A(n_56739), .B(n_339276229), .C(n_339376230), .D
		(n_27577), .Z(n_193274800));
	notech_nao3 i_195353409(.A(n_193074798), .B(n_193274800), .C(n_178674654
		), .Z(n_193374801));
	notech_ao4 i_194853414(.A(n_57346), .B(n_2656), .C(n_339176228), .D(\nbus_11276[12] 
		), .Z(n_193474802));
	notech_ao4 i_194453418(.A(n_171658004), .B(n_327576114), .C(n_238768192)
		, .D(n_56139), .Z(n_193774805));
	notech_ao4 i_194353419(.A(n_56730), .B(n_339276229), .C(n_339376230), .D
		(n_27576), .Z(n_193974807));
	notech_nao3 i_194653416(.A(n_193774805), .B(n_193974807), .C(n_177874646
		), .Z(n_194074808));
	notech_ao4 i_194153421(.A(n_57347), .B(n_2656), .C(n_339176228), .D(n_55469
		), .Z(n_194174809));
	notech_or4 i_193953423(.A(n_56465), .B(n_56431), .C(n_177074638), .D(n_29010
		), .Z(n_194474812));
	notech_ao4 i_193753425(.A(n_319431581), .B(n_56139), .C(n_174358031), .D
		(n_194474812), .Z(n_194574813));
	notech_ao4 i_193653426(.A(n_164274510), .B(nbus_11273[10]), .C(n_174258030
		), .D(n_327576114), .Z(n_194674814));
	notech_ao4 i_193453428(.A(n_57348), .B(n_2656), .C(n_164374511), .D(\nbus_11276[10] 
		), .Z(n_194874816));
	notech_and3 i_193553427(.A(n_154070859), .B(n_194874816), .C(n_176374631
		), .Z(n_195074818));
	notech_or4 i_185253507(.A(n_56465), .B(n_355988238), .C(n_54594), .D(n_29010
		), .Z(n_195174819));
	notech_ao4 i_185053509(.A(n_319431581), .B(n_56043), .C(n_174358031), .D
		(n_195174819), .Z(n_195274820));
	notech_ao4 i_184953510(.A(n_54562), .B(nbus_11273[10]), .C(n_364788148),
		 .D(n_174258030), .Z(n_195374821));
	notech_ao4 i_184753512(.A(n_54455), .B(n_57348), .C(\nbus_11276[10] ), .D
		(n_54547), .Z(n_195574823));
	notech_and3 i_184853511(.A(n_154070859), .B(n_195574823), .C(n_175674624
		), .Z(n_195774825));
	notech_ao4 i_184353516(.A(n_322231609), .B(n_309618873), .C(n_251061538)
		, .D(n_308418861), .Z(n_195874826));
	notech_ao4 i_184253517(.A(n_55404), .B(n_57334), .C(n_29137), .D(n_55405
		), .Z(n_196074828));
	notech_nand3 i_184553514(.A(n_175574623), .B(n_195874826), .C(n_196074828
		), .Z(n_196174829));
	notech_ao4 i_184053519(.A(n_55064), .B(nbus_11273[24]), .C(n_55062), .D(\nbus_11276[24] 
		), .Z(n_196274830));
	notech_ao4 i_174353615(.A(n_177164109), .B(n_354188267), .C(n_177264110)
		, .D(n_354088268), .Z(n_196574833));
	notech_ao4 i_174153617(.A(n_59168), .B(n_27534), .C(n_59193), .D(n_26757
		), .Z(n_196774835));
	notech_and4 i_174553613(.A(n_196774835), .B(n_174774615), .C(n_196574833
		), .D(n_174474612), .Z(n_196974837));
	notech_ao4 i_173853620(.A(n_55308), .B(\nbus_11276[15] ), .C(n_55307), .D
		(n_56766), .Z(n_197074838));
	notech_ao4 i_173653622(.A(n_53993), .B(n_29356), .C(n_55427), .D(n_29087
		), .Z(n_197274840));
	notech_and4 i_174053618(.A(n_197274840), .B(n_197074838), .C(n_173874606
		), .D(n_174174609), .Z(n_197474842));
	notech_ao4 i_172353635(.A(n_169157979), .B(n_354188267), .C(n_169057978)
		, .D(n_354088268), .Z(n_197574843));
	notech_ao4 i_172153637(.A(n_59163), .B(n_27531), .C(n_59193), .D(n_26753
		), .Z(n_197774845));
	notech_and4 i_172553633(.A(n_197774845), .B(n_173574603), .C(n_197574843
		), .D(n_173274600), .Z(n_197974847));
	notech_ao4 i_171853640(.A(n_55308), .B(n_55542), .C(n_55307), .D(n_56739
		), .Z(n_198074848));
	notech_ao4 i_171653642(.A(n_53993), .B(n_29355), .C(n_55427), .D(n_29084
		), .Z(n_198274850));
	notech_and4 i_172053638(.A(n_198274850), .B(n_198074848), .C(n_172674594
		), .D(n_172974597), .Z(n_198474852));
	notech_ao4 i_169053668(.A(n_161857906), .B(n_354188267), .C(n_161957907)
		, .D(n_354088268), .Z(n_198574853));
	notech_ao4 i_168853670(.A(n_59159), .B(n_27527), .C(n_59193), .D(n_26748
		), .Z(n_198774855));
	notech_and4 i_169253666(.A(n_198774855), .B(n_172374591), .C(n_198574853
		), .D(n_172074588), .Z(n_198974857));
	notech_ao4 i_168553673(.A(n_55308), .B(\nbus_11276[8] ), .C(n_55307), .D
		(n_56703), .Z(n_199074858));
	notech_ao4 i_168353675(.A(n_53993), .B(n_29354), .C(n_55427), .D(n_29045
		), .Z(n_199274860));
	notech_and4 i_168753671(.A(n_199274860), .B(n_199074858), .C(n_171474582
		), .D(n_171774585), .Z(n_199474862));
	notech_ao4 i_166653692(.A(n_166457952), .B(n_2326), .C(n_55873), .D(n_187874746
		), .Z(n_199574863));
	notech_ao4 i_166553693(.A(n_55727), .B(n_27578), .C(n_2193), .D(n_27532)
		, .Z(n_199774865));
	notech_and3 i_166853690(.A(n_199574863), .B(n_199774865), .C(n_171174579
		), .Z(n_199874866));
	notech_ao4 i_166353695(.A(n_55310), .B(n_55552), .C(n_26548), .D(n_56748
		), .Z(n_199974867));
	notech_ao4 i_166253696(.A(n_55354), .B(n_29037), .C(n_55156), .D(n_57345
		), .Z(n_200074868));
	notech_ao4 i_165153707(.A(n_163874506), .B(n_29080), .C(n_56730), .D(n_163774505
		), .Z(n_200374871));
	notech_ao4 i_165053708(.A(n_171658004), .B(n_2326), .C(n_238768192), .D(n_55873
		), .Z(n_200474872));
	notech_ao4 i_164853710(.A(n_55253), .B(n_251834144), .C(n_171758005), .D
		(n_248534111), .Z(n_200674874));
	notech_and4 i_165353705(.A(n_200674874), .B(n_200474872), .C(n_200374871
		), .D(n_169774565), .Z(n_200874876));
	notech_ao4 i_164553713(.A(n_27530), .B(n_2193), .C(n_55282), .D(n_186374731
		), .Z(n_200974877));
	notech_ao4 i_164353715(.A(n_57347), .B(n_55156), .C(n_55469), .D(n_55310
		), .Z(n_201174879));
	notech_and4 i_164753711(.A(n_201174879), .B(n_200974877), .C(n_169174559
		), .D(n_169474562), .Z(n_201374881));
	notech_ao4 i_154553812(.A(n_318231569), .B(n_166557953), .C(n_318031567)
		, .D(n_166457952), .Z(n_201474882));
	notech_ao4 i_154453813(.A(n_54944), .B(n_56748), .C(n_54943), .D(n_55552
		), .Z(n_201674884));
	notech_nand3 i_154853810(.A(n_168874556), .B(n_201474882), .C(n_201674884
		), .Z(n_201774885));
	notech_ao4 i_154253815(.A(n_54902), .B(n_29037), .C(n_55726), .D(n_27578
		), .Z(n_201874886));
	notech_ao4 i_146153894(.A(n_174358031), .B(n_320565522), .C(n_174258030)
		, .D(n_320665523), .Z(n_202174889));
	notech_ao4 i_146053895(.A(n_55381), .B(\nbus_11276[10] ), .C(n_322131608
		), .D(n_320465521), .Z(n_202274890));
	notech_ao4 i_145853897(.A(n_55519), .B(n_57348), .C(n_55382), .D(n_56721
		), .Z(n_202474892));
	notech_and4 i_146353892(.A(n_202474892), .B(n_202274890), .C(n_202174889
		), .D(n_167674544), .Z(n_202674894));
	notech_ao4 i_145553900(.A(n_59193), .B(n_26695), .C(n_55738), .D(n_27575
		), .Z(n_202774895));
	notech_ao4 i_145353902(.A(n_55977), .B(n_28424), .C(n_56024), .D(n_29352
		), .Z(n_202974897));
	notech_and4 i_145753898(.A(n_202974897), .B(n_202774895), .C(n_167074538
		), .D(n_167374541), .Z(n_203174899));
	notech_ao4 i_141753931(.A(n_166457952), .B(n_333669135), .C(n_55888), .D
		(n_187874746), .Z(n_203274900));
	notech_ao4 i_141653932(.A(n_56748), .B(n_54946), .C(n_27578), .D(n_55725
		), .Z(n_203474902));
	notech_ao4 i_141353935(.A(n_57345), .B(n_54852), .C(n_54945), .D(n_55552
		), .Z(n_203674904));
	notech_and4 i_141553933(.A(n_53844), .B(n_203674904), .C(n_166274530), .D
		(n_26408), .Z(n_203974907));
	notech_ao4 i_126954077(.A(n_322231609), .B(n_352265811), .C(n_251061538)
		, .D(n_352865817), .Z(n_204074908));
	notech_ao4 i_126854078(.A(n_57334), .B(n_351865807), .C(n_29137), .D(n_351765806
		), .Z(n_204274910));
	notech_ao4 i_126554081(.A(n_55143), .B(nbus_11273[24]), .C(n_55142), .D(\nbus_11276[24] 
		), .Z(n_204474912));
	notech_and4 i_126754079(.A(n_204474912), .B(n_26375), .C(n_165174519), .D
		(n_165474522), .Z(n_204774915));
	notech_and3 i_22729(.A(n_55658), .B(n_238758633), .C(n_322288468), .Z(n_34533
		));
	notech_nand2 i_25651721(.A(n_323488456), .B(n_26516), .Z(n_204874916));
	notech_or2 i_26251715(.A(n_55580), .B(n_56043), .Z(n_204974917));
	notech_or4 i_87351145(.A(n_56196), .B(n_274288715), .C(n_2688), .D(n_55820
		), .Z(n_205074918));
	notech_or2 i_87051148(.A(n_55756), .B(n_27561), .Z(n_205574923));
	notech_nao3 i_87151147(.A(n_62409), .B(opc[0]), .C(n_279739585), .Z(n_205674924
		));
	notech_nao3 i_87251146(.A(opc_10[0]), .B(n_62431), .C(n_275539543), .Z(n_205774925
		));
	notech_and4 i_120652(.A(n_205774925), .B(n_41726130), .C(n_209174959), .D
		(n_205074918), .Z(n_19785));
	notech_and3 i_185452042(.A(n_322088470), .B(n_54455), .C(n_204874916), .Z
		(n_54631));
	notech_nand3 i_181852041(.A(n_97522962), .B(n_54431), .C(n_355976395), .Z
		(n_54661));
	notech_and2 i_59652040(.A(n_353465823), .B(n_204974917), .Z(n_55753));
	notech_or4 i_105050975(.A(n_204788866), .B(n_56074), .C(n_2688), .D(n_55820
		), .Z(n_205874926));
	notech_nand2 i_104450981(.A(n_54661), .B(opa[0]), .Z(n_206374931));
	notech_nao3 i_104850977(.A(n_62433), .B(opc[0]), .C(n_356276398), .Z(n_206474932
		));
	notech_nao3 i_104950976(.A(opc_10[0]), .B(n_62431), .C(n_356376399), .Z(n_206574933
		));
	notech_and4 i_120940(.A(n_41726130), .B(n_209874966), .C(n_205874926), .D
		(n_206574933), .Z(n_8979));
	notech_nand3 i_114150887(.A(n_273688719), .B(n_59945), .C(read_data[0]),
		 .Z(n_207274940));
	notech_ao3 i_114350885(.A(n_62409), .B(opc[0]), .C(n_249434120), .Z(n_207374941
		));
	notech_nao3 i_121292(.A(n_210674974), .B(n_210974976), .C(n_207374941), 
		.Z(n_20601));
	notech_or4 i_129950739(.A(n_56074), .B(n_206288851), .C(n_2688), .D(n_55820
		), .Z(n_207674944));
	notech_nao3 i_129750741(.A(n_62423), .B(opc[0]), .C(n_248634112), .Z(n_208274950
		));
	notech_nao3 i_129850740(.A(opc_10[0]), .B(n_62431), .C(n_259336748), .Z(n_208374951
		));
	notech_and4 i_121836(.A(n_211574982), .B(n_207674944), .C(n_208374951), 
		.D(n_41726130), .Z(n_12401));
	notech_nand2 i_138957960(.A(n_54822), .B(n_151174379), .Z(n_208474952)
		);
	notech_ao4 i_87551143(.A(n_54655), .B(\nbus_11276[0] ), .C(n_54656), .D(nbus_11273
		[0]), .Z(n_208774955));
	notech_ao4 i_87451144(.A(n_54438), .B(n_28986), .C(n_2699), .D(n_54469),
		 .Z(n_208874956));
	notech_and4 i_87851140(.A(n_208874956), .B(n_208774955), .C(n_205574923)
		, .D(n_205674924), .Z(n_209174959));
	notech_ao4 i_105150974(.A(n_356176397), .B(n_28986), .C(n_356076396), .D
		(n_2699), .Z(n_209474962));
	notech_ao4 i_105250973(.A(n_55753), .B(n_27561), .C(n_54631), .D(\nbus_11276[0] 
		), .Z(n_209574963));
	notech_and4 i_105550970(.A(n_209574963), .B(n_209474962), .C(n_206374931
		), .D(n_206474932), .Z(n_209874966));
	notech_ao4 i_114550883(.A(n_55518), .B(n_2699), .C(n_26341), .D(n_26891)
		, .Z(n_210174969));
	notech_ao4 i_114650882(.A(n_55270), .B(nbus_11273[0]), .C(n_55355), .D(n_28986
		), .Z(n_210374971));
	notech_ao4 i_114750881(.A(n_55740), .B(n_27561), .C(n_55380), .D(\nbus_11276[0] 
		), .Z(n_210474972));
	notech_and4 i_115150878(.A(n_210474972), .B(n_210374971), .C(n_210174969
		), .D(n_207274940), .Z(n_210674974));
	notech_ao4 i_115350876(.A(n_43626149), .B(n_249534121), .C(n_55685), .D(n_2688
		), .Z(n_210974976));
	notech_ao4 i_130350736(.A(n_55342), .B(n_26405), .C(n_54922), .D(\nbus_11276[0] 
		), .Z(n_211074977));
	notech_ao4 i_130150738(.A(n_54695), .B(n_2699), .C(n_1031), .D(n_59945),
		 .Z(n_211174978));
	notech_ao4 i_130250737(.A(n_54923), .B(nbus_11273[0]), .C(n_54749), .D(n_28986
		), .Z(n_211274979));
	notech_and4 i_130650733(.A(n_211274979), .B(n_211174978), .C(n_211074977
		), .D(n_208274950), .Z(n_211574982));
	notech_or2 i_45848722(.A(n_55070), .B(n_56901), .Z(n_212274989));
	notech_nao3 i_46148719(.A(opc_10[30]), .B(n_62417), .C(n_306621953), .Z(n_212374990
		));
	notech_or4 i_46048720(.A(n_56196), .B(n_274288715), .C(n_54367), .D(n_271188744
		), .Z(n_212474991));
	notech_or2 i_45948721(.A(n_55396), .B(n_270988746), .Z(n_212574992));
	notech_and4 i_3120682(.A(n_228075137), .B(n_101523002), .C(n_212474991),
		 .D(n_212574992), .Z(n_19965));
	notech_or4 i_58148608(.A(n_204788866), .B(n_56074), .C(n_54367), .D(n_270688747
		), .Z(n_212674993));
	notech_or2 i_57548614(.A(n_121623203), .B(nbus_11326[29]), .Z(n_212774994
		));
	notech_or2 i_58048609(.A(n_97522962), .B(n_56892), .Z(n_213274999));
	notech_nao3 i_58248607(.A(opc_10[29]), .B(n_62417), .C(n_121723204), .Z(n_213375000
		));
	notech_nand3 i_3020969(.A(n_228875145), .B(n_213375000), .C(n_212674993)
		, .Z(n_9153));
	notech_nor2 i_76748429(.A(n_354969318), .B(n_271088745), .Z(n_213475001)
		);
	notech_or2 i_76448432(.A(n_55562), .B(n_58951), .Z(n_213775004));
	notech_nor2 i_76548431(.A(n_354669316), .B(n_56943), .Z(n_213875005));
	notech_and2 i_76648430(.A(n_354869317), .B(\regs_13_14[31] ), .Z(n_213975006
		));
	notech_nor2 i_77048426(.A(n_113313527), .B(nbus_11326[31]), .Z(n_214075007
		));
	notech_ao3 i_76948427(.A(opc_10[31]), .B(n_62417), .C(n_113113525), .Z(n_214175008
		));
	notech_nor2 i_76848428(.A(n_354569315), .B(n_271288743), .Z(n_214275009)
		);
	notech_or4 i_3221323(.A(n_214175008), .B(n_229475151), .C(n_214275009), 
		.D(n_213475001), .Z(n_20787));
	notech_nor2 i_78648412(.A(n_270988746), .B(n_354969318), .Z(n_214475010)
		);
	notech_or2 i_78248415(.A(n_55562), .B(n_56901), .Z(n_214775013));
	notech_nor2 i_78348414(.A(n_354669316), .B(\nbus_11276[30] ), .Z(n_214875014
		));
	notech_and2 i_78448413(.A(\regs_13_14[30] ), .B(n_354869317), .Z(n_214975015
		));
	notech_nor2 i_79248409(.A(n_113313527), .B(nbus_11326[30]), .Z(n_215075016
		));
	notech_ao3 i_78848410(.A(opc_10[30]), .B(n_62417), .C(n_113113525), .Z(n_215175017
		));
	notech_nor2 i_78748411(.A(n_271188744), .B(n_354569315), .Z(n_215275018)
		);
	notech_or4 i_3121322(.A(n_215175017), .B(n_230175158), .C(n_215275018), 
		.D(n_214475010), .Z(n_20781));
	notech_or2 i_90948302(.A(n_55219), .B(n_56901), .Z(n_215875023));
	notech_nao3 i_91248299(.A(opc_10[30]), .B(n_62417), .C(n_308718864), .Z(n_215975024
		));
	notech_or4 i_91148300(.A(n_274288715), .B(n_206288851), .C(n_55523), .D(n_271188744
		), .Z(n_216075025));
	notech_or2 i_91048301(.A(n_55554), .B(n_270988746), .Z(n_216175026));
	notech_and4 i_3121610(.A(n_230875165), .B(n_101523002), .C(n_216075025),
		 .D(n_216175026), .Z(n_13295));
	notech_or4 i_92848284(.A(n_274288715), .B(n_206288851), .C(n_54367), .D(n_270688747
		), .Z(n_216275027));
	notech_or2 i_92248290(.A(n_308318860), .B(n_59104), .Z(n_216375028));
	notech_or2 i_92748285(.A(n_55219), .B(n_56892), .Z(n_216875033));
	notech_nao3 i_92948283(.A(opc_10[29]), .B(n_62417), .C(n_263575474), .Z(n_216975034
		));
	notech_nand3 i_3021609(.A(n_231675173), .B(n_216275027), .C(n_216975034)
		, .Z(n_13289));
	notech_or4 i_139047846(.A(n_244656264), .B(n_1844), .C(n_59945), .D(nbus_11326
		[26]), .Z(n_217075035));
	notech_nand3 i_2716836(.A(n_231975176), .B(n_231875175), .C(n_232575182)
		, .Z(n_9837));
	notech_or4 i_142847810(.A(n_244656264), .B(n_1844), .C(n_59945), .D(nbus_11326
		[24]), .Z(n_218175044));
	notech_nand3 i_2516834(.A(n_232875184), .B(n_232775183), .C(n_233675190)
		, .Z(n_9827));
	notech_or4 i_172447528(.A(n_57445), .B(n_59863), .C(n_2792), .D(n_27549)
		, .Z(n_219275053));
	notech_nand2 i_173647517(.A(\opc_5[10] ), .B(n_26596), .Z(n_220375064)
		);
	notech_nand3 i_1116820(.A(n_233775191), .B(n_234775201), .C(n_233975193)
		, .Z(n_9757));
	notech_or4 i_177547480(.A(n_57445), .B(n_59863), .C(n_2792), .D(n_27546)
		, .Z(n_220475065));
	notech_nand2 i_178647469(.A(\opc_5[8] ), .B(n_26596), .Z(n_221575076));
	notech_nand3 i_916818(.A(n_234875202), .B(n_235975212), .C(n_235075204),
		 .Z(n_9747));
	notech_nand2 i_184547410(.A(n_149823485), .B(n_321888472), .Z(n_221675077
		));
	notech_ao3 i_2849131(.A(n_321988471), .B(n_208358369), .C(n_208258368), 
		.Z(n_221875079));
	notech_nao3 i_2749132(.A(n_236175214), .B(n_236375216), .C(n_26343), .Z(n_222575085
		));
	notech_nor2 i_186747388(.A(opc[3]), .B(n_222775087), .Z(n_222675086));
	notech_ao4 i_2649133(.A(n_236075213), .B(opc[2]), .C(n_21822205), .D(n_2708
		), .Z(n_222775087));
	notech_or2 i_185447401(.A(n_54735), .B(n_55469), .Z(n_222875088));
	notech_nao3 i_186347392(.A(mul64[35]), .B(n_59863), .C(n_55389), .Z(n_223775097
		));
	notech_nao3 i_186547390(.A(\opc_1[3] ), .B(n_26596), .C(n_213758422), .Z
		(n_223875098));
	notech_and3 i_186447391(.A(rep_en3), .B(n_213458419), .C(n_4728), .Z(n_223975099
		));
	notech_and2 i_186647389(.A(opc[3]), .B(n_222575085), .Z(n_224075100));
	notech_or4 i_416813(.A(n_223975099), .B(n_224075100), .C(n_222675086), .D
		(n_26344), .Z(n_9722));
	notech_nao3 i_188447373(.A(opc[1]), .B(opc[0]), .C(n_21822205), .Z(n_224175101
		));
	notech_nor2 i_189847359(.A(opc[2]), .B(n_224375103), .Z(n_224275102));
	notech_and2 i_2949130(.A(n_236075213), .B(n_224175101), .Z(n_224375103)
		);
	notech_or2 i_188547372(.A(n_54735), .B(n_55438), .Z(n_224475104));
	notech_nao3 i_189447363(.A(mul64[34]), .B(n_59863), .C(n_55389), .Z(n_225375113
		));
	notech_nao3 i_189747360(.A(\opc_1[2] ), .B(n_26596), .C(n_213758422), .Z
		(n_225475114));
	notech_and3 i_189547362(.A(rep_en3), .B(n_213458419), .C(n_4727), .Z(n_225575115
		));
	notech_and2 i_189647361(.A(opc[2]), .B(n_236275215), .Z(n_225675116));
	notech_or4 i_316812(.A(n_225575115), .B(n_225675116), .C(n_224275102), .D
		(n_26345), .Z(n_9717));
	notech_nor2 i_195847299(.A(opc[0]), .B(n_225875118), .Z(n_225775117));
	notech_ao3 i_3549126(.A(n_21822205), .B(n_208358369), .C(n_208258368), .Z
		(n_225875118));
	notech_nand2 i_3449127(.A(n_54884), .B(n_321988471), .Z(n_225975119));
	notech_or2 i_194647311(.A(n_54735), .B(n_55413), .Z(n_226075120));
	notech_nao3 i_195547302(.A(mul64[32]), .B(n_59863), .C(n_55389), .Z(n_227275129
		));
	notech_nao3 i_195747300(.A(\opc_1[0] ), .B(n_26596), .C(n_213758422), .Z
		(n_227375130));
	notech_and2 i_195947298(.A(n_225975119), .B(opc[0]), .Z(n_227475131));
	notech_and3 i_195647301(.A(rep_en3), .B(n_4725), .C(n_213458419), .Z(n_227575132
		));
	notech_or4 i_116810(.A(n_227475131), .B(n_227575132), .C(n_225775117), .D
		(n_26346), .Z(n_9707));
	notech_ao4 i_46348717(.A(n_55719), .B(n_27599), .C(n_55397), .D(n_28997)
		, .Z(n_227675133));
	notech_ao4 i_46248718(.A(n_55071), .B(n_55234), .C(n_303521922), .D(nbus_11326
		[30]), .Z(n_227775134));
	notech_and4 i_46648714(.A(n_227775134), .B(n_227675133), .C(n_212274989)
		, .D(n_212374990), .Z(n_228075137));
	notech_and2 i_58348606(.A(n_262736782), .B(n_212774994), .Z(n_228375140)
		);
	notech_ao4 i_58448605(.A(n_57329), .B(n_55402), .C(n_322088470), .D(\nbus_11276[29] 
		), .Z(n_228575142));
	notech_ao4 i_58548604(.A(n_262936784), .B(n_56043), .C(n_55403), .D(n_28977
		), .Z(n_228675143));
	notech_and4 i_58948601(.A(n_228675143), .B(n_228575142), .C(n_213274999)
		, .D(n_228375140), .Z(n_228875145));
	notech_ao4 i_77148425(.A(n_55776), .B(n_27601), .C(n_2193), .D(n_27554),
		 .Z(n_229075147));
	notech_nand2 i_77248424(.A(n_229075147), .B(n_213775004), .Z(n_229175148
		));
	notech_or4 i_77548421(.A(n_213875005), .B(n_229175148), .C(n_213975006),
		 .D(n_214075007), .Z(n_229475151));
	notech_ao4 i_79348408(.A(n_55776), .B(n_27599), .C(n_2193), .D(n_27553),
		 .Z(n_229775154));
	notech_nand2 i_79448407(.A(n_229775154), .B(n_214775013), .Z(n_229875155
		));
	notech_or4 i_79748404(.A(n_214875014), .B(n_229875155), .C(n_214975015),
		 .D(n_215075016), .Z(n_230175158));
	notech_ao4 i_91448297(.A(n_55773), .B(n_27599), .C(n_55555), .D(n_28997)
		, .Z(n_230475161));
	notech_ao4 i_91348298(.A(n_55218), .B(n_55234), .C(n_308318860), .D(nbus_11326
		[30]), .Z(n_230575162));
	notech_and4 i_91748294(.A(n_230575162), .B(n_230475161), .C(n_215875023)
		, .D(n_215975024), .Z(n_230875165));
	notech_and2 i_93048282(.A(n_262736782), .B(n_216375028), .Z(n_231175168)
		);
	notech_ao4 i_93148281(.A(n_240675259), .B(n_57329), .C(n_55218), .D(n_55249
		), .Z(n_231375170));
	notech_ao4 i_93248280(.A(n_262936784), .B(n_55864), .C(n_240575258), .D(n_28977
		), .Z(n_231475171));
	notech_and4 i_93548277(.A(n_231475171), .B(n_231375170), .C(n_216875033)
		, .D(n_231175168), .Z(n_231675173));
	notech_ao4 i_140147835(.A(n_2247), .B(n_29357), .C(n_2313), .D(n_28926),
		 .Z(n_231875175));
	notech_ao4 i_140247834(.A(n_329546800), .B(n_29358), .C(n_2248), .D(nbus_11348
		[26]), .Z(n_231975176));
	notech_ao4 i_140347833(.A(n_231547139), .B(nbus_11326[2]), .C(n_2249), .D
		(n_29359), .Z(n_232175178));
	notech_ao4 i_140047836(.A(n_2314), .B(\nbus_11276[26] ), .C(n_55009), .D
		(n_28077), .Z(n_232375180));
	notech_and4 i_140747830(.A(n_2312), .B(n_232375180), .C(n_232175178), .D
		(n_217075035), .Z(n_232575182));
	notech_ao4 i_143947799(.A(n_2313), .B(n_28924), .C(n_2314), .D(\nbus_11276[24] 
		), .Z(n_232775183));
	notech_ao4 i_144047798(.A(n_2248), .B(nbus_11348[24]), .C(n_2247), .D(n_29360
		), .Z(n_232875184));
	notech_ao4 i_144147797(.A(n_2249), .B(n_29362), .C(n_329546800), .D(n_29361
		), .Z(n_233075186));
	notech_ao4 i_143847800(.A(n_231547139), .B(nbus_11326[0]), .C(n_55009), 
		.D(n_28075), .Z(n_233475188));
	notech_and4 i_144447794(.A(n_2312), .B(n_233475188), .C(n_233075186), .D
		(n_218175044), .Z(n_233675190));
	notech_ao4 i_174347511(.A(n_329546800), .B(n_29364), .C(n_2248), .D(nbus_11348
		[10]), .Z(n_233775191));
	notech_and4 i_174447510(.A(n_57312), .B(n_2186), .C(n_219275053), .D(n_220375064
		), .Z(n_233975193));
	notech_ao4 i_173947515(.A(n_54735), .B(nbus_11326[26]), .C(n_2311), .D(n_29339
		), .Z(n_234175195));
	notech_ao4 i_174047514(.A(n_55009), .B(n_28061), .C(n_54884), .D(n_55289
		), .Z(n_234275196));
	notech_ao4 i_174147513(.A(n_2314), .B(n_55438), .C(n_231547139), .D(nbus_11326
		[18]), .Z(n_234475198));
	notech_ao4 i_174247512(.A(n_2247), .B(n_29363), .C(n_2313), .D(n_28910),
		 .Z(n_234575199));
	notech_and4 i_174847506(.A(n_234575199), .B(n_234475198), .C(n_234275196
		), .D(n_234175195), .Z(n_234775201));
	notech_ao4 i_179247463(.A(n_329546800), .B(n_29368), .C(n_2248), .D(nbus_11348
		[8]), .Z(n_234875202));
	notech_and4 i_179347462(.A(n_57312), .B(n_2186), .C(n_220475065), .D(n_221575076
		), .Z(n_235075204));
	notech_ao4 i_178847467(.A(n_54735), .B(nbus_11326[24]), .C(n_2311), .D(n_29335
		), .Z(n_235275206));
	notech_ao4 i_178947466(.A(n_55009), .B(n_28059), .C(n_54884), .D(\nbus_11276[0] 
		), .Z(n_235375207));
	notech_ao4 i_179047465(.A(n_2314), .B(n_55413), .C(n_231547139), .D(nbus_11326
		[16]), .Z(n_235675209));
	notech_ao4 i_179147464(.A(n_2247), .B(n_29367), .C(n_2313), .D(n_28908),
		 .Z(n_235775210));
	notech_and4 i_179747458(.A(n_235775210), .B(n_235675209), .C(n_235375207
		), .D(n_235275206), .Z(n_235975212));
	notech_ao4 i_187949158(.A(n_26342), .B(n_149823485), .C(n_57430), .D(n_2249
		), .Z(n_236075213));
	notech_ao4 i_184747408(.A(n_21822205), .B(n_110723094), .C(n_1968), .D(n_1844
		), .Z(n_236175214));
	notech_nand2 i_198849157(.A(n_236175214), .B(n_221675077), .Z(n_236275215
		));
	notech_mux2 i_185047405(.S(opc[2]), .A(n_21822205), .B(n_221875079), .Z(n_236375216
		));
	notech_ao4 i_187247384(.A(n_2313), .B(n_28904), .C(n_2314), .D(n_55277),
		 .Z(n_236475217));
	notech_ao4 i_187347383(.A(n_2248), .B(nbus_11348[3]), .C(n_2247), .D(n_29369
		), .Z(n_236575218));
	notech_and3 i_186847387(.A(n_57312), .B(n_2186), .C(n_222875088), .Z(n_236775220
		));
	notech_ao4 i_186947386(.A(n_2311), .B(n_29325), .C(n_2246), .D(n_27539),
		 .Z(n_236975222));
	notech_ao4 i_187147385(.A(n_231547139), .B(nbus_11326[27]), .C(n_55009),
		 .D(n_28054), .Z(n_237075223));
	notech_and4 i_187747379(.A(n_237075223), .B(n_236975222), .C(n_223775097
		), .D(n_236775220), .Z(n_237275225));
	notech_and4 i_188047377(.A(n_236575218), .B(n_236475217), .C(n_237275225
		), .D(n_223875098), .Z(n_237475227));
	notech_ao4 i_190247355(.A(n_2313), .B(n_28903), .C(n_2314), .D(n_55289),
		 .Z(n_237775230));
	notech_ao4 i_190347354(.A(n_2248), .B(nbus_11348[2]), .C(n_2247), .D(n_29370
		), .Z(n_237875231));
	notech_and3 i_189947358(.A(n_57312), .B(n_2186), .C(n_224475104), .Z(n_238075233
		));
	notech_ao4 i_190047357(.A(n_2311), .B(n_29323), .C(n_2246), .D(n_27538),
		 .Z(n_238275235));
	notech_ao4 i_190147356(.A(n_231547139), .B(nbus_11326[26]), .C(n_55009),
		 .D(n_28053), .Z(n_238375236));
	notech_and4 i_190747350(.A(n_238375236), .B(n_238275235), .C(n_225375113
		), .D(n_238075233), .Z(n_238575238));
	notech_and4 i_190947348(.A(n_237875231), .B(n_237775230), .C(n_238575238
		), .D(n_225475114), .Z(n_238775240));
	notech_ao4 i_196347294(.A(n_2313), .B(n_28901), .C(n_2314), .D(\nbus_11276[0] 
		), .Z(n_239075243));
	notech_ao4 i_196447293(.A(n_2248), .B(nbus_11348[0]), .C(n_29371), .D(n_2247
		), .Z(n_239175244));
	notech_and3 i_196047297(.A(n_57312), .B(n_2186), .C(n_226075120), .Z(n_239375246
		));
	notech_ao4 i_196147296(.A(n_2311), .B(n_29320), .C(n_2246), .D(n_27535),
		 .Z(n_239575248));
	notech_ao4 i_196247295(.A(n_231547139), .B(nbus_11326[24]), .C(n_55009),
		 .D(n_28051), .Z(n_239675249));
	notech_and4 i_196847289(.A(n_239675249), .B(n_239575248), .C(n_227275129
		), .D(n_239375246), .Z(n_239875251));
	notech_and4 i_197047287(.A(n_239175244), .B(n_239075243), .C(n_239875251
		), .D(n_227375130), .Z(n_240075253));
	notech_and4 i_2345350(.A(n_55667), .B(n_55975), .C(n_293161935), .D(n_293761941
		), .Z(n_240475257));
	notech_ao3 i_102445409(.A(n_54748), .B(n_54902), .C(n_46842), .Z(n_240575258
		));
	notech_and3 i_102545410(.A(n_54740), .B(n_46844), .C(n_54872), .Z(n_240675259
		));
	notech_nand3 i_6945308(.A(n_54124), .B(tsc[23]), .C(n_59863), .Z(n_240975262
		));
	notech_or2 i_6845309(.A(n_351665805), .B(nbus_11326[23]), .Z(n_241275265
		));
	notech_or2 i_6345314(.A(n_308921976), .B(n_351865807), .Z(n_241775270)
		);
	notech_nand3 i_9645281(.A(n_54124), .B(tsc[27]), .C(n_59863), .Z(n_241875271
		));
	notech_or2 i_9545282(.A(n_351665805), .B(nbus_11326[27]), .Z(n_242175274
		));
	notech_or2 i_9045287(.A(n_308621973), .B(n_351865807), .Z(n_242875279)
		);
	notech_or2 i_41644967(.A(n_308318860), .B(nbus_11326[25]), .Z(n_242975280
		));
	notech_or2 i_42344960(.A(n_308318860), .B(nbus_11326[26]), .Z(n_244075287
		));
	notech_or2 i_43044953(.A(n_308318860), .B(nbus_11326[27]), .Z(n_244975294
		));
	notech_or2 i_44344946(.A(n_308318860), .B(nbus_11326[28]), .Z(n_245675301
		));
	notech_nao3 i_56944821(.A(n_2464), .B(n_55450), .C(n_54015), .Z(n_246975310
		));
	notech_or2 i_56644824(.A(n_353988269), .B(nbus_11273[25]), .Z(n_247475313
		));
	notech_nand3 i_56344827(.A(n_59193), .B(n_59945), .C(read_data[25]), .Z(n_247775316
		));
	notech_or2 i_56044830(.A(n_308821975), .B(n_354788261), .Z(n_248075319)
		);
	notech_nao3 i_58144809(.A(n_2466), .B(n_55450), .C(n_54015), .Z(n_248375322
		));
	notech_or2 i_57844812(.A(n_353988269), .B(nbus_11273[26]), .Z(n_248675325
		));
	notech_nand3 i_57544815(.A(n_59193), .B(n_59945), .C(read_data[26]), .Z(n_248975328
		));
	notech_or2 i_57244818(.A(n_308721974), .B(n_354788261), .Z(n_249275331)
		);
	notech_nao3 i_60544785(.A(n_2470), .B(n_55450), .C(n_54015), .Z(n_249575334
		));
	notech_or2 i_60244788(.A(n_353488274), .B(nbus_11326[28]), .Z(n_249875337
		));
	notech_or2 i_59944791(.A(n_354888260), .B(n_29219), .Z(n_250175340));
	notech_nand3 i_59644794(.A(n_59193), .B(n_59945), .C(read_data[28]), .Z(n_250475343
		));
	notech_nor2 i_65344737(.A(n_55424), .B(nbus_11326[23]), .Z(n_250575344)
		);
	notech_or2 i_64844742(.A(n_308921976), .B(n_55404), .Z(n_251275351));
	notech_nor2 i_66144729(.A(n_55424), .B(nbus_11326[25]), .Z(n_251375352)
		);
	notech_or4 i_65644734(.A(n_56196), .B(n_58656), .C(n_54367), .D(n_308421971
		), .Z(n_252075359));
	notech_nor2 i_66944721(.A(n_55424), .B(nbus_11326[26]), .Z(n_252175360)
		);
	notech_or4 i_66444726(.A(n_56196), .B(n_58656), .C(n_55798), .D(n_308321970
		), .Z(n_252875367));
	notech_nor2 i_67744713(.A(n_55424), .B(nbus_11326[27]), .Z(n_252975368)
		);
	notech_or4 i_67244718(.A(n_56196), .B(n_58656), .C(n_55794), .D(n_308221969
		), .Z(n_253675375));
	notech_nor2 i_68644705(.A(n_55424), .B(nbus_11326[28]), .Z(n_253775376)
		);
	notech_or2 i_68144710(.A(n_55062), .B(\nbus_11276[28] ), .Z(n_254475383)
		);
	notech_nor2 i_77444617(.A(n_2672), .B(nbus_11326[23]), .Z(n_254575384)
		);
	notech_or2 i_76944622(.A(n_308921976), .B(n_2655), .Z(n_255275391));
	notech_nor2 i_78244609(.A(n_2672), .B(nbus_11326[25]), .Z(n_255375392)
		);
	notech_or4 i_77744614(.A(n_204788866), .B(n_56158), .C(n_55794), .D(n_308421971
		), .Z(n_256075399));
	notech_nor2 i_79044601(.A(n_2672), .B(nbus_11326[26]), .Z(n_256175400)
		);
	notech_or4 i_78544606(.A(n_204788866), .B(n_56158), .C(n_55794), .D(n_308321970
		), .Z(n_256875407));
	notech_nor2 i_79844593(.A(n_2672), .B(nbus_11326[27]), .Z(n_256975408)
		);
	notech_or4 i_79344598(.A(n_204788866), .B(n_56158), .C(n_55798), .D(n_308221969
		), .Z(n_257675415));
	notech_nor2 i_80644585(.A(n_2672), .B(nbus_11326[28]), .Z(n_257775416)
		);
	notech_or2 i_80144590(.A(n_55069), .B(\nbus_11276[28] ), .Z(n_258475423)
		);
	notech_nor2 i_81444577(.A(n_55070), .B(nbus_11273[23]), .Z(n_258575424)
		);
	notech_or2 i_80944582(.A(n_308521972), .B(n_309921986), .Z(n_259275431)
		);
	notech_nor2 i_81744574(.A(n_56057), .B(\nbus_11276[23] ), .Z(n_259675435
		));
	notech_or2 i_82544566(.A(n_55070), .B(nbus_11273[25]), .Z(n_259775436)
		);
	notech_or2 i_83844553(.A(n_55070), .B(nbus_11273[26]), .Z(n_260475443)
		);
	notech_or4 i_84244549(.A(n_60782), .B(n_60729), .C(n_54761), .D(n_29156)
		, .Z(n_261575454));
	notech_or2 i_85144540(.A(n_55070), .B(nbus_11273[27]), .Z(n_261675455)
		);
	notech_or4 i_85544536(.A(n_60782), .B(n_60729), .C(n_54761), .D(n_29154)
		, .Z(n_262775466));
	notech_or2 i_86444527(.A(n_55070), .B(nbus_11273[28]), .Z(n_262875467)
		);
	notech_or2 i_4645331(.A(n_240475257), .B(n_294261946), .Z(n_263575474)
		);
	notech_ao4 i_187943554(.A(n_55965), .B(n_304221929), .C(n_303521922), .D
		(nbus_11326[28]), .Z(n_263675475));
	notech_ao4 i_187843555(.A(n_57330), .B(n_55396), .C(n_343565725), .D(n_306621953
		), .Z(n_263775476));
	notech_ao4 i_187643557(.A(n_55071), .B(\nbus_11276[28] ), .C(n_29219), .D
		(n_55397), .Z(n_263975478));
	notech_and3 i_187743556(.A(n_263975478), .B(n_26249), .C(n_262875467), .Z
		(n_264175480));
	notech_ao4 i_187043563(.A(n_304121928), .B(n_55965), .C(n_303521922), .D
		(nbus_11326[27]), .Z(n_264275481));
	notech_ao4 i_186943564(.A(n_308621973), .B(n_55396), .C(n_286061878), .D
		(n_306621953), .Z(n_264375482));
	notech_ao4 i_186743566(.A(n_55071), .B(\nbus_11276[27] ), .C(n_29154), .D
		(n_55397), .Z(n_264575484));
	notech_ao4 i_187343560(.A(n_59863), .B(n_27550), .C(n_101213406), .D(n_308621973
		), .Z(n_264675485));
	notech_ao4 i_187243561(.A(n_98113375), .B(nbus_11273[27]), .C(n_56057), 
		.D(\nbus_11276[27] ), .Z(n_264875487));
	notech_nand3 i_45345374(.A(n_264675485), .B(n_264875487), .C(n_262775466
		), .Z(n_264975488));
	notech_ao3 i_186843565(.A(n_264575484), .B(n_261675455), .C(n_264975488)
		, .Z(n_265175490));
	notech_ao4 i_186143572(.A(n_55965), .B(n_304021927), .C(n_303521922), .D
		(nbus_11326[26]), .Z(n_265275491));
	notech_ao4 i_186043573(.A(n_308721974), .B(n_55396), .C(n_288561889), .D
		(n_306621953), .Z(n_265375492));
	notech_ao4 i_185843575(.A(n_55071), .B(\nbus_11276[26] ), .C(n_29156), .D
		(n_55397), .Z(n_265575494));
	notech_ao4 i_186443569(.A(n_59863), .B(n_27549), .C(n_101213406), .D(n_308721974
		), .Z(n_265675495));
	notech_ao4 i_186343570(.A(n_98113375), .B(nbus_11273[26]), .C(n_56216), 
		.D(\nbus_11276[26] ), .Z(n_265875497));
	notech_nand3 i_44145376(.A(n_265675495), .B(n_265875497), .C(n_261575454
		), .Z(n_265975498));
	notech_and3 i_185943574(.A(n_265575494), .B(n_26413), .C(n_260475443), .Z
		(n_266175500));
	notech_ao4 i_185243581(.A(n_303921926), .B(n_55965), .C(n_303521922), .D
		(nbus_11326[25]), .Z(n_266275501));
	notech_ao4 i_185143582(.A(n_308821975), .B(n_55396), .C(n_268264999), .D
		(n_306621953), .Z(n_266375502));
	notech_ao4 i_184943584(.A(n_55071), .B(\nbus_11276[25] ), .C(n_29215), .D
		(n_55397), .Z(n_266575504));
	notech_and3 i_185043583(.A(n_266575504), .B(n_26308), .C(n_259775436), .Z
		(n_266775506));
	notech_ao4 i_184243591(.A(n_270765024), .B(n_306621953), .C(n_303521922)
		, .D(nbus_11326[23]), .Z(n_266875507));
	notech_ao4 i_184143592(.A(n_29152), .B(n_55397), .C(n_308921976), .D(n_55396
		), .Z(n_267075509));
	notech_nand3 i_184443589(.A(n_266875507), .B(n_267075509), .C(n_259275431
		), .Z(n_267175510));
	notech_ao4 i_183943594(.A(n_55071), .B(\nbus_11276[23] ), .C(n_27590), .D
		(n_55719), .Z(n_267275511));
	notech_ao4 i_184643587(.A(n_101413408), .B(n_29152), .C(n_101213406), .D
		(n_308921976), .Z(n_267375512));
	notech_ao4 i_184543588(.A(n_27545), .B(n_59863), .C(n_98113375), .D(nbus_11273
		[23]), .Z(n_267575514));
	notech_nao3 i_68045373(.A(n_267375512), .B(n_267575514), .C(n_259675435)
		, .Z(n_267675515));
	notech_ao4 i_183543598(.A(n_57330), .B(n_2655), .C(n_307421961), .D(n_56139
		), .Z(n_267975518));
	notech_ao4 i_183443599(.A(n_29219), .B(n_26444), .C(n_55068), .D(nbus_11273
		[28]), .Z(n_268175520));
	notech_nand3 i_183743596(.A(n_267975518), .B(n_268175520), .C(n_258475423
		), .Z(n_268275521));
	notech_ao4 i_183243601(.A(n_343565725), .B(n_2694), .C(n_57306), .D(n_2674
		), .Z(n_268375522));
	notech_ao4 i_182843605(.A(n_286061878), .B(n_2694), .C(n_56139), .D(n_303621923
		), .Z(n_268675525));
	notech_ao4 i_182743606(.A(n_29154), .B(n_26444), .C(n_308621973), .D(n_2655
		), .Z(n_268875527));
	notech_nand3 i_183043603(.A(n_268675525), .B(n_268875527), .C(n_257675415
		), .Z(n_268975528));
	notech_ao4 i_182543608(.A(n_55068), .B(nbus_11273[27]), .C(n_55069), .D(\nbus_11276[27] 
		), .Z(n_269075529));
	notech_ao4 i_182143612(.A(n_288561889), .B(n_2694), .C(n_307621963), .D(n_56139
		), .Z(n_269375532));
	notech_ao4 i_182043613(.A(n_29156), .B(n_26444), .C(n_308721974), .D(n_2655
		), .Z(n_269575534));
	notech_nand3 i_182343610(.A(n_269375532), .B(n_269575534), .C(n_256875407
		), .Z(n_269675535));
	notech_ao4 i_181843615(.A(n_55068), .B(nbus_11273[26]), .C(n_55069), .D(\nbus_11276[26] 
		), .Z(n_269775536));
	notech_ao4 i_181443619(.A(n_268264999), .B(n_2694), .C(n_307521962), .D(n_56139
		), .Z(n_270075539));
	notech_ao4 i_181343620(.A(n_29215), .B(n_26444), .C(n_308821975), .D(n_2655
		), .Z(n_270275541));
	notech_nand3 i_181643617(.A(n_270075539), .B(n_270275541), .C(n_256075399
		), .Z(n_270375542));
	notech_ao4 i_181143622(.A(n_55068), .B(nbus_11273[25]), .C(n_55069), .D(\nbus_11276[25] 
		), .Z(n_270475543));
	notech_ao4 i_180743626(.A(n_308521972), .B(n_2674), .C(n_270765024), .D(n_2694
		), .Z(n_270775546));
	notech_ao4 i_180643627(.A(n_29152), .B(n_26444), .C(n_27590), .D(n_55717
		), .Z(n_270975548));
	notech_nand3 i_180943624(.A(n_270775546), .B(n_270975548), .C(n_255275391
		), .Z(n_271075549));
	notech_ao4 i_180443629(.A(nbus_11273[23]), .B(n_55068), .C(n_55069), .D(\nbus_11276[23] 
		), .Z(n_271175550));
	notech_ao4 i_172943703(.A(n_57330), .B(n_55404), .C(n_307421961), .D(n_56382
		), .Z(n_271475553));
	notech_ao4 i_172843704(.A(n_29219), .B(n_55405), .C(n_55064), .D(nbus_11273
		[28]), .Z(n_271675555));
	notech_nand3 i_173143701(.A(n_271475553), .B(n_271675555), .C(n_254475383
		), .Z(n_271775556));
	notech_ao4 i_172643706(.A(n_343565725), .B(n_308418861), .C(n_57306), .D
		(n_309618873), .Z(n_271875557));
	notech_ao4 i_172243710(.A(n_286061878), .B(n_308418861), .C(n_56382), .D
		(n_303621923), .Z(n_272175560));
	notech_ao4 i_172143711(.A(n_29154), .B(n_55405), .C(n_308621973), .D(n_55404
		), .Z(n_272375562));
	notech_nand3 i_172443708(.A(n_272175560), .B(n_272375562), .C(n_253675375
		), .Z(n_272475563));
	notech_ao4 i_171943713(.A(n_55064), .B(nbus_11273[27]), .C(n_55062), .D(\nbus_11276[27] 
		), .Z(n_272575564));
	notech_ao4 i_171543717(.A(n_288561889), .B(n_308418861), .C(n_307621963)
		, .D(n_56382), .Z(n_272875567));
	notech_ao4 i_171443718(.A(n_29156), .B(n_55405), .C(n_308721974), .D(n_55404
		), .Z(n_273075569));
	notech_nand3 i_171743715(.A(n_272875567), .B(n_273075569), .C(n_252875367
		), .Z(n_273175570));
	notech_ao4 i_171243720(.A(n_55064), .B(nbus_11273[26]), .C(n_55062), .D(\nbus_11276[26] 
		), .Z(n_273275571));
	notech_ao4 i_170743724(.A(n_268264999), .B(n_308418861), .C(n_307521962)
		, .D(n_56382), .Z(n_273575574));
	notech_ao4 i_170643725(.A(n_29215), .B(n_55405), .C(n_308821975), .D(n_55404
		), .Z(n_273775576));
	notech_nand3 i_170943722(.A(n_273575574), .B(n_273775576), .C(n_252075359
		), .Z(n_273875577));
	notech_ao4 i_170443727(.A(n_55064), .B(nbus_11273[25]), .C(n_55062), .D(\nbus_11276[25] 
		), .Z(n_273975578));
	notech_ao4 i_170043731(.A(n_308521972), .B(n_309618873), .C(n_270765024)
		, .D(n_308418861), .Z(n_274275581));
	notech_ao4 i_169943732(.A(n_29152), .B(n_55405), .C(n_27590), .D(n_55720
		), .Z(n_274475583));
	notech_nand3 i_170243729(.A(n_274275581), .B(n_274475583), .C(n_251275351
		), .Z(n_274575584));
	notech_ao4 i_169743734(.A(nbus_11273[23]), .B(n_55064), .C(n_55062), .D(\nbus_11276[23] 
		), .Z(n_274675585));
	notech_ao4 i_165843773(.A(n_59193), .B(n_26771), .C(n_57330), .D(n_354788261
		), .Z(n_274975588));
	notech_ao4 i_165643775(.A(n_353988269), .B(nbus_11273[28]), .C(n_354488264
		), .D(\nbus_11276[28] ), .Z(n_275175590));
	notech_and4 i_166043771(.A(n_275175590), .B(n_274975588), .C(n_250175340
		), .D(n_250475343), .Z(n_275375592));
	notech_ao4 i_165343778(.A(n_354988259), .B(n_343565725), .C(n_57306), .D
		(n_354388265), .Z(n_275475593));
	notech_ao4 i_165143780(.A(n_53993), .B(n_29374), .C(n_5538), .D(n_27596)
		, .Z(n_275675595));
	notech_and4 i_165543776(.A(n_275675595), .B(n_275475593), .C(n_249575334
		), .D(n_249875337), .Z(n_275875597));
	notech_ao4 i_163843793(.A(n_308321970), .B(n_354388265), .C(n_354988259)
		, .D(n_288561889), .Z(n_275975598));
	notech_ao4 i_163643795(.A(n_5538), .B(n_27594), .C(n_59195), .D(n_26769)
		, .Z(n_276175600));
	notech_and4 i_164043791(.A(n_276175600), .B(n_275975598), .C(n_248975328
		), .D(n_249275331), .Z(n_276375602));
	notech_ao4 i_163343798(.A(n_354488264), .B(\nbus_11276[26] ), .C(n_354888260
		), .D(n_29156), .Z(n_276475603));
	notech_ao4 i_163143800(.A(n_53993), .B(n_29373), .C(n_353488274), .D(nbus_11326
		[26]), .Z(n_276675605));
	notech_and4 i_163543796(.A(n_276675605), .B(n_276475603), .C(n_248375322
		), .D(n_248675325), .Z(n_276875607));
	notech_ao4 i_162843803(.A(n_308421971), .B(n_354388265), .C(n_268264999)
		, .D(n_354988259), .Z(n_276975608));
	notech_ao4 i_162643805(.A(n_5538), .B(n_27593), .C(n_59195), .D(n_26767)
		, .Z(n_277175610));
	notech_and4 i_163043801(.A(n_277175610), .B(n_276975608), .C(n_247775316
		), .D(n_248075319), .Z(n_277375612));
	notech_ao4 i_162343808(.A(n_354488264), .B(\nbus_11276[25] ), .C(n_354888260
		), .D(n_29215), .Z(n_277475613));
	notech_ao4 i_162143810(.A(n_53993), .B(n_29372), .C(n_353488274), .D(nbus_11326
		[25]), .Z(n_277675615));
	notech_and4 i_162543806(.A(n_277675615), .B(n_277475613), .C(n_246975310
		), .D(n_247475313), .Z(n_277875617));
	notech_ao4 i_152243903(.A(n_55906), .B(n_304221929), .C(n_343565725), .D
		(n_263575474), .Z(n_277975618));
	notech_ao4 i_152143904(.A(n_57330), .B(n_240675259), .C(n_240575258), .D
		(n_29219), .Z(n_278075619));
	notech_ao4 i_151943906(.A(n_55219), .B(n_56883), .C(n_55218), .D(\nbus_11276[28] 
		), .Z(n_278275621));
	notech_and3 i_152043905(.A(n_278275621), .B(n_26249), .C(n_245675301), .Z
		(n_278475623));
	notech_ao4 i_151643909(.A(n_304121928), .B(n_55906), .C(n_286061878), .D
		(n_263575474), .Z(n_278575624));
	notech_ao4 i_151543910(.A(n_240575258), .B(n_29154), .C(n_308621973), .D
		(n_240675259), .Z(n_278675625));
	notech_ao4 i_151343912(.A(n_55219), .B(n_56874), .C(n_55218), .D(\nbus_11276[27] 
		), .Z(n_278875627));
	notech_ao3 i_151443911(.A(n_278875627), .B(n_244975294), .C(n_264975488)
		, .Z(n_279075629));
	notech_ao4 i_151043915(.A(n_55906), .B(n_304021927), .C(n_288561889), .D
		(n_263575474), .Z(n_279175630));
	notech_ao4 i_150943916(.A(n_240575258), .B(n_29156), .C(n_308721974), .D
		(n_240675259), .Z(n_279275631));
	notech_ao4 i_150743918(.A(n_55219), .B(n_56865), .C(n_55218), .D(\nbus_11276[26] 
		), .Z(n_279475633));
	notech_and3 i_150843917(.A(n_279475633), .B(n_26413), .C(n_244075287), .Z
		(n_279675635));
	notech_ao4 i_150443921(.A(n_303921926), .B(n_55906), .C(n_268264999), .D
		(n_263575474), .Z(n_279775636));
	notech_ao4 i_150343922(.A(n_29215), .B(n_240575258), .C(n_308821975), .D
		(n_240675259), .Z(n_279875637));
	notech_ao4 i_150143924(.A(n_55219), .B(n_56856), .C(n_55218), .D(\nbus_11276[25] 
		), .Z(n_280075639));
	notech_and3 i_150243923(.A(n_280075639), .B(n_26308), .C(n_242975280), .Z
		(n_280275641));
	notech_ao4 i_117444244(.A(n_308221969), .B(n_352265811), .C(n_286061878)
		, .D(n_352865817), .Z(n_280375642));
	notech_ao4 i_117344245(.A(n_351765806), .B(n_29154), .C(n_351165800), .D
		(n_27595), .Z(n_280575644));
	notech_ao4 i_117044248(.A(n_55143), .B(n_56874), .C(n_55142), .D(\nbus_11276[27] 
		), .Z(n_280775646));
	notech_and4 i_117244246(.A(n_280775646), .B(n_241875271), .C(n_242175274
		), .D(n_26412), .Z(n_281075649));
	notech_ao4 i_114844268(.A(n_308521972), .B(n_352265811), .C(n_270765024)
		, .D(n_352865817), .Z(n_281175650));
	notech_ao4 i_114744269(.A(n_29152), .B(n_351765806), .C(n_351165800), .D
		(n_27590), .Z(n_281375652));
	notech_ao4 i_114444272(.A(n_55143), .B(nbus_11273[23]), .C(n_55142), .D(\nbus_11276[23] 
		), .Z(n_281575654));
	notech_and4 i_114644270(.A(n_281575654), .B(n_240975262), .C(n_241275265
		), .D(n_26414), .Z(n_281875657));
	notech_nand3 i_2942213(.A(n_54128), .B(tsc[18]), .C(n_59863), .Z(n_281975658
		));
	notech_or2 i_2842214(.A(n_351665805), .B(nbus_11326[18]), .Z(n_282275661
		));
	notech_or2 i_2042219(.A(n_311318890), .B(n_351865807), .Z(n_282775666)
		);
	notech_nand3 i_3842204(.A(n_54128), .B(tsc[19]), .C(n_59865), .Z(n_282875667
		));
	notech_or2 i_3742205(.A(n_351665805), .B(nbus_11326[19]), .Z(n_283175670
		));
	notech_or2 i_3242210(.A(n_311218889), .B(n_351865807), .Z(n_283675675)
		);
	notech_nand3 i_4742195(.A(n_54128), .B(tsc[20]), .C(n_59863), .Z(n_283775676
		));
	notech_or2 i_4642196(.A(n_351665805), .B(nbus_11326[20]), .Z(n_284075679
		));
	notech_or2 i_4142201(.A(n_311118888), .B(n_351865807), .Z(n_284575684)
		);
	notech_nand3 i_5642186(.A(n_54128), .B(tsc[21]), .C(n_59863), .Z(n_284675685
		));
	notech_or2 i_5542187(.A(n_351665805), .B(nbus_11326[21]), .Z(n_284975688
		));
	notech_or2 i_5042192(.A(n_311018887), .B(n_351865807), .Z(n_285475693)
		);
	notech_nand3 i_6542177(.A(n_54128), .B(tsc[22]), .C(n_59863), .Z(n_285575694
		));
	notech_or2 i_6442178(.A(n_351665805), .B(nbus_11326[22]), .Z(n_285875697
		));
	notech_or2 i_5942183(.A(n_26618), .B(n_351865807), .Z(n_286375702));
	notech_or2 i_26641977(.A(n_303421921), .B(nbus_11326[22]), .Z(n_286675705
		));
	notech_or2 i_26141982(.A(n_26618), .B(n_55556), .Z(n_287175710));
	notech_or2 i_39541852(.A(n_55555), .B(n_29174), .Z(n_287275711));
	notech_or4 i_39041857(.A(n_56158), .B(n_206288851), .C(n_310418881), .D(n_55523
		), .Z(n_287975718));
	notech_or2 i_60441647(.A(n_123423221), .B(nbus_11326[22]), .Z(n_288075719
		));
	notech_or2 i_59941652(.A(n_26618), .B(n_2702), .Z(n_288775726));
	notech_nor2 i_61241639(.A(n_55062), .B(\nbus_11276[18] ), .Z(n_288875727
		));
	notech_or2 i_60741644(.A(n_311318890), .B(n_55404), .Z(n_289575734));
	notech_nor2 i_62041631(.A(n_55062), .B(\nbus_11276[19] ), .Z(n_289675735
		));
	notech_or2 i_61541636(.A(n_311218889), .B(n_55404), .Z(n_290375742));
	notech_nor2 i_62841623(.A(n_55062), .B(\nbus_11276[20] ), .Z(n_290475743
		));
	notech_or2 i_62341628(.A(n_311118888), .B(n_55404), .Z(n_291175750));
	notech_nor2 i_63741615(.A(n_55062), .B(\nbus_11276[21] ), .Z(n_291275751
		));
	notech_or2 i_63241620(.A(n_311018887), .B(n_55404), .Z(n_291975758));
	notech_or2 i_64541607(.A(n_55062), .B(\nbus_11276[22] ), .Z(n_292075759)
		);
	notech_or2 i_64041612(.A(n_26618), .B(n_55404), .Z(n_292775766));
	notech_or2 i_68541572(.A(n_26618), .B(n_353365822), .Z(n_293575774));
	notech_nor2 i_73841519(.A(n_2672), .B(nbus_11326[18]), .Z(n_293675775)
		);
	notech_or2 i_73341524(.A(n_311318890), .B(n_2655), .Z(n_294375782));
	notech_nor2 i_74641511(.A(n_2672), .B(nbus_11326[19]), .Z(n_294475783)
		);
	notech_or2 i_74141516(.A(n_311218889), .B(n_2655), .Z(n_295175790));
	notech_nor2 i_75441503(.A(n_2672), .B(nbus_11326[20]), .Z(n_295275791)
		);
	notech_or2 i_74941508(.A(n_311118888), .B(n_2655), .Z(n_295975798));
	notech_nor2 i_76241495(.A(n_2672), .B(nbus_11326[21]), .Z(n_296075799)
		);
	notech_or2 i_75741500(.A(n_311018887), .B(n_2655), .Z(n_296775806));
	notech_or2 i_77041487(.A(n_2672), .B(nbus_11326[22]), .Z(n_296875807));
	notech_or2 i_76541492(.A(n_26618), .B(n_2655), .Z(n_297575814));
	notech_nor2 i_77841479(.A(n_303521922), .B(nbus_11326[18]), .Z(n_297675815
		));
	notech_or2 i_77341484(.A(n_311318890), .B(n_55396), .Z(n_298375822));
	notech_nor2 i_79041467(.A(n_303521922), .B(nbus_11326[19]), .Z(n_298475823
		));
	notech_or2 i_78541472(.A(n_311218889), .B(n_55396), .Z(n_299175830));
	notech_nor2 i_79341464(.A(n_56216), .B(\nbus_11276[19] ), .Z(n_299575834
		));
	notech_nor2 i_80441455(.A(n_303521922), .B(nbus_11326[20]), .Z(n_299675835
		));
	notech_or2 i_79941460(.A(n_311118888), .B(n_55396), .Z(n_300375842));
	notech_nor2 i_81841443(.A(n_303521922), .B(nbus_11326[21]), .Z(n_300475843
		));
	notech_or2 i_81141448(.A(n_311018887), .B(n_55396), .Z(n_301175850));
	notech_nor2 i_82141440(.A(n_56216), .B(\nbus_11276[21] ), .Z(n_301575854
		));
	notech_or2 i_83041431(.A(n_303521922), .B(nbus_11326[22]), .Z(n_301675855
		));
	notech_or2 i_82541436(.A(n_26618), .B(n_55396), .Z(n_302375862));
	notech_nor2 i_83341428(.A(n_56216), .B(\nbus_11276[22] ), .Z(n_302775866
		));
	notech_ao4 i_186940423(.A(n_310418881), .B(n_309921986), .C(n_305565372)
		, .D(n_306621953), .Z(n_302875867));
	notech_ao4 i_186840424(.A(n_29174), .B(n_55397), .C(n_55719), .D(n_27589
		), .Z(n_303075869));
	notech_and3 i_187140421(.A(n_302875867), .B(n_303075869), .C(n_302375862
		), .Z(n_303175870));
	notech_ao4 i_186640426(.A(n_55070), .B(nbus_11273[22]), .C(n_55071), .D(\nbus_11276[22] 
		), .Z(n_303275871));
	notech_ao4 i_187340419(.A(n_101413408), .B(n_29174), .C(n_26618), .D(n_101213406
		), .Z(n_303375872));
	notech_ao4 i_187240420(.A(n_27542), .B(n_59863), .C(n_98113375), .D(nbus_11273
		[22]), .Z(n_303575874));
	notech_ao3 i_67942245(.A(n_303375872), .B(n_303575874), .C(n_302775866),
		 .Z(n_303675875));
	notech_ao4 i_185940433(.A(n_310518882), .B(n_309921986), .C(n_312662130)
		, .D(n_306621953), .Z(n_303975878));
	notech_ao4 i_185840434(.A(n_29172), .B(n_55397), .C(n_55719), .D(n_27588
		), .Z(n_304175880));
	notech_nand3 i_186140431(.A(n_303975878), .B(n_304175880), .C(n_301175850
		), .Z(n_304275881));
	notech_ao4 i_185640436(.A(n_55070), .B(nbus_11273[21]), .C(n_55071), .D(\nbus_11276[21] 
		), .Z(n_304375882));
	notech_ao4 i_186340429(.A(n_101413408), .B(n_29172), .C(n_311018887), .D
		(n_101213406), .Z(n_304475883));
	notech_ao4 i_186240430(.A(n_27541), .B(n_59863), .C(n_98113375), .D(nbus_11273
		[21]), .Z(n_304675885));
	notech_nao3 i_67842246(.A(n_304475883), .B(n_304675885), .C(n_301575854)
		, .Z(n_304775886));
	notech_ao4 i_184940443(.A(n_310618883), .B(n_309921986), .C(n_315162155)
		, .D(n_306621953), .Z(n_305075889));
	notech_ao4 i_184840444(.A(n_29169), .B(n_55397), .C(n_55719), .D(n_27586
		), .Z(n_305275891));
	notech_nand3 i_185140441(.A(n_305075889), .B(n_305275891), .C(n_300375842
		), .Z(n_305375892));
	notech_ao4 i_184640446(.A(n_55070), .B(nbus_11273[20]), .C(n_55071), .D(\nbus_11276[20] 
		), .Z(n_305475893));
	notech_ao4 i_183940453(.A(n_310718884), .B(n_309921986), .C(n_308065397)
		, .D(n_306621953), .Z(n_305775896));
	notech_ao4 i_183840454(.A(n_29167), .B(n_55397), .C(n_55719), .D(n_27585
		), .Z(n_305975898));
	notech_nand3 i_184140451(.A(n_305775896), .B(n_305975898), .C(n_299175830
		), .Z(n_306075899));
	notech_ao4 i_183640456(.A(n_55070), .B(nbus_11273[19]), .C(n_55071), .D(\nbus_11276[19] 
		), .Z(n_306175900));
	notech_ao4 i_184340449(.A(n_101413408), .B(n_29167), .C(n_311218889), .D
		(n_101213406), .Z(n_306275901));
	notech_ao4 i_184240450(.A(n_27539), .B(n_59863), .C(n_98113375), .D(nbus_11273
		[19]), .Z(n_306475903));
	notech_nao3 i_67642248(.A(n_306275901), .B(n_306475903), .C(n_299575834)
		, .Z(n_306575904));
	notech_ao4 i_182940463(.A(n_310818885), .B(n_309921986), .C(n_310565422)
		, .D(n_306621953), .Z(n_306875907));
	notech_ao4 i_182840464(.A(n_29165), .B(n_55397), .C(n_55719), .D(n_27584
		), .Z(n_307075909));
	notech_nand3 i_183140461(.A(n_306875907), .B(n_307075909), .C(n_298375822
		), .Z(n_307175910));
	notech_ao4 i_182640466(.A(n_55070), .B(nbus_11273[18]), .C(n_55071), .D(\nbus_11276[18] 
		), .Z(n_307275911));
	notech_ao4 i_182240470(.A(n_310418881), .B(n_2674), .C(n_305565372), .D(n_2694
		), .Z(n_307575914));
	notech_ao4 i_182140471(.A(n_29174), .B(n_26444), .C(n_55717), .D(n_27589
		), .Z(n_307775916));
	notech_and3 i_182440468(.A(n_307575914), .B(n_307775916), .C(n_297575814
		), .Z(n_307875917));
	notech_ao4 i_181940473(.A(n_55068), .B(nbus_11273[22]), .C(n_55069), .D(\nbus_11276[22] 
		), .Z(n_307975918));
	notech_ao4 i_181540477(.A(n_310518882), .B(n_2674), .C(n_312662130), .D(n_2694
		), .Z(n_308275921));
	notech_ao4 i_181440478(.A(n_29172), .B(n_26444), .C(n_55717), .D(n_27588
		), .Z(n_308475923));
	notech_nand3 i_181740475(.A(n_308275921), .B(n_308475923), .C(n_296775806
		), .Z(n_308575924));
	notech_ao4 i_181240480(.A(n_55068), .B(nbus_11273[21]), .C(n_55069), .D(\nbus_11276[21] 
		), .Z(n_308675925));
	notech_ao4 i_180840484(.A(n_310618883), .B(n_2674), .C(n_315162155), .D(n_2694
		), .Z(n_308975928));
	notech_ao4 i_180740485(.A(n_29169), .B(n_26444), .C(n_55717), .D(n_27586
		), .Z(n_309175930));
	notech_nand3 i_181040482(.A(n_308975928), .B(n_309175930), .C(n_295975798
		), .Z(n_309275931));
	notech_ao4 i_180540487(.A(n_55068), .B(nbus_11273[20]), .C(n_55069), .D(\nbus_11276[20] 
		), .Z(n_309375932));
	notech_ao4 i_180140491(.A(n_310718884), .B(n_2674), .C(n_308065397), .D(n_2694
		), .Z(n_309675935));
	notech_ao4 i_180040492(.A(n_29167), .B(n_26444), .C(n_55717), .D(n_27585
		), .Z(n_309875937));
	notech_nand3 i_180340489(.A(n_309675935), .B(n_309875937), .C(n_295175790
		), .Z(n_309975938));
	notech_ao4 i_179840494(.A(n_55068), .B(nbus_11273[19]), .C(n_55069), .D(\nbus_11276[19] 
		), .Z(n_310075939));
	notech_ao4 i_179440498(.A(n_310818885), .B(n_2674), .C(n_310565422), .D(n_2694
		), .Z(n_310375942));
	notech_ao4 i_179340499(.A(n_29165), .B(n_26444), .C(n_55717), .D(n_27584
		), .Z(n_310575944));
	notech_nand3 i_179640496(.A(n_310375942), .B(n_310575944), .C(n_294375782
		), .Z(n_310675945));
	notech_ao4 i_179140501(.A(n_55068), .B(nbus_11273[18]), .C(n_55069), .D(\nbus_11276[18] 
		), .Z(n_310775946));
	notech_ao4 i_175240540(.A(n_310418881), .B(n_121523202), .C(n_305565372)
		, .D(n_121723204), .Z(n_311075949));
	notech_ao4 i_175140541(.A(n_353165820), .B(n_29174), .C(n_353465823), .D
		(n_27589), .Z(n_311275951));
	notech_and3 i_175440538(.A(n_311075949), .B(n_311275951), .C(n_293575774
		), .Z(n_311375952));
	notech_ao4 i_174940543(.A(n_353265821), .B(nbus_11273[22]), .C(n_26572),
		 .D(\nbus_11276[22] ), .Z(n_311475953));
	notech_ao4 i_174840544(.A(n_27542), .B(n_59856), .C(n_121623203), .D(nbus_11326
		[22]), .Z(n_311575954));
	notech_ao4 i_171640575(.A(n_310418881), .B(n_309618873), .C(n_305565372)
		, .D(n_308418861), .Z(n_311775956));
	notech_ao4 i_171540576(.A(n_29174), .B(n_55405), .C(n_55720), .D(n_27589
		), .Z(n_311975958));
	notech_and3 i_171840573(.A(n_311775956), .B(n_311975958), .C(n_292775766
		), .Z(n_312075959));
	notech_ao4 i_171240578(.A(n_55064), .B(nbus_11273[22]), .C(n_55424), .D(nbus_11326
		[22]), .Z(n_312175960));
	notech_ao4 i_170840582(.A(n_310518882), .B(n_309618873), .C(n_312662130)
		, .D(n_308418861), .Z(n_312475963));
	notech_ao4 i_170740583(.A(n_29172), .B(n_55405), .C(n_55720), .D(n_27588
		), .Z(n_312675965));
	notech_nand3 i_171040580(.A(n_312475963), .B(n_312675965), .C(n_291975758
		), .Z(n_312775966));
	notech_ao4 i_170540585(.A(n_55064), .B(nbus_11273[21]), .C(n_55424), .D(nbus_11326
		[21]), .Z(n_312875967));
	notech_ao4 i_170140589(.A(n_310618883), .B(n_309618873), .C(n_315162155)
		, .D(n_308418861), .Z(n_313175970));
	notech_ao4 i_170040590(.A(n_29169), .B(n_55405), .C(n_55720), .D(n_27586
		), .Z(n_313375972));
	notech_nand3 i_170340587(.A(n_313175970), .B(n_313375972), .C(n_291175750
		), .Z(n_313475973));
	notech_ao4 i_169840592(.A(n_55064), .B(nbus_11273[20]), .C(n_55424), .D(nbus_11326
		[20]), .Z(n_313575974));
	notech_ao4 i_169440596(.A(n_310718884), .B(n_309618873), .C(n_308065397)
		, .D(n_308418861), .Z(n_313875977));
	notech_ao4 i_169340597(.A(n_29167), .B(n_55405), .C(n_55720), .D(n_27585
		), .Z(n_314075979));
	notech_nand3 i_169640594(.A(n_313875977), .B(n_314075979), .C(n_290375742
		), .Z(n_314175980));
	notech_ao4 i_169140599(.A(n_55064), .B(nbus_11273[19]), .C(n_55424), .D(nbus_11326
		[19]), .Z(n_314275981));
	notech_ao4 i_168740603(.A(n_310818885), .B(n_309618873), .C(n_310565422)
		, .D(n_308418861), .Z(n_314575984));
	notech_ao4 i_168640604(.A(n_29165), .B(n_55405), .C(n_55720), .D(n_27584
		), .Z(n_314775986));
	notech_nand3 i_168940601(.A(n_314575984), .B(n_314775986), .C(n_289575734
		), .Z(n_314875987));
	notech_ao4 i_168440606(.A(n_55064), .B(nbus_11273[18]), .C(n_55424), .D(nbus_11326
		[18]), .Z(n_314975988));
	notech_ao4 i_168040610(.A(n_310418881), .B(n_123223219), .C(n_123623223)
		, .D(n_305565372), .Z(n_315275991));
	notech_ao4 i_167940611(.A(n_26450), .B(n_29174), .C(n_181471126), .D(n_27589
		), .Z(n_315475993));
	notech_and3 i_168240608(.A(n_315275991), .B(n_315475993), .C(n_288775726
		), .Z(n_315575994));
	notech_ao4 i_167740613(.A(n_55073), .B(nbus_11273[22]), .C(n_55072), .D(\nbus_11276[22] 
		), .Z(n_315675995));
	notech_ao4 i_150340780(.A(n_308718864), .B(n_305565372), .C(n_308318860)
		, .D(nbus_11326[22]), .Z(n_315975998));
	notech_ao4 i_150240781(.A(n_55773), .B(n_27589), .C(n_26618), .D(n_55554
		), .Z(n_316176000));
	notech_and3 i_150540778(.A(n_315975998), .B(n_316176000), .C(n_287975718
		), .Z(n_316276001));
	notech_ao4 i_150040783(.A(n_55219), .B(n_56829), .C(n_55218), .D(\nbus_11276[22] 
		), .Z(n_316376002));
	notech_ao4 i_133340943(.A(n_310418881), .B(n_322631613), .C(n_305565372)
		, .D(n_322931616), .Z(n_316676005));
	notech_ao4 i_133240944(.A(n_55557), .B(n_29174), .C(n_55772), .D(n_27589
		), .Z(n_316876007));
	notech_ao4 i_132940947(.A(n_55220), .B(n_56829), .C(n_55221), .D(n_55647
		), .Z(n_317076009));
	notech_and4 i_133140945(.A(n_53844), .B(n_303675875), .C(n_317076009), .D
		(n_286675705), .Z(n_317376012));
	notech_ao4 i_114341128(.A(n_310418881), .B(n_352265811), .C(n_305565372)
		, .D(n_352865817), .Z(n_317476013));
	notech_ao4 i_114241129(.A(n_351765806), .B(n_29174), .C(n_351165800), .D
		(n_27589), .Z(n_317676015));
	notech_ao4 i_113941132(.A(n_55143), .B(n_56829), .C(n_55142), .D(n_55647
		), .Z(n_317876017));
	notech_and4 i_114141130(.A(n_303675875), .B(n_317876017), .C(n_285575694
		), .D(n_285875697), .Z(n_318176020));
	notech_ao4 i_113541136(.A(n_310518882), .B(n_352265811), .C(n_312662130)
		, .D(n_352865817), .Z(n_318276021));
	notech_ao4 i_113441137(.A(n_351765806), .B(n_29172), .C(n_351165800), .D
		(n_27588), .Z(n_318476023));
	notech_ao4 i_113141140(.A(n_55143), .B(nbus_11273[21]), .C(n_54148), .D(\nbus_11276[21] 
		), .Z(n_318676025));
	notech_and4 i_113341138(.A(n_318676025), .B(n_26416), .C(n_284675685), .D
		(n_284975688), .Z(n_318976028));
	notech_ao4 i_112741144(.A(n_310618883), .B(n_352265811), .C(n_315162155)
		, .D(n_352865817), .Z(n_319076029));
	notech_ao4 i_112641145(.A(n_351765806), .B(n_29169), .C(n_351165800), .D
		(n_27586), .Z(n_319276031));
	notech_ao4 i_112341148(.A(n_55143), .B(nbus_11273[20]), .C(n_54148), .D(\nbus_11276[20] 
		), .Z(n_319476033));
	notech_and4 i_112541146(.A(n_319476033), .B(n_283775676), .C(n_284075679
		), .D(n_26491), .Z(n_319776036));
	notech_ao4 i_111941152(.A(n_310718884), .B(n_352265811), .C(n_308065397)
		, .D(n_352865817), .Z(n_319876037));
	notech_ao4 i_111841153(.A(n_351765806), .B(n_29167), .C(n_351165800), .D
		(n_27585), .Z(n_320076039));
	notech_ao4 i_111541156(.A(n_55143), .B(nbus_11273[19]), .C(n_54148), .D(\nbus_11276[19] 
		), .Z(n_320276041));
	notech_and4 i_111741154(.A(n_320276041), .B(n_26417), .C(n_282875667), .D
		(n_283175670), .Z(n_320576044));
	notech_ao4 i_111141160(.A(n_310818885), .B(n_352265811), .C(n_310565422)
		, .D(n_352865817), .Z(n_320676045));
	notech_ao4 i_111041161(.A(n_351765806), .B(n_29165), .C(n_351165800), .D
		(n_27584), .Z(n_320876047));
	notech_ao4 i_110741164(.A(n_55143), .B(nbus_11273[18]), .C(n_54148), .D(\nbus_11276[18] 
		), .Z(n_321076049));
	notech_and4 i_110941162(.A(n_321076049), .B(n_26492), .C(n_281975658), .D
		(n_282275661), .Z(n_321376052));
	notech_mux2 i_1511672(.S(n_60138), .A(n_570), .B(add_len_pc32[14]), .Z(\add_len_pc[14] 
		));
	notech_or2 i_82238300(.A(n_271888737), .B(n_55264), .Z(n_323276071));
	notech_nand2 i_82038302(.A(sav_epc[14]), .B(n_60595), .Z(n_323976078));
	notech_nand2 i_82138301(.A(\add_len_pc[14] ), .B(n_55819), .Z(n_324076079
		));
	notech_or4 i_82338299(.A(n_56104), .B(n_205088863), .C(n_55940), .D(n_272188734
		), .Z(n_324176080));
	notech_nand3 i_1520634(.A(n_340576242), .B(n_323276071), .C(n_340476241)
		, .Z(n_20195));
	notech_nor2 i_84038282(.A(n_101213406), .B(n_271988736), .Z(n_324476083)
		);
	notech_or4 i_84838274(.A(n_56196), .B(n_56158), .C(n_56376), .D(n_27582)
		, .Z(n_325276091));
	notech_nao3 i_85138271(.A(opc_10[16]), .B(n_62417), .C(n_306621953), .Z(n_325376092
		));
	notech_nor2 i_85038272(.A(n_272088735), .B(n_309921986), .Z(n_325476093)
		);
	notech_nor2 i_84938273(.A(n_55396), .B(n_271988736), .Z(n_325576094));
	notech_or4 i_1720668(.A(n_82113215), .B(n_325476093), .C(n_325576094), .D
		(n_26389), .Z(n_19881));
	notech_or2 i_1455283(.A(n_151860600), .B(n_163674504), .Z(n_325676095)
		);
	notech_or2 i_1155286(.A(n_151860600), .B(n_55987), .Z(n_325776096));
	notech_nao3 i_87738249(.A(n_62423), .B(opc[14]), .C(n_325676095), .Z(n_326276101
		));
	notech_nao3 i_87838248(.A(opc_10[14]), .B(n_62417), .C(n_325776096), .Z(n_326376102
		));
	notech_nor2 i_87638250(.A(n_54445), .B(n_271888737), .Z(n_326476103));
	notech_nor2 i_87938247(.A(n_80913203), .B(n_55965), .Z(n_326576104));
	notech_or4 i_1520666(.A(n_5990), .B(n_326476103), .C(n_26391), .D(n_326576104
		), .Z(n_19869));
	notech_or4 i_89438234(.A(n_204788866), .B(n_56158), .C(n_56375), .D(n_27582
		), .Z(n_327076109));
	notech_nao3 i_89738231(.A(opc_10[16]), .B(n_62417), .C(n_2694), .Z(n_327176110
		));
	notech_nor2 i_89638232(.A(n_2674), .B(n_272088735), .Z(n_327276111));
	notech_nor2 i_89538233(.A(n_271988736), .B(n_2655), .Z(n_327376112));
	notech_or4 i_1720732(.A(n_82113215), .B(n_327276111), .C(n_327376112), .D
		(n_26393), .Z(n_19533));
	notech_or4 i_133960569(.A(n_56465), .B(n_56431), .C(n_137574243), .D(n_29010
		), .Z(n_327476113));
	notech_or4 i_133160571(.A(n_56465), .B(n_56431), .C(n_29010), .D(n_55986
		), .Z(n_327576114));
	notech_nao3 i_91538217(.A(n_62409), .B(opc[14]), .C(n_327476113), .Z(n_328076119
		));
	notech_nao3 i_91838216(.A(opc_10[14]), .B(n_62417), .C(n_327576114), .Z(n_328176120
		));
	notech_nor2 i_91338218(.A(n_2656), .B(n_271888737), .Z(n_328276121));
	notech_nor2 i_92138215(.A(n_56139), .B(n_80913203), .Z(n_328376122));
	notech_or4 i_1520730(.A(n_5990), .B(n_328276121), .C(n_26394), .D(n_328376122
		), .Z(n_19521));
	notech_nor2 i_97538168(.A(n_353165820), .B(n_28987), .Z(n_328476123));
	notech_or4 i_98238161(.A(n_204788866), .B(n_56074), .C(n_55794), .D(n_2648
		), .Z(n_328576124));
	notech_or4 i_97938164(.A(n_204788866), .B(n_56074), .C(n_56363), .D(n_27583
		), .Z(n_328676125));
	notech_nor2 i_98038163(.A(n_121623203), .B(nbus_11326[17]), .Z(n_328776126
		));
	notech_ao3 i_98138162(.A(opc_10[17]), .B(n_62417), .C(n_121723204), .Z(n_328876127
		));
	notech_nor2 i_97838165(.A(n_2700), .B(n_353365822), .Z(n_328976128));
	notech_and2 i_97638167(.A(opb[17]), .B(n_353065819), .Z(n_329076129));
	notech_nor2 i_97738166(.A(n_353265821), .B(nbus_11273[17]), .Z(n_329176130
		));
	notech_or4 i_1820957(.A(n_329076129), .B(n_344376279), .C(n_329176130), 
		.D(n_328476123), .Z(n_9081));
	notech_nor2 i_99138152(.A(n_353165820), .B(n_29004), .Z(n_329276131));
	notech_or2 i_99638147(.A(n_121623203), .B(nbus_11326[16]), .Z(n_329476133
		));
	notech_ao3 i_99738146(.A(opc_10[16]), .B(n_62431), .C(n_121723204), .Z(n_329576134
		));
	notech_nor2 i_99838145(.A(n_121523202), .B(n_272088735), .Z(n_329676135)
		);
	notech_nor2 i_99538148(.A(n_271988736), .B(n_353365822), .Z(n_329776136)
		);
	notech_and2 i_99238151(.A(opb[16]), .B(n_353065819), .Z(n_329876137));
	notech_nor2 i_99338150(.A(n_353265821), .B(nbus_11273[16]), .Z(n_329976138
		));
	notech_or4 i_1720956(.A(n_329876137), .B(n_345076286), .C(n_329976138), 
		.D(n_329276131), .Z(n_9075));
	notech_or4 i_110838038(.A(n_56196), .B(n_58656), .C(n_56363), .D(n_27582
		), .Z(n_330476143));
	notech_nao3 i_111138035(.A(opc_10[16]), .B(n_62415), .C(n_308418861), .Z
		(n_330576144));
	notech_nor2 i_111038036(.A(n_272088735), .B(n_309618873), .Z(n_330676145
		));
	notech_nor2 i_110938037(.A(n_55404), .B(n_271988736), .Z(n_330776146));
	notech_or4 i_1720988(.A(n_82113215), .B(n_330676145), .C(n_330776146), .D
		(n_26396), .Z(n_16795));
	notech_or2 i_136337789(.A(n_55218), .B(\nbus_11276[17] ), .Z(n_331476153
		));
	notech_or2 i_136437788(.A(n_55554), .B(n_2700), .Z(n_331576154));
	notech_nand3 i_1821597(.A(n_346576301), .B(n_43426147), .C(n_331576154),
		 .Z(n_13217));
	notech_or4 i_137737775(.A(n_56158), .B(n_206288851), .C(n_56363), .D(n_27582
		), .Z(n_332076159));
	notech_nao3 i_138037772(.A(opc_10[16]), .B(n_62431), .C(n_308718864), .Z
		(n_332176160));
	notech_nor2 i_137937773(.A(n_272088735), .B(n_309518872), .Z(n_332276161
		));
	notech_nor2 i_137837774(.A(n_55554), .B(n_271988736), .Z(n_332376162));
	notech_or4 i_1721596(.A(n_82113215), .B(n_332276161), .C(n_332376162), .D
		(n_26397), .Z(n_13211));
	notech_or2 i_146537690(.A(n_55556), .B(n_2700), .Z(n_333176170));
	notech_nand3 i_1821853(.A(n_348076316), .B(n_333176170), .C(n_43426147),
		 .Z(n_12503));
	notech_or4 i_147937676(.A(n_56074), .B(n_206288851), .C(n_56363), .D(n_27582
		), .Z(n_333676175));
	notech_nao3 i_148237673(.A(opc_10[16]), .B(n_62431), .C(n_322931616), .Z
		(n_333776176));
	notech_nor2 i_148137674(.A(n_272088735), .B(n_322631613), .Z(n_333876177
		));
	notech_nor2 i_148037675(.A(n_55556), .B(n_271988736), .Z(n_333976178));
	notech_or4 i_1721852(.A(n_82113215), .B(n_333876177), .C(n_333976178), .D
		(n_26398), .Z(n_12497));
	notech_nand2 i_162237533(.A(add_src[15]), .B(n_26579), .Z(n_335076189)
		);
	notech_or2 i_162337532(.A(n_356476400), .B(n_2320), .Z(n_335176190));
	notech_or4 i_162537530(.A(n_260988754), .B(n_260888755), .C(n_2318), .D(n_28845
		), .Z(n_335476193));
	notech_nand3 i_1616185(.A(n_350476340), .B(n_349076326), .C(n_348976325)
		, .Z(n_14182));
	notech_or2 i_221036952(.A(n_351865807), .B(n_2700), .Z(n_336776204));
	notech_nand3 i_1817244(.A(n_351276348), .B(n_43426147), .C(n_336776204),
		 .Z(n_15876));
	notech_nao3 i_222836934(.A(opc_10[16]), .B(n_62431), .C(n_352865817), .Z
		(n_337476211));
	notech_nor2 i_222736935(.A(n_352265811), .B(n_272088735), .Z(n_337576212
		));
	notech_nor2 i_222636936(.A(n_271988736), .B(n_351865807), .Z(n_337676213
		));
	notech_or4 i_1717243(.A(n_337576212), .B(n_337676213), .C(n_82113215), .D
		(n_26400), .Z(n_15870));
	notech_ao4 i_22238871(.A(n_56240), .B(n_27730), .C(n_2261), .D(n_29206),
		 .Z(n_337776214));
	notech_ao4 i_22338870(.A(n_56178), .B(n_28000), .C(n_197114365), .D(n_27833
		), .Z(n_337876215));
	notech_ao4 i_22438869(.A(n_56415), .B(n_27968), .C(n_57343), .D(n_27764)
		, .Z(n_338076217));
	notech_ao4 i_22538868(.A(n_56182), .B(n_27934), .C(n_56310), .D(n_27621)
		, .Z(n_338176218));
	notech_and4 i_23538859(.A(n_338176218), .B(n_338076217), .C(n_337876215)
		, .D(n_337776214), .Z(n_338376220));
	notech_ao4 i_22638867(.A(n_60484), .B(n_27902), .C(n_56183), .D(n_29205)
		, .Z(n_338476221));
	notech_ao4 i_22838866(.A(n_56186), .B(n_27866), .C(n_56290), .D(n_27658)
		, .Z(n_338576222));
	notech_and2 i_23338861(.A(n_338576222), .B(n_338476221), .Z(n_338676223)
		);
	notech_ao4 i_22938865(.A(n_59224), .B(n_28034), .C(n_56270), .D(n_27698)
		, .Z(n_338776224));
	notech_ao4 i_23038864(.A(n_2262), .B(n_27801), .C(n_57373), .D(n_27385),
		 .Z(n_338876225));
	notech_and2 i_95260674(.A(n_55069), .B(n_2654), .Z(n_339176228));
	notech_and2 i_95160675(.A(n_55068), .B(n_2649), .Z(n_339276229));
	notech_and2 i_60060704(.A(n_55717), .B(n_137674244), .Z(n_339376230));
	notech_and2 i_95455344(.A(n_55487), .B(n_55071), .Z(n_339476231));
	notech_and2 i_95355345(.A(n_55070), .B(n_55488), .Z(n_339576232));
	notech_and2 i_59955358(.A(n_55719), .B(n_165074518), .Z(n_339676233));
	notech_ao4 i_82638296(.A(n_354269312), .B(n_55566), .C(n_55263), .D(n_29006
		), .Z(n_339776234));
	notech_ao4 i_82738295(.A(n_353969310), .B(n_27579), .C(n_56757), .D(n_26434
		), .Z(n_339976236));
	notech_ao4 i_82838294(.A(n_58922), .B(n_29375), .C(n_55492), .D(n_27533)
		, .Z(n_340076237));
	notech_and4 i_83138291(.A(n_340076237), .B(n_339976236), .C(n_339776234)
		, .D(n_323976078), .Z(n_340276239));
	notech_and3 i_83338289(.A(n_340276239), .B(n_324076079), .C(n_324176080)
		, .Z(n_340476241));
	notech_ao4 i_83438288(.A(n_354369313), .B(n_82713221), .C(n_354469314), 
		.D(n_82813222), .Z(n_340576242));
	notech_ao4 i_84138281(.A(\nbus_11276[16] ), .B(n_56216), .C(n_56775), .D
		(n_98113375), .Z(n_340776244));
	notech_ao4 i_84238280(.A(n_59856), .B(n_27535), .C(n_101413408), .D(n_29004
		), .Z(n_340876245));
	notech_nand2 i_84338279(.A(n_340876245), .B(n_340776244), .Z(n_340976246
		));
	notech_or2 i_67339080(.A(n_324476083), .B(n_340976246), .Z(n_82113215)
		);
	notech_ao4 i_85338269(.A(n_55397), .B(n_29004), .C(\nbus_11276[16] ), .D
		(n_55071), .Z(n_341076247));
	notech_ao4 i_85238270(.A(n_55070), .B(n_56775), .C(n_303521922), .D(nbus_11326
		[16]), .Z(n_341176248));
	notech_and4 i_85638266(.A(n_325276091), .B(n_341176248), .C(n_341076247)
		, .D(n_325376092), .Z(n_341476251));
	notech_ao4 i_88038246(.A(n_339476231), .B(n_55566), .C(n_54433), .D(n_29006
		), .Z(n_341776254));
	notech_ao4 i_88138245(.A(n_339676233), .B(n_27579), .C(n_339576232), .D(n_56757
		), .Z(n_341876255));
	notech_and4 i_88438242(.A(n_341876255), .B(n_341776254), .C(n_326276101)
		, .D(n_326376102), .Z(n_342176258));
	notech_ao4 i_89938229(.A(n_29004), .B(n_26444), .C(n_55069), .D(n_55590)
		, .Z(n_342576261));
	notech_ao4 i_89838230(.A(n_55068), .B(n_56775), .C(n_2672), .D(nbus_11326
		[16]), .Z(n_342676262));
	notech_and4 i_90238226(.A(n_327076109), .B(n_342676262), .C(n_342576261)
		, .D(n_327176110), .Z(n_342976265));
	notech_ao4 i_92238214(.A(n_339176228), .B(n_55566), .C(n_2653), .D(n_29006
		), .Z(n_343276268));
	notech_ao4 i_92438213(.A(n_339376230), .B(n_27579), .C(n_339276229), .D(n_56757
		), .Z(n_343376269));
	notech_and4 i_92738210(.A(n_343376269), .B(n_343276268), .C(n_328076119)
		, .D(n_328176120), .Z(n_343676272));
	notech_nand3 i_98438159(.A(n_272488731), .B(n_328576124), .C(n_328676125
		), .Z(n_344076276));
	notech_or4 i_98738156(.A(n_328776126), .B(n_344076276), .C(n_328876127),
		 .D(n_328976128), .Z(n_344376279));
	notech_ao4 i_99938144(.A(n_59856), .B(n_27535), .C(n_353465823), .D(n_27582
		), .Z(n_344676282));
	notech_nand2 i_100038143(.A(n_344676282), .B(n_329476133), .Z(n_344776283
		));
	notech_or4 i_100338140(.A(n_329576134), .B(n_344776283), .C(n_329676135)
		, .D(n_329776136), .Z(n_345076286));
	notech_ao4 i_111338033(.A(n_55405), .B(n_29004), .C(n_55062), .D(n_55590
		), .Z(n_345376289));
	notech_ao4 i_111238034(.A(n_55064), .B(n_56775), .C(n_55424), .D(n_58987
		), .Z(n_345476290));
	notech_and4 i_111638030(.A(n_330476143), .B(n_345476290), .C(n_345376289
		), .D(n_330576144), .Z(n_345776293));
	notech_ao4 i_136537787(.A(n_308318860), .B(nbus_11326[17]), .C(n_63826342
		), .D(n_308718864), .Z(n_346076296));
	notech_ao4 i_136637786(.A(n_2648), .B(n_309518872), .C(n_55773), .D(n_27583
		), .Z(n_346276298));
	notech_ao4 i_136737785(.A(n_55219), .B(nbus_11273[17]), .C(n_55555), .D(n_28987
		), .Z(n_346376299));
	notech_and4 i_137037782(.A(n_346376299), .B(n_346276298), .C(n_346076296
		), .D(n_331476153), .Z(n_346576301));
	notech_ao4 i_138237770(.A(n_55555), .B(n_29004), .C(n_55218), .D(n_55590
		), .Z(n_346776303));
	notech_ao4 i_138137771(.A(n_55219), .B(n_56775), .C(n_308318860), .D(n_58987
		), .Z(n_346876304));
	notech_and4 i_138537767(.A(n_346876304), .B(n_346776303), .C(n_332076159
		), .D(n_332176160), .Z(n_347176307));
	notech_ao4 i_146637689(.A(n_1031), .B(n_59945), .C(n_322931616), .D(n_63826342
		), .Z(n_347476310));
	notech_ao4 i_146737688(.A(n_55772), .B(n_27583), .C(n_303421921), .D(nbus_11326
		[17]), .Z(n_347576311));
	notech_ao4 i_146837687(.A(n_55557), .B(n_28987), .C(n_2648), .D(n_322631613
		), .Z(n_347776313));
	notech_ao4 i_146937686(.A(n_55221), .B(\nbus_11276[17] ), .C(n_55220), .D
		(nbus_11273[17]), .Z(n_347876314));
	notech_and4 i_147237683(.A(n_347876314), .B(n_347776313), .C(n_347576311
		), .D(n_347476310), .Z(n_348076316));
	notech_ao4 i_148437671(.A(n_55557), .B(n_29004), .C(n_55221), .D(n_55590
		), .Z(n_348276318));
	notech_ao4 i_148337672(.A(n_55220), .B(n_56775), .C(n_303421921), .D(n_58987
		), .Z(n_348376319));
	notech_and4 i_148737668(.A(n_333676175), .B(n_348376319), .C(n_348276318
		), .D(n_333776176), .Z(n_348676322));
	notech_ao4 i_164437511(.A(n_89713291), .B(n_28594), .C(n_89513289), .D(n_27601
		), .Z(n_348976325));
	notech_ao4 i_164237513(.A(n_272288733), .B(n_55578), .C(n_88813282), .D(n_28411
		), .Z(n_349076326));
	notech_ao4 i_163437521(.A(n_55526), .B(n_28593), .C(n_55366), .D(n_28789
		), .Z(n_349176327));
	notech_and4 i_163837517(.A(n_330946790), .B(n_349176327), .C(n_54719), .D
		(n_335076189), .Z(n_349476330));
	notech_ao4 i_163037525(.A(n_54884), .B(n_56943), .C(n_54735), .D(nbus_11326
		[7]), .Z(n_349576331));
	notech_ao4 i_163137524(.A(n_2156), .B(n_28816), .C(n_2323), .D(n_27581),
		 .Z(n_349676332));
	notech_ao4 i_163237523(.A(n_2319), .B(n_29031), .C(n_2322), .D(n_56766),
		 .Z(n_349876334));
	notech_ao4 i_163337522(.A(n_55243), .B(n_27534), .C(n_2164), .D(nbus_11326
		[15]), .Z(n_349976335));
	notech_and4 i_163937516(.A(n_349976335), .B(n_349876334), .C(n_349676332
		), .D(n_349576331), .Z(n_350176337));
	notech_and4 i_164337512(.A(n_350176337), .B(n_349476330), .C(n_335176190
		), .D(n_335476193), .Z(n_350476340));
	notech_ao4 i_221136951(.A(n_352865817), .B(n_63826342), .C(n_107626780),
		 .D(n_28711), .Z(n_350676342));
	notech_ao4 i_221236950(.A(n_351165800), .B(n_27583), .C(n_351665805), .D
		(nbus_11326[17]), .Z(n_350776343));
	notech_ao4 i_221336949(.A(n_351765806), .B(n_28987), .C(n_352265811), .D
		(n_2648), .Z(n_350976345));
	notech_ao4 i_221436948(.A(n_54148), .B(\nbus_11276[17] ), .C(n_55143), .D
		(nbus_11273[17]), .Z(n_351076346));
	notech_and4 i_221736945(.A(n_351076346), .B(n_350976345), .C(n_350776343
		), .D(n_350676342), .Z(n_351276348));
	notech_ao4 i_223136931(.A(n_351165800), .B(n_27582), .C(n_351765806), .D
		(n_29004), .Z(n_351476350));
	notech_ao4 i_222936933(.A(n_351665805), .B(n_58987), .C(n_107626780), .D
		(n_28710), .Z(n_351576351));
	notech_ao4 i_223036932(.A(n_54148), .B(n_55590), .C(n_55143), .D(n_56775
		), .Z(n_351676352));
	notech_and4 i_223436928(.A(n_351676352), .B(n_351576351), .C(n_351476350
		), .D(n_337476211), .Z(n_351976355));
	notech_or4 i_5935639(.A(n_272588730), .B(n_273188724), .C(n_59945), .D(n_55578
		), .Z(n_352276358));
	notech_nand3 i_72332887(.A(n_205988854), .B(n_2182), .C(n_354476380), .Z
		(n_352376359));
	notech_and2 i_15232727(.A(n_354376379), .B(n_2823), .Z(n_352476360));
	notech_and4 i_15332726(.A(n_2236), .B(n_354276378), .C(n_55843), .D(n_354676382
		), .Z(n_352576361));
	notech_and2 i_45832489(.A(n_2107), .B(n_54689), .Z(n_352676362));
	notech_nor2 i_45932488(.A(n_2265), .B(n_613), .Z(n_352776363));
	notech_or4 i_27432648(.A(n_2647), .B(n_59370), .C(n_272788728), .D(n_60474
		), .Z(n_353176367));
	notech_or4 i_27332649(.A(n_26862), .B(n_59159), .C(n_26497), .D(write_ack
		), .Z(n_353476370));
	notech_or4 i_28463(.A(n_2793), .B(n_26629), .C(n_59159), .D(n_29130), .Z
		(n_353776373));
	notech_nao3 i_145431662(.A(n_27566), .B(n_27565), .C(opd[2]), .Z(n_353976375
		));
	notech_ao4 i_6732797(.A(n_2647), .B(n_2179), .C(n_273388722), .D(n_26600
		), .Z(n_354276378));
	notech_ao4 i_137732848(.A(n_57458), .B(n_57441), .C(read_ack), .D(n_2824
		), .Z(n_354376379));
	notech_ao4 i_118231897(.A(n_2209), .B(n_352676362), .C(n_55280), .D(n_60474
		), .Z(n_354476380));
	notech_and3 i_81032217(.A(n_57380), .B(n_57423), .C(n_57414), .Z(n_354676382
		));
	notech_ao4 i_80632221(.A(n_60474), .B(n_352576361), .C(n_494), .D(n_352476360
		), .Z(n_354976385));
	notech_and4 i_80832219(.A(n_1914), .B(n_353176367), .C(n_354976385), .D(n_353476370
		), .Z(n_355276388));
	notech_or4 i_80332224(.A(n_26620), .B(n_26543), .C(n_26420), .D(n_352376359
		), .Z(n_355476390));
	notech_or4 i_16741(.A(n_170914103), .B(n_2793), .C(n_2823), .D(n_29130),
		 .Z(n_355776393));
	notech_nand3 i_54889(.A(n_55642), .B(n_125874126), .C(n_1918), .Z(\nbus_11354[0] 
		));
	notech_ao3 i_173861856(.A(n_167260754), .B(n_167060752), .C(n_167160753)
		, .Z(n_197061044));
	notech_and4 i_820659(.A(n_132574193), .B(n_132774195), .C(n_133174199), 
		.D(n_131974187), .Z(n_19827));
	notech_and4 i_820723(.A(n_133274200), .B(n_133474202), .C(n_133874206), 
		.D(n_131174179), .Z(n_19479));
	notech_and4 i_720722(.A(n_133974207), .B(n_134174209), .C(n_134574213), 
		.D(n_130374171), .Z(n_19473));
	notech_and4 i_520720(.A(n_134674214), .B(n_134874216), .C(n_135274220), 
		.D(n_129574163), .Z(n_19461));
	notech_and4 i_820947(.A(n_135374221), .B(n_135574223), .C(n_135974227), 
		.D(n_128774155), .Z(n_9021));
	notech_and4 i_720946(.A(n_136074228), .B(n_136274230), .C(n_136674234), 
		.D(n_127974147), .Z(n_9015));
	notech_and4 i_520944(.A(n_136774235), .B(n_136974237), .C(n_137374241), 
		.D(n_127174139), .Z(n_9003));
	notech_or2 i_191163545(.A(n_151860600), .B(n_126274130), .Z(n_279739585)
		);
	notech_or2 i_4163506(.A(n_151860600), .B(n_56005), .Z(n_275539543));
	notech_and3 i_182563589(.A(n_55071), .B(n_126174129), .C(n_54445), .Z(n_54655
		));
	notech_ao3 i_182463590(.A(n_55070), .B(n_54433), .C(n_126074128), .Z(n_54656
		));
	notech_and2 i_59363600(.A(n_55719), .B(n_126374131), .Z(n_55756));
	notech_ao4 i_174361851(.A(n_263436789), .B(n_182360897), .C(n_148160563)
		, .D(n_145860540), .Z(n_196861042));
	notech_or4 i_174461850(.A(n_54528), .B(instrc[124]), .C(instrc[126]), .D
		(n_60563), .Z(n_196761041));
	notech_ao3 i_150360654(.A(n_54853), .B(n_55220), .C(n_47685), .Z(n_54923
		));
	notech_and3 i_150460653(.A(n_54852), .B(n_47687), .C(n_55221), .Z(n_54922
		));
	notech_and4 i_189860639(.A(n_55658), .B(n_238758633), .C(n_322288468), .D
		(n_323388457), .Z(n_54594));
	notech_and3 i_193760630(.A(n_97522962), .B(n_355976395), .C(n_356176397)
		, .Z(n_54562));
	notech_and2 i_195560622(.A(n_128967109), .B(n_356076396), .Z(n_54547));
	notech_and4 i_3020681(.A(n_262736782), .B(n_144874316), .C(n_143674304),
		 .D(n_144774315), .Z(n_19959));
	notech_or4 i_920660(.A(n_145974327), .B(n_26324), .C(n_145474322), .D(n_26323
		), .Z(n_19833));
	notech_and4 i_3020745(.A(n_262736782), .B(n_146674334), .C(n_141574283),
		 .D(n_146574333), .Z(n_19611));
	notech_or4 i_1020725(.A(n_185167671), .B(n_140874276), .C(n_147274340), 
		.D(n_26325), .Z(n_19491));
	notech_and4 i_920724(.A(n_147674344), .B(n_147874346), .C(n_140774275), 
		.D(n_148274350), .Z(n_19485));
	notech_nand2 i_521168(.A(n_149374361), .B(n_148874356), .Z(n_13491));
	notech_and4 i_821555(.A(n_138174249), .B(n_149974367), .C(n_150274370), 
		.D(n_149874366), .Z(n_16392));
	notech_nao3 i_137560562(.A(n_56487), .B(n_268064997), .C(n_55976), .Z(n_259336748
		));
	notech_ao4 i_173961855(.A(n_196361037), .B(n_183160905), .C(n_196261036)
		, .D(n_179960880), .Z(n_196461038));
	notech_nand3 i_174661848(.A(n_29034), .B(n_28972), .C(n_29026), .Z(n_196361037
		));
	notech_nao3 i_174761847(.A(n_29032), .B(n_28970), .C(n_176360845), .Z(n_196261036
		));
	notech_ao4 i_174061854(.A(n_196061034), .B(n_190460978), .C(n_195961033)
		, .D(n_194061014), .Z(n_196161035));
	notech_nand2 i_174861846(.A(n_29019), .B(n_29022), .Z(n_196061034));
	notech_nao3 i_174961845(.A(n_29033), .B(n_26528), .C(instrc[102]), .Z(n_195961033
		));
	notech_and4 i_175661838(.A(n_54769), .B(n_195661030), .C(n_195461028), .D
		(n_195361027), .Z(n_195861032));
	notech_nand2 i_62157979(.A(n_55772), .B(n_151274380), .Z(n_55729));
	notech_ao4 i_175161843(.A(n_184760921), .B(n_1529), .C(n_191060984), .D(n_1916
		), .Z(n_195661030));
	notech_and2 i_80557919(.A(n_57375), .B(n_57376), .Z(n_55546));
	notech_and4 i_820979(.A(n_157674444), .B(n_158174449), .C(n_158374451), 
		.D(n_158874456), .Z(n_16741));
	notech_nand2 i_821299(.A(n_159874466), .B(n_159374461), .Z(n_20643));
	notech_and4 i_521296(.A(n_154974417), .B(n_160374471), .C(n_160574473), 
		.D(n_160274470), .Z(n_20625));
	notech_and4 i_821587(.A(n_154474412), .B(n_160774475), .C(n_160974477), 
		.D(n_161374481), .Z(n_13157));
	notech_and4 i_821843(.A(n_161474482), .B(n_161674484), .C(n_162074488), 
		.D(n_153674404), .Z(n_12443));
	notech_and4 i_721842(.A(n_162174489), .B(n_162374491), .C(n_162874496), 
		.D(n_152874396), .Z(n_12437));
	notech_and4 i_521840(.A(n_162974497), .B(n_163174499), .C(n_163574503), 
		.D(n_152074388), .Z(n_12425));
	notech_or2 i_62657895(.A(n_252034146), .B(n_26599), .Z(n_251834144));
	notech_or2 i_63757894(.A(n_55820), .B(n_2675), .Z(n_251734143));
	notech_nao3 i_131657863(.A(n_56487), .B(n_268064997), .C(n_150774375), .Z
		(n_248634112));
	notech_ao4 i_188657853(.A(n_55854), .B(n_55400), .C(n_1135), .D(n_28983)
		, .Z(n_247634102));
	notech_ao4 i_175361841(.A(n_148060562), .B(n_1025), .C(n_185560929), .D(n_56183
		), .Z(n_195461028));
	notech_ao4 i_175461840(.A(n_56382), .B(n_148160563), .C(n_147960561), .D
		(n_146260544), .Z(n_195361027));
	notech_and4 i_175861836(.A(n_194961023), .B(n_146360545), .C(n_168660768
		), .D(n_168560767), .Z(n_195161025));
	notech_mux2 i_108955330(.S(opa[7]), .A(n_186274730), .B(n_186174729), .Z
		(n_55282));
	notech_mux2 i_112055329(.S(opa[31]), .A(n_186274730), .B(n_186174729), .Z
		(n_55252));
	notech_mux2 i_111955328(.S(opa[15]), .A(n_186274730), .B(n_186174729), .Z
		(n_55253));
	notech_or4 i_2520676(.A(n_252861556), .B(n_185374721), .C(n_186774735), 
		.D(n_26328), .Z(n_19929));
	notech_and4 i_1620667(.A(n_363088165), .B(n_184574713), .C(n_187574743),
		 .D(n_187474742), .Z(n_19875));
	notech_or4 i_1420665(.A(n_188774755), .B(n_183274700), .C(n_188274750), 
		.D(n_26329), .Z(n_19863));
	notech_or4 i_1320664(.A(n_189974767), .B(n_181974687), .C(n_189474762), 
		.D(n_26332), .Z(n_19857));
	notech_or4 i_1220663(.A(n_239168196), .B(n_181174679), .C(n_190574773), 
		.D(n_26333), .Z(n_19851));
	notech_or4 i_2520740(.A(n_252861556), .B(n_180374671), .C(n_191274780), 
		.D(n_26334), .Z(n_19581));
	notech_and4 i_1620731(.A(n_363088165), .B(n_192074788), .C(n_179574663),
		 .D(n_191974787), .Z(n_19527));
	notech_or4 i_1420729(.A(n_188774755), .B(n_178774655), .C(n_192674794), 
		.D(n_26335), .Z(n_19515));
	notech_or4 i_1320728(.A(n_189974767), .B(n_177974647), .C(n_193374801), 
		.D(n_26336), .Z(n_19509));
	notech_or4 i_1220727(.A(n_239168196), .B(n_177174639), .C(n_194074808), 
		.D(n_26337), .Z(n_19503));
	notech_nand3 i_1120726(.A(n_194674814), .B(n_194574813), .C(n_195074818)
		, .Z(n_19497));
	notech_nand3 i_1120950(.A(n_195374821), .B(n_195274820), .C(n_195774825)
		, .Z(n_9039));
	notech_or4 i_2520996(.A(n_252861556), .B(n_174874616), .C(n_196174829), 
		.D(n_26338), .Z(n_16843));
	notech_nand2 i_1621179(.A(n_197474842), .B(n_196974837), .Z(n_13557));
	notech_nand2 i_1321176(.A(n_198474852), .B(n_197974847), .Z(n_13539));
	notech_nand2 i_921172(.A(n_199474862), .B(n_198974857), .Z(n_13515));
	notech_nand3 i_1421305(.A(n_200074868), .B(n_199974867), .C(n_199874866)
		, .Z(n_20679));
	notech_nand2 i_1221303(.A(n_201374881), .B(n_200874876), .Z(n_20667));
	notech_or4 i_1421593(.A(n_188774755), .B(n_168174549), .C(n_201774885), 
		.D(n_26340), .Z(n_13193));
	notech_nand2 i_1121718(.A(n_203174899), .B(n_202674894), .Z(n_12827));
	notech_and4 i_1421849(.A(n_203274900), .B(n_203474902), .C(n_203974907),
		 .D(n_166774535), .Z(n_12479));
	notech_and4 i_2517251(.A(n_165974527), .B(n_204074908), .C(n_204274910),
		 .D(n_204774915), .Z(n_15918));
	notech_ao4 i_176361831(.A(n_1025), .B(n_182360897), .C(n_148160563), .D(n_146260544
		), .Z(n_194961023));
	notech_or4 i_176461830(.A(n_54527), .B(n_29032), .C(instrc[126]), .D(n_60563
		), .Z(n_194861022));
	notech_and4 i_176161833(.A(n_168760769), .B(n_168860770), .C(n_168960771
		), .D(n_169060772), .Z(n_194761021));
	notech_and3 i_252052056(.A(n_55667), .B(n_238958635), .C(n_34533), .Z(n_355876394
		));
	notech_nand2 i_12440(.A(n_322188469), .B(n_323488456), .Z(n_355976395)
		);
	notech_nand2 i_208752018(.A(n_26516), .B(n_26411), .Z(n_356076396));
	notech_nand2 i_210452017(.A(n_322188469), .B(n_26411), .Z(n_356176397)
		);
	notech_or4 i_28406(.A(n_56465), .B(n_355988238), .C(n_355876394), .D(n_29010
		), .Z(n_356276398));
	notech_or4 i_28409(.A(n_56465), .B(n_355988238), .C(n_323388457), .D(n_29010
		), .Z(n_356376399));
	notech_or4 i_205163587(.A(n_1916), .B(n_148560567), .C(n_56005), .D(n_59235
		), .Z(n_54469));
	notech_or2 i_209063585(.A(n_54523), .B(n_56005), .Z(n_54438));
	notech_nand3 i_2920680(.A(n_263775476), .B(n_263675475), .C(n_264175480)
		, .Z(n_19953));
	notech_nand3 i_2820679(.A(n_264375482), .B(n_264275481), .C(n_265175490)
		, .Z(n_19947));
	notech_nand3 i_2720678(.A(n_265375492), .B(n_265275491), .C(n_266175500)
		, .Z(n_19941));
	notech_nand3 i_2620677(.A(n_266375502), .B(n_266275501), .C(n_266775506)
		, .Z(n_19935));
	notech_or4 i_2420675(.A(n_267675515), .B(n_258575424), .C(n_267175510), 
		.D(n_26347), .Z(n_19923));
	notech_or4 i_2920744(.A(n_313168930), .B(n_257775416), .C(n_268275521), 
		.D(n_26348), .Z(n_19605));
	notech_or4 i_2820743(.A(n_264975488), .B(n_256975408), .C(n_268975528), 
		.D(n_26349), .Z(n_19599));
	notech_or4 i_2720742(.A(n_265975498), .B(n_256175400), .C(n_269675535), 
		.D(n_26350), .Z(n_19593));
	notech_or4 i_2620741(.A(n_173971058), .B(n_255375392), .C(n_270375542), 
		.D(n_26351), .Z(n_19587));
	notech_or4 i_2420739(.A(n_267675515), .B(n_254575384), .C(n_271075549), 
		.D(n_26352), .Z(n_19575));
	notech_or4 i_2921000(.A(n_313168930), .B(n_253775376), .C(n_271775556), 
		.D(n_26353), .Z(n_16867));
	notech_or4 i_2820999(.A(n_264975488), .B(n_252975368), .C(n_272475563), 
		.D(n_26354), .Z(n_16861));
	notech_or4 i_2720998(.A(n_265975498), .B(n_252175360), .C(n_273175570), 
		.D(n_26355), .Z(n_16855));
	notech_or4 i_2620997(.A(n_173971058), .B(n_251375352), .C(n_273875577), 
		.D(n_26356), .Z(n_16849));
	notech_or4 i_2420995(.A(n_267675515), .B(n_250575344), .C(n_274575584), 
		.D(n_26357), .Z(n_16837));
	notech_nand2 i_2921192(.A(n_275875597), .B(n_275375592), .Z(n_13635));
	notech_nand2 i_2721190(.A(n_276875607), .B(n_276375602), .Z(n_13623));
	notech_nand2 i_2621189(.A(n_277875617), .B(n_277375612), .Z(n_13617));
	notech_nand3 i_2921608(.A(n_278075619), .B(n_277975618), .C(n_278475623)
		, .Z(n_13283));
	notech_nand3 i_2821607(.A(n_278675625), .B(n_278575624), .C(n_279075629)
		, .Z(n_13277));
	notech_nand3 i_2721606(.A(n_279275631), .B(n_279175630), .C(n_279675635)
		, .Z(n_13271));
	notech_nand3 i_2621605(.A(n_279875637), .B(n_279775636), .C(n_280275641)
		, .Z(n_13265));
	notech_and4 i_2817254(.A(n_280375642), .B(n_280575644), .C(n_242875279),
		 .D(n_281075649), .Z(n_15936));
	notech_and4 i_2417250(.A(n_281175650), .B(n_281375652), .C(n_241775270),
		 .D(n_281875657), .Z(n_15912));
	notech_or2 i_43145380(.A(n_56363), .B(n_27594), .Z(n_307621963));
	notech_or2 i_3545342(.A(n_56369), .B(n_27595), .Z(n_303621923));
	notech_ao4 i_3145346(.A(n_56369), .B(n_27594), .C(n_308321970), .D(n_55794
		), .Z(n_304021927));
	notech_ao4 i_2645348(.A(n_56363), .B(n_27596), .C(n_57306), .D(n_55794),
		 .Z(n_304221929));
	notech_nand2 i_176961825(.A(instrc[103]), .B(n_29025), .Z(n_194061014)
		);
	notech_ao3 i_177261822(.A(n_169560777), .B(n_193861012), .C(n_169460776)
		, .Z(n_193961013));
	notech_and4 i_2320674(.A(n_303675875), .B(n_303275871), .C(n_301675855),
		 .D(n_303175870), .Z(n_19917));
	notech_or4 i_2220673(.A(n_304775886), .B(n_300475843), .C(n_304275881), 
		.D(n_26358), .Z(n_19911));
	notech_or4 i_2120672(.A(n_320179591), .B(n_299675835), .C(n_305375892), 
		.D(n_26359), .Z(n_19905));
	notech_or4 i_2020671(.A(n_306575904), .B(n_298475823), .C(n_306075899), 
		.D(n_26360), .Z(n_19899));
	notech_or4 i_1920670(.A(n_320579595), .B(n_297675815), .C(n_307175910), 
		.D(n_26363), .Z(n_19893));
	notech_and4 i_2320738(.A(n_303675875), .B(n_307975918), .C(n_296875807),
		 .D(n_307875917), .Z(n_19569));
	notech_or4 i_2220737(.A(n_304775886), .B(n_296075799), .C(n_308575924), 
		.D(n_26364), .Z(n_19563));
	notech_or4 i_2120736(.A(n_320179591), .B(n_295275791), .C(n_309275931), 
		.D(n_26365), .Z(n_19557));
	notech_or4 i_2020735(.A(n_306575904), .B(n_294475783), .C(n_309975938), 
		.D(n_26366), .Z(n_19551));
	notech_or4 i_1920734(.A(n_320579595), .B(n_293675775), .C(n_310675945), 
		.D(n_26368), .Z(n_19545));
	notech_nand3 i_2320962(.A(n_311575954), .B(n_311475953), .C(n_311375952)
		, .Z(n_9111));
	notech_and4 i_2320994(.A(n_303675875), .B(n_312175960), .C(n_292075759),
		 .D(n_312075959), .Z(n_16831));
	notech_or4 i_2220993(.A(n_304775886), .B(n_291275751), .C(n_312775966), 
		.D(n_26370), .Z(n_16825));
	notech_or4 i_2120992(.A(n_320179591), .B(n_290475743), .C(n_313475973), 
		.D(n_26371), .Z(n_16819));
	notech_or4 i_2020991(.A(n_306575904), .B(n_289675735), .C(n_314175980), 
		.D(n_26372), .Z(n_16813));
	notech_or4 i_1920990(.A(n_320579595), .B(n_288875727), .C(n_314875987), 
		.D(n_26373), .Z(n_16807));
	notech_and4 i_2321058(.A(n_303675875), .B(n_315675995), .C(n_288075719),
		 .D(n_315575994), .Z(n_13947));
	notech_and4 i_2321602(.A(n_303675875), .B(n_316376002), .C(n_287275711),
		 .D(n_316276001), .Z(n_13247));
	notech_and4 i_2321858(.A(n_316676005), .B(n_316876007), .C(n_317376012),
		 .D(n_287175710), .Z(n_12533));
	notech_and4 i_2317249(.A(n_317476013), .B(n_317676015), .C(n_318176020),
		 .D(n_286375702), .Z(n_15906));
	notech_and4 i_2217248(.A(n_318276021), .B(n_318476023), .C(n_285475693),
		 .D(n_318976028), .Z(n_15900));
	notech_and4 i_2117247(.A(n_319076029), .B(n_319276031), .C(n_284575684),
		 .D(n_319776036), .Z(n_15894));
	notech_and4 i_2017246(.A(n_319876037), .B(n_320076039), .C(n_283675675),
		 .D(n_320576044), .Z(n_15888));
	notech_and4 i_1917245(.A(n_320676045), .B(n_320876047), .C(n_282775666),
		 .D(n_321376052), .Z(n_15882));
	notech_nand2 i_165242237(.A(read_data[22]), .B(n_59945), .Z(n_308218859)
		);
	notech_nand2 i_165742235(.A(read_data[21]), .B(n_59944), .Z(n_308018857)
		);
	notech_ao4 i_177061824(.A(n_323688454), .B(n_60474), .C(n_56043), .D(n_148160563
		), .Z(n_193861012));
	notech_and4 i_92629150(.A(n_338876225), .B(n_338776224), .C(n_338376220)
		, .D(n_338676223), .Z(n_356476400));
	notech_ao4 i_177661818(.A(n_56186), .B(n_26524), .C(n_56100), .D(n_26523
		), .Z(n_193561009));
	notech_and2 i_32321(.A(n_54725), .B(n_352276358), .Z(n_330946790));
	notech_or4 i_153933167(.A(n_59159), .B(n_275388704), .C(n_273688719), .D
		(n_26418), .Z(n_54892));
	notech_or4 i_52734(.A(n_170914103), .B(n_2793), .C(n_55641), .D(n_29130)
		, .Z(n_57461));
	notech_ao3 i_5383(.A(sema_rw), .B(n_26590), .C(n_2222), .Z(n_51730));
	notech_ao4 i_177761817(.A(n_135360435), .B(n_26530), .C(n_170860790), .D
		(n_26538), .Z(n_193461008));
	notech_ao4 i_177961815(.A(n_170960791), .B(n_26525), .C(n_171060792), .D
		(n_26529), .Z(n_193261006));
	notech_nand2 i_7063477(.A(n_29033), .B(n_28971), .Z(n_193161005));
	notech_ao4 i_178061814(.A(n_171160793), .B(n_26532), .C(n_192961003), .D
		(n_192761001), .Z(n_193061004));
	notech_nand3 i_178661808(.A(n_182960903), .B(n_29034), .C(n_28972), .Z(n_192961003
		));
	notech_nand2 i_5263495(.A(n_29034), .B(n_28972), .Z(n_192861002));
	notech_nand2 i_178761807(.A(instrc[93]), .B(instrc[95]), .Z(n_192761001)
		);
	notech_or4 i_226952(.A(n_355476390), .B(n_51730), .C(n_26619), .D(n_26401
		), .Z(n_14902));
	notech_or4 i_1330759(.A(opd[0]), .B(opd[1]), .C(opd[3]), .D(n_353976375)
		, .Z(n_2265));
	notech_or2 i_5395(.A(n_2175), .B(n_352776363), .Z(n_2224));
	notech_ao4 i_178861806(.A(n_56100), .B(n_182360897), .C(n_148160563), .D
		(n_192260996), .Z(n_192560999));
	notech_and2 i_109132987(.A(n_2271), .B(n_2269), .Z(n_55280));
	notech_ao4 i_177361821(.A(n_147960561), .B(n_146560547), .C(n_191060984)
		, .D(n_191960993), .Z(n_192360997));
	notech_and2 i_4463503(.A(n_146960551), .B(n_54507), .Z(n_192260996));
	notech_nand3 i_179061804(.A(instrc[123]), .B(n_28566), .C(instrc[121]), 
		.Z(n_191960993));
	notech_nand2 i_112663549(.A(n_29032), .B(n_28970), .Z(n_191760991));
	notech_nao3 i_179561799(.A(n_26380), .B(n_2822), .C(n_353776373), .Z(n_191560989
		));
	notech_and4 i_180261793(.A(n_191160985), .B(n_190860982), .C(n_171860800
		), .D(n_172160803), .Z(n_191360987));
	notech_nand2 i_25187228(.A(over_seg[5]), .B(n_60138), .Z(n_56076));
	notech_ao4 i_179861797(.A(n_1913), .B(n_191060984), .C(n_148060562), .D(n_324669045
		), .Z(n_191160985));
	notech_or4 i_69263559(.A(tcmp), .B(n_1900), .C(n_60474), .D(n_60532), .Z
		(n_191060984));
	notech_ao4 i_180061795(.A(n_56009), .B(n_148160563), .C(n_147960561), .D
		(n_147160553), .Z(n_190860982));
	notech_ao4 i_180361792(.A(n_190260976), .B(n_190460978), .C(n_189960973)
		, .D(n_190160975), .Z(n_190560979));
	notech_nand3 i_15163400(.A(instrc[99]), .B(n_29013), .C(n_26531), .Z(n_190460978
		));
	notech_nand2 i_8963458(.A(instrc[96]), .B(instrc[97]), .Z(n_190260976)
		);
	notech_nand3 i_15463397(.A(instrc[88]), .B(n_184460918), .C(instrc[89]),
		 .Z(n_190160975));
	notech_nand2 i_7463473(.A(instrc[91]), .B(n_29014), .Z(n_189960973));
	notech_and2 i_7263475(.A(instrc[107]), .B(n_29008), .Z(n_189760971));
	notech_nand2 i_9363454(.A(instrc[104]), .B(instrc[105]), .Z(n_189660970)
		);
	notech_and4 i_180861788(.A(n_172560807), .B(n_172860810), .C(n_172760809
		), .D(n_26517), .Z(n_189560969));
	notech_ao4 i_181061786(.A(n_324669045), .B(n_182360897), .C(n_148160563)
		, .D(n_147160553), .Z(n_189360967));
	notech_nand2 i_6363484(.A(instrc[124]), .B(n_28970), .Z(n_188960963));
	notech_nand2 i_9263455(.A(instrc[92]), .B(n_28972), .Z(n_188660960));
	notech_nand2 i_11363436(.A(instrc[100]), .B(n_28971), .Z(n_188460958));
	notech_and4 i_181961777(.A(n_188160955), .B(n_187960953), .C(n_173360815
		), .D(n_173660818), .Z(n_188360957));
	notech_ao4 i_181561781(.A(n_148060562), .B(n_56101), .C(n_56310), .D(n_185560929
		), .Z(n_188160955));
	notech_ao4 i_181761779(.A(n_147960561), .B(n_147560557), .C(n_187860952)
		, .D(n_183960913), .Z(n_187960953));
	notech_nao3 i_14363408(.A(n_184460918), .B(n_29023), .C(instrc[88]), .Z(n_187860952
		));
	notech_ao3 i_182161775(.A(n_173860820), .B(n_173760819), .C(n_173960821)
		, .Z(n_187660950));
	notech_ao4 i_182861770(.A(n_56101), .B(n_182360897), .C(n_148160563), .D
		(n_147560557), .Z(n_187260946));
	notech_and4 i_182661772(.A(n_174160823), .B(n_174060822), .C(n_26522), .D
		(n_174260824), .Z(n_186960943));
	notech_and4 i_184161757(.A(n_186060934), .B(n_185060924), .C(n_174860830
		), .D(n_175160833), .Z(n_186260936));
	notech_ao4 i_183761761(.A(n_148060562), .B(n_151860600), .C(n_185560929)
		, .D(n_56178), .Z(n_186060934));
	notech_or2 i_14963402(.A(n_26523), .B(n_177860860), .Z(n_185960933));
	notech_and4 i_20363569(.A(n_56425), .B(n_179660877), .C(n_27557), .D(all_cnt
		[1]), .Z(n_185860932));
	notech_or2 i_119663548(.A(n_26524), .B(n_177860860), .Z(n_185560929));
	notech_and4 i_20263570(.A(n_176860850), .B(n_56415), .C(n_27557), .D(n_27556
		), .Z(n_185460928));
	notech_ao4 i_183961759(.A(n_147960561), .B(n_148260564), .C(n_183960913)
		, .D(n_184660920), .Z(n_185060924));
	notech_or2 i_22655(.A(tcmp), .B(n_135860440), .Z(n_184960923));
	notech_or2 i_65363560(.A(tcmp), .B(n_54865), .Z(n_184760921));
	notech_nand3 i_14863403(.A(n_184460918), .B(instrc[88]), .C(n_29023), .Z
		(n_184660920));
	notech_nor2 i_2063527(.A(n_177860860), .B(n_26525), .Z(n_184460918));
	notech_and4 i_20863564(.A(n_334962247), .B(all_cnt[1]), .C(all_cnt[2]), 
		.D(n_176860850), .Z(n_184360917));
	notech_nand2 i_8263465(.A(instrc[90]), .B(n_29017), .Z(n_184060914));
	notech_nand2 i_14463407(.A(instrc[90]), .B(instrc[91]), .Z(n_183960913)
		);
	notech_and4 i_184361755(.A(n_182460898), .B(n_175360835), .C(n_175260834
		), .D(n_148360565), .Z(n_183760911));
	notech_or4 i_9163456(.A(tcmp), .B(n_1900), .C(n_60474), .D(n_59235), .Z(n_183460908
		));
	notech_or4 i_6263485(.A(tcmp), .B(n_60595), .C(n_59944), .D(n_1900), .Z(n_183360907
		));
	notech_nand2 i_9463453(.A(n_183060904), .B(instrc[95]), .Z(n_183160905)
		);
	notech_and2 i_2263525(.A(n_182960903), .B(n_26535), .Z(n_183060904));
	notech_and4 i_20763565(.A(n_334662244), .B(n_179660877), .C(all_cnt[1]),
		 .D(all_cnt[2]), .Z(n_182960903));
	notech_and2 i_5963488(.A(instrc[94]), .B(n_29026), .Z(n_182660900));
	notech_ao4 i_185661742(.A(n_151860600), .B(n_182360897), .C(n_148260564)
		, .D(n_148160563), .Z(n_182460898));
	notech_or2 i_2563522(.A(n_181560891), .B(n_60512), .Z(n_182360897));
	notech_nao3 i_179663547(.A(instrc[126]), .B(n_62395), .C(instrc[125]), .Z
		(n_182060895));
	notech_ao4 i_186061738(.A(n_2263), .B(n_26384), .C(n_148560567), .D(n_26316
		), .Z(n_181860893));
	notech_or2 i_76763556(.A(tcmp), .B(n_135760439), .Z(n_181560891));
	notech_or4 i_184661752(.A(n_175760839), .B(n_175660838), .C(n_26527), .D
		(n_175560837), .Z(n_181160889));
	notech_nand2 i_2363524(.A(n_180460885), .B(n_26535), .Z(n_180560886));
	notech_and4 i_20563567(.A(n_341962313), .B(n_179660877), .C(all_cnt[2]),
		 .D(n_27556), .Z(n_180460885));
	notech_nand2 i_1863529(.A(instrc[102]), .B(n_29025), .Z(n_180160882));
	notech_or2 i_12963422(.A(instrc[125]), .B(n_29028), .Z(n_179960880));
	notech_and4 i_20163571(.A(n_56583), .B(n_179660877), .C(n_27557), .D(n_27556
		), .Z(n_179860879));
	notech_and2 i_10863440(.A(n_27558), .B(n_27555), .Z(n_179660877));
	notech_or2 i_2863519(.A(instrc[125]), .B(instrc[127]), .Z(n_179460876)
		);
	notech_and2 i_100863550(.A(n_55325), .B(n_149060572), .Z(n_179260874));
	notech_nand2 i_13063421(.A(instrc[124]), .B(instrc[126]), .Z(n_179160873
		));
	notech_nand2 i_2163526(.A(n_178760869), .B(n_26535), .Z(n_178860870));
	notech_and4 i_20663566(.A(n_334762245), .B(n_176860850), .C(all_cnt[2]),
		 .D(n_27556), .Z(n_178760869));
	notech_nand2 i_8163466(.A(instrc[98]), .B(n_29022), .Z(n_178460866));
	notech_nand2 i_11663434(.A(instrc[104]), .B(n_29122), .Z(n_178060862));
	notech_and2 i_1963528(.A(n_177060852), .B(n_26535), .Z(n_177960861));
	notech_or4 i_76863555(.A(n_26629), .B(n_177660858), .C(n_2792), .D(n_190388902
		), .Z(n_177860860));
	notech_or2 i_3463513(.A(n_177560857), .B(n_177460856), .Z(n_177660858)
		);
	notech_nao3 i_3363514(.A(n_26625), .B(n_57444), .C(n_2594), .Z(n_177560857
		));
	notech_or4 i_1563532(.A(n_4737261), .B(n_177260854), .C(n_26496), .D(n_275888699
		), .Z(n_177460856));
	notech_nand2 i_1063537(.A(n_57441), .B(n_2824), .Z(n_177260854));
	notech_and4 i_20463568(.A(n_334862246), .B(n_176860850), .C(all_cnt[1]),
		 .D(n_27557), .Z(n_177060852));
	notech_and2 i_10963439(.A(all_cnt[0]), .B(n_27558), .Z(n_176860850));
	notech_and2 i_8063467(.A(n_29120), .B(n_29122), .Z(n_176660848));
	notech_ao4 i_75463557(.A(n_26530), .B(n_177860860), .C(n_994), .D(n_171460796
		), .Z(n_176360845));
	notech_nand3 i_12063431(.A(instrc[102]), .B(n_29025), .C(instrc[103]), .Z
		(n_176260844));
	notech_and4 i_100762575(.A(n_26531), .B(instrc[96]), .C(n_26533), .D(instrc
		[99]), .Z(n_175760839));
	notech_and4 i_100662576(.A(n_57162), .B(instrc[107]), .C(n_177960861), .D
		(n_26534), .Z(n_175660838));
	notech_ao3 i_101062573(.A(instrc[100]), .B(n_26528), .C(n_176260844), .Z
		(n_175560837));
	notech_or4 i_100962574(.A(n_176360845), .B(n_179960880), .C(n_29032), .D
		(n_28970), .Z(n_175460836));
	notech_or4 i_101262571(.A(n_183360907), .B(n_323888452), .C(n_59235), .D
		(n_28566), .Z(n_175360835));
	notech_or4 i_101162572(.A(n_183160905), .B(n_28972), .C(instrc[93]), .D(n_29034
		), .Z(n_175260834));
	notech_or2 i_101662567(.A(n_55965), .B(n_148160563), .Z(n_175160833));
	notech_or4 i_101962564(.A(n_56449), .B(n_56431), .C(n_184760921), .D(n_60512
		), .Z(n_174860830));
	notech_and4 i_99062592(.A(n_57162), .B(instrc[107]), .C(n_177960861), .D
		(n_176660848), .Z(n_174360825));
	notech_or4 i_98962593(.A(instrc[96]), .B(n_29016), .C(n_178460866), .D(n_178860870
		), .Z(n_174260824));
	notech_nao3 i_99262590(.A(n_29033), .B(n_26528), .C(n_176260844), .Z(n_174160823
		));
	notech_or4 i_99162591(.A(n_176360845), .B(n_179960880), .C(n_28970), .D(instrc
		[124]), .Z(n_174060822));
	notech_ao4 i_99562587(.A(n_56177), .B(n_56158), .C(n_147660558), .D(n_26521
		), .Z(n_173960821));
	notech_or4 i_99462588(.A(n_183360907), .B(n_323888452), .C(n_59235), .D(instrc
		[120]), .Z(n_173860820));
	notech_or4 i_99362589(.A(n_183160905), .B(n_28972), .C(instrc[93]), .D(instrc
		[92]), .Z(n_173760819));
	notech_or2 i_99862584(.A(n_56139), .B(n_148160563), .Z(n_173660818));
	notech_or4 i_100162581(.A(n_2349), .B(n_56431), .C(n_184760921), .D(n_60512
		), .Z(n_173360815));
	notech_or4 i_97362609(.A(n_183160905), .B(n_29034), .C(instrc[94]), .D(n_29026
		), .Z(n_172860810));
	notech_or4 i_97262610(.A(n_188460958), .B(n_29025), .C(n_29029), .D(n_180560886
		), .Z(n_172760809));
	notech_ao4 i_97562607(.A(n_56196), .B(n_56074), .C(n_147260554), .D(n_26518
		), .Z(n_172660808));
	notech_or4 i_97462608(.A(n_176360845), .B(n_29032), .C(instrc[126]), .D(n_221961291
		), .Z(n_172560807));
	notech_nao3 i_97862604(.A(n_177960861), .B(n_189760971), .C(n_189660970)
		, .Z(n_172460806));
	notech_or2 i_98162601(.A(n_56182), .B(n_185560929), .Z(n_172160803));
	notech_or4 i_98462598(.A(n_56449), .B(n_355988238), .C(n_184760921), .D(n_60512
		), .Z(n_171860800));
	notech_or4 i_14263409(.A(n_2603), .B(n_26615), .C(n_26377), .D(n_26536),
		 .Z(n_171560797));
	notech_and2 i_5563492(.A(n_54761), .B(n_179260874), .Z(n_171460796));
	notech_or4 i_15863393(.A(n_29022), .B(instrc[96]), .C(n_29016), .D(instrc
		[98]), .Z(n_171160793));
	notech_or4 i_15663395(.A(n_29025), .B(n_29029), .C(instrc[100]), .D(instrc
		[102]), .Z(n_171060792));
	notech_or4 i_15063401(.A(n_29023), .B(instrc[88]), .C(n_29017), .D(instrc
		[90]), .Z(n_170960791));
	notech_or4 i_14763404(.A(n_29122), .B(instrc[104]), .C(n_29040), .D(n_57162
		), .Z(n_170860790));
	notech_or4 i_95362628(.A(n_221961291), .B(n_191760991), .C(n_994), .D(n_171460796
		), .Z(n_169960781));
	notech_or4 i_95262629(.A(n_26496), .B(n_171560797), .C(n_4737261), .D(n_191560989
		), .Z(n_169860780));
	notech_or4 i_95762624(.A(n_170914103), .B(n_2793), .C(n_177460856), .D(n_146760549
		), .Z(n_169560777));
	notech_ao4 i_95662625(.A(n_56172), .B(n_56074), .C(n_146860550), .D(n_26515
		), .Z(n_169460776));
	notech_nao3 i_93662645(.A(instrc[96]), .B(n_29022), .C(n_190460978), .Z(n_169060772
		));
	notech_or4 i_93562646(.A(n_188460958), .B(n_29029), .C(instrc[101]), .D(n_180560886
		), .Z(n_168960771));
	notech_or4 i_93862643(.A(n_183160905), .B(n_29034), .C(instrc[94]), .D(instrc
		[93]), .Z(n_168860770));
	notech_or4 i_93762644(.A(n_176360845), .B(n_179960880), .C(instrc[126]),
		 .D(n_29032), .Z(n_168760769));
	notech_nand3 i_94162640(.A(n_177960861), .B(n_189760971), .C(n_26534), .Z
		(n_168660768));
	notech_nao3 i_94062641(.A(instrc[91]), .B(n_29014), .C(n_184660920), .Z(n_168560767
		));
	notech_nand3 i_92462657(.A(n_177960861), .B(n_189760971), .C(n_176660848
		), .Z(n_167260754));
	notech_ao4 i_92362658(.A(n_56172), .B(n_58656), .C(n_145960541), .D(n_26495
		), .Z(n_167160753));
	notech_or4 i_92262659(.A(n_1909), .B(n_60532), .C(n_183360907), .D(instrc
		[121]), .Z(n_167060752));
	notech_or4 i_92762654(.A(n_59259), .B(n_59268), .C(n_56172), .D(n_148160563
		), .Z(n_166960751));
	notech_or4 i_93062651(.A(n_263436789), .B(tcmp), .C(n_54865), .D(n_60512
		), .Z(n_166660748));
	notech_and4 i_7663471(.A(n_260261630), .B(n_259861626), .C(n_54893), .D(n_322762231
		), .Z(n_166360745));
	notech_or4 i_91762664(.A(n_166360745), .B(n_179160873), .C(n_60563), .D(n_198661060
		), .Z(n_166260744));
	notech_or2 i_15563396(.A(tcmp), .B(n_60512), .Z(n_166160743));
	notech_and4 i_90662675(.A(instrc[102]), .B(instrc[101]), .C(instrc[100])
		, .D(n_198161055), .Z(n_166060742));
	notech_ao3 i_90562676(.A(instrc[92]), .B(instrc[94]), .C(n_197861052), .Z
		(n_165960741));
	notech_nor2 i_90862673(.A(tcmp), .B(n_145660538), .Z(n_165860740));
	notech_and4 i_90762674(.A(n_26531), .B(n_29016), .C(instrc[98]), .D(n_26460
		), .Z(n_165760739));
	notech_nor2 i_91162670(.A(n_323062234), .B(n_185960933), .Z(n_165660738)
		);
	notech_or4 i_89262689(.A(n_221961291), .B(n_26530), .C(n_29032), .D(n_28970
		), .Z(n_164860730));
	notech_and4 i_89162690(.A(n_177060852), .B(n_57162), .C(instrc[107]), .D
		(n_26461), .Z(n_164760729));
	notech_and4 i_88862693(.A(n_198061054), .B(instrc[100]), .C(instrc[103])
		, .D(n_180460885), .Z(n_164460726));
	notech_and4 i_88762694(.A(n_182960903), .B(instrc[93]), .C(instrc[94]), 
		.D(n_202261096), .Z(n_164360725));
	notech_and4 i_89062691(.A(instrc[88]), .B(instrc[89]), .C(n_184360917), 
		.D(n_26526), .Z(n_164260724));
	notech_and4 i_88962692(.A(n_178760869), .B(n_26460), .C(instrc[98]), .D(instrc
		[99]), .Z(n_164160723));
	notech_nao3 i_89962682(.A(n_59141), .B(n_26242), .C(n_28975), .Z(n_163860720
		));
	notech_ao4 i_89862683(.A(n_200761081), .B(n_201361087), .C(n_59141), .D(n_145260534
		), .Z(n_163760719));
	notech_and2 i_89562686(.A(n_55006), .B(n_200861082), .Z(n_163560717));
	notech_ao4 i_30023(.A(n_201661090), .B(n_59944), .C(n_2191), .D(n_26887)
		, .Z(n_163460716));
	notech_ao3 i_88562695(.A(n_135460436), .B(n_26606), .C(n_494), .Z(n_163360715
		));
	notech_nand3 i_15263399(.A(instrc[126]), .B(n_29032), .C(\opcode[0] ), .Z
		(n_163260714));
	notech_and4 i_7863469(.A(n_317388516), .B(n_317288517), .C(n_55222), .D(n_319188498
		), .Z(n_163160713));
	notech_or4 i_88462696(.A(n_60563), .B(n_135060432), .C(n_163160713), .D(n_198661060
		), .Z(n_163060712));
	notech_nand2 i_27018(.A(instrc[94]), .B(n_29034), .Z(n_162960711));
	notech_ao3 i_87462706(.A(instrc[90]), .B(n_29017), .C(n_203561109), .Z(n_162860710
		));
	notech_and4 i_87362707(.A(n_198161055), .B(instrc[102]), .C(n_29033), .D
		(instrc[101]), .Z(n_162760709));
	notech_nor2 i_87662704(.A(n_59141), .B(n_144860530), .Z(n_162660708));
	notech_ao3 i_87562705(.A(n_198461058), .B(instrc[98]), .C(n_137360455), 
		.Z(n_162560707));
	notech_nor2 i_87962701(.A(n_137960461), .B(n_199861072), .Z(n_162460706)
		);
	notech_or4 i_88262698(.A(instrc[123]), .B(n_183460908), .C(n_28567), .D(instrc
		[120]), .Z(n_162160703));
	notech_ao3 i_85762723(.A(n_28567), .B(n_26558), .C(n_183460908), .Z(n_161560697
		));
	notech_or4 i_85662724(.A(instrc[127]), .B(instrc[125]), .C(n_176360845),
		 .D(n_179160873), .Z(n_161460696));
	notech_and4 i_85962721(.A(n_183060904), .B(n_29030), .C(instrc[92]), .D(n_182660900
		), .Z(n_161360695));
	notech_and4 i_85862722(.A(instrc[96]), .B(instrc[98]), .C(n_29022), .D(n_198461058
		), .Z(n_161260694));
	notech_ao3 i_86262718(.A(instrc[90]), .B(n_29017), .C(n_184660920), .Z(n_161160693
		));
	notech_and4 i_86062720(.A(instrc[102]), .B(n_198161055), .C(n_29025), .D
		(instrc[100]), .Z(n_161060692));
	notech_or2 i_86562715(.A(n_55906), .B(n_148160563), .Z(n_160960691));
	notech_or4 i_86862712(.A(n_56431), .B(n_231461383), .C(n_184760921), .D(n_60511
		), .Z(n_160660688));
	notech_nand2 i_82362756(.A(n_55992), .B(n_26542), .Z(n_160160683));
	notech_ao4 i_82262757(.A(n_141960501), .B(n_26476), .C(n_26427), .D(n_207661150
		), .Z(n_160060682));
	notech_nand3 i_82162758(.A(n_26772), .B(n_60532), .C(n_141360495), .Z(n_159960681
		));
	notech_and4 i_81762762(.A(n_26377), .B(n_57458), .C(n_26478), .D(n_141160493
		), .Z(n_158660668));
	notech_nao3 i_80162776(.A(instrc[124]), .B(n_28970), .C(n_199961073), .Z
		(n_157660658));
	notech_or4 i_78662789(.A(n_2689), .B(n_59141), .C(n_60512), .D(n_54865),
		 .Z(n_155360635));
	notech_ao4 i_75662817(.A(n_139260474), .B(n_26476), .C(n_26549), .D(n_219361266
		), .Z(n_155260634));
	notech_ao3 i_75562818(.A(n_141360495), .B(n_59235), .C(n_273888717), .Z(n_155160633
		));
	notech_and4 i_76462809(.A(n_184360917), .B(instrc[88]), .C(n_29023), .D(n_26469
		), .Z(n_154860630));
	notech_and4 i_76362810(.A(instrc[96]), .B(n_29022), .C(n_178760869), .D(n_217461247
		), .Z(n_154760629));
	notech_or4 i_76662807(.A(n_188460958), .B(n_26529), .C(instrc[101]), .D(instrc
		[103]), .Z(n_154660628));
	notech_and4 i_76562808(.A(n_177060852), .B(n_26534), .C(n_29040), .D(n_29008
		), .Z(n_154560627));
	notech_nor2 i_77162804(.A(n_57373), .B(n_26524), .Z(n_154460626));
	notech_ao3 i_77062805(.A(n_56458), .B(n_195658242), .C(n_26523), .Z(n_154360625
		));
	notech_and4 i_76962806(.A(n_182960903), .B(n_29026), .C(n_29030), .D(n_26459
		), .Z(n_154260624));
	notech_or4 i_75262820(.A(n_177560857), .B(n_177460856), .C(n_2205), .D(n_26544
		), .Z(n_154160623));
	notech_or4 i_9307(.A(n_214461218), .B(n_215061224), .C(opa[6]), .D(n_1845
		), .Z(n_153760619));
	notech_nao3 i_73362839(.A(n_183060904), .B(n_29030), .C(n_196361037), .Z
		(n_153460616));
	notech_or2 i_73262840(.A(n_213261206), .B(n_196061034), .Z(n_153360615)
		);
	notech_or4 i_73562837(.A(instrc[127]), .B(instrc[125]), .C(n_176360845),
		 .D(n_191760991), .Z(n_153260614));
	notech_or4 i_73462838(.A(n_193161005), .B(instrc[103]), .C(n_180560886),
		 .D(instrc[101]), .Z(n_153160613));
	notech_or4 i_73762835(.A(instrc[104]), .B(instrc[105]), .C(n_57162), .D(n_199761071
		), .Z(n_153060612));
	notech_ao4 i_73662836(.A(n_58656), .B(n_56108), .C(n_138460466), .D(n_26464
		), .Z(n_152960611));
	notech_or4 i_74462828(.A(n_114626850), .B(n_229364616), .C(n_184760921),
		 .D(n_60512), .Z(n_152260604));
	notech_nand3 i_36179(.A(n_56583), .B(n_135360435), .C(n_221861290), .Z(n_152160603
		));
	notech_nand3 i_36324(.A(n_56100), .B(n_56425), .C(n_135260434), .Z(n_152060602
		));
	notech_or4 i_36322(.A(n_56458), .B(n_355988238), .C(n_56440), .D(n_26382
		), .Z(n_151960601));
	notech_nao3 i_22563563(.A(n_56469), .B(n_56458), .C(n_56431), .Z(n_151860600
		));
	notech_or4 i_36320(.A(n_26251), .B(n_26382), .C(n_26384), .D(n_26550), .Z
		(n_151760599));
	notech_or4 i_36389(.A(n_29008), .B(n_26385), .C(n_29040), .D(instrc[105]
		), .Z(n_151260594));
	notech_nand2 i_71862854(.A(n_137960461), .B(n_29008), .Z(n_151160593));
	notech_nand2 i_36461(.A(n_341962313), .B(n_135560437), .Z(n_151060592)
		);
	notech_or4 i_36531(.A(n_29013), .B(n_26386), .C(n_29016), .D(instrc[97])
		, .Z(n_150960591));
	notech_nand2 i_70462867(.A(n_137360455), .B(n_29013), .Z(n_150860590));
	notech_nand3 i_36605(.A(instrc[94]), .B(n_29026), .C(instrc[95]), .Z(n_150760589
		));
	notech_or4 i_36602(.A(instrc[92]), .B(instrc[94]), .C(n_29026), .D(n_29030
		), .Z(n_150660588));
	notech_nand2 i_69762874(.A(n_29026), .B(n_28972), .Z(n_150560587));
	notech_or4 i_36669(.A(n_29014), .B(n_26388), .C(n_29017), .D(instrc[89])
		, .Z(n_150460586));
	notech_or4 i_38163184(.A(n_56369), .B(n_58483), .C(n_60595), .D(n_27583)
		, .Z(n_150160583));
	notech_or2 i_38463181(.A(n_353988269), .B(n_56784), .Z(n_149860580));
	notech_or2 i_38763178(.A(n_354488264), .B(\nbus_11276[17] ), .Z(n_149560577
		));
	notech_or4 i_103062553(.A(n_58945), .B(n_273288723), .C(n_2260), .D(n_54520
		), .Z(n_149060572));
	notech_ao4 i_180663546(.A(n_59380), .B(n_62431), .C(n_2264), .D(n_26384)
		, .Z(n_148560567));
	notech_or4 i_102362560(.A(n_54523), .B(n_182060895), .C(n_29032), .D(n_29028
		), .Z(n_148460566));
	notech_or4 i_102262561(.A(n_59141), .B(n_2250), .C(n_151860600), .D(n_60512
		), .Z(n_148360565));
	notech_and2 i_2663521(.A(n_148460566), .B(n_135160433), .Z(n_148260564)
		);
	notech_and2 i_363544(.A(n_134960431), .B(n_181560891), .Z(n_148160563)
		);
	notech_ao4 i_96963551(.A(n_177860860), .B(n_26523), .C(n_184960923), .D(n_60512
		), .Z(n_148060562));
	notech_and2 i_463543(.A(n_184960923), .B(n_184760921), .Z(n_147960561)
		);
	notech_or4 i_100562577(.A(n_182060895), .B(n_2650), .C(instrc[124]), .D(n_29028
		), .Z(n_147760559));
	notech_ao3 i_100462578(.A(n_62409), .B(n_26550), .C(n_134960431), .Z(n_147660558
		));
	notech_and2 i_3563512(.A(n_147760559), .B(n_54508), .Z(n_147560557));
	notech_or4 i_98862594(.A(n_54525), .B(n_221961291), .C(n_60563), .D(n_188960963
		), .Z(n_147360555));
	notech_ao3 i_98762595(.A(n_62409), .B(n_26241), .C(n_134960431), .Z(n_147260554
		));
	notech_and2 i_4363504(.A(n_147360555), .B(n_54494), .Z(n_147160553));
	notech_or4 i_96262619(.A(n_191760991), .B(n_221961291), .C(n_60563), .D(n_26410
		), .Z(n_146960551));
	notech_ao3 i_96162620(.A(n_62433), .B(n_26251), .C(n_134960431), .Z(n_146860550
		));
	notech_and4 i_16663385(.A(n_193561009), .B(n_193461008), .C(n_193261006)
		, .D(n_193061004), .Z(n_146760549));
	notech_and2 i_16463387(.A(n_192260996), .B(n_323288458), .Z(n_146560547)
		);
	notech_or4 i_95062631(.A(n_1025), .B(n_59141), .C(n_2250), .D(n_60507), 
		.Z(n_146360545));
	notech_ao4 i_4563502(.A(n_56183), .B(n_1023), .C(n_179960880), .D(n_194861022
		), .Z(n_146260544));
	notech_ao3 i_93362648(.A(n_62427), .B(n_26304), .C(n_134960431), .Z(n_145960541
		));
	notech_ao4 i_4663501(.A(n_997), .B(n_56290), .C(n_196761041), .D(n_179960880
		), .Z(n_145860540));
	notech_and4 i_16963382(.A(n_166260744), .B(n_323762241), .C(n_353488274)
		, .D(n_199161065), .Z(n_145660538));
	notech_or2 i_90262679(.A(n_2261), .B(n_59141), .Z(n_145360535));
	notech_and3 i_90162680(.A(n_54505), .B(n_56223), .C(n_200961083), .Z(n_145260534
		));
	notech_and2 i_89762684(.A(n_200761081), .B(n_26887), .Z(n_144960531));
	notech_and4 i_17063381(.A(n_55133), .B(n_204061114), .C(n_323731624), .D
		(n_320388486), .Z(n_144860530));
	notech_or4 i_87262708(.A(n_182060895), .B(n_293061934), .C(n_29032), .D(instrc
		[127]), .Z(n_144760529));
	notech_or4 i_87162709(.A(n_56431), .B(n_231461383), .C(n_134960431), .D(n_60504
		), .Z(n_144660528));
	notech_and2 i_3663511(.A(n_144760529), .B(n_312462128), .Z(n_144560527)
		);
	notech_mux2 i_9563452(.S(all_cnt[2]), .A(n_56415), .B(n_334762245), .Z(n_143160513
		));
	notech_nao3 i_84562735(.A(all_cnt[0]), .B(n_27556), .C(n_143160513), .Z(n_143060512
		));
	notech_or2 i_84462736(.A(n_2822), .B(n_29130), .Z(n_142960511));
	notech_mux4 i_13963412(.S0(all_cnt[1]), .S1(all_cnt[2]), .A(n_56583), .B
		(n_56425), .C(n_341962313), .D(n_334662244), .Z(n_142860510));
	notech_and2 i_14163410(.A(n_207161145), .B(n_143060512), .Z(n_142760509)
		);
	notech_nand2 i_17263379(.A(n_142960511), .B(n_207261146), .Z(n_142660508
		));
	notech_ao3 i_84162739(.A(n_61175), .B(n_142660508), .C(n_494), .Z(n_142560507
		));
	notech_or4 i_83262748(.A(n_135060432), .B(n_54935), .C(n_179460876), .D(n_60563
		), .Z(n_142460506));
	notech_or4 i_83062749(.A(n_60752), .B(n_60739), .C(n_60779), .D(n_179260874
		), .Z(n_142360505));
	notech_or4 i_82962750(.A(n_60779), .B(n_60729), .C(n_1900), .D(n_54520),
		 .Z(n_142260504));
	notech_nor2 i_82662753(.A(n_56363), .B(n_26583), .Z(n_141960501));
	notech_and2 i_2463523(.A(n_101413408), .B(n_142360505), .Z(n_141860500)
		);
	notech_and3 i_5763490(.A(n_55820), .B(n_55580), .C(n_56363), .Z(n_141760499
		));
	notech_ao4 i_13163420(.A(n_55523), .B(n_306062064), .C(n_55794), .D(n_26477
		), .Z(n_141660498));
	notech_nand2 i_2763520(.A(n_101213406), .B(n_142260504), .Z(n_141360495)
		);
	notech_or4 i_17663375(.A(n_212061194), .B(n_211761191), .C(n_210761181),
		 .D(n_211461188), .Z(n_141160493));
	notech_and4 i_17463377(.A(n_208361157), .B(n_159960681), .C(n_160160683)
		, .D(n_26475), .Z(n_140960491));
	notech_ao4 i_17363378(.A(n_57458), .B(n_57441), .C(n_171560797), .D(n_142960511
		), .Z(n_140860490));
	notech_or4 i_81062767(.A(n_243964756), .B(n_59141), .C(n_2250), .D(n_60504
		), .Z(n_140660488));
	notech_ao4 i_4763500(.A(n_57343), .B(n_243664753), .C(n_198661060), .D(n_212961203
		), .Z(n_140560487));
	notech_and2 i_17763374(.A(n_140660488), .B(n_213061204), .Z(n_140460486)
		);
	notech_or4 i_78962786(.A(n_56458), .B(n_1189), .C(n_134960431), .D(n_60504
		), .Z(n_140060482));
	notech_ao4 i_4863499(.A(n_1076), .B(n_197114365), .C(n_215661230), .D(n_198661060
		), .Z(n_139960481));
	notech_and2 i_17863373(.A(n_140060482), .B(n_215761231), .Z(n_139860480)
		);
	notech_or4 i_76262811(.A(n_188960963), .B(n_54938), .C(n_179460876), .D(n_60563
		), .Z(n_139560477));
	notech_nor2 i_75962814(.A(n_56363), .B(n_26500), .Z(n_139260474));
	notech_ao4 i_13263419(.A(n_55523), .B(n_323788453), .C(n_55794), .D(n_26466
		), .Z(n_139160473));
	notech_or4 i_19263359(.A(n_154360625), .B(n_154260624), .C(n_218561258),
		 .D(n_154460626), .Z(n_138860470));
	notech_ao3 i_19163360(.A(n_219561268), .B(n_26465), .C(n_155160633), .Z(n_138760469
		));
	notech_ao4 i_13363418(.A(n_207461148), .B(n_141860500), .C(n_217361246),
		 .D(n_26530), .Z(n_138660468));
	notech_ao3 i_74762825(.A(n_62423), .B(n_26237), .C(n_134960431), .Z(n_138460466
		));
	notech_ao4 i_4963498(.A(n_212964463), .B(n_60484), .C(n_220561278), .D(n_179460876
		), .Z(n_138360465));
	notech_nand2 i_3163516(.A(instrc[105]), .B(n_29120), .Z(n_137960461));
	notech_and3 i_18463367(.A(n_189660970), .B(n_151160593), .C(instrc[107])
		, .Z(n_137760459));
	notech_and2 i_71062861(.A(n_29025), .B(n_28971), .Z(n_137560457));
	notech_and2 i_70962862(.A(instrc[100]), .B(n_180160882), .Z(n_137460456)
		);
	notech_nand2 i_3063517(.A(instrc[97]), .B(n_29019), .Z(n_137360455));
	notech_and3 i_18363368(.A(n_190260976), .B(n_150860590), .C(instrc[99]),
		 .Z(n_137160453));
	notech_and3 i_18263369(.A(n_188660960), .B(n_150560587), .C(instrc[95]),
		 .Z(n_136860450));
	notech_nand2 i_2963518(.A(instrc[89]), .B(n_29020), .Z(n_136660448));
	notech_and2 i_18163370(.A(n_223361304), .B(instrc[91]), .Z(n_136460446)
		);
	notech_or2 i_68062890(.A(n_55852), .B(n_26312), .Z(n_136060442));
	notech_or2 i_67862892(.A(n_56063), .B(n_26312), .Z(n_135960441));
	notech_and3 i_19463357(.A(n_55845), .B(n_55846), .C(n_55847), .Z(n_135860440
		));
	notech_and3 i_19363358(.A(n_56345), .B(n_2239), .C(n_2241), .Z(n_135760439
		));
	notech_or4 i_8663461(.A(n_198061054), .B(n_29029), .C(n_137460456), .D(n_137560457
		), .Z(n_135560437));
	notech_or4 i_7763470(.A(n_164760729), .B(n_203261106), .C(n_26486), .D(n_26485
		), .Z(n_135460436));
	notech_nao3 i_5463493(.A(instrc[125]), .B(instrc[127]), .C(n_191760991),
		 .Z(n_135360435));
	notech_nand2 i_5063497(.A(n_151860600), .B(n_56101), .Z(n_135260434));
	notech_or2 i_3863509(.A(n_148560567), .B(n_56178), .Z(n_135160433));
	notech_nand2 i_3763510(.A(instrc[126]), .B(n_29032), .Z(n_135060432));
	notech_or2 i_58163561(.A(n_59141), .B(n_2250), .Z(n_134960431));
	notech_nand2 i_54539(.A(n_46243), .B(n_201561089), .Z(n_134860430));
	notech_nao3 i_149864221(.A(n_26712), .B(n_26629), .C(n_275088707), .Z(n_134560427
		));
	notech_or4 i_149964220(.A(n_275888699), .B(n_275388704), .C(n_26540), .D
		(n_26629), .Z(n_134460426));
	notech_or4 i_90464796(.A(n_275288705), .B(n_2550), .C(n_106813462), .D(n_60474
		), .Z(n_134360425));
	notech_ao4 i_90964791(.A(n_26887), .B(n_134560427), .C(n_177560857), .D(n_134460426
		), .Z(n_134060422));
	notech_ao4 i_10568174(.A(n_2645), .B(n_273188724), .C(n_2647), .D(n_2830
		), .Z(n_133860420));
	notech_ao4 i_5868216(.A(n_54880), .B(n_133660418), .C(n_132960411), .D(n_54968
		), .Z(n_133760419));
	notech_or4 i_5768217(.A(n_60780), .B(n_60729), .C(n_60595), .D(n_56104),
		 .Z(n_133660418));
	notech_or4 i_668268(.A(n_2647), .B(tss_esp0), .C(n_58945), .D(n_272788728
		), .Z(n_133360415));
	notech_nand2 i_10268175(.A(n_133360415), .B(n_133860420), .Z(n_133260414
		));
	notech_or4 i_54737(.A(n_132760409), .B(n_132860410), .C(n_26494), .D(n_26552
		), .Z(\nbus_11353[2] ));
	notech_and3 i_368271(.A(n_56574), .B(n_56112), .C(n_57448), .Z(n_132960411
		));
	notech_and4 i_5368221(.A(n_57448), .B(n_26326), .C(n_26621), .D(n_26508)
		, .Z(n_132860410));
	notech_and3 i_5268222(.A(n_59195), .B(n_59856), .C(n_134860430), .Z(n_132760409
		));
	notech_ao4 i_107869185(.A(n_56160), .B(n_29125), .C(n_170960791), .D(n_27329
		), .Z(n_132660408));
	notech_ao4 i_107969184(.A(n_27362), .B(n_150460586), .C(n_334962247), .D
		(n_26979), .Z(n_132560407));
	notech_ao4 i_117769087(.A(n_56147), .B(n_29126), .C(n_150660588), .D(n_27310
		), .Z(n_132460406));
	notech_ao4 i_117869086(.A(n_150760589), .B(n_27342), .C(n_334662244), .D
		(n_26941), .Z(n_132360405));
	notech_ao4 i_122669039(.A(n_56150), .B(n_29127), .C(n_171160793), .D(n_27317
		), .Z(n_132260404));
	notech_ao4 i_122769038(.A(n_27350), .B(n_150960591), .C(n_334762245), .D
		(n_26955), .Z(n_132160403));
	notech_ao4 i_129068975(.A(n_151060592), .B(n_29128), .C(n_171060792), .D
		(n_27316), .Z(n_132060402));
	notech_ao4 i_129168974(.A(n_176260844), .B(n_27349), .C(n_341962313), .D
		(n_26953), .Z(n_131960401));
	notech_ao4 i_138368883(.A(n_56153), .B(n_29129), .C(n_27297), .D(n_170860790
		), .Z(n_131860400));
	notech_ao4 i_138468882(.A(n_27333), .B(n_151260594), .C(n_334862246), .D
		(n_26923), .Z(n_131760399));
	notech_ao4 i_150768759(.A(n_152160603), .B(n_29049), .C(n_135360435), .D
		(n_27298), .Z(n_131660398));
	notech_ao4 i_150868758(.A(n_21051), .B(n_27334), .C(n_56583), .D(n_26925
		), .Z(n_131560397));
	notech_or4 i_55632973(.A(n_60780), .B(n_60731), .C(n_275288705), .D(n_205588858
		), .Z(n_55793));
	notech_and2 i_71032978(.A(n_54813), .B(n_313088558), .Z(n_55640));
	notech_and4 i_163332979(.A(n_314688543), .B(n_314488544), .C(n_332088392
		), .D(n_57382), .Z(n_54813));
	notech_ao4 i_123032853(.A(n_48510), .B(n_316088529), .C(n_315988530), .D
		(n_310588583), .Z(n_2186));
	notech_nand2 i_99932875(.A(n_26712), .B(n_57445), .Z(n_2208));
	notech_or4 i_155232997(.A(n_275288705), .B(n_2550), .C(n_59944), .D(n_2826
		), .Z(n_54881));
	notech_or2 i_137033005(.A(n_206688847), .B(n_55226), .Z(n_55018));
	notech_nand2 i_155733048(.A(n_26629), .B(n_59944), .Z(n_54877));
	notech_ao4 i_57833137(.A(n_321731604), .B(n_26616), .C(n_314988540), .D(n_55226
		), .Z(n_55771));
	notech_mux2 i_138033138(.S(n_57451), .A(n_29124), .B(n_2593), .Z(n_55008
		));
	notech_and2 i_71333139(.A(n_315088539), .B(n_314888541), .Z(n_55637));
	notech_or4 i_5254(.A(n_56117), .B(n_2572), .C(n_272788728), .D(n_59945),
		 .Z(n_51840));
	notech_or4 i_2145(.A(n_2260), .B(n_272988726), .C(\opcode[1] ), .D(\opcode[0] 
		), .Z(n_57382));
	notech_and3 i_139033172(.A(n_54777), .B(n_57382), .C(n_57391), .Z(n_54998
		));
	notech_ao4 i_47644(.A(n_29123), .B(n_55637), .C(n_271039498), .D(n_312788561
		), .Z(\nbus_11286[5] ));
	notech_nand3 i_216171(.A(n_309588593), .B(n_309088598), .C(n_309988589),
		 .Z(n_14098));
	notech_nand3 i_816177(.A(n_307788611), .B(n_306988618), .C(n_307388614),
		 .Z(n_14134));
	notech_xor2 i_104135764(.A(n_27518), .B(opz[0]), .Z(n_55328));
	notech_nand2 i_5739036(.A(instrc[123]), .B(n_28567), .Z(n_323888452));
	notech_nand3 i_33122(.A(n_56458), .B(n_195658242), .C(n_62431), .Z(n_323788453
		));
	notech_or4 i_28228(.A(n_2831), .B(n_62395), .C(n_62437), .D(n_106813462)
		, .Z(n_323688454));
	notech_nand2 i_209839107(.A(n_322188469), .B(n_323588455), .Z(n_54431)
		);
	notech_nand2 i_36539085(.A(n_55667), .B(n_238958635), .Z(n_323588455));
	notech_nand2 i_206939108(.A(n_323588455), .B(n_26516), .Z(n_54455));
	notech_or4 i_200439109(.A(n_1909), .B(n_216658447), .C(n_28567), .D(n_60532
		), .Z(n_54507));
	notech_nand2 i_35939110(.A(n_55658), .B(n_238758633), .Z(n_323488456));
	notech_ao4 i_34739111(.A(n_56574), .B(n_2044), .C(n_55820), .D(n_26576),
		 .Z(n_323388457));
	notech_or4 i_28209(.A(n_56458), .B(n_355988238), .C(n_56440), .D(n_60504
		), .Z(n_323288458));
	notech_or2 i_22739112(.A(n_355988238), .B(n_2349), .Z(n_56100));
	notech_or2 i_26939(.A(instrc[123]), .B(n_28566), .Z(n_323188459));
	notech_nand2 i_86039114(.A(n_322188469), .B(n_107113465), .Z(n_323088460
		));
	notech_nand2 i_86139115(.A(n_107113465), .B(n_26516), .Z(n_322988461));
	notech_and4 i_91639144(.A(n_266858912), .B(n_266758911), .C(n_266358907)
		, .D(n_266658910), .Z(n_322788463));
	notech_and4 i_91439145(.A(n_264058884), .B(n_263958883), .C(n_263558879)
		, .D(n_263858882), .Z(n_322688464));
	notech_ao3 i_91329142(.A(n_262858872), .B(n_221058483), .C(n_221158484),
		 .Z(n_322488466));
	notech_and2 i_19188(.A(opb[0]), .B(n_59856), .Z(n_322388467));
	notech_ao4 i_35339086(.A(n_2044), .B(n_54520), .C(n_56363), .D(n_26576),
		 .Z(n_322288468));
	notech_nao3 i_198139154(.A(n_56260), .B(n_216758448), .C(n_216558446), .Z
		(n_322188469));
	notech_ao4 i_137933140(.A(n_57423), .B(n_59945), .C(n_26616), .D(n_2208)
		, .Z(n_55009));
	notech_and2 i_41633129(.A(n_55292), .B(n_54735), .Z(n_55933));
	notech_nand2 i_131439155(.A(n_322188469), .B(n_26559), .Z(n_97522962));
	notech_and2 i_96045401(.A(n_54431), .B(n_323088460), .Z(n_55403));
	notech_and2 i_96145402(.A(n_54455), .B(n_322988461), .Z(n_55402));
	notech_or2 i_8639007(.A(n_55794), .B(n_56043), .Z(n_121523202));
	notech_or4 i_8039013(.A(n_355988238), .B(n_2349), .C(n_60504), .D(n_322288468
		), .Z(n_121623203));
	notech_or4 i_8339010(.A(n_56458), .B(n_355988238), .C(n_216358445), .D(n_56440
		), .Z(n_121723204));
	notech_and2 i_33538(.A(n_57312), .B(n_2186), .Z(n_2312));
	notech_or4 i_31435692(.A(n_60752), .B(n_60739), .C(n_60779), .D(n_55389)
		, .Z(n_329546800));
	notech_nand3 i_33632912(.A(n_26556), .B(n_59945), .C(n_2797), .Z(n_2248)
		);
	notech_nao3 i_33732911(.A(n_26556), .B(n_59944), .C(n_2797), .Z(n_2247)
		);
	notech_or2 i_33523(.A(n_57451), .B(n_59856), .Z(n_2313));
	notech_or4 i_33522(.A(n_60752), .B(n_60739), .C(n_60779), .D(n_54998), .Z
		(n_2314));
	notech_or4 i_33518(.A(n_275288705), .B(n_60494), .C(n_2253), .D(n_59944)
		, .Z(n_231547139));
	notech_nand2 i_33678(.A(n_55159), .B(n_59856), .Z(n_2311));
	notech_or4 i_42032910(.A(n_2582), .B(n_2599), .C(n_59856), .D(n_2792), .Z
		(n_2246));
	notech_nao3 i_4745330(.A(n_56458), .B(n_195658242), .C(n_215558439), .Z(n_302421911
		));
	notech_or4 i_4945328(.A(n_59259), .B(n_59268), .C(n_59281), .D(n_55088),
		 .Z(n_302221909));
	notech_or2 i_89545429(.A(n_215558439), .B(n_54938), .Z(n_55459));
	notech_and3 i_121332854(.A(n_54719), .B(n_313388555), .C(n_54725), .Z(n_2187
		));
	notech_ao4 i_93839106(.A(n_323688454), .B(n_59935), .C(n_322288468), .D(n_54507
		), .Z(n_322088470));
	notech_or4 i_30632913(.A(n_273488721), .B(n_59856), .C(n_2792), .D(n_26611
		), .Z(n_2249));
	notech_nand3 i_208549159(.A(rep_en2), .B(n_2770), .C(n_26596), .Z(n_321988471
		));
	notech_or2 i_48649182(.A(n_208258368), .B(n_26560), .Z(n_321888472));
	notech_or4 i_47049183(.A(rep_en2), .B(rep_en3), .C(n_213358418), .D(n_26890
		), .Z(n_21822205));
	notech_or2 i_30207(.A(n_54707), .B(\eflags[10] ), .Z(n_321788473));
	notech_or2 i_30209(.A(n_54707), .B(n_55450), .Z(n_321688474));
	notech_nao3 i_33206(.A(n_56458), .B(n_195658242), .C(n_216158443), .Z(n_321588475
		));
	notech_or2 i_33124(.A(n_316988520), .B(n_323788453), .Z(n_131123298));
	notech_or2 i_31395(.A(n_56478), .B(n_56469), .Z(n_114626850));
	notech_and3 i_56839148(.A(n_317188518), .B(n_217058450), .C(n_55690), .Z
		(n_3214));
	notech_and4 i_91739151(.A(n_317988510), .B(n_55265), .C(n_55978), .D(n_318788502
		), .Z(n_321388476));
	notech_and4 i_91939152(.A(n_318088509), .B(n_55257), .C(n_318688503), .D
		(n_55979), .Z(n_321288477));
	notech_and4 i_91529143(.A(n_265458898), .B(n_265358897), .C(n_264958893)
		, .D(n_265258896), .Z(n_321188478));
	notech_and2 i_24351993(.A(n_56458), .B(n_195658242), .Z(n_321088479));
	notech_nao3 i_24451992(.A(n_28966), .B(n_56440), .C(n_55522), .Z(n_320988480
		));
	notech_or2 i_158151968(.A(n_57373), .B(n_183258118), .Z(n_320888481));
	notech_or2 i_152451969(.A(n_182758113), .B(n_56270), .Z(n_320788482));
	notech_or4 i_120451972(.A(n_56458), .B(n_56469), .C(n_55522), .D(n_187758163
		), .Z(n_320688483));
	notech_ao4 i_52651987(.A(n_56112), .B(n_204988864), .C(n_2239), .D(n_26500
		), .Z(n_320588484));
	notech_and2 i_30485(.A(n_317588514), .B(n_317488515), .Z(n_320388486));
	notech_or4 i_30479(.A(n_56458), .B(n_55522), .C(n_317788512), .D(n_56469
		), .Z(n_320188488));
	notech_or4 i_124252069(.A(instrc[115]), .B(instrc[112]), .C(n_2250), .D(n_59250
		), .Z(n_320088489));
	notech_and2 i_30395(.A(n_320088489), .B(n_319488495), .Z(n_319988490));
	notech_or2 i_115052011(.A(n_317888511), .B(n_317788512), .Z(n_55222));
	notech_or4 i_113452012(.A(n_2740), .B(n_182758113), .C(n_317788512), .D(n_59235
		), .Z(n_55238));
	notech_nand2 i_27030(.A(n_28966), .B(n_56440), .Z(n_319888491));
	notech_mux2 i_711664(.S(n_60138), .A(n_562), .B(add_len_pc32[6]), .Z(n_319788492
		));
	notech_mux2 i_511662(.S(n_60138), .A(n_560), .B(add_len_pc32[4]), .Z(n_319688493
		));
	notech_and4 i_142752032(.A(n_196958255), .B(n_196858254), .C(n_196458250
		), .D(n_196758253), .Z(n_319588494));
	notech_or4 i_10728(.A(instrc[115]), .B(instrc[112]), .C(n_2239), .D(n_59250
		), .Z(n_319488495));
	notech_ao4 i_52151988(.A(n_204988864), .B(n_56112), .C(n_2239), .D(n_26581
		), .Z(n_319388496));
	notech_and2 i_57552043(.A(n_317088519), .B(n_319988490), .Z(n_319288497)
		);
	notech_or2 i_10725(.A(n_319388496), .B(n_317888511), .Z(n_319188498));
	notech_and3 i_85152044(.A(n_317388516), .B(n_317288517), .C(n_319188498)
		, .Z(n_319088499));
	notech_or4 i_10723(.A(n_2740), .B(n_182758113), .C(n_319388496), .D(n_59235
		), .Z(n_318988500));
	notech_and3 i_85252045(.A(n_317588514), .B(n_317488515), .C(n_318988500)
		, .Z(n_318888501));
	notech_or2 i_7534(.A(n_320588484), .B(n_54938), .Z(n_318788502));
	notech_or2 i_7532(.A(n_320588484), .B(n_320888481), .Z(n_318688503));
	notech_or4 i_33314(.A(n_60595), .B(n_59856), .C(n_273688719), .D(n_28140
		), .Z(n_318588504));
	notech_or4 i_33340(.A(n_60596), .B(n_59845), .C(n_273688719), .D(n_60138
		), .Z(n_318488505));
	notech_or2 i_174852081(.A(n_316988520), .B(n_54938), .Z(n_318388506));
	notech_or2 i_171452080(.A(n_316988520), .B(n_320888481), .Z(n_318288507)
		);
	notech_or2 i_154052063(.A(n_55825), .B(n_320888481), .Z(n_318088509));
	notech_or2 i_153252064(.A(n_55825), .B(n_54938), .Z(n_317988510));
	notech_and3 i_149152065(.A(n_56260), .B(n_182858114), .C(n_182658112), .Z
		(n_317888511));
	notech_or4 i_126352067(.A(n_59259), .B(n_59268), .C(n_59277), .D(n_2250)
		, .Z(n_131423301));
	notech_ao4 i_51952070(.A(n_56574), .B(n_204988864), .C(n_2241), .D(n_26581
		), .Z(n_317788512));
	notech_ao4 i_52252071(.A(n_56574), .B(n_204988864), .C(n_2241), .D(n_26500
		), .Z(n_317688513));
	notech_or4 i_140352082(.A(n_2740), .B(n_182758113), .C(n_55829), .D(n_59235
		), .Z(n_317588514));
	notech_or4 i_170452083(.A(n_2740), .B(n_182758113), .C(n_316888521), .D(n_59235
		), .Z(n_317488515));
	notech_ao4 i_52052013(.A(n_204988864), .B(n_56104), .C(n_56345), .D(n_26581
		), .Z(n_55829));
	notech_or2 i_141052084(.A(n_317888511), .B(n_55829), .Z(n_317388516));
	notech_or2 i_168452085(.A(n_317888511), .B(n_316888521), .Z(n_317288517)
		);
	notech_or4 i_66252086(.A(instrc[115]), .B(instrc[112]), .C(n_2241), .D(n_59250
		), .Z(n_55688));
	notech_or4 i_65452088(.A(n_59259), .B(n_59268), .C(n_59277), .D(n_56345)
		, .Z(n_317188518));
	notech_or4 i_65952090(.A(instrc[115]), .B(n_59290), .C(n_56345), .D(n_59250
		), .Z(n_317088519));
	notech_ao4 i_38352091(.A(n_56059), .B(n_60596), .C(n_2250), .D(n_26500),
		 .Z(n_316988520));
	notech_ao4 i_38152092(.A(n_60596), .B(n_56059), .C(n_26581), .D(n_2250),
		 .Z(n_316888521));
	notech_and4 i_1116660(.A(n_181758104), .B(n_181658103), .C(n_181558102),
		 .D(n_182158107), .Z(n_11752));
	notech_nand2 i_1216661(.A(n_180858095), .B(n_180358090), .Z(n_11758));
	notech_nand2 i_1316662(.A(n_179758085), .B(n_179258080), .Z(n_11764));
	notech_nand2 i_1416663(.A(n_178658074), .B(n_178158069), .Z(n_11770));
	notech_nand2 i_1616665(.A(n_177558063), .B(n_177058058), .Z(n_11782));
	notech_nand2 i_920628(.A(n_176358051), .B(n_175858046), .Z(n_20159));
	notech_nand2 i_1120630(.A(n_175358041), .B(n_174858036), .Z(n_20171));
	notech_nand2 i_1220631(.A(n_172758015), .B(n_172258010), .Z(n_20177));
	notech_nand2 i_1320632(.A(n_170157989), .B(n_169657984), .Z(n_20183));
	notech_nand2 i_1420633(.A(n_167557963), .B(n_167057958), .Z(n_20189));
	notech_and4 i_143655318(.A(n_166157949), .B(n_166057948), .C(n_165657944
		), .D(n_165957947), .Z(n_321831605));
	notech_and4 i_143555319(.A(n_168757975), .B(n_168657974), .C(n_168257970
		), .D(n_168557973), .Z(n_321931606));
	notech_and4 i_143455320(.A(n_171358001), .B(n_171258000), .C(n_170857996
		), .D(n_171157999), .Z(n_322031607));
	notech_and4 i_143355321(.A(n_173958027), .B(n_173858026), .C(n_173458022
		), .D(n_173758025), .Z(n_322131608));
	notech_mux2 i_1411671(.S(n_60138), .A(n_569), .B(add_len_pc32[13]), .Z(\add_len_pc[13] 
		));
	notech_mux2 i_1311670(.S(n_60138), .A(n_568), .B(add_len_pc32[12]), .Z(\add_len_pc[12] 
		));
	notech_mux2 i_1211669(.S(n_60138), .A(n_567), .B(add_len_pc32[11]), .Z(\add_len_pc[11] 
		));
	notech_mux2 i_1111668(.S(n_60138), .A(n_566), .B(add_len_pc32[10]), .Z(\add_len_pc[10] 
		));
	notech_mux2 i_911666(.S(n_60138), .A(n_564), .B(add_len_pc32[8]), .Z(\add_len_pc[8] 
		));
	notech_or4 i_45552016(.A(n_56574), .B(n_60596), .C(n_59935), .D(n_1900),
		 .Z(n_316788522));
	notech_nand3 i_57052015(.A(n_56056), .B(n_59195), .C(n_59845), .Z(n_316688523
		));
	notech_mux2 i_162333126(.S(n_59931), .A(n_311388575), .B(n_273688719), .Z
		(n_54822));
	notech_nand2 i_26786(.A(opc_10[6]), .B(n_62431), .Z(n_316588524));
	notech_nand2 i_26787(.A(n_62423), .B(opc[6]), .Z(n_316488525));
	notech_nand2 i_26868(.A(n_62433), .B(opc[4]), .Z(n_316388526));
	notech_nand2 i_26867(.A(opc_10[4]), .B(n_62431), .Z(n_316288527));
	notech_ao4 i_56233149(.A(n_54881), .B(n_26600), .C(n_2105), .D(n_59931),
		 .Z(n_55787));
	notech_ao3 i_56133148(.A(n_55943), .B(n_54762), .C(n_313488554), .Z(n_55788
		));
	notech_ao4 i_55733147(.A(n_57445), .B(n_59845), .C(n_315488535), .D(n_315388536
		), .Z(n_55792));
	notech_mux2 i_50133146(.S(n_59931), .A(n_57419), .B(n_315588534), .Z(n_55848
		));
	notech_mux2 i_50033145(.S(n_59935), .A(n_57420), .B(n_275788700), .Z(n_55849
		));
	notech_ao4 i_127557869(.A(n_55854), .B(n_55289), .C(n_1135), .D(n_29050)
		, .Z(n_249234118));
	notech_ao4 i_127457870(.A(n_55854), .B(n_59753), .C(n_1135), .D(n_29049)
		, .Z(n_249334119));
	notech_and2 i_116757873(.A(n_55270), .B(n_55302), .Z(n_249634122));
	notech_and2 i_116557874(.A(n_55355), .B(n_120357491), .Z(n_249734123));
	notech_and2 i_77457897(.A(n_121357501), .B(n_55841), .Z(n_252034146));
	notech_nand2 i_1717563(.A(n_141957707), .B(n_141457702), .Z(n_20939));
	notech_and4 i_216651(.A(n_140557693), .B(n_140457692), .C(n_140857696), 
		.D(n_140357691), .Z(n_11698));
	notech_and4 i_316652(.A(n_139357681), .B(n_139257680), .C(n_139657684), 
		.D(n_139157679), .Z(n_11704));
	notech_and4 i_516654(.A(n_138157669), .B(n_138057668), .C(n_125757545), 
		.D(n_138457672), .Z(n_11716));
	notech_and4 i_616655(.A(n_137057658), .B(n_136957657), .C(n_137357661), 
		.D(n_136857656), .Z(n_11722));
	notech_and4 i_716656(.A(n_135857646), .B(n_135757645), .C(n_136157649), 
		.D(n_135657644), .Z(n_11728));
	notech_and4 i_816657(.A(n_134657634), .B(n_134557633), .C(n_129357581), 
		.D(n_134957637), .Z(n_11734));
	notech_nand2 i_721298(.A(n_133957627), .B(n_133457622), .Z(n_20637));
	notech_ao4 i_126457918(.A(n_1845), .B(n_56574), .C(n_56104), .D(n_326546823
		), .Z(n_55115));
	notech_or2 i_117457872(.A(n_2255), .B(n_55961), .Z(n_249534121));
	notech_or2 i_120157871(.A(n_2255), .B(n_120857496), .Z(n_249434120));
	notech_or4 i_56657896(.A(calc_sz[3]), .B(calc_sz[0]), .C(n_260888755), .D
		(n_252034146), .Z(n_251934145));
	notech_nand3 i_17068(.A(n_26599), .B(n_56104), .C(n_57448), .Z(n_253034156
		));
	notech_and3 i_110257967(.A(n_26246), .B(n_132157609), .C(n_54711), .Z(n_55270
		));
	notech_or4 i_106857968(.A(n_205588858), .B(n_59370), .C(n_253034156), .D
		(n_59935), .Z(n_55302));
	notech_ao4 i_100957972(.A(n_54530), .B(n_55961), .C(n_56574), .D(n_55353
		), .Z(n_55355));
	notech_and2 i_98357973(.A(n_54718), .B(n_132357611), .Z(n_55380));
	notech_ao4 i_83557974(.A(n_54505), .B(n_55961), .C(n_55920), .D(eval_flag
		), .Z(n_55518));
	notech_and2 i_61057981(.A(n_46041), .B(n_55776), .Z(n_55740));
	notech_and4 i_143155327(.A(n_164757935), .B(n_164657934), .C(n_164257930
		), .D(n_164557933), .Z(n_57300));
	notech_or2 i_130160573(.A(n_323062234), .B(n_111757405), .Z(n_260436759)
		);
	notech_or2 i_117560580(.A(n_323062234), .B(n_56038), .Z(n_261136766));
	notech_and4 i_416653(.A(n_119357481), .B(n_119257480), .C(n_119157479), 
		.D(n_119657484), .Z(n_11710));
	notech_nand2 i_916658(.A(n_118557473), .B(n_118057468), .Z(n_11740));
	notech_and4 i_1016659(.A(n_117157459), .B(n_117057458), .C(n_114657434),
		 .D(n_117457462), .Z(n_11746));
	notech_and4 i_106660668(.A(n_55584), .B(n_56022), .C(n_54781), .D(n_115857446
		), .Z(n_55304));
	notech_and4 i_105360670(.A(n_225661327), .B(n_224461315), .C(n_54893), .D
		(n_316688523), .Z(n_55316));
	notech_or4 i_47560593(.A(n_60779), .B(n_60731), .C(n_1135), .D(n_60596),
		 .Z(n_262436779));
	notech_and2 i_94260681(.A(n_54710), .B(n_262436779), .Z(n_55421));
	notech_and2 i_94060682(.A(n_54774), .B(n_316788522), .Z(n_55422));
	notech_and2 i_39860714(.A(n_45486), .B(n_5538), .Z(n_55951));
	notech_ao3 i_118031899(.A(fsm[4]), .B(fsm[1]), .C(n_2585), .Z(n_316188528
		));
	notech_or2 i_119131888(.A(n_58904), .B(nbus_11326[15]), .Z(n_316088529)
		);
	notech_or4 i_119231887(.A(n_58945), .B(n_60494), .C(n_59935), .D(n_106813462
		), .Z(n_315988530));
	notech_and3 i_119431885(.A(sign_div), .B(opd[31]), .C(n_59935), .Z(n_315788532
		));
	notech_nand3 i_129931802(.A(n_57445), .B(n_275788700), .C(n_26377), .Z(n_315588534
		));
	notech_nand2 i_130031801(.A(n_275188706), .B(n_55641), .Z(n_315488535)
		);
	notech_nao3 i_168532827(.A(n_57441), .B(n_59935), .C(n_4737261), .Z(n_315388536
		));
	notech_ao4 i_143631679(.A(n_206688847), .B(n_55771), .C(n_55008), .D(n_190388902
		), .Z(n_315088539));
	notech_nand2 i_143831677(.A(n_57430), .B(n_26806), .Z(n_314988540));
	notech_ao4 i_143731678(.A(n_170914103), .B(n_2157), .C(n_55018), .D(n_213758422
		), .Z(n_314888541));
	notech_and4 i_144231673(.A(n_54777), .B(n_305088637), .C(n_328246806), .D
		(n_2983), .Z(n_314688543));
	notech_and4 i_144731668(.A(n_314288546), .B(n_2269), .C(n_2271), .D(n_313988549
		), .Z(n_314488544));
	notech_ao4 i_144631669(.A(n_56117), .B(n_106813462), .C(n_2253), .D(n_275488703
		), .Z(n_314288546));
	notech_or2 i_66132339(.A(n_55389), .B(n_55324), .Z(n_313988549));
	notech_ao4 i_60032395(.A(n_28140), .B(n_28413), .C(n_312388565), .D(n_26609
		), .Z(n_313488554));
	notech_or2 i_48732472(.A(n_310988579), .B(n_55578), .Z(n_313388555));
	notech_nao3 i_65832342(.A(pipe_mul[1]), .B(n_55159), .C(pipe_mul[0]), .Z
		(n_313088558));
	notech_or2 i_65432345(.A(n_2647), .B(n_2195), .Z(n_312988559));
	notech_and2 i_11032769(.A(n_312988559), .B(n_55640), .Z(n_312788561));
	notech_nor2 i_60132394(.A(n_55525), .B(n_59931), .Z(n_312388565));
	notech_and3 i_11932760(.A(n_57374), .B(n_1900), .C(n_57378), .Z(n_311588573
		));
	notech_ao4 i_11832761(.A(n_2258), .B(n_206188852), .C(n_26887), .D(n_311588573
		), .Z(n_311388575));
	notech_ao4 i_15932720(.A(n_58904), .B(n_48510), .C(n_2253), .D(n_55332),
		 .Z(n_310988579));
	notech_mux2 i_16032719(.S(n_56112), .A(n_56766), .B(n_58951), .Z(n_310588583
		));
	notech_or4 i_55532895(.A(n_2585), .B(n_2584), .C(n_315388536), .D(n_26613
		), .Z(n_310388585));
	notech_or4 i_55432896(.A(n_60752), .B(n_60739), .C(n_60779), .D(n_55838)
		, .Z(n_310288586));
	notech_or4 i_55232897(.A(n_4737261), .B(n_26377), .C(n_59845), .D(n_55641
		), .Z(n_310188587));
	notech_and3 i_205333715(.A(n_300188677), .B(n_309688592), .C(n_309888590
		), .Z(n_309988589));
	notech_ao4 i_205033718(.A(n_2987), .B(n_28590), .C(n_2323), .D(n_55331),
		 .Z(n_309888590));
	notech_ao4 i_205133717(.A(n_2156), .B(n_28802), .C(n_2319), .D(n_28555),
		 .Z(n_309688592));
	notech_and4 i_205833710(.A(n_309388595), .B(n_309188597), .C(n_300488675
		), .D(n_300788672), .Z(n_309588593));
	notech_ao4 i_205433714(.A(n_2164), .B(nbus_11326[1]), .C(n_54884), .D(nbus_11326
		[9]), .Z(n_309388595));
	notech_ao4 i_205633712(.A(n_55619), .B(n_28612), .C(n_2322), .D(n_56649)
		, .Z(n_309188597));
	notech_and4 i_207033699(.A(n_308688602), .B(n_308888600), .C(n_308588603
		), .D(n_301288669), .Z(n_309088598));
	notech_ao4 i_206133708(.A(n_55292), .B(\nbus_11276[9] ), .C(n_298688685)
		, .D(n_55328), .Z(n_308888600));
	notech_ao4 i_206233707(.A(n_2990), .B(n_27520), .C(n_2985), .D(n_357479919
		), .Z(n_308688602));
	notech_and4 i_206933700(.A(n_308388605), .B(n_308188607), .C(n_3015), .D
		(n_301888666), .Z(n_308588603));
	notech_ao4 i_206533704(.A(n_304188646), .B(n_27537), .C(n_304688641), .D
		(n_28404), .Z(n_308388605));
	notech_ao4 i_206733702(.A(n_304588642), .B(n_28831), .C(n_2213), .D(n_2984
		), .Z(n_308188607));
	notech_ao4 i_207233697(.A(n_26573), .B(n_29122), .C(n_60484), .D(n_27518
		), .Z(n_307988609));
	notech_and4 i_207633693(.A(n_330946790), .B(n_302488663), .C(n_307488613
		), .D(n_3021), .Z(n_307788611));
	notech_ao4 i_207433695(.A(n_2156), .B(n_28808), .C(n_2319), .D(n_28561),
		 .Z(n_307488613));
	notech_and3 i_208033689(.A(n_307088617), .B(n_307288615), .C(n_302988658
		), .Z(n_307388614));
	notech_ao4 i_207733692(.A(n_89513289), .B(n_27590), .C(nbus_11326[7]), .D
		(n_2164), .Z(n_307288615));
	notech_ao4 i_207833691(.A(n_55366), .B(n_28781), .C(n_55619), .D(n_28618
		), .Z(n_307088617));
	notech_and4 i_209033679(.A(n_306188626), .B(n_306388624), .C(n_303988648
		), .D(n_306888619), .Z(n_306988618));
	notech_ao3 i_208533684(.A(n_306588622), .B(n_306788620), .C(n_303488653)
		, .Z(n_306888619));
	notech_ao4 i_208233687(.A(n_88913283), .B(n_28837), .C(n_88813282), .D(n_28409
		), .Z(n_306788620));
	notech_ao4 i_208333686(.A(n_57351), .B(n_2320), .C(n_27526), .D(n_2990),
		 .Z(n_306588622));
	notech_ao4 i_208633683(.A(n_2989), .B(n_55400), .C(n_27534), .D(n_304288645
		), .Z(n_306388624));
	notech_ao4 i_208733682(.A(n_304088647), .B(n_27554), .C(n_2988), .D(n_28571
		), .Z(n_306188626));
	notech_or4 i_3335665(.A(fsm[3]), .B(fsm[0]), .C(n_60780), .D(n_57448), .Z
		(n_305988628));
	notech_nand2 i_3735661(.A(n_57448), .B(n_59845), .Z(n_305888629));
	notech_ao4 i_217733592(.A(n_1968), .B(n_2253), .C(n_1844), .D(n_2198), .Z
		(n_305588632));
	notech_and3 i_4235656(.A(mask8b[2]), .B(n_59931), .C(n_26862), .Z(n_305388634
		));
	notech_and4 i_7035628(.A(n_327246816), .B(n_54899), .C(n_48299), .D(n_304988638
		), .Z(n_305288635));
	notech_and2 i_115835686(.A(n_327246816), .B(n_54899), .Z(n_305088637));
	notech_ao4 i_4635652(.A(n_2253), .B(n_299688682), .C(n_1844), .D(n_56117
		), .Z(n_304988638));
	notech_or4 i_8135617(.A(n_59370), .B(n_60494), .C(n_274488713), .D(n_305888629
		), .Z(n_304688641));
	notech_or4 i_8335615(.A(n_59370), .B(n_60494), .C(n_274488713), .D(n_305988628
		), .Z(n_304588642));
	notech_nao3 i_7535623(.A(n_305388634), .B(mask8b[0]), .C(mask8b[1]), .Z(n_304288645
		));
	notech_nao3 i_8035618(.A(mask8b[1]), .B(n_305388634), .C(mask8b[0]), .Z(n_304188646
		));
	notech_nand3 i_8235616(.A(mask8b[1]), .B(n_305388634), .C(mask8b[0]), .Z
		(n_304088647));
	notech_or2 i_105634690(.A(n_304188646), .B(n_27545), .Z(n_303988648));
	notech_nor2 i_106134685(.A(n_2322), .B(n_57326), .Z(n_303488653));
	notech_or4 i_106634680(.A(n_244656264), .B(n_1844), .C(n_59931), .D(nbus_11326
		[15]), .Z(n_302988658));
	notech_nao3 i_107134675(.A(imm[39]), .B(n_26795), .C(n_2198), .Z(n_302488663
		));
	notech_or2 i_107234674(.A(n_2323), .B(n_27570), .Z(n_3021));
	notech_or2 i_103034714(.A(n_304088647), .B(n_27548), .Z(n_301888666));
	notech_or2 i_103334711(.A(n_304288645), .B(n_27528), .Z(n_3015));
	notech_or2 i_103734708(.A(n_57357), .B(n_2320), .Z(n_301288669));
	notech_nand2 i_104334703(.A(resb_shiftbox[1]), .B(n_26578), .Z(n_300788672
		));
	notech_or4 i_104634700(.A(n_275288705), .B(n_272588730), .C(n_59931), .D
		(n_27583), .Z(n_300488675));
	notech_nao3 i_104934697(.A(imm[33]), .B(n_26795), .C(n_2198), .Z(n_300188677
		));
	notech_and3 i_3835660(.A(n_274588712), .B(n_244656264), .C(n_56117), .Z(n_299688682
		));
	notech_nao3 i_113334614(.A(n_305388634), .B(n_27064), .C(mask8b[0]), .Z(n_2992
		));
	notech_or4 i_107334673(.A(n_1909), .B(n_2213), .C(n_28567), .D(n_60532),
		 .Z(n_2991));
	notech_and2 i_161135754(.A(n_55243), .B(n_2992), .Z(n_2990));
	notech_and4 i_40535753(.A(n_272288733), .B(n_54735), .C(n_305588632), .D
		(n_54910), .Z(n_2989));
	notech_and2 i_9235606(.A(n_55526), .B(n_2991), .Z(n_2988));
	notech_nao3 i_145939077(.A(n_239058636), .B(instrc[107]), .C(n_190688899
		), .Z(n_2987));
	notech_or2 i_32485(.A(n_57373), .B(n_2213), .Z(n_298688685));
	notech_and2 i_127935757(.A(n_272888727), .B(n_305288635), .Z(n_2985));
	notech_and3 i_9335605(.A(n_55087), .B(n_307988609), .C(n_56415), .Z(n_2984
		));
	notech_or4 i_5835640(.A(n_60494), .B(n_1844), .C(n_62395), .D(n_62437), 
		.Z(n_2983));
	notech_ao4 i_214937013(.A(n_89713291), .B(n_28589), .C(n_89513289), .D(n_27582
		), .Z(n_298288686));
	notech_ao4 i_214737015(.A(n_259158835), .B(n_2213), .C(n_2987), .D(n_28588
		), .Z(n_2980));
	notech_and4 i_214537017(.A(n_2970), .B(n_2969), .C(n_2968), .D(n_2974), 
		.Z(n_2976));
	notech_and3 i_214237020(.A(n_2972), .B(n_260658850), .C(n_260758851), .Z
		(n_2974));
	notech_ao4 i_213137031(.A(n_304688641), .B(n_28403), .C(n_304588642), .D
		(n_28830), .Z(n_2972));
	notech_ao4 i_213737025(.A(n_55619), .B(n_28611), .C(n_55366), .D(n_28769
		), .Z(n_2970));
	notech_ao4 i_213637026(.A(n_2164), .B(nbus_11326[0]), .C(n_2319), .D(n_28554
		), .Z(n_2969));
	notech_and4 i_214337019(.A(n_2966), .B(n_2965), .C(n_2963), .D(n_2962), 
		.Z(n_2968));
	notech_ao4 i_213537027(.A(n_2322), .B(nbus_11273[0]), .C(n_2156), .D(n_28801
		), .Z(n_2966));
	notech_ao4 i_213437028(.A(n_2323), .B(n_55342), .C(n_54884), .D(nbus_11326
		[8]), .Z(n_2965));
	notech_ao4 i_213337029(.A(n_55292), .B(n_55413), .C(n_304288645), .D(n_27527
		), .Z(n_2963));
	notech_ao4 i_213237030(.A(n_2990), .B(n_27519), .C(n_27546), .D(n_304088647
		), .Z(n_2962));
	notech_and4 i_210337059(.A(n_2956), .B(n_2959), .C(n_258458828), .D(n_258158825
		), .Z(n_2960));
	notech_ao4 i_210137061(.A(n_89513289), .B(n_27584), .C(n_88913283), .D(n_28832
		), .Z(n_2959));
	notech_and4 i_209637065(.A(n_2946), .B(n_2945), .C(n_2944), .D(n_2955), 
		.Z(n_2956));
	notech_and4 i_209537066(.A(n_2953), .B(n_2952), .C(n_2950), .D(n_2949), 
		.Z(n_2955));
	notech_ao4 i_208937072(.A(n_2164), .B(nbus_11326[2]), .C(n_2319), .D(n_28556
		), .Z(n_2953));
	notech_ao4 i_208837073(.A(n_2322), .B(n_56658), .C(n_2156), .D(n_28803),
		 .Z(n_2952));
	notech_ao4 i_208737074(.A(n_2323), .B(n_55299), .C(n_54884), .D(nbus_11326
		[10]), .Z(n_2950));
	notech_ao4 i_208637075(.A(n_55292), .B(n_55438), .C(n_304288645), .D(n_27529
		), .Z(n_2949));
	notech_ao4 i_208537076(.A(n_2989), .B(n_55289), .C(n_2990), .D(n_27521),
		 .Z(n_2946));
	notech_ao4 i_208437077(.A(n_304088647), .B(n_27549), .C(n_304188646), .D
		(n_27538), .Z(n_2945));
	notech_ao4 i_209037071(.A(n_55619), .B(n_28613), .C(n_55366), .D(n_28770
		), .Z(n_2944));
	notech_ao4 i_209937063(.A(n_256658810), .B(n_2213), .C(n_298688685), .D(n_123281220
		), .Z(n_2942));
	notech_ao4 i_205337107(.A(n_89713291), .B(n_28586), .C(n_89513289), .D(n_27585
		), .Z(n_2938));
	notech_ao4 i_205237108(.A(n_88913283), .B(n_28833), .C(n_88813282), .D(n_28405
		), .Z(n_2937));
	notech_and4 i_205137109(.A(n_255458798), .B(n_2932), .C(n_255558799), .D
		(n_255658800), .Z(n_2935));
	notech_and4 i_204837112(.A(n_2922), .B(n_2921), .C(n_2920), .D(n_2931), 
		.Z(n_2932));
	notech_and4 i_204737113(.A(n_2929), .B(n_2928), .C(n_2926), .D(n_2925), 
		.Z(n_2931));
	notech_ao4 i_204137119(.A(n_2164), .B(nbus_11326[3]), .C(n_2319), .D(n_28557
		), .Z(n_2929));
	notech_ao4 i_204037120(.A(n_2322), .B(nbus_11273[3]), .C(n_2156), .D(n_28804
		), .Z(n_2928));
	notech_ao4 i_203937121(.A(n_2323), .B(n_27564), .C(n_54884), .D(nbus_11326
		[11]), .Z(n_2926));
	notech_ao4 i_203837122(.A(n_55292), .B(n_55469), .C(n_304288645), .D(n_27530
		), .Z(n_2925));
	notech_ao4 i_203737123(.A(n_2989), .B(n_55277), .C(n_2990), .D(n_27522),
		 .Z(n_2922));
	notech_ao4 i_203637124(.A(n_304088647), .B(n_27550), .C(n_304188646), .D
		(n_27539), .Z(n_2921));
	notech_ao4 i_204237118(.A(n_55619), .B(n_28614), .C(n_55366), .D(n_28775
		), .Z(n_2920));
	notech_ao4 i_201037150(.A(n_88913283), .B(n_28834), .C(n_88813282), .D(n_28406
		), .Z(n_2918));
	notech_and4 i_200937151(.A(n_255458798), .B(n_2913), .C(n_2916), .D(n_253358777
		), .Z(n_2917));
	notech_ao4 i_200837152(.A(n_2987), .B(n_28583), .C(n_2320), .D(n_321188478
		), .Z(n_2916));
	notech_and4 i_200537155(.A(n_2903), .B(n_2902), .C(n_2901), .D(n_2912), 
		.Z(n_2913));
	notech_and4 i_200337156(.A(n_2910), .B(n_2909), .C(n_2907), .D(n_2906), 
		.Z(n_2912));
	notech_ao4 i_199737162(.A(n_2164), .B(nbus_11326[4]), .C(n_2319), .D(n_28558
		), .Z(n_2910));
	notech_ao4 i_199637163(.A(n_2322), .B(nbus_11273[4]), .C(n_2156), .D(n_28805
		), .Z(n_2909));
	notech_ao4 i_199537164(.A(n_2323), .B(n_58548), .C(n_54884), .D(nbus_11326
		[12]), .Z(n_2907));
	notech_ao4 i_199437165(.A(n_55292), .B(n_55542), .C(n_304288645), .D(n_27531
		), .Z(n_2906));
	notech_ao4 i_199337166(.A(n_2989), .B(\nbus_11276[4] ), .C(n_2990), .D(n_27523
		), .Z(n_2903));
	notech_ao4 i_199237167(.A(n_304088647), .B(n_27551), .C(n_304188646), .D
		(n_27540), .Z(n_2902));
	notech_ao4 i_199837161(.A(n_55619), .B(n_28615), .C(n_55366), .D(n_28778
		), .Z(n_2901));
	notech_ao4 i_201137149(.A(n_89713291), .B(n_28584), .C(n_89513289), .D(n_27586
		), .Z(n_2899));
	notech_ao4 i_196537193(.A(n_88913283), .B(n_28835), .C(n_88813282), .D(n_28407
		), .Z(n_289788687));
	notech_and4 i_196437194(.A(n_2893), .B(n_255458798), .C(n_251358757), .D
		(n_251458758), .Z(n_2896));
	notech_and4 i_196137197(.A(n_2883), .B(n_2882), .C(n_2881), .D(n_2892), 
		.Z(n_2893));
	notech_and4 i_196037198(.A(n_2890), .B(n_2889), .C(n_2887), .D(n_2886), 
		.Z(n_2892));
	notech_ao4 i_195437204(.A(n_2164), .B(nbus_11326[5]), .C(n_2319), .D(n_28559
		), .Z(n_2890));
	notech_ao4 i_195337205(.A(n_2322), .B(n_56685), .C(n_2156), .D(n_28806),
		 .Z(n_2889));
	notech_ao4 i_195237206(.A(n_2323), .B(n_27566), .C(n_54884), .D(nbus_11326
		[13]), .Z(n_2887));
	notech_ao4 i_195137207(.A(n_55292), .B(n_55552), .C(n_304288645), .D(n_27532
		), .Z(n_2886));
	notech_ao4 i_195037208(.A(n_2989), .B(n_55375), .C(n_2990), .D(n_27524),
		 .Z(n_2883));
	notech_ao4 i_194937209(.A(n_304088647), .B(n_27552), .C(n_304188646), .D
		(n_27541), .Z(n_2882));
	notech_ao4 i_195537203(.A(n_55619), .B(n_28616), .C(n_55366), .D(n_28779
		), .Z(n_2881));
	notech_ao4 i_196637192(.A(n_89713291), .B(n_28582), .C(n_89513289), .D(n_27588
		), .Z(n_2880));
	notech_ao4 i_192537233(.A(n_88913283), .B(n_28836), .C(n_88813282), .D(n_28408
		), .Z(n_287888688));
	notech_and4 i_192437234(.A(n_255458798), .B(n_2860), .C(n_249358737), .D
		(n_249458738), .Z(n_2865));
	notech_and4 i_192037237(.A(n_2843), .B(n_2842), .C(n_283859082), .D(n_2859
		), .Z(n_2860));
	notech_and4 i_191937238(.A(n_2852), .B(n_2851), .C(n_2848), .D(n_2847), 
		.Z(n_2859));
	notech_ao4 i_191337244(.A(n_54884), .B(nbus_11326[14]), .C(n_55619), .D(n_28617
		), .Z(n_2852));
	notech_ao4 i_191237245(.A(n_55366), .B(n_28780), .C(n_2164), .D(nbus_11326
		[6]), .Z(n_2851));
	notech_ao4 i_191137246(.A(n_2319), .B(n_28560), .C(n_2322), .D(nbus_11273
		[6]), .Z(n_2848));
	notech_ao4 i_191037247(.A(n_2156), .B(n_28807), .C(n_2323), .D(n_27568),
		 .Z(n_2847));
	notech_ao4 i_190937248(.A(n_2989), .B(\nbus_11276[6] ), .C(n_2990), .D(n_27525
		), .Z(n_2843));
	notech_ao4 i_190837249(.A(n_304088647), .B(n_27553), .C(n_27542), .D(n_304188646
		), .Z(n_2842));
	notech_ao4 i_191437243(.A(n_304288645), .B(n_27533), .C(n_55292), .D(n_55566
		), .Z(n_283859082));
	notech_ao4 i_192637232(.A(n_89713291), .B(n_28580), .C(n_89513289), .D(n_27589
		), .Z(n_283759081));
	notech_and4 i_188437273(.A(n_283259076), .B(n_247758721), .C(n_247358717
		), .D(n_247458718), .Z(n_283559079));
	notech_and4 i_188037277(.A(n_282359067), .B(n_282259066), .C(n_283059074
		), .D(n_36812763), .Z(n_283259076));
	notech_and4 i_187837279(.A(n_282859072), .B(n_282759071), .C(n_282559069
		), .D(n_247258716), .Z(n_283059074));
	notech_ao4 i_187237285(.A(n_2319), .B(n_29021), .C(n_2322), .D(n_56703),
		 .Z(n_282859072));
	notech_ao4 i_187137286(.A(n_2156), .B(n_28809), .C(n_2323), .D(n_27571),
		 .Z(n_282759071));
	notech_ao4 i_187037287(.A(n_54884), .B(\nbus_11276[24] ), .C(n_54735), .D
		(nbus_11326[0]), .Z(n_282559069));
	notech_ao4 i_187437283(.A(n_55526), .B(n_28579), .C(n_55366), .D(n_28782
		), .Z(n_282359067));
	notech_ao4 i_187337284(.A(n_55243), .B(n_27527), .C(n_2164), .D(nbus_11326
		[8]), .Z(n_282259066));
	notech_ao4 i_188337274(.A(n_89513289), .B(n_27592), .C(n_88913283), .D(n_28838
		), .Z(n_282159065));
	notech_and4 i_181637341(.A(n_281659060), .B(n_246058704), .C(n_245658700
		), .D(n_245758701), .Z(n_281959063));
	notech_and4 i_181237345(.A(n_280759051), .B(n_280659050), .C(n_281459058
		), .D(n_36812763), .Z(n_281659060));
	notech_and4 i_181037347(.A(n_281259056), .B(n_281159055), .C(n_280959053
		), .D(n_245558699), .Z(n_281459058));
	notech_ao4 i_180437353(.A(n_2319), .B(n_29015), .C(n_2322), .D(n_56721),
		 .Z(n_281259056));
	notech_ao4 i_180337354(.A(n_2156), .B(n_28811), .C(n_2323), .D(n_27575),
		 .Z(n_281159055));
	notech_ao4 i_180237355(.A(n_54884), .B(n_59337), .C(n_54735), .D(nbus_11326
		[2]), .Z(n_280959053));
	notech_ao4 i_180637351(.A(n_55526), .B(n_28578), .C(n_55366), .D(n_28784
		), .Z(n_280759051));
	notech_ao4 i_180537352(.A(n_55243), .B(n_27529), .C(n_2164), .D(nbus_11326
		[10]), .Z(n_280659050));
	notech_ao4 i_181537342(.A(n_89513289), .B(n_27594), .C(n_88913283), .D(n_28840
		), .Z(n_280559049));
	notech_and4 i_178237375(.A(n_280059044), .B(n_244358687), .C(n_243958683
		), .D(n_244058684), .Z(n_280359047));
	notech_and4 i_177837379(.A(n_279159035), .B(n_279059034), .C(n_279859042
		), .D(n_36812763), .Z(n_280059044));
	notech_and4 i_177637381(.A(n_279659040), .B(n_279559039), .C(n_279359037
		), .D(n_243858682), .Z(n_279859042));
	notech_ao4 i_176937387(.A(n_2319), .B(n_29018), .C(n_2322), .D(n_56730),
		 .Z(n_279659040));
	notech_ao4 i_176837388(.A(n_2156), .B(n_28812), .C(n_2323), .D(n_27576),
		 .Z(n_279559039));
	notech_ao4 i_1065658(.A(n_276588692), .B(n_56076), .C(n_58895), .D(n_2777
		), .Z(n_121477614));
	notech_or4 i_91064790(.A(n_275888699), .B(n_2205), .C(n_177560857), .D(n_26540
		), .Z(n_121777617));
	notech_or4 i_25363307(.A(n_56074), .B(n_56108), .C(n_55820), .D(n_319588494
		), .Z(n_121977619));
	notech_nand3 i_25263308(.A(n_54128), .B(tsc[36]), .C(n_59856), .Z(n_122277622
		));
	notech_or2 i_24763313(.A(n_2665), .B(n_55365), .Z(n_122777627));
	notech_nao3 i_31263249(.A(n_62427), .B(opc[9]), .C(n_320565522), .Z(n_123077630
		));
	notech_or2 i_30963252(.A(n_55382), .B(n_56712), .Z(n_123377633));
	notech_or4 i_30663255(.A(n_56158), .B(n_56108), .C(n_56345), .D(n_57299)
		, .Z(n_123677636));
	notech_or4 i_32563236(.A(n_59159), .B(n_26604), .C(n_26377), .D(n_27537)
		, .Z(n_124377643));
	notech_or2 i_32263239(.A(n_308518862), .B(nbus_11326[17]), .Z(n_124677646
		));
	notech_or2 i_31963242(.A(n_2700), .B(n_55442), .Z(n_124977649));
	notech_or2 i_35963205(.A(n_54748), .B(n_29063), .Z(n_125477654));
	notech_or2 i_35363210(.A(n_54921), .B(nbus_11273[4]), .Z(n_126177661));
	notech_ao3 i_74962823(.A(n_26564), .B(n_26418), .C(n_275388704), .Z(n_126277662
		));
	notech_ao4 i_117262415(.A(n_139770716), .B(n_55906), .C(n_55730), .D(n_58548
		), .Z(n_126577665));
	notech_ao4 i_117162416(.A(n_316288527), .B(n_248434110), .C(n_54920), .D
		(n_55365), .Z(n_126777667));
	notech_ao4 i_116962418(.A(n_54740), .B(n_321188478), .C(n_316388526), .D
		(n_248734113), .Z(n_126977669));
	notech_and3 i_117062417(.A(n_137970698), .B(n_126977669), .C(n_125477654
		), .Z(n_127177671));
	notech_ao4 i_114462443(.A(n_54066), .B(n_26957), .C(n_59195), .D(n_26702
		), .Z(n_127277672));
	notech_ao4 i_114362444(.A(n_2648), .B(n_55780), .C(n_55135), .D(n_27583)
		, .Z(n_127377673));
	notech_ao4 i_114162446(.A(n_55443), .B(n_28987), .C(n_55536), .D(n_56784
		), .Z(n_127577675));
	notech_and4 i_114662441(.A(n_127577675), .B(n_127377673), .C(n_127277672
		), .D(n_124977649), .Z(n_127777677));
	notech_ao4 i_113862449(.A(n_63826342), .B(n_308618863), .C(n_55535), .D(n_55600
		), .Z(n_127877678));
	notech_ao4 i_113662451(.A(n_54080), .B(n_28431), .C(n_54092), .D(n_29378
		), .Z(n_128077680));
	notech_and4 i_114062447(.A(n_128077680), .B(n_127877678), .C(n_124377643
		), .D(n_124677646), .Z(n_128277682));
	notech_ao4 i_113362454(.A(n_54066), .B(n_26941), .C(n_59195), .D(n_26694
		), .Z(n_128377683));
	notech_ao4 i_113262455(.A(n_54080), .B(n_28423), .C(n_54092), .D(n_29377
		), .Z(n_128477684));
	notech_ao4 i_113062457(.A(n_55738), .B(n_27574), .C(n_262536780), .D(n_27528
		), .Z(n_128677686));
	notech_and4 i_113562452(.A(n_123677636), .B(n_128677686), .C(n_128477684
		), .D(n_128377683), .Z(n_128877688));
	notech_ao4 i_112762460(.A(n_57349), .B(n_55519), .C(n_55520), .D(n_29048
		), .Z(n_128977689));
	notech_ao4 i_112262462(.A(n_352969301), .B(n_320665523), .C(n_55381), .D
		(n_55425), .Z(n_129177691));
	notech_and4 i_112962458(.A(n_123077630), .B(n_129177691), .C(n_128977689
		), .D(n_123377633), .Z(n_129377693));
	notech_ao4 i_107662508(.A(n_2666), .B(n_56676), .C(n_2687), .D(n_58548),
		 .Z(n_129477694));
	notech_ao4 i_107562509(.A(n_316388526), .B(n_2697), .C(n_316288527), .D(n_54606
		), .Z(n_129677696));
	notech_ao4 i_107262512(.A(n_2667), .B(n_29063), .C(n_321188478), .D(n_2668
		), .Z(n_129877698));
	notech_and4 i_107462510(.A(n_121977619), .B(n_129877698), .C(n_137377773
		), .D(n_122277622), .Z(n_130177701));
	notech_nand3 i_63359962(.A(n_59195), .B(n_59931), .C(read_data[6]), .Z(n_130277702
		));
	notech_nand3 i_17360382(.A(n_54124), .B(tsc[9]), .C(n_59856), .Z(n_130577705
		));
	notech_or2 i_17060385(.A(n_350965798), .B(n_57349), .Z(n_130877708));
	notech_or2 i_16760388(.A(n_350865797), .B(n_29048), .Z(n_131177711));
	notech_nand3 i_24060317(.A(n_54124), .B(tsc[38]), .C(n_59845), .Z(n_131477714
		));
	notech_or4 i_23660320(.A(n_56074), .B(n_56108), .C(n_55820), .D(n_57320)
		, .Z(n_131777717));
	notech_or2 i_23360323(.A(n_2666), .B(nbus_11273[6]), .Z(n_132077720));
	notech_nor2 i_28760271(.A(n_55085), .B(n_55888), .Z(n_132177721));
	notech_nor2 i_41460157(.A(n_161857906), .B(n_318231569), .Z(n_132877728)
		);
	notech_or2 i_40960162(.A(n_54943), .B(n_55413), .Z(n_133577735));
	notech_or4 i_50160078(.A(n_182758113), .B(n_56270), .C(n_317788512), .D(n_57352
		), .Z(n_134077740));
	notech_or2 i_49860081(.A(n_319288497), .B(n_27568), .Z(n_134377743));
	notech_or2 i_49560084(.A(n_318888501), .B(\nbus_11276[6] ), .Z(n_134677746
		));
	notech_nao3 i_54260040(.A(n_3404), .B(n_55450), .C(n_54707), .Z(n_135177751
		));
	notech_or2 i_53960043(.A(n_270688747), .B(n_302821915), .Z(n_135477754)
		);
	notech_or2 i_53660046(.A(n_271688739), .B(n_56892), .Z(n_135777757));
	notech_or4 i_71859882(.A(n_59370), .B(n_58895), .C(n_59931), .D(nbus_11326
		[9]), .Z(n_135877758));
	notech_or2 i_71359887(.A(n_54564), .B(n_55425), .Z(n_136577765));
	notech_or2 i_80959801(.A(n_54445), .B(n_57349), .Z(n_136677766));
	notech_or4 i_80359807(.A(n_56449), .B(n_56431), .C(n_353069302), .D(n_231778707
		), .Z(n_137177771));
	notech_and2 i_80459806(.A(n_215478548), .B(opb[9]), .Z(n_137277772));
	notech_mux2 i_31981(.S(n_59931), .A(n_249261520), .B(n_27523), .Z(n_137377773
		));
	notech_ao4 i_166059019(.A(n_325776096), .B(n_352969301), .C(n_56712), .D
		(n_215378547), .Z(n_137677776));
	notech_ao4 i_165859021(.A(n_54433), .B(n_29048), .C(n_55965), .D(n_55085
		), .Z(n_137877778));
	notech_nand3 i_165959020(.A(n_137877778), .B(n_26240), .C(n_136677766), 
		.Z(n_138077780));
	notech_or4 i_158859089(.A(n_56487), .B(n_56478), .C(n_56449), .D(n_353069302
		), .Z(n_138177781));
	notech_ao4 i_158559092(.A(n_178971108), .B(n_352969301), .C(n_54595), .D
		(n_138177781), .Z(n_138277782));
	notech_ao4 i_158459093(.A(n_54459), .B(n_29048), .C(n_54566), .D(n_56712
		), .Z(n_138477784));
	notech_ao4 i_158259095(.A(n_55085), .B(n_56382), .C(n_54441), .D(n_57349
		), .Z(n_138677786));
	notech_and3 i_158359094(.A(n_138677786), .B(n_26240), .C(n_135877758), .Z
		(n_138877788));
	notech_ao4 i_134759306(.A(n_271588740), .B(n_55249), .C(n_59193), .D(n_26739
		), .Z(n_139077790));
	notech_ao4 i_134559308(.A(n_55314), .B(n_28977), .C(n_57329), .D(n_55313
		), .Z(n_139277792));
	notech_and4 i_134959304(.A(n_139277792), .B(n_139077790), .C(n_135477754
		), .D(n_135777757), .Z(n_139477794));
	notech_ao4 i_134259311(.A(n_55133), .B(n_59104), .C(n_110923096), .D(n_302321910
		), .Z(n_139577795));
	notech_ao4 i_134059313(.A(n_320088489), .B(n_27597), .C(n_321688474), .D
		(n_29381), .Z(n_139777797));
	notech_and4 i_134459309(.A(n_139777797), .B(n_139577795), .C(n_45527), .D
		(n_135177751), .Z(n_139977799));
	notech_ao4 i_131059339(.A(n_320188488), .B(n_316588524), .C(n_59193), .D
		(n_26722), .Z(n_140077800));
	notech_ao4 i_130859341(.A(n_320688483), .B(n_316488525), .C(n_319088499)
		, .D(nbus_11273[6]), .Z(n_140277802));
	notech_and4 i_131259337(.A(n_140277802), .B(n_140077800), .C(n_134377743
		), .D(n_134677746), .Z(n_140477804));
	notech_ao4 i_130359344(.A(n_55222), .B(n_29068), .C(n_55688), .D(n_57320
		), .Z(n_140577805));
	notech_ao4 i_130059346(.A(n_321688474), .B(n_29380), .C(n_321788473), .D
		(n_29379), .Z(n_140777807));
	notech_and4 i_130259345(.A(n_144577845), .B(n_183678231), .C(n_140777807
		), .D(n_130277702), .Z(n_140877808));
	notech_ao4 i_122959414(.A(n_54944), .B(n_56703), .C(n_54902), .D(n_29045
		), .Z(n_141077810));
	notech_ao4 i_122859415(.A(n_27571), .B(n_55726), .C(n_57350), .D(n_54872
		), .Z(n_141277812));
	notech_nand3 i_123159412(.A(n_141077810), .B(n_141277812), .C(n_133577735
		), .Z(n_141377813));
	notech_ao4 i_122559417(.A(n_161957907), .B(n_318031567), .C(n_157974447)
		, .D(n_55906), .Z(n_141477814));
	notech_nao3 i_107559559(.A(n_56487), .B(n_268064997), .C(n_353069302), .Z
		(n_141777817));
	notech_ao4 i_107359561(.A(n_333669135), .B(n_352969301), .C(n_217778571)
		, .D(n_141777817), .Z(n_141877818));
	notech_ao4 i_107259562(.A(n_54946), .B(n_56712), .C(n_54945), .D(n_55425
		), .Z(n_141977819));
	notech_nand2 i_107459560(.A(n_141977819), .B(n_141877818), .Z(n_142077820
		));
	notech_ao4 i_107059564(.A(n_54852), .B(n_57349), .C(n_54853), .D(n_29048
		), .Z(n_142177821));
	notech_ao4 i_102259607(.A(n_2665), .B(\nbus_11276[6] ), .C(n_316588524),
		 .D(n_54606), .Z(n_142477824));
	notech_ao4 i_102059609(.A(n_2687), .B(n_27568), .C(n_316488525), .D(n_2697
		), .Z(n_142677826));
	notech_and4 i_102459605(.A(n_131777717), .B(n_142677826), .C(n_142477824
		), .D(n_132077720), .Z(n_142877828));
	notech_ao4 i_101759612(.A(n_57352), .B(n_2668), .C(n_2667), .D(n_29068),
		 .Z(n_142977829));
	notech_and4 i_101959610(.A(n_53844), .B(n_142977829), .C(n_54470), .D(n_131477714
		), .Z(n_143277832));
	notech_ao4 i_96159667(.A(n_336065662), .B(n_352969301), .C(n_353069302),
		 .D(n_26422), .Z(n_143377833));
	notech_ao4 i_95959669(.A(n_54572), .B(n_55425), .C(n_54573), .D(n_56712)
		, .Z(n_143577835));
	notech_and4 i_96359665(.A(n_143577835), .B(n_143377833), .C(n_130877708)
		, .D(n_131177711), .Z(n_143777837));
	notech_ao4 i_95659672(.A(n_61624), .B(nbus_11326[9]), .C(n_55085), .D(n_56023
		), .Z(n_143877838));
	notech_and4 i_95859670(.A(n_143877838), .B(n_55876), .C(n_130577705), .D
		(n_26240), .Z(n_144177841));
	notech_and2 i_66857892(.A(n_183578230), .B(n_183478229), .Z(n_144277842)
		);
	notech_or2 i_68557888(.A(n_55820), .B(n_57320), .Z(n_144377843));
	notech_or2 i_85257063(.A(n_316688523), .B(nbus_11273[6]), .Z(n_144577845
		));
	notech_ao4 i_188557854(.A(n_55854), .B(n_55387), .C(n_1135), .D(n_29068)
		, .Z(n_144677846));
	notech_and4 i_89557020(.A(n_55667), .B(n_293761941), .C(n_293161935), .D
		(n_55973), .Z(n_144977849));
	notech_or2 i_92656991(.A(n_55580), .B(n_55906), .Z(n_145077850));
	notech_ao3 i_7257786(.A(n_26763), .B(Daddrs_8[1]), .C(n_1908), .Z(n_145377853
		));
	notech_ao3 i_6957789(.A(n_316188528), .B(n_5154), .C(n_315388536), .Z(n_145677856
		));
	notech_and3 i_6557792(.A(n_361879963), .B(Daddrgs[1]), .C(n_59856), .Z(n_145977859
		));
	notech_or4 i_6057797(.A(n_60780), .B(n_60731), .C(n_358179926), .D(n_55331
		), .Z(n_146077860));
	notech_or4 i_6157796(.A(n_244656264), .B(n_2572), .C(n_274988708), .D(n_357479919
		), .Z(n_146177861));
	notech_or2 i_6257795(.A(n_55849), .B(n_28415), .Z(n_146277862));
	notech_ao3 i_8657773(.A(n_26763), .B(Daddrs_8[2]), .C(n_1908), .Z(n_146577865
		));
	notech_ao3 i_8357776(.A(n_316188528), .B(n_5155), .C(n_315388536), .Z(n_146877868
		));
	notech_and3 i_8057779(.A(n_361879963), .B(Daddrgs[2]), .C(n_59856), .Z(n_147177871
		));
	notech_nao3 i_9957760(.A(n_26763), .B(Daddrs_8[3]), .C(n_1908), .Z(n_147877878
		));
	notech_nao3 i_9657763(.A(n_6355), .B(n_59854), .C(n_55838), .Z(n_148177881
		));
	notech_nand3 i_9357766(.A(n_26498), .B(n_6356), .C(n_59854), .Z(n_148477884
		));
	notech_nao3 i_11257747(.A(n_26763), .B(Daddrs_8[4]), .C(n_1908), .Z(n_149177891
		));
	notech_nao3 i_10957750(.A(n_316188528), .B(n_5157), .C(n_315388536), .Z(n_149477894
		));
	notech_nand3 i_10657753(.A(n_361879963), .B(Daddrgs[4]), .C(n_59854), .Z
		(n_149777897));
	notech_nao3 i_12557734(.A(n_26763), .B(Daddrs_8[5]), .C(n_1908), .Z(n_150477904
		));
	notech_nao3 i_12257737(.A(n_6359), .B(n_59854), .C(n_55838), .Z(n_150777907
		));
	notech_nand3 i_11957740(.A(n_26498), .B(n_6360), .C(n_59854), .Z(n_151077910
		));
	notech_nao3 i_13857721(.A(n_26763), .B(Daddrs_8[6]), .C(n_1908), .Z(n_151777917
		));
	notech_nao3 i_13557724(.A(n_6361), .B(n_59854), .C(n_55838), .Z(n_152077920
		));
	notech_nand3 i_13257727(.A(n_26498), .B(n_6362), .C(n_59854), .Z(n_152377923
		));
	notech_nao3 i_15157708(.A(n_26763), .B(Daddrs_8[7]), .C(n_1908), .Z(n_153077930
		));
	notech_nao3 i_14857711(.A(n_6363), .B(n_59854), .C(n_55838), .Z(n_153377933
		));
	notech_nand3 i_14557714(.A(n_26498), .B(n_6364), .C(n_59854), .Z(n_153677936
		));
	notech_nao3 i_16457695(.A(n_26763), .B(Daddrs_8[8]), .C(n_1908), .Z(n_154377943
		));
	notech_nao3 i_16157698(.A(n_316188528), .B(n_5161), .C(n_315388536), .Z(n_154677946
		));
	notech_nand3 i_15857701(.A(Daddrgs[8]), .B(n_59854), .C(n_361879963), .Z
		(n_154977949));
	notech_nao3 i_17757682(.A(n_26763), .B(Daddrs_8[9]), .C(n_1908), .Z(n_155677956
		));
	notech_nand2 i_17457685(.A(Daddrs_1[9]), .B(n_26468), .Z(n_155977959));
	notech_nao3 i_17157688(.A(n_6367), .B(n_59856), .C(n_55838), .Z(n_156277962
		));
	notech_nao3 i_18957670(.A(n_26763), .B(Daddrs_8[10]), .C(n_1908), .Z(n_156977969
		));
	notech_nand2 i_18657673(.A(Daddrs_1[10]), .B(n_26468), .Z(n_157277972)
		);
	notech_nao3 i_18357676(.A(n_6369), .B(n_59856), .C(n_55838), .Z(n_157577975
		));
	notech_nand3 i_18057679(.A(n_26498), .B(n_6370), .C(n_59856), .Z(n_157877978
		));
	notech_nao3 i_20157658(.A(n_26763), .B(Daddrs_8[11]), .C(n_1908), .Z(n_158177981
		));
	notech_nand2 i_19857661(.A(Daddrs_1[11]), .B(n_26468), .Z(n_158477984)
		);
	notech_nao3 i_19557664(.A(n_6371), .B(n_59856), .C(n_55838), .Z(n_158777987
		));
	notech_nand3 i_19257667(.A(n_26498), .B(n_6372), .C(n_59854), .Z(n_159077990
		));
	notech_nao3 i_21357646(.A(n_26763), .B(Daddrs_8[12]), .C(n_1908), .Z(n_159377993
		));
	notech_nand2 i_21057649(.A(Daddrs_1[12]), .B(n_26468), .Z(n_159677996)
		);
	notech_nao3 i_20757652(.A(n_6373), .B(n_59854), .C(n_55838), .Z(n_159977999
		));
	notech_nand3 i_20457655(.A(n_26498), .B(n_6374), .C(n_59854), .Z(n_160278002
		));
	notech_nao3 i_22557634(.A(n_26763), .B(Daddrs_8[13]), .C(n_1908), .Z(n_160578005
		));
	notech_nand2 i_22257637(.A(Daddrs_1[13]), .B(n_26468), .Z(n_160878008)
		);
	notech_nao3 i_21957640(.A(n_6375), .B(n_59854), .C(n_55838), .Z(n_161178011
		));
	notech_nand3 i_21657643(.A(n_26498), .B(n_6376), .C(n_59854), .Z(n_161478014
		));
	notech_nao3 i_23857622(.A(n_26763), .B(Daddrs_8[14]), .C(n_1908), .Z(n_161778017
		));
	notech_nand2 i_23557625(.A(Daddrs_1[14]), .B(n_26468), .Z(n_162078020)
		);
	notech_nao3 i_23157628(.A(n_6377), .B(n_59789), .C(n_55838), .Z(n_162378023
		));
	notech_nand3 i_22857631(.A(n_26498), .B(n_6378), .C(n_59789), .Z(n_162678026
		));
	notech_nao3 i_25157610(.A(n_26763), .B(Daddrs_8[15]), .C(n_1908), .Z(n_162978029
		));
	notech_nand2 i_24857613(.A(Daddrs_1[15]), .B(n_26468), .Z(n_163278032)
		);
	notech_nao3 i_24457616(.A(n_6379), .B(n_59789), .C(n_55838), .Z(n_163578035
		));
	notech_nand3 i_24157619(.A(n_26498), .B(n_6380), .C(n_59789), .Z(n_163878038
		));
	notech_nao3 i_27557586(.A(n_26763), .B(Daddrs_8[17]), .C(n_1908), .Z(n_164178041
		));
	notech_nand2 i_27257589(.A(Daddrs_1[17]), .B(n_26468), .Z(n_164478044)
		);
	notech_nao3 i_26957592(.A(n_6383), .B(n_59789), .C(n_55838), .Z(n_164778047
		));
	notech_nand3 i_26657595(.A(n_26498), .B(n_6384), .C(n_59789), .Z(n_165078050
		));
	notech_nao3 i_28757574(.A(n_26763), .B(Daddrs_8[18]), .C(n_1908), .Z(n_165378053
		));
	notech_nand2 i_28457577(.A(Daddrs_1[18]), .B(n_26468), .Z(n_165678056)
		);
	notech_nao3 i_28157580(.A(n_6385), .B(n_59789), .C(n_55838), .Z(n_165978059
		));
	notech_nand3 i_27857583(.A(n_26498), .B(n_6386), .C(n_59789), .Z(n_166278062
		));
	notech_nao3 i_30057562(.A(n_26763), .B(Daddrs_8[19]), .C(n_55149), .Z(n_166578065
		));
	notech_nand2 i_29757565(.A(Daddrs_1[19]), .B(n_26468), .Z(n_166878068)
		);
	notech_nao3 i_29457568(.A(n_6387), .B(n_59789), .C(n_55838), .Z(n_167178071
		));
	notech_nand3 i_29057571(.A(n_26498), .B(n_6388), .C(n_59789), .Z(n_167478074
		));
	notech_nao3 i_31357550(.A(n_55040), .B(Daddrs_8[20]), .C(n_55149), .Z(n_167778077
		));
	notech_nand2 i_31057553(.A(Daddrs_1[20]), .B(n_26468), .Z(n_168078080)
		);
	notech_nao3 i_30757556(.A(n_6389), .B(n_59800), .C(n_58886), .Z(n_168378083
		));
	notech_nand3 i_30357559(.A(n_58591), .B(n_6390), .C(n_59800), .Z(n_168678086
		));
	notech_nao3 i_32557538(.A(n_55040), .B(Daddrs_8[21]), .C(n_55149), .Z(n_168978089
		));
	notech_nand2 i_32257541(.A(Daddrs_1[21]), .B(n_26468), .Z(n_169278092)
		);
	notech_nao3 i_31957544(.A(n_6391), .B(n_59800), .C(n_58886), .Z(n_169578095
		));
	notech_nand3 i_31657547(.A(n_58591), .B(n_6392), .C(n_59800), .Z(n_169878098
		));
	notech_nao3 i_33757526(.A(n_55040), .B(Daddrs_8[22]), .C(n_55149), .Z(n_170178101
		));
	notech_nand2 i_33457529(.A(Daddrs_1[22]), .B(n_54701), .Z(n_170478104)
		);
	notech_nao3 i_33157532(.A(n_6393), .B(n_59800), .C(n_58886), .Z(n_170778107
		));
	notech_nand3 i_32857535(.A(n_58591), .B(n_6394), .C(n_59789), .Z(n_171078110
		));
	notech_nao3 i_35157514(.A(n_55040), .B(Daddrs_8[23]), .C(n_55149), .Z(n_171378113
		));
	notech_nand2 i_34757517(.A(Daddrs_1[23]), .B(n_54701), .Z(n_171678116)
		);
	notech_nao3 i_34357520(.A(n_6395), .B(n_59789), .C(n_58886), .Z(n_171978119
		));
	notech_nand3 i_34057523(.A(n_58591), .B(n_6396), .C(n_59800), .Z(n_172278122
		));
	notech_nao3 i_36957502(.A(n_55040), .B(Daddrs_8[24]), .C(n_55149), .Z(n_172578125
		));
	notech_nand2 i_36557505(.A(Daddrs_1[24]), .B(n_54701), .Z(n_172878128)
		);
	notech_nao3 i_36157508(.A(n_6397), .B(n_59789), .C(n_58886), .Z(n_173178131
		));
	notech_nand3 i_35657511(.A(n_58591), .B(n_6398), .C(n_59789), .Z(n_173478134
		));
	notech_nao3 i_38157490(.A(n_55040), .B(Daddrs_8[25]), .C(n_55149), .Z(n_173778137
		));
	notech_nand2 i_37857493(.A(Daddrs_1[25]), .B(n_54701), .Z(n_174078140)
		);
	notech_nao3 i_37557496(.A(n_6399), .B(n_59809), .C(n_58886), .Z(n_174378143
		));
	notech_nand3 i_37257499(.A(n_58591), .B(n_6400), .C(n_59809), .Z(n_174678146
		));
	notech_nao3 i_39357478(.A(n_55040), .B(Daddrs_8[26]), .C(n_55149), .Z(n_174978149
		));
	notech_nand2 i_39057481(.A(Daddrs_1[26]), .B(n_54701), .Z(n_175278152)
		);
	notech_nao3 i_38757484(.A(n_6401), .B(n_59809), .C(n_58886), .Z(n_175578155
		));
	notech_nand3 i_38457487(.A(n_58591), .B(n_6402), .C(n_59809), .Z(n_175878158
		));
	notech_nao3 i_40557466(.A(n_55040), .B(Daddrs_8[27]), .C(n_55149), .Z(n_176178161
		));
	notech_nand2 i_40257469(.A(Daddrs_1[27]), .B(n_54701), .Z(n_176478164)
		);
	notech_nao3 i_39957472(.A(n_6403), .B(n_59809), .C(n_58886), .Z(n_176778167
		));
	notech_nand3 i_39657475(.A(n_58591), .B(n_6404), .C(n_59809), .Z(n_177078170
		));
	notech_nao3 i_41757454(.A(n_55040), .B(Daddrs_8[28]), .C(n_55149), .Z(n_177378173
		));
	notech_nand2 i_41457457(.A(Daddrs_1[28]), .B(n_54701), .Z(n_177678176)
		);
	notech_nao3 i_41157460(.A(n_6405), .B(n_59809), .C(n_58886), .Z(n_177978179
		));
	notech_nand3 i_40857463(.A(n_58591), .B(n_6406), .C(n_59809), .Z(n_178278182
		));
	notech_nao3 i_42957442(.A(n_55040), .B(Daddrs_8[29]), .C(n_55149), .Z(n_178578185
		));
	notech_nand2 i_42657445(.A(Daddrs_1[29]), .B(n_54701), .Z(n_178878188)
		);
	notech_nao3 i_42357448(.A(n_6407), .B(n_59809), .C(n_58886), .Z(n_179178191
		));
	notech_nand3 i_42057451(.A(n_58591), .B(n_6408), .C(n_59809), .Z(n_179478194
		));
	notech_nao3 i_44757430(.A(n_55040), .B(Daddrs_8[30]), .C(n_1908), .Z(n_179778197
		));
	notech_nand2 i_44157433(.A(Daddrs_1[30]), .B(n_54701), .Z(n_180078200)
		);
	notech_nao3 i_43857436(.A(n_6409), .B(n_59789), .C(n_58886), .Z(n_180378203
		));
	notech_nand3 i_43357439(.A(n_58591), .B(n_6410), .C(n_59809), .Z(n_180978206
		));
	notech_or4 i_59457290(.A(n_56240), .B(n_294061944), .C(n_55975), .D(n_57352
		), .Z(n_181078207));
	notech_or2 i_58857295(.A(n_55906), .B(n_144377843), .Z(n_181778214));
	notech_or4 i_78057133(.A(n_59370), .B(n_58895), .C(n_59931), .D(nbus_11326
		[6]), .Z(n_181878215));
	notech_nand2 i_77957134(.A(n_55752), .B(opd[6]), .Z(n_182178218));
	notech_or4 i_77257139(.A(n_59259), .B(n_59268), .C(n_56196), .D(n_144377843
		), .Z(n_182878223));
	notech_ao4 i_170156256(.A(n_55810), .B(nbus_11273[6]), .C(n_144677846), 
		.D(n_59931), .Z(n_183478229));
	notech_ao4 i_170056257(.A(n_27525), .B(n_59789), .C(n_55920), .D(n_57352
		), .Z(n_183578230));
	notech_ao4 i_168456273(.A(n_316788522), .B(n_57352), .C(n_144677846), .D
		(n_60474), .Z(n_183678231));
	notech_ao4 i_158856369(.A(n_247334099), .B(n_316488525), .C(n_247234098)
		, .D(n_316588524), .Z(n_183778232));
	notech_ao4 i_158756370(.A(n_54458), .B(n_57352), .C(n_54435), .D(n_29068
		), .Z(n_183978234));
	notech_ao4 i_158456373(.A(n_54565), .B(n_56694), .C(n_54563), .D(n_55387
		), .Z(n_184178236));
	notech_and4 i_158656371(.A(n_144277842), .B(n_184178236), .C(n_181878215
		), .D(n_182178218), .Z(n_184478239));
	notech_ao4 i_140956540(.A(n_316488525), .B(n_248734113), .C(n_316588524)
		, .D(n_248434110), .Z(n_184578240));
	notech_ao4 i_140856541(.A(n_56694), .B(n_54921), .C(n_54920), .D(n_55387
		), .Z(n_184778242));
	notech_ao4 i_140656543(.A(n_29068), .B(n_54748), .C(n_27568), .D(n_55730
		), .Z(n_184978244));
	notech_and4 i_140756542(.A(n_183578230), .B(n_183478229), .C(n_184978244
		), .D(n_181078207), .Z(n_185178246));
	notech_ao4 i_125756674(.A(n_55848), .B(n_27983), .C(n_55849), .D(n_28444
		), .Z(n_185278247));
	notech_ao4 i_125556676(.A(n_310188587), .B(n_28498), .C(n_358079925), .D
		(n_27294), .Z(n_185478249));
	notech_and4 i_125956672(.A(n_185478249), .B(n_185278247), .C(n_180378203
		), .D(n_180978206), .Z(n_185678251));
	notech_ao4 i_125256679(.A(n_55793), .B(n_59050), .C(n_310388585), .D(n_29415
		), .Z(n_185778252));
	notech_ao4 i_125056681(.A(n_55787), .B(n_55234), .C(n_55788), .D(n_27599
		), .Z(n_185978254));
	notech_and4 i_125456677(.A(n_185978254), .B(n_185778252), .C(n_180078200
		), .D(n_179778197), .Z(n_186178256));
	notech_ao4 i_124756684(.A(n_55848), .B(n_27982), .C(n_55849), .D(n_28443
		), .Z(n_186278257));
	notech_ao4 i_124556686(.A(n_310188587), .B(n_28497), .C(n_358079925), .D
		(n_27293), .Z(n_186478259));
	notech_and4 i_124956682(.A(n_186478259), .B(n_186278257), .C(n_179178191
		), .D(n_179478194), .Z(n_186678261));
	notech_ao4 i_124256689(.A(n_55793), .B(n_59104), .C(n_310388585), .D(n_29414
		), .Z(n_186778262));
	notech_ao4 i_124056691(.A(n_55787), .B(n_55249), .C(n_55788), .D(n_27597
		), .Z(n_186978264));
	notech_and4 i_124456687(.A(n_186978264), .B(n_186778262), .C(n_178878188
		), .D(n_178578185), .Z(n_187178266));
	notech_ao4 i_123756694(.A(n_55848), .B(n_27981), .C(n_55849), .D(n_28442
		), .Z(n_187278267));
	notech_ao4 i_123556696(.A(n_310188587), .B(n_28496), .C(n_358079925), .D
		(n_27292), .Z(n_187478269));
	notech_and4 i_123956692(.A(n_187478269), .B(n_187278267), .C(n_177978179
		), .D(n_178278182), .Z(n_187678271));
	notech_ao4 i_123256699(.A(n_55793), .B(nbus_11326[28]), .C(n_310388585),
		 .D(n_29413), .Z(n_187778272));
	notech_ao4 i_123056701(.A(n_55787), .B(n_55261), .C(n_55788), .D(n_27596
		), .Z(n_187978274));
	notech_and4 i_123456697(.A(n_187978274), .B(n_187778272), .C(n_177678176
		), .D(n_177378173), .Z(n_188178276));
	notech_ao4 i_122756704(.A(n_55848), .B(n_27980), .C(n_55849), .D(n_28441
		), .Z(n_188278277));
	notech_ao4 i_122556706(.A(n_310188587), .B(n_28495), .C(n_358079925), .D
		(n_27291), .Z(n_188478279));
	notech_and4 i_122956702(.A(n_188478279), .B(n_188278277), .C(n_176778167
		), .D(n_177078170), .Z(n_188678281));
	notech_ao4 i_122256709(.A(n_55793), .B(nbus_11326[27]), .C(n_310388585),
		 .D(n_29412), .Z(n_188778282));
	notech_ao4 i_122056711(.A(n_55787), .B(n_59328), .C(n_55788), .D(n_27595
		), .Z(n_188978284));
	notech_and4 i_122456707(.A(n_188978284), .B(n_188778282), .C(n_176478164
		), .D(n_176178161), .Z(n_189178286));
	notech_ao4 i_121756714(.A(n_55848), .B(n_27979), .C(n_55849), .D(n_28440
		), .Z(n_189278287));
	notech_ao4 i_121556716(.A(n_310188587), .B(n_28494), .C(n_358079925), .D
		(n_27290), .Z(n_189478289));
	notech_and4 i_121956712(.A(n_189478289), .B(n_189278287), .C(n_175578155
		), .D(n_175878158), .Z(n_189678291));
	notech_ao4 i_121256719(.A(n_55793), .B(n_59068), .C(n_310388585), .D(n_29411
		), .Z(n_189778292));
	notech_ao4 i_121056721(.A(n_55787), .B(n_59337), .C(n_55788), .D(n_27594
		), .Z(n_189978294));
	notech_and4 i_121456717(.A(n_189978294), .B(n_189778292), .C(n_175278152
		), .D(n_174978149), .Z(n_190178296));
	notech_ao4 i_120756724(.A(n_55848), .B(n_27978), .C(n_55849), .D(n_28439
		), .Z(n_190278297));
	notech_ao4 i_120556726(.A(n_310188587), .B(n_28493), .C(n_358079925), .D
		(n_27289), .Z(n_190478299));
	notech_and4 i_120956722(.A(n_190478299), .B(n_190278297), .C(n_174378143
		), .D(n_174678146), .Z(n_190678301));
	notech_ao4 i_120256729(.A(n_55793), .B(nbus_11326[25]), .C(n_310388585),
		 .D(n_29410), .Z(n_190778302));
	notech_ao4 i_119956731(.A(n_55787), .B(n_59346), .C(n_55788), .D(n_27593
		), .Z(n_190978304));
	notech_and4 i_120456727(.A(n_190978304), .B(n_190778302), .C(n_174078140
		), .D(n_173778137), .Z(n_191178306));
	notech_ao4 i_119656734(.A(n_55848), .B(n_27977), .C(n_55849), .D(n_28438
		), .Z(n_191278307));
	notech_ao4 i_119456736(.A(n_310188587), .B(n_28492), .C(n_358079925), .D
		(n_27288), .Z(n_191478309));
	notech_and4 i_119856732(.A(n_191478309), .B(n_191278307), .C(n_173178131
		), .D(n_173478134), .Z(n_191678311));
	notech_ao4 i_119156739(.A(n_55793), .B(nbus_11326[24]), .C(n_310388585),
		 .D(n_29409), .Z(n_191778312));
	notech_ao4 i_118956741(.A(n_55787), .B(n_56207), .C(n_55788), .D(n_27592
		), .Z(n_191978314));
	notech_and4 i_119356737(.A(n_191978314), .B(n_191778312), .C(n_172878128
		), .D(n_172578125), .Z(n_192178316));
	notech_ao4 i_118656744(.A(n_55848), .B(n_27976), .C(n_55849), .D(n_28437
		), .Z(n_192278317));
	notech_ao4 i_118456746(.A(n_310188587), .B(n_28491), .C(n_358079925), .D
		(n_27287), .Z(n_192478319));
	notech_and4 i_118856742(.A(n_192478319), .B(n_192278317), .C(n_171978119
		), .D(n_172278122), .Z(n_192678321));
	notech_ao4 i_118156749(.A(n_55793), .B(nbus_11326[23]), .C(n_310388585),
		 .D(n_29408), .Z(n_192778322));
	notech_ao4 i_117956751(.A(n_55787), .B(\nbus_11276[23] ), .C(n_55788), .D
		(n_27590), .Z(n_192978324));
	notech_and4 i_118356747(.A(n_192978324), .B(n_192778322), .C(n_171678116
		), .D(n_171378113), .Z(n_193178326));
	notech_ao4 i_117656754(.A(n_55848), .B(n_27975), .C(n_55849), .D(n_28436
		), .Z(n_193278327));
	notech_ao4 i_117356756(.A(n_310188587), .B(n_28490), .C(n_358079925), .D
		(n_27286), .Z(n_193478329));
	notech_and4 i_117856752(.A(n_193478329), .B(n_193278327), .C(n_170778107
		), .D(n_171078110), .Z(n_193678331));
	notech_ao4 i_117056759(.A(n_55793), .B(nbus_11326[22]), .C(n_310388585),
		 .D(n_29407), .Z(n_193778332));
	notech_ao4 i_116856761(.A(n_55787), .B(n_55647), .C(n_55788), .D(n_27589
		), .Z(n_193978334));
	notech_and4 i_117256757(.A(n_193978334), .B(n_193778332), .C(n_170478104
		), .D(n_170178101), .Z(n_194178336));
	notech_ao4 i_116356764(.A(n_55848), .B(n_27974), .C(n_55849), .D(n_28435
		), .Z(n_194278337));
	notech_ao4 i_116156766(.A(n_310188587), .B(n_28489), .C(n_358079925), .D
		(n_27285), .Z(n_194478339));
	notech_and4 i_116656762(.A(n_194478339), .B(n_194278337), .C(n_169578095
		), .D(n_169878098), .Z(n_194678341));
	notech_ao4 i_115856769(.A(n_55793), .B(nbus_11326[21]), .C(n_310388585),
		 .D(n_29406), .Z(n_194778342));
	notech_ao4 i_115556771(.A(n_55787), .B(\nbus_11276[21] ), .C(n_55788), .D
		(n_27588), .Z(n_194978344));
	notech_and4 i_116056767(.A(n_194978344), .B(n_194778342), .C(n_169278092
		), .D(n_168978089), .Z(n_195178346));
	notech_ao4 i_115256774(.A(n_55848), .B(n_27973), .C(n_55849), .D(n_28434
		), .Z(n_195278347));
	notech_ao4 i_115056776(.A(n_310188587), .B(n_28488), .C(n_358079925), .D
		(n_27284), .Z(n_195478349));
	notech_and4 i_115456772(.A(n_195478349), .B(n_195278347), .C(n_168378083
		), .D(n_168678086), .Z(n_195678351));
	notech_ao4 i_114756779(.A(n_55793), .B(nbus_11326[20]), .C(n_310388585),
		 .D(n_29405), .Z(n_195778352));
	notech_ao4 i_114556781(.A(n_55787), .B(\nbus_11276[20] ), .C(n_55788), .D
		(n_27586), .Z(n_195978354));
	notech_and4 i_114956777(.A(n_195978354), .B(n_195778352), .C(n_168078080
		), .D(n_167778077), .Z(n_196178356));
	notech_ao4 i_114256784(.A(n_55848), .B(n_27972), .C(n_55849), .D(n_28433
		), .Z(n_196278357));
	notech_ao4 i_114056786(.A(n_310188587), .B(n_28487), .C(n_358079925), .D
		(n_27283), .Z(n_196478359));
	notech_and4 i_114456782(.A(n_196478359), .B(n_196278357), .C(n_167178071
		), .D(n_167478074), .Z(n_196678361));
	notech_ao4 i_113756789(.A(n_55793), .B(nbus_11326[19]), .C(n_310388585),
		 .D(n_29404), .Z(n_196778362));
	notech_ao4 i_113556791(.A(n_55787), .B(\nbus_11276[19] ), .C(n_55788), .D
		(n_27585), .Z(n_196978364));
	notech_and4 i_113956787(.A(n_196978364), .B(n_196778362), .C(n_166878068
		), .D(n_166578065), .Z(n_197178366));
	notech_ao4 i_113256794(.A(n_55848), .B(n_27971), .C(n_55849), .D(n_28432
		), .Z(n_197278367));
	notech_ao4 i_113056796(.A(n_310188587), .B(n_28486), .C(n_358079925), .D
		(n_27282), .Z(n_197478369));
	notech_and4 i_113456792(.A(n_197478369), .B(n_197278367), .C(n_165978059
		), .D(n_166278062), .Z(n_197678371));
	notech_ao4 i_112756799(.A(n_55793), .B(nbus_11326[18]), .C(n_310388585),
		 .D(n_29403), .Z(n_197778372));
	notech_ao4 i_112556801(.A(n_55787), .B(\nbus_11276[18] ), .C(n_55788), .D
		(n_27584), .Z(n_197978374));
	notech_and4 i_112956797(.A(n_197978374), .B(n_197778372), .C(n_165678056
		), .D(n_165378053), .Z(n_198178376));
	notech_ao4 i_112256804(.A(n_55848), .B(n_27970), .C(n_55849), .D(n_28431
		), .Z(n_198278377));
	notech_ao4 i_112056806(.A(n_310188587), .B(n_28481), .C(n_358079925), .D
		(n_27281), .Z(n_198478379));
	notech_and4 i_112456802(.A(n_198478379), .B(n_198278377), .C(n_164778047
		), .D(n_165078050), .Z(n_198678381));
	notech_ao4 i_111756809(.A(n_55793), .B(nbus_11326[17]), .C(n_310388585),
		 .D(n_29402), .Z(n_198778382));
	notech_ao4 i_111556811(.A(n_55787), .B(n_55600), .C(n_55788), .D(n_27583
		), .Z(n_198978384));
	notech_and4 i_111956807(.A(n_198978384), .B(n_198778382), .C(n_164478044
		), .D(n_164178041), .Z(n_199178386));
	notech_ao4 i_110056824(.A(n_55848), .B(n_27968), .C(n_55849), .D(n_28429
		), .Z(n_199278387));
	notech_ao4 i_109856826(.A(n_310188587), .B(n_28476), .C(n_58523), .D(n_27279
		), .Z(n_199478389));
	notech_and4 i_110356822(.A(n_199478389), .B(n_199278387), .C(n_163578035
		), .D(n_163878038), .Z(n_199678391));
	notech_ao4 i_109556829(.A(n_55793), .B(nbus_11326[15]), .C(n_54714), .D(n_29401
		), .Z(n_199778392));
	notech_ao4 i_109356831(.A(n_55787), .B(n_55578), .C(n_55788), .D(n_27581
		), .Z(n_199978394));
	notech_and4 i_109756827(.A(n_199978394), .B(n_199778392), .C(n_163278032
		), .D(n_162978029), .Z(n_200178396));
	notech_ao4 i_109056834(.A(n_55848), .B(n_27967), .C(n_54659), .D(n_28428
		), .Z(n_200278397));
	notech_ao4 i_108856836(.A(n_310188587), .B(n_28475), .C(n_58523), .D(n_27278
		), .Z(n_200478399));
	notech_and4 i_109256832(.A(n_200478399), .B(n_200278397), .C(n_162378023
		), .D(n_162678026), .Z(n_200678401));
	notech_ao4 i_108556839(.A(n_55793), .B(nbus_11326[14]), .C(n_54714), .D(n_29400
		), .Z(n_200778402));
	notech_ao4 i_108356841(.A(n_54771), .B(n_55566), .C(n_54742), .D(n_27579
		), .Z(n_200978404));
	notech_and4 i_108756837(.A(n_200978404), .B(n_200778402), .C(n_162078020
		), .D(n_161778017), .Z(n_201178406));
	notech_ao4 i_108056844(.A(n_54674), .B(n_27966), .C(n_54659), .D(n_28427
		), .Z(n_201278407));
	notech_ao4 i_107856846(.A(n_54685), .B(n_28474), .C(n_58523), .D(n_27277
		), .Z(n_201478409));
	notech_and4 i_108256842(.A(n_201478409), .B(n_201278407), .C(n_161178011
		), .D(n_161478014), .Z(n_201678411));
	notech_ao4 i_107556849(.A(n_54727), .B(nbus_11326[13]), .C(n_54714), .D(n_29399
		), .Z(n_201778412));
	notech_ao4 i_107356851(.A(n_54771), .B(n_55552), .C(n_54742), .D(n_27578
		), .Z(n_201978414));
	notech_and4 i_107756847(.A(n_201978414), .B(n_201778412), .C(n_160878008
		), .D(n_160578005), .Z(n_202178416));
	notech_ao4 i_107056854(.A(n_54674), .B(n_27965), .C(n_54659), .D(n_28426
		), .Z(n_202278417));
	notech_ao4 i_106756856(.A(n_54685), .B(n_28470), .C(n_58523), .D(n_27276
		), .Z(n_202478419));
	notech_and4 i_107256852(.A(n_202478419), .B(n_202278417), .C(n_159977999
		), .D(n_160278002), .Z(n_202678421));
	notech_ao4 i_106456859(.A(n_54727), .B(nbus_11326[12]), .C(n_54714), .D(n_29398
		), .Z(n_202778422));
	notech_ao4 i_106256861(.A(n_54771), .B(n_55542), .C(n_54742), .D(n_27577
		), .Z(n_202978424));
	notech_and4 i_106656857(.A(n_202978424), .B(n_202778422), .C(n_159677996
		), .D(n_159377993), .Z(n_203178426));
	notech_ao4 i_105856864(.A(n_54674), .B(n_27964), .C(n_54659), .D(n_28425
		), .Z(n_203278427));
	notech_ao4 i_105656866(.A(n_54685), .B(n_28469), .C(n_58523), .D(n_27275
		), .Z(n_203478429));
	notech_and4 i_106156862(.A(n_203478429), .B(n_203278427), .C(n_158777987
		), .D(n_159077990), .Z(n_203678431));
	notech_ao4 i_105356869(.A(n_54727), .B(nbus_11326[11]), .C(n_54714), .D(n_29397
		), .Z(n_203778432));
	notech_ao4 i_105156871(.A(n_54771), .B(n_55469), .C(n_54742), .D(n_27576
		), .Z(n_203978434));
	notech_and4 i_105556867(.A(n_203978434), .B(n_203778432), .C(n_158477984
		), .D(n_158177981), .Z(n_204178436));
	notech_ao4 i_104856874(.A(n_54674), .B(n_27963), .C(n_54659), .D(n_28424
		), .Z(n_204278437));
	notech_ao4 i_104656876(.A(n_54685), .B(n_28468), .C(n_58523), .D(n_27274
		), .Z(n_204478439));
	notech_and4 i_105056872(.A(n_204478439), .B(n_204278437), .C(n_157577975
		), .D(n_157877978), .Z(n_204678441));
	notech_ao4 i_104356879(.A(n_54727), .B(nbus_11326[10]), .C(n_54714), .D(n_29396
		), .Z(n_204778442));
	notech_ao4 i_104156881(.A(n_54771), .B(n_55438), .C(n_54742), .D(n_27575
		), .Z(n_204978444));
	notech_and4 i_104556877(.A(n_204978444), .B(n_204778442), .C(n_157277972
		), .D(n_156977969), .Z(n_205178446));
	notech_ao4 i_103856884(.A(n_54659), .B(n_28423), .C(n_55684), .D(n_27570
		), .Z(n_205278447));
	notech_ao4 i_103756885(.A(n_2234), .B(n_29395), .C(n_54674), .D(n_27962)
		, .Z(n_205378448));
	notech_ao4 i_103556887(.A(n_54685), .B(n_28467), .C(n_58523), .D(n_27273
		), .Z(n_205578450));
	notech_and4 i_104056882(.A(n_205578450), .B(n_205378448), .C(n_205278447
		), .D(n_156277962), .Z(n_205778452));
	notech_ao4 i_103256890(.A(n_54727), .B(nbus_11326[9]), .C(n_54714), .D(n_29394
		), .Z(n_205878453));
	notech_ao4 i_103056892(.A(n_54771), .B(n_55425), .C(n_54742), .D(n_27574
		), .Z(n_206078455));
	notech_and4 i_103456888(.A(n_206078455), .B(n_205878453), .C(n_155977959
		), .D(n_155677956), .Z(n_206278457));
	notech_ao4 i_102756895(.A(n_54742), .B(n_27571), .C(n_55684), .D(n_27568
		), .Z(n_206378458));
	notech_ao4 i_102656896(.A(n_54659), .B(n_28422), .C(n_54771), .D(n_55413
		), .Z(n_206478459));
	notech_ao4 i_102456898(.A(n_2234), .B(n_29393), .C(n_54674), .D(n_27961)
		, .Z(n_206678461));
	notech_and4 i_102956893(.A(n_206678461), .B(n_206478459), .C(n_206378458
		), .D(n_154977949), .Z(n_206878463));
	notech_ao4 i_102156901(.A(n_310288586), .B(n_29392), .C(n_54685), .D(n_28466
		), .Z(n_206978464));
	notech_ao4 i_101956903(.A(n_55792), .B(n_28453), .C(n_54727), .D(nbus_11326
		[8]), .Z(n_207178466));
	notech_and4 i_102356899(.A(n_207178466), .B(n_206978464), .C(n_154377943
		), .D(n_154677946), .Z(n_207378468));
	notech_ao4 i_101656906(.A(n_54771), .B(n_55400), .C(n_55684), .D(n_27566
		), .Z(n_207478469));
	notech_ao4 i_101556907(.A(n_54727), .B(nbus_11326[7]), .C(n_54742), .D(n_27570
		), .Z(n_207578470));
	notech_ao4 i_101356909(.A(n_54674), .B(n_27960), .C(n_54659), .D(n_28421
		), .Z(n_207778472));
	notech_and4 i_101856904(.A(n_207778472), .B(n_207578470), .C(n_207478469
		), .D(n_153677936), .Z(n_207978474));
	notech_ao4 i_100756912(.A(n_54685), .B(n_28464), .C(n_58523), .D(n_27272
		), .Z(n_208078475));
	notech_ao4 i_100556914(.A(n_55792), .B(n_28452), .C(n_54714), .D(n_29391
		), .Z(n_208278477));
	notech_and4 i_101156910(.A(n_208278477), .B(n_208078475), .C(n_153377933
		), .D(n_153077930), .Z(n_208478479));
	notech_ao4 i_100256917(.A(n_54771), .B(n_55387), .C(n_55684), .D(n_58548
		), .Z(n_208578480));
	notech_ao4 i_100156918(.A(n_54742), .B(n_27568), .C(n_54727), .D(nbus_11326
		[6]), .Z(n_208678481));
	notech_ao4 i_99956920(.A(n_54674), .B(n_27959), .C(n_54659), .D(n_28420)
		, .Z(n_208878483));
	notech_and4 i_100456915(.A(n_208878483), .B(n_208678481), .C(n_208578480
		), .D(n_152377923), .Z(n_209078485));
	notech_ao4 i_99656923(.A(n_54685), .B(n_28463), .C(n_58523), .D(n_27271)
		, .Z(n_209178486));
	notech_ao4 i_99456925(.A(n_55792), .B(n_28451), .C(n_54714), .D(n_29390)
		, .Z(n_209378488));
	notech_and4 i_99856921(.A(n_209378488), .B(n_209178486), .C(n_152077920)
		, .D(n_151777917), .Z(n_209578490));
	notech_ao4 i_99156928(.A(n_54771), .B(n_55375), .C(n_55684), .D(n_27564)
		, .Z(n_209678491));
	notech_ao4 i_99056929(.A(nbus_11326[5]), .B(n_54727), .C(n_27566), .D(n_54742
		), .Z(n_209778492));
	notech_ao4 i_98856931(.A(n_54674), .B(n_27958), .C(n_54659), .D(n_28419)
		, .Z(n_209978494));
	notech_and4 i_99356926(.A(n_209978494), .B(n_209778492), .C(n_209678491)
		, .D(n_151077910), .Z(n_210178496));
	notech_ao4 i_98556934(.A(n_54685), .B(n_28462), .C(n_358079925), .D(n_27270
		), .Z(n_210278497));
	notech_ao4 i_98256936(.A(n_55792), .B(n_28450), .C(n_310388585), .D(n_29389
		), .Z(n_210478499));
	notech_and4 i_98756932(.A(n_210478499), .B(n_210278497), .C(n_150777907)
		, .D(n_150477904), .Z(n_210678501));
	notech_ao4 i_97956939(.A(n_54771), .B(n_55365), .C(n_55684), .D(n_55299)
		, .Z(n_210778502));
	notech_ao4 i_97856940(.A(n_54659), .B(n_28418), .C(n_54742), .D(n_58548)
		, .Z(n_210878503));
	notech_ao4 i_97656942(.A(n_2234), .B(n_29388), .C(n_54674), .D(n_27957),
		 .Z(n_211078505));
	notech_and4 i_98156937(.A(n_211078505), .B(n_210878503), .C(n_210778502)
		, .D(n_149777897), .Z(n_211278507));
	notech_ao4 i_97356945(.A(n_310288586), .B(n_29387), .C(n_54685), .D(n_28461
		), .Z(n_211378508));
	notech_ao4 i_97156947(.A(n_55792), .B(n_28449), .C(n_54727), .D(nbus_11326
		[4]), .Z(n_211578510));
	notech_and4 i_97556943(.A(n_211578510), .B(n_211378508), .C(n_149177891)
		, .D(n_149477894), .Z(n_211778512));
	notech_ao4 i_96856950(.A(n_54771), .B(n_55277), .C(n_55684), .D(n_55331)
		, .Z(n_211878513));
	notech_ao4 i_96756951(.A(n_54727), .B(nbus_11326[3]), .C(n_54742), .D(n_27564
		), .Z(n_211978514));
	notech_ao4 i_96556953(.A(n_54674), .B(n_27956), .C(n_54659), .D(n_28417)
		, .Z(n_212178516));
	notech_and4 i_97056948(.A(n_212178516), .B(n_211978514), .C(n_211878513)
		, .D(n_148477884), .Z(n_212378518));
	notech_ao4 i_96256956(.A(n_54685), .B(n_28460), .C(n_58523), .D(n_27269)
		, .Z(n_212478519));
	notech_ao4 i_96056958(.A(n_55792), .B(n_28448), .C(n_54714), .D(n_29386)
		, .Z(n_212678521));
	notech_and4 i_96456954(.A(n_212678521), .B(n_212478519), .C(n_148177881)
		, .D(n_147877878), .Z(n_212878523));
	notech_ao4 i_95756961(.A(n_54771), .B(\nbus_11276[2] ), .C(n_55684), .D(n_55342
		), .Z(n_212978524));
	notech_ao4 i_95656962(.A(n_54659), .B(n_28416), .C(n_54742), .D(n_55299)
		, .Z(n_213078525));
	notech_nand2 i_95856960(.A(n_213078525), .B(n_212978524), .Z(n_213178526
		));
	notech_ao4 i_95356964(.A(n_2234), .B(n_29385), .C(n_54674), .D(n_27955),
		 .Z(n_213278527));
	notech_ao4 i_95056967(.A(n_310288586), .B(n_29384), .C(n_54685), .D(n_28459
		), .Z(n_213578530));
	notech_ao4 i_94856969(.A(n_55792), .B(n_28447), .C(n_54727), .D(nbus_11326
		[2]), .Z(n_213778532));
	notech_or4 i_95256965(.A(n_146577865), .B(n_146877868), .C(n_26430), .D(n_26429
		), .Z(n_213978534));
	notech_nand3 i_94456973(.A(n_146177861), .B(n_146077860), .C(n_146277862
		), .Z(n_214478538));
	notech_ao4 i_94156976(.A(n_2234), .B(n_29383), .C(n_54674), .D(n_27954),
		 .Z(n_214578539));
	notech_ao4 i_93856979(.A(n_310288586), .B(n_29382), .C(n_54685), .D(n_28457
		), .Z(n_214878542));
	notech_ao4 i_93656981(.A(n_55792), .B(n_28446), .C(n_54727), .D(nbus_11326
		[1]), .Z(n_215078544));
	notech_or4 i_94056977(.A(n_145377853), .B(n_145677856), .C(n_26433), .D(n_26432
		), .Z(n_215278546));
	notech_ao3 i_194960625(.A(n_55070), .B(n_54438), .C(n_126074128), .Z(n_215378547
		));
	notech_nand3 i_195260624(.A(n_55071), .B(n_126174129), .C(n_54469), .Z(n_215478548
		));
	notech_or2 i_16855137(.A(n_55534), .B(nbus_11273[24]), .Z(n_216378557)
		);
	notech_or2 i_16555140(.A(n_321388476), .B(n_29137), .Z(n_216678560));
	notech_nand2 i_16255143(.A(sav_ecx[24]), .B(n_60596), .Z(n_216978563));
	notech_nao3 i_22655079(.A(opc_10[10]), .B(n_62431), .C(n_333669135), .Z(n_217678570
		));
	notech_and3 i_128460663(.A(n_55976), .B(n_258664903), .C(n_55974), .Z(n_217778571
		));
	notech_nor2 i_24655059(.A(n_54853), .B(n_29084), .Z(n_217878572));
	notech_ao3 i_24155064(.A(n_62427), .B(opc[12]), .C(n_333569134), .Z(n_218578579
		));
	notech_or2 i_28355022(.A(n_54066), .B(n_26939), .Z(n_219078582));
	notech_or4 i_28055025(.A(n_59159), .B(n_26604), .C(n_26377), .D(n_27527)
		, .Z(n_219378585));
	notech_or2 i_27755028(.A(n_55520), .B(n_29045), .Z(n_219678588));
	notech_or2 i_30954996(.A(n_54066), .B(n_26945), .Z(n_220378595));
	notech_or4 i_30654999(.A(n_59159), .B(n_26604), .C(n_26377), .D(n_27530)
		, .Z(n_220678598));
	notech_or2 i_30355002(.A(n_55520), .B(n_29080), .Z(n_221078601));
	notech_or2 i_33554970(.A(n_54066), .B(n_26949), .Z(n_221778608));
	notech_or4 i_33254973(.A(n_59159), .B(n_26604), .C(n_26377), .D(n_27532)
		, .Z(n_222078611));
	notech_or2 i_32954976(.A(n_55520), .B(n_29037), .Z(n_222378614));
	notech_or2 i_36154944(.A(n_54066), .B(n_26971), .Z(n_223078621));
	notech_or2 i_35854947(.A(n_308518862), .B(nbus_11326[24]), .Z(n_223378624
		));
	notech_or2 i_35554950(.A(n_57334), .B(n_55442), .Z(n_223678627));
	notech_or2 i_36854937(.A(n_57348), .B(n_54872), .Z(n_224178632));
	notech_nor2 i_37654929(.A(n_57347), .B(n_54872), .Z(n_224878639));
	notech_or4 i_37154934(.A(n_322031607), .B(n_55852), .C(n_56158), .D(n_59277
		), .Z(n_225578646));
	notech_nor2 i_38454921(.A(n_57346), .B(n_54872), .Z(n_225678647));
	notech_or4 i_37954926(.A(n_321931606), .B(n_55852), .C(n_56158), .D(n_59277
		), .Z(n_226378654));
	notech_or4 i_40054905(.A(n_57293), .B(n_55852), .C(n_56158), .D(n_59277)
		, .Z(n_226478655));
	notech_or2 i_39554910(.A(n_54943), .B(n_55578), .Z(n_227278662));
	notech_nor2 i_40854897(.A(n_308318860), .B(n_59086), .Z(n_227378663));
	notech_or4 i_40354902(.A(n_56158), .B(n_59277), .C(n_56363), .D(n_27592)
		, .Z(n_228078670));
	notech_nao3 i_49954809(.A(n_3395), .B(\eflags[10] ), .C(n_54707), .Z(n_228378673
		));
	notech_or2 i_49654812(.A(n_271688739), .B(n_56847), .Z(n_228678676));
	notech_or2 i_49354815(.A(n_355688241), .B(n_29137), .Z(n_228978679));
	notech_nand2 i_49054818(.A(sav_esi[24]), .B(n_60596), .Z(n_229278682));
	notech_or4 i_55454755(.A(n_56196), .B(n_56363), .C(n_59250), .D(n_27592)
		, .Z(n_230178691));
	notech_nor2 i_70654617(.A(n_123423221), .B(n_59086), .Z(n_230278692));
	notech_or4 i_70154622(.A(n_56172), .B(n_58656), .C(n_56363), .D(n_27592)
		, .Z(n_230978699));
	notech_nand2 i_91454417(.A(opb[10]), .B(n_215478548), .Z(n_231078700));
	notech_or4 i_90854423(.A(n_56449), .B(n_56431), .C(n_231778707), .D(n_174358031
		), .Z(n_231578705));
	notech_nao3 i_90954422(.A(opc_10[10]), .B(n_62431), .C(n_325776096), .Z(n_231678706
		));
	notech_and4 i_190260636(.A(n_55658), .B(n_135960441), .C(n_55999), .D(n_56005
		), .Z(n_231778707));
	notech_or2 i_113154213(.A(n_55263), .B(n_29087), .Z(n_232078710));
	notech_nand2 i_112854216(.A(n_354069311), .B(opa[15]), .Z(n_232378713)
		);
	notech_nao3 i_112554219(.A(n_205688857), .B(n_6809), .C(n_205588858), .Z
		(n_232678716));
	notech_nand2 i_112254222(.A(\add_len_pc[15] ), .B(n_55819), .Z(n_232978719
		));
	notech_or2 i_114354201(.A(n_2212), .B(n_59086), .Z(n_233278722));
	notech_or2 i_114054204(.A(n_55587), .B(n_57334), .Z(n_233578725));
	notech_nao3 i_113754207(.A(n_6818), .B(n_205688857), .C(n_205588858), .Z
		(n_233878728));
	notech_nand2 i_113454210(.A(\add_len_pc[24] ), .B(n_55819), .Z(n_234178731
		));
	notech_ao4 i_215653207(.A(n_55811), .B(n_322231609), .C(n_2211), .D(n_251061538
		), .Z(n_234278732));
	notech_ao4 i_215453209(.A(n_55842), .B(n_27592), .C(n_59195), .D(n_26790
		), .Z(n_234478734));
	notech_and4 i_215853205(.A(n_234478734), .B(n_234278732), .C(n_233878728
		), .D(n_234178731), .Z(n_234678736));
	notech_ao4 i_215153212(.A(n_55597), .B(n_29137), .C(n_55492), .D(n_27546
		), .Z(n_234778737));
	notech_ao4 i_214953214(.A(n_55567), .B(n_56847), .C(n_55568), .D(n_56207
		), .Z(n_234978739));
	notech_and4 i_215353210(.A(n_234978739), .B(n_234778737), .C(n_233578725
		), .D(n_233278722), .Z(n_235178741));
	notech_ao4 i_214653217(.A(n_354469314), .B(n_177164109), .C(n_354369313)
		, .D(n_177264110), .Z(n_235278742));
	notech_ao4 i_214453219(.A(n_59195), .B(n_26780), .C(n_55693), .D(n_57293
		), .Z(n_235478744));
	notech_and4 i_214853215(.A(n_235478744), .B(n_235278742), .C(n_232678716
		), .D(n_232978719), .Z(n_235678746));
	notech_ao4 i_214153222(.A(n_353969310), .B(n_27581), .C(n_55492), .D(n_27534
		), .Z(n_235778747));
	notech_ao4 i_213953224(.A(n_55264), .B(n_356476400), .C(n_354269312), .D
		(n_55578), .Z(n_235978749));
	notech_and4 i_214353220(.A(n_235978749), .B(n_235778747), .C(n_232078710
		), .D(n_232378713), .Z(n_236178751));
	notech_ao4 i_197953384(.A(n_54433), .B(n_29077), .C(n_319431581), .D(n_55965
		), .Z(n_236478754));
	notech_and3 i_198153382(.A(n_231578705), .B(n_236478754), .C(n_231678706
		), .Z(n_236578755));
	notech_ao4 i_197753386(.A(n_215378547), .B(n_56721), .C(n_57348), .D(n_54445
		), .Z(n_236678756));
	notech_ao4 i_179553563(.A(n_123223219), .B(n_322231609), .C(n_123623223)
		, .D(n_251061538), .Z(n_236978759));
	notech_ao4 i_179453564(.A(n_2702), .B(n_57334), .C(n_29137), .D(n_26450)
		, .Z(n_237178761));
	notech_nand3 i_179753561(.A(n_230978699), .B(n_236978759), .C(n_237178761
		), .Z(n_237278762));
	notech_ao4 i_179253566(.A(n_55073), .B(n_56847), .C(n_55072), .D(n_56207
		), .Z(n_237378763));
	notech_ao4 i_168053678(.A(n_322231609), .B(n_354569315), .C(n_113113525)
		, .D(n_251061538), .Z(n_237678766));
	notech_ao4 i_167953679(.A(n_29137), .B(n_26571), .C(n_2193), .D(n_27546)
		, .Z(n_237878768));
	notech_and3 i_168253676(.A(n_237678766), .B(n_237878768), .C(n_230178691
		), .Z(n_237978769));
	notech_ao4 i_167753681(.A(n_354669316), .B(n_56207), .C(n_57334), .D(n_354969318
		), .Z(n_238078770));
	notech_ao4 i_167653682(.A(n_113313527), .B(n_59086), .C(n_55562), .D(n_56847
		), .Z(n_238178771));
	notech_ao4 i_163253726(.A(n_322231609), .B(n_355788240), .C(n_353788271)
		, .D(n_251061538), .Z(n_238378773));
	notech_ao4 i_163053728(.A(n_27546), .B(n_59159), .C(n_320088489), .D(n_27592
		), .Z(n_238578775));
	notech_and4 i_163453724(.A(n_238578775), .B(n_238378773), .C(n_228978679
		), .D(n_229278682), .Z(n_238778777));
	notech_ao4 i_162753731(.A(n_271588740), .B(n_56207), .C(n_57334), .D(n_355488242
		), .Z(n_238878778));
	notech_ao4 i_162553733(.A(n_54024), .B(n_29421), .C(n_55133), .D(n_59086
		), .Z(n_239078780));
	notech_and4 i_162953729(.A(n_239078780), .B(n_238878778), .C(n_228378673
		), .D(n_228678676), .Z(n_239278782));
	notech_ao4 i_156053798(.A(n_322231609), .B(n_309518872), .C(n_251061538)
		, .D(n_308718864), .Z(n_239378783));
	notech_ao4 i_155953799(.A(n_55554), .B(n_57334), .C(n_55555), .D(n_29137
		), .Z(n_239578785));
	notech_nand3 i_156253796(.A(n_239378783), .B(n_239578785), .C(n_228078670
		), .Z(n_239678786));
	notech_ao4 i_155753801(.A(n_55219), .B(n_56847), .C(n_55218), .D(n_56207
		), .Z(n_239778787));
	notech_ao4 i_155353805(.A(n_177164109), .B(n_318231569), .C(n_177264110)
		, .D(n_318031567), .Z(n_240078790));
	notech_ao4 i_155253806(.A(n_55726), .B(n_27581), .C(n_54944), .D(n_56766
		), .Z(n_240278792));
	notech_and3 i_155553803(.A(n_240078790), .B(n_240278792), .C(n_227278662
		), .Z(n_240378793));
	notech_ao4 i_155053808(.A(n_356476400), .B(n_54872), .C(n_54902), .D(n_29087
		), .Z(n_240478794));
	notech_ao4 i_153853819(.A(n_169157979), .B(n_318231569), .C(n_169057978)
		, .D(n_318031567), .Z(n_240778797));
	notech_ao4 i_153753820(.A(n_56739), .B(n_54944), .C(n_54943), .D(n_55542
		), .Z(n_240978799));
	notech_nand3 i_154053817(.A(n_226378654), .B(n_240778797), .C(n_240978799
		), .Z(n_241078800));
	notech_ao4 i_153553822(.A(n_54902), .B(n_29084), .C(n_55726), .D(n_27577
		), .Z(n_241178801));
	notech_ao4 i_153153826(.A(n_171758005), .B(n_318231569), .C(n_171658004)
		, .D(n_318031567), .Z(n_241478804));
	notech_ao4 i_153053827(.A(n_54944), .B(n_56730), .C(n_54943), .D(n_55469
		), .Z(n_241678806));
	notech_nand3 i_153353824(.A(n_225578646), .B(n_241478804), .C(n_241678806
		), .Z(n_241778807));
	notech_ao4 i_152853829(.A(n_54902), .B(n_29080), .C(n_55726), .D(n_27576
		), .Z(n_241878808));
	notech_ao4 i_152553832(.A(n_174358031), .B(n_318231569), .C(n_174258030)
		, .D(n_318031567), .Z(n_242178811));
	notech_ao4 i_152453833(.A(n_54943), .B(n_55438), .C(n_319431581), .D(n_55906
		), .Z(n_242278812));
	notech_ao4 i_152253835(.A(n_54902), .B(n_29077), .C(n_54944), .D(n_56721
		), .Z(n_242478814));
	notech_and3 i_152353834(.A(n_154070859), .B(n_242478814), .C(n_224178632
		), .Z(n_242678816));
	notech_ao4 i_151853839(.A(n_322231609), .B(n_55780), .C(n_251061538), .D
		(n_308618863), .Z(n_242778817));
	notech_ao4 i_151753840(.A(n_55135), .B(n_27592), .C(n_59195), .D(n_26709
		), .Z(n_242878818));
	notech_ao4 i_151553842(.A(n_55443), .B(n_29137), .C(n_262536780), .D(n_27546
		), .Z(n_243078820));
	notech_and4 i_152053837(.A(n_243078820), .B(n_242878818), .C(n_242778817
		), .D(n_223678627), .Z(n_243278822));
	notech_ao4 i_151253845(.A(n_55536), .B(n_56847), .C(n_55535), .D(n_56207
		), .Z(n_243378823));
	notech_ao4 i_151053847(.A(n_54080), .B(n_28438), .C(n_54092), .D(n_29420
		), .Z(n_243578825));
	notech_and4 i_151453843(.A(n_243578825), .B(n_243378823), .C(n_223078621
		), .D(n_223378624), .Z(n_243778827));
	notech_ao4 i_149653861(.A(n_166557953), .B(n_320565522), .C(n_166457952)
		, .D(n_320665523), .Z(n_243878828));
	notech_ao4 i_149553862(.A(n_55381), .B(n_55552), .C(n_321831605), .D(n_320465521
		), .Z(n_243978829));
	notech_ao4 i_149353864(.A(n_55519), .B(n_57345), .C(n_55382), .D(n_56748
		), .Z(n_244178831));
	notech_and4 i_149853859(.A(n_244178831), .B(n_243978829), .C(n_243878828
		), .D(n_222378614), .Z(n_244378833));
	notech_ao4 i_149053867(.A(n_59176), .B(n_26699), .C(n_55738), .D(n_27578
		), .Z(n_244478834));
	notech_ao4 i_148853869(.A(n_54080), .B(n_28427), .C(n_54092), .D(n_29419
		), .Z(n_244678836));
	notech_and4 i_149253865(.A(n_244678836), .B(n_244478834), .C(n_221778608
		), .D(n_222078611), .Z(n_244878838));
	notech_ao4 i_147253883(.A(n_171758005), .B(n_320565522), .C(n_171658004)
		, .D(n_320665523), .Z(n_244978839));
	notech_ao4 i_147153884(.A(n_55381), .B(n_55469), .C(n_320465521), .D(n_322031607
		), .Z(n_245078840));
	notech_ao4 i_146953886(.A(n_55519), .B(n_57347), .C(n_55382), .D(n_56730
		), .Z(n_245278842));
	notech_and4 i_147453881(.A(n_245278842), .B(n_245078840), .C(n_244978839
		), .D(n_221078601), .Z(n_245478844));
	notech_ao4 i_146653889(.A(n_59176), .B(n_26696), .C(n_55738), .D(n_27576
		), .Z(n_245578845));
	notech_ao4 i_146453891(.A(n_54080), .B(n_28425), .C(n_54092), .D(n_29418
		), .Z(n_245778847));
	notech_and4 i_146853887(.A(n_245778847), .B(n_245578845), .C(n_220378595
		), .D(n_220678598), .Z(n_245978849));
	notech_ao4 i_145053905(.A(n_161857906), .B(n_320565522), .C(n_161957907)
		, .D(n_320665523), .Z(n_246078850));
	notech_ao4 i_144953906(.A(n_55381), .B(n_55413), .C(n_57300), .D(n_320465521
		), .Z(n_246178851));
	notech_ao4 i_144653908(.A(n_57350), .B(n_55519), .C(n_55382), .D(n_56703
		), .Z(n_246378853));
	notech_and4 i_145253903(.A(n_246378853), .B(n_246178851), .C(n_246078850
		), .D(n_219678588), .Z(n_246578855));
	notech_ao4 i_144353911(.A(n_59176), .B(n_26693), .C(n_27571), .D(n_55738
		), .Z(n_246678856));
	notech_ao4 i_144153913(.A(n_54080), .B(n_28422), .C(n_54092), .D(n_29417
		), .Z(n_246878858));
	notech_and4 i_144553909(.A(n_246878858), .B(n_246678856), .C(n_219078582
		), .D(n_219378585), .Z(n_247078860));
	notech_ao4 i_140953939(.A(n_169057978), .B(n_333669135), .C(n_189074758)
		, .D(n_55888), .Z(n_247178861));
	notech_ao4 i_140853940(.A(n_54946), .B(n_56739), .C(n_55725), .D(n_27577
		), .Z(n_247378863));
	notech_nao3 i_141153937(.A(n_247178861), .B(n_247378863), .C(n_218578579
		), .Z(n_247478864));
	notech_ao4 i_140653942(.A(n_57346), .B(n_54852), .C(n_54945), .D(n_55542
		), .Z(n_247578865));
	notech_nao3 i_139753951(.A(n_56487), .B(n_268064997), .C(n_217778571), .Z
		(n_247878868));
	notech_ao4 i_139453954(.A(n_319431581), .B(n_55888), .C(n_174358031), .D
		(n_247878868), .Z(n_247978869));
	notech_ao4 i_139353955(.A(n_54945), .B(n_55438), .C(n_54946), .D(n_56721
		), .Z(n_248178871));
	notech_and3 i_139653952(.A(n_247978869), .B(n_248178871), .C(n_217678570
		), .Z(n_248278872));
	notech_ao4 i_139153957(.A(n_54853), .B(n_29077), .C(n_57348), .D(n_54852
		), .Z(n_248378873));
	notech_ao4 i_133554013(.A(n_322231609), .B(n_3214), .C(n_251061538), .D(n_321588475
		), .Z(n_248678876));
	notech_ao4 i_133354015(.A(n_170914103), .B(n_27546), .C(n_131423301), .D
		(n_27592), .Z(n_248878878));
	notech_and4 i_133754011(.A(n_248878878), .B(n_248678876), .C(n_216678560
		), .D(n_216978563), .Z(n_249078880));
	notech_ao4 i_133054018(.A(n_55533), .B(n_56207), .C(n_57334), .D(n_321288477
		), .Z(n_249178881));
	notech_ao4 i_132954019(.A(n_55131), .B(n_29416), .C(n_131123298), .D(n_59086
		), .Z(n_249378883));
	notech_or4 i_125550781(.A(n_2688), .B(n_55827), .C(n_56163), .D(n_59277)
		, .Z(n_249578885));
	notech_or2 i_125250784(.A(n_55730), .B(n_55342), .Z(n_250078890));
	notech_nao3 i_125350783(.A(n_62423), .B(opc[0]), .C(n_248734113), .Z(n_250178891
		));
	notech_or4 i_125450782(.A(n_55975), .B(n_28051), .C(n_60504), .D(n_294261946
		), .Z(n_250278892));
	notech_and4 i_121580(.A(n_41726130), .B(n_250778897), .C(n_249578885), .D
		(n_250278892), .Z(n_13115));
	notech_ao4 i_125750779(.A(n_54920), .B(n_55356), .C(n_54921), .D(nbus_11273
		[0]), .Z(n_250378893));
	notech_ao4 i_125650780(.A(n_54748), .B(n_28986), .C(n_2699), .D(n_54740)
		, .Z(n_250478894));
	notech_and4 i_126050776(.A(n_250478894), .B(n_250378893), .C(n_250078890
		), .D(n_250178891), .Z(n_250778897));
	notech_or2 i_49448690(.A(n_55068), .B(n_56901), .Z(n_251478904));
	notech_nao3 i_49748687(.A(opc_10[30]), .B(n_62415), .C(n_2694), .Z(n_251578905
		));
	notech_or4 i_49648688(.A(n_56172), .B(n_56163), .C(n_55794), .D(n_271188744
		), .Z(n_251678906));
	notech_or2 i_49548689(.A(n_2655), .B(n_270988746), .Z(n_251778907));
	notech_and4 i_3120746(.A(n_256478954), .B(n_101523002), .C(n_251678906),
		 .D(n_251778907), .Z(n_19617));
	notech_or2 i_121248017(.A(n_2320), .B(n_271088745), .Z(n_251878908));
	notech_and3 i_120148028(.A(n_2219), .B(resb_shift4box[31]), .C(n_274788710
		), .Z(n_251978909));
	notech_and4 i_3216201(.A(n_256878958), .B(n_256778957), .C(n_257678966),
		 .D(n_251878908), .Z(n_14278));
	notech_and2 i_179947456(.A(opc[4]), .B(n_253178921), .Z(n_253078920));
	notech_or4 i_2249136(.A(opc[3]), .B(opc[2]), .C(opc[0]), .D(opc[1]), .Z(n_253178921
		));
	notech_or2 i_180547450(.A(n_271488741), .B(n_253778927), .Z(n_253678926)
		);
	notech_xor2 i_2049138(.A(opc[4]), .B(n_257878968), .Z(n_253778927));
	notech_ao4 i_180447451(.A(n_253078920), .B(n_270388750), .C(n_26445), .D
		(n_26553), .Z(n_254078930));
	notech_ao3 i_1949139(.A(n_257978969), .B(n_253678926), .C(n_254078930), 
		.Z(n_254378933));
	notech_xor2 i_1849140(.A(n_55541), .B(opc[4]), .Z(n_254578935));
	notech_ao3 i_182147434(.A(n_26712), .B(n_57445), .C(n_254778937), .Z(n_254678936
		));
	notech_ao4 i_1749141(.A(n_275988698), .B(n_254578935), .C(n_276088697), 
		.D(n_254378933), .Z(n_254778937));
	notech_or2 i_181147444(.A(n_54735), .B(n_55542), .Z(n_254878938));
	notech_or4 i_182047435(.A(n_60780), .B(n_60729), .C(n_55365), .D(n_54998
		), .Z(n_255778947));
	notech_or4 i_182247433(.A(n_56117), .B(n_58904), .C(n_59931), .D(n_57326
		), .Z(n_255878948));
	notech_and4 i_182347432(.A(read_data[20]), .B(n_59931), .C(n_26712), .D(n_26611
		), .Z(n_255978949));
	notech_or4 i_516814(.A(n_255978949), .B(n_254678936), .C(n_26447), .D(n_26446
		), .Z(n_9727));
	notech_ao4 i_49948685(.A(n_55717), .B(n_27599), .C(n_28997), .D(n_26444)
		, .Z(n_256078950));
	notech_ao4 i_49848686(.A(n_55069), .B(n_55234), .C(n_2672), .D(n_59050),
		 .Z(n_256178951));
	notech_and4 i_50248682(.A(n_256178951), .B(n_256078950), .C(n_251478904)
		, .D(n_251578905), .Z(n_256478954));
	notech_ao4 i_121748012(.A(n_2323), .B(n_27601), .C(n_55243), .D(n_27554)
		, .Z(n_256778957));
	notech_ao4 i_121848011(.A(n_2319), .B(n_29029), .C(n_2322), .D(n_58951),
		 .Z(n_256878958));
	notech_ao4 i_121448015(.A(n_55526), .B(n_28595), .C(n_55366), .D(n_28800
		), .Z(n_257178961));
	notech_ao3 i_121948010(.A(n_2187), .B(n_257178961), .C(n_251978909), .Z(n_257278962
		));
	notech_ao4 i_121548014(.A(n_2318), .B(n_28855), .C(n_55619), .D(n_28642)
		, .Z(n_257378963));
	notech_ao4 i_121648013(.A(n_55933), .B(n_56943), .C(n_2164), .D(n_59095)
		, .Z(n_257478964));
	notech_and3 i_122248007(.A(n_257478964), .B(n_257378963), .C(n_257278962
		), .Z(n_257678966));
	notech_or4 i_2549134(.A(nbus_11326[1]), .B(nbus_11326[0]), .C(nbus_11326
		[2]), .D(nbus_11326[3]), .Z(n_257878968));
	notech_ao4 i_180647449(.A(n_271388742), .B(n_29423), .C(n_26889), .D(n_29422
		), .Z(n_257978969));
	notech_ao4 i_182847427(.A(n_231547139), .B(nbus_11326[28]), .C(n_55009),
		 .D(n_28055), .Z(n_258178971));
	notech_ao4 i_182947426(.A(n_2247), .B(n_29424), .C(n_2313), .D(n_28905),
		 .Z(n_258278972));
	notech_ao4 i_183047425(.A(n_329546800), .B(n_29425), .C(n_2248), .D(nbus_11348
		[4]), .Z(n_258478974));
	notech_and4 i_183547420(.A(n_258478974), .B(n_258278972), .C(n_258178971
		), .D(n_255778947), .Z(n_258678976));
	notech_ao4 i_182747428(.A(n_54884), .B(nbus_11326[4]), .C(n_2311), .D(n_29327
		), .Z(n_259078980));
	notech_and4 i_183447421(.A(n_2186), .B(n_259078980), .C(n_255878948), .D
		(n_254878938), .Z(n_259278982));
	notech_or2 i_11445263(.A(n_55534), .B(n_56838), .Z(n_259978989));
	notech_or4 i_11145266(.A(n_60596), .B(n_59789), .C(n_26629), .D(n_27545)
		, .Z(n_260278992));
	notech_or2 i_10845269(.A(n_308921976), .B(n_321288477), .Z(n_260578995)
		);
	notech_nor2 i_28445094(.A(n_55557), .B(n_29152), .Z(n_260678996));
	notech_or4 i_27945099(.A(n_56074), .B(n_59277), .C(n_55523), .D(n_308521972
		), .Z(n_261379003));
	notech_or2 i_34645034(.A(n_54066), .B(n_26969), .Z(n_261679006));
	notech_or2 i_34345037(.A(n_308518862), .B(nbus_11326[23]), .Z(n_261979009
		));
	notech_or2 i_34045040(.A(n_55443), .B(n_29152), .Z(n_262279012));
	notech_or2 i_35945021(.A(n_54066), .B(n_26973), .Z(n_262979019));
	notech_or2 i_35645024(.A(n_308518862), .B(nbus_11326[25]), .Z(n_263279022
		));
	notech_or2 i_35345027(.A(n_354688262), .B(n_29215), .Z(n_263579025));
	notech_or2 i_37245008(.A(n_54066), .B(n_26975), .Z(n_264279032));
	notech_or2 i_36945011(.A(n_308518862), .B(n_59068), .Z(n_264579035));
	notech_or2 i_36645014(.A(n_354688262), .B(n_29156), .Z(n_264879038));
	notech_or2 i_38844995(.A(n_54066), .B(n_26977), .Z(n_265579045));
	notech_or2 i_38544998(.A(n_308518862), .B(n_59059), .Z(n_265879048));
	notech_or2 i_38245001(.A(n_354688262), .B(n_29154), .Z(n_266179051));
	notech_or2 i_40144982(.A(n_54066), .B(n_26979), .Z(n_266879058));
	notech_or4 i_39844985(.A(n_56363), .B(n_55992), .C(n_60596), .D(n_27596)
		, .Z(n_267179061));
	notech_or2 i_39544988(.A(n_57306), .B(n_110123088), .Z(n_267479064));
	notech_nor2 i_40944974(.A(n_308318860), .B(nbus_11326[23]), .Z(n_267979069
		));
	notech_or2 i_40444979(.A(n_308921976), .B(n_55554), .Z(n_268679076));
	notech_nao3 i_45644934(.A(n_3393), .B(\eflags[10] ), .C(n_54046), .Z(n_268979079
		));
	notech_or2 i_45244937(.A(n_271688739), .B(n_56838), .Z(n_269279082));
	notech_nand3 i_44944940(.A(n_59176), .B(n_59936), .C(read_data[23]), .Z(n_269579085
		));
	notech_or2 i_44644943(.A(n_308921976), .B(n_355488242), .Z(n_269879088)
		);
	notech_nao3 i_46844922(.A(n_3397), .B(\eflags[10] ), .C(n_54046), .Z(n_270179091
		));
	notech_or2 i_46544925(.A(n_271688739), .B(n_56856), .Z(n_270479094));
	notech_or4 i_46244928(.A(n_56363), .B(n_56097), .C(n_60596), .D(n_27593)
		, .Z(n_270779097));
	notech_or2 i_45944931(.A(n_308821975), .B(n_55313), .Z(n_271079100));
	notech_nao3 i_48044910(.A(n_3399), .B(\eflags[10] ), .C(n_54046), .Z(n_271379103
		));
	notech_or2 i_47744913(.A(n_271688739), .B(n_56865), .Z(n_271679106));
	notech_or4 i_47444916(.A(n_56369), .B(n_56097), .C(n_60579), .D(n_27594)
		, .Z(n_271979109));
	notech_or2 i_47144919(.A(n_308721974), .B(n_55313), .Z(n_272279112));
	notech_nao3 i_49244898(.A(n_3401), .B(\eflags[10] ), .C(n_54046), .Z(n_272579115
		));
	notech_or2 i_48944901(.A(n_271688739), .B(n_56874), .Z(n_272879118));
	notech_or4 i_48644904(.A(n_56369), .B(n_56092), .C(n_60579), .D(n_27595)
		, .Z(n_273179121));
	notech_or2 i_48344907(.A(n_308621973), .B(n_55313), .Z(n_273479124));
	notech_nao3 i_50444886(.A(n_3403), .B(\eflags[10] ), .C(n_54046), .Z(n_273779127
		));
	notech_or2 i_50144889(.A(n_55133), .B(nbus_11326[28]), .Z(n_274079130)
		);
	notech_nand3 i_49844892(.A(n_59176), .B(n_59936), .C(read_data[28]), .Z(n_274379133
		));
	notech_or2 i_49544895(.A(n_55314), .B(n_29219), .Z(n_274679136));
	notech_or2 i_50744883(.A(n_308921976), .B(n_354969318), .Z(n_275579145)
		);
	notech_ao4 i_158143847(.A(n_308521972), .B(n_354569315), .C(n_270765024)
		, .D(n_113113525), .Z(n_275679146));
	notech_ao4 i_158043848(.A(n_2193), .B(n_27545), .C(n_27590), .D(n_55776)
		, .Z(n_275879148));
	notech_and3 i_158343845(.A(n_275679146), .B(n_275879148), .C(n_275579145
		), .Z(n_275979149));
	notech_ao4 i_157743850(.A(n_354669316), .B(n_59319), .C(n_29152), .D(n_26571
		), .Z(n_276079150));
	notech_ao4 i_157643851(.A(n_113313527), .B(nbus_11326[23]), .C(n_55562),
		 .D(n_56838), .Z(n_276179151));
	notech_ao4 i_157343854(.A(n_57306), .B(n_302821915), .C(n_343565725), .D
		(n_302321910), .Z(n_276379153));
	notech_ao4 i_157143856(.A(n_59176), .B(n_26738), .C(n_57330), .D(n_55313
		), .Z(n_276579155));
	notech_and4 i_157543852(.A(n_276579155), .B(n_276379153), .C(n_274379133
		), .D(n_274679136), .Z(n_276779157));
	notech_ao4 i_156843859(.A(n_271688739), .B(n_56883), .C(n_271588740), .D
		(n_55261), .Z(n_276879158));
	notech_ao4 i_156643861(.A(n_54024), .B(n_29436), .C(n_320088489), .D(n_27596
		), .Z(n_277079160));
	notech_and4 i_157043857(.A(n_277079160), .B(n_276879158), .C(n_273779127
		), .D(n_274079130), .Z(n_277279162));
	notech_ao4 i_156343864(.A(n_308221969), .B(n_302821915), .C(n_286061878)
		, .D(n_302321910), .Z(n_277379163));
	notech_ao4 i_156143866(.A(n_59174), .B(n_26737), .C(n_55314), .D(n_29154
		), .Z(n_277579165));
	notech_and4 i_156543862(.A(n_277579165), .B(n_277379163), .C(n_273479124
		), .D(n_273179121), .Z(n_277779167));
	notech_ao4 i_155743869(.A(n_271588740), .B(n_59328), .C(n_59159), .D(n_27550
		), .Z(n_277879168));
	notech_ao4 i_155543871(.A(n_54024), .B(n_29435), .C(n_55133), .D(n_59059
		), .Z(n_278079170));
	notech_and4 i_156043867(.A(n_278079170), .B(n_277879168), .C(n_272579115
		), .D(n_272879118), .Z(n_278279172));
	notech_ao4 i_155243874(.A(n_302821915), .B(n_308321970), .C(n_288561889)
		, .D(n_302321910), .Z(n_278379173));
	notech_ao4 i_155043876(.A(n_59174), .B(n_26735), .C(n_55314), .D(n_29156
		), .Z(n_278579175));
	notech_and4 i_155443872(.A(n_278579175), .B(n_278379173), .C(n_272279112
		), .D(n_271979109), .Z(n_278779177));
	notech_ao4 i_154743879(.A(n_271588740), .B(n_59337), .C(n_59159), .D(n_27549
		), .Z(n_278879178));
	notech_ao4 i_154543881(.A(n_54024), .B(n_29434), .C(n_55133), .D(n_59068
		), .Z(n_279079180));
	notech_and4 i_154943877(.A(n_279079180), .B(n_278879178), .C(n_271379103
		), .D(n_271679106), .Z(n_279279182));
	notech_ao4 i_154243884(.A(n_308421971), .B(n_302821915), .C(n_268264999)
		, .D(n_302321910), .Z(n_279379183));
	notech_ao4 i_154043886(.A(n_59174), .B(n_26734), .C(n_55314), .D(n_29215
		), .Z(n_279579185));
	notech_and4 i_154443882(.A(n_279579185), .B(n_279379183), .C(n_271079100
		), .D(n_270779097), .Z(n_279779187));
	notech_ao4 i_153743889(.A(n_271588740), .B(n_59346), .C(n_59159), .D(n_27548
		), .Z(n_279879188));
	notech_ao4 i_153543891(.A(n_54024), .B(n_29433), .C(n_55133), .D(nbus_11326
		[25]), .Z(n_280079190));
	notech_and4 i_153943887(.A(n_280079190), .B(n_279879188), .C(n_270179091
		), .D(n_270479094), .Z(n_280279192));
	notech_ao4 i_153243894(.A(n_308521972), .B(n_355788240), .C(n_270765024)
		, .D(n_353788271), .Z(n_280379193));
	notech_ao4 i_152943896(.A(n_320088489), .B(n_27590), .C(n_59174), .D(n_26733
		), .Z(n_280579195));
	notech_and4 i_153443892(.A(n_280579195), .B(n_280379193), .C(n_269579085
		), .D(n_269879088), .Z(n_280779197));
	notech_ao4 i_152643899(.A(n_271588740), .B(n_59319), .C(n_355688241), .D
		(n_29152), .Z(n_280879198));
	notech_ao4 i_152443901(.A(n_54024), .B(n_29432), .C(n_55133), .D(n_59041
		), .Z(n_281079200));
	notech_and4 i_152843897(.A(n_281079200), .B(n_280879198), .C(n_268979079
		), .D(n_269279082), .Z(n_281279202));
	notech_ao4 i_149743928(.A(n_308521972), .B(n_309518872), .C(n_270765024)
		, .D(n_308718864), .Z(n_281379203));
	notech_ao4 i_149643929(.A(n_55555), .B(n_29152), .C(n_55773), .D(n_27590
		), .Z(n_281579205));
	notech_nand3 i_149943926(.A(n_281379203), .B(n_281579205), .C(n_268679076
		), .Z(n_281679206));
	notech_ao4 i_149443931(.A(n_56838), .B(n_55219), .C(n_55218), .D(n_59319
		), .Z(n_281779207));
	notech_ao4 i_149043935(.A(n_59174), .B(n_26715), .C(n_57330), .D(n_354588263
		), .Z(n_282079210));
	notech_ao4 i_148943936(.A(n_55535), .B(n_55261), .C(n_262536780), .D(n_27551
		), .Z(n_282179211));
	notech_ao4 i_148643938(.A(n_354688262), .B(n_29219), .C(n_55536), .D(n_56883
		), .Z(n_282379213));
	notech_and4 i_149243933(.A(n_282379213), .B(n_282179211), .C(n_282079210
		), .D(n_267479064), .Z(n_282579215));
	notech_ao4 i_148343941(.A(n_308518862), .B(n_59077), .C(n_343565725), .D
		(n_110323090), .Z(n_282679216));
	notech_ao4 i_148143943(.A(n_54080), .B(n_28442), .C(n_54092), .D(n_29431
		), .Z(n_282879218));
	notech_and4 i_148543939(.A(n_282879218), .B(n_282679216), .C(n_266879058
		), .D(n_267179061), .Z(n_283079220));
	notech_ao4 i_147843946(.A(n_308221969), .B(n_110123088), .C(n_286061878)
		, .D(n_110323090), .Z(n_283179221));
	notech_ao4 i_147743947(.A(n_59174), .B(n_26713), .C(n_308621973), .D(n_354588263
		), .Z(n_283279222));
	notech_ao4 i_147543949(.A(n_262536780), .B(n_27550), .C(n_55135), .D(n_27595
		), .Z(n_283479224));
	notech_and4 i_148043944(.A(n_283479224), .B(n_283279222), .C(n_283179221
		), .D(n_266179051), .Z(n_283679226));
	notech_ao4 i_147243952(.A(n_55536), .B(n_56874), .C(n_55535), .D(n_59328
		), .Z(n_283779227));
	notech_ao4 i_147043954(.A(n_54080), .B(n_28441), .C(n_54092), .D(n_29430
		), .Z(n_283979229));
	notech_and4 i_147443950(.A(n_283979229), .B(n_283779227), .C(n_265579045
		), .D(n_265879048), .Z(n_284179231));
	notech_ao4 i_146743957(.A(n_308321970), .B(n_110123088), .C(n_288561889)
		, .D(n_110323090), .Z(n_284279232));
	notech_ao4 i_146643958(.A(n_59176), .B(n_26711), .C(n_308721974), .D(n_354588263
		), .Z(n_284379233));
	notech_ao4 i_146443960(.A(n_262536780), .B(n_27549), .C(n_55135), .D(n_27594
		), .Z(n_284579235));
	notech_and4 i_146943955(.A(n_284579235), .B(n_284379233), .C(n_284279232
		), .D(n_264879038), .Z(n_284779237));
	notech_ao4 i_146143963(.A(n_55536), .B(n_56865), .C(n_55535), .D(n_59337
		), .Z(n_284879238));
	notech_ao4 i_145943965(.A(n_54080), .B(n_28440), .C(n_54092), .D(n_29429
		), .Z(n_285079240));
	notech_and4 i_146343961(.A(n_285079240), .B(n_284879238), .C(n_264279032
		), .D(n_264579035), .Z(n_285279242));
	notech_ao4 i_145643968(.A(n_308421971), .B(n_110123088), .C(n_268264999)
		, .D(n_110323090), .Z(n_285379243));
	notech_ao4 i_145543969(.A(n_59176), .B(n_26710), .C(n_308821975), .D(n_354588263
		), .Z(n_285479244));
	notech_ao4 i_145343971(.A(n_262536780), .B(n_27548), .C(n_55135), .D(n_27593
		), .Z(n_285679246));
	notech_and4 i_145843966(.A(n_285679246), .B(n_285479244), .C(n_285379243
		), .D(n_263579025), .Z(n_285879248));
	notech_ao4 i_144743974(.A(n_55536), .B(n_56856), .C(n_55535), .D(n_59346
		), .Z(n_285979249));
	notech_ao4 i_144443976(.A(n_54080), .B(n_28439), .C(n_54092), .D(n_29428
		), .Z(n_286179251));
	notech_and4 i_145243972(.A(n_286179251), .B(n_285979249), .C(n_262979019
		), .D(n_263279022), .Z(n_286379253));
	notech_ao4 i_144143979(.A(n_308521972), .B(n_55780), .C(n_270765024), .D
		(n_308618863), .Z(n_286479254));
	notech_ao4 i_144043980(.A(n_59176), .B(n_26708), .C(n_308921976), .D(n_55442
		), .Z(n_286579255));
	notech_ao4 i_143843982(.A(n_262536780), .B(n_27545), .C(n_55135), .D(n_27590
		), .Z(n_286779257));
	notech_and4 i_144343977(.A(n_286779257), .B(n_286579255), .C(n_286479254
		), .D(n_262279012), .Z(n_286979259));
	notech_ao4 i_143543985(.A(n_55536), .B(n_56838), .C(n_55535), .D(n_59319
		), .Z(n_287079260));
	notech_ao4 i_143343987(.A(n_54080), .B(n_28437), .C(n_56024), .D(n_29427
		), .Z(n_287279262));
	notech_and4 i_143743983(.A(n_287279262), .B(n_287079260), .C(n_261679006
		), .D(n_261979009), .Z(n_287479264));
	notech_ao4 i_134244078(.A(n_322931616), .B(n_270765024), .C(n_303421921)
		, .D(n_59041), .Z(n_287579265));
	notech_ao4 i_134144079(.A(n_55220), .B(n_56838), .C(n_55556), .D(n_308921976
		), .Z(n_287779267));
	notech_nand3 i_134444076(.A(n_287579265), .B(n_287779267), .C(n_261379003
		), .Z(n_287879268));
	notech_ao4 i_133944081(.A(n_55772), .B(n_27590), .C(n_55221), .D(n_59319
		), .Z(n_287979269));
	notech_ao4 i_119144227(.A(n_308521972), .B(n_3214), .C(n_270765024), .D(n_321588475
		), .Z(n_288279272));
	notech_ao4 i_118944229(.A(n_131423301), .B(n_27590), .C(n_59176), .D(n_26658
		), .Z(n_288479274));
	notech_and4 i_119344225(.A(n_288479274), .B(n_288279272), .C(n_260278992
		), .D(n_260578995), .Z(n_288679276));
	notech_ao4 i_118644232(.A(n_55533), .B(n_59319), .C(n_321388476), .D(n_29152
		), .Z(n_288779277));
	notech_ao4 i_118544233(.A(n_55131), .B(n_29426), .C(n_131123298), .D(n_59041
		), .Z(n_288979279));
	notech_or2 i_8542157(.A(n_55534), .B(nbus_11273[19]), .Z(n_289579285));
	notech_or4 i_8242160(.A(n_60579), .B(n_59809), .C(n_59771), .D(n_27539),
		 .Z(n_289879288));
	notech_or2 i_7942163(.A(n_311218889), .B(n_321288477), .Z(n_290179291)
		);
	notech_or2 i_9642146(.A(n_55534), .B(nbus_11273[20]), .Z(n_290679296));
	notech_or4 i_9342149(.A(n_60579), .B(n_59809), .C(n_59771), .D(n_27540),
		 .Z(n_290979299));
	notech_or2 i_9042152(.A(n_311118888), .B(n_321288477), .Z(n_291279302)
		);
	notech_or2 i_10742135(.A(n_55534), .B(nbus_11273[21]), .Z(n_291779307)
		);
	notech_or4 i_10442138(.A(n_60579), .B(n_59809), .C(n_59771), .D(n_27541)
		, .Z(n_292079310));
	notech_or2 i_10142141(.A(n_311018887), .B(n_321288477), .Z(n_292379313)
		);
	notech_or2 i_11842124(.A(n_55534), .B(n_56829), .Z(n_292879318));
	notech_or4 i_11542127(.A(n_60579), .B(n_59809), .C(n_59771), .D(n_27542)
		, .Z(n_293179321));
	notech_or2 i_11242130(.A(n_26618), .B(n_321288477), .Z(n_293479324));
	notech_or2 i_23342009(.A(n_303421921), .B(nbus_11326[18]), .Z(n_293779327
		));
	notech_or2 i_22842014(.A(n_311318890), .B(n_55556), .Z(n_294279332));
	notech_or2 i_24242001(.A(n_303421921), .B(nbus_11326[19]), .Z(n_294579335
		));
	notech_or2 i_23642006(.A(n_311218889), .B(n_55556), .Z(n_295079340));
	notech_nor2 i_25041993(.A(n_303421921), .B(nbus_11326[20]), .Z(n_295179341
		));
	notech_or2 i_24541998(.A(n_311118888), .B(n_55556), .Z(n_295879348));
	notech_or2 i_25841985(.A(n_303421921), .B(nbus_11326[21]), .Z(n_296179351
		));
	notech_or2 i_25341990(.A(n_311018887), .B(n_55556), .Z(n_296679356));
	notech_or2 i_27941964(.A(n_54066), .B(n_26959), .Z(n_296979359));
	notech_or4 i_27641967(.A(n_59159), .B(n_26604), .C(n_26377), .D(n_27538)
		, .Z(n_297279362));
	notech_or2 i_27341970(.A(n_55536), .B(nbus_11273[18]), .Z(n_297579365)
		);
	notech_or2 i_29241951(.A(n_54066), .B(n_26961), .Z(n_298279372));
	notech_or4 i_28941954(.A(n_59159), .B(n_26604), .C(n_26377), .D(n_27539)
		, .Z(n_298579375));
	notech_or2 i_28641957(.A(n_55536), .B(n_56802), .Z(n_298879378));
	notech_or2 i_30541938(.A(n_54066), .B(n_26963), .Z(n_299579385));
	notech_or4 i_30241941(.A(n_59159), .B(n_26604), .C(n_26377), .D(n_27540)
		, .Z(n_299879388));
	notech_or2 i_29941944(.A(n_55536), .B(nbus_11273[20]), .Z(n_300179391)
		);
	notech_or2 i_31841925(.A(n_54066), .B(n_26965), .Z(n_300879398));
	notech_or4 i_31541928(.A(n_59163), .B(n_26604), .C(n_26377), .D(n_27541)
		, .Z(n_301179401));
	notech_or2 i_31241931(.A(n_55536), .B(n_56820), .Z(n_301479404));
	notech_or2 i_33141912(.A(n_54066), .B(n_26967), .Z(n_302179411));
	notech_or4 i_32841915(.A(n_59163), .B(n_26604), .C(n_26377), .D(n_27542)
		, .Z(n_302479414));
	notech_or2 i_32541918(.A(n_55536), .B(n_56829), .Z(n_302779417));
	notech_nor2 i_33941904(.A(n_55555), .B(n_29165), .Z(n_303279422));
	notech_or4 i_33441909(.A(n_56163), .B(n_59277), .C(n_55523), .D(n_310818885
		), .Z(n_303979429));
	notech_nor2 i_36741876(.A(n_55555), .B(n_29167), .Z(n_304079430));
	notech_or4 i_36241881(.A(n_56163), .B(n_59277), .C(n_55523), .D(n_310718884
		), .Z(n_304779437));
	notech_nor2 i_37741868(.A(n_55555), .B(n_29169), .Z(n_304879438));
	notech_or4 i_37041873(.A(n_56163), .B(n_59277), .C(n_55523), .D(n_310618883
		), .Z(n_305579445));
	notech_nor2 i_38741860(.A(n_55555), .B(n_29172), .Z(n_305679446));
	notech_or4 i_38241865(.A(n_56163), .B(n_59277), .C(n_55523), .D(n_310518882
		), .Z(n_306379453));
	notech_nao3 i_40841840(.A(n_3383), .B(\eflags[10] ), .C(n_54046), .Z(n_306679456
		));
	notech_or2 i_40541843(.A(n_271688739), .B(n_56793), .Z(n_306979459));
	notech_nand3 i_40141846(.A(n_59179), .B(n_59936), .C(read_data[18]), .Z(n_307279462
		));
	notech_or2 i_39841849(.A(n_311318890), .B(n_355488242), .Z(n_307579465)
		);
	notech_nao3 i_42041828(.A(n_3385), .B(n_55460), .C(n_54046), .Z(n_307879468
		));
	notech_or2 i_41741831(.A(n_271688739), .B(n_56802), .Z(n_308179471));
	notech_nand3 i_41441834(.A(n_59179), .B(n_59936), .C(read_data[19]), .Z(n_308479474
		));
	notech_or2 i_41141837(.A(n_311218889), .B(n_355488242), .Z(n_308779477)
		);
	notech_nao3 i_43241816(.A(n_3387), .B(n_55460), .C(n_54707), .Z(n_309079480
		));
	notech_or2 i_42941819(.A(n_271688739), .B(n_56811), .Z(n_309379483));
	notech_nand3 i_42641822(.A(n_59179), .B(n_59936), .C(read_data[20]), .Z(n_309679486
		));
	notech_or2 i_42341825(.A(n_311118888), .B(n_355488242), .Z(n_309979489)
		);
	notech_nao3 i_44441804(.A(n_3389), .B(n_55460), .C(n_54046), .Z(n_310279492
		));
	notech_or2 i_44141807(.A(n_271688739), .B(n_56820), .Z(n_310579495));
	notech_nand3 i_43841810(.A(n_59176), .B(n_59936), .C(read_data[21]), .Z(n_310879498
		));
	notech_or2 i_43541813(.A(n_311018887), .B(n_355488242), .Z(n_311179501)
		);
	notech_nao3 i_45641792(.A(n_3391), .B(n_55460), .C(n_54046), .Z(n_311479504
		));
	notech_or2 i_45341795(.A(n_271688739), .B(n_56829), .Z(n_311779507));
	notech_nand3 i_45041798(.A(n_59176), .B(n_59936), .C(read_data[22]), .Z(n_312079510
		));
	notech_or2 i_44741801(.A(n_26618), .B(n_355488242), .Z(n_312379513));
	notech_or2 i_48641762(.A(n_311018887), .B(n_354969318), .Z(n_313279522)
		);
	notech_or2 i_49541753(.A(n_26618), .B(n_354969318), .Z(n_314179531));
	notech_nor2 i_57141679(.A(n_123423221), .B(nbus_11326[18]), .Z(n_314279532
		));
	notech_or2 i_56541684(.A(n_311318890), .B(n_2702), .Z(n_314979539));
	notech_nor2 i_58041671(.A(n_123423221), .B(nbus_11326[19]), .Z(n_315079540
		));
	notech_or2 i_57441676(.A(n_311218889), .B(n_2702), .Z(n_315779547));
	notech_nor2 i_58841663(.A(n_123423221), .B(nbus_11326[20]), .Z(n_315879548
		));
	notech_or2 i_58341668(.A(n_311118888), .B(n_2702), .Z(n_316579555));
	notech_nor2 i_59641655(.A(n_123423221), .B(nbus_11326[21]), .Z(n_316679556
		));
	notech_or2 i_59141660(.A(n_311018887), .B(n_2702), .Z(n_317379563));
	notech_or2 i_64841604(.A(n_353365822), .B(n_311318890), .Z(n_318179571)
		);
	notech_or2 i_66441588(.A(n_353365822), .B(n_311118888), .Z(n_318979579)
		);
	notech_nor2 i_78141476(.A(n_56216), .B(n_55609), .Z(n_319379583));
	notech_nor2 i_80741452(.A(n_56057), .B(\nbus_11276[20] ), .Z(n_319779587
		));
	notech_ao4 i_185340439(.A(n_101413408), .B(n_29169), .C(n_101213406), .D
		(n_311118888), .Z(n_319879588));
	notech_ao4 i_185240440(.A(n_98113375), .B(n_56811), .C(n_27540), .D(n_59809
		), .Z(n_320079590));
	notech_nao3 i_67742247(.A(n_319879588), .B(n_320079590), .C(n_319779587)
		, .Z(n_320179591));
	notech_ao4 i_183340459(.A(n_101413408), .B(n_29165), .C(n_101213406), .D
		(n_311318890), .Z(n_320279592));
	notech_ao4 i_183240460(.A(n_27538), .B(n_59791), .C(n_98113375), .D(n_56793
		), .Z(n_320479594));
	notech_nao3 i_67542249(.A(n_320279592), .B(n_320479594), .C(n_319379583)
		, .Z(n_320579595));
	notech_ao4 i_173840554(.A(n_121523202), .B(n_310618883), .C(n_121723204)
		, .D(n_315162155), .Z(n_320679596));
	notech_ao4 i_173740555(.A(n_353165820), .B(n_29169), .C(n_353465823), .D
		(n_27586), .Z(n_320879598));
	notech_and3 i_174040552(.A(n_320679596), .B(n_320879598), .C(n_318979579
		), .Z(n_320979599));
	notech_ao4 i_173540557(.A(n_353265821), .B(n_56811), .C(n_26572), .D(n_55631
		), .Z(n_321079600));
	notech_ao4 i_173440558(.A(n_121623203), .B(nbus_11326[20]), .C(n_27540),
		 .D(n_59791), .Z(n_321179601));
	notech_ao4 i_172440568(.A(n_121523202), .B(n_310818885), .C(n_121723204)
		, .D(n_310565422), .Z(n_321379603));
	notech_ao4 i_172340569(.A(n_353165820), .B(n_29165), .C(n_353465823), .D
		(n_27584), .Z(n_321579605));
	notech_and3 i_172640566(.A(n_321379603), .B(n_321579605), .C(n_318179571
		), .Z(n_321679606));
	notech_ao4 i_172040571(.A(n_353265821), .B(n_56793), .C(n_26572), .D(n_55609
		), .Z(n_321779607));
	notech_ao4 i_171940572(.A(n_27538), .B(n_59791), .C(n_121623203), .D(n_58969
		), .Z(n_321879608));
	notech_ao4 i_167340617(.A(n_310518882), .B(n_123223219), .C(n_312662130)
		, .D(n_123623223), .Z(n_322079610));
	notech_ao4 i_167240618(.A(n_29172), .B(n_26450), .C(n_181471126), .D(n_27588
		), .Z(n_322279612));
	notech_nand3 i_167540615(.A(n_322079610), .B(n_322279612), .C(n_317379563
		), .Z(n_322379613));
	notech_ao4 i_167040620(.A(n_55073), .B(n_56820), .C(n_55072), .D(\nbus_11276[21] 
		), .Z(n_322479614));
	notech_ao4 i_166640624(.A(n_310618883), .B(n_123223219), .C(n_315162155)
		, .D(n_123623223), .Z(n_322779617));
	notech_ao4 i_166540625(.A(n_29169), .B(n_26450), .C(n_181471126), .D(n_27586
		), .Z(n_322979619));
	notech_nand3 i_166840622(.A(n_322779617), .B(n_322979619), .C(n_316579555
		), .Z(n_323079620));
	notech_ao4 i_166240627(.A(n_55073), .B(n_56811), .C(n_55072), .D(n_55631
		), .Z(n_323179621));
	notech_ao4 i_165840631(.A(n_310718884), .B(n_123223219), .C(n_308065397)
		, .D(n_123623223), .Z(n_323479624));
	notech_ao4 i_165640632(.A(n_29167), .B(n_26450), .C(n_181471126), .D(n_27585
		), .Z(n_323679626));
	notech_nand3 i_166040629(.A(n_323479624), .B(n_323679626), .C(n_315779547
		), .Z(n_323779627));
	notech_ao4 i_165340634(.A(n_55073), .B(n_56802), .C(n_55072), .D(n_55620
		), .Z(n_323879628));
	notech_ao4 i_164840638(.A(n_310818885), .B(n_123223219), .C(n_310565422)
		, .D(n_123623223), .Z(n_324179631));
	notech_ao4 i_164740639(.A(n_29165), .B(n_26450), .C(n_181471126), .D(n_27584
		), .Z(n_324379633));
	notech_nand3 i_165040636(.A(n_324179631), .B(n_324379633), .C(n_314979539
		), .Z(n_324479634));
	notech_ao4 i_164540641(.A(n_55073), .B(n_56793), .C(n_55072), .D(n_55609
		), .Z(n_324579635));
	notech_ao4 i_159140695(.A(n_310418881), .B(n_354569315), .C(n_305565372)
		, .D(n_113113525), .Z(n_324879638));
	notech_ao4 i_159040696(.A(n_2193), .B(n_27542), .C(n_55776), .D(n_27589)
		, .Z(n_325079640));
	notech_and3 i_159340693(.A(n_324879638), .B(n_325079640), .C(n_314179531
		), .Z(n_325179641));
	notech_ao4 i_158840698(.A(n_354669316), .B(n_55647), .C(n_29174), .D(n_26571
		), .Z(n_325279642));
	notech_ao4 i_158740699(.A(n_113313527), .B(n_59032), .C(n_55562), .D(n_56829
		), .Z(n_325379643));
	notech_ao4 i_158440702(.A(n_310518882), .B(n_354569315), .C(n_312662130)
		, .D(n_113113525), .Z(n_325579645));
	notech_ao4 i_158340703(.A(n_58514), .B(n_27541), .C(n_55776), .D(n_27588
		), .Z(n_325779647));
	notech_and3 i_158640700(.A(n_325579645), .B(n_325779647), .C(n_313279522
		), .Z(n_325879648));
	notech_ao4 i_158040705(.A(n_354669316), .B(n_59310), .C(n_29172), .D(n_26571
		), .Z(n_325979649));
	notech_ao4 i_157940706(.A(n_113313527), .B(nbus_11326[21]), .C(n_55562),
		 .D(n_56820), .Z(n_326079650));
	notech_ao4 i_155440730(.A(n_310418881), .B(n_355788240), .C(n_305565372)
		, .D(n_353788271), .Z(n_326279652));
	notech_ao4 i_155240732(.A(n_320088489), .B(n_27589), .C(n_59176), .D(n_26732
		), .Z(n_326479654));
	notech_and4 i_155640728(.A(n_326479654), .B(n_326279652), .C(n_312079510
		), .D(n_312379513), .Z(n_326679656));
	notech_ao4 i_154940735(.A(n_271588740), .B(n_55647), .C(n_355688241), .D
		(n_29174), .Z(n_326779657));
	notech_ao4 i_154740737(.A(n_54024), .B(n_29452), .C(n_55133), .D(n_59032
		), .Z(n_326979659));
	notech_and4 i_155140733(.A(n_326979659), .B(n_326779657), .C(n_311479504
		), .D(n_311779507), .Z(n_327179661));
	notech_ao4 i_154440740(.A(n_310518882), .B(n_355788240), .C(n_312662130)
		, .D(n_353788271), .Z(n_327279662));
	notech_ao4 i_154240742(.A(n_320088489), .B(n_27588), .C(n_59176), .D(n_26731
		), .Z(n_327479664));
	notech_and4 i_154640738(.A(n_327479664), .B(n_327279662), .C(n_310879498
		), .D(n_311179501), .Z(n_327679666));
	notech_ao4 i_153940745(.A(n_271588740), .B(n_59310), .C(n_355688241), .D
		(n_29172), .Z(n_327779667));
	notech_ao4 i_153740747(.A(n_54024), .B(n_29451), .C(n_55133), .D(n_58996
		), .Z(n_327979669));
	notech_and4 i_154140743(.A(n_327979669), .B(n_327779667), .C(n_310279492
		), .D(n_310579495), .Z(n_328179671));
	notech_ao4 i_153440750(.A(n_310618883), .B(n_355788240), .C(n_315162155)
		, .D(n_353788271), .Z(n_328279672));
	notech_ao4 i_153240752(.A(n_320088489), .B(n_27586), .C(n_59176), .D(n_26730
		), .Z(n_328479674));
	notech_and4 i_153640748(.A(n_328479674), .B(n_328279672), .C(n_309679486
		), .D(n_309979489), .Z(n_328679676));
	notech_ao4 i_152940755(.A(n_271588740), .B(n_55631), .C(n_355688241), .D
		(n_29169), .Z(n_328779677));
	notech_ao4 i_152640757(.A(n_54024), .B(n_29450), .C(n_55133), .D(nbus_11326
		[20]), .Z(n_328979679));
	notech_and4 i_153140753(.A(n_328979679), .B(n_328779677), .C(n_309079480
		), .D(n_309379483), .Z(n_329179681));
	notech_ao4 i_152340760(.A(n_310718884), .B(n_355788240), .C(n_308065397)
		, .D(n_353788271), .Z(n_329279682));
	notech_ao4 i_152140762(.A(n_320088489), .B(n_27585), .C(n_59176), .D(n_26729
		), .Z(n_329479684));
	notech_and4 i_152540758(.A(n_329479684), .B(n_329279682), .C(n_308479474
		), .D(n_308779477), .Z(n_329679686));
	notech_ao4 i_151840765(.A(n_271588740), .B(n_55620), .C(n_355688241), .D
		(n_29167), .Z(n_329779687));
	notech_ao4 i_151640767(.A(n_54024), .B(n_29449), .C(n_55133), .D(nbus_11326
		[19]), .Z(n_329979689));
	notech_and4 i_152040763(.A(n_329979689), .B(n_329779687), .C(n_307879468
		), .D(n_308179471), .Z(n_330179691));
	notech_ao4 i_151340770(.A(n_310818885), .B(n_355788240), .C(n_310565422)
		, .D(n_353788271), .Z(n_330279692));
	notech_ao4 i_151140772(.A(n_320088489), .B(n_27584), .C(n_59174), .D(n_26728
		), .Z(n_330479694));
	notech_and4 i_151540768(.A(n_330479694), .B(n_330279692), .C(n_307279462
		), .D(n_307579465), .Z(n_330679696));
	notech_ao4 i_150840775(.A(n_271588740), .B(n_55609), .C(n_355688241), .D
		(n_29165), .Z(n_330779697));
	notech_ao4 i_150640777(.A(n_54024), .B(n_29448), .C(n_55133), .D(n_58969
		), .Z(n_330979699));
	notech_and4 i_151040773(.A(n_330979699), .B(n_330779697), .C(n_306679456
		), .D(n_306979459), .Z(n_331179701));
	notech_ao4 i_149640787(.A(n_312662130), .B(n_308718864), .C(n_308318860)
		, .D(n_58996), .Z(n_331279702));
	notech_ao4 i_149540788(.A(n_55773), .B(n_27588), .C(n_311018887), .D(n_55554
		), .Z(n_331479704));
	notech_nand3 i_149840785(.A(n_331279702), .B(n_331479704), .C(n_306379453
		), .Z(n_331579705));
	notech_ao4 i_149340790(.A(n_55219), .B(n_56820), .C(n_55218), .D(n_59310
		), .Z(n_331679706));
	notech_ao4 i_148840794(.A(n_315162155), .B(n_308718864), .C(n_308318860)
		, .D(n_59005), .Z(n_331979709));
	notech_ao4 i_148740795(.A(n_55773), .B(n_27586), .C(n_311118888), .D(n_55554
		), .Z(n_332179711));
	notech_nand3 i_149140792(.A(n_331979709), .B(n_332179711), .C(n_305579445
		), .Z(n_332279712));
	notech_ao4 i_148540797(.A(n_55219), .B(n_56811), .C(n_55218), .D(n_55631
		), .Z(n_332379713));
	notech_ao4 i_148140801(.A(n_308065397), .B(n_308718864), .C(n_308318860)
		, .D(nbus_11326[19]), .Z(n_332679716));
	notech_ao4 i_148040802(.A(n_55773), .B(n_27585), .C(n_311218889), .D(n_55554
		), .Z(n_332879718));
	notech_nand3 i_148340799(.A(n_332679716), .B(n_332879718), .C(n_304779437
		), .Z(n_332979719));
	notech_ao4 i_147840804(.A(n_55219), .B(n_56802), .C(n_55218), .D(n_55620
		), .Z(n_333079720));
	notech_ao4 i_139540881(.A(n_310565422), .B(n_308718864), .C(n_308318860)
		, .D(n_58969), .Z(n_333379723));
	notech_ao4 i_139440882(.A(n_55773), .B(n_27584), .C(n_311318890), .D(n_55554
		), .Z(n_333579725));
	notech_nand3 i_139740879(.A(n_333379723), .B(n_333579725), .C(n_303979429
		), .Z(n_333679726));
	notech_ao4 i_139240884(.A(n_55219), .B(n_56793), .C(n_55218), .D(n_55609
		), .Z(n_333779727));
	notech_ao4 i_138840888(.A(n_305565372), .B(n_308618863), .C(n_308518862)
		, .D(n_59032), .Z(n_334079730));
	notech_ao4 i_138740889(.A(n_26618), .B(n_55442), .C(n_310418881), .D(n_55780
		), .Z(n_334179731));
	notech_ao4 i_138540891(.A(n_55535), .B(n_55647), .C(n_55443), .D(n_29174
		), .Z(n_334379733));
	notech_and4 i_139040886(.A(n_334379733), .B(n_334179731), .C(n_334079730
		), .D(n_302779417), .Z(n_334579735));
	notech_ao4 i_138240894(.A(n_55135), .B(n_27589), .C(n_59172), .D(n_26707
		), .Z(n_334679736));
	notech_ao4 i_138040896(.A(n_54080), .B(n_28436), .C(n_54092), .D(n_29447
		), .Z(n_334879738));
	notech_and4 i_138440892(.A(n_334879738), .B(n_334679736), .C(n_302179411
		), .D(n_302479414), .Z(n_335079740));
	notech_ao4 i_137740899(.A(n_312662130), .B(n_308618863), .C(n_308518862)
		, .D(n_58996), .Z(n_335179741));
	notech_ao4 i_137640900(.A(n_311018887), .B(n_55442), .C(n_55780), .D(n_310518882
		), .Z(n_335279742));
	notech_ao4 i_137440902(.A(n_55535), .B(n_59310), .C(n_55443), .D(n_29172
		), .Z(n_335479744));
	notech_and4 i_137940897(.A(n_335479744), .B(n_335279742), .C(n_335179741
		), .D(n_301479404), .Z(n_335679746));
	notech_ao4 i_137140905(.A(n_55135), .B(n_27588), .C(n_59172), .D(n_26706
		), .Z(n_335779747));
	notech_ao4 i_136940907(.A(n_54080), .B(n_28435), .C(n_54092), .D(n_29444
		), .Z(n_336179749));
	notech_and4 i_137340903(.A(n_336179749), .B(n_335779747), .C(n_300879398
		), .D(n_301179401), .Z(n_336379751));
	notech_ao4 i_136640910(.A(n_315162155), .B(n_308618863), .C(n_308518862)
		, .D(n_59005), .Z(n_336479752));
	notech_ao4 i_136540911(.A(n_311118888), .B(n_55442), .C(n_55780), .D(n_310618883
		), .Z(n_336579753));
	notech_ao4 i_136340913(.A(n_55535), .B(n_55631), .C(n_29169), .D(n_55443
		), .Z(n_336779755));
	notech_and4 i_136840908(.A(n_336779755), .B(n_336579753), .C(n_336479752
		), .D(n_300179391), .Z(n_336979757));
	notech_ao4 i_136040916(.A(n_55135), .B(n_27586), .C(n_59172), .D(n_26705
		), .Z(n_337079758));
	notech_ao4 i_135840918(.A(n_54080), .B(n_28434), .C(n_54092), .D(n_29443
		), .Z(n_337279760));
	notech_and4 i_136240914(.A(n_337279760), .B(n_337079758), .C(n_299579385
		), .D(n_299879388), .Z(n_337479762));
	notech_ao4 i_135540921(.A(n_308065397), .B(n_308618863), .C(n_308518862)
		, .D(n_59014), .Z(n_337579763));
	notech_ao4 i_135440922(.A(n_311218889), .B(n_55442), .C(n_55780), .D(n_310718884
		), .Z(n_337679764));
	notech_ao4 i_135240924(.A(n_55535), .B(n_55620), .C(n_55443), .D(n_29167
		), .Z(n_337879766));
	notech_and4 i_135740919(.A(n_337879766), .B(n_337679764), .C(n_337579763
		), .D(n_298879378), .Z(n_338079768));
	notech_ao4 i_134940927(.A(n_55135), .B(n_27585), .C(n_59172), .D(n_26704
		), .Z(n_338179769));
	notech_ao4 i_134740929(.A(n_54080), .B(n_28433), .C(n_54092), .D(n_29442
		), .Z(n_340779771));
	notech_and4 i_135140925(.A(n_340779771), .B(n_338179769), .C(n_298279372
		), .D(n_298579375), .Z(n_340979773));
	notech_ao4 i_134440932(.A(n_310565422), .B(n_308618863), .C(n_308518862)
		, .D(n_58969), .Z(n_341079774));
	notech_ao4 i_134340933(.A(n_311318890), .B(n_55442), .C(n_55780), .D(n_310818885
		), .Z(n_341179775));
	notech_ao4 i_134140935(.A(n_55535), .B(n_55609), .C(n_55443), .D(n_29165
		), .Z(n_341379777));
	notech_and4 i_134640930(.A(n_341379777), .B(n_341179775), .C(n_341079774
		), .D(n_297579365), .Z(n_341579779));
	notech_ao4 i_133840938(.A(n_55135), .B(n_27584), .C(n_59172), .D(n_26703
		), .Z(n_341679780));
	notech_ao4 i_133640940(.A(n_54080), .B(n_28432), .C(n_54092), .D(n_29441
		), .Z(n_341879782));
	notech_and4 i_134040936(.A(n_341879782), .B(n_341679780), .C(n_296979359
		), .D(n_297279362), .Z(n_342079784));
	notech_ao4 i_132540951(.A(n_310518882), .B(n_322631613), .C(n_312662130)
		, .D(n_322931616), .Z(n_342179785));
	notech_ao4 i_132440952(.A(n_55557), .B(n_29172), .C(n_55772), .D(n_27588
		), .Z(n_342679787));
	notech_ao4 i_132040955(.A(n_55220), .B(n_56820), .C(n_55221), .D(n_59310
		), .Z(n_342979789));
	notech_and4 i_132340953(.A(n_53844), .B(n_342979789), .C(n_296179351), .D
		(n_26416), .Z(n_344479792));
	notech_ao4 i_131640959(.A(n_310618883), .B(n_322631613), .C(n_315162155)
		, .D(n_322931616), .Z(n_344579793));
	notech_ao4 i_131540960(.A(n_55557), .B(n_29169), .C(n_55772), .D(n_27586
		), .Z(n_344779795));
	notech_nand3 i_131840957(.A(n_344579793), .B(n_344779795), .C(n_295879348
		), .Z(n_344879796));
	notech_ao4 i_131340962(.A(n_55220), .B(n_56811), .C(n_55221), .D(n_55631
		), .Z(n_344979797));
	notech_ao4 i_130940966(.A(n_310718884), .B(n_322631613), .C(n_308065397)
		, .D(n_322931616), .Z(n_345279800));
	notech_ao4 i_130840967(.A(n_55557), .B(n_29167), .C(n_55772), .D(n_27585
		), .Z(n_345479802));
	notech_ao4 i_130540970(.A(n_55220), .B(n_56802), .C(n_55221), .D(n_55620
		), .Z(n_345679804));
	notech_and4 i_130740968(.A(n_53844), .B(n_345679804), .C(n_294579335), .D
		(n_26417), .Z(n_345979807));
	notech_ao4 i_130140974(.A(n_310818885), .B(n_322631613), .C(n_310565422)
		, .D(n_322931616), .Z(n_346079808));
	notech_ao4 i_130040975(.A(n_55557), .B(n_29165), .C(n_55772), .D(n_27584
		), .Z(n_346279810));
	notech_ao4 i_129740978(.A(n_55220), .B(n_56793), .C(n_55221), .D(n_55609
		), .Z(n_346479812));
	notech_and4 i_129940976(.A(n_53844), .B(n_346479812), .C(n_293779327), .D
		(n_26492), .Z(n_346779815));
	notech_ao4 i_119441080(.A(n_310418881), .B(n_3214), .C(n_305565372), .D(n_321588475
		), .Z(n_346879816));
	notech_ao4 i_119241082(.A(n_131423301), .B(n_27589), .C(n_59172), .D(n_26657
		), .Z(n_347079818));
	notech_and4 i_119641078(.A(n_347079818), .B(n_346879816), .C(n_293179321
		), .D(n_293479324), .Z(n_347279820));
	notech_ao4 i_118941085(.A(n_55533), .B(n_55647), .C(n_321388476), .D(n_29174
		), .Z(n_347379821));
	notech_ao4 i_118741087(.A(n_55131), .B(n_29440), .C(n_131123298), .D(n_59032
		), .Z(n_347579823));
	notech_and4 i_119141083(.A(n_54860), .B(n_347579823), .C(n_347379821), .D
		(n_292879318), .Z(n_347779825));
	notech_ao4 i_118441090(.A(n_310518882), .B(n_3214), .C(n_312662130), .D(n_321588475
		), .Z(n_347879826));
	notech_ao4 i_118241092(.A(n_131423301), .B(n_27588), .C(n_59172), .D(n_26655
		), .Z(n_348079828));
	notech_and4 i_118641088(.A(n_348079828), .B(n_347879826), .C(n_292079310
		), .D(n_292379313), .Z(n_348279830));
	notech_ao4 i_117941095(.A(n_55533), .B(n_59310), .C(n_321388476), .D(n_29172
		), .Z(n_348379831));
	notech_ao4 i_117741097(.A(n_55131), .B(n_29439), .C(n_131123298), .D(n_58996
		), .Z(n_348579833));
	notech_and4 i_118141093(.A(n_54860), .B(n_348579833), .C(n_348379831), .D
		(n_291779307), .Z(n_348779835));
	notech_ao4 i_117441100(.A(n_310618883), .B(n_3214), .C(n_315162155), .D(n_321588475
		), .Z(n_348879836));
	notech_ao4 i_117241102(.A(n_131423301), .B(n_27586), .C(n_59172), .D(n_26654
		), .Z(n_349079838));
	notech_and4 i_117641098(.A(n_349079838), .B(n_348879836), .C(n_290979299
		), .D(n_291279302), .Z(n_349279840));
	notech_ao4 i_116941105(.A(n_55533), .B(n_55631), .C(n_321388476), .D(n_29169
		), .Z(n_349379841));
	notech_ao4 i_116841106(.A(n_55131), .B(n_29438), .C(n_131123298), .D(n_59005
		), .Z(n_349579843));
	notech_ao4 i_116541109(.A(n_310718884), .B(n_3214), .C(n_308065397), .D(n_321588475
		), .Z(n_349779845));
	notech_ao4 i_116341111(.A(n_131423301), .B(n_27585), .C(n_59172), .D(n_26653
		), .Z(n_349979847));
	notech_and4 i_116741107(.A(n_349979847), .B(n_349779845), .C(n_289879288
		), .D(n_290179291), .Z(n_350179849));
	notech_ao4 i_116041114(.A(n_55533), .B(n_55620), .C(n_321388476), .D(n_29167
		), .Z(n_350279850));
	notech_ao4 i_115941115(.A(n_55131), .B(n_29437), .C(n_131123298), .D(n_59014
		), .Z(n_350479852));
	notech_or2 i_124537906(.A(n_354969318), .B(n_2700), .Z(n_350679854));
	notech_nand2 i_1821309(.A(n_354579893), .B(n_350679854), .Z(n_20703));
	notech_or2 i_157537580(.A(n_2320), .B(n_2700), .Z(n_351579863));
	notech_and3 i_156437591(.A(n_2219), .B(resb_shift4box[17]), .C(n_274788710
		), .Z(n_351679864));
	notech_and4 i_1816187(.A(n_354779895), .B(n_354679894), .C(n_355579903),
		 .D(n_351579863), .Z(n_14194));
	notech_or2 i_159937556(.A(n_271988736), .B(n_2320), .Z(n_352779875));
	notech_and3 i_158837567(.A(resb_shift4box[16]), .B(n_274788710), .C(n_2219
		), .Z(n_352879876));
	notech_and4 i_1716186(.A(n_355879906), .B(n_355779905), .C(n_356779914),
		 .D(n_352779875), .Z(n_14188));
	notech_ao4 i_124637905(.A(n_63826342), .B(n_113113525), .C(n_58514), .D(n_27537
		), .Z(n_353979887));
	notech_ao4 i_124737904(.A(n_55776), .B(n_27583), .C(n_58978), .D(n_113313527
		), .Z(n_354079888));
	notech_ao4 i_124837903(.A(n_26571), .B(n_28987), .C(n_354569315), .D(n_2648
		), .Z(n_354279890));
	notech_ao4 i_124937902(.A(n_354669316), .B(n_55600), .C(n_55562), .D(n_56784
		), .Z(n_354379891));
	notech_and4 i_125237899(.A(n_354379891), .B(n_354279890), .C(n_354079888
		), .D(n_353979887), .Z(n_354579893));
	notech_ao4 i_158037575(.A(n_2323), .B(n_27583), .C(n_2164), .D(n_58978),
		 .Z(n_354679894));
	notech_ao4 i_158137574(.A(n_55933), .B(n_55600), .C(n_2322), .D(n_56784)
		, .Z(n_354779895));
	notech_ao4 i_157737578(.A(n_55366), .B(n_28791), .C(n_2319), .D(n_29023)
		, .Z(n_355079898));
	notech_ao3 i_158237573(.A(n_2187), .B(n_355079898), .C(n_351679864), .Z(n_355179899
		));
	notech_ao4 i_157837577(.A(n_55619), .B(n_28628), .C(n_55526), .D(n_28596
		), .Z(n_355279900));
	notech_ao4 i_157937576(.A(n_55243), .B(n_27537), .C(n_2318), .D(n_28847)
		, .Z(n_355379901));
	notech_and3 i_158537570(.A(n_355379901), .B(n_355279900), .C(n_355179899
		), .Z(n_355579903));
	notech_ao4 i_160437551(.A(n_55243), .B(n_27535), .C(n_55933), .D(n_55590
		), .Z(n_355779905));
	notech_ao4 i_160537550(.A(n_2319), .B(n_29020), .C(n_2323), .D(n_27582),
		 .Z(n_355879906));
	notech_ao4 i_160137554(.A(n_55526), .B(n_28592), .C(n_55366), .D(n_28790
		), .Z(n_356179909));
	notech_ao3 i_160637549(.A(n_2187), .B(n_356179909), .C(n_352879876), .Z(n_356279910
		));
	notech_ao4 i_160237553(.A(n_2318), .B(n_28846), .C(n_55619), .D(n_28627)
		, .Z(n_356379911));
	notech_ao4 i_160337552(.A(n_2322), .B(n_56775), .C(n_2164), .D(n_58987),
		 .Z(n_356479912));
	notech_and3 i_160937546(.A(n_356479912), .B(n_356379911), .C(n_356279910
		), .Z(n_356779914));
	notech_and2 i_13335572(.A(n_336165663), .B(n_2822), .Z(n_357179916));
	notech_nand2 i_117034579(.A(n_1862), .B(n_55656), .Z(n_357279917));
	notech_nor2 i_15835569(.A(n_494), .B(n_357179916), .Z(n_357379918));
	notech_or4 i_19213(.A(fsm[3]), .B(fsm[0]), .C(n_60780), .D(n_59753), .Z(n_357479919
		));
	notech_nor2 i_120234550(.A(n_360779952), .B(n_357379918), .Z(n_357579920
		));
	notech_and4 i_119834552(.A(n_2224), .B(n_276188696), .C(n_26419), .D(n_54892
		), .Z(n_357979924));
	notech_nand2 i_54532898(.A(n_361879963), .B(n_59791), .Z(n_358079925));
	notech_and3 i_66733151(.A(n_354276378), .B(n_361379958), .C(n_2268), .Z(n_358179926
		));
	notech_and4 i_15132728(.A(n_2823), .B(n_2822), .C(n_55641), .D(n_362079965
		), .Z(n_358279927));
	notech_and2 i_23232684(.A(Daddrs_1[0]), .B(n_54701), .Z(n_358579930));
	notech_ao3 i_22732687(.A(n_55040), .B(Daddrs_8[0]), .C(n_55149), .Z(n_358879933
		));
	notech_and3 i_22432690(.A(n_361879963), .B(Daddrgs[0]), .C(n_59791), .Z(n_359179936
		));
	notech_or4 i_21432695(.A(n_60780), .B(n_60731), .C(n_55342), .D(n_358179926
		), .Z(n_359279937));
	notech_or4 i_21532694(.A(n_274988708), .B(n_1901), .C(n_55356), .D(n_59936
		), .Z(n_359379938));
	notech_ao3 i_22032693(.A(n_316188528), .B(n_5153), .C(n_315388536), .Z(n_359479939
		));
	notech_or2 i_25832663(.A(n_54771), .B(n_56943), .Z(n_359779942));
	notech_or2 i_25232666(.A(n_54674), .B(n_27984), .Z(n_360079945));
	notech_or4 i_24932669(.A(n_275288705), .B(n_205588858), .C(n_59936), .D(n_59095
		), .Z(n_360379948));
	notech_nao3 i_24532672(.A(Daddrs_3[31]), .B(n_26613), .C(n_315388536), .Z
		(n_360679951));
	notech_and3 i_5398(.A(n_59172), .B(n_59795), .C(n_357279917), .Z(n_360779952
		));
	notech_or4 i_27532647(.A(n_190388902), .B(n_613), .C(n_2265), .D(n_57451
		), .Z(n_360979954));
	notech_or4 i_27632646(.A(n_2793), .B(n_58514), .C(n_358279927), .D(n_60579
		), .Z(n_361079955));
	notech_or4 i_60632391(.A(n_272688729), .B(n_272988726), .C(n_26600), .D(n_26593
		), .Z(n_361379958));
	notech_and3 i_118531894(.A(n_364988146), .B(over_seg[5]), .C(n_60138), .Z
		(n_361879963));
	notech_mux2 i_82332204(.S(read_ack), .A(n_57434), .B(n_2824), .Z(n_362079965
		));
	notech_ao4 i_81432213(.A(n_2209), .B(n_352676362), .C(n_58523), .D(n_60579
		), .Z(n_362379968));
	notech_nand3 i_81632211(.A(n_360979954), .B(n_362379968), .C(n_361079955
		), .Z(n_362479969));
	notech_ao4 i_78032242(.A(n_310288586), .B(n_29457), .C(n_54714), .D(n_29456
		), .Z(n_362779972));
	notech_ao4 i_77832244(.A(n_2234), .B(n_29455), .C(n_27295), .D(n_58523),
		 .Z(n_362979974));
	notech_and4 i_78532240(.A(n_362979974), .B(n_362779972), .C(n_360379948)
		, .D(n_360679951), .Z(n_363179976));
	notech_ao4 i_77532247(.A(n_54659), .B(n_28445), .C(n_54642), .D(n_28455)
		, .Z(n_363279977));
	notech_ao4 i_77332249(.A(n_54742), .B(n_27601), .C(n_55792), .D(n_28454)
		, .Z(n_363479979));
	notech_and4 i_77732245(.A(n_363479979), .B(n_363279977), .C(n_359779942)
		, .D(n_360079945), .Z(n_363679981));
	notech_nao3 i_74432276(.A(n_359379938), .B(n_359279937), .C(n_359479939)
		, .Z(n_363979984));
	notech_ao4 i_74132279(.A(n_54685), .B(n_28456), .C(n_310288586), .D(n_29454
		), .Z(n_364079985));
	notech_ao4 i_73732282(.A(n_54727), .B(nbus_11326[0]), .C(n_2234), .D(n_29453
		), .Z(n_364379988));
	notech_ao4 i_73532284(.A(n_54674), .B(n_27953), .C(n_54659), .D(n_28414)
		, .Z(n_364579990));
	notech_or4 i_74032280(.A(n_358879933), .B(n_358579930), .C(n_26472), .D(n_26471
		), .Z(n_364779992));
	notech_nand3 i_106388441(.A(over_seg[5]), .B(n_60138), .C(n_364988146), 
		.Z(n_364888147));
	notech_nand2 i_128788442(.A(n_276588692), .B(n_273388722), .Z(n_364988146
		));
	notech_or4 i_106788443(.A(n_60780), .B(n_60731), .C(n_60579), .D(n_365188144
		), .Z(n_365088145));
	notech_ao3 i_12888444(.A(n_58886), .B(n_364888147), .C(n_58591), .Z(n_365188144
		));
	notech_or2 i_106488447(.A(n_276488693), .B(read_ack), .Z(n_365488141));
	notech_nand3 i_526955(.A(n_276188696), .B(n_365788138), .C(n_365088145),
		 .Z(n_14920));
	notech_ao4 i_106888448(.A(n_494), .B(n_366088135), .C(n_57458), .D(n_54770
		), .Z(n_365588140));
	notech_and4 i_107088450(.A(n_55763), .B(n_365588140), .C(n_2406), .D(n_365488141
		), .Z(n_365788138));
	notech_nand2 i_54742(.A(n_163460716), .B(n_121777617), .Z(\nbus_11353[12] 
		));
	notech_ao4 i_53386(.A(n_55642), .B(n_56076), .C(n_121477614), .D(n_60474
		), .Z(n_18859));
	notech_nao3 i_48863(.A(n_219961272), .B(n_270739495), .C(n_126277662), .Z
		(\nbus_11305[16] ));
	notech_and4 i_521584(.A(n_126577665), .B(n_126777667), .C(n_127177671), 
		.D(n_126177661), .Z(n_13139));
	notech_nand2 i_1821725(.A(n_128277682), .B(n_127777677), .Z(n_12869));
	notech_nand2 i_1021717(.A(n_129377693), .B(n_128877688), .Z(n_12821));
	notech_and4 i_521904(.A(n_129477694), .B(n_129677696), .C(n_130177701), 
		.D(n_122777627), .Z(n_12073));
	notech_nand2 i_205060618(.A(read_data[6]), .B(n_59936), .Z(n_54470));
	notech_or4 i_1020661(.A(n_26423), .B(n_137277772), .C(n_138077780), .D(n_26424
		), .Z(n_19839));
	notech_and4 i_1020981(.A(n_138277782), .B(n_138477784), .C(n_136577765),
		 .D(n_138877788), .Z(n_16753));
	notech_nand2 i_3021577(.A(n_139977799), .B(n_139477794), .Z(n_16524));
	notech_and4 i_721554(.A(n_134077740), .B(n_140577805), .C(n_140877808), 
		.D(n_140477804), .Z(n_16386));
	notech_or4 i_921588(.A(n_132877728), .B(n_145974327), .C(n_141377813), .D
		(n_26425), .Z(n_13163));
	notech_or4 i_1021845(.A(n_185167671), .B(n_132177721), .C(n_142077820), 
		.D(n_26426), .Z(n_12455));
	notech_nand2 i_721906(.A(n_143277832), .B(n_142877828), .Z(n_12085));
	notech_nand2 i_1017236(.A(n_144177841), .B(n_143777837), .Z(n_15828));
	notech_ao4 i_176737389(.A(n_55122), .B(n_59328), .C(n_55111), .D(nbus_11326
		[3]), .Z(n_279359037));
	notech_and2 i_62057980(.A(n_55773), .B(n_145077850), .Z(n_55730));
	notech_ao4 i_177137385(.A(n_55526), .B(n_28577), .C(n_55102), .D(n_28785
		), .Z(n_279159035));
	notech_and4 i_720978(.A(n_182878223), .B(n_183778232), .C(n_183978234), 
		.D(n_184478239), .Z(n_16735));
	notech_and4 i_721586(.A(n_181778214), .B(n_184578240), .C(n_184778242), 
		.D(n_185178246), .Z(n_13151));
	notech_nand2 i_3117577(.A(n_186178256), .B(n_185678251), .Z(n_21023));
	notech_nand2 i_3017576(.A(n_187178266), .B(n_186678261), .Z(n_21017));
	notech_nand2 i_2917575(.A(n_188178276), .B(n_187678271), .Z(n_21011));
	notech_nand2 i_2817574(.A(n_189178286), .B(n_188678281), .Z(n_21005));
	notech_nand2 i_2717573(.A(n_190178296), .B(n_189678291), .Z(n_20999));
	notech_nand2 i_2617572(.A(n_191178306), .B(n_190678301), .Z(n_20993));
	notech_nand2 i_2517571(.A(n_192178316), .B(n_191678311), .Z(n_20987));
	notech_nand2 i_2417570(.A(n_193178326), .B(n_192678321), .Z(n_20981));
	notech_nand2 i_2317569(.A(n_194178336), .B(n_193678331), .Z(n_20975));
	notech_nand2 i_2217568(.A(n_195178346), .B(n_194678341), .Z(n_20969));
	notech_nand2 i_2117567(.A(n_196178356), .B(n_195678351), .Z(n_20963));
	notech_nand2 i_2017566(.A(n_197178366), .B(n_196678361), .Z(n_20957));
	notech_nand2 i_1917565(.A(n_198178376), .B(n_197678371), .Z(n_20951));
	notech_nand2 i_1817564(.A(n_199178386), .B(n_198678381), .Z(n_20945));
	notech_nand2 i_1617562(.A(n_200178396), .B(n_199678391), .Z(n_20933));
	notech_nand2 i_1517561(.A(n_201178406), .B(n_200678401), .Z(n_20927));
	notech_nand2 i_1417560(.A(n_202178416), .B(n_201678411), .Z(n_20921));
	notech_nand2 i_1317559(.A(n_203178426), .B(n_202678421), .Z(n_20915));
	notech_nand2 i_1217558(.A(n_204178436), .B(n_203678431), .Z(n_20909));
	notech_nand2 i_1117557(.A(n_205178446), .B(n_204678441), .Z(n_20903));
	notech_nand2 i_1017556(.A(n_206278457), .B(n_205778452), .Z(n_20897));
	notech_nand2 i_917555(.A(n_206878463), .B(n_207378468), .Z(n_20891));
	notech_nand2 i_817554(.A(n_208478479), .B(n_207978474), .Z(n_20885));
	notech_nand2 i_717553(.A(n_209578490), .B(n_209078485), .Z(n_20879));
	notech_nand2 i_617552(.A(n_210678501), .B(n_210178496), .Z(n_20873));
	notech_nand2 i_517551(.A(n_211278507), .B(n_211778512), .Z(n_20867));
	notech_nand2 i_417550(.A(n_212878523), .B(n_212378518), .Z(n_20861));
	notech_or4 i_317549(.A(n_147177871), .B(n_213178526), .C(n_213978534), .D
		(n_26428), .Z(n_20855));
	notech_or4 i_217548(.A(n_145977859), .B(n_214478538), .C(n_215278546), .D
		(n_26431), .Z(n_20849));
	notech_or2 i_130257864(.A(n_144977849), .B(n_294261946), .Z(n_248734113)
		);
	notech_ao4 i_177037386(.A(n_55243), .B(n_27530), .C(n_2164), .D(nbus_11326
		[11]), .Z(n_279059034));
	notech_ao4 i_178137376(.A(n_89513289), .B(n_27595), .C(n_88913283), .D(n_28841
		), .Z(n_278959033));
	notech_mux2 i_1611673(.S(n_60138), .A(n_571), .B(add_len_pc32[15]), .Z(\add_len_pc[15] 
		));
	notech_mux2 i_2511682(.S(n_60138), .A(regs_14[24]), .B(add_len_pc32[24])
		, .Z(\add_len_pc[24] ));
	notech_nand2 i_2520644(.A(n_235178741), .B(n_234678736), .Z(n_20255));
	notech_nand2 i_1620635(.A(n_236178751), .B(n_235678746), .Z(n_20201));
	notech_and4 i_1120662(.A(n_154070859), .B(n_236678756), .C(n_231078700),
		 .D(n_236578755), .Z(n_19845));
	notech_or4 i_2521060(.A(n_252861556), .B(n_230278692), .C(n_237278762), 
		.D(n_26436), .Z(n_13959));
	notech_nand3 i_2521316(.A(n_238178771), .B(n_238078770), .C(n_237978769)
		, .Z(n_20745));
	notech_nand2 i_2521572(.A(n_239278782), .B(n_238778777), .Z(n_16494));
	notech_or4 i_2521604(.A(n_252861556), .B(n_227378663), .C(n_239678786), 
		.D(n_26438), .Z(n_13259));
	notech_and4 i_1621595(.A(n_363088165), .B(n_226478655), .C(n_240478794),
		 .D(n_240378793), .Z(n_13205));
	notech_or4 i_1321592(.A(n_189974767), .B(n_225678647), .C(n_241078800), 
		.D(n_26439), .Z(n_13187));
	notech_or4 i_1221591(.A(n_239168196), .B(n_224878639), .C(n_241778807), 
		.D(n_26440), .Z(n_13181));
	notech_nand3 i_1121590(.A(n_242278812), .B(n_242178811), .C(n_242678816)
		, .Z(n_13175));
	notech_nand2 i_2521732(.A(n_243778827), .B(n_243278822), .Z(n_12911));
	notech_nand2 i_1421721(.A(n_244878838), .B(n_244378833), .Z(n_12845));
	notech_nand2 i_1221719(.A(n_245978849), .B(n_245478844), .Z(n_12833));
	notech_nand2 i_921716(.A(n_247078860), .B(n_246578855), .Z(n_12815));
	notech_or4 i_1321848(.A(n_189974767), .B(n_217878572), .C(n_247478864), 
		.D(n_26441), .Z(n_12473));
	notech_and4 i_1121846(.A(n_53844), .B(n_248378873), .C(n_154070859), .D(n_248278872
		), .Z(n_12461));
	notech_and4 i_2516674(.A(n_249178881), .B(n_249378883), .C(n_249078880),
		 .D(n_216378557), .Z(n_11836));
	notech_and4 i_174737409(.A(n_278459028), .B(n_242658670), .C(n_242258666
		), .D(n_242358667), .Z(n_278759031));
	notech_and2 i_18085(.A(opb[4]), .B(n_59795), .Z(n_365988136));
	notech_nand3 i_2421315(.A(n_276179151), .B(n_276079150), .C(n_275979149)
		, .Z(n_20739));
	notech_nand2 i_2921576(.A(n_277279162), .B(n_276779157), .Z(n_16518));
	notech_nand2 i_2821575(.A(n_278279172), .B(n_277779167), .Z(n_16512));
	notech_nand2 i_2721574(.A(n_279279182), .B(n_278779177), .Z(n_16506));
	notech_nand2 i_2621573(.A(n_280279192), .B(n_279779187), .Z(n_16500));
	notech_nand2 i_2421571(.A(n_281279202), .B(n_280779197), .Z(n_16488));
	notech_or4 i_2421603(.A(n_267675515), .B(n_267979069), .C(n_281679206), 
		.D(n_26448), .Z(n_13253));
	notech_nand2 i_2921736(.A(n_283079220), .B(n_282579215), .Z(n_12935));
	notech_nand2 i_2821735(.A(n_284179231), .B(n_283679226), .Z(n_12929));
	notech_nand2 i_2721734(.A(n_285279242), .B(n_284779237), .Z(n_12923));
	notech_nand2 i_2621733(.A(n_286379253), .B(n_285879248), .Z(n_12917));
	notech_nand2 i_2421731(.A(n_287479264), .B(n_286979259), .Z(n_12905));
	notech_or4 i_2421859(.A(n_267675515), .B(n_260678996), .C(n_287879268), 
		.D(n_26449), .Z(n_12539));
	notech_and4 i_2416673(.A(n_288779277), .B(n_288979279), .C(n_288679276),
		 .D(n_259978989), .Z(n_11830));
	notech_and4 i_174337413(.A(n_277559019), .B(n_277459018), .C(n_278259026
		), .D(n_36812763), .Z(n_278459028));
	notech_and4 i_174137415(.A(n_278059024), .B(n_277959023), .C(n_277759021
		), .D(n_242158665), .Z(n_278259026));
	notech_ao4 i_173537421(.A(n_55181), .B(n_29035), .C(n_55170), .D(n_56739
		), .Z(n_278059024));
	notech_nand3 i_2120960(.A(n_321179601), .B(n_321079600), .C(n_320979599)
		, .Z(n_9099));
	notech_nand3 i_1920958(.A(n_321879608), .B(n_321779607), .C(n_321679606)
		, .Z(n_9087));
	notech_or4 i_2221057(.A(n_304775886), .B(n_316679556), .C(n_322379613), 
		.D(n_26451), .Z(n_13941));
	notech_or4 i_2121056(.A(n_320179591), .B(n_315879548), .C(n_323079620), 
		.D(n_26452), .Z(n_13935));
	notech_or4 i_2021055(.A(n_306575904), .B(n_315079540), .C(n_323779627), 
		.D(n_26453), .Z(n_13929));
	notech_or4 i_1921054(.A(n_320579595), .B(n_314279532), .C(n_324479634), 
		.D(n_26454), .Z(n_13923));
	notech_nand3 i_2321314(.A(n_325379643), .B(n_325279642), .C(n_325179641)
		, .Z(n_20733));
	notech_nand3 i_2221313(.A(n_326079650), .B(n_325979649), .C(n_325879648)
		, .Z(n_20727));
	notech_nand2 i_2321570(.A(n_327179661), .B(n_326679656), .Z(n_16482));
	notech_nand2 i_2221569(.A(n_328179671), .B(n_327679666), .Z(n_16476));
	notech_nand2 i_2121568(.A(n_329179681), .B(n_328679676), .Z(n_16470));
	notech_nand2 i_2021567(.A(n_330179691), .B(n_329679686), .Z(n_16464));
	notech_nand2 i_1921566(.A(n_331179701), .B(n_330679696), .Z(n_16458));
	notech_or4 i_2221601(.A(n_304775886), .B(n_305679446), .C(n_331579705), 
		.D(n_26455), .Z(n_13241));
	notech_or4 i_2121600(.A(n_320179591), .B(n_304879438), .C(n_332279712), 
		.D(n_26456), .Z(n_13235));
	notech_or4 i_2021599(.A(n_306575904), .B(n_304079430), .C(n_332979719), 
		.D(n_26457), .Z(n_13229));
	notech_or4 i_1921598(.A(n_320579595), .B(n_303279422), .C(n_333679726), 
		.D(n_26458), .Z(n_13223));
	notech_nand2 i_2321730(.A(n_335079740), .B(n_334579735), .Z(n_12899));
	notech_nand2 i_2221729(.A(n_336379751), .B(n_335679746), .Z(n_12893));
	notech_nand2 i_2121728(.A(n_337479762), .B(n_336979757), .Z(n_12887));
	notech_nand2 i_2021727(.A(n_340979773), .B(n_338079768), .Z(n_12881));
	notech_nand2 i_1921726(.A(n_342079784), .B(n_341579779), .Z(n_12875));
	notech_and4 i_2221857(.A(n_342179785), .B(n_342679787), .C(n_344479792),
		 .D(n_296679356), .Z(n_12527));
	notech_or4 i_2121856(.A(n_320179591), .B(n_295179341), .C(n_344879796), 
		.D(n_26462), .Z(n_12521));
	notech_and4 i_2021855(.A(n_345279800), .B(n_345479802), .C(n_345979807),
		 .D(n_295079340), .Z(n_12515));
	notech_and4 i_1921854(.A(n_346079808), .B(n_346279810), .C(n_346779815),
		 .D(n_294279332), .Z(n_12509));
	notech_nand2 i_2316672(.A(n_347779825), .B(n_347279820), .Z(n_11824));
	notech_nand2 i_2216671(.A(n_348779835), .B(n_348279830), .Z(n_11818));
	notech_and4 i_2116670(.A(n_349379841), .B(n_349579843), .C(n_349279840),
		 .D(n_290679296), .Z(n_11812));
	notech_and4 i_2016669(.A(n_350279850), .B(n_350479852), .C(n_350179849),
		 .D(n_289579285), .Z(n_11806));
	notech_nand2 i_166442234(.A(read_data[18]), .B(n_59936), .Z(n_307918856)
		);
	notech_ao4 i_173437422(.A(n_2156), .B(n_28813), .C(n_55136), .D(n_27577)
		, .Z(n_277959023));
	notech_and4 i_326953(.A(n_1914), .B(n_357579920), .C(n_357979924), .D(n_54784
		), .Z(n_14908));
	notech_ao4 i_173337423(.A(n_55122), .B(n_55261), .C(n_55111), .D(nbus_11326
		[4]), .Z(n_277759021));
	notech_or4 i_151533150(.A(instrc[110]), .B(instrc[111]), .C(n_28562), .D
		(n_28563), .Z(n_54913));
	notech_or4 i_426954(.A(n_26620), .B(n_360779952), .C(n_362479969), .D(n_26232
		), .Z(n_14914));
	notech_nand2 i_3217578(.A(n_363679981), .B(n_363179976), .Z(n_21029));
	notech_or4 i_117547(.A(n_359179936), .B(n_363979984), .C(n_26470), .D(n_364779992
		), .Z(n_20843));
	notech_and2 i_138188455(.A(n_353688272), .B(n_275888699), .Z(n_366088135
		));
	notech_ao4 i_173737419(.A(n_55526), .B(n_28576), .C(n_55102), .D(n_28786
		), .Z(n_277559019));
	notech_ao4 i_173637420(.A(n_55243), .B(n_27531), .C(n_55192), .D(nbus_11326
		[12]), .Z(n_277459018));
	notech_ao4 i_174637410(.A(n_89513289), .B(n_27596), .C(n_88913283), .D(n_28842
		), .Z(n_277359017));
	notech_and4 i_171337443(.A(n_276859012), .B(n_240758653), .C(n_240358649
		), .D(n_240458650), .Z(n_277159015));
	notech_and4 i_170937447(.A(n_275959003), .B(n_275859002), .C(n_276659010
		), .D(n_36812763), .Z(n_276859012));
	notech_and4 i_170737449(.A(n_276459008), .B(n_276359007), .C(n_276159005
		), .D(n_240258648), .Z(n_276659010));
	notech_ao4 i_170137455(.A(n_55181), .B(n_29027), .C(n_55170), .D(n_56748
		), .Z(n_276459008));
	notech_ao4 i_170037456(.A(n_55161), .B(n_28814), .C(n_55136), .D(n_27578
		), .Z(n_276359007));
	notech_ao4 i_169937457(.A(n_55122), .B(n_55249), .C(n_55111), .D(nbus_11326
		[5]), .Z(n_276159005));
	notech_ao4 i_170337453(.A(n_55526), .B(n_28573), .C(n_55102), .D(n_28787
		), .Z(n_275959003));
	notech_ao4 i_170237454(.A(n_55243), .B(n_27532), .C(n_55192), .D(nbus_11326
		[13]), .Z(n_275859002));
	notech_ao4 i_171237444(.A(n_89513289), .B(n_27597), .C(n_88913283), .D(n_28843
		), .Z(n_275759001));
	notech_nand3 i_3939053(.A(n_56060), .B(n_238758633), .C(n_323388457), .Z
		(n_107113465));
	notech_ao4 i_60938499(.A(n_2262), .B(n_27799), .C(n_57373), .D(n_27383),
		 .Z(n_275258996));
	notech_ao4 i_60838500(.A(n_59224), .B(n_28032), .C(n_56270), .D(n_27696)
		, .Z(n_275158995));
	notech_and2 i_61238496(.A(n_274958993), .B(n_274858992), .Z(n_275058994)
		);
	notech_ao4 i_60738501(.A(n_56186), .B(n_27863), .C(n_56290), .D(n_27655)
		, .Z(n_274958993));
	notech_ao4 i_60638502(.A(n_60484), .B(n_27900), .C(n_56183), .D(n_29099)
		, .Z(n_274858992));
	notech_and4 i_61438494(.A(n_274558989), .B(n_274458988), .C(n_274258986)
		, .D(n_274158985), .Z(n_274758991));
	notech_ao4 i_60538503(.A(n_56182), .B(n_27932), .C(n_56310), .D(n_27619)
		, .Z(n_274558989));
	notech_ao4 i_60438504(.A(n_56415), .B(n_27966), .C(n_57343), .D(n_27761)
		, .Z(n_274458988));
	notech_ao4 i_60338505(.A(n_56226), .B(n_27998), .C(n_197114365), .D(n_27831
		), .Z(n_274258986));
	notech_ao4 i_60138506(.A(n_56240), .B(n_27728), .C(n_2261), .D(n_29100),
		 .Z(n_274158985));
	notech_ao4 i_57738530(.A(n_2262), .B(n_27798), .C(n_57373), .D(n_27382),
		 .Z(n_273858982));
	notech_ao4 i_57638531(.A(n_59224), .B(n_28031), .C(n_56270), .D(n_27695)
		, .Z(n_273758981));
	notech_and2 i_58038527(.A(n_273558979), .B(n_273458978), .Z(n_273658980)
		);
	notech_ao4 i_57538532(.A(n_56276), .B(n_27862), .C(n_56285), .D(n_27654)
		, .Z(n_273558979));
	notech_ao4 i_57438533(.A(n_60479), .B(n_27899), .C(n_56183), .D(n_29096)
		, .Z(n_273458978));
	notech_and4 i_58238525(.A(n_273158975), .B(n_273058974), .C(n_272858972)
		, .D(n_272758971), .Z(n_273358977));
	notech_ao4 i_57338534(.A(n_56182), .B(n_27931), .C(n_56310), .D(n_27618)
		, .Z(n_273158975));
	notech_ao4 i_57238535(.A(n_56415), .B(n_27965), .C(n_57343), .D(n_27760)
		, .Z(n_273058974));
	notech_ao4 i_57138536(.A(n_56226), .B(n_27997), .C(n_57358), .D(n_27830)
		, .Z(n_272858972));
	notech_ao4 i_57038537(.A(n_56235), .B(n_27727), .C(n_2261), .D(n_29097),
		 .Z(n_272758971));
	notech_ao4 i_54438561(.A(n_56255), .B(n_27797), .C(n_57371), .D(n_27381)
		, .Z(n_272458968));
	notech_ao4 i_54338562(.A(n_59219), .B(n_28030), .C(n_56265), .D(n_27694)
		, .Z(n_272358967));
	notech_and2 i_54738558(.A(n_272158965), .B(n_272058964), .Z(n_272258966)
		);
	notech_ao4 i_54238563(.A(n_56276), .B(n_27861), .C(n_56285), .D(n_27653)
		, .Z(n_272158965));
	notech_ao4 i_54138564(.A(n_60479), .B(n_27898), .C(n_56395), .D(n_29093)
		, .Z(n_272058964));
	notech_and4 i_54938556(.A(n_271758961), .B(n_271658960), .C(n_271458958)
		, .D(n_271358957), .Z(n_271958963));
	notech_ao4 i_54038565(.A(n_56296), .B(n_27930), .C(n_56305), .D(n_27617)
		, .Z(n_271758961));
	notech_ao4 i_53938566(.A(n_56415), .B(n_27964), .C(n_57338), .D(n_27758)
		, .Z(n_271658960));
	notech_ao4 i_53838567(.A(n_56226), .B(n_27996), .C(n_57358), .D(n_27829)
		, .Z(n_271458958));
	notech_ao4 i_53738568(.A(n_56235), .B(n_27726), .C(n_56246), .D(n_29094)
		, .Z(n_271358957));
	notech_ao4 i_51338592(.A(n_56255), .B(n_27796), .C(n_57367), .D(n_27380)
		, .Z(n_271058954));
	notech_ao4 i_51238593(.A(n_59219), .B(n_28029), .C(n_56265), .D(n_27693)
		, .Z(n_270958953));
	notech_and2 i_51638589(.A(n_270758951), .B(n_270658950), .Z(n_270858952)
		);
	notech_ao4 i_51138594(.A(n_56276), .B(n_27860), .C(n_56285), .D(n_27652)
		, .Z(n_270758951));
	notech_ao4 i_51038595(.A(n_60479), .B(n_27897), .C(n_29090), .D(n_56395)
		, .Z(n_270658950));
	notech_and4 i_51838587(.A(n_270358947), .B(n_270258946), .C(n_270058944)
		, .D(n_269958943), .Z(n_270558949));
	notech_ao4 i_50938596(.A(n_56296), .B(n_27929), .C(n_56305), .D(n_27616)
		, .Z(n_270358947));
	notech_ao4 i_50838597(.A(n_56415), .B(n_27963), .C(n_57338), .D(n_27757)
		, .Z(n_270258946));
	notech_ao4 i_50738598(.A(n_56226), .B(n_27995), .C(n_27828), .D(n_57358)
		, .Z(n_270058944));
	notech_ao4 i_50638599(.A(n_56235), .B(n_27725), .C(n_55450), .D(n_56246)
		, .Z(n_269958943));
	notech_ao4 i_48238623(.A(n_56255), .B(n_27794), .C(n_57367), .D(n_27378)
		, .Z(n_269658940));
	notech_ao4 i_48138624(.A(n_59219), .B(n_28027), .C(n_56265), .D(n_27691)
		, .Z(n_269558939));
	notech_and2 i_48538620(.A(n_269358937), .B(n_269258936), .Z(n_269458938)
		);
	notech_ao4 i_48038625(.A(n_56276), .B(n_27858), .C(n_56285), .D(n_27649)
		, .Z(n_269358937));
	notech_ao4 i_47938626(.A(n_60479), .B(n_27895), .C(n_56395), .D(n_29101)
		, .Z(n_269258936));
	notech_and4 i_48738618(.A(n_268958933), .B(n_268858932), .C(n_268658930)
		, .D(n_268558929), .Z(n_269158935));
	notech_ao4 i_47838627(.A(n_56296), .B(n_27927), .C(n_56305), .D(n_27614)
		, .Z(n_268958933));
	notech_ao4 i_47738628(.A(n_56415), .B(n_27961), .C(n_57338), .D(n_27755)
		, .Z(n_268858932));
	notech_ao4 i_47638629(.A(n_27993), .B(n_56226), .C(n_57358), .D(n_27826)
		, .Z(n_268658930));
	notech_ao4 i_47538630(.A(n_56235), .B(n_27723), .C(n_29102), .D(n_56246)
		, .Z(n_268558929));
	notech_ao4 i_45138654(.A(n_56255), .B(n_27792), .C(n_57367), .D(n_27376)
		, .Z(n_268258926));
	notech_ao4 i_45038655(.A(n_59219), .B(n_28025), .C(n_56265), .D(n_27689)
		, .Z(n_268158925));
	notech_and2 i_45438651(.A(n_267958923), .B(n_267858922), .Z(n_268058924)
		);
	notech_ao4 i_44938656(.A(n_56276), .B(n_27856), .C(n_56285), .D(n_27646)
		, .Z(n_267958923));
	notech_ao4 i_44838657(.A(n_60479), .B(n_27893), .C(n_56395), .D(n_29105)
		, .Z(n_267858922));
	notech_and4 i_45638649(.A(n_267558919), .B(n_267458918), .C(n_267258916)
		, .D(n_267158915), .Z(n_267758921));
	notech_ao4 i_44638658(.A(n_56296), .B(n_27925), .C(n_56305), .D(n_27612)
		, .Z(n_267558919));
	notech_ao4 i_44538659(.A(n_56415), .B(n_27959), .C(n_57338), .D(n_27753)
		, .Z(n_267458918));
	notech_ao4 i_44438660(.A(n_56226), .B(n_27991), .C(n_27824), .D(n_57358)
		, .Z(n_267258916));
	notech_ao4 i_44338661(.A(n_56235), .B(n_27721), .C(n_56246), .D(n_29106)
		, .Z(n_267158915));
	notech_ao4 i_41738685(.A(n_56255), .B(n_27791), .C(n_57367), .D(n_27375)
		, .Z(n_266858912));
	notech_ao4 i_41638686(.A(n_59219), .B(n_28024), .C(n_56265), .D(n_27688)
		, .Z(n_266758911));
	notech_and2 i_42038682(.A(n_266558909), .B(n_266458908), .Z(n_266658910)
		);
	notech_ao4 i_41538687(.A(n_56276), .B(n_27855), .C(n_56285), .D(n_27644)
		, .Z(n_266558909));
	notech_ao4 i_41438688(.A(n_60479), .B(n_27891), .C(n_56395), .D(n_29119)
		, .Z(n_266458908));
	notech_and4 i_42238680(.A(n_266158905), .B(n_266058904), .C(n_265858902)
		, .D(n_265758901), .Z(n_266358907));
	notech_ao4 i_41338689(.A(n_56296), .B(n_27924), .C(n_56305), .D(n_27611)
		, .Z(n_266158905));
	notech_ao4 i_41238690(.A(n_56415), .B(n_27958), .C(n_57338), .D(n_27752)
		, .Z(n_266058904));
	notech_ao4 i_41138691(.A(n_56226), .B(n_27990), .C(n_27823), .D(n_57358)
		, .Z(n_265858902));
	notech_ao4 i_41038692(.A(n_56235), .B(n_27720), .C(n_56246), .D(n_29118)
		, .Z(n_265758901));
	notech_ao4 i_38638716(.A(n_56255), .B(n_27790), .C(n_57367), .D(n_27374)
		, .Z(n_265458898));
	notech_ao4 i_38538717(.A(n_59219), .B(n_28023), .C(n_56265), .D(n_27687)
		, .Z(n_265358897));
	notech_and2 i_38938713(.A(n_265158895), .B(n_265058894), .Z(n_265258896)
		);
	notech_ao4 i_38438718(.A(n_56276), .B(n_27854), .C(n_56285), .D(n_27643)
		, .Z(n_265158895));
	notech_ao4 i_38338719(.A(n_60479), .B(n_27889), .C(n_56395), .D(n_29103)
		, .Z(n_265058894));
	notech_and4 i_39138711(.A(n_264758891), .B(n_264658890), .C(n_264458888)
		, .D(n_264358887), .Z(n_264958893));
	notech_ao4 i_38238720(.A(n_56296), .B(n_27923), .C(n_56305), .D(n_27610)
		, .Z(n_264758891));
	notech_ao4 i_38138721(.A(n_56415), .B(n_27957), .C(n_57338), .D(n_27751)
		, .Z(n_264658890));
	notech_ao4 i_38038722(.A(n_56226), .B(n_27989), .C(n_27822), .D(n_57358)
		, .Z(n_264458888));
	notech_ao4 i_37938723(.A(n_56235), .B(n_27719), .C(n_56246), .D(n_29104)
		, .Z(n_264358887));
	notech_ao4 i_34938747(.A(n_56255), .B(n_27789), .C(n_57367), .D(n_27373)
		, .Z(n_264058884));
	notech_ao4 i_34838748(.A(n_59219), .B(n_28022), .C(n_56265), .D(n_27686)
		, .Z(n_263958883));
	notech_and2 i_35238744(.A(n_263758881), .B(n_263658880), .Z(n_263858882)
		);
	notech_ao4 i_34638749(.A(n_56276), .B(n_27853), .C(n_56285), .D(n_27642)
		, .Z(n_263758881));
	notech_ao4 i_34538750(.A(n_60479), .B(n_27888), .C(n_56395), .D(n_29117)
		, .Z(n_263658880));
	notech_and4 i_35538742(.A(n_263358877), .B(n_263258876), .C(n_263058874)
		, .D(n_262958873), .Z(n_263558879));
	notech_ao4 i_34438751(.A(n_56296), .B(n_27922), .C(n_56305), .D(n_27609)
		, .Z(n_263358877));
	notech_ao4 i_34338752(.A(n_56415), .B(n_27956), .C(n_57338), .D(n_27750)
		, .Z(n_263258876));
	notech_ao4 i_34238753(.A(n_56226), .B(n_27988), .C(n_27821), .D(n_57358)
		, .Z(n_263058874));
	notech_ao4 i_34138754(.A(n_56235), .B(n_27718), .C(n_29116), .D(n_56246)
		, .Z(n_262958873));
	notech_ao4 i_32138773(.A(instrc[120]), .B(n_220758481), .C(n_220658480),
		 .D(n_59235), .Z(n_262858872));
	notech_ao4 i_29738797(.A(n_323888452), .B(n_217658456), .C(n_323188459),
		 .D(n_217558455), .Z(n_262558869));
	notech_and2 i_7339020(.A(instrc[123]), .B(instrc[121]), .Z(n_262058864)
		);
	notech_and4 i_116170(.A(n_2976), .B(n_2980), .C(n_298288686), .D(n_260858852
		), .Z(n_14092));
	notech_or2 i_212537037(.A(n_2320), .B(n_2699), .Z(n_260858852));
	notech_or4 i_212637036(.A(n_60780), .B(n_60726), .C(n_2985), .D(n_55356)
		, .Z(n_260758851));
	notech_or2 i_212437038(.A(n_304188646), .B(n_27535), .Z(n_260658850));
	notech_and4 i_9438999(.A(n_55087), .B(n_57338), .C(n_259058834), .D(n_258858832
		), .Z(n_259158835));
	notech_nand2 i_210637056(.A(opz[0]), .B(n_2796), .Z(n_259058834));
	notech_nand2 i_112239156(.A(n_56395), .B(n_56296), .Z(n_258958833));
	notech_nand2 i_210737055(.A(instrc[104]), .B(n_258958833), .Z(n_258858832
		));
	notech_and4 i_316172(.A(n_258758831), .B(n_2942), .C(n_2960), .D(n_256458808
		), .Z(n_14104));
	notech_nao3 i_208137080(.A(imm[34]), .B(n_26795), .C(n_2198), .Z(n_258758831
		));
	notech_nao3 i_207737084(.A(n_57448), .B(nbus_138[2]), .C(n_2318), .Z(n_258458828
		));
	notech_nao3 i_207937082(.A(n_239058636), .B(imm[2]), .C(n_2213), .Z(n_258158825
		));
	notech_and4 i_9339000(.A(n_55087), .B(n_56235), .C(n_256358807), .D(n_256258806
		), .Z(n_256658810));
	notech_or2 i_207637085(.A(n_2320), .B(n_322488466), .Z(n_256458808));
	notech_nand3 i_205737103(.A(opz[2]), .B(n_59230), .C(n_26772), .Z(n_256358807
		));
	notech_nand2 i_205837102(.A(n_57162), .B(n_258958833), .Z(n_256258806)
		);
	notech_and4 i_416173(.A(n_2938), .B(n_2937), .C(n_2935), .D(n_256158805)
		, .Z(n_14110));
	notech_or4 i_203437126(.A(n_55087), .B(n_2213), .C(n_28567), .D(n_26499)
		, .Z(n_256158805));
	notech_nao3 i_203137129(.A(n_239058636), .B(imm[3]), .C(n_2213), .Z(n_255658800
		));
	notech_or2 i_202837132(.A(n_2320), .B(n_322688464), .Z(n_255558799));
	notech_or2 i_6239031(.A(n_2213), .B(n_216258444), .Z(n_255458798));
	notech_nand3 i_516174(.A(n_2918), .B(n_2917), .C(n_2899), .Z(n_14116));
	notech_or4 i_199037169(.A(n_55087), .B(n_2213), .C(n_48760), .D(n_28567)
		, .Z(n_253358777));
	notech_nand3 i_616175(.A(n_289788687), .B(n_2880), .C(n_2896), .Z(n_14122
		));
	notech_nao3 i_194637212(.A(n_239058636), .B(imm[5]), .C(n_2213), .Z(n_251458758
		));
	notech_or2 i_194337215(.A(n_2320), .B(n_322788463), .Z(n_251358757));
	notech_nand3 i_716176(.A(n_287888688), .B(n_2865), .C(n_283759081), .Z(n_14128
		));
	notech_nao3 i_190537252(.A(imm[6]), .B(n_239058636), .C(n_2213), .Z(n_249458738
		));
	notech_or2 i_190237255(.A(n_2320), .B(n_57352), .Z(n_249358737));
	notech_and4 i_91729144(.A(n_268258926), .B(n_268158925), .C(n_267758921)
		, .D(n_268058924), .Z(n_57352));
	notech_nao3 i_188737270(.A(n_56079), .B(n_59230), .C(n_273888717), .Z(n_247858722
		));
	notech_nand3 i_916178(.A(n_283559079), .B(n_282159065), .C(n_246158705),
		 .Z(n_14140));
	notech_nao3 i_186837289(.A(imm[40]), .B(n_26795), .C(n_2198), .Z(n_247758721
		));
	notech_nao3 i_186537292(.A(n_57448), .B(nbus_138[8]), .C(n_2318), .Z(n_247458718
		));
	notech_or2 i_186437293(.A(n_57350), .B(n_2320), .Z(n_247358717));
	notech_nand2 i_186337294(.A(add_src[8]), .B(n_26579), .Z(n_247258716));
	notech_nand2 i_186937288(.A(opb[8]), .B(n_272388732), .Z(n_246158705));
	notech_and4 i_91929145(.A(n_269658940), .B(n_269558939), .C(n_269158935)
		, .D(n_269458938), .Z(n_57350));
	notech_nand3 i_1116180(.A(n_281959063), .B(n_280559049), .C(n_244458688)
		, .Z(n_14152));
	notech_nao3 i_180037357(.A(imm[42]), .B(n_26795), .C(n_2198), .Z(n_246058704
		));
	notech_nao3 i_179737360(.A(n_57448), .B(nbus_138[10]), .C(n_2318), .Z(n_245758701
		));
	notech_or2 i_179637361(.A(n_2320), .B(n_57348), .Z(n_245658700));
	notech_nand2 i_179537362(.A(add_src[10]), .B(n_26579), .Z(n_245558699)
		);
	notech_nand2 i_180137356(.A(n_272388732), .B(opb[10]), .Z(n_244458688)
		);
	notech_and4 i_92129146(.A(n_271058954), .B(n_270958953), .C(n_270558949)
		, .D(n_270858952), .Z(n_57348));
	notech_nand3 i_1216181(.A(n_280359047), .B(n_278959033), .C(n_242758671)
		, .Z(n_14158));
	notech_nao3 i_176537391(.A(imm[43]), .B(n_26795), .C(n_2198), .Z(n_244358687
		));
	notech_nao3 i_176237394(.A(n_57448), .B(nbus_138[11]), .C(n_2318), .Z(n_244058684
		));
	notech_or2 i_176137395(.A(n_2320), .B(n_57347), .Z(n_243958683));
	notech_nand2 i_176037396(.A(add_src[11]), .B(n_26579), .Z(n_243858682)
		);
	notech_nand2 i_176637390(.A(n_272388732), .B(opb[11]), .Z(n_242758671)
		);
	notech_and4 i_92229147(.A(n_272458968), .B(n_272358967), .C(n_271958963)
		, .D(n_272258966), .Z(n_57347));
	notech_nand3 i_1316182(.A(n_278759031), .B(n_277359017), .C(n_240858654)
		, .Z(n_14164));
	notech_nao3 i_173137425(.A(imm[44]), .B(n_26795), .C(n_2198), .Z(n_242658670
		));
	notech_nao3 i_172837428(.A(n_57448), .B(nbus_138[12]), .C(n_2318), .Z(n_242358667
		));
	notech_or2 i_172737429(.A(n_55075), .B(n_57346), .Z(n_242258666));
	notech_nand2 i_172637430(.A(add_src[12]), .B(n_26579), .Z(n_242158665)
		);
	notech_nand2 i_173237424(.A(n_272388732), .B(opb[12]), .Z(n_240858654)
		);
	notech_and4 i_92339143(.A(n_273858982), .B(n_273758981), .C(n_273358977)
		, .D(n_273658980), .Z(n_57346));
	notech_nand3 i_1416183(.A(n_277159015), .B(n_275759001), .C(n_239158637)
		, .Z(n_14170));
	notech_nao3 i_169737459(.A(imm[45]), .B(n_26795), .C(n_2198), .Z(n_240758653
		));
	notech_nao3 i_169437462(.A(n_57448), .B(nbus_138[13]), .C(n_2318), .Z(n_240458650
		));
	notech_or2 i_169337463(.A(n_55075), .B(n_57345), .Z(n_240358649));
	notech_nand2 i_169237464(.A(add_src[13]), .B(n_26579), .Z(n_240258648)
		);
	notech_nand2 i_169837458(.A(n_272388732), .B(opb[13]), .Z(n_239158637)
		);
	notech_and4 i_92429148(.A(n_275258996), .B(n_275158995), .C(n_274758991)
		, .D(n_275058994), .Z(n_57345));
	notech_nand3 i_72138393(.A(n_56276), .B(n_56265), .C(n_56285), .Z(n_239058636
		));
	notech_or2 i_65938453(.A(n_55852), .B(n_26576), .Z(n_238958635));
	notech_or2 i_64538466(.A(n_56063), .B(n_26576), .Z(n_238758633));
	notech_and4 i_31838776(.A(instrc[120]), .B(regs_11[2]), .C(n_59230), .D(n_262058864
		), .Z(n_221158484));
	notech_or2 i_31738777(.A(n_60525), .B(n_220958482), .Z(n_221058483));
	notech_ao4 i_8939004(.A(n_323888452), .B(n_220558479), .C(n_323188459), 
		.D(n_220358477), .Z(n_220958482));
	notech_and3 i_9039003(.A(n_219658471), .B(n_219458470), .C(n_218958467),
		 .Z(n_220758481));
	notech_and2 i_9139002(.A(n_262558869), .B(n_217758457), .Z(n_220658480)
		);
	notech_mux2 i_6639027(.S(instrc[120]), .A(n_27641), .B(n_29115), .Z(n_220558479
		));
	notech_mux2 i_6439029(.S(instrc[121]), .A(n_27372), .B(n_27749), .Z(n_220358477
		));
	notech_nao3 i_30638788(.A(instrc[121]), .B(n_219258469), .C(instrc[123])
		, .Z(n_219658471));
	notech_nao3 i_30438790(.A(n_218858466), .B(n_28567), .C(instrc[123]), .Z
		(n_219458470));
	notech_mux2 i_5839035(.S(n_60525), .A(regs_2[2]), .B(regs_6[2]), .Z(n_219258469
		));
	notech_mux2 i_5939034(.S(n_60525), .A(regs_10[2]), .B(regs_14[2]), .Z(n_219158468
		));
	notech_nand3 i_30538789(.A(instrc[123]), .B(instrc[121]), .C(n_219158468
		), .Z(n_218958467));
	notech_mux2 i_6339030(.S(n_60525), .A(regs_0[2]), .B(regs_4[2]), .Z(n_218858466
		));
	notech_nand3 i_29538799(.A(instrc[120]), .B(n_262058864), .C(\eflags[2] 
		), .Z(n_217758457));
	notech_mux2 i_6739026(.S(instrc[120]), .A(n_27608), .B(n_27987), .Z(n_217658456
		));
	notech_mux2 i_6539028(.S(instrc[121]), .A(n_27717), .B(n_28021), .Z(n_217558455
		));
	notech_or4 i_7537(.A(n_59259), .B(n_59268), .C(n_59277), .D(n_2239), .Z(n_217058450
		));
	notech_or2 i_110752073(.A(n_317688513), .B(n_54938), .Z(n_55265));
	notech_or2 i_111552072(.A(n_317688513), .B(n_320888481), .Z(n_55257));
	notech_nand3 i_24238852(.A(n_62433), .B(n_59380), .C(n_56100), .Z(n_216758448
		));
	notech_ao4 i_8839005(.A(n_59380), .B(n_62415), .C(n_2264), .D(n_26251), 
		.Z(n_216658447));
	notech_and2 i_24338851(.A(n_56276), .B(n_26557), .Z(n_216558446));
	notech_ao3 i_4639046(.A(n_55667), .B(n_238958635), .C(n_107113465), .Z(n_216358445
		));
	notech_and3 i_4239050(.A(n_56305), .B(n_1934), .C(n_247858722), .Z(n_216258444
		));
	notech_and3 i_5039042(.A(n_320588484), .B(n_55825), .C(n_317688513), .Z(n_216158443
		));
	notech_or4 i_66052087(.A(n_59259), .B(n_59268), .C(n_59281), .D(n_2241),
		 .Z(n_55690));
	notech_ao4 i_202143412(.A(n_60579), .B(n_55667), .C(n_303321920), .D(n_26500
		), .Z(n_215958441));
	notech_and3 i_246645371(.A(n_54900), .B(n_215958441), .C(n_54851), .Z(n_215558439
		));
	notech_nao3 i_194247315(.A(n_215058434), .B(n_209958385), .C(n_209858384
		), .Z(n_215258436));
	notech_and3 i_194047317(.A(n_214158426), .B(n_214058425), .C(n_214958433
		), .Z(n_215058434));
	notech_and4 i_193947318(.A(n_214758431), .B(n_214658430), .C(n_209758383
		), .D(n_214358428), .Z(n_214958433));
	notech_ao4 i_193347324(.A(n_231547139), .B(n_59023), .C(n_55009), .D(n_28052
		), .Z(n_214758431));
	notech_ao4 i_193247325(.A(n_2311), .B(n_29113), .C(n_2246), .D(n_27537),
		 .Z(n_214658430));
	notech_and3 i_193147326(.A(n_57312), .B(n_2186), .C(n_208858374), .Z(n_214358428
		));
	notech_ao4 i_193547322(.A(n_2248), .B(nbus_11348[1]), .C(n_2247), .D(n_29114
		), .Z(n_214158426));
	notech_ao4 i_193447323(.A(n_2313), .B(n_28902), .C(n_2314), .D(n_59753),
		 .Z(n_214058425));
	notech_nand2 i_184047415(.A(n_57430), .B(rep_en1), .Z(n_213758422));
	notech_nor2 i_203049154(.A(rep_en2), .B(n_213358418), .Z(n_213458419));
	notech_nand3 i_201649155(.A(n_57430), .B(n_26889), .C(n_26596), .Z(n_213358418
		));
	notech_and4 i_129247940(.A(n_212258407), .B(n_212158406), .C(n_212758412
		), .D(n_207958365), .Z(n_212958414));
	notech_and4 i_129047942(.A(n_54860), .B(n_212458409), .C(n_207858364), .D
		(n_207158357), .Z(n_212758412));
	notech_ao4 i_128747945(.A(n_318388506), .B(n_56901), .C(n_318288507), .D
		(n_55234), .Z(n_212458409));
	notech_ao4 i_128647946(.A(n_28997), .B(n_55459), .C(n_131423301), .D(n_27599
		), .Z(n_212258407));
	notech_ao4 i_128547947(.A(n_170914103), .B(n_27553), .C(n_131123298), .D
		(n_59050), .Z(n_212158406));
	notech_and3 i_124947983(.A(n_211758402), .B(n_211658401), .C(n_211558400
		), .Z(n_211958404));
	notech_ao4 i_124247989(.A(n_55933), .B(n_55234), .C(n_55192), .D(n_59050
		), .Z(n_211758402));
	notech_ao4 i_124147990(.A(n_2318), .B(n_28854), .C(n_55619), .D(n_28641)
		, .Z(n_211658401));
	notech_ao3 i_124547986(.A(n_2187), .B(n_211458399), .C(n_206058346), .Z(n_211558400
		));
	notech_ao4 i_124047991(.A(n_55526), .B(n_28572), .C(n_55102), .D(n_28799
		), .Z(n_211458399));
	notech_ao4 i_124447987(.A(n_55181), .B(n_28971), .C(n_55170), .D(n_56901
		), .Z(n_211158396));
	notech_ao4 i_124347988(.A(n_55136), .B(n_27599), .C(n_55243), .D(n_27553
		), .Z(n_211058395));
	notech_and4 i_55548634(.A(n_210358389), .B(n_210258388), .C(n_205558341)
		, .D(n_205658342), .Z(n_210758392));
	notech_ao4 i_55248637(.A(n_97522962), .B(n_58951), .C(n_55403), .D(n_28996
		), .Z(n_210358389));
	notech_ao4 i_55048638(.A(n_322088470), .B(n_56943), .C(n_121623203), .D(n_59095
		), .Z(n_210258388));
	notech_or4 i_216811(.A(n_210158387), .B(n_210058386), .C(n_215258436), .D
		(n_208558371), .Z(n_9712));
	notech_ao4 i_192847329(.A(n_208258368), .B(n_26560), .C(n_110723094), .D
		(n_26421), .Z(n_210158387));
	notech_ao3 i_192947328(.A(opc[0]), .B(nbus_11326[1]), .C(n_21822205), .Z
		(n_210058386));
	notech_nand3 i_192547332(.A(rep_en3), .B(n_213458419), .C(n_4726), .Z(n_209958385
		));
	notech_and4 i_192647331(.A(n_57430), .B(rep_en1), .C(\opc_1[1] ), .D(n_26596
		), .Z(n_209858384));
	notech_nao3 i_192447333(.A(mul64[33]), .B(n_59795), .C(n_55389), .Z(n_209758383
		));
	notech_or2 i_191547342(.A(n_55111), .B(n_55425), .Z(n_208858374));
	notech_nand3 i_3349128(.A(n_55122), .B(n_321988471), .C(n_208458370), .Z
		(n_208658372));
	notech_and2 i_192747330(.A(opc[1]), .B(n_208658372), .Z(n_208558371));
	notech_or2 i_191347344(.A(n_59113), .B(n_21822205), .Z(n_208458370));
	notech_or4 i_184347412(.A(rep_en2), .B(n_213358418), .C(rep_en3), .D(rep_en4
		), .Z(n_208358369));
	notech_and4 i_184247413(.A(n_57430), .B(rep_en2), .C(n_26596), .D(n_26889
		), .Z(n_208258368));
	notech_and4 i_3116680(.A(n_212958414), .B(n_208158367), .C(n_208058366),
		 .D(n_82622813), .Z(n_11872));
	notech_or4 i_128147951(.A(n_57367), .B(n_183258118), .C(n_270988746), .D
		(n_215558439), .Z(n_208158367));
	notech_or2 i_128247950(.A(n_271188744), .B(n_302221909), .Z(n_208058366)
		);
	notech_nao3 i_128347949(.A(opc_10[30]), .B(n_62415), .C(n_302421911), .Z
		(n_207958365));
	notech_nand2 i_128047952(.A(sav_ecx[30]), .B(n_60583), .Z(n_207858364)
		);
	notech_nand3 i_127347959(.A(\regs_1_0[30] ), .B(n_26554), .C(n_59771), .Z
		(n_207158357));
	notech_and4 i_3116200(.A(n_211158396), .B(n_211058395), .C(n_211958404),
		 .D(n_205958345), .Z(n_14272));
	notech_and3 i_122548004(.A(n_2219), .B(resb_shift4box[30]), .C(n_274788710
		), .Z(n_206058346));
	notech_or2 i_123847993(.A(n_55075), .B(n_270988746), .Z(n_205958345));
	notech_or4 i_3220971(.A(n_102723014), .B(n_205758343), .C(n_205858344), 
		.D(n_26602), .Z(n_9165));
	notech_nor2 i_54548642(.A(n_55402), .B(n_271088745), .Z(n_205858344));
	notech_nor2 i_54748641(.A(n_121523202), .B(n_271288743), .Z(n_205758343)
		);
	notech_nao3 i_54848640(.A(opc_10[31]), .B(n_62415), .C(n_121723204), .Z(n_205658342
		));
	notech_or4 i_54948639(.A(n_56172), .B(n_56074), .C(n_56369), .D(n_27601)
		, .Z(n_205558341));
	notech_and4 i_148950566(.A(n_204358329), .B(n_195258238), .C(n_195058236
		), .D(n_204658332), .Z(n_204858334));
	notech_and3 i_148750568(.A(n_16825881), .B(n_194958235), .C(n_195158237)
		, .Z(n_204658332));
	notech_and4 i_148250571(.A(n_204058326), .B(n_194658232), .C(n_194758233
		), .D(n_194858234), .Z(n_204358329));
	notech_ao4 i_147950574(.A(n_59172), .B(n_26632), .C(n_27519), .D(n_170914103
		), .Z(n_204058326));
	notech_nand3 i_146050593(.A(n_203558321), .B(n_203458320), .C(n_193858224
		), .Z(n_203758323));
	notech_ao4 i_145450599(.A(n_131123298), .B(n_58978), .C(n_55131), .D(n_29112
		), .Z(n_203558321));
	notech_ao4 i_145750596(.A(n_131423301), .B(n_27583), .C(n_170914103), .D
		(n_27537), .Z(n_203458320));
	notech_nand2 i_145950594(.A(n_203258318), .B(n_203158317), .Z(n_203358319
		));
	notech_ao4 i_145650597(.A(n_321388476), .B(n_28987), .C(n_321288477), .D
		(n_2700), .Z(n_203258318));
	notech_ao4 i_145550598(.A(n_55533), .B(n_55600), .C(n_55534), .D(n_56784
		), .Z(n_203158317));
	notech_nand3 i_124350792(.A(n_202658312), .B(n_192658212), .C(n_202158307
		), .Z(n_202858314));
	notech_and4 i_124050794(.A(n_202358309), .B(n_192458210), .C(n_202258308
		), .D(n_192058206), .Z(n_202658312));
	notech_ao4 i_123450800(.A(n_59172), .B(n_26716), .C(n_59163), .D(n_27519
		), .Z(n_202358309));
	notech_ao4 i_123750797(.A(n_320188488), .B(n_43626149), .C(n_54024), .D(n_29111
		), .Z(n_202258308));
	notech_and3 i_123950795(.A(n_16825881), .B(n_192158207), .C(n_192558211)
		, .Z(n_202158307));
	notech_and2 i_69951983(.A(n_201958305), .B(n_191558201), .Z(n_16825881)
		);
	notech_ao4 i_122150813(.A(n_2693), .B(n_60474), .C(n_316788522), .D(n_2699
		), .Z(n_201958305));
	notech_ao4 i_113250895(.A(n_43626149), .B(n_261136766), .C(n_2688), .D(n_5577
		), .Z(n_201858304));
	notech_and4 i_113050897(.A(n_201358299), .B(n_201258298), .C(n_191158197
		), .D(n_201158297), .Z(n_201658302));
	notech_ao4 i_112350904(.A(n_53993), .B(n_29110), .C(n_262236777), .D(n_29109
		), .Z(n_201358299));
	notech_ao4 i_112650901(.A(n_59163), .B(n_27519), .C(n_55951), .D(n_55342
		), .Z(n_201258298));
	notech_and2 i_112850899(.A(n_201058296), .B(n_200958295), .Z(n_201158297
		));
	notech_ao4 i_112550902(.A(n_55304), .B(n_55356), .C(n_55316), .D(n_58960
		), .Z(n_201058296));
	notech_ao4 i_112450903(.A(n_55421), .B(n_28986), .C(n_55422), .D(n_2699)
		, .Z(n_200958295));
	notech_and4 i_70851301(.A(n_189758183), .B(n_189658182), .C(n_200458290)
		, .D(n_190058186), .Z(n_200758293));
	notech_and3 i_70451305(.A(n_200258288), .B(n_200158287), .C(n_189558181)
		, .Z(n_200458290));
	notech_ao4 i_70151308(.A(n_58922), .B(n_29108), .C(n_55492), .D(n_27523)
		, .Z(n_200258288));
	notech_ao4 i_70251307(.A(n_321188478), .B(n_55216), .C(n_55236), .D(n_29063
		), .Z(n_200158287));
	notech_ao4 i_70751302(.A(n_2691), .B(n_55365), .C(n_2690), .D(n_58548), 
		.Z(n_200058286));
	notech_ao4 i_70951300(.A(n_316388526), .B(n_55426267), .C(n_319588494), 
		.D(n_55687), .Z(n_199958285));
	notech_and4 i_65651347(.A(n_188558171), .B(n_188458170), .C(n_199458280)
		, .D(n_188858174), .Z(n_199758283));
	notech_and3 i_65151351(.A(n_199258278), .B(n_199158277), .C(n_188358169)
		, .Z(n_199458280));
	notech_ao4 i_64851354(.A(n_58922), .B(n_29107), .C(n_55492), .D(n_27525)
		, .Z(n_199258278));
	notech_ao4 i_64951353(.A(n_57352), .B(n_55216), .C(n_55236), .D(n_29068)
		, .Z(n_199158277));
	notech_ao4 i_65551348(.A(n_2691), .B(n_55387), .C(n_2690), .D(n_27568), 
		.Z(n_199058276));
	notech_ao4 i_65751346(.A(n_316488525), .B(n_55426267), .C(n_57320), .D(n_55687
		), .Z(n_198958275));
	notech_nao3 i_120251974(.A(n_56458), .B(n_195658242), .C(n_187858164), .Z
		(n_198858274));
	notech_nao3 i_33422(.A(n_56460), .B(n_195658242), .C(n_317688513), .Z(n_198758273
		));
	notech_ao4 i_48351505(.A(n_58483), .B(n_28025), .C(n_55873), .D(n_29106)
		, .Z(n_198358269));
	notech_ao4 i_48251506(.A(n_55965), .B(n_27991), .C(n_55992), .D(n_27959)
		, .Z(n_198258268));
	notech_and2 i_48651502(.A(n_198058266), .B(n_197958265), .Z(n_198158267)
		);
	notech_ao4 i_48151507(.A(n_56009), .B(n_27925), .C(n_56023), .D(n_27893)
		, .Z(n_198058266));
	notech_ao4 i_48051508(.A(n_56043), .B(n_27856), .C(n_55866), .D(n_27824)
		, .Z(n_197958265));
	notech_and4 i_48851500(.A(n_197658262), .B(n_197558261), .C(n_197358259)
		, .D(n_197258258), .Z(n_197858264));
	notech_ao4 i_47951509(.A(n_55940), .B(n_27792), .C(n_55888), .D(n_27753)
		, .Z(n_197658262));
	notech_ao4 i_47851510(.A(n_55906), .B(n_27721), .C(n_55924), .D(n_27376)
		, .Z(n_197558261));
	notech_ao4 i_47751511(.A(n_56092), .B(n_27689), .C(n_56126), .D(n_27646)
		, .Z(n_197358259));
	notech_ao4 i_47651512(.A(n_56139), .B(n_27612), .C(n_56382), .D(n_29105)
		, .Z(n_197258258));
	notech_ao4 i_41451573(.A(n_58483), .B(n_28023), .C(n_55873), .D(n_29104)
		, .Z(n_196958255));
	notech_ao4 i_41351574(.A(n_55965), .B(n_27989), .C(n_55992), .D(n_27957)
		, .Z(n_196858254));
	notech_and2 i_41751570(.A(n_196658252), .B(n_196558251), .Z(n_196758253)
		);
	notech_ao4 i_41251575(.A(n_56009), .B(n_27923), .C(n_56023), .D(n_27889)
		, .Z(n_196658252));
	notech_ao4 i_41151576(.A(n_56043), .B(n_27854), .C(n_55866), .D(n_27822)
		, .Z(n_196558251));
	notech_and4 i_41951568(.A(n_196258248), .B(n_196158247), .C(n_195958245)
		, .D(n_195858244), .Z(n_196458250));
	notech_ao4 i_41051577(.A(n_55934), .B(n_27790), .C(n_55888), .D(n_27751)
		, .Z(n_196258248));
	notech_ao4 i_40951578(.A(n_55906), .B(n_27719), .C(n_55919), .D(n_27374)
		, .Z(n_196158247));
	notech_ao4 i_40851579(.A(n_56092), .B(n_27687), .C(n_56126), .D(n_27643)
		, .Z(n_195958245));
	notech_ao4 i_40751580(.A(n_56139), .B(n_27610), .C(n_56382), .D(n_29103)
		, .Z(n_195858244));
	notech_nor2 i_16551808(.A(n_114626850), .B(n_56487), .Z(n_195658242));
	notech_or4 i_116650(.A(n_195358239), .B(n_195458240), .C(n_194158227), .D
		(n_26603), .Z(n_11692));
	notech_nor2 i_147150582(.A(n_194058226), .B(n_55356), .Z(n_195458240));
	notech_nor2 i_146950584(.A(n_55265), .B(n_28986), .Z(n_195358239));
	notech_or2 i_147050583(.A(n_2699), .B(n_55257), .Z(n_195258238));
	notech_or4 i_147650577(.A(n_56574), .B(n_56354), .C(n_55919), .D(n_2688)
		, .Z(n_195158237));
	notech_nao3 i_147850575(.A(n_62427), .B(n_59113), .C(n_198858274), .Z(n_195058236
		));
	notech_nao3 i_147750576(.A(opc_10[0]), .B(n_62415), .C(n_198758273), .Z(n_194958235
		));
	notech_or2 i_147450579(.A(n_194358229), .B(n_55342), .Z(n_194858234));
	notech_nao3 i_147550578(.A(n_4675), .B(n_60138), .C(n_58496), .Z(n_194758233
		));
	notech_nao3 i_147350580(.A(\regs_1[0] ), .B(n_28140), .C(n_58496), .Z(n_194658232
		));
	notech_and3 i_61452051(.A(n_131423301), .B(n_317188518), .C(n_217058450)
		, .Z(n_194358229));
	notech_and3 i_84852052(.A(n_318788502), .B(n_317988510), .C(n_318388506)
		, .Z(n_194258228));
	notech_nor2 i_147250581(.A(n_194258228), .B(n_58960), .Z(n_194158227));
	notech_and3 i_84952053(.A(n_318688503), .B(n_318088509), .C(n_318288507)
		, .Z(n_194058226));
	notech_or4 i_1816667(.A(n_203758323), .B(n_203358319), .C(n_193958225), 
		.D(n_192958215), .Z(n_11794));
	notech_ao3 i_145350600(.A(opc_10[17]), .B(n_62415), .C(n_321588475), .Z(n_193958225
		));
	notech_nand2 i_145150602(.A(sav_ecx[17]), .B(n_60583), .Z(n_193858224)
		);
	notech_nor2 i_145250601(.A(n_3214), .B(n_2648), .Z(n_192958215));
	notech_or4 i_121548(.A(n_192758213), .B(n_202858314), .C(n_192858214), .D
		(n_191858204), .Z(n_16350));
	notech_nor2 i_122450810(.A(n_318888501), .B(n_55356), .Z(n_192858214));
	notech_nor2 i_123050804(.A(n_55222), .B(n_28986), .Z(n_192758213));
	notech_or4 i_122950805(.A(n_182758113), .B(n_56265), .C(n_317788512), .D
		(n_2699), .Z(n_192658212));
	notech_nao3 i_123350801(.A(n_62423), .B(n_59113), .C(n_320688483), .Z(n_192558211
		));
	notech_or4 i_123150803(.A(n_56569), .B(n_56354), .C(n_56092), .D(n_2688)
		, .Z(n_192458210));
	notech_nao3 i_122750807(.A(n_3347), .B(n_55460), .C(n_54046), .Z(n_192158207
		));
	notech_or2 i_122650808(.A(n_319288497), .B(n_27561), .Z(n_192058206));
	notech_nor2 i_122550809(.A(n_319088499), .B(n_58960), .Z(n_191858204));
	notech_or2 i_121950815(.A(n_316688523), .B(n_58960), .Z(n_191558201));
	notech_nao3 i_121164(.A(n_201858304), .B(n_201658302), .C(n_191258198), 
		.Z(n_13467));
	notech_ao3 i_112150906(.A(n_62427), .B(n_59113), .C(n_260436759), .Z(n_191258198
		));
	notech_nand2 i_111950908(.A(sav_edi[0]), .B(n_60583), .Z(n_191158197));
	notech_nand3 i_520624(.A(n_200058286), .B(n_199958285), .C(n_200758293),
		 .Z(n_20135));
	notech_nand2 i_69751311(.A(opa[4]), .B(n_2692), .Z(n_190058186));
	notech_nao3 i_70051309(.A(opc_10[4]), .B(n_62415), .C(n_54526258), .Z(n_189758183
		));
	notech_nand2 i_69451314(.A(n_319688493), .B(n_55819), .Z(n_189658182));
	notech_nand2 i_69251316(.A(sav_epc[4]), .B(n_60583), .Z(n_189558181));
	notech_nand3 i_720626(.A(n_199058276), .B(n_198958275), .C(n_199758283),
		 .Z(n_20147));
	notech_nand2 i_64551357(.A(n_2692), .B(opa[6]), .Z(n_188858174));
	notech_nao3 i_64751355(.A(opc_10[6]), .B(n_62415), .C(n_54526258), .Z(n_188558171
		));
	notech_nand2 i_64251360(.A(n_319788492), .B(n_55819), .Z(n_188458170));
	notech_nand2 i_64051362(.A(sav_epc[6]), .B(n_60583), .Z(n_188358169));
	notech_and4 i_142952030(.A(n_198358269), .B(n_198258268), .C(n_197858264
		), .D(n_198158267), .Z(n_57320));
	notech_and3 i_55351441(.A(n_320588484), .B(n_55825), .C(n_316988520), .Z
		(n_187858164));
	notech_and3 i_54951445(.A(n_316888521), .B(n_319388496), .C(n_55829), .Z
		(n_187758163));
	notech_or4 i_176352014(.A(n_60780), .B(n_60719), .C(n_183958125), .D(n_60579
		), .Z(n_54707));
	notech_ao4 i_25451723(.A(n_272688729), .B(n_274988708), .C(n_273288723),
		 .D(n_2251), .Z(n_183958125));
	notech_ao4 i_52452005(.A(n_204988864), .B(n_56104), .C(n_56345), .D(n_26500
		), .Z(n_55825));
	notech_and3 i_148552066(.A(n_56260), .B(n_183358119), .C(n_183158117), .Z
		(n_54938));
	notech_nao3 i_16751806(.A(n_62429), .B(n_59380), .C(n_321088479), .Z(n_183358119
		));
	notech_ao4 i_83951982(.A(n_59380), .B(n_62401), .C(n_2264), .D(n_321088479
		), .Z(n_183258118));
	notech_nand2 i_16851805(.A(n_57367), .B(n_26562), .Z(n_183158117));
	notech_nand3 i_15551818(.A(n_62433), .B(n_59380), .C(n_320988480), .Z(n_182858114
		));
	notech_ao4 i_84451980(.A(n_59380), .B(n_62419), .C(n_2264), .D(n_26561),
		 .Z(n_182758113));
	notech_nand2 i_15651817(.A(n_56265), .B(n_26563), .Z(n_182658112));
	notech_and3 i_127354073(.A(n_176558053), .B(n_176458052), .C(n_54860), .Z
		(n_182158107));
	notech_ao4 i_127454072(.A(n_318488505), .B(n_29079), .C(n_318588504), .D
		(n_29078), .Z(n_181758104));
	notech_ao4 i_127554071(.A(n_317988510), .B(n_29077), .C(n_57348), .D(n_318088509
		), .Z(n_181658103));
	notech_and4 i_128454062(.A(n_181358100), .B(n_181258099), .C(n_181058097
		), .D(n_180958096), .Z(n_181558102));
	notech_ao4 i_127854068(.A(n_55500), .B(n_55438), .C(n_55501), .D(n_56721
		), .Z(n_181358100));
	notech_ao4 i_127954067(.A(n_55739), .B(n_27575), .C(n_170914103), .D(n_27529
		), .Z(n_181258099));
	notech_ao4 i_128154065(.A(n_59172), .B(n_26644), .C(n_317188518), .D(n_322131608
		), .Z(n_181058097));
	notech_ao4 i_128254064(.A(n_174358031), .B(n_260936764), .C(n_174258030)
		, .D(n_261036765), .Z(n_180958096));
	notech_and4 i_129054057(.A(n_180658093), .B(n_180458091), .C(n_144857736
		), .D(n_145157739), .Z(n_180858095));
	notech_ao4 i_128654061(.A(n_318588504), .B(n_29081), .C(n_55431), .D(n_29080
		), .Z(n_180658093));
	notech_ao4 i_128854059(.A(n_55317), .B(n_55469), .C(n_55318), .D(nbus_11273
		[11]), .Z(n_180458091));
	notech_and4 i_129654052(.A(n_180158088), .B(n_179858086), .C(n_145457742
		), .D(n_145757745), .Z(n_180358090));
	notech_ao4 i_129154056(.A(n_170914103), .B(n_27530), .C(n_59174), .D(n_26645
		), .Z(n_180158088));
	notech_ao4 i_129354054(.A(n_171758005), .B(n_260936764), .C(n_171658004)
		, .D(n_261036765), .Z(n_179858086));
	notech_and4 i_130154047(.A(n_54860), .B(n_179558083), .C(n_179358081), .D
		(n_146257750), .Z(n_179758085));
	notech_ao4 i_129754051(.A(n_318488505), .B(n_29083), .C(n_318588504), .D
		(n_29082), .Z(n_179558083));
	notech_ao4 i_129954049(.A(n_55430), .B(n_57346), .C(n_55317), .D(n_55542
		), .Z(n_179358081));
	notech_and4 i_130754041(.A(n_179058078), .B(n_178858076), .C(n_178758075
		), .D(n_146557753), .Z(n_179258080));
	notech_ao4 i_130254046(.A(n_55739), .B(n_27577), .C(n_170914103), .D(n_27531
		), .Z(n_179058078));
	notech_ao4 i_130454044(.A(n_59174), .B(n_26647), .C(n_317188518), .D(n_321931606
		), .Z(n_178858076));
	notech_ao4 i_130554043(.A(n_169157979), .B(n_260936764), .C(n_169057978)
		, .D(n_261036765), .Z(n_178758075));
	notech_and4 i_131254036(.A(n_54860), .B(n_178458072), .C(n_178258070), .D
		(n_147457762), .Z(n_178658074));
	notech_ao4 i_130854040(.A(n_318488505), .B(n_29086), .C(n_318588504), .D
		(n_29085), .Z(n_178458072));
	notech_ao4 i_131054038(.A(n_55430), .B(n_57345), .C(n_55317), .D(n_55552
		), .Z(n_178258070));
	notech_and4 i_131854030(.A(n_177958067), .B(n_177758065), .C(n_177658064
		), .D(n_147757765), .Z(n_178158069));
	notech_ao4 i_131354035(.A(n_55739), .B(n_27578), .C(n_59150), .D(n_27532
		), .Z(n_177958067));
	notech_ao4 i_131554033(.A(n_59174), .B(n_26648), .C(n_317188518), .D(n_321831605
		), .Z(n_177758065));
	notech_ao4 i_131654032(.A(n_166557953), .B(n_260936764), .C(n_166457952)
		, .D(n_261036765), .Z(n_177658064));
	notech_and4 i_132354025(.A(n_177358061), .B(n_177158059), .C(n_148457772
		), .D(n_148757775), .Z(n_177558063));
	notech_ao4 i_131954029(.A(n_318588504), .B(n_29088), .C(n_29087), .D(n_55431
		), .Z(n_177358061));
	notech_ao4 i_132154027(.A(n_55317), .B(n_55578), .C(n_55318), .D(n_56766
		), .Z(n_177158059));
	notech_and4 i_132854020(.A(n_176858056), .B(n_176658054), .C(n_149057778
		), .D(n_149357781), .Z(n_177058058));
	notech_ao4 i_132454024(.A(n_59150), .B(n_27534), .C(n_59174), .D(n_26649
		), .Z(n_176858056));
	notech_ao4 i_132654022(.A(n_177164109), .B(n_260936764), .C(n_177264110)
		, .D(n_261036765), .Z(n_176658054));
	notech_ao4 i_2055278(.A(n_55791), .B(n_55438), .C(n_55790), .D(n_56721),
		 .Z(n_176558053));
	notech_ao4 i_1955279(.A(n_55789), .B(n_29077), .C(n_57348), .D(n_55786),
		 .Z(n_176458052));
	notech_and4 i_203753326(.A(n_176158049), .B(n_175958047), .C(n_149657784
		), .D(n_149957787), .Z(n_176358051));
	notech_ao4 i_203353330(.A(n_55264), .B(n_57350), .C(n_354269312), .D(n_55413
		), .Z(n_176158049));
	notech_ao4 i_203553328(.A(n_353969310), .B(n_27571), .C(n_55492), .D(n_27527
		), .Z(n_175958047));
	notech_and4 i_204253321(.A(n_175658044), .B(n_175458042), .C(n_150257790
		), .D(n_150557793), .Z(n_175858046));
	notech_ao4 i_203853325(.A(n_26774), .B(n_59174), .C(n_55693), .D(n_57300
		), .Z(n_175658044));
	notech_ao4 i_204053323(.A(n_161857906), .B(n_354469314), .C(n_161957907)
		, .D(n_354369313), .Z(n_175458042));
	notech_and4 i_204753316(.A(n_175158039), .B(n_174958037), .C(n_150857796
		), .D(n_151157799), .Z(n_175358041));
	notech_ao4 i_204353320(.A(n_55264), .B(n_57348), .C(n_354269312), .D(n_55438
		), .Z(n_175158039));
	notech_ao4 i_204553318(.A(n_353969310), .B(n_27575), .C(n_55492), .D(n_27529
		), .Z(n_174958037));
	notech_and4 i_205253311(.A(n_174658034), .B(n_174458032), .C(n_151457802
		), .D(n_151757805), .Z(n_174858036));
	notech_ao4 i_204853315(.A(n_59174), .B(n_26775), .C(n_26435), .D(n_29089
		), .Z(n_174658034));
	notech_ao4 i_205053313(.A(n_354469314), .B(n_174358031), .C(n_354369313)
		, .D(n_174258030), .Z(n_174458032));
	notech_nand2 i_1655313(.A(n_62433), .B(opc[10]), .Z(n_174358031));
	notech_nand2 i_5655306(.A(opc_10[10]), .B(n_62403), .Z(n_174258030));
	notech_ao4 i_205353310(.A(n_56382), .B(n_29090), .C(n_56139), .D(n_27616
		), .Z(n_173958027));
	notech_ao4 i_205453309(.A(n_56126), .B(n_27652), .C(n_56092), .D(n_27693
		), .Z(n_173858026));
	notech_and2 i_205853305(.A(n_173658024), .B(n_173558023), .Z(n_173758025
		));
	notech_ao4 i_205653307(.A(n_55919), .B(n_27380), .C(n_55906), .D(n_27725
		), .Z(n_173658024));
	notech_ao4 i_205753306(.A(n_55888), .B(n_27757), .C(n_55934), .D(n_27796
		), .Z(n_173558023));
	notech_and4 i_206653297(.A(n_173258020), .B(n_173158019), .C(n_172958017
		), .D(n_172858016), .Z(n_173458022));
	notech_ao4 i_206053303(.A(n_55866), .B(n_27828), .C(n_56043), .D(n_27860
		), .Z(n_173258020));
	notech_ao4 i_206153302(.A(n_56023), .B(n_27897), .C(n_56009), .D(n_27929
		), .Z(n_173158019));
	notech_ao4 i_206353300(.A(n_55992), .B(n_27963), .C(n_55965), .D(n_27995
		), .Z(n_172958017));
	notech_ao4 i_206453299(.A(n_55873), .B(n_55450), .C(n_58483), .D(n_28029
		), .Z(n_172858016));
	notech_and4 i_207153292(.A(n_172558013), .B(n_172358011), .C(n_153657824
		), .D(n_153957827), .Z(n_172758015));
	notech_ao4 i_206753296(.A(n_55264), .B(n_57347), .C(n_354269312), .D(n_55469
		), .Z(n_172558013));
	notech_ao4 i_206953294(.A(n_353969310), .B(n_27576), .C(n_55492), .D(n_27530
		), .Z(n_172358011));
	notech_and4 i_207653287(.A(n_172058008), .B(n_171858006), .C(n_154257830
		), .D(n_154557833), .Z(n_172258010));
	notech_ao4 i_207253291(.A(n_59172), .B(n_26777), .C(n_26435), .D(n_29092
		), .Z(n_172058008));
	notech_ao4 i_207453289(.A(n_354469314), .B(n_171758005), .C(n_354369313)
		, .D(n_171658004), .Z(n_171858006));
	notech_nand2 i_3755311(.A(n_62433), .B(opc[11]), .Z(n_171758005));
	notech_nand2 i_5555307(.A(opc_10[11]), .B(n_62403), .Z(n_171658004));
	notech_ao4 i_207753286(.A(n_56382), .B(n_29093), .C(n_56139), .D(n_27617
		), .Z(n_171358001));
	notech_nand2 i_13170130(.A(imm[1]), .B(n_316783142), .Z(n_109081078));
	notech_and3 i_47285(.A(n_42082), .B(n_206482046), .C(n_54862), .Z(n_9223
		));
	notech_ao4 i_47440(.A(n_271039498), .B(n_117781165), .C(n_29123), .D(n_54892
		), .Z(\nbus_11284[0] ));
	notech_ao4 i_46581(.A(n_107542794), .B(n_366088135), .C(n_271039498), .D
		(n_2781), .Z(\nbus_11275[0] ));
	notech_or4 i_4968225(.A(n_60780), .B(n_60721), .C(n_60579), .D(n_55006),
		 .Z(n_109681084));
	notech_nand3 i_54739(.A(n_55634), .B(n_206841699), .C(n_109681084), .Z(\nbus_11353[8] 
		));
	notech_nao3 i_54735(.A(n_206841699), .B(n_54968), .C(n_132760409), .Z(\nbus_11353[0] 
		));
	notech_ao4 i_46791(.A(n_335262250), .B(n_29123), .C(n_271039498), .D(n_55280
		), .Z(\nbus_11277[0] ));
	notech_ao4 i_52903(.A(n_29123), .B(n_117981167), .C(n_55280), .D(n_271039498
		), .Z(\nbus_11342[0] ));
	notech_or4 i_7668198(.A(n_260988754), .B(n_260888755), .C(n_244656264), 
		.D(n_2826), .Z(n_109981087));
	notech_ao3 i_568269(.A(n_2223), .B(n_109981087), .C(n_58591), .Z(n_110281090
		));
	notech_or2 i_8268192(.A(n_110481092), .B(n_29123), .Z(n_110381091));
	notech_ao4 i_468270(.A(n_59150), .B(n_118081168), .C(n_2205), .D(n_38340
		), .Z(n_110481092));
	notech_nand2 i_55072(.A(n_118381171), .B(n_110381091), .Z(\nbus_11355[16] 
		));
	notech_and2 i_8768187(.A(n_110881096), .B(n_118481172), .Z(n_110781095)
		);
	notech_or4 i_868266(.A(n_26380), .B(n_55771), .C(n_333188381), .D(n_59771
		), .Z(n_110881096));
	notech_ao4 i_47646(.A(n_54813), .B(n_271039498), .C(n_110781095), .D(n_118581173
		), .Z(\nbus_11286[16] ));
	notech_ao4 i_47645(.A(n_55640), .B(n_271039498), .C(n_110781095), .D(n_118581173
		), .Z(\nbus_11286[8] ));
	notech_ao4 i_6327543(.A(n_54513), .B(n_28705), .C(n_54491), .D(n_28707),
		 .Z(n_8622));
	notech_ao4 i_6227542(.A(n_54513), .B(n_28704), .C(n_54491), .D(n_28706),
		 .Z(n_8617));
	notech_ao4 i_6127541(.A(n_54491), .B(n_28705), .C(n_54513), .D(n_28703),
		 .Z(n_8612));
	notech_ao4 i_6027540(.A(n_54513), .B(n_28702), .C(n_54491), .D(n_28704),
		 .Z(n_8607));
	notech_ao4 i_5927539(.A(n_54513), .B(n_28701), .C(n_54492), .D(n_28703),
		 .Z(n_8602));
	notech_ao4 i_5827538(.A(n_54513), .B(n_28700), .C(n_54492), .D(n_28702),
		 .Z(n_8597));
	notech_ao4 i_5727537(.A(n_54513), .B(n_28699), .C(n_54491), .D(n_28701),
		 .Z(n_8592));
	notech_ao4 i_5627536(.A(n_54513), .B(n_28698), .C(n_54491), .D(n_28700),
		 .Z(n_8587));
	notech_ao4 i_5527535(.A(n_54513), .B(n_28697), .C(n_54491), .D(n_28699),
		 .Z(n_8582));
	notech_ao4 i_5427534(.A(n_54513), .B(n_28696), .C(n_54491), .D(n_28698),
		 .Z(n_8577));
	notech_ao4 i_5327533(.A(n_54513), .B(n_28695), .C(n_54491), .D(n_28697),
		 .Z(n_8572));
	notech_ao4 i_5227532(.A(n_54513), .B(n_28694), .C(n_54491), .D(n_28696),
		 .Z(n_8567));
	notech_ao4 i_5127531(.A(n_54513), .B(n_28693), .C(n_54491), .D(n_28695),
		 .Z(n_8562));
	notech_ao4 i_5027530(.A(n_54513), .B(n_28692), .C(n_54491), .D(n_28694),
		 .Z(n_8557));
	notech_ao4 i_4927529(.A(n_54513), .B(n_28691), .C(n_54491), .D(n_28693),
		 .Z(n_8552));
	notech_ao4 i_4827528(.A(n_54513), .B(n_28690), .C(n_54491), .D(n_28692),
		 .Z(n_8547));
	notech_ao4 i_4727527(.A(n_54513), .B(n_28689), .C(n_54492), .D(n_28691),
		 .Z(n_8542));
	notech_ao4 i_4627526(.A(n_54514), .B(n_28688), .C(n_54492), .D(n_28690),
		 .Z(n_8537));
	notech_ao4 i_4527525(.A(n_54514), .B(n_28687), .C(n_54492), .D(n_28689),
		 .Z(n_8532));
	notech_ao4 i_4427524(.A(n_54514), .B(n_28686), .C(n_54492), .D(n_28688),
		 .Z(n_8527));
	notech_ao4 i_4327523(.A(n_54514), .B(n_28685), .C(n_54492), .D(n_28687),
		 .Z(n_8522));
	notech_ao4 i_4227522(.A(n_54514), .B(n_28684), .C(n_54492), .D(n_28686),
		 .Z(n_8517));
	notech_ao4 i_4127521(.A(n_54514), .B(n_28683), .C(n_54492), .D(n_28685),
		 .Z(n_8512));
	notech_ao4 i_4027520(.A(n_54514), .B(n_28682), .C(n_54492), .D(n_28684),
		 .Z(n_8507));
	notech_ao4 i_3927519(.A(n_54514), .B(n_28681), .C(n_54492), .D(n_28683),
		 .Z(n_8502));
	notech_ao4 i_3827518(.A(n_54514), .B(n_28680), .C(n_54492), .D(n_28682),
		 .Z(n_8497));
	notech_ao4 i_3727517(.A(n_54514), .B(n_28679), .C(n_54492), .D(n_28681),
		 .Z(n_8492));
	notech_ao4 i_3627516(.A(n_54514), .B(n_28678), .C(n_54492), .D(n_28680),
		 .Z(n_8487));
	notech_ao4 i_3527515(.A(n_54514), .B(n_28677), .C(n_54492), .D(n_28679),
		 .Z(n_8482));
	notech_ao4 i_3427514(.A(n_54514), .B(n_28676), .C(n_54492), .D(n_28678),
		 .Z(n_8477));
	notech_ao4 i_1268262(.A(n_275788700), .B(n_118681174), .C(n_26496), .D(n_258636741
		), .Z(n_117581163));
	notech_ao4 i_8228(.A(n_117581163), .B(n_275588702), .C(n_60583), .D(n_59935
		), .Z(n_10127));
	notech_nao3 i_2268252(.A(n_2042), .B(n_26785), .C(n_2179), .Z(n_117781165
		));
	notech_or4 i_7468200(.A(n_275088707), .B(n_57451), .C(n_59163), .D(n_29124
		), .Z(n_117981167));
	notech_or4 i_8068194(.A(n_275388704), .B(n_2835), .C(n_29130), .D(n_57444
		), .Z(n_118081168));
	notech_nao3 i_8468190(.A(n_57445), .B(n_26399), .C(n_346288346), .Z(n_118281170
		));
	notech_ao4 i_8568189(.A(n_107542794), .B(n_118281170), .C(n_271039498), 
		.D(n_110281090), .Z(n_118381171));
	notech_ao4 i_8868186(.A(n_55008), .B(n_275088707), .C(n_2157), .D(n_59771
		), .Z(n_118481172));
	notech_nand3 i_8968185(.A(n_59172), .B(n_59935), .C(n_61175), .Z(n_118581173
		));
	notech_nand3 i_147466821(.A(n_349988309), .B(n_349488314), .C(n_26554), 
		.Z(n_118681174));
	notech_and2 i_2765641(.A(n_328083255), .B(n_327783252), .Z(n_118781175)
		);
	notech_ao4 i_2665642(.A(n_328083255), .B(n_328183256), .C(n_325783232), 
		.D(n_27564), .Z(n_118881176));
	notech_or2 i_63965060(.A(n_54492), .B(n_28644), .Z(n_119081178));
	notech_ao4 i_149465670(.A(n_2271), .B(n_59935), .C(opb[31]), .D(n_172781715
		), .Z(n_119181179));
	notech_or2 i_77264928(.A(n_54492), .B(n_28677), .Z(n_119381181));
	notech_ao4 i_2065648(.A(n_119881186), .B(n_29485), .C(n_28569), .D(n_169181679
		), .Z(n_119481182));
	notech_mux2 i_2165647(.S(mul64[15]), .A(n_29486), .B(n_29487), .Z(n_119581183
		));
	notech_ao4 i_2365645(.A(n_272788728), .B(mul64[7]), .C(n_62403), .D(\opcode[3] 
		), .Z(n_119881186));
	notech_ao3 i_85464846(.A(n_26390), .B(imm[31]), .C(n_56114), .Z(n_120381191
		));
	notech_ao3 i_85564845(.A(n_26390), .B(imm[30]), .C(n_56114), .Z(n_120481192
		));
	notech_ao3 i_85664844(.A(n_26390), .B(imm[29]), .C(n_56108), .Z(n_120581193
		));
	notech_ao3 i_85764843(.A(n_26390), .B(imm[28]), .C(n_56108), .Z(n_120681194
		));
	notech_ao3 i_85864842(.A(n_26390), .B(imm[27]), .C(n_56108), .Z(n_120781195
		));
	notech_ao3 i_85964841(.A(n_26390), .B(imm[26]), .C(n_56108), .Z(n_120881196
		));
	notech_ao3 i_86064840(.A(n_26390), .B(imm[25]), .C(n_56108), .Z(n_120981197
		));
	notech_ao3 i_86164839(.A(n_26390), .B(imm[24]), .C(n_56108), .Z(n_121081198
		));
	notech_ao3 i_86264838(.A(n_26390), .B(imm[23]), .C(n_56108), .Z(n_121181199
		));
	notech_ao3 i_86364837(.A(n_26390), .B(imm[22]), .C(n_56108), .Z(n_121281200
		));
	notech_ao3 i_86464836(.A(n_58645), .B(imm[21]), .C(n_56108), .Z(n_121381201
		));
	notech_ao3 i_86564835(.A(n_58645), .B(imm[20]), .C(n_56108), .Z(n_121481202
		));
	notech_ao3 i_86664834(.A(n_58645), .B(imm[19]), .C(n_56108), .Z(n_121581203
		));
	notech_ao3 i_86764833(.A(n_58645), .B(imm[18]), .C(n_56114), .Z(n_121681204
		));
	notech_ao3 i_86864832(.A(n_58645), .B(imm[17]), .C(n_56114), .Z(n_121781205
		));
	notech_ao3 i_87064830(.A(n_58645), .B(imm[15]), .C(n_56114), .Z(n_121881206
		));
	notech_ao3 i_87164829(.A(n_58645), .B(imm[14]), .C(n_56114), .Z(n_121981207
		));
	notech_ao3 i_87264828(.A(n_58645), .B(imm[13]), .C(n_56120), .Z(n_122081208
		));
	notech_ao3 i_87364827(.A(n_58645), .B(imm[12]), .C(n_56120), .Z(n_122181209
		));
	notech_ao3 i_87464826(.A(n_58645), .B(imm[11]), .C(n_56114), .Z(n_122281210
		));
	notech_ao3 i_87564825(.A(n_58645), .B(imm[10]), .C(n_56114), .Z(n_122381211
		));
	notech_ao3 i_87664824(.A(n_58645), .B(imm[9]), .C(n_56114), .Z(n_122481212
		));
	notech_nand2 i_87764823(.A(imm[6]), .B(n_316783142), .Z(n_122581213));
	notech_or2 i_87864822(.A(n_26577), .B(n_28571), .Z(n_122681214));
	notech_or2 i_87964821(.A(n_26577), .B(n_28581), .Z(n_122781215));
	notech_or2 i_88064820(.A(n_26577), .B(n_28583), .Z(n_122881216));
	notech_or2 i_88264818(.A(n_26577), .B(n_28585), .Z(n_122981217));
	notech_nao3 i_88364817(.A(n_58645), .B(n_57432), .C(n_56172), .Z(n_123081218
		));
	notech_or2 i_88464816(.A(n_26577), .B(n_28587), .Z(n_123181219));
	notech_xor2 i_2965639(.A(opz[2]), .B(n_1899), .Z(n_123281220));
	notech_or2 i_88864812(.A(n_26577), .B(n_28588), .Z(n_123381221));
	notech_and2 i_2865640(.A(n_56023), .B(n_55924), .Z(n_123481222));
	notech_ao4 i_1165657(.A(n_1910), .B(n_26497), .C(n_494), .D(n_57442), .Z
		(n_123581223));
	notech_and3 i_965659(.A(n_46243), .B(n_54880), .C(n_46244), .Z(n_123781225
		));
	notech_and4 i_365662(.A(n_57415), .B(n_57417), .C(n_57387), .D(n_57402),
		 .Z(n_123881226));
	notech_or4 i_465661(.A(n_26506), .B(n_26598), .C(n_166281650), .D(n_166381651
		), .Z(n_123981227));
	notech_nand2 i_565660(.A(n_57378), .B(n_57374), .Z(n_124081228));
	notech_or2 i_14365527(.A(n_317383148), .B(n_28611), .Z(n_124481232));
	notech_nand3 i_14065530(.A(n_26785), .B(n_5801), .C(n_312883103), .Z(n_124781235
		));
	notech_or2 i_15865512(.A(n_328583260), .B(n_55299), .Z(n_125481242));
	notech_nao3 i_15165519(.A(n_5812), .B(n_59795), .C(n_57382), .Z(n_126181249
		));
	notech_nand2 i_18565485(.A(opd[4]), .B(n_328983264), .Z(n_128281270));
	notech_or4 i_18265488(.A(n_260988754), .B(n_260888755), .C(n_312083095),
		 .D(n_28735), .Z(n_128581273));
	notech_nao3 i_17965491(.A(n_5820), .B(n_26680), .C(n_55332), .Z(n_128881276
		));
	notech_nao3 i_19565476(.A(n_57448), .B(nbus_144[6]), .C(n_312083095), .Z
		(n_129781285));
	notech_or2 i_18965481(.A(n_311783092), .B(nbus_11326[6]), .Z(n_130281290
		));
	notech_nao3 i_20565466(.A(n_57448), .B(nbus_144[9]), .C(n_312083095), .Z
		(n_130781295));
	notech_or2 i_20065471(.A(n_311783092), .B(nbus_11326[9]), .Z(n_131281300
		));
	notech_nao3 i_21565456(.A(n_57448), .B(nbus_144[10]), .C(n_312083095), .Z
		(n_131781305));
	notech_or2 i_21065461(.A(n_311783092), .B(nbus_11326[10]), .Z(n_132281310
		));
	notech_nao3 i_22565446(.A(n_57448), .B(nbus_144[11]), .C(n_312083095), .Z
		(n_132781315));
	notech_or2 i_22065451(.A(n_311783092), .B(nbus_11326[11]), .Z(n_133281320
		));
	notech_nao3 i_23565436(.A(n_57448), .B(nbus_144[12]), .C(n_312083095), .Z
		(n_133781325));
	notech_or2 i_23065441(.A(n_311783092), .B(nbus_11326[12]), .Z(n_134281330
		));
	notech_nao3 i_24565426(.A(n_57448), .B(nbus_144[13]), .C(n_312083095), .Z
		(n_134781335));
	notech_or2 i_24065431(.A(n_311783092), .B(nbus_11326[13]), .Z(n_135281340
		));
	notech_nao3 i_25565416(.A(n_57438), .B(nbus_144[14]), .C(n_312083095), .Z
		(n_135781345));
	notech_or2 i_25065421(.A(n_311783092), .B(nbus_11326[14]), .Z(n_136281350
		));
	notech_nao3 i_28665406(.A(n_57438), .B(nbus_144[15]), .C(n_312083095), .Z
		(n_136781355));
	notech_or2 i_26665411(.A(n_311783092), .B(nbus_11326[15]), .Z(n_137281360
		));
	notech_ao4 i_30065392(.A(n_312283097), .B(n_125170570), .C(n_55484), .D(n_121781205
		), .Z(n_138181369));
	notech_ao4 i_31165383(.A(n_312283097), .B(n_125170570), .C(n_55484), .D(n_121681204
		), .Z(n_139081378));
	notech_ao4 i_32065374(.A(n_312283097), .B(n_125170570), .C(n_55484), .D(n_121581203
		), .Z(n_139981387));
	notech_ao4 i_33065365(.A(n_312283097), .B(n_125170570), .C(n_55484), .D(n_121481202
		), .Z(n_140881396));
	notech_ao4 i_33965356(.A(n_312283097), .B(n_125170570), .C(n_55484), .D(n_121381201
		), .Z(n_141781405));
	notech_ao4 i_34865347(.A(n_312283097), .B(n_125170570), .C(n_55484), .D(n_121281200
		), .Z(n_142681414));
	notech_ao4 i_35765338(.A(n_312283097), .B(n_125170570), .C(n_55484), .D(n_121181199
		), .Z(n_143581423));
	notech_ao4 i_36665329(.A(n_312283097), .B(n_125170570), .C(n_55484), .D(n_121081198
		), .Z(n_144481432));
	notech_ao4 i_37565320(.A(n_312283097), .B(n_125170570), .C(n_55484), .D(n_120981197
		), .Z(n_145381441));
	notech_ao4 i_38465311(.A(n_312283097), .B(n_125170570), .C(n_55484), .D(n_120881196
		), .Z(n_146281450));
	notech_ao4 i_39365302(.A(n_312283097), .B(n_125170570), .C(n_55484), .D(n_120781195
		), .Z(n_147181459));
	notech_ao4 i_40265293(.A(n_312283097), .B(n_125170570), .C(n_55484), .D(n_120681194
		), .Z(n_148081468));
	notech_ao4 i_41165284(.A(n_312283097), .B(n_125170570), .C(n_55484), .D(n_120581193
		), .Z(n_148981477));
	notech_ao4 i_42265275(.A(n_312283097), .B(n_125170570), .C(n_55484), .D(n_120481192
		), .Z(n_149881486));
	notech_nao3 i_43765260(.A(n_5958), .B(n_59791), .C(n_57382), .Z(n_150381491
		));
	notech_or2 i_43465263(.A(n_311783092), .B(n_59095), .Z(n_150681494));
	notech_or4 i_43165266(.A(n_2269), .B(n_59935), .C(n_56943), .D(opc[31]),
		 .Z(n_150981497));
	notech_or4 i_84164859(.A(n_170581693), .B(n_172281710), .C(n_170281690),
		 .D(n_169981687), .Z(n_164081628));
	notech_and4 i_84264858(.A(n_26652), .B(n_580), .C(mul64[31]), .D(n_26792
		), .Z(n_164181629));
	notech_nor2 i_84364857(.A(n_2386), .B(n_119481182), .Z(n_164281630));
	notech_ao4 i_2265646(.A(n_2768), .B(mul64[31]), .C(n_272988726), .D(n_2837
		), .Z(n_164381631));
	notech_nand2 i_88764813(.A(opz[2]), .B(n_26501), .Z(n_164781635));
	notech_and2 i_89364807(.A(n_26604), .B(n_26590), .Z(n_165281640));
	notech_and2 i_89864802(.A(read_ack), .B(n_26504), .Z(n_165381641));
	notech_or4 i_89764803(.A(n_60773), .B(n_60721), .C(n_55644), .D(n_60583)
		, .Z(n_165681644));
	notech_ao3 i_90764793(.A(n_26621), .B(n_26782), .C(n_55247), .Z(n_165981647
		));
	notech_and3 i_91364787(.A(n_59172), .B(n_59791), .C(n_124081228), .Z(n_166281650
		));
	notech_nand2 i_61765677(.A(n_54862), .B(n_54892), .Z(n_166381651));
	notech_ao4 i_150164218(.A(n_26887), .B(n_26505), .C(n_123881226), .D(n_60474
		), .Z(n_166781655));
	notech_ao4 i_149364224(.A(n_58940), .B(n_2005), .C(n_60463), .D(n_123781225
		), .Z(n_166981657));
	notech_ao4 i_148264234(.A(n_55642), .B(n_56076), .C(n_2176), .D(sema_rw)
		, .Z(n_167181659));
	notech_nand2 i_148464233(.A(n_167181659), .B(n_165681644), .Z(n_167281660
		));
	notech_ao4 i_147364240(.A(n_55642), .B(n_26600), .C(n_123581223), .D(n_29376
		), .Z(n_167781665));
	notech_ao3 i_147264241(.A(n_52420), .B(n_59174), .C(n_51730), .Z(n_168081668
		));
	notech_ao4 i_147064243(.A(n_316383138), .B(n_29120), .C(n_123481222), .D
		(n_27517), .Z(n_168181669));
	notech_and3 i_163065665(.A(n_326183236), .B(n_168181669), .C(n_55888), .Z
		(n_168381671));
	notech_ao4 i_146664246(.A(n_316383138), .B(n_29008), .C(n_55924), .D(n_123281220
		), .Z(n_168481672));
	notech_and4 i_163165664(.A(n_326183236), .B(n_168481672), .C(n_55906), .D
		(n_164781635), .Z(n_168781675));
	notech_and2 i_149665669(.A(n_317283147), .B(n_123081218), .Z(n_168881676
		));
	notech_ao4 i_146464248(.A(n_55919), .B(n_26587), .C(n_48760), .D(n_55934
		), .Z(n_168981677));
	notech_and3 i_162065666(.A(n_168981677), .B(n_56139), .C(n_327546813), .Z
		(n_169081678));
	notech_nand3 i_142664286(.A(n_576), .B(n_62403), .C(n_28975), .Z(n_169181679
		));
	notech_nand3 i_145564257(.A(n_29459), .B(n_29458), .C(n_29460), .Z(n_169381681
		));
	notech_or4 i_145264260(.A(mul64[51]), .B(mul64[48]), .C(mul64[61]), .D(mul64
		[58]), .Z(n_169881686));
	notech_or4 i_145764255(.A(mul64[59]), .B(mul64[56]), .C(n_169381681), .D
		(n_169881686), .Z(n_169981687));
	notech_or4 i_144864264(.A(mul64[52]), .B(mul64[55]), .C(mul64[50]), .D(mul64
		[53]), .Z(n_170281690));
	notech_or4 i_144564267(.A(mul64[33]), .B(mul64[35]), .C(mul64[54]), .D(mul64
		[57]), .Z(n_170581693));
	notech_or4 i_144064272(.A(mul64[34]), .B(mul64[32]), .C(mul64[37]), .D(mul64
		[36]), .Z(n_171081698));
	notech_or4 i_143764275(.A(mul64[41]), .B(mul64[40]), .C(mul64[38]), .D(mul64
		[39]), .Z(n_171381701));
	notech_or4 i_143364279(.A(mul64[44]), .B(mul64[45]), .C(mul64[43]), .D(mul64
		[42]), .Z(n_171781705));
	notech_or4 i_143064282(.A(n_164381631), .B(mul64[49]), .C(mul64[46]), .D
		(mul64[47]), .Z(n_172081708));
	notech_or4 i_144264270(.A(n_172081708), .B(n_171081698), .C(n_171781705)
		, .D(n_171381701), .Z(n_172281710));
	notech_ao4 i_142364289(.A(n_2775), .B(n_29486), .C(n_2774), .D(n_119581183
		), .Z(n_172681714));
	notech_or4 i_117065674(.A(fsm[3]), .B(fsm[0]), .C(n_60761), .D(n_2269), 
		.Z(n_172781715));
	notech_or4 i_32965679(.A(n_60761), .B(n_60719), .C(n_2269), .D(n_56943),
		 .Z(n_172881716));
	notech_ao4 i_141564297(.A(n_54514), .B(n_28675), .C(n_172881716), .D(n_29597
		), .Z(n_172981717));
	notech_ao4 i_141464298(.A(n_172881716), .B(n_29596), .C(n_207041701), .D
		(\nbus_11276[31] ), .Z(n_173081718));
	notech_ao4 i_141364299(.A(n_54491), .B(n_28676), .C(n_54514), .D(n_28674
		), .Z(n_173181719));
	notech_ao4 i_141264300(.A(n_172881716), .B(n_29595), .C(n_119181179), .D
		(n_55234), .Z(n_173281720));
	notech_ao4 i_141164301(.A(n_54514), .B(n_28673), .C(n_54486), .D(n_28675
		), .Z(n_173381721));
	notech_ao4 i_141064302(.A(n_172881716), .B(n_29594), .C(n_119181179), .D
		(n_55249), .Z(n_173481722));
	notech_ao4 i_140964303(.A(n_54486), .B(n_28674), .C(n_54514), .D(n_28672
		), .Z(n_173581723));
	notech_ao4 i_140864304(.A(n_172881716), .B(n_29593), .C(n_119181179), .D
		(n_55261), .Z(n_173681724));
	notech_ao4 i_140764305(.A(n_54481), .B(n_28673), .C(n_54514), .D(n_28671
		), .Z(n_173781725));
	notech_ao4 i_140664306(.A(n_172881716), .B(n_29592), .C(n_119181179), .D
		(n_59328), .Z(n_173881726));
	notech_ao4 i_140564307(.A(n_54481), .B(n_28672), .C(n_54513), .D(n_28670
		), .Z(n_173981727));
	notech_ao4 i_140464308(.A(n_172881716), .B(n_29591), .C(n_119181179), .D
		(n_59337), .Z(n_174081728));
	notech_ao4 i_140364309(.A(n_54486), .B(n_28671), .C(n_54498), .D(n_28669
		), .Z(n_174181729));
	notech_ao4 i_140264310(.A(n_172881716), .B(n_29590), .C(n_119181179), .D
		(n_59346), .Z(n_174281730));
	notech_ao4 i_140164311(.A(n_54486), .B(n_28670), .C(n_54498), .D(n_28668
		), .Z(n_174381731));
	notech_ao4 i_140064312(.A(n_172881716), .B(n_29589), .C(n_119181179), .D
		(\nbus_11276[24] ), .Z(n_174481732));
	notech_ao4 i_139964313(.A(n_54486), .B(n_28669), .C(n_54498), .D(n_28667
		), .Z(n_174581733));
	notech_ao4 i_139864314(.A(n_172881716), .B(n_29588), .C(n_119181179), .D
		(n_59319), .Z(n_174681734));
	notech_ao4 i_139764315(.A(n_54486), .B(n_28668), .C(n_54498), .D(n_28666
		), .Z(n_174781735));
	notech_ao4 i_139664316(.A(n_172881716), .B(n_29587), .C(n_119181179), .D
		(n_55647), .Z(n_174881736));
	notech_ao4 i_139564317(.A(n_54481), .B(n_28667), .C(n_54498), .D(n_28665
		), .Z(n_174981737));
	notech_ao4 i_139464318(.A(n_172881716), .B(n_29586), .C(n_119181179), .D
		(n_59310), .Z(n_175081738));
	notech_ao4 i_139364319(.A(n_54481), .B(n_28666), .C(n_54498), .D(n_28664
		), .Z(n_175181739));
	notech_ao4 i_139264320(.A(n_172881716), .B(n_29585), .C(n_119181179), .D
		(n_55631), .Z(n_175281740));
	notech_ao4 i_139164321(.A(n_54481), .B(n_28665), .C(n_54498), .D(n_28663
		), .Z(n_175381741));
	notech_ao4 i_139064322(.A(n_172881716), .B(n_29584), .C(n_119181179), .D
		(n_55620), .Z(n_175481742));
	notech_ao4 i_138964323(.A(n_54481), .B(n_28664), .C(n_54498), .D(n_28662
		), .Z(n_175581743));
	notech_ao4 i_138864324(.A(n_172881716), .B(n_29583), .C(n_119181179), .D
		(n_55609), .Z(n_175681744));
	notech_ao4 i_138764325(.A(n_54481), .B(n_28663), .C(n_54498), .D(n_28661
		), .Z(n_175781745));
	notech_ao4 i_138664326(.A(n_172881716), .B(n_29582), .C(n_119181179), .D
		(n_55600), .Z(n_175881746));
	notech_ao4 i_138564327(.A(n_54481), .B(n_28662), .C(n_54498), .D(n_28660
		), .Z(n_175981747));
	notech_ao4 i_138464328(.A(n_172881716), .B(n_29581), .C(n_119181179), .D
		(n_55590), .Z(n_176081748));
	notech_ao4 i_138364329(.A(n_54481), .B(n_28661), .C(n_54498), .D(n_28659
		), .Z(n_176181749));
	notech_ao4 i_138264330(.A(n_54344), .B(n_29580), .C(n_119181179), .D(n_55578
		), .Z(n_176281750));
	notech_ao4 i_138164331(.A(n_54481), .B(n_28660), .C(n_54498), .D(n_28658
		), .Z(n_176381751));
	notech_ao4 i_138064332(.A(n_54344), .B(n_29579), .C(n_54335), .D(n_55566
		), .Z(n_176481752));
	notech_ao4 i_137964333(.A(n_54486), .B(n_28659), .C(n_54498), .D(n_28657
		), .Z(n_176581753));
	notech_ao4 i_137864334(.A(n_54344), .B(n_29578), .C(n_54335), .D(n_55552
		), .Z(n_176681754));
	notech_ao4 i_137764335(.A(n_54486), .B(n_28658), .C(n_54498), .D(n_28656
		), .Z(n_176781755));
	notech_ao4 i_137664336(.A(n_54344), .B(n_29577), .C(n_54335), .D(n_55542
		), .Z(n_176881756));
	notech_ao4 i_137564337(.A(n_54486), .B(n_28657), .C(n_54498), .D(n_28655
		), .Z(n_176981757));
	notech_ao4 i_137464338(.A(n_54344), .B(n_29576), .C(n_54335), .D(n_55469
		), .Z(n_177081758));
	notech_ao4 i_137364339(.A(n_54486), .B(n_28656), .C(n_54498), .D(n_28654
		), .Z(n_177181759));
	notech_ao4 i_137264340(.A(n_54344), .B(n_29575), .C(n_54335), .D(n_55438
		), .Z(n_177281760));
	notech_ao4 i_137164341(.A(n_54491), .B(n_28655), .C(n_54498), .D(n_28653
		), .Z(n_177381761));
	notech_ao4 i_137064342(.A(n_54344), .B(n_29574), .C(n_54335), .D(n_55425
		), .Z(n_177481762));
	notech_ao4 i_136964343(.A(n_54491), .B(n_28654), .C(n_54498), .D(n_28652
		), .Z(n_177581763));
	notech_ao4 i_136864344(.A(n_54344), .B(n_29573), .C(n_54335), .D(n_55413
		), .Z(n_177681764));
	notech_ao4 i_136764345(.A(n_54486), .B(n_28653), .C(n_54504), .D(n_28651
		), .Z(n_177781765));
	notech_ao4 i_136064346(.A(n_54344), .B(n_29572), .C(n_54335), .D(n_55400
		), .Z(n_177881766));
	notech_ao4 i_135864347(.A(n_54486), .B(n_28652), .C(n_54504), .D(n_28650
		), .Z(n_177981767));
	notech_ao4 i_135764348(.A(n_54344), .B(n_29571), .C(n_54335), .D(n_55387
		), .Z(n_178081768));
	notech_ao4 i_135664349(.A(n_54486), .B(n_28651), .C(n_54504), .D(n_28649
		), .Z(n_178181769));
	notech_ao4 i_135564350(.A(n_172881716), .B(n_29570), .C(n_54335), .D(n_55375
		), .Z(n_178281770));
	notech_ao4 i_135464351(.A(n_54486), .B(n_28650), .C(n_54504), .D(n_28648
		), .Z(n_178381771));
	notech_ao4 i_135364352(.A(n_54344), .B(n_29569), .C(n_54335), .D(n_55365
		), .Z(n_178481772));
	notech_ao4 i_135264353(.A(n_54486), .B(n_28649), .C(n_54504), .D(n_28647
		), .Z(n_178581773));
	notech_ao4 i_135164354(.A(n_54344), .B(n_29568), .C(n_54335), .D(\nbus_11276[3] 
		), .Z(n_178681774));
	notech_ao4 i_135064355(.A(n_54486), .B(n_28648), .C(n_54504), .D(n_28645
		), .Z(n_178781775));
	notech_ao4 i_134964356(.A(n_54344), .B(n_29567), .C(n_54335), .D(n_55289
		), .Z(n_178881776));
	notech_ao4 i_134864357(.A(n_54486), .B(n_28647), .C(n_54504), .D(n_28644
		), .Z(n_178981777));
	notech_ao4 i_134764358(.A(n_54344), .B(n_29566), .C(n_54335), .D(n_59753
		), .Z(n_179081778));
	notech_ao4 i_134664359(.A(n_54486), .B(n_28645), .C(n_54504), .D(n_28643
		), .Z(n_179181779));
	notech_ao4 i_133864367(.A(n_54344), .B(n_29565), .C(n_54335), .D(n_55356
		), .Z(n_179281780));
	notech_or4 i_30565680(.A(n_60761), .B(n_60719), .C(n_2269), .D(n_59095),
		 .Z(n_179381781));
	notech_ao4 i_127064434(.A(n_27554), .B(n_126470583), .C(n_207341704), .D
		(n_28642), .Z(n_179481782));
	notech_ao4 i_126864436(.A(n_207841709), .B(n_28866), .C(n_54388), .D(opb
		[31]), .Z(n_179681784));
	notech_and4 i_127264432(.A(n_179681784), .B(n_179481782), .C(n_150681494
		), .D(n_150981497), .Z(n_179881786));
	notech_ao4 i_126564439(.A(n_312083095), .B(n_28767), .C(n_311683091), .D
		(n_58951), .Z(n_179981787));
	notech_ao4 i_126464440(.A(n_311583090), .B(n_29564), .C(n_311483089), .D
		(n_29563), .Z(n_180181789));
	notech_ao4 i_126164443(.A(n_126470583), .B(n_27553), .C(n_207341704), .D
		(n_28641), .Z(n_180481791));
	notech_ao4 i_126064444(.A(n_311683091), .B(nbus_11273[30]), .C(n_311783092
		), .D(n_59050), .Z(n_180781793));
	notech_ao3 i_126364441(.A(n_180481791), .B(n_180781793), .C(n_149881486)
		, .Z(n_180881794));
	notech_ao4 i_125864446(.A(n_311383088), .B(n_29562), .C(n_312083095), .D
		(n_28766), .Z(n_180981795));
	notech_ao4 i_125764447(.A(n_311583090), .B(n_29561), .C(n_311483089), .D
		(n_29560), .Z(n_181081796));
	notech_ao4 i_125464450(.A(n_126470583), .B(n_27552), .C(n_207341704), .D
		(n_28640), .Z(n_181281798));
	notech_ao4 i_125364451(.A(n_311683091), .B(n_56892), .C(n_311783092), .D
		(n_59104), .Z(n_181481800));
	notech_ao3 i_125664448(.A(n_181281798), .B(n_181481800), .C(n_148981477)
		, .Z(n_181581801));
	notech_ao4 i_125164453(.A(n_311383088), .B(n_29559), .C(n_312083095), .D
		(n_28764), .Z(n_181681802));
	notech_ao4 i_125064454(.A(n_311583090), .B(n_29558), .C(n_311483089), .D
		(n_29557), .Z(n_181981803));
	notech_ao4 i_124764457(.A(n_126470583), .B(n_27551), .C(n_207341704), .D
		(n_28639), .Z(n_182181805));
	notech_ao4 i_124664458(.A(n_311683091), .B(n_56883), .C(n_311783092), .D
		(n_59077), .Z(n_182381807));
	notech_ao3 i_124964455(.A(n_182181805), .B(n_182381807), .C(n_148081468)
		, .Z(n_182681808));
	notech_ao4 i_124464460(.A(n_311383088), .B(n_29556), .C(n_312083095), .D
		(n_28763), .Z(n_182781809));
	notech_ao4 i_124364461(.A(n_311583090), .B(n_29555), .C(n_311483089), .D
		(n_29554), .Z(n_182881810));
	notech_ao4 i_124064464(.A(n_126470583), .B(n_27550), .C(n_207341704), .D
		(n_28638), .Z(n_183081812));
	notech_ao4 i_123964465(.A(n_311683091), .B(n_56874), .C(n_311783092), .D
		(n_59059), .Z(n_183281814));
	notech_ao3 i_124264462(.A(n_183081812), .B(n_183281814), .C(n_147181459)
		, .Z(n_183381815));
	notech_ao4 i_123764467(.A(n_311383088), .B(n_29553), .C(n_54519), .D(n_28758
		), .Z(n_183481816));
	notech_ao4 i_123664468(.A(n_311583090), .B(n_29552), .C(n_311483089), .D
		(n_29551), .Z(n_183581817));
	notech_ao4 i_123364471(.A(n_126470583), .B(n_27549), .C(n_207341704), .D
		(n_28637), .Z(n_183781819));
	notech_ao4 i_123264472(.A(n_311683091), .B(n_56865), .C(n_311783092), .D
		(n_59068), .Z(n_183981821));
	notech_ao3 i_123564469(.A(n_183781819), .B(n_183981821), .C(n_146281450)
		, .Z(n_184081822));
	notech_ao4 i_123064474(.A(n_311383088), .B(n_29550), .C(n_54519), .D(n_28757
		), .Z(n_184181823));
	notech_ao4 i_122964475(.A(n_311583090), .B(n_29549), .C(n_311483089), .D
		(n_29548), .Z(n_184281824));
	notech_ao4 i_122664478(.A(n_126470583), .B(n_27548), .C(n_207341704), .D
		(n_28636), .Z(n_184481826));
	notech_ao4 i_122564479(.A(n_311683091), .B(n_56856), .C(n_311783092), .D
		(n_59023), .Z(n_184681828));
	notech_ao3 i_122864476(.A(n_184481826), .B(n_184681828), .C(n_145381441)
		, .Z(n_184781829));
	notech_ao4 i_122364481(.A(n_311383088), .B(n_29547), .C(n_54519), .D(n_28756
		), .Z(n_184881830));
	notech_ao4 i_122264482(.A(n_311583090), .B(n_29546), .C(n_311483089), .D
		(n_29545), .Z(n_184981831));
	notech_ao4 i_121964485(.A(n_126470583), .B(n_27546), .C(n_207341704), .D
		(n_28635), .Z(n_185181833));
	notech_ao4 i_121864486(.A(n_311683091), .B(n_56847), .C(n_54416), .D(n_59086
		), .Z(n_185381835));
	notech_ao3 i_122164483(.A(n_185181833), .B(n_185381835), .C(n_144481432)
		, .Z(n_185481836));
	notech_ao4 i_121664488(.A(n_311383088), .B(n_29544), .C(n_54519), .D(n_28755
		), .Z(n_185581837));
	notech_ao4 i_121564489(.A(n_311583090), .B(n_29543), .C(n_311483089), .D
		(n_29542), .Z(n_185681838));
	notech_ao4 i_121264492(.A(n_126470583), .B(n_27545), .C(n_207341704), .D
		(n_28634), .Z(n_185881840));
	notech_ao4 i_121164493(.A(n_311683091), .B(n_56838), .C(n_54416), .D(n_59041
		), .Z(n_186081842));
	notech_ao3 i_121464490(.A(n_185881840), .B(n_186081842), .C(n_143581423)
		, .Z(n_186181843));
	notech_ao4 i_120964495(.A(n_311383088), .B(n_29541), .C(n_54519), .D(n_28754
		), .Z(n_186281844));
	notech_ao4 i_120864496(.A(n_311583090), .B(n_29540), .C(n_311483089), .D
		(n_29539), .Z(n_186381845));
	notech_ao4 i_120564499(.A(n_126470583), .B(n_27542), .C(n_207341704), .D
		(n_28633), .Z(n_186581847));
	notech_ao4 i_120464500(.A(n_311683091), .B(n_56829), .C(n_54416), .D(n_59032
		), .Z(n_186781849));
	notech_ao3 i_120764497(.A(n_186581847), .B(n_186781849), .C(n_142681414)
		, .Z(n_186881850));
	notech_ao4 i_120264502(.A(n_311383088), .B(n_29538), .C(n_54519), .D(n_28753
		), .Z(n_186981851));
	notech_ao4 i_120164503(.A(n_311583090), .B(n_29537), .C(n_311483089), .D
		(n_29536), .Z(n_187081852));
	notech_ao4 i_119864506(.A(n_126470583), .B(n_27541), .C(n_207341704), .D
		(n_28632), .Z(n_187281854));
	notech_ao4 i_119764507(.A(n_311683091), .B(n_56820), .C(n_54416), .D(n_58996
		), .Z(n_187481856));
	notech_ao3 i_120064504(.A(n_187281854), .B(n_187481856), .C(n_141781405)
		, .Z(n_187581857));
	notech_ao4 i_119564509(.A(n_311383088), .B(n_29535), .C(n_54519), .D(n_28752
		), .Z(n_187681858));
	notech_ao4 i_119464510(.A(n_311583090), .B(n_29534), .C(n_311483089), .D
		(n_29533), .Z(n_187781859));
	notech_ao4 i_119164513(.A(n_126470583), .B(n_27540), .C(n_207341704), .D
		(n_28631), .Z(n_187981861));
	notech_ao4 i_119064514(.A(n_311683091), .B(n_56811), .C(n_54416), .D(n_59005
		), .Z(n_188181863));
	notech_ao3 i_119364511(.A(n_187981861), .B(n_188181863), .C(n_140881396)
		, .Z(n_188281864));
	notech_ao4 i_118864516(.A(n_311383088), .B(n_29532), .C(n_54519), .D(n_28751
		), .Z(n_188381865));
	notech_ao4 i_118764517(.A(n_311583090), .B(n_29531), .C(n_311483089), .D
		(n_29530), .Z(n_188481866));
	notech_ao4 i_118464520(.A(n_126470583), .B(n_27539), .C(n_207341704), .D
		(n_28630), .Z(n_188681868));
	notech_ao4 i_118364521(.A(n_311683091), .B(n_56802), .C(n_54416), .D(n_59014
		), .Z(n_188881870));
	notech_ao3 i_118664518(.A(n_188681868), .B(n_188881870), .C(n_139981387)
		, .Z(n_188981871));
	notech_ao4 i_118164523(.A(n_311383088), .B(n_29529), .C(n_54519), .D(n_28750
		), .Z(n_189081872));
	notech_ao4 i_118064524(.A(n_311583090), .B(n_29528), .C(n_311483089), .D
		(n_29527), .Z(n_189181873));
	notech_ao4 i_117764527(.A(n_126470583), .B(n_27538), .C(n_207341704), .D
		(n_28629), .Z(n_189381875));
	notech_ao4 i_117664528(.A(n_311683091), .B(n_56793), .C(n_54416), .D(n_58969
		), .Z(n_189581877));
	notech_ao3 i_117964525(.A(n_189381875), .B(n_189581877), .C(n_139081378)
		, .Z(n_189681878));
	notech_ao4 i_117464530(.A(n_311383088), .B(n_29526), .C(n_54519), .D(n_28749
		), .Z(n_189781879));
	notech_ao4 i_117364531(.A(n_311583090), .B(n_29525), .C(n_311483089), .D
		(n_29524), .Z(n_189881880));
	notech_ao4 i_116964534(.A(n_126470583), .B(n_27537), .C(n_207341704), .D
		(n_28628), .Z(n_190081882));
	notech_ao4 i_116864535(.A(n_311683091), .B(n_56784), .C(n_54416), .D(n_58978
		), .Z(n_190281884));
	notech_ao3 i_117264532(.A(n_190081882), .B(n_190281884), .C(n_138181369)
		, .Z(n_190381885));
	notech_ao4 i_116664537(.A(n_54449), .B(n_29523), .C(n_54519), .D(n_28748
		), .Z(n_190481886));
	notech_ao4 i_116564538(.A(n_311583090), .B(n_29522), .C(n_54472), .D(n_29521
		), .Z(n_190581887));
	notech_ao4 i_115464548(.A(n_312183096), .B(n_27534), .C(n_28865), .D(n_307583050
		), .Z(n_190781889));
	notech_ao4 i_115364549(.A(n_54449), .B(n_29520), .C(n_54427), .D(n_56766
		), .Z(n_190981891));
	notech_and3 i_115664546(.A(n_190781889), .B(n_190981891), .C(n_137281360
		), .Z(n_191081892));
	notech_ao4 i_115064552(.A(n_54405), .B(n_29519), .C(n_54472), .D(n_29518
		), .Z(n_191181893));
	notech_ao4 i_114964553(.A(n_307183046), .B(n_28626), .C(n_311983094), .D
		(n_28746), .Z(n_191381895));
	notech_ao4 i_114664556(.A(n_312183096), .B(n_27533), .C(n_28864), .D(n_307583050
		), .Z(n_191581897));
	notech_ao4 i_114564557(.A(n_54449), .B(n_29517), .C(n_54427), .D(n_56757
		), .Z(n_191781899));
	notech_and3 i_114864554(.A(n_191581897), .B(n_191781899), .C(n_136281350
		), .Z(n_191881900));
	notech_ao4 i_114264560(.A(n_54405), .B(n_29516), .C(n_54472), .D(n_29515
		), .Z(n_191981901));
	notech_ao4 i_114164561(.A(n_307183046), .B(n_28625), .C(n_311983094), .D
		(n_28745), .Z(n_192181903));
	notech_ao4 i_113864564(.A(n_312183096), .B(n_27532), .C(n_28863), .D(n_307583050
		), .Z(n_192381905));
	notech_ao4 i_113764565(.A(n_54449), .B(n_29514), .C(n_54427), .D(n_56748
		), .Z(n_192581907));
	notech_and3 i_114064562(.A(n_192381905), .B(n_192581907), .C(n_135281340
		), .Z(n_192681908));
	notech_ao4 i_113464568(.A(n_54405), .B(n_29513), .C(n_54472), .D(n_29512
		), .Z(n_192781909));
	notech_ao4 i_113364569(.A(n_307183046), .B(n_28624), .C(n_311983094), .D
		(n_28744), .Z(n_192981911));
	notech_ao4 i_113064572(.A(n_312183096), .B(n_27531), .C(n_28862), .D(n_307583050
		), .Z(n_193181913));
	notech_ao4 i_112964573(.A(n_54449), .B(n_29511), .C(n_56739), .D(n_54427
		), .Z(n_193381915));
	notech_and3 i_113264570(.A(n_134281330), .B(n_193181913), .C(n_193381915
		), .Z(n_193481916));
	notech_ao4 i_112664576(.A(n_54405), .B(n_29510), .C(n_54472), .D(n_29509
		), .Z(n_193581917));
	notech_ao4 i_112564577(.A(n_307183046), .B(n_28623), .C(n_311983094), .D
		(n_28743), .Z(n_193781919));
	notech_ao4 i_112264580(.A(n_312183096), .B(n_27530), .C(n_28861), .D(n_307583050
		), .Z(n_193981921));
	notech_ao4 i_112164581(.A(n_54449), .B(n_29508), .C(n_54427), .D(n_56730
		), .Z(n_194181923));
	notech_and3 i_112464578(.A(n_133281320), .B(n_193981921), .C(n_194181923
		), .Z(n_194281924));
	notech_ao4 i_111864584(.A(n_54405), .B(n_29507), .C(n_54472), .D(n_29506
		), .Z(n_194381925));
	notech_ao4 i_111764585(.A(n_307183046), .B(n_28622), .C(n_311983094), .D
		(n_28742), .Z(n_194581927));
	notech_ao4 i_111464588(.A(n_312183096), .B(n_27529), .C(n_28860), .D(n_307583050
		), .Z(n_194781929));
	notech_ao4 i_111364589(.A(n_54449), .B(n_29505), .C(n_54427), .D(nbus_11273
		[10]), .Z(n_194981931));
	notech_and3 i_111664586(.A(n_194781929), .B(n_194981931), .C(n_132281310
		), .Z(n_195081932));
	notech_ao4 i_111064592(.A(n_54405), .B(n_29504), .C(n_54472), .D(n_29503
		), .Z(n_195181933));
	notech_ao4 i_110964593(.A(n_307183046), .B(n_28621), .C(n_311983094), .D
		(n_28741), .Z(n_195381935));
	notech_ao4 i_110664596(.A(n_312183096), .B(n_27528), .C(n_28859), .D(n_307583050
		), .Z(n_195581937));
	notech_ao4 i_110564597(.A(n_54449), .B(n_29502), .C(n_54427), .D(n_56712
		), .Z(n_195781939));
	notech_and3 i_110864594(.A(n_131281300), .B(n_195581937), .C(n_195781939
		), .Z(n_195881940));
	notech_ao4 i_110264600(.A(n_54405), .B(n_29501), .C(n_54472), .D(n_29500
		), .Z(n_195981941));
	notech_ao4 i_110164601(.A(n_307183046), .B(n_28620), .C(n_311983094), .D
		(n_28740), .Z(n_196181943));
	notech_ao4 i_109864604(.A(n_312183096), .B(n_27525), .C(n_307583050), .D
		(n_28857), .Z(n_196381945));
	notech_ao4 i_109764605(.A(n_54449), .B(n_29499), .C(n_54427), .D(n_56694
		), .Z(n_196581947));
	notech_and3 i_110064602(.A(n_196381945), .B(n_196581947), .C(n_130281290
		), .Z(n_196681948));
	notech_ao4 i_109464608(.A(n_54405), .B(n_29498), .C(n_54472), .D(n_29497
		), .Z(n_196781949));
	notech_ao4 i_109364609(.A(n_307183046), .B(n_28617), .C(n_311983094), .D
		(n_28737), .Z(n_196981951));
	notech_ao4 i_109064612(.A(n_318383158), .B(n_169081678), .C(n_118881176)
		, .D(opd[4]), .Z(n_197181953));
	notech_ao4 i_108964613(.A(n_54416), .B(nbus_11326[4]), .C(n_316483139), 
		.D(n_27523), .Z(n_197281954));
	notech_ao4 i_108764615(.A(n_311383088), .B(n_29496), .C(n_54427), .D(n_56676
		), .Z(n_197481956));
	notech_and4 i_109264610(.A(n_197481956), .B(n_197281954), .C(n_197181953
		), .D(n_128881276), .Z(n_197681958));
	notech_ao4 i_108464618(.A(n_311883093), .B(n_28727), .C(n_54405), .D(n_29495
		), .Z(n_197781959));
	notech_ao4 i_108264620(.A(n_316683141), .B(n_28583), .C(n_317383148), .D
		(n_28615), .Z(n_197981961));
	notech_and4 i_108664616(.A(n_197981961), .B(n_197781959), .C(n_128281270
		), .D(n_128581273), .Z(n_198181963));
	notech_ao4 i_107964623(.A(n_58895), .B(n_55149), .C(n_318383158), .D(n_168881676
		), .Z(n_198281964));
	notech_ao4 i_107864624(.A(n_54416), .B(nbus_11326[3]), .C(n_316483139), 
		.D(n_27522), .Z(n_198381965));
	notech_ao4 i_107664626(.A(n_54449), .B(n_29494), .C(n_54427), .D(n_56667
		), .Z(n_198581967));
	notech_ao4 i_107564627(.A(n_54405), .B(n_29493), .C(n_54472), .D(n_29492
		), .Z(n_198681968));
	notech_and4 i_108164621(.A(n_198681968), .B(n_198581967), .C(n_198381965
		), .D(n_198281964), .Z(n_198881970));
	notech_ao4 i_107264630(.A(n_311983094), .B(n_28734), .C(n_311883093), .D
		(n_28726), .Z(n_198981971));
	notech_mux2 i_107164631(.S(opd[3]), .A(n_325783232), .B(n_328783262), .Z
		(n_199081972));
	notech_ao4 i_106964633(.A(n_316683141), .B(n_28585), .C(n_317383148), .D
		(n_28614), .Z(n_199281974));
	notech_and4 i_107464628(.A(n_328283257), .B(n_199281974), .C(n_198981971
		), .D(n_199081972), .Z(n_199481976));
	notech_ao4 i_106664636(.A(n_318383158), .B(n_168781675), .C(opd[2]), .D(n_118781175
		), .Z(n_199581977));
	notech_ao4 i_106564637(.A(n_316483139), .B(n_27521), .C(n_58895), .D(n_1967
		), .Z(n_199681978));
	notech_ao4 i_106364639(.A(n_54427), .B(n_56658), .C(n_54416), .D(nbus_11326
		[2]), .Z(n_199881980));
	notech_and4 i_106864634(.A(n_199881980), .B(n_199681978), .C(n_199581977
		), .D(n_126181249), .Z(n_200081982));
	notech_ao4 i_106064642(.A(n_54405), .B(n_29491), .C(n_54472), .D(n_29490
		), .Z(n_200181983));
	notech_ao4 i_105964643(.A(n_311983094), .B(n_28733), .C(n_311883093), .D
		(n_28725), .Z(n_200281984));
	notech_ao4 i_105764645(.A(n_316683141), .B(n_28587), .C(n_317383148), .D
		(n_28613), .Z(n_200481986));
	notech_and4 i_106264640(.A(n_200481986), .B(n_200281984), .C(n_200181983
		), .D(n_125481242), .Z(n_200681988));
	notech_ao4 i_105464648(.A(n_316483139), .B(n_27519), .C(n_318383158), .D
		(n_168381671), .Z(n_200781989));
	notech_ao4 i_105364649(.A(n_54427), .B(n_58960), .C(n_54416), .D(nbus_11326
		[0]), .Z(n_200881990));
	notech_ao4 i_105164651(.A(n_54472), .B(n_29489), .C(n_54449), .D(n_29488
		), .Z(n_201081992));
	notech_and4 i_105664646(.A(n_201081992), .B(n_200881990), .C(n_200781989
		), .D(n_124781235), .Z(n_201281994));
	notech_ao4 i_104864654(.A(n_311983094), .B(n_28731), .C(n_311883093), .D
		(n_28723), .Z(n_201381995));
	notech_ao4 i_104664656(.A(n_327883253), .B(opd[0]), .C(n_316683141), .D(n_28588
		), .Z(n_201581997));
	notech_and4 i_105064652(.A(n_201581997), .B(n_201381995), .C(n_316583140
		), .D(n_124481232), .Z(n_201781999));
	notech_ao3 i_67762893(.A(n_58645), .B(imm[8]), .C(n_56114), .Z(n_201882000
		));
	notech_and2 i_18063371(.A(n_202282004), .B(n_55210), .Z(n_202082002));
	notech_or4 i_73162841(.A(n_274588712), .B(n_2572), .C(n_272988726), .D(tcmp
		), .Z(n_202282004));
	notech_mux2 i_15963392(.S(reps[2]), .A(n_2168), .B(n_325883233), .Z(n_202482006
		));
	notech_ao3 i_16063391(.A(n_206482046), .B(n_270739495), .C(n_26543), .Z(n_202682008
		));
	notech_or4 i_21463345(.A(n_260988754), .B(n_260888755), .C(n_54519), .D(n_28739
		), .Z(n_203382015));
	notech_nao3 i_20963350(.A(n_5840), .B(n_26680), .C(n_55332), .Z(n_203882020
		));
	notech_or4 i_46263103(.A(n_59370), .B(n_58895), .C(n_59935), .D(nbus_11326
		[4]), .Z(n_203982021));
	notech_or2 i_46163104(.A(n_54435), .B(n_29063), .Z(n_204282024));
	notech_or2 i_45663109(.A(n_54565), .B(n_56676), .Z(n_204782029));
	notech_or4 i_65162918(.A(n_56196), .B(n_56163), .C(n_55827), .D(n_319588494
		), .Z(n_204882030));
	notech_or2 i_64662923(.A(n_54438), .B(n_29063), .Z(n_205582037));
	notech_or2 i_66762903(.A(n_144377843), .B(n_55965), .Z(n_205682038));
	notech_or2 i_66262908(.A(n_54438), .B(n_29068), .Z(n_206382045));
	notech_and3 i_25616(.A(n_55745), .B(n_54874), .C(n_1960), .Z(n_206482046
		));
	notech_ao4 i_145162141(.A(n_316488525), .B(n_279739585), .C(n_316588524)
		, .D(n_275539543), .Z(n_206682048));
	notech_ao4 i_145062142(.A(n_54655), .B(n_55387), .C(n_57352), .D(n_54469
		), .Z(n_206882050));
	notech_ao4 i_144862144(.A(n_27568), .B(n_55756), .C(n_54656), .D(n_56694
		), .Z(n_207082052));
	notech_and4 i_144962143(.A(n_183578230), .B(n_183478229), .C(n_205682038
		), .D(n_207082052), .Z(n_207282054));
	notech_ao4 i_143862154(.A(n_279739585), .B(n_316388526), .C(n_275539543)
		, .D(n_316288527), .Z(n_207382055));
	notech_ao4 i_143762155(.A(n_54655), .B(n_55365), .C(n_54469), .D(n_321188478
		), .Z(n_207582057));
	notech_ao4 i_143562157(.A(n_55756), .B(n_27565), .C(n_54656), .D(n_56676
		), .Z(n_207782059));
	notech_and3 i_143662156(.A(n_137970698), .B(n_204882030), .C(n_207782059
		), .Z(n_207982061));
	notech_ao4 i_126762322(.A(n_139770716), .B(n_56382), .C(n_58548), .D(n_26539
		), .Z(n_208082062));
	notech_ao4 i_126662323(.A(n_316288527), .B(n_247234098), .C(n_54563), .D
		(n_55365), .Z(n_208282064));
	notech_ao4 i_126362326(.A(n_321188478), .B(n_54458), .C(n_316388526), .D
		(n_247334099), .Z(n_208482066));
	notech_and4 i_126562324(.A(n_208482066), .B(n_137970698), .C(n_203982021
		), .D(n_204282024), .Z(n_208782069));
	notech_ao4 i_104162542(.A(n_54449), .B(n_29599), .C(n_28858), .D(n_307583050
		), .Z(n_208882070));
	notech_ao4 i_104062543(.A(n_54427), .B(n_56703), .C(n_54405), .D(n_29598
		), .Z(n_209082072));
	notech_and3 i_104462540(.A(n_208882070), .B(n_209082072), .C(n_203882020
		), .Z(n_209182073));
	notech_ao4 i_103762546(.A(n_311883093), .B(n_28730), .C(n_54416), .D(nbus_11326
		[8]), .Z(n_209282074));
	notech_ao4 i_103662547(.A(n_307183046), .B(n_28619), .C(n_312183096), .D
		(n_27527), .Z(n_209482076));
	notech_nand3 i_18260373(.A(n_54124), .B(tsc[29]), .C(n_59791), .Z(n_209682078
		));
	notech_nand2 i_18160374(.A(n_351965808), .B(opc[29]), .Z(n_209982081));
	notech_or2 i_17660379(.A(n_55143), .B(n_56892), .Z(n_210482086));
	notech_ao3 i_47860101(.A(n_62411), .B(opc[4]), .C(n_320688483), .Z(n_210982091
		));
	notech_or2 i_47460104(.A(n_319088499), .B(n_56676), .Z(n_211282094));
	notech_ao4 i_128559360(.A(n_59163), .B(n_27523), .C(n_59174), .D(n_26720
		), .Z(n_211782099));
	notech_ao4 i_128359361(.A(n_55688), .B(n_319588494), .C(n_319288497), .D
		(n_58548), .Z(n_211882100));
	notech_ao4 i_128159363(.A(n_55222), .B(n_29063), .C(n_55238), .D(n_321188478
		), .Z(n_212082102));
	notech_and4 i_128759358(.A(n_212082102), .B(n_211882100), .C(n_211782099
		), .D(n_211282094), .Z(n_212282104));
	notech_ao4 i_127859366(.A(n_320188488), .B(n_316288527), .C(n_318888501)
		, .D(\nbus_11276[4] ), .Z(n_212382105));
	notech_ao4 i_127659368(.A(n_321688474), .B(n_29601), .C(n_54024), .D(n_29600
		), .Z(n_212582107));
	notech_nand3 i_127759367(.A(n_169564033), .B(n_174464082), .C(n_212582107
		), .Z(n_212682108));
	notech_ao4 i_96959659(.A(n_55142), .B(n_55249), .C(n_56023), .D(n_262936784
		), .Z(n_212882110));
	notech_ao4 i_96859660(.A(n_28977), .B(n_26565), .C(n_57329), .D(n_352165810
		), .Z(n_213082112));
	notech_ao4 i_96559663(.A(n_352965818), .B(n_110923096), .C(n_270688747),
		 .D(n_352365812), .Z(n_213282114));
	notech_and4 i_96759661(.A(n_262736782), .B(n_213282114), .C(n_209682078)
		, .D(n_209982081), .Z(n_213582117));
	notech_and2 i_93556982(.A(n_253034156), .B(n_26589), .Z(n_213682118));
	notech_nand3 i_71457193(.A(n_59780), .B(n_59936), .C(read_data[8]), .Z(n_214182123
		));
	notech_nand2 i_70957198(.A(n_55268), .B(opa[8]), .Z(n_214682128));
	notech_ao4 i_149056461(.A(n_157974447), .B(n_55947), .C(n_161857906), .D
		(n_248534111), .Z(n_214782129));
	notech_ao4 i_148956462(.A(n_55354), .B(n_29045), .C(n_55310), .D(n_55413
		), .Z(n_214982131));
	notech_and3 i_149256459(.A(n_214782129), .B(n_214982131), .C(n_214682128
		), .Z(n_215082132));
	notech_ao4 i_148656465(.A(n_54822), .B(n_29102), .C(n_55727), .D(n_27571
		), .Z(n_215182133));
	notech_ao4 i_148556466(.A(n_161957907), .B(n_2326), .C(n_55156), .D(n_57350
		), .Z(n_215382135));
	notech_or2 i_26255043(.A(n_54853), .B(n_29087), .Z(n_215582137));
	notech_or4 i_25755048(.A(n_56081), .B(n_59281), .C(n_57293), .D(n_55852)
		, .Z(n_216282144));
	notech_or4 i_50054808(.A(n_55522), .B(n_56449), .C(n_324883223), .D(n_174358031
		), .Z(n_216982151));
	notech_or2 i_50154807(.A(n_319431581), .B(n_55947), .Z(n_217082152));
	notech_or4 i_50254806(.A(n_55958), .B(n_2255), .C(n_28061), .D(n_60504),
		 .Z(n_217182153));
	notech_nao3 i_52654782(.A(n_62411), .B(opc[12]), .C(n_248534111), .Z(n_218182162
		));
	notech_or4 i_54554764(.A(n_57293), .B(n_55858), .C(n_56196), .D(n_59250)
		, .Z(n_219082171));
	notech_or4 i_80254523(.A(n_56172), .B(n_56081), .C(n_56369), .D(n_27592)
		, .Z(n_219882179));
	notech_ao4 i_188653474(.A(n_121523202), .B(n_322231609), .C(n_121723204)
		, .D(n_251061538), .Z(n_219982180));
	notech_ao4 i_188553475(.A(n_57334), .B(n_353365822), .C(n_353165820), .D
		(n_29137), .Z(n_220182182));
	notech_and3 i_188853472(.A(n_219882179), .B(n_219982180), .C(n_220182182
		), .Z(n_220282183));
	notech_ao4 i_188253477(.A(n_353265821), .B(n_56847), .C(n_56207), .D(n_26572
		), .Z(n_220382184));
	notech_ao4 i_188153478(.A(n_27546), .B(n_59791), .C(n_121623203), .D(n_59086
		), .Z(n_220482185));
	notech_ao4 i_167353685(.A(n_248534111), .B(n_177164109), .C(n_2326), .D(n_177264110
		), .Z(n_220782187));
	notech_ao4 i_167253686(.A(n_55727), .B(n_27581), .C(n_202067840), .D(n_27534
		), .Z(n_220982189));
	notech_and3 i_167553683(.A(n_219082171), .B(n_220782187), .C(n_220982189
		), .Z(n_221082190));
	notech_ao4 i_167053688(.A(n_55310), .B(n_55578), .C(n_26548), .D(nbus_11273
		[15]), .Z(n_221182191));
	notech_ao4 i_166953689(.A(n_55354), .B(n_29087), .C(n_356476400), .D(n_55156
		), .Z(n_221282192));
	notech_ao4 i_165953699(.A(n_2326), .B(n_169057978), .C(n_55947), .D(n_189074758
		), .Z(n_221482194));
	notech_ao4 i_165853700(.A(n_55727), .B(n_27577), .C(n_58514), .D(n_27531
		), .Z(n_221782196));
	notech_and3 i_166153697(.A(n_221482194), .B(n_221782196), .C(n_218182162
		), .Z(n_221882197));
	notech_ao4 i_165653702(.A(n_55310), .B(n_55542), .C(n_56739), .D(n_26548
		), .Z(n_221982198));
	notech_ao4 i_165553703(.A(n_55354), .B(n_29084), .C(n_55156), .D(n_57346
		), .Z(n_222082199));
	notech_ao4 i_163853720(.A(n_58514), .B(n_27529), .C(n_54822), .D(n_55450
		), .Z(n_222682204));
	notech_and4 i_164153717(.A(n_216982151), .B(n_222682204), .C(n_217082152
		), .D(n_217182153), .Z(n_222782205));
	notech_ao4 i_163653722(.A(n_55438), .B(n_317783152), .C(n_317883153), .D
		(n_56721), .Z(n_222882206));
	notech_ao4 i_163553723(.A(n_317683151), .B(n_29077), .C(n_57348), .D(n_55156
		), .Z(n_222982207));
	notech_ao4 i_142453924(.A(n_177164109), .B(n_333569134), .C(n_177264110)
		, .D(n_333669135), .Z(n_223182209));
	notech_ao4 i_142353925(.A(n_54946), .B(n_56766), .C(n_55725), .D(n_27581
		), .Z(n_223382211));
	notech_and3 i_142653922(.A(n_216282144), .B(n_223182209), .C(n_223382211
		), .Z(n_223482212));
	notech_ao4 i_142153927(.A(n_356476400), .B(n_54852), .C(n_54945), .D(\nbus_11276[15] 
		), .Z(n_223582213));
	notech_nand2 i_5349109(.A(rep_en5), .B(n_26445), .Z(n_223982217));
	notech_or2 i_5649106(.A(n_224182219), .B(n_55018), .Z(n_224082218));
	notech_and4 i_1049148(.A(n_271488741), .B(n_57430), .C(n_223982217), .D(n_270488749
		), .Z(n_224182219));
	notech_and2 i_949149(.A(n_224082218), .B(n_55637), .Z(n_224382221));
	notech_ao4 i_47643(.A(n_29123), .B(n_224382221), .C(n_55640), .D(n_271039498
		), .Z(\nbus_11286[0] ));
	notech_or4 i_140947828(.A(n_244656264), .B(n_1844), .C(n_59936), .D(n_59023
		), .Z(n_224482222));
	notech_nand3 i_2616835(.A(n_238282357), .B(n_238182356), .C(n_238882363)
		, .Z(n_9832));
	notech_or4 i_144647792(.A(n_244656264), .B(n_1844), .C(n_59936), .D(n_59041
		), .Z(n_225382231));
	notech_nand3 i_2416833(.A(n_239082365), .B(n_238982364), .C(n_239682371)
		, .Z(n_9822));
	notech_or4 i_146747774(.A(n_244656264), .B(n_1844), .C(n_59935), .D(n_59032
		), .Z(n_226382240));
	notech_nand3 i_2316832(.A(n_239882373), .B(n_239782372), .C(n_240482379)
		, .Z(n_9817));
	notech_or4 i_148647756(.A(n_244656264), .B(n_1844), .C(n_59935), .D(n_58996
		), .Z(n_227382249));
	notech_nand3 i_2216831(.A(n_240682381), .B(n_240582380), .C(n_241282387)
		, .Z(n_9812));
	notech_or4 i_150447738(.A(n_57383), .B(n_57404), .C(n_59889), .D(n_59005
		), .Z(n_228282258));
	notech_nand3 i_2116830(.A(n_241482389), .B(n_241382388), .C(n_242082395)
		, .Z(n_9807));
	notech_or4 i_152347720(.A(n_57383), .B(n_57404), .C(n_59889), .D(n_59014
		), .Z(n_229182267));
	notech_nand3 i_2016829(.A(n_242282397), .B(n_242182396), .C(n_242882403)
		, .Z(n_9802));
	notech_or4 i_154247702(.A(n_57383), .B(n_57404), .C(n_59885), .D(n_58969
		), .Z(n_230082276));
	notech_nand3 i_1916828(.A(n_243082405), .B(n_242982404), .C(n_243682411)
		, .Z(n_9797));
	notech_or4 i_156047684(.A(n_57383), .B(n_57404), .C(n_59885), .D(n_58978
		), .Z(n_230982285));
	notech_nand3 i_1816827(.A(n_243882413), .B(n_243782412), .C(n_244482419)
		, .Z(n_9792));
	notech_nand3 i_159747648(.A(n_55159), .B(n_59791), .C(mul64[31]), .Z(n_231982294
		));
	notech_or4 i_160847637(.A(n_57445), .B(n_59791), .C(n_2792), .D(n_27554)
		, .Z(n_233082305));
	notech_nand3 i_1616825(.A(n_244582420), .B(n_245582430), .C(n_244782422)
		, .Z(n_9782));
	notech_nand3 i_162147624(.A(n_55159), .B(n_59791), .C(mul64[30]), .Z(n_233182306
		));
	notech_or4 i_163247613(.A(n_57445), .B(n_59791), .C(n_2792), .D(n_27553)
		, .Z(n_234282317));
	notech_nand3 i_1516824(.A(n_245682431), .B(n_246682441), .C(n_245882433)
		, .Z(n_9777));
	notech_or4 i_167147576(.A(n_57445), .B(n_59791), .C(n_2792), .D(n_27551)
		, .Z(n_234382318));
	notech_nand2 i_168347565(.A(\opc_5[12] ), .B(n_26596), .Z(n_235482329)
		);
	notech_nand3 i_1316822(.A(n_246782442), .B(n_247782452), .C(n_246982444)
		, .Z(n_9767));
	notech_or4 i_169847552(.A(n_57445), .B(n_59791), .C(n_2792), .D(n_27550)
		, .Z(n_235582330));
	notech_nand2 i_171147541(.A(\opc_5[11] ), .B(n_26596), .Z(n_236682341)
		);
	notech_nand3 i_1216821(.A(n_247882453), .B(n_248882463), .C(n_248082455)
		, .Z(n_9762));
	notech_or4 i_175047504(.A(n_57445), .B(n_59795), .C(n_2792), .D(n_27548)
		, .Z(n_236782342));
	notech_nand2 i_176147493(.A(\opc_5[9] ), .B(n_26596), .Z(n_237882353));
	notech_nand3 i_1016819(.A(n_248982464), .B(n_249982474), .C(n_249182466)
		, .Z(n_9752));
	notech_ao4 i_142147817(.A(n_2313), .B(n_28925), .C(n_2314), .D(n_59346),
		 .Z(n_238182356));
	notech_ao4 i_142247816(.A(n_2248), .B(nbus_11348[25]), .C(n_2247), .D(n_29602
		), .Z(n_238282357));
	notech_ao4 i_142347815(.A(n_2249), .B(n_29603), .C(n_56627), .D(n_29464)
		, .Z(n_238482359));
	notech_ao4 i_142047818(.A(n_231547139), .B(nbus_11326[1]), .C(n_55009), 
		.D(n_28076), .Z(n_238682361));
	notech_and4 i_142647812(.A(n_2312), .B(n_238682361), .C(n_238482359), .D
		(n_224482222), .Z(n_238882363));
	notech_ao4 i_146047781(.A(n_2313), .B(n_28923), .C(n_2314), .D(n_59319),
		 .Z(n_238982364));
	notech_ao4 i_146147780(.A(n_2248), .B(nbus_11348[23]), .C(n_2247), .D(n_29604
		), .Z(n_239082365));
	notech_ao4 i_146247779(.A(n_2249), .B(n_29605), .C(n_56627), .D(n_29465)
		, .Z(n_239282367));
	notech_ao4 i_145947782(.A(n_231547139), .B(nbus_11326[15]), .C(n_55009),
		 .D(n_28074), .Z(n_239482369));
	notech_and4 i_146547776(.A(n_2312), .B(n_239482369), .C(n_239282367), .D
		(n_225382231), .Z(n_239682371));
	notech_ao4 i_147847763(.A(n_2313), .B(n_28922), .C(n_2314), .D(n_55647),
		 .Z(n_239782372));
	notech_ao4 i_147947762(.A(n_2248), .B(nbus_11348[22]), .C(n_2247), .D(n_29606
		), .Z(n_239882373));
	notech_ao4 i_148047761(.A(n_2249), .B(n_29607), .C(n_56627), .D(n_29470)
		, .Z(n_240082375));
	notech_ao4 i_147747764(.A(n_231547139), .B(nbus_11326[14]), .C(n_55009),
		 .D(n_28073), .Z(n_240282377));
	notech_and4 i_148347758(.A(n_2312), .B(n_240282377), .C(n_240082375), .D
		(n_226382240), .Z(n_240482379));
	notech_ao4 i_149747745(.A(n_2313), .B(n_28921), .C(n_2314), .D(n_59310),
		 .Z(n_240582380));
	notech_ao4 i_149847744(.A(n_2248), .B(nbus_11348[21]), .C(n_2247), .D(n_29608
		), .Z(n_240682381));
	notech_ao4 i_149947743(.A(n_2249), .B(n_29609), .C(n_56631), .D(n_29471)
		, .Z(n_240882383));
	notech_ao4 i_149647746(.A(n_231547139), .B(nbus_11326[13]), .C(n_55009),
		 .D(n_28072), .Z(n_241082385));
	notech_and4 i_150247740(.A(n_2312), .B(n_241082385), .C(n_240882383), .D
		(n_227382249), .Z(n_241282387));
	notech_ao4 i_151547727(.A(n_2313), .B(n_28920), .C(n_2314), .D(n_55631),
		 .Z(n_241382388));
	notech_ao4 i_151647726(.A(n_2248), .B(nbus_11348[20]), .C(n_2247), .D(n_29610
		), .Z(n_241482389));
	notech_ao4 i_151747725(.A(n_2249), .B(n_29611), .C(n_56631), .D(n_29472)
		, .Z(n_241682391));
	notech_ao4 i_151447728(.A(n_231547139), .B(nbus_11326[12]), .C(n_55009),
		 .D(n_28071), .Z(n_241882393));
	notech_and4 i_152147722(.A(n_2312), .B(n_241882393), .C(n_241682391), .D
		(n_228282258), .Z(n_242082395));
	notech_ao4 i_153547709(.A(n_2313), .B(n_28919), .C(n_2314), .D(n_55620),
		 .Z(n_242182396));
	notech_ao4 i_153647708(.A(n_2248), .B(nbus_11348[19]), .C(n_2247), .D(n_29612
		), .Z(n_242282397));
	notech_ao4 i_153747707(.A(n_2249), .B(n_29614), .C(n_56627), .D(n_29473)
		, .Z(n_242482399));
	notech_ao4 i_153447710(.A(n_231547139), .B(nbus_11326[11]), .C(n_55009),
		 .D(n_28070), .Z(n_242682401));
	notech_and4 i_154047704(.A(n_2312), .B(n_242682401), .C(n_242482399), .D
		(n_229182267), .Z(n_242882403));
	notech_ao4 i_155347691(.A(n_54887), .B(n_28918), .C(n_2314), .D(n_55609)
		, .Z(n_242982404));
	notech_ao4 i_155447690(.A(n_54926), .B(nbus_11348[18]), .C(n_54908), .D(n_29615
		), .Z(n_243082405));
	notech_ao4 i_155547689(.A(n_2249), .B(n_29616), .C(n_56627), .D(n_29475)
		, .Z(n_243282407));
	notech_ao4 i_155247692(.A(n_54847), .B(nbus_11326[10]), .C(n_54836), .D(n_28069
		), .Z(n_243482409));
	notech_and4 i_155847686(.A(n_2312), .B(n_243482409), .C(n_243282407), .D
		(n_230082276), .Z(n_243682411));
	notech_ao4 i_157247673(.A(n_54887), .B(n_28917), .C(n_54863), .D(n_55600
		), .Z(n_243782412));
	notech_ao4 i_157347672(.A(n_54926), .B(nbus_11348[17]), .C(n_54908), .D(n_29617
		), .Z(n_243882413));
	notech_ao4 i_157447671(.A(n_54940), .B(n_29618), .C(n_56627), .D(n_29476
		), .Z(n_244082415));
	notech_ao4 i_157147674(.A(n_54847), .B(nbus_11326[9]), .C(n_54836), .D(n_28068
		), .Z(n_244282417));
	notech_and4 i_157747668(.A(n_2312), .B(n_244282417), .C(n_244082415), .D
		(n_230982285), .Z(n_244482419));
	notech_ao4 i_161447631(.A(n_55111), .B(n_59095), .C(n_54940), .D(n_29621
		), .Z(n_244582420));
	notech_and4 i_161547630(.A(n_57312), .B(n_2186), .C(n_231982294), .D(n_233082305
		), .Z(n_244782422));
	notech_ao4 i_161047635(.A(n_54836), .B(n_28066), .C(n_55122), .D(n_55400
		), .Z(n_244982424));
	notech_ao4 i_161147634(.A(n_54863), .B(n_55578), .C(n_54847), .D(n_59041
		), .Z(n_245082425));
	notech_ao4 i_161247633(.A(n_54908), .B(n_29619), .C(n_54887), .D(n_28915
		), .Z(n_245282427));
	notech_ao4 i_161347632(.A(n_56627), .B(n_29477), .C(n_54926), .D(nbus_11348
		[15]), .Z(n_245382428));
	notech_and4 i_161947626(.A(n_245382428), .B(n_245282427), .C(n_245082425
		), .D(n_244982424), .Z(n_245582430));
	notech_ao4 i_163847607(.A(n_55111), .B(n_59050), .C(n_54940), .D(n_29623
		), .Z(n_245682431));
	notech_and4 i_163947606(.A(n_57312), .B(n_2186), .C(n_233182306), .D(n_234282317
		), .Z(n_245882433));
	notech_ao4 i_163447611(.A(n_54836), .B(n_28065), .C(n_55122), .D(n_55387
		), .Z(n_246082435));
	notech_ao4 i_163547610(.A(n_54863), .B(n_55566), .C(n_54847), .D(n_59032
		), .Z(n_246182436));
	notech_ao4 i_163647609(.A(n_54908), .B(n_29622), .C(n_54887), .D(n_28914
		), .Z(n_246382438));
	notech_ao4 i_163747608(.A(n_56627), .B(n_29478), .C(n_54926), .D(nbus_11348
		[14]), .Z(n_246482439));
	notech_and4 i_164347602(.A(n_246482439), .B(n_246382438), .C(n_246182436
		), .D(n_246082435), .Z(n_246682441));
	notech_ao4 i_168947559(.A(n_56627), .B(n_29479), .C(n_54926), .D(nbus_11348
		[12]), .Z(n_246782442));
	notech_and4 i_169147558(.A(n_57312), .B(n_2186), .C(n_234382318), .D(n_235482329
		), .Z(n_246982444));
	notech_ao4 i_168547563(.A(n_55111), .B(n_59077), .C(n_2311), .D(n_29343)
		, .Z(n_247182446));
	notech_ao4 i_168647562(.A(n_54836), .B(n_28063), .C(n_55122), .D(n_55365
		), .Z(n_247282447));
	notech_ao4 i_168747561(.A(n_54863), .B(n_55542), .C(n_54847), .D(n_59005
		), .Z(n_247482449));
	notech_ao4 i_168847560(.A(n_54908), .B(n_29624), .C(n_54887), .D(n_28912
		), .Z(n_247582450));
	notech_and4 i_169547554(.A(n_247582450), .B(n_247482449), .C(n_247282447
		), .D(n_247182446), .Z(n_247782452));
	notech_ao4 i_171747535(.A(n_56631), .B(n_29480), .C(n_54926), .D(nbus_11348
		[11]), .Z(n_247882453));
	notech_and4 i_171847534(.A(n_57312), .B(n_2186), .C(n_235582330), .D(n_236682341
		), .Z(n_248082455));
	notech_ao4 i_171347539(.A(n_55111), .B(n_59059), .C(n_2311), .D(n_29341)
		, .Z(n_248282457));
	notech_ao4 i_171447538(.A(n_54836), .B(n_28062), .C(n_55122), .D(n_55277
		), .Z(n_248382458));
	notech_ao4 i_171547537(.A(n_54863), .B(n_55469), .C(n_54847), .D(n_59014
		), .Z(n_248582460));
	notech_ao4 i_171647536(.A(n_54908), .B(n_29625), .C(n_54887), .D(n_28911
		), .Z(n_248682461));
	notech_and4 i_172247530(.A(n_248682461), .B(n_248582460), .C(n_248382458
		), .D(n_248282457), .Z(n_248882463));
	notech_ao4 i_176747487(.A(n_56631), .B(n_29481), .C(n_54926), .D(nbus_11348
		[9]), .Z(n_248982464));
	notech_and4 i_176847486(.A(n_57312), .B(n_2186), .C(n_236782342), .D(n_237882353
		), .Z(n_249182466));
	notech_ao4 i_176347491(.A(n_55111), .B(n_59023), .C(n_2311), .D(n_29337)
		, .Z(n_249382468));
	notech_ao4 i_176447490(.A(n_54836), .B(n_28060), .C(n_55122), .D(\nbus_11276[1] 
		), .Z(n_249482469));
	notech_ao4 i_176547489(.A(n_54863), .B(n_55425), .C(n_54847), .D(n_58978
		), .Z(n_249682471));
	notech_ao4 i_176647488(.A(n_54908), .B(n_29628), .C(n_54887), .D(n_28909
		), .Z(n_249782472));
	notech_and4 i_177347482(.A(n_249782472), .B(n_249682471), .C(n_249482469
		), .D(n_249382468), .Z(n_249982474));
	notech_nand3 i_7845299(.A(n_54128), .B(tsc[25]), .C(n_59800), .Z(n_250282477
		));
	notech_nand2 i_7745300(.A(opc[25]), .B(n_351965808), .Z(n_250582480));
	notech_or4 i_7245305(.A(n_58656), .B(n_56114), .C(n_55798), .D(n_308421971
		), .Z(n_251082485));
	notech_nand3 i_8745290(.A(n_54128), .B(tsc[26]), .C(n_59800), .Z(n_251182486
		));
	notech_nand2 i_8645291(.A(n_351965808), .B(opc[26]), .Z(n_251482489));
	notech_or4 i_8145296(.A(n_58656), .B(n_56114), .C(n_55798), .D(n_308321970
		), .Z(n_251982494));
	notech_nand3 i_10545272(.A(tsc[28]), .B(n_59800), .C(n_54128), .Z(n_252082495
		));
	notech_nand2 i_10445273(.A(n_351965808), .B(opc[28]), .Z(n_252382498));
	notech_or2 i_9945278(.A(n_54148), .B(n_55261), .Z(n_252882503));
	notech_or4 i_17045207(.A(n_2740), .B(n_2213), .C(n_59230), .D(n_28605), 
		.Z(n_253382508));
	notech_or2 i_16745210(.A(n_55192), .B(n_59041), .Z(n_253682511));
	notech_nand2 i_18245195(.A(resb_shiftbox[25]), .B(n_26578), .Z(n_254582520
		));
	notech_nand3 i_17945198(.A(n_1969), .B(nbus_137[25]), .C(n_59800), .Z(n_254882523
		));
	notech_or4 i_19445183(.A(n_2740), .B(n_2213), .C(n_59230), .D(n_28602), 
		.Z(n_255782532));
	notech_or2 i_19145186(.A(n_55192), .B(n_59068), .Z(n_256082535));
	notech_or4 i_20645171(.A(n_2740), .B(n_2213), .C(n_59230), .D(n_28600), 
		.Z(n_256982544));
	notech_or2 i_20345174(.A(n_55192), .B(n_59059), .Z(n_257282547));
	notech_nand2 i_21845159(.A(resb_shiftbox[28]), .B(n_26578), .Z(n_258182556
		));
	notech_nand3 i_21545162(.A(n_1969), .B(nbus_137[28]), .C(n_59800), .Z(n_258482559
		));
	notech_or2 i_23045147(.A(n_55170), .B(n_56892), .Z(n_259382568));
	notech_or2 i_22745150(.A(n_55243), .B(n_27552), .Z(n_259682571));
	notech_or2 i_31245068(.A(n_55347), .B(n_29215), .Z(n_260182576));
	notech_or2 i_31545065(.A(n_304021927), .B(n_55888), .Z(n_261482589));
	notech_or2 i_32645054(.A(n_55347), .B(n_29154), .Z(n_261582590));
	notech_or2 i_32945051(.A(n_304221929), .B(n_55888), .Z(n_262882603));
	notech_or2 i_68944702(.A(n_308921976), .B(n_353365822), .Z(n_266882643)
		);
	notech_nor2 i_70244689(.A(n_121623203), .B(n_59023), .Z(n_266982644));
	notech_or4 i_69744694(.A(n_56172), .B(n_56081), .C(n_55798), .D(n_308421971
		), .Z(n_267682651));
	notech_nor2 i_71044681(.A(n_121623203), .B(n_59068), .Z(n_267782652));
	notech_or4 i_70544686(.A(n_56172), .B(n_56081), .C(n_55798), .D(n_308321970
		), .Z(n_268482659));
	notech_nor2 i_71844673(.A(n_121623203), .B(n_59059), .Z(n_268582660));
	notech_or4 i_71344678(.A(n_56172), .B(n_56081), .C(n_55798), .D(n_308221969
		), .Z(n_269282667));
	notech_nor2 i_72644665(.A(n_121623203), .B(n_59077), .Z(n_269382668));
	notech_or2 i_72144670(.A(n_55402), .B(n_57330), .Z(n_270082675));
	notech_ao4 i_176443668(.A(n_55403), .B(n_29219), .C(n_56043), .D(n_307421961
		), .Z(n_270182676));
	notech_ao4 i_176343669(.A(n_322088470), .B(n_55261), .C(n_97522962), .D(n_56883
		), .Z(n_270382678));
	notech_nand3 i_176643666(.A(n_270182676), .B(n_270382678), .C(n_270082675
		), .Z(n_270482679));
	notech_ao4 i_176143671(.A(n_343565725), .B(n_121723204), .C(n_121523202)
		, .D(n_57306), .Z(n_270582680));
	notech_ao4 i_175743675(.A(n_286061878), .B(n_121723204), .C(n_56043), .D
		(n_303621923), .Z(n_270882683));
	notech_ao4 i_175643676(.A(n_55403), .B(n_29154), .C(n_55402), .D(n_308621973
		), .Z(n_271082685));
	notech_nand3 i_175943673(.A(n_270882683), .B(n_271082685), .C(n_269282667
		), .Z(n_271182686));
	notech_ao4 i_175443678(.A(n_322088470), .B(n_59328), .C(n_97522962), .D(n_56874
		), .Z(n_271282687));
	notech_ao4 i_175043682(.A(n_288561889), .B(n_121723204), .C(n_56043), .D
		(n_307621963), .Z(n_271582690));
	notech_ao4 i_174943683(.A(n_55403), .B(n_29156), .C(n_55402), .D(n_308721974
		), .Z(n_271782692));
	notech_nand3 i_175243680(.A(n_271582690), .B(n_271782692), .C(n_268482659
		), .Z(n_271882693));
	notech_ao4 i_174743685(.A(n_322088470), .B(n_59337), .C(n_97522962), .D(n_56865
		), .Z(n_271982694));
	notech_ao4 i_174343689(.A(n_268264999), .B(n_121723204), .C(n_56043), .D
		(n_307521962), .Z(n_272282697));
	notech_ao4 i_174243690(.A(n_55403), .B(n_29215), .C(n_308821975), .D(n_55402
		), .Z(n_272482699));
	notech_nand3 i_174543687(.A(n_272282697), .B(n_272482699), .C(n_267682651
		), .Z(n_272582700));
	notech_ao4 i_174043692(.A(n_322088470), .B(n_59346), .C(n_97522962), .D(n_56856
		), .Z(n_272682701));
	notech_ao4 i_173643696(.A(n_121523202), .B(n_308521972), .C(n_121723204)
		, .D(n_270765024), .Z(n_272982704));
	notech_ao4 i_173543697(.A(n_353165820), .B(n_29152), .C(n_27590), .D(n_353465823
		), .Z(n_273182706));
	notech_and3 i_173843694(.A(n_272982704), .B(n_273182706), .C(n_266882643
		), .Z(n_273282707));
	notech_ao4 i_173343699(.A(n_353265821), .B(n_56838), .C(\nbus_11276[23] 
		), .D(n_26572), .Z(n_273382708));
	notech_ao4 i_173243700(.A(n_27545), .B(n_59800), .C(n_121623203), .D(nbus_11326
		[23]), .Z(n_273482709));
	notech_ao4 i_160943822(.A(n_304221929), .B(n_55947), .C(n_302721914), .D
		(n_343565725), .Z(n_273682711));
	notech_ao4 i_160843823(.A(n_55269), .B(n_57330), .C(n_55447), .D(n_55261
		), .Z(n_273782712));
	notech_ao4 i_160643825(.A(n_58514), .B(n_27551), .C(n_55267), .D(n_29219
		), .Z(n_273982714));
	notech_ao4 i_160543826(.A(n_113313527), .B(n_59077), .C(n_55562), .D(n_56883
		), .Z(n_274082715));
	notech_ao4 i_160343828(.A(n_55947), .B(n_304121928), .C(n_302721914), .D
		(n_286061878), .Z(n_274282717));
	notech_ao4 i_160243829(.A(n_55447), .B(n_59328), .C(n_55269), .D(n_308621973
		), .Z(n_274382718));
	notech_ao4 i_160043831(.A(n_58514), .B(n_27550), .C(n_55267), .D(n_29154
		), .Z(n_274582720));
	notech_ao4 i_159943832(.A(n_113313527), .B(n_59059), .C(n_55562), .D(n_56874
		), .Z(n_274682721));
	notech_ao4 i_159743834(.A(n_304021927), .B(n_55947), .C(n_302721914), .D
		(n_288561889), .Z(n_274882723));
	notech_ao4 i_159643835(.A(n_55447), .B(n_59337), .C(n_55269), .D(n_308721974
		), .Z(n_274982724));
	notech_ao4 i_159443837(.A(n_58514), .B(n_27549), .C(n_55267), .D(n_29156
		), .Z(n_275182726));
	notech_ao4 i_159343838(.A(n_113313527), .B(n_59068), .C(n_55562), .D(n_56865
		), .Z(n_275282727));
	notech_ao4 i_159143840(.A(n_55947), .B(n_303921926), .C(n_268264999), .D
		(n_302721914), .Z(n_275482729));
	notech_ao4 i_159043841(.A(n_55447), .B(n_59346), .C(n_308821975), .D(n_55269
		), .Z(n_275582730));
	notech_ao4 i_158543843(.A(n_58514), .B(n_27548), .C(n_55267), .D(n_29215
		), .Z(n_275782732));
	notech_ao4 i_158443844(.A(n_113313527), .B(n_59023), .C(n_55562), .D(n_56856
		), .Z(n_275882733));
	notech_ao4 i_143043990(.A(n_303421921), .B(n_59077), .C(n_343565725), .D
		(n_302621913), .Z(n_276082735));
	notech_ao4 i_142943991(.A(n_55221), .B(\nbus_11276[28] ), .C(n_55220), .D
		(n_56883), .Z(n_276282737));
	notech_ao4 i_142743993(.A(n_55346), .B(n_57330), .C(n_55347), .D(n_29219
		), .Z(n_276482739));
	notech_and3 i_142843992(.A(n_53844), .B(n_276482739), .C(n_26249), .Z(n_276682741
		));
	notech_ao4 i_142443996(.A(n_303421921), .B(n_59059), .C(n_286061878), .D
		(n_302621913), .Z(n_276782742));
	notech_ao4 i_142343997(.A(n_55346), .B(n_308621973), .C(n_55888), .D(n_304121928
		), .Z(n_276882743));
	notech_ao4 i_142143999(.A(n_55221), .B(n_59328), .C(n_55220), .D(n_56874
		), .Z(n_277082745));
	notech_ao3 i_142243998(.A(n_277082745), .B(n_261582590), .C(n_264975488)
		, .Z(n_277282747));
	notech_ao4 i_141744003(.A(n_303421921), .B(nbus_11326[26]), .C(n_288561889
		), .D(n_302621913), .Z(n_277382748));
	notech_ao4 i_141644004(.A(n_55220), .B(n_56865), .C(n_55346), .D(n_308721974
		), .Z(n_277582750));
	notech_ao4 i_141444006(.A(n_55347), .B(n_29156), .C(n_55221), .D(n_59337
		), .Z(n_277782752));
	notech_and3 i_141544005(.A(n_53844), .B(n_277782752), .C(n_26413), .Z(n_277982754
		));
	notech_ao4 i_141144009(.A(n_303421921), .B(n_59023), .C(n_268264999), .D
		(n_302621913), .Z(n_278082755));
	notech_ao4 i_141044010(.A(n_55346), .B(n_308821975), .C(n_55893), .D(n_303921926
		), .Z(n_278182756));
	notech_ao4 i_140844012(.A(n_55221), .B(n_59346), .C(n_55220), .D(n_56856
		), .Z(n_278382758));
	notech_and3 i_140944011(.A(n_278382758), .B(n_26308), .C(n_260182576), .Z
		(n_278582760));
	notech_ao4 i_129644123(.A(n_2318), .B(n_28853), .C(n_55075), .D(n_57329)
		, .Z(n_278682761));
	notech_ao4 i_129544124(.A(n_55619), .B(n_28640), .C(n_55933), .D(n_55249
		), .Z(n_278782762));
	notech_ao4 i_129344126(.A(n_55102), .B(n_28798), .C(n_55526), .D(n_28598
		), .Z(n_278982764));
	notech_and4 i_129844121(.A(n_278982764), .B(n_278782762), .C(n_278682761
		), .D(n_259682571), .Z(n_279182766));
	notech_ao4 i_128944129(.A(n_55181), .B(n_29025), .C(n_55192), .D(n_59104
		), .Z(n_279282767));
	notech_ao4 i_128744131(.A(n_55136), .B(n_27597), .C(n_55161), .D(n_28829
		), .Z(n_279482769));
	notech_and4 i_129244127(.A(n_2187), .B(n_279482769), .C(n_279282767), .D
		(n_259382568), .Z(n_279682771));
	notech_ao4 i_128444134(.A(n_55204), .B(n_27551), .C(n_55075), .D(n_57330
		), .Z(n_279782772));
	notech_ao4 i_128344135(.A(n_55170), .B(n_56883), .C(n_55933), .D(n_55261
		), .Z(n_279882773));
	notech_ao4 i_128144137(.A(n_55136), .B(n_27596), .C(n_55192), .D(n_59077
		), .Z(n_280082775));
	notech_and4 i_128644132(.A(n_280082775), .B(n_279882773), .C(n_279782772
		), .D(n_258482559), .Z(n_280282777));
	notech_ao4 i_127844140(.A(n_55526), .B(n_28599), .C(n_55091), .D(n_28639
		), .Z(n_280382778));
	notech_ao4 i_127644142(.A(n_55161), .B(n_28828), .C(n_55181), .D(n_29033
		), .Z(n_280582780));
	notech_and4 i_128044138(.A(n_2187), .B(n_280582780), .C(n_280382778), .D
		(n_258182556), .Z(n_280782782));
	notech_ao4 i_127344145(.A(n_55181), .B(n_29016), .C(n_308621973), .D(n_55075
		), .Z(n_280882783));
	notech_ao4 i_127244146(.A(n_55204), .B(n_27550), .C(n_55136), .D(n_27595
		), .Z(n_280982784));
	notech_ao4 i_127044148(.A(n_55170), .B(n_56874), .C(n_55933), .D(\nbus_11276[27] 
		), .Z(n_281182786));
	notech_and4 i_127544143(.A(n_281182786), .B(n_280982784), .C(n_280882783
		), .D(n_257282547), .Z(n_281382788));
	notech_ao4 i_126744151(.A(n_55091), .B(n_28638), .C(n_2318), .D(n_28852)
		, .Z(n_281482789));
	notech_ao4 i_126544153(.A(n_55161), .B(n_28827), .C(n_55102), .D(n_28797
		), .Z(n_281682791));
	notech_and4 i_126944149(.A(n_2187), .B(n_281682791), .C(n_281482789), .D
		(n_256982544), .Z(n_281882793));
	notech_ao4 i_126244156(.A(n_55181), .B(n_29013), .C(n_55075), .D(n_308721974
		), .Z(n_281982794));
	notech_ao4 i_126144157(.A(n_55204), .B(n_27549), .C(n_55136), .D(n_27594
		), .Z(n_282082795));
	notech_ao4 i_125944159(.A(n_55170), .B(n_56865), .C(n_55933), .D(\nbus_11276[26] 
		), .Z(n_282282797));
	notech_and4 i_126444154(.A(n_282282797), .B(n_282082795), .C(n_281982794
		), .D(n_256082535), .Z(n_282482799));
	notech_ao4 i_125644162(.A(n_55091), .B(n_28637), .C(n_2318), .D(n_28851)
		, .Z(n_282582800));
	notech_ao4 i_125444164(.A(n_55161), .B(n_28826), .C(n_55102), .D(n_28796
		), .Z(n_282782802));
	notech_and4 i_125844160(.A(n_2187), .B(n_282782802), .C(n_282582800), .D
		(n_255782532), .Z(n_282982804));
	notech_ao4 i_125144167(.A(n_55136), .B(n_27593), .C(n_55075), .D(n_308821975
		), .Z(n_283082805));
	notech_ao4 i_125044168(.A(n_55933), .B(\nbus_11276[25] ), .C(n_55204), .D
		(n_27548), .Z(n_283182806));
	notech_ao4 i_124844170(.A(n_55192), .B(nbus_11326[25]), .C(n_55170), .D(n_56856
		), .Z(n_283382808));
	notech_and4 i_125344165(.A(n_283382808), .B(n_283182806), .C(n_283082805
		), .D(n_254882523), .Z(n_283582810));
	notech_ao4 i_124544173(.A(n_55526), .B(n_28603), .C(n_55091), .D(n_28636
		), .Z(n_283682811));
	notech_ao4 i_124344175(.A(n_55161), .B(n_28825), .C(n_55181), .D(n_29022
		), .Z(n_283882813));
	notech_and4 i_124744171(.A(n_2187), .B(n_283882813), .C(n_283682811), .D
		(n_254582520), .Z(n_284082815));
	notech_ao4 i_124044178(.A(n_55181), .B(n_29030), .C(n_308921976), .D(n_55075
		), .Z(n_284182816));
	notech_ao4 i_123944179(.A(n_55204), .B(n_27545), .C(n_55136), .D(n_27590
		), .Z(n_284282817));
	notech_ao4 i_123744181(.A(n_55170), .B(n_56838), .C(n_55933), .D(n_59319
		), .Z(n_284482819));
	notech_and4 i_124244176(.A(n_284482819), .B(n_284282817), .C(n_284182816
		), .D(n_253682511), .Z(n_284682821));
	notech_ao4 i_123444184(.A(n_55091), .B(n_28634), .C(n_2318), .D(n_28850)
		, .Z(n_284782822));
	notech_ao4 i_123244186(.A(n_55161), .B(n_28823), .C(n_55102), .D(n_28794
		), .Z(n_284982824));
	notech_and4 i_123644182(.A(n_2187), .B(n_284982824), .C(n_284782822), .D
		(n_253382508), .Z(n_285182826));
	notech_ao4 i_118244236(.A(n_57330), .B(n_352165810), .C(n_56023), .D(n_307421961
		), .Z(n_285282827));
	notech_ao4 i_118144237(.A(n_29219), .B(n_26565), .C(n_55143), .D(n_56883
		), .Z(n_285482829));
	notech_ao4 i_117844240(.A(n_343565725), .B(n_352965818), .C(n_57306), .D
		(n_352365812), .Z(n_285682831));
	notech_and4 i_118044238(.A(n_285682831), .B(n_252082495), .C(n_252382498
		), .D(n_26249), .Z(n_285982834));
	notech_ao4 i_116644252(.A(n_288561889), .B(n_352965818), .C(n_307621963)
		, .D(n_56023), .Z(n_286082835));
	notech_ao4 i_116544253(.A(n_29156), .B(n_26565), .C(n_308721974), .D(n_352165810
		), .Z(n_286282837));
	notech_ao4 i_116244256(.A(n_55143), .B(n_56865), .C(n_54148), .D(n_59337
		), .Z(n_286482839));
	notech_and4 i_116444254(.A(n_286482839), .B(n_251182486), .C(n_251482489
		), .D(n_26413), .Z(n_286782842));
	notech_ao4 i_115844260(.A(n_268264999), .B(n_352965818), .C(n_307521962)
		, .D(n_56023), .Z(n_286882843));
	notech_ao4 i_115744261(.A(n_29215), .B(n_26565), .C(n_308821975), .D(n_352165810
		), .Z(n_287082845));
	notech_ao4 i_115444264(.A(n_55143), .B(n_56856), .C(n_54148), .D(n_59346
		), .Z(n_287282847));
	notech_and4 i_115644262(.A(n_287282847), .B(n_250282477), .C(n_250582480
		), .D(n_26308), .Z(n_287582850));
	notech_nand2 i_13042112(.A(resb_shiftbox[18]), .B(n_26578), .Z(n_288082855
		));
	notech_nand3 i_12742115(.A(n_1969), .B(nbus_137[18]), .C(n_59800), .Z(n_288382858
		));
	notech_or4 i_14242100(.A(n_2740), .B(n_2213), .C(n_59230), .D(n_28609), 
		.Z(n_289282867));
	notech_or2 i_13942103(.A(n_55192), .B(n_59014), .Z(n_289582870));
	notech_nand2 i_15442088(.A(resb_shiftbox[20]), .B(n_26578), .Z(n_290482879
		));
	notech_nand3 i_15142091(.A(n_1969), .B(nbus_137[20]), .C(n_59800), .Z(n_290782882
		));
	notech_or4 i_16642076(.A(n_2740), .B(n_2213), .C(n_59230), .D(n_28607), 
		.Z(n_291682891));
	notech_or2 i_16342079(.A(n_55192), .B(n_58996), .Z(n_291982894));
	notech_nand2 i_17842064(.A(resb_shiftbox[22]), .B(n_26578), .Z(n_292882903
		));
	notech_nand3 i_17542067(.A(nbus_137[22]), .B(n_1969), .C(n_59800), .Z(n_293182906
		));
	notech_or2 i_45941789(.A(n_354969318), .B(n_311318890), .Z(n_294482919)
		);
	notech_or2 i_46841780(.A(n_354969318), .B(n_311218889), .Z(n_295382928)
		);
	notech_or2 i_47741771(.A(n_354969318), .B(n_311118888), .Z(n_296282937)
		);
	notech_or2 i_65641596(.A(n_311218889), .B(n_353365822), .Z(n_297082945)
		);
	notech_or2 i_67241580(.A(n_311018887), .B(n_353365822), .Z(n_297882953)
		);
	notech_ao4 i_174540547(.A(n_310518882), .B(n_121523202), .C(n_121723204)
		, .D(n_312662130), .Z(n_297982954));
	notech_ao4 i_174440548(.A(n_353165820), .B(n_29172), .C(n_353465823), .D
		(n_27588), .Z(n_298182956));
	notech_and3 i_174740545(.A(n_297982954), .B(n_298182956), .C(n_297882953
		), .Z(n_298282957));
	notech_ao4 i_174240550(.A(n_353265821), .B(n_56820), .C(n_59310), .D(n_26572
		), .Z(n_298382958));
	notech_ao4 i_174140551(.A(n_27541), .B(n_59795), .C(n_121623203), .D(nbus_11326
		[21]), .Z(n_298482959));
	notech_ao4 i_173140561(.A(n_310718884), .B(n_121523202), .C(n_121723204)
		, .D(n_308065397), .Z(n_298682961));
	notech_ao4 i_173040562(.A(n_353165820), .B(n_29167), .C(n_353465823), .D
		(n_27585), .Z(n_298882963));
	notech_and3 i_173340559(.A(n_298682961), .B(n_298882963), .C(n_297082945
		), .Z(n_298982964));
	notech_ao4 i_172840564(.A(n_353265821), .B(n_56802), .C(n_55620), .D(n_26572
		), .Z(n_299082965));
	notech_ao4 i_172740565(.A(n_27539), .B(n_59795), .C(n_121623203), .D(n_59014
		), .Z(n_299182966));
	notech_ao4 i_157640709(.A(n_310618883), .B(n_354569315), .C(n_113113525)
		, .D(n_315162155), .Z(n_299382968));
	notech_ao4 i_157540710(.A(n_58514), .B(n_27540), .C(n_55776), .D(n_27586
		), .Z(n_299582970));
	notech_and3 i_157840707(.A(n_299382968), .B(n_299582970), .C(n_296282937
		), .Z(n_299682971));
	notech_ao4 i_157340712(.A(n_354669316), .B(n_55631), .C(n_29169), .D(n_26571
		), .Z(n_299782972));
	notech_ao4 i_157240713(.A(n_113313527), .B(n_59005), .C(n_55562), .D(n_56811
		), .Z(n_299882973));
	notech_ao4 i_156940716(.A(n_310718884), .B(n_354569315), .C(n_308065397)
		, .D(n_113113525), .Z(n_300082975));
	notech_ao4 i_156840717(.A(n_58514), .B(n_27539), .C(n_55776), .D(n_27585
		), .Z(n_300282977));
	notech_and3 i_157140714(.A(n_300082975), .B(n_300282977), .C(n_295382928
		), .Z(n_300382978));
	notech_ao4 i_156640719(.A(n_354669316), .B(n_55620), .C(n_29167), .D(n_26571
		), .Z(n_300482979));
	notech_ao4 i_156540720(.A(n_113313527), .B(nbus_11326[19]), .C(n_55562),
		 .D(n_56802), .Z(n_300582980));
	notech_ao4 i_156140723(.A(n_310818885), .B(n_354569315), .C(n_113113525)
		, .D(n_310565422), .Z(n_300782982));
	notech_ao4 i_156040724(.A(n_58514), .B(n_27538), .C(n_55776), .D(n_27584
		), .Z(n_300982984));
	notech_and3 i_156440721(.A(n_300782982), .B(n_300982984), .C(n_294482919
		), .Z(n_301082985));
	notech_ao4 i_155840726(.A(n_354669316), .B(n_55609), .C(n_29165), .D(n_26571
		), .Z(n_301182986));
	notech_ao4 i_155740727(.A(n_113313527), .B(n_58969), .C(n_55562), .D(n_56793
		), .Z(n_301282987));
	notech_ao4 i_125041025(.A(n_55136), .B(n_27589), .C(n_26618), .D(n_55075
		), .Z(n_301482989));
	notech_ao4 i_124941026(.A(n_55933), .B(n_55647), .C(n_55204), .D(n_27542
		), .Z(n_301582990));
	notech_ao4 i_124741028(.A(n_55192), .B(nbus_11326[22]), .C(n_55170), .D(n_56829
		), .Z(n_301782992));
	notech_and4 i_125241023(.A(n_301782992), .B(n_301582990), .C(n_301482989
		), .D(n_293182906), .Z(n_301982994));
	notech_ao4 i_124441031(.A(n_55526), .B(n_28606), .C(n_55091), .D(n_28633
		), .Z(n_302082995));
	notech_ao4 i_124241033(.A(n_55161), .B(n_28822), .C(n_55181), .D(n_28972
		), .Z(n_302282997));
	notech_and4 i_124641029(.A(n_2187), .B(n_302282997), .C(n_302082995), .D
		(n_292882903), .Z(n_302482999));
	notech_ao4 i_123941036(.A(n_55181), .B(n_29026), .C(n_311018887), .D(n_55075
		), .Z(n_302583000));
	notech_ao4 i_123841037(.A(n_55204), .B(n_27541), .C(n_55136), .D(n_27588
		), .Z(n_302683001));
	notech_ao4 i_123541039(.A(n_55170), .B(n_56820), .C(n_55933), .D(n_59310
		), .Z(n_302883003));
	notech_and4 i_124141034(.A(n_302883003), .B(n_302683001), .C(n_302583000
		), .D(n_291982894), .Z(n_303083005));
	notech_ao4 i_123241042(.A(n_55091), .B(n_28632), .C(n_2318), .D(n_28849)
		, .Z(n_303183006));
	notech_ao4 i_123041044(.A(n_55161), .B(n_28821), .C(n_55102), .D(n_28793
		), .Z(n_303383008));
	notech_and4 i_123441040(.A(n_2187), .B(n_303383008), .C(n_303183006), .D
		(n_291682891), .Z(n_303583010));
	notech_ao4 i_122741047(.A(n_55136), .B(n_27586), .C(n_311118888), .D(n_55075
		), .Z(n_303683011));
	notech_ao4 i_122641048(.A(n_55933), .B(n_55631), .C(n_55204), .D(n_27540
		), .Z(n_303783012));
	notech_ao4 i_122441050(.A(n_55192), .B(nbus_11326[20]), .C(n_55170), .D(n_56811
		), .Z(n_303983014));
	notech_and4 i_122941045(.A(n_303983014), .B(n_303783012), .C(n_303683011
		), .D(n_290782882), .Z(n_304183016));
	notech_ao4 i_122141053(.A(n_55526), .B(n_28608), .C(n_55091), .D(n_28631
		), .Z(n_304283017));
	notech_ao4 i_121941055(.A(n_2156), .B(n_28819), .C(n_55181), .D(n_29034)
		, .Z(n_304483019));
	notech_and4 i_122341051(.A(n_2187), .B(n_304483019), .C(n_304283017), .D
		(n_290482879), .Z(n_304683021));
	notech_ao4 i_121641058(.A(n_55181), .B(n_29017), .C(n_311218889), .D(n_55075
		), .Z(n_304783022));
	notech_ao4 i_121541059(.A(n_55204), .B(n_27539), .C(n_55136), .D(n_27585
		), .Z(n_304883023));
	notech_ao4 i_121341061(.A(n_55170), .B(n_56802), .C(n_55933), .D(n_55620
		), .Z(n_305083025));
	notech_and4 i_121841056(.A(n_305083025), .B(n_304883023), .C(n_304783022
		), .D(n_289582870), .Z(n_305283027));
	notech_ao4 i_121041064(.A(n_55091), .B(n_28630), .C(n_2318), .D(n_28848)
		, .Z(n_305383028));
	notech_ao4 i_120841066(.A(n_55161), .B(n_28818), .C(n_55366), .D(n_28792
		), .Z(n_305583030));
	notech_and4 i_121241062(.A(n_2187), .B(n_305583030), .C(n_305383028), .D
		(n_289282867), .Z(n_305783032));
	notech_ao4 i_120541069(.A(n_55136), .B(n_27584), .C(n_311318890), .D(n_55075
		), .Z(n_305883033));
	notech_ao4 i_120441070(.A(n_55933), .B(n_55609), .C(n_55204), .D(n_27538
		), .Z(n_305983034));
	notech_ao4 i_120241072(.A(n_55192), .B(nbus_11326[18]), .C(n_55170), .D(n_56793
		), .Z(n_306183036));
	notech_and4 i_120741067(.A(n_306183036), .B(n_305983034), .C(n_305883033
		), .D(n_288382858), .Z(n_306383038));
	notech_ao4 i_119941075(.A(n_55526), .B(n_28610), .C(n_55091), .D(n_28629
		), .Z(n_306483039));
	notech_ao4 i_119741077(.A(n_55161), .B(n_28817), .C(n_55181), .D(n_29014
		), .Z(n_306683041));
	notech_and4 i_120141073(.A(n_2187), .B(n_306683041), .C(n_306483039), .D
		(n_288082855), .Z(n_306883043));
	notech_or4 i_5635642(.A(fsm[3]), .B(fsm[0]), .C(n_60761), .D(n_57414), .Z
		(n_306983044));
	notech_ao4 i_83235759(.A(n_59795), .B(n_274788710), .C(n_58483), .D(n_307583050
		), .Z(n_307183046));
	notech_and2 i_102234722(.A(imm[7]), .B(n_307383048), .Z(n_307283047));
	notech_nand2 i_6235636(.A(n_56043), .B(n_56092), .Z(n_307383048));
	notech_nor2 i_32635758(.A(n_312283097), .B(n_327083245), .Z(n_307583050)
		);
	notech_or4 i_118734562(.A(calc_sz[3]), .B(calc_sz[0]), .C(n_260888755), 
		.D(n_54775), .Z(n_307683051));
	notech_or2 i_99234752(.A(n_54847), .B(n_59050), .Z(n_308583060));
	notech_nand3 i_100534739(.A(n_4699), .B(n_26556), .C(n_315788532), .Z(n_309883073
		));
	notech_or4 i_101934725(.A(n_260988754), .B(n_260888755), .C(n_54519), .D
		(n_28738), .Z(n_310783082));
	notech_ao4 i_101234732(.A(n_312283097), .B(n_327083245), .C(n_55484), .D
		(n_307283047), .Z(n_311083085));
	notech_nao3 i_101334731(.A(n_5837), .B(n_59795), .C(n_57382), .Z(n_311183086
		));
	notech_nao3 i_101434730(.A(n_5835), .B(n_26680), .C(n_55332), .Z(n_311283087
		));
	notech_or4 i_32781(.A(fsm[3]), .B(fsm[0]), .C(n_60761), .D(n_57382), .Z(n_311383088
		));
	notech_or4 i_32773(.A(n_58940), .B(n_60494), .C(n_59885), .D(n_2826), .Z
		(n_311483089));
	notech_nand2 i_32776(.A(n_26785), .B(n_312883103), .Z(n_311583090));
	notech_or4 i_32774(.A(n_2831), .B(n_2572), .C(n_274988708), .D(n_1041), 
		.Z(n_311683091));
	notech_or4 i_32767(.A(n_273188724), .B(n_60494), .C(n_57404), .D(n_59889
		), .Z(n_311783092));
	notech_nao3 i_32919(.A(n_57438), .B(n_26680), .C(n_1968), .Z(n_311883093
		));
	notech_or4 i_32914(.A(calc_sz[3]), .B(calc_sz[0]), .C(n_260888755), .D(n_54519
		), .Z(n_311983094));
	notech_or4 i_7935619(.A(n_59370), .B(n_2550), .C(n_59889), .D(n_2826), .Z
		(n_312083095));
	notech_or4 i_32916(.A(n_2582), .B(n_2599), .C(n_26296), .D(n_59795), .Z(n_312183096
		));
	notech_nand2 i_32769(.A(n_55195), .B(n_306983044), .Z(n_312283097));
	notech_ao4 i_222333546(.A(n_280372114), .B(n_55389), .C(n_57438), .D(n_54811
		), .Z(n_312683101));
	notech_nor2 i_221033559(.A(n_1968), .B(n_273288723), .Z(n_312883103));
	notech_ao4 i_199833770(.A(n_54427), .B(n_57326), .C(n_54405), .D(n_29641
		), .Z(n_313283107));
	notech_and4 i_200133767(.A(n_313283107), .B(n_311183086), .C(n_311283087
		), .D(n_26575), .Z(n_313383108));
	notech_ao4 i_199533773(.A(n_311883093), .B(n_28729), .C(n_54416), .D(nbus_11326
		[7]), .Z(n_313483109));
	notech_ao4 i_199433774(.A(n_307183046), .B(n_28618), .C(n_27526), .D(n_312183096
		), .Z(n_313683111));
	notech_ao4 i_199133777(.A(n_54735), .B(n_55578), .C(n_56631), .D(n_29482
		), .Z(n_313883113));
	notech_ao4 i_199033778(.A(n_55122), .B(nbus_11326[7]), .C(n_54863), .D(n_55400
		), .Z(n_313983114));
	notech_ao4 i_198833780(.A(n_54926), .B(nbus_11348[7]), .C(n_2246), .D(n_27545
		), .Z(n_314183116));
	notech_and4 i_199333775(.A(n_314183116), .B(n_313983114), .C(n_313883113
		), .D(n_309883073), .Z(n_314383118));
	notech_ao4 i_198533783(.A(n_54847), .B(n_59095), .C(n_54887), .D(n_28907
		), .Z(n_314483119));
	notech_ao4 i_198433784(.A(n_54836), .B(n_28058), .C(n_2311), .D(n_29333)
		, .Z(n_314583120));
	notech_ao4 i_198233786(.A(n_325083225), .B(n_29638), .C(n_324983224), .D
		(n_29634), .Z(n_314783122));
	notech_and4 i_198733781(.A(n_2312), .B(n_314783122), .C(n_314583120), .D
		(n_314483119), .Z(n_314983124));
	notech_ao4 i_197933789(.A(n_55122), .B(nbus_11326[6]), .C(n_56631), .D(n_29483
		), .Z(n_315083125));
	notech_ao4 i_197833790(.A(n_54908), .B(n_29633), .C(n_54926), .D(nbus_11348
		[6]), .Z(n_315183126));
	notech_ao4 i_197633792(.A(n_54863), .B(\nbus_11276[6] ), .C(n_54887), .D
		(n_28906), .Z(n_315383128));
	notech_and4 i_198133787(.A(n_308583060), .B(n_315383128), .C(n_315183126
		), .D(n_315083125), .Z(n_315583130));
	notech_ao4 i_197333795(.A(n_2246), .B(n_27542), .C(n_2311), .D(n_29331),
		 .Z(n_315683131));
	notech_ao4 i_197233796(.A(n_55111), .B(n_55566), .C(n_54836), .D(n_28057
		), .Z(n_315783132));
	notech_ao4 i_197033798(.A(n_325083225), .B(n_29632), .C(n_324983224), .D
		(n_29630), .Z(n_315983134));
	notech_and4 i_197533793(.A(n_2312), .B(n_315983134), .C(n_315783132), .D
		(n_315683131), .Z(n_316183136));
	notech_or2 i_21632923(.A(n_275688701), .B(n_59795), .Z(n_316283137));
	notech_nand3 i_22932920(.A(n_59299), .B(n_59290), .C(n_318583160), .Z(n_316383138
		));
	notech_nao3 i_47432908(.A(n_57451), .B(n_275688701), .C(n_312183096), .Z
		(n_316483139));
	notech_or2 i_7720(.A(n_54504), .B(opd[0]), .Z(n_316583140));
	notech_or2 i_134332850(.A(n_318383158), .B(n_26577), .Z(n_316683141));
	notech_nand3 i_9233174(.A(n_56126), .B(n_56092), .C(n_56049), .Z(n_316783142
		));
	notech_nand2 i_169132826(.A(n_275688701), .B(n_59889), .Z(n_316883143)
		);
	notech_and4 i_163533136(.A(n_326683241), .B(n_55992), .C(n_326183236), .D
		(n_326483239), .Z(n_316983144));
	notech_ao4 i_14932730(.A(n_328283257), .B(opd[4]), .C(n_331283287), .D(n_325783232
		), .Z(n_317083145));
	notech_and4 i_15032729(.A(n_328683261), .B(n_328883263), .C(n_331383288)
		, .D(n_328583260), .Z(n_317183146));
	notech_ao3 i_121433135(.A(n_56139), .B(n_327546813), .C(n_49223), .Z(n_317283147
		));
	notech_ao4 i_92833134(.A(n_58483), .B(n_318383158), .C(n_54486), .D(n_326983244
		), .Z(n_317383148));
	notech_ao4 i_122833122(.A(n_55958), .B(n_54530), .C(n_56104), .D(n_327583250
		), .Z(n_317683151));
	notech_and3 i_150133124(.A(n_54718), .B(n_55527), .C(n_325983234), .Z(n_317783152
		));
	notech_and3 i_150833125(.A(n_326083235), .B(n_55562), .C(n_55528), .Z(n_317883153
		));
	notech_nor2 i_36933133(.A(n_312283097), .B(n_318483159), .Z(n_318383158)
		);
	notech_and3 i_58732407(.A(n_57451), .B(n_275688701), .C(n_327083245), .Z
		(n_318483159));
	notech_nand2 i_59232403(.A(n_56081), .B(n_58656), .Z(n_318583160));
	notech_nao3 i_31732618(.A(opc_14[5]), .B(n_59889), .C(n_57451), .Z(n_319483169
		));
	notech_nao3 i_34032597(.A(n_5807), .B(n_59795), .C(n_57382), .Z(n_320783182
		));
	notech_nao3 i_33232603(.A(opd[0]), .B(n_55331), .C(n_54504), .Z(n_321083185
		));
	notech_or2 i_33332602(.A(n_316683141), .B(n_28590), .Z(n_321183186));
	notech_or4 i_36432573(.A(n_260988754), .B(n_260888755), .C(n_54519), .D(n_28736
		), .Z(n_321483189));
	notech_or2 i_36132576(.A(n_54427), .B(n_56685), .Z(n_321783192));
	notech_nao3 i_35832579(.A(n_5827), .B(n_59795), .C(n_57382), .Z(n_322083195
		));
	notech_nand2 i_37932559(.A(add_src[24]), .B(n_26579), .Z(n_323183206));
	notech_nor2 i_37632562(.A(n_55170), .B(n_56847), .Z(n_323483209));
	notech_ao3 i_37032568(.A(instrc[96]), .B(n_26760), .C(n_1967), .Z(n_323783212
		));
	notech_nand3 i_37132567(.A(nbus_137[24]), .B(n_1969), .C(n_59795), .Z(n_323883213
		));
	notech_or4 i_39632546(.A(n_55522), .B(n_1976), .C(n_353069302), .D(n_324883223
		), .Z(n_324583220));
	notech_nand3 i_39732545(.A(n_59780), .B(n_59889), .C(read_data[9]), .Z(n_324683221
		));
	notech_or4 i_39832544(.A(n_55958), .B(n_2255), .C(n_28060), .D(n_60504),
		 .Z(n_324783222));
	notech_and3 i_128633127(.A(n_55961), .B(n_55959), .C(n_55960), .Z(n_324883223
		));
	notech_nand2 i_33766(.A(rep_en1), .B(n_26596), .Z(n_324983224));
	notech_nand2 i_33765(.A(n_26889), .B(n_26596), .Z(n_325083225));
	notech_or2 i_33008(.A(n_327783252), .B(n_55299), .Z(n_325783232));
	notech_or4 i_25592(.A(n_272988726), .B(n_2647), .C(n_60563), .D(n_59380)
		, .Z(n_325883233));
	notech_or2 i_54832437(.A(n_56034), .B(eval_flag), .Z(n_325983234));
	notech_or4 i_55132434(.A(n_60761), .B(n_60719), .C(n_2216), .D(n_26599),
		 .Z(n_326083235));
	notech_nao3 i_23133101(.A(n_59299), .B(n_59268), .C(n_59290), .Z(n_326183236
		));
	notech_or4 i_59032404(.A(n_59259), .B(n_59268), .C(n_59281), .D(n_55328)
		, .Z(n_326483239));
	notech_ao4 i_129531805(.A(n_27518), .B(n_56023), .C(n_316383138), .D(n_29122
		), .Z(n_326683241));
	notech_nand2 i_128931807(.A(n_57451), .B(n_26296), .Z(n_326983244));
	notech_and3 i_18809(.A(n_274788710), .B(n_59885), .C(n_57445), .Z(n_327083245
		));
	notech_or4 i_126231833(.A(fsm[3]), .B(fsm[0]), .C(n_60761), .D(n_55334),
		 .Z(n_327583250));
	notech_nao3 i_159732986(.A(opd[0]), .B(opd[1]), .C(n_54504), .Z(n_327783252
		));
	notech_nao3 i_43232909(.A(n_275688701), .B(n_59885), .C(n_57451), .Z(n_327883253
		));
	notech_or4 i_142232984(.A(n_57451), .B(n_54486), .C(opd[0]), .D(opd[1]),
		 .Z(n_328083255));
	notech_nand2 i_120331877(.A(n_27564), .B(n_55299), .Z(n_328183256));
	notech_or4 i_176432983(.A(opd[0]), .B(n_327883253), .C(n_328183256), .D(opd
		[1]), .Z(n_328283257));
	notech_mux2 i_90032882(.S(opd[0]), .A(n_54504), .B(n_327883253), .Z(n_328383258
		));
	notech_mux2 i_120231878(.S(opd[1]), .A(n_54504), .B(n_327883253), .Z(n_328483259
		));
	notech_and2 i_116332982(.A(n_328383258), .B(n_328483259), .Z(n_328583260
		));
	notech_mux2 i_120131879(.S(opd[2]), .A(n_54504), .B(n_327883253), .Z(n_328683261
		));
	notech_and2 i_129632981(.A(n_328683261), .B(n_328583260), .Z(n_328783262
		));
	notech_mux2 i_120031880(.S(opd[3]), .A(n_54504), .B(n_327883253), .Z(n_328883263
		));
	notech_nand3 i_150932980(.A(n_328683261), .B(n_328583260), .C(n_328883263
		), .Z(n_328983264));
	notech_ao4 i_101232033(.A(n_55156), .B(n_57349), .C(n_55085), .D(n_55947
		), .Z(n_329483269));
	notech_and4 i_101832030(.A(n_329483269), .B(n_324683221), .C(n_324783222
		), .D(n_324583220), .Z(n_329583270));
	notech_ao4 i_100932035(.A(n_317783152), .B(n_55425), .C(n_317683151), .D
		(n_29048), .Z(n_329683271));
	notech_ao4 i_100832036(.A(n_29265), .B(n_54822), .C(n_317883153), .D(nbus_11273
		[9]), .Z(n_329783272));
	notech_ao4 i_93432103(.A(n_55192), .B(nbus_11326[24]), .C(n_55161), .D(n_28824
		), .Z(n_330283277));
	notech_nao3 i_93632101(.A(n_330283277), .B(n_323883213), .C(n_323783212)
		, .Z(n_330383278));
	notech_ao4 i_93232105(.A(n_55075), .B(n_57334), .C(n_55526), .D(n_28604)
		, .Z(n_330483279));
	notech_ao4 i_92932108(.A(n_55933), .B(n_56207), .C(n_55136), .D(n_27592)
		, .Z(n_330783282));
	notech_ao4 i_92632110(.A(n_55204), .B(n_27546), .C(n_55102), .D(n_28795)
		, .Z(n_330983284));
	notech_and4 i_93132106(.A(n_330983284), .B(n_330783282), .C(n_2187), .D(n_323183206
		), .Z(n_331183286));
	notech_nand2 i_92432111(.A(opd[4]), .B(opd[3]), .Z(n_331283287));
	notech_mux2 i_92332112(.S(opd[4]), .A(n_54504), .B(n_327883253), .Z(n_331383288
		));
	notech_mux2 i_91932115(.S(opd[5]), .A(n_317083145), .B(n_317183146), .Z(n_331483289
		));
	notech_ao4 i_91832116(.A(n_316483139), .B(n_27524), .C(n_316683141), .D(n_28581
		), .Z(n_331583290));
	notech_ao4 i_91632118(.A(n_317383148), .B(n_28616), .C(n_318383158), .D(n_317283147
		), .Z(n_331783292));
	notech_and4 i_92132113(.A(n_331783292), .B(n_331583290), .C(n_331483289)
		, .D(n_322083195), .Z(n_331983294));
	notech_ao4 i_91332121(.A(n_54405), .B(n_29648), .C(n_54472), .D(n_29647)
		, .Z(n_332083295));
	notech_ao4 i_91132123(.A(n_311883093), .B(n_28728), .C(n_54416), .D(nbus_11326
		[5]), .Z(n_332283297));
	notech_and4 i_91532119(.A(n_332283297), .B(n_332083295), .C(n_321483189)
		, .D(n_321783192), .Z(n_332483299));
	notech_ao4 i_90132133(.A(n_27520), .B(n_316483139), .C(n_328383258), .D(n_55331
		), .Z(n_332783302));
	notech_and3 i_90332131(.A(n_332783302), .B(n_321183186), .C(n_321083185)
		, .Z(n_332883303));
	notech_ao4 i_89832135(.A(n_317383148), .B(n_28612), .C(n_318383158), .D(n_316983144
		), .Z(n_332983304));
	notech_ao4 i_89532138(.A(n_54405), .B(n_29646), .C(n_54472), .D(n_29645)
		, .Z(n_333283307));
	notech_ao4 i_89432139(.A(n_54416), .B(nbus_11326[1]), .C(n_54427), .D(n_56649
		), .Z(n_333383308));
	notech_ao4 i_89232141(.A(n_311983094), .B(n_28732), .C(n_311883093), .D(n_28724
		), .Z(n_333583310));
	notech_and4 i_89732136(.A(n_328083255), .B(n_333583310), .C(n_333383308)
		, .D(n_333283307), .Z(n_333783312));
	notech_ao4 i_84832184(.A(n_54908), .B(n_29644), .C(n_2246), .D(n_27541),
		 .Z(n_333883313));
	notech_ao4 i_84732185(.A(n_29643), .B(n_324983224), .C(n_54926), .D(nbus_11348
		[5]), .Z(n_333983314));
	notech_ao4 i_84532187(.A(n_2311), .B(n_29329), .C(n_325083225), .D(n_29642
		), .Z(n_334183316));
	notech_and4 i_85032182(.A(n_334183316), .B(n_333983314), .C(n_333883313)
		, .D(n_319483169), .Z(n_334383318));
	notech_ao4 i_84232190(.A(n_54847), .B(n_59104), .C(\nbus_11276[5] ), .D(n_54863
		), .Z(n_334483319));
	notech_ao4 i_84132191(.A(n_55111), .B(n_55552), .C(n_55122), .D(nbus_11326
		[5]), .Z(n_334583320));
	notech_ao4 i_83932193(.A(n_56631), .B(n_29484), .C(n_54836), .D(n_28056)
		, .Z(n_334783322));
	notech_and4 i_84432188(.A(n_334783322), .B(n_334583320), .C(n_334483319)
		, .D(n_2312), .Z(n_334983324));
	notech_nand2 i_136070265(.A(n_316983144), .B(n_109081078), .Z(nbus_11313
		[1]));
	notech_or4 i_25037(.A(n_55248), .B(n_60583), .C(n_59885), .D(n_29123), .Z
		(n_335083325));
	notech_or4 i_103268291(.A(n_2793), .B(n_59771), .C(n_59163), .D(n_29123)
		, .Z(n_107542794));
	notech_nor2 i_19168(.A(n_54504), .B(n_28706), .Z(n_335283327));
	notech_nao3 i_47925(.A(n_54733), .B(n_206482046), .C(n_166381651), .Z(n_10174
		));
	notech_ao4 i_54741(.A(n_134060422), .B(n_59163), .C(n_59885), .D(n_201661090
		), .Z(\nbus_11353[10] ));
	notech_or4 i_54740(.A(n_165981647), .B(n_26511), .C(n_26494), .D(n_26509
		), .Z(\nbus_11353[9] ));
	notech_or4 i_53445(.A(n_60577), .B(n_165381641), .C(n_26510), .D(n_167281660
		), .Z(n_18922));
	notech_or4 i_48649(.A(n_166381651), .B(n_1919), .C(n_1915), .D(n_26511),
		 .Z(n_11472));
	notech_nao3 i_47881(.A(n_167781665), .B(n_168081668), .C(n_165281640), .Z
		(n_10124));
	notech_nand2 i_135965726(.A(n_168381671), .B(n_123381221), .Z(nbus_11313
		[0]));
	notech_nand2 i_136165725(.A(n_168781675), .B(n_123181219), .Z(nbus_11313
		[2]));
	notech_nand2 i_136265724(.A(n_168881676), .B(n_122981217), .Z(nbus_11313
		[3]));
	notech_nand2 i_136365723(.A(n_169081678), .B(n_122881216), .Z(nbus_11313
		[4]));
	notech_nand2 i_136465722(.A(n_317283147), .B(n_122781215), .Z(nbus_11313
		[5]));
	notech_nand2 i_136665721(.A(n_317283147), .B(n_122681214), .Z(nbus_11313
		[7]));
	notech_or4 i_155565720(.A(n_28975), .B(n_274588712), .C(n_2572), .D(n_62403
		), .Z(n_57417));
	notech_or4 i_158065719(.A(n_60540), .B(n_274588712), .C(n_2572), .D(n_60503
		), .Z(n_57415));
	notech_nand2 i_136565714(.A(n_317283147), .B(n_122581213), .Z(nbus_11313
		[6]));
	notech_or2 i_27865713(.A(n_55484), .B(n_122481212), .Z(nbus_11313[9]));
	notech_or2 i_28065712(.A(n_55484), .B(n_122381211), .Z(nbus_11313[10])
		);
	notech_or2 i_26065711(.A(n_55484), .B(n_122281210), .Z(nbus_11313[11])
		);
	notech_or2 i_26765710(.A(n_55478), .B(n_122181209), .Z(nbus_11313[12])
		);
	notech_or2 i_27265709(.A(n_55478), .B(n_122081208), .Z(nbus_11313[13])
		);
	notech_or2 i_27565708(.A(n_55478), .B(n_121981207), .Z(nbus_11313[14])
		);
	notech_or2 i_26165707(.A(n_55478), .B(n_121881206), .Z(nbus_11313[15])
		);
	notech_or2 i_148065705(.A(n_55478), .B(n_121781205), .Z(nbus_11313[17])
		);
	notech_or2 i_148165704(.A(n_55478), .B(n_121681204), .Z(nbus_11313[18])
		);
	notech_or2 i_26265703(.A(n_55478), .B(n_121581203), .Z(nbus_11313[19])
		);
	notech_or2 i_26965702(.A(n_55478), .B(n_121481202), .Z(nbus_11313[20])
		);
	notech_or2 i_27365701(.A(n_55478), .B(n_121381201), .Z(nbus_11313[21])
		);
	notech_or2 i_27665700(.A(n_55478), .B(n_121281200), .Z(nbus_11313[22])
		);
	notech_or2 i_26365699(.A(n_55478), .B(n_121181199), .Z(nbus_11313[23])
		);
	notech_or2 i_27065698(.A(n_55478), .B(n_121081198), .Z(nbus_11313[24])
		);
	notech_or2 i_27965697(.A(n_55478), .B(n_120981197), .Z(nbus_11313[25])
		);
	notech_or2 i_28165696(.A(n_55478), .B(n_120881196), .Z(nbus_11313[26])
		);
	notech_or2 i_26465695(.A(n_55478), .B(n_120781195), .Z(nbus_11313[27])
		);
	notech_or2 i_27165694(.A(n_55478), .B(n_120681194), .Z(nbus_11313[28])
		);
	notech_or2 i_27465693(.A(n_55478), .B(n_120581193), .Z(nbus_11313[29])
		);
	notech_or2 i_27765692(.A(n_55478), .B(n_120481192), .Z(nbus_11313[30])
		);
	notech_or2 i_26565691(.A(n_55478), .B(n_120381191), .Z(nbus_11313[31])
		);
	notech_ao4 i_207853285(.A(n_56130), .B(n_27653), .C(n_56092), .D(n_27694
		), .Z(n_171258000));
	notech_or4 i_6376(.A(n_164181629), .B(n_164281630), .C(n_26519), .D(n_26520
		), .Z(n_8721));
	notech_nand2 i_3327513(.A(n_172981717), .B(n_119381181), .Z(n_8472));
	notech_nand2 i_3227512(.A(n_173181719), .B(n_173081718), .Z(n_8467));
	notech_nand2 i_3127511(.A(n_173381721), .B(n_173281720), .Z(n_8462));
	notech_nand2 i_3027510(.A(n_173581723), .B(n_173481722), .Z(n_8457));
	notech_nand2 i_2927509(.A(n_173781725), .B(n_173681724), .Z(n_8452));
	notech_nand2 i_2827508(.A(n_173981727), .B(n_173881726), .Z(n_8447));
	notech_nand2 i_2727507(.A(n_174181729), .B(n_174081728), .Z(n_8442));
	notech_nand2 i_2627506(.A(n_174381731), .B(n_174281730), .Z(n_8437));
	notech_nand2 i_2527505(.A(n_174581733), .B(n_174481732), .Z(n_8432));
	notech_nand2 i_2427504(.A(n_174781735), .B(n_174681734), .Z(n_8427));
	notech_nand2 i_2327503(.A(n_174981737), .B(n_174881736), .Z(n_8422));
	notech_nand2 i_2227502(.A(n_175181739), .B(n_175081738), .Z(n_8417));
	notech_nand2 i_2127501(.A(n_175381741), .B(n_175281740), .Z(n_8412));
	notech_nand2 i_2027500(.A(n_175581743), .B(n_175481742), .Z(n_8407));
	notech_nand2 i_1927499(.A(n_175781745), .B(n_175681744), .Z(n_8402));
	notech_nand2 i_1827498(.A(n_175981747), .B(n_175881746), .Z(n_8397));
	notech_nand2 i_1727497(.A(n_176181749), .B(n_176081748), .Z(n_8392));
	notech_nand2 i_1627496(.A(n_176381751), .B(n_176281750), .Z(n_8387));
	notech_nand2 i_1527495(.A(n_176581753), .B(n_176481752), .Z(n_8382));
	notech_nand2 i_1427494(.A(n_176781755), .B(n_176681754), .Z(n_8377));
	notech_nand2 i_1327493(.A(n_176981757), .B(n_176881756), .Z(n_8372));
	notech_nand2 i_1227492(.A(n_177181759), .B(n_177081758), .Z(n_8367));
	notech_nand2 i_1127491(.A(n_177381761), .B(n_177281760), .Z(n_8362));
	notech_nand2 i_1027490(.A(n_177581763), .B(n_177481762), .Z(n_8357));
	notech_nand2 i_927489(.A(n_177781765), .B(n_177681764), .Z(n_8352));
	notech_nand2 i_827488(.A(n_177981767), .B(n_177881766), .Z(n_8347));
	notech_nand2 i_727487(.A(n_178181769), .B(n_178081768), .Z(n_8342));
	notech_nand2 i_627486(.A(n_178381771), .B(n_178281770), .Z(n_8337));
	notech_nand2 i_527485(.A(n_178581773), .B(n_178481772), .Z(n_8332));
	notech_nand2 i_427484(.A(n_178781775), .B(n_178681774), .Z(n_8327));
	notech_nand2 i_327483(.A(n_178981777), .B(n_178881776), .Z(n_8322));
	notech_nand2 i_227482(.A(n_179181779), .B(n_179081778), .Z(n_8317));
	notech_nand2 i_127481(.A(n_179281780), .B(n_119081178), .Z(n_8312));
	notech_and4 i_3216233(.A(n_179981787), .B(n_180181789), .C(n_179881786),
		 .D(n_150381491), .Z(n_21277));
	notech_nand3 i_3116232(.A(n_181081796), .B(n_180981795), .C(n_180881794)
		, .Z(n_21272));
	notech_nand3 i_3016231(.A(n_181981803), .B(n_181681802), .C(n_181581801)
		, .Z(n_21267));
	notech_nand3 i_2916230(.A(n_182881810), .B(n_182781809), .C(n_182681808)
		, .Z(n_21262));
	notech_nand3 i_2816229(.A(n_183581817), .B(n_183481816), .C(n_183381815)
		, .Z(n_21257));
	notech_nand3 i_2716228(.A(n_184281824), .B(n_184181823), .C(n_184081822)
		, .Z(n_21252));
	notech_nand3 i_2616227(.A(n_184981831), .B(n_184881830), .C(n_184781829)
		, .Z(n_21247));
	notech_nand3 i_2516226(.A(n_185681838), .B(n_185581837), .C(n_185481836)
		, .Z(n_21242));
	notech_nand3 i_2416225(.A(n_186381845), .B(n_186281844), .C(n_186181843)
		, .Z(n_21237));
	notech_nand3 i_2316224(.A(n_187081852), .B(n_186981851), .C(n_186881850)
		, .Z(n_21232));
	notech_nand3 i_2216223(.A(n_187781859), .B(n_187681858), .C(n_187581857)
		, .Z(n_21227));
	notech_nand3 i_2116222(.A(n_188481866), .B(n_188381865), .C(n_188281864)
		, .Z(n_21222));
	notech_nand3 i_2016221(.A(n_189181873), .B(n_189081872), .C(n_188981871)
		, .Z(n_21217));
	notech_nand3 i_1916220(.A(n_189881880), .B(n_189781879), .C(n_189681878)
		, .Z(n_21212));
	notech_nand3 i_1816219(.A(n_190581887), .B(n_190481886), .C(n_190381885)
		, .Z(n_21207));
	notech_and4 i_1616217(.A(n_191181893), .B(n_191381895), .C(n_136781355),
		 .D(n_191081892), .Z(n_21197));
	notech_and4 i_1516216(.A(n_191981901), .B(n_192181903), .C(n_135781345),
		 .D(n_191881900), .Z(n_21192));
	notech_and4 i_1416215(.A(n_192781909), .B(n_192981911), .C(n_134781335),
		 .D(n_192681908), .Z(n_21187));
	notech_and4 i_1316214(.A(n_193581917), .B(n_193781919), .C(n_133781325),
		 .D(n_193481916), .Z(n_21182));
	notech_and4 i_1216213(.A(n_194381925), .B(n_194581927), .C(n_132781315),
		 .D(n_194281924), .Z(n_21177));
	notech_and4 i_1116212(.A(n_195181933), .B(n_195381935), .C(n_131781305),
		 .D(n_195081932), .Z(n_21172));
	notech_and4 i_1016211(.A(n_195981941), .B(n_196181943), .C(n_130781295),
		 .D(n_195881940), .Z(n_21167));
	notech_and4 i_716208(.A(n_196781949), .B(n_196981951), .C(n_129781285), 
		.D(n_196681948), .Z(n_21152));
	notech_nand2 i_516206(.A(n_198181963), .B(n_197681958), .Z(n_21142));
	notech_nand2 i_416205(.A(n_199481976), .B(n_198881970), .Z(n_21137));
	notech_nand2 i_316204(.A(n_200681988), .B(n_200081982), .Z(n_21132));
	notech_nand2 i_116202(.A(n_201781999), .B(n_201281994), .Z(n_21122));
	notech_and2 i_208253281(.A(n_171057998), .B(n_170957997), .Z(n_171157999
		));
	notech_and2 i_103365675(.A(n_57415), .B(n_57417), .Z(n_207241703));
	notech_ao4 i_208053283(.A(n_55919), .B(n_27381), .C(n_55910), .D(n_27726
		), .Z(n_171057998));
	notech_ao4 i_208153282(.A(n_55893), .B(n_27758), .C(n_55934), .D(n_27797
		), .Z(n_170957997));
	notech_and4 i_209053273(.A(n_170657994), .B(n_170557993), .C(n_170357991
		), .D(n_170257990), .Z(n_170857996));
	notech_ao4 i_46273(.A(n_202682008), .B(n_29123), .C(n_271039498), .D(n_202482006
		), .Z(n_7487));
	notech_ao4 i_53106(.A(n_275788700), .B(n_107542794), .C(n_271039498), .D
		(n_202082002), .Z(\nbus_11345[0] ));
	notech_or2 i_26663579(.A(n_55478), .B(n_201882000), .Z(nbus_11313[8]));
	notech_and4 i_720658(.A(n_206682048), .B(n_206882050), .C(n_207282054), 
		.D(n_206382045), .Z(n_19821));
	notech_and4 i_520656(.A(n_207382055), .B(n_207582057), .C(n_207982061), 
		.D(n_205582037), .Z(n_19809));
	notech_and4 i_520976(.A(n_208082062), .B(n_208282064), .C(n_208782069), 
		.D(n_204782029), .Z(n_16723));
	notech_and4 i_916210(.A(n_209282074), .B(n_209482076), .C(n_203382015), 
		.D(n_209182073), .Z(n_21162));
	notech_or4 i_8763460(.A(n_60761), .B(n_60721), .C(n_60577), .D(n_29123),
		 .Z(n_271039498));
	notech_ao4 i_208453279(.A(n_55866), .B(n_27829), .C(n_56049), .D(n_27861
		), .Z(n_170657994));
	notech_or4 i_521552(.A(n_210982091), .B(n_212682108), .C(n_26547), .D(n_26546
		), .Z(n_16374));
	notech_and4 i_3017256(.A(n_212882110), .B(n_213082112), .C(n_213582117),
		 .D(n_210482086), .Z(n_15948));
	notech_or4 i_54738(.A(n_132860410), .B(n_132760409), .C(n_213682118), .D
		(n_26494), .Z(\nbus_11353[6] ));
	notech_and4 i_921300(.A(n_215182133), .B(n_215382135), .C(n_214182123), 
		.D(n_215082132), .Z(n_20649));
	notech_nand3 i_2520964(.A(n_220482185), .B(n_220382184), .C(n_220282183)
		, .Z(n_9123));
	notech_nand3 i_1621307(.A(n_221282192), .B(n_221182191), .C(n_221082190)
		, .Z(n_20691));
	notech_nand3 i_1321304(.A(n_222082199), .B(n_221982198), .C(n_221882197)
		, .Z(n_20673));
	notech_nand3 i_1121302(.A(n_222982207), .B(n_222882206), .C(n_222782205)
		, .Z(n_20661));
	notech_and4 i_1621851(.A(n_363088165), .B(n_223582213), .C(n_215582137),
		 .D(n_223482212), .Z(n_12491));
	notech_or4 i_2920968(.A(n_313168930), .B(n_269382668), .C(n_270482679), 
		.D(n_26566), .Z(n_9147));
	notech_or4 i_2820967(.A(n_264975488), .B(n_268582660), .C(n_271182686), 
		.D(n_26567), .Z(n_9141));
	notech_or4 i_2720966(.A(n_265975498), .B(n_267782652), .C(n_271882693), 
		.D(n_26568), .Z(n_9135));
	notech_or4 i_2620965(.A(n_173971058), .B(n_266982644), .C(n_272582700), 
		.D(n_26569), .Z(n_9129));
	notech_nand3 i_2420963(.A(n_273482709), .B(n_273382708), .C(n_273282707)
		, .Z(n_9117));
	notech_and4 i_2921320(.A(n_274082715), .B(n_273982714), .C(n_273782712),
		 .D(n_273682711), .Z(n_20769));
	notech_and4 i_2821319(.A(n_274682721), .B(n_274582720), .C(n_274382718),
		 .D(n_274282717), .Z(n_20763));
	notech_and4 i_2721318(.A(n_275282727), .B(n_275182726), .C(n_274982724),
		 .D(n_274882723), .Z(n_20757));
	notech_and4 i_2621317(.A(n_275882733), .B(n_275782732), .C(n_275582730),
		 .D(n_275482729), .Z(n_20751));
	notech_and4 i_2921864(.A(n_276082735), .B(n_276282737), .C(n_262882603),
		 .D(n_276682741), .Z(n_12569));
	notech_nand3 i_2821863(.A(n_276882743), .B(n_276782742), .C(n_277282747)
		, .Z(n_12563));
	notech_and4 i_2721862(.A(n_277382748), .B(n_277582750), .C(n_261482589),
		 .D(n_277982754), .Z(n_12557));
	notech_nand3 i_2621861(.A(n_278182756), .B(n_278082755), .C(n_278582760)
		, .Z(n_12551));
	notech_nand2 i_3016199(.A(n_279682771), .B(n_279182766), .Z(n_14266));
	notech_nand2 i_2916198(.A(n_280782782), .B(n_280282777), .Z(n_14260));
	notech_nand2 i_2816197(.A(n_281882793), .B(n_281382788), .Z(n_14254));
	notech_nand2 i_2716196(.A(n_282982804), .B(n_282482799), .Z(n_14248));
	notech_nand2 i_2616195(.A(n_284082815), .B(n_283582810), .Z(n_14242));
	notech_nand2 i_2416193(.A(n_285182826), .B(n_284682821), .Z(n_14230));
	notech_and4 i_2917255(.A(n_285282827), .B(n_285482829), .C(n_252882503),
		 .D(n_285982834), .Z(n_15942));
	notech_and4 i_2717253(.A(n_251982494), .B(n_286082835), .C(n_286282837),
		 .D(n_286782842), .Z(n_15930));
	notech_and4 i_2617252(.A(n_286882843), .B(n_287082845), .C(n_287582850),
		 .D(n_251082485), .Z(n_15924));
	notech_ao4 i_3045347(.A(n_56369), .B(n_27595), .C(n_55798), .D(n_308221969
		), .Z(n_304121928));
	notech_ao4 i_3245345(.A(n_27593), .B(n_56369), .C(n_55798), .D(n_308421971
		), .Z(n_303921926));
	notech_nand3 i_2220961(.A(n_298482959), .B(n_298382958), .C(n_298282957)
		, .Z(n_9105));
	notech_nand3 i_2020959(.A(n_299182966), .B(n_299082965), .C(n_298982964)
		, .Z(n_9093));
	notech_nand3 i_2121312(.A(n_299882973), .B(n_299782972), .C(n_299682971)
		, .Z(n_20721));
	notech_nand3 i_2021311(.A(n_300582980), .B(n_300482979), .C(n_300382978)
		, .Z(n_20715));
	notech_nand3 i_1921310(.A(n_301282987), .B(n_301182986), .C(n_301082985)
		, .Z(n_20709));
	notech_nand2 i_2316192(.A(n_302482999), .B(n_301982994), .Z(n_14224));
	notech_nand2 i_2216191(.A(n_303583010), .B(n_303083005), .Z(n_14218));
	notech_nand2 i_2116190(.A(n_304683021), .B(n_304183016), .Z(n_14212));
	notech_nand2 i_2016189(.A(n_305783032), .B(n_305283027), .Z(n_14206));
	notech_nand2 i_1916188(.A(n_306883043), .B(n_306383038), .Z(n_14200));
	notech_nand3 i_50598(.A(n_334588367), .B(n_334488368), .C(n_307683051), 
		.Z(\nbus_11314[16] ));
	notech_and4 i_52598(.A(n_282272133), .B(n_312683101), .C(n_187771188), .D
		(n_55645), .Z(\nbus_11339[16] ));
	notech_and2 i_8017(.A(n_56079), .B(n_26500), .Z(n_49223));
	notech_or4 i_173335714(.A(n_273188724), .B(n_2550), .C(n_274988708), .D(n_2399
		), .Z(n_57402));
	notech_or4 i_205935713(.A(n_2831), .B(n_274488713), .C(\opcode[0] ), .D(n_59380
		), .Z(n_57387));
	notech_and4 i_816209(.A(n_313483109), .B(n_313683111), .C(n_310783082), 
		.D(n_313383108), .Z(n_21157));
	notech_nand2 i_816817(.A(n_314983124), .B(n_314383118), .Z(n_9742));
	notech_nand2 i_716816(.A(n_316183136), .B(n_315583130), .Z(n_9737));
	notech_or4 i_1535672(.A(n_59259), .B(n_59268), .C(n_56196), .D(n_29008),
		 .Z(n_327546813));
	notech_ao4 i_208553278(.A(n_56023), .B(n_27898), .C(n_56013), .D(n_27930
		), .Z(n_170557993));
	notech_ao4 i_208753276(.A(n_55992), .B(n_27964), .C(n_55965), .D(n_27996
		), .Z(n_170357991));
	notech_ao4 i_208853275(.A(n_55947), .B(n_29094), .C(n_58483), .D(n_28030
		), .Z(n_170257990));
	notech_and4 i_209553268(.A(n_169957987), .B(n_169757985), .C(n_156457852
		), .D(n_156757855), .Z(n_170157989));
	notech_ao4 i_209153272(.A(n_55264), .B(n_57346), .C(n_354269312), .D(n_55542
		), .Z(n_169957987));
	notech_ao4 i_209353270(.A(n_353969310), .B(n_27577), .C(n_55492), .D(n_27531
		), .Z(n_169757985));
	notech_nand3 i_1021301(.A(n_329783272), .B(n_329683271), .C(n_329583270)
		, .Z(n_20655));
	notech_or4 i_2516194(.A(n_323483209), .B(n_330383278), .C(n_26584), .D(n_26585
		), .Z(n_14236));
	notech_nand2 i_616207(.A(n_332483299), .B(n_331983294), .Z(n_21147));
	notech_and4 i_216203(.A(n_332983304), .B(n_333783312), .C(n_320783182), 
		.D(n_332883303), .Z(n_21127));
	notech_nand2 i_616815(.A(n_334983324), .B(n_334383318), .Z(n_9732));
	notech_and4 i_210053263(.A(n_169457982), .B(n_169257980), .C(n_157057858
		), .D(n_157357861), .Z(n_169657984));
	notech_ao4 i_209653267(.A(n_59174), .B(n_26778), .C(n_26435), .D(n_29095
		), .Z(n_169457982));
	notech_ao4 i_209853265(.A(n_354469314), .B(n_169157979), .C(n_354369313)
		, .D(n_169057978), .Z(n_169257980));
	notech_nand2 i_955315(.A(n_62411), .B(opc[12]), .Z(n_169157979));
	notech_nand2 i_5455308(.A(opc_10[12]), .B(n_62403), .Z(n_169057978));
	notech_ao4 i_210153262(.A(n_56386), .B(n_29096), .C(n_56139), .D(n_27618
		), .Z(n_168757975));
	notech_ao4 i_210253261(.A(n_56130), .B(n_27654), .C(n_56092), .D(n_27695
		), .Z(n_168657974));
	notech_and2 i_210653257(.A(n_168457972), .B(n_168357971), .Z(n_168557973
		));
	notech_ao4 i_210453259(.A(n_55919), .B(n_27382), .C(n_55910), .D(n_27727
		), .Z(n_168457972));
	notech_ao4 i_210553258(.A(n_55893), .B(n_27760), .C(n_55934), .D(n_27798
		), .Z(n_168357971));
	notech_and4 i_211453249(.A(n_168057968), .B(n_167957967), .C(n_167757965
		), .D(n_167657964), .Z(n_168257970));
	notech_ao4 i_210853255(.A(n_55866), .B(n_27830), .C(n_56049), .D(n_27862
		), .Z(n_168057968));
	notech_ao4 i_210953254(.A(n_56033), .B(n_27899), .C(n_56013), .D(n_27931
		), .Z(n_167957967));
	notech_ao4 i_211153252(.A(n_55992), .B(n_27965), .C(n_55972), .D(n_27997
		), .Z(n_167757965));
	notech_ao4 i_211253251(.A(n_55947), .B(n_29097), .C(n_58487), .D(n_28031
		), .Z(n_167657964));
	notech_and4 i_211953244(.A(n_167357961), .B(n_167157959), .C(n_159257880
		), .D(n_159557883), .Z(n_167557963));
	notech_ao4 i_211553248(.A(n_55264), .B(n_57345), .C(n_354269312), .D(n_55552
		), .Z(n_167357961));
	notech_ao4 i_211753246(.A(n_27578), .B(n_353969310), .C(n_55492), .D(n_27532
		), .Z(n_167157959));
	notech_and4 i_212453239(.A(n_166857956), .B(n_166657954), .C(n_159857886
		), .D(n_160157889), .Z(n_167057958));
	notech_ao4 i_212053243(.A(n_59183), .B(n_26779), .C(n_26435), .D(n_29098
		), .Z(n_166857956));
	notech_ao4 i_212253241(.A(n_354469314), .B(n_166557953), .C(n_354369313)
		, .D(n_166457952), .Z(n_166657954));
	notech_nand2 i_755316(.A(n_62423), .B(opc[13]), .Z(n_166557953));
	notech_nand2 i_5355309(.A(opc_10[13]), .B(n_62403), .Z(n_166457952));
	notech_ao4 i_212553238(.A(n_56386), .B(n_29099), .C(n_56144), .D(n_27619
		), .Z(n_166157949));
	notech_ao4 i_212653237(.A(n_56130), .B(n_27655), .C(n_56092), .D(n_27696
		), .Z(n_166057948));
	notech_and2 i_213053233(.A(n_165857946), .B(n_165757945), .Z(n_165957947
		));
	notech_ao4 i_212853235(.A(n_55919), .B(n_27383), .C(n_55910), .D(n_27728
		), .Z(n_165857946));
	notech_ao4 i_212953234(.A(n_55893), .B(n_27761), .C(n_55934), .D(n_27799
		), .Z(n_165757945));
	notech_and4 i_213853225(.A(n_165457942), .B(n_165357941), .C(n_165157939
		), .D(n_165057938), .Z(n_165657944));
	notech_ao4 i_213253231(.A(n_55879), .B(n_27831), .C(n_56049), .D(n_27863
		), .Z(n_165457942));
	notech_ao4 i_213353230(.A(n_56033), .B(n_27900), .C(n_56013), .D(n_27932
		), .Z(n_165357941));
	notech_ao4 i_213553228(.A(n_55992), .B(n_27966), .C(n_55972), .D(n_27998
		), .Z(n_165157939));
	notech_ao4 i_213653227(.A(n_55947), .B(n_29100), .C(n_58487), .D(n_28032
		), .Z(n_165057938));
	notech_ao4 i_218053183(.A(n_56386), .B(n_29101), .C(n_56144), .D(n_27614
		), .Z(n_164757935));
	notech_ao4 i_218153182(.A(n_56130), .B(n_27649), .C(n_56092), .D(n_27691
		), .Z(n_164657934));
	notech_and2 i_218553178(.A(n_164457932), .B(n_164357931), .Z(n_164557933
		));
	notech_ao4 i_218353180(.A(n_55919), .B(n_27378), .C(n_55910), .D(n_27723
		), .Z(n_164457932));
	notech_ao4 i_218453179(.A(n_55893), .B(n_27755), .C(n_55934), .D(n_27794
		), .Z(n_164357931));
	notech_and4 i_219353170(.A(n_164057928), .B(n_163957927), .C(n_163757925
		), .D(n_163657924), .Z(n_164257930));
	notech_ao4 i_218753176(.A(n_27826), .B(n_55879), .C(n_56049), .D(n_27858
		), .Z(n_164057928));
	notech_ao4 i_218853175(.A(n_56033), .B(n_27895), .C(n_56013), .D(n_27927
		), .Z(n_163957927));
	notech_ao4 i_219053173(.A(n_55992), .B(n_27961), .C(n_55972), .D(n_27993
		), .Z(n_163757925));
	notech_ao4 i_219153172(.A(n_55947), .B(n_29102), .C(n_58487), .D(n_28027
		), .Z(n_163657924));
	notech_nand2 i_1855280(.A(opc_10[8]), .B(n_62403), .Z(n_161957907));
	notech_nand2 i_1755281(.A(n_62409), .B(opc[8]), .Z(n_161857906));
	notech_or4 i_109254250(.A(n_56172), .B(n_59250), .C(n_56345), .D(n_321831605
		), .Z(n_160157889));
	notech_nao3 i_109554247(.A(n_205688857), .B(n_6807), .C(n_205588858), .Z
		(n_159857886));
	notech_nand2 i_109854244(.A(opa[13]), .B(n_354069311), .Z(n_159557883)
		);
	notech_or2 i_110154241(.A(n_55263), .B(n_29037), .Z(n_159257880));
	notech_or4 i_106354278(.A(n_56177), .B(n_59250), .C(n_56345), .D(n_321931606
		), .Z(n_157357861));
	notech_nao3 i_106654275(.A(n_205688857), .B(n_6806), .C(n_58931), .Z(n_157057858
		));
	notech_nand2 i_106954272(.A(opa[12]), .B(n_354069311), .Z(n_156757855)
		);
	notech_or2 i_107254269(.A(n_55263), .B(n_29084), .Z(n_156457852));
	notech_or4 i_103354306(.A(n_56177), .B(n_59250), .C(n_56345), .D(n_322031607
		), .Z(n_154557833));
	notech_nao3 i_103654303(.A(n_205688857), .B(n_6805), .C(n_58931), .Z(n_154257830
		));
	notech_nand2 i_103954300(.A(n_354069311), .B(opa[11]), .Z(n_153957827)
		);
	notech_or2 i_104254297(.A(n_55263), .B(n_29080), .Z(n_153657824));
	notech_or4 i_100554334(.A(n_56104), .B(n_56354), .C(n_55934), .D(n_322131608
		), .Z(n_151757805));
	notech_nao3 i_100854331(.A(n_205688857), .B(n_6804), .C(n_58931), .Z(n_151457802
		));
	notech_nand2 i_101154328(.A(opa[10]), .B(n_354069311), .Z(n_151157799)
		);
	notech_or2 i_101454325(.A(n_55263), .B(n_29077), .Z(n_150857796));
	notech_nand2 i_99354346(.A(\add_len_pc[8] ), .B(n_55819), .Z(n_150557793
		));
	notech_nao3 i_99654343(.A(n_205688857), .B(n_6802), .C(n_58931), .Z(n_150257790
		));
	notech_nand2 i_99954340(.A(opa[8]), .B(n_354069311), .Z(n_149957787));
	notech_or2 i_100254337(.A(n_55263), .B(n_29045), .Z(n_149657784));
	notech_or4 i_15055155(.A(n_58660), .B(n_59281), .C(n_56345), .D(n_57293)
		, .Z(n_149357781));
	notech_or2 i_15355152(.A(n_55739), .B(n_27581), .Z(n_149057778));
	notech_or2 i_15655149(.A(n_356476400), .B(n_55430), .Z(n_148757775));
	notech_nao3 i_15955146(.A(\regs_1[15] ), .B(n_28140), .C(n_58496), .Z(n_148457772
		));
	notech_or2 i_14255163(.A(n_55318), .B(n_56748), .Z(n_147757765));
	notech_or2 i_14555160(.A(n_55431), .B(n_29037), .Z(n_147457762));
	notech_or2 i_13055175(.A(n_55318), .B(n_56739), .Z(n_146557753));
	notech_or2 i_13355172(.A(n_55431), .B(n_29084), .Z(n_146257750));
	notech_or4 i_11455191(.A(n_58660), .B(n_59281), .C(n_56345), .D(n_322031607
		), .Z(n_145757745));
	notech_or2 i_11755188(.A(n_55739), .B(n_27576), .Z(n_145457742));
	notech_or2 i_12055185(.A(n_55430), .B(n_57347), .Z(n_145157739));
	notech_nao3 i_12355182(.A(\regs_1[11] ), .B(n_28140), .C(n_58496), .Z(n_144857736
		));
	notech_and4 i_110956817(.A(n_141757705), .B(n_141557703), .C(n_122257510
		), .D(n_121957507), .Z(n_141957707));
	notech_ao4 i_110556821(.A(n_54771), .B(n_55590), .C(n_54742), .D(n_27582
		), .Z(n_141757705));
	notech_ao4 i_110756819(.A(n_54727), .B(n_58987), .C(n_29051), .D(n_54714
		), .Z(n_141557703));
	notech_and4 i_111456812(.A(n_141257700), .B(n_141057698), .C(n_122557513
		), .D(n_122857516), .Z(n_141457702));
	notech_ao4 i_111056816(.A(n_54685), .B(n_28478), .C(n_58523), .D(n_27280
		), .Z(n_141257700));
	notech_ao4 i_111256814(.A(n_54674), .B(n_27969), .C(n_54659), .D(n_28430
		), .Z(n_141057698));
	notech_and4 i_128756651(.A(n_120457492), .B(n_132957617), .C(n_54860), .D
		(n_122957517), .Z(n_140857696));
	notech_ao4 i_128956650(.A(n_318588504), .B(n_29053), .C(n_59150), .D(n_27520
		), .Z(n_140557693));
	notech_ao4 i_129056649(.A(n_57325), .B(n_55690), .C(n_353869309), .D(n_198858274
		), .Z(n_140457692));
	notech_and4 i_129856641(.A(n_140157689), .B(n_139957687), .C(n_139857686
		), .D(n_123657524), .Z(n_140357691));
	notech_ao4 i_129356646(.A(n_57357), .B(n_55257), .C(n_55265), .D(n_29049
		), .Z(n_140157689));
	notech_ao4 i_129556644(.A(n_194058226), .B(n_59753), .C(n_194358229), .D
		(n_55331), .Z(n_139957687));
	notech_ao4 i_129656643(.A(n_194258228), .B(n_56649), .C(n_59183), .D(n_26633
		), .Z(n_139857686));
	notech_and4 i_130056639(.A(n_132857616), .B(n_54860), .C(n_120557493), .D
		(n_124157529), .Z(n_139657684));
	notech_ao4 i_130156638(.A(n_29056), .B(n_318588504), .C(n_353569307), .D
		(n_198858274), .Z(n_139357681));
	notech_ao4 i_130356637(.A(n_353469306), .B(n_198758273), .C(n_59150), .D
		(n_27521), .Z(n_139257680));
	notech_and4 i_131156629(.A(n_124857536), .B(n_138957677), .C(n_138757675
		), .D(n_138657674), .Z(n_139157679));
	notech_ao4 i_130656634(.A(n_194358229), .B(n_55299), .C(n_194258228), .D
		(nbus_11273[2]), .Z(n_138957677));
	notech_ao4 i_130856632(.A(n_322488466), .B(n_55257), .C(n_55265), .D(n_29050
		), .Z(n_138757675));
	notech_ao4 i_130956631(.A(n_194058226), .B(n_55289), .C(n_59183), .D(n_26634
		), .Z(n_138657674));
	notech_and3 i_131856627(.A(n_169564033), .B(n_174464082), .C(n_138357671
		), .Z(n_138457672));
	notech_ao4 i_131456628(.A(n_318488505), .B(n_29059), .C(n_318588504), .D
		(n_29058), .Z(n_138357671));
	notech_ao4 i_131956626(.A(n_316288527), .B(n_198758273), .C(n_59150), .D
		(n_27523), .Z(n_138157669));
	notech_and4 i_132756618(.A(n_126057548), .B(n_137857666), .C(n_137657664
		), .D(n_137557663), .Z(n_138057668));
	notech_ao4 i_132256623(.A(n_194358229), .B(n_58548), .C(n_194258228), .D
		(n_56676), .Z(n_137857666));
	notech_ao4 i_132456621(.A(n_321188478), .B(n_55257), .C(n_55265), .D(n_29063
		), .Z(n_137657664));
	notech_ao4 i_132556620(.A(n_194058226), .B(n_55365), .C(n_59183), .D(n_26636
		), .Z(n_137557663));
	notech_and4 i_132956616(.A(n_132757615), .B(n_132657614), .C(n_54860), .D
		(n_126557553), .Z(n_137357661));
	notech_ao4 i_133056615(.A(n_318588504), .B(n_29064), .C(n_351265801), .D
		(n_198758273), .Z(n_137057658));
	notech_ao4 i_133156614(.A(n_57321), .B(n_55690), .C(n_27566), .D(n_194358229
		), .Z(n_136957657));
	notech_and4 i_134056606(.A(n_136657654), .B(n_136457652), .C(n_136357651
		), .D(n_127257560), .Z(n_136857656));
	notech_ao4 i_133456611(.A(n_29065), .B(n_55265), .C(n_322788463), .D(n_55257
		), .Z(n_136657654));
	notech_ao4 i_133656609(.A(n_59150), .B(n_27524), .C(n_351365802), .D(n_198858274
		), .Z(n_136457652));
	notech_ao4 i_133756608(.A(n_194058226), .B(n_55375), .C(n_59183), .D(n_26637
		), .Z(n_136357651));
	notech_and4 i_134256604(.A(n_144577845), .B(n_183678231), .C(n_54860), .D
		(n_127757565), .Z(n_136157649));
	notech_ao4 i_134356603(.A(n_318588504), .B(n_29066), .C(n_59150), .D(n_27525
		), .Z(n_135857646));
	notech_ao4 i_134456602(.A(n_57320), .B(n_55690), .C(n_316588524), .D(n_198758273
		), .Z(n_135757645));
	notech_and4 i_135256594(.A(n_135457642), .B(n_135257640), .C(n_135157639
		), .D(n_128457572), .Z(n_135657644));
	notech_ao4 i_134756599(.A(n_194358229), .B(n_27568), .C(n_194258228), .D
		(n_56694), .Z(n_135457642));
	notech_ao4 i_134956597(.A(n_57352), .B(n_55257), .C(n_55265), .D(n_29068
		), .Z(n_135257640));
	notech_ao4 i_135056596(.A(n_194058226), .B(n_55387), .C(n_59183), .D(n_26638
		), .Z(n_135157639));
	notech_and3 i_135456592(.A(n_150874376), .B(n_158074448), .C(n_134857636
		), .Z(n_134957637));
	notech_ao4 i_135356593(.A(n_2675), .B(n_55690), .C(n_318488505), .D(n_29076
		), .Z(n_134857636));
	notech_ao4 i_135556591(.A(n_2680), .B(n_198858274), .C(n_2679), .D(n_198758273
		), .Z(n_134657634));
	notech_and4 i_136356583(.A(n_134357631), .B(n_134157629), .C(n_134057628
		), .D(n_129657584), .Z(n_134557633));
	notech_ao4 i_135856588(.A(n_194258228), .B(n_57326), .C(n_57351), .D(n_55257
		), .Z(n_134357631));
	notech_ao4 i_136056586(.A(n_59150), .B(n_27526), .C(n_55265), .D(n_28983
		), .Z(n_134157629));
	notech_ao4 i_136156585(.A(n_194058226), .B(n_55400), .C(n_59181), .D(n_26640
		), .Z(n_134057628));
	notech_and4 i_146756482(.A(n_133757625), .B(n_133557623), .C(n_130357591
		), .D(n_130657594), .Z(n_133957627));
	notech_ao4 i_146356486(.A(n_54822), .B(n_27146), .C(n_55740), .D(n_27568
		), .Z(n_133757625));
	notech_ao4 i_146556484(.A(n_55518), .B(n_57352), .C(n_55380), .D(n_55387
		), .Z(n_133557623));
	notech_and4 i_147456477(.A(n_130957597), .B(n_133257620), .C(n_131257600
		), .D(n_133057618), .Z(n_133457622));
	notech_ao4 i_146856481(.A(n_249734123), .B(n_29068), .C(n_249534121), .D
		(n_316588524), .Z(n_133257620));
	notech_ao4 i_147056479(.A(n_252034146), .B(n_120157489), .C(n_56694), .D
		(n_249634122), .Z(n_133057618));
	notech_ao4 i_167756280(.A(n_316688523), .B(n_56649), .C(n_249334119), .D
		(n_60463), .Z(n_132957617));
	notech_ao4 i_167856279(.A(n_322488466), .B(n_316788522), .C(n_249234118)
		, .D(n_60463), .Z(n_132857616));
	notech_ao4 i_168056277(.A(n_316688523), .B(n_56685), .C(n_262436779), .D
		(n_29065), .Z(n_132757615));
	notech_ao4 i_168156276(.A(n_322788463), .B(n_316788522), .C(n_132557613)
		, .D(n_55854), .Z(n_132657614));
	notech_or4 i_168256275(.A(n_60761), .B(n_60721), .C(n_60577), .D(n_55375
		), .Z(n_132557613));
	notech_ao4 i_172556233(.A(n_54505), .B(n_250234128), .C(n_2327), .D(n_55854
		), .Z(n_132357611));
	notech_or4 i_91557002(.A(n_57378), .B(eval_flag), .C(n_59885), .D(n_121457502
		), .Z(n_132157609));
	notech_or4 i_67357226(.A(n_56449), .B(n_120857496), .C(n_316488525), .D(n_55522
		), .Z(n_131257600));
	notech_or4 i_67657223(.A(n_260988754), .B(n_260888755), .C(n_252034146),
		 .D(n_57433), .Z(n_130957597));
	notech_or4 i_67957220(.A(n_56196), .B(n_59250), .C(n_55827), .D(n_57320)
		, .Z(n_130657594));
	notech_nand3 i_68257217(.A(n_59780), .B(n_59885), .C(read_data[6]), .Z(n_130357591
		));
	notech_or2 i_53757343(.A(n_194358229), .B(n_27570), .Z(n_129657584));
	notech_nao3 i_54157340(.A(n_4682), .B(n_60138), .C(n_58496), .Z(n_129357581
		));
	notech_nao3 i_52557355(.A(n_62423), .B(opc[6]), .C(n_198858274), .Z(n_128457572
		));
	notech_nao3 i_53057350(.A(\regs_1[6] ), .B(n_28140), .C(n_58496), .Z(n_127757565
		));
	notech_or2 i_51257367(.A(n_194258228), .B(n_56685), .Z(n_127257560));
	notech_nao3 i_51757362(.A(\regs_1[5] ), .B(n_28140), .C(n_58496), .Z(n_126557553
		));
	notech_or4 i_50057379(.A(n_56569), .B(n_56354), .C(n_55924), .D(n_319588494
		), .Z(n_126057548));
	notech_nao3 i_50357376(.A(n_62409), .B(opc[4]), .C(n_198858274), .Z(n_125757545
		));
	notech_or4 i_48657391(.A(n_56569), .B(n_56354), .C(n_55924), .D(n_57324)
		, .Z(n_124857536));
	notech_nao3 i_49257386(.A(\regs_1[2] ), .B(n_28140), .C(n_58496), .Z(n_124157529
		));
	notech_nao3 i_47457403(.A(opc_10[1]), .B(n_62419), .C(n_198758273), .Z(n_123657524
		));
	notech_nao3 i_47957398(.A(\regs_1[1] ), .B(n_28140), .C(n_58496), .Z(n_122957517
		));
	notech_nand3 i_25457607(.A(n_6382), .B(n_58591), .C(n_59795), .Z(n_122857516
		));
	notech_nao3 i_25757604(.A(n_6381), .B(n_59809), .C(n_58886), .Z(n_122557513
		));
	notech_nand2 i_26057601(.A(Daddrs_1[16]), .B(n_54701), .Z(n_122257510)
		);
	notech_nao3 i_26357598(.A(Daddrs_8[16]), .B(n_55040), .C(n_55149), .Z(n_121957507
		));
	notech_ao3 i_2257835(.A(n_56112), .B(n_56104), .C(n_56569), .Z(n_121457502
		));
	notech_or4 i_89257023(.A(n_60767), .B(n_60721), .C(n_58931), .D(n_273188724
		), .Z(n_121357501));
	notech_and3 i_84857067(.A(n_55958), .B(n_55960), .C(n_55959), .Z(n_120857496
		));
	notech_or2 i_83857077(.A(n_316688523), .B(n_56658), .Z(n_120557493));
	notech_or2 i_83457080(.A(n_57357), .B(n_316788522), .Z(n_120457492));
	notech_or2 i_70657201(.A(n_56569), .B(n_55302), .Z(n_120357491));
	notech_or4 i_68457215(.A(n_327446814), .B(n_1845), .C(n_56560), .D(opa[7
		]), .Z(n_120257490));
	notech_and2 i_4357814(.A(n_120257490), .B(n_55115), .Z(n_120157489));
	notech_and4 i_97359655(.A(n_191467734), .B(n_54860), .C(n_191367733), .D
		(n_111857406), .Z(n_119657484));
	notech_ao4 i_97459654(.A(n_318588504), .B(n_29041), .C(n_353269304), .D(n_198758273
		), .Z(n_119357481));
	notech_ao4 i_97559653(.A(n_57323), .B(n_55690), .C(n_194358229), .D(n_27564
		), .Z(n_119257480));
	notech_and4 i_98459645(.A(n_118957477), .B(n_118757475), .C(n_118657474)
		, .D(n_112557413), .Z(n_119157479));
	notech_ao4 i_97859650(.A(n_55265), .B(n_29043), .C(n_322688464), .D(n_55257
		), .Z(n_118957477));
	notech_ao4 i_98159648(.A(n_59150), .B(n_27522), .C(n_353369305), .D(n_198858274
		), .Z(n_118757475));
	notech_ao4 i_98259647(.A(n_194058226), .B(n_55277), .C(n_59181), .D(n_26635
		), .Z(n_118657474));
	notech_and4 i_98959640(.A(n_118357471), .B(n_113557423), .C(n_118157469)
		, .D(n_113257420), .Z(n_118557473));
	notech_ao4 i_98559644(.A(n_318588504), .B(n_29044), .C(n_59150), .D(n_27527
		), .Z(n_118357471));
	notech_ao4 i_98759642(.A(n_59181), .B(n_26641), .C(n_55739), .D(n_27571)
		, .Z(n_118157469));
	notech_and4 i_99459635(.A(n_117857466), .B(n_117657464), .C(n_113857426)
		, .D(n_114157429), .Z(n_118057468));
	notech_ao4 i_99059639(.A(n_55430), .B(n_57350), .C(n_55318), .D(n_56703)
		, .Z(n_117857466));
	notech_ao4 i_99259637(.A(n_161957907), .B(n_261036765), .C(n_161857906),
		 .D(n_260936764), .Z(n_117657464));
	notech_and3 i_99659633(.A(n_116357451), .B(n_116257450), .C(n_117357461)
		, .Z(n_117457462));
	notech_ao4 i_99559634(.A(n_318488505), .B(n_29047), .C(n_318588504), .D(n_29046
		), .Z(n_117357461));
	notech_ao4 i_99759632(.A(n_29048), .B(n_317988510), .C(n_57349), .D(n_318088509
		), .Z(n_117157459));
	notech_and4 i_100559624(.A(n_114957437), .B(n_116857456), .C(n_116657454
		), .D(n_116557453), .Z(n_117057458));
	notech_ao4 i_100059629(.A(n_59183), .B(n_26643), .C(n_55739), .D(n_27574
		), .Z(n_116857456));
	notech_ao4 i_100259627(.A(n_55501), .B(n_56712), .C(n_55500), .D(n_55425
		), .Z(n_116657454));
	notech_ao4 i_100359626(.A(n_352969301), .B(n_261036765), .C(n_353069302)
		, .D(n_260936764), .Z(n_116557453));
	notech_ao4 i_133759315(.A(n_55425), .B(n_55791), .C(n_56712), .D(n_55790
		), .Z(n_116357451));
	notech_ao4 i_133859314(.A(n_55789), .B(n_29048), .C(n_57349), .D(n_55786
		), .Z(n_116257450));
	notech_or4 i_85659758(.A(n_26190), .B(n_55524), .C(n_60577), .D(n_59885)
		, .Z(n_115857446));
	notech_or4 i_21360342(.A(n_58660), .B(n_59281), .C(n_56345), .D(n_57299)
		, .Z(n_114957437));
	notech_or4 i_21660339(.A(n_60577), .B(n_59817), .C(n_59771), .D(n_27528)
		, .Z(n_114657434));
	notech_or2 i_19760358(.A(n_55317), .B(n_55413), .Z(n_114157429));
	notech_or2 i_20060355(.A(n_55431), .B(n_29045), .Z(n_113857426));
	notech_or4 i_20360352(.A(n_58660), .B(n_59281), .C(n_56345), .D(n_57300)
		, .Z(n_113557423));
	notech_nao3 i_20660349(.A(\regs_1[8] ), .B(n_28140), .C(n_58496), .Z(n_113257420
		));
	notech_or2 i_18960366(.A(n_194258228), .B(n_56667), .Z(n_112557413));
	notech_nao3 i_19460361(.A(\regs_1[3] ), .B(n_28140), .C(n_58496), .Z(n_111857406
		));
	notech_and2 i_83859772(.A(n_56040), .B(n_261436769), .Z(n_111757405));
	notech_ao4 i_120267092(.A(n_27341992), .B(n_27347), .C(n_57345), .D(n_26595
		), .Z(n_111657404));
	notech_ao4 i_120167093(.A(n_28442003), .B(n_27314), .C(n_56415), .D(n_26949
		), .Z(n_111557403));
	notech_ao4 i_119567099(.A(n_27341992), .B(n_27346), .C(n_57346), .D(n_26595
		), .Z(n_111457402));
	notech_ao4 i_119467100(.A(n_28442003), .B(n_27313), .C(n_56415), .D(n_26947
		), .Z(n_111357401));
	notech_ao4 i_118867106(.A(n_27341992), .B(n_27345), .C(n_57347), .D(n_26595
		), .Z(n_111257400));
	notech_ao4 i_118767107(.A(n_28442003), .B(n_27312), .C(n_56409), .D(n_26945
		), .Z(n_111157399));
	notech_ao4 i_118167113(.A(n_27341992), .B(n_27343), .C(n_26595), .D(n_57348
		), .Z(n_111057398));
	notech_ao4 i_118067114(.A(n_28442003), .B(n_27311), .C(n_56409), .D(n_26943
		), .Z(n_110957397));
	notech_ao4 i_116767127(.A(n_27341992), .B(n_27341), .C(n_57350), .D(n_26595
		), .Z(n_110857396));
	notech_ao4 i_116667128(.A(n_28442003), .B(n_27309), .C(n_56404), .D(n_26939
		), .Z(n_110757395));
	notech_ao4 i_115367141(.A(n_27341992), .B(n_27339), .C(n_26595), .D(n_57352
		), .Z(n_110657394));
	notech_ao4 i_115267142(.A(n_28442003), .B(n_27307), .C(n_56404), .D(n_26935
		), .Z(n_110557393));
	notech_nand2 i_1417816(.A(n_111657404), .B(n_111557403), .Z(write_data_26
		[13]));
	notech_nand2 i_1317815(.A(n_111457402), .B(n_111357401), .Z(write_data_26
		[12]));
	notech_nand2 i_1217814(.A(n_111257400), .B(n_111157399), .Z(write_data_26
		[11]));
	notech_nand2 i_1117813(.A(n_111057398), .B(n_110957397), .Z(write_data_26
		[10]));
	notech_nand2 i_917811(.A(n_110857396), .B(n_110757395), .Z(write_data_26
		[8]));
	notech_nand2 i_717809(.A(n_110657394), .B(n_110557393), .Z(write_data_26
		[6]));
	notech_or4 i_116(.A(n_272788728), .B(n_260788756), .C(n_60767), .D(n_60721
		), .Z(n_2838));
	notech_or4 i_107(.A(n_2385), .B(n_2361), .C(n_273188724), .D(n_2550), .Z
		(n_2837));
	notech_nand3 i_23448(.A(n_276288695), .B(n_26625), .C(n_274788710), .Z(n_2835
		));
	notech_or4 i_17357(.A(n_275288705), .B(n_2550), .C(n_274488713), .D(n_59885
		), .Z(n_2834));
	notech_or4 i_17356(.A(n_273188724), .B(n_2550), .C(n_274488713), .D(n_59885
		), .Z(n_2833));
	notech_nand2 i_1908(.A(vliw_pc[3]), .B(n_27268), .Z(n_2832));
	notech_or2 i_1194(.A(n_26663), .B(n_2340), .Z(n_2831));
	notech_or4 i_1169(.A(n_60563), .B(n_62437), .C(n_60503), .D(\opcode[3] )
		, .Z(n_2830));
	notech_nand2 i_899(.A(n_57445), .B(n_275788700), .Z(n_4737261));
	notech_or2 i_505(.A(n_275388704), .B(n_2835), .Z(n_2828));
	notech_nao3 i_258(.A(n_62411), .B(n_26867), .C(n_60540), .Z(n_2826));
	notech_or4 i_220(.A(n_2341), .B(n_2385), .C(n_2562), .D(n_272788728), .Z
		(n_2825));
	notech_nao3 i_46372(.A(fsm[2]), .B(n_244556263), .C(n_2584), .Z(n_2824)
		);
	notech_or4 i_46375(.A(n_2584), .B(n_27265), .C(fsm[0]), .D(fsm[2]), .Z(n_2823
		));
	notech_or4 i_46377(.A(fsm[0]), .B(n_2582), .C(n_27264), .D(n_27265), .Z(n_2822
		));
	notech_and2 i_580(.A(n_2822), .B(n_2823), .Z(n_2821));
	notech_or4 i_46374(.A(n_2582), .B(n_27265), .C(n_27262), .D(fsm[2]), .Z(n_55641
		));
	notech_or4 i_34646(.A(n_2831), .B(n_2572), .C(n_54689), .D(n_59885), .Z(n_2820
		));
	notech_nand3 i_34643(.A(n_57438), .B(n_26295), .C(n_59817), .Z(n_2819)
		);
	notech_or4 i_34641(.A(n_274488713), .B(n_274588712), .C(n_57438), .D(n_59885
		), .Z(n_2818));
	notech_nao3 i_34640(.A(n_57438), .B(n_59817), .C(n_57409), .Z(n_2817));
	notech_or4 i_34635(.A(calc_sz[3]), .B(calc_sz[0]), .C(n_260888755), .D(n_2805
		), .Z(n_2816));
	notech_or4 i_34634(.A(calc_sz[3]), .B(calc_sz[0]), .C(n_260888755), .D(n_2834
		), .Z(n_2815));
	notech_or4 i_34631(.A(n_272788728), .B(n_260788756), .C(n_57438), .D(n_59890
		), .Z(n_2814));
	notech_or4 i_34629(.A(calc_sz[3]), .B(calc_sz[2]), .C(n_260688757), .D(n_2838
		), .Z(n_2813));
	notech_or4 i_34622(.A(n_60767), .B(n_60721), .C(n_59364), .D(n_2610), .Z
		(n_2812));
	notech_nao3 i_34620(.A(n_57438), .B(n_59817), .C(n_57412), .Z(n_2811));
	notech_nao3 i_34290(.A(n_2575), .B(n_244056258), .C(n_2797), .Z(n_2810)
		);
	notech_or2 i_34287(.A(n_275988698), .B(n_2596), .Z(n_2809));
	notech_nand3 i_34286(.A(n_2797), .B(n_2575), .C(n_244056258), .Z(n_2808)
		);
	notech_or4 i_34281(.A(n_57383), .B(n_57367), .C(n_106813462), .D(n_59890
		), .Z(n_2807));
	notech_or4 i_34279(.A(n_2801), .B(n_60525), .C(n_2739), .D(n_59890), .Z(n_2806
		));
	notech_or4 i_34274(.A(n_58940), .B(n_2550), .C(n_274488713), .D(n_59890)
		, .Z(n_2805));
	notech_or4 i_34270(.A(fsm[3]), .B(fsm[0]), .C(n_60767), .D(n_2227), .Z(n_2804
		));
	notech_or4 i_34262(.A(n_2740), .B(n_2801), .C(n_60525), .D(n_59890), .Z(n_2803
		));
	notech_or4 i_34255(.A(n_2796), .B(n_2801), .C(n_59890), .D(n_26315), .Z(n_2802
		));
	notech_or4 i_34252(.A(n_2550), .B(n_60563), .C(n_62437), .D(n_106813462)
		, .Z(n_2801));
	notech_or4 i_34249(.A(n_60767), .B(n_60721), .C(n_58940), .D(n_2610), .Z
		(n_280088689));
	notech_or4 i_34247(.A(fsm[3]), .B(fsm[0]), .C(n_60761), .D(n_2798), .Z(n_2799
		));
	notech_or4 i_34246(.A(n_275288705), .B(n_2550), .C(n_274988708), .D(n_2399
		), .Z(n_2798));
	notech_or4 i_1142(.A(n_60767), .B(n_60721), .C(n_272588730), .D(n_58940)
		, .Z(n_55230));
	notech_or4 i_970(.A(fsm[3]), .B(fsm[0]), .C(n_60767), .D(n_57390), .Z(n_55393
		));
	notech_or4 i_413(.A(n_60761), .B(n_60719), .C(n_273288723), .D(n_2386), 
		.Z(n_55936));
	notech_or4 i_1141(.A(n_60761), .B(n_60719), .C(n_273188724), .D(n_2610),
		 .Z(n_55231));
	notech_nand2 i_210044(.A(sign_div), .B(opd[31]), .Z(n_2797));
	notech_nand2 i_1225(.A(n_57367), .B(n_60479), .Z(n_2796));
	notech_or4 i_29814(.A(fsm[3]), .B(fsm[0]), .C(n_60762), .D(n_57413), .Z(n_2795
		));
	notech_nand2 i_210004(.A(rep_en2), .B(n_2770), .Z(n_57430));
	notech_nao3 i_1647(.A(n_26867), .B(n_2573), .C(n_2550), .Z(n_57413));
	notech_or2 i_2054(.A(n_2388), .B(n_2831), .Z(n_57388));
	notech_nao3 i_1751(.A(n_60540), .B(n_62419), .C(n_260788756), .Z(n_57399
		));
	notech_or4 i_1654(.A(n_2550), .B(n_274488713), .C(n_62395), .D(n_62437),
		 .Z(n_57412));
	notech_or4 i_1671(.A(n_60540), .B(n_275488703), .C(n_62419), .D(n_2586),
		 .Z(n_57409));
	notech_or4 i_1666(.A(n_60540), .B(n_274588712), .C(n_62419), .D(n_2586),
		 .Z(n_57410));
	notech_nand2 i_810(.A(nbus_11326[3]), .B(nbus_11326[2]), .Z(n_55541));
	notech_nand2 i_29518(.A(n_2771), .B(n_59817), .Z(n_2794));
	notech_or4 i_25513(.A(n_275088707), .B(n_2835), .C(n_2792), .D(n_26612),
		 .Z(n_2793));
	notech_nand2 i_25505(.A(n_57451), .B(n_2593), .Z(n_2792));
	notech_or4 i_46368(.A(n_2582), .B(n_27262), .C(fsm[3]), .D(fsm[2]), .Z(n_57444
		));
	notech_or4 i_46378(.A(n_2582), .B(n_27265), .C(n_27264), .D(n_27262), .Z
		(n_57434));
	notech_nao3 i_46370(.A(n_244556263), .B(fsm[2]), .C(n_2582), .Z(n_57442)
		);
	notech_or4 i_46367(.A(fsm[1]), .B(n_60719), .C(n_27266), .D(fsm[2]), .Z(n_57445
		));
	notech_or4 i_46371(.A(fsm[3]), .B(fsm[0]), .C(n_2584), .D(n_27264), .Z(n_57441
		));
	notech_nao3 i_127961(.A(n_2512), .B(n_227588798), .C(n_228888785), .Z(\opcode[0] 
		));
	notech_nand3 i_1871(.A(vliw_pc[1]), .B(vliw_pc[0]), .C(vliw_pc[2]), .Z(n_2790
		));
	notech_nand2 i_232(.A(vliw_pc[1]), .B(vliw_pc[0]), .Z(n_2789));
	notech_or4 i_6397(.A(n_272988726), .B(n_2588), .C(n_60563), .D(n_59380),
		 .Z(n_2788));
	notech_or4 i_1792(.A(n_2588), .B(n_60563), .C(n_62437), .D(n_272788728),
		 .Z(n_2787));
	notech_or4 i_418(.A(n_60762), .B(n_60719), .C(n_54899), .D(nbus_11273[7]
		), .Z(n_2786));
	notech_mux2 i_1003(.S(n_59890), .A(n_57418), .B(n_276288695), .Z(n_2785)
		);
	notech_and2 i_1004(.A(n_55195), .B(n_26616), .Z(n_2784));
	notech_ao4 i_1005(.A(n_57388), .B(n_59890), .C(n_276088697), .D(n_2596),
		 .Z(n_2783));
	notech_or4 i_1683(.A(n_2647), .B(n_60558), .C(n_62437), .D(n_272788728),
		 .Z(n_2782));
	notech_and3 i_1090(.A(n_2772), .B(n_2395), .C(n_2782), .Z(n_2781));
	notech_or2 i_509(.A(n_2777), .B(n_58895), .Z(n_2779));
	notech_or4 i_1589(.A(fsm[3]), .B(n_60735), .C(n_60761), .D(n_57388), .Z(n_2778
		));
	notech_and2 i_1378(.A(n_275288705), .B(n_273188724), .Z(n_2777));
	notech_or4 i_2119(.A(n_59355), .B(n_2647), .C(n_59380), .D(n_62395), .Z(n_2776
		));
	notech_nao3 i_1695(.A(n_28975), .B(n_60503), .C(n_2221), .Z(n_2775));
	notech_nao3 i_1712(.A(n_26785), .B(n_26792), .C(n_57383), .Z(n_2774));
	notech_and2 i_807(.A(n_274588712), .B(n_57383), .Z(n_2773));
	notech_or4 i_2089(.A(n_2647), .B(n_62395), .C(n_62437), .D(n_59958), .Z(n_2772
		));
	notech_nao3 i_330(.A(n_55389), .B(n_2387), .C(n_55159), .Z(n_2771));
	notech_nand3 i_979(.A(nbus_11326[3]), .B(nbus_11326[2]), .C(nbus_11326[4
		]), .Z(n_2770));
	notech_or4 i_1701(.A(n_273188724), .B(n_2550), .C(n_272988726), .D(n_2399
		), .Z(n_2769));
	notech_or4 i_1717(.A(n_273188724), .B(n_2550), .C(n_2399), .D(n_59958), 
		.Z(n_2768));
	notech_and2 i_897(.A(n_2394), .B(n_55525), .Z(n_276588692));
	notech_ao4 i_92970267(.A(n_494), .B(n_57434), .C(n_170914103), .D(n_57444
		), .Z(n_276488693));
	notech_nand3 i_46365(.A(n_206788846), .B(n_60748), .C(n_27262), .Z(n_276288695
		));
	notech_ao4 i_1132(.A(n_494), .B(n_57442), .C(n_2781), .D(n_60463), .Z(n_276188696
		));
	notech_nand3 i_32087(.A(n_26616), .B(n_57430), .C(n_59890), .Z(n_276088697
		));
	notech_nao3 i_32063(.A(n_26616), .B(n_59890), .C(n_57430), .Z(n_275988698
		));
	notech_or4 i_46373(.A(n_2582), .B(n_27265), .C(n_60735), .D(fsm[2]), .Z(n_275888699
		));
	notech_or4 i_46369(.A(n_60735), .B(n_2582), .C(n_60748), .D(n_27264), .Z
		(n_275788700));
	notech_nand3 i_7532790(.A(n_28975), .B(n_62419), .C(n_1942), .Z(n_2107)
		);
	notech_nao3 i_46360(.A(fsm[1]), .B(n_244356261), .C(n_60719), .Z(n_275688701
		));
	notech_or4 i_6832796(.A(n_2591), .B(n_275688701), .C(n_275588702), .D(n_59159
		), .Z(n_2113));
	notech_and4 i_46358(.A(fsm[1]), .B(n_244556263), .C(n_27264), .D(n_27266
		), .Z(n_275588702));
	notech_or4 i_177232822(.A(n_60577), .B(n_59828), .C(n_26862), .D(n_26497
		), .Z(n_2155));
	notech_nao3 i_167932828(.A(n_276288695), .B(n_274788710), .C(n_26625), .Z
		(n_2161));
	notech_or4 i_8132788(.A(n_59364), .B(n_2550), .C(n_2572), .D(n_59355), .Z
		(n_2105));
	notech_nand3 i_46361(.A(fsm[1]), .B(n_244356261), .C(n_244556263), .Z(n_57451
		));
	notech_or4 i_157232842(.A(n_275088707), .B(n_57451), .C(n_60577), .D(n_59828
		), .Z(n_2175));
	notech_or4 i_1118(.A(n_2793), .B(n_60577), .C(n_59817), .D(n_59771), .Z(n_494
		));
	notech_or4 i_157032843(.A(n_2793), .B(n_2222), .C(n_59771), .D(n_59159),
		 .Z(n_2176));
	notech_or4 i_134632849(.A(n_273288723), .B(n_275288705), .C(n_2258), .D(n_60463
		), .Z(n_2182));
	notech_nand3 i_119532857(.A(n_2575), .B(n_244056258), .C(n_57451), .Z(n_2190
		));
	notech_or4 i_115532858(.A(n_275388704), .B(n_60577), .C(n_59828), .D(n_59780
		), .Z(n_2191));
	notech_and2 i_113132862(.A(n_2196), .B(n_206488849), .Z(n_2195));
	notech_nao3 i_215(.A(n_62395), .B(n_62437), .C(n_2550), .Z(n_275488703)
		);
	notech_or2 i_499(.A(n_275088707), .B(n_2792), .Z(n_275388704));
	notech_nand2 i_197(.A(n_62395), .B(n_62437), .Z(n_275288705));
	notech_or4 i_46376(.A(n_2584), .B(n_27265), .C(n_27262), .D(fsm[2]), .Z(n_275188706
		));
	notech_or4 i_71932888(.A(n_2601), .B(n_2585), .C(n_2584), .D(n_2603), .Z
		(n_2222));
	notech_and2 i_139232891(.A(n_2195), .B(n_1950), .Z(n_2226));
	notech_nao3 i_25502(.A(n_275688701), .B(n_26497), .C(n_2591), .Z(n_275088707
		));
	notech_or4 i_21832921(.A(n_2038), .B(n_2035), .C(n_2031), .D(n_2028), .Z
		(n_22579221));
	notech_or2 i_172832929(.A(n_2221), .B(n_59355), .Z(n_2269));
	notech_nand2 i_94(.A(\opcode[3] ), .B(n_60503), .Z(n_274988708));
	notech_and4 i_162732975(.A(n_2406), .B(n_55763), .C(n_276488693), .D(n_54764
		), .Z(n_54818));
	notech_and4 i_70632976(.A(n_58886), .B(n_199688883), .C(n_211888826), .D
		(n_2779), .Z(n_55644));
	notech_ao4 i_52932901(.A(n_2251), .B(n_59958), .C(n_58931), .D(n_59762),
		 .Z(n_2236));
	notech_or2 i_172332930(.A(n_2386), .B(n_59355), .Z(n_2271));
	notech_or4 i_179832990(.A(n_2831), .B(n_2572), .C(n_273188724), .D(n_59958
		), .Z(n_57393));
	notech_or4 i_151832992(.A(n_60748), .B(n_60735), .C(n_60761), .D(n_192288896
		), .Z(n_54910));
	notech_or2 i_92532880(.A(n_190688899), .B(n_29040), .Z(n_2213));
	notech_nao3 i_46364(.A(fsm[1]), .B(n_27266), .C(n_2585), .Z(n_274788710)
		);
	notech_nand2 i_30832995(.A(n_59890), .B(n_26296), .Z(n_56041));
	notech_or4 i_153732996(.A(n_2831), .B(n_2572), .C(n_58940), .D(n_273288723
		), .Z(n_54894));
	notech_or4 i_32060(.A(n_28975), .B(n_2831), .C(n_2572), .D(n_62419), .Z(n_274688711
		));
	notech_nao3 i_213(.A(n_62437), .B(n_60558), .C(n_60490), .Z(n_274588712)
		);
	notech_nand3 i_2155(.A(n_62437), .B(n_60558), .C(n_55040), .Z(n_2268));
	notech_ao4 i_50632999(.A(n_273188724), .B(n_1911), .C(n_2260), .D(n_222356214
		), .Z(n_55843));
	notech_or4 i_30081(.A(n_28975), .B(n_60503), .C(n_59380), .D(\opcode[0] 
		), .Z(n_2325));
	notech_or4 i_102932872(.A(n_275388704), .B(n_60577), .C(n_59817), .D(n_59771
		), .Z(n_2205));
	notech_or4 i_29851(.A(n_60748), .B(n_60735), .C(n_60761), .D(eval_flag),
		 .Z(n_2327));
	notech_or2 i_2007(.A(n_1936), .B(n_56246), .Z(n_54505));
	notech_nao3 i_23532919(.A(n_56487), .B(n_56478), .C(n_56449), .Z(n_2255)
		);
	notech_nao3 i_1335(.A(n_60503), .B(n_26867), .C(n_28975), .Z(n_274488713
		));
	notech_nao3 i_126033006(.A(n_2174), .B(n_1984), .C(n_1985), .Z(n_57431)
		);
	notech_or4 i_155932844(.A(n_60761), .B(n_60719), .C(n_1900), .D(n_56551)
		, .Z(n_2177));
	notech_or2 i_1853(.A(n_59268), .B(n_28565), .Z(n_274388714));
	notech_nand2 i_1830(.A(n_59272), .B(n_28565), .Z(n_274288715));
	notech_or2 i_1812(.A(n_59272), .B(n_59263), .Z(n_274188716));
	notech_nao3 i_25725(.A(instrc[121]), .B(n_28566), .C(instrc[123]), .Z(n_2740
		));
	notech_nao3 i_25733(.A(n_28567), .B(n_28566), .C(instrc[123]), .Z(n_2739
		));
	notech_nao3 i_25722(.A(n_28567), .B(instrc[120]), .C(instrc[123]), .Z(n_273888717
		));
	notech_or4 i_49432904(.A(calc_sz[3]), .B(calc_sz[2]), .C(n_260688757), .D
		(n_56354), .Z(n_2239));
	notech_or2 i_49232906(.A(n_56569), .B(n_56354), .Z(n_2241));
	notech_or2 i_49332905(.A(n_56354), .B(n_56547), .Z(n_2240));
	notech_nand2 i_2031(.A(n_56487), .B(n_56478), .Z(n_2145));
	notech_nand3 i_129233040(.A(instrc[123]), .B(n_28566), .C(n_60525), .Z(n_55087
		));
	notech_or2 i_29532914(.A(n_56375), .B(n_60579), .Z(n_2250));
	notech_nao3 i_21933043(.A(calc_sz[1]), .B(calc_sz[0]), .C(n_2605), .Z(n_56107
		));
	notech_or4 i_145732846(.A(n_28975), .B(n_62419), .C(n_60558), .D(n_59380
		), .Z(n_2179));
	notech_nand3 i_98632876(.A(n_26785), .B(n_2042), .C(n_26621), .Z(n_2209)
		);
	notech_or4 i_152033049(.A(n_59364), .B(n_60490), .C(n_2572), .D(n_59958)
		, .Z(n_57419));
	notech_or4 i_151333050(.A(n_58940), .B(n_60490), .C(n_2572), .D(n_59958)
		, .Z(n_57420));
	notech_or4 i_25932915(.A(n_60490), .B(n_2572), .C(\opcode[0] ), .D(n_62437
		), .Z(n_2251));
	notech_nand2 i_199(.A(n_60558), .B(n_59375), .Z(n_273788718));
	notech_or4 i_103132871(.A(n_60762), .B(n_60719), .C(n_2647), .D(n_60577)
		, .Z(n_2204));
	notech_or4 i_2183(.A(n_28975), .B(n_2260), .C(n_59364), .D(n_62419), .Z(n_57376
		));
	notech_nao3 i_2171(.A(n_2042), .B(n_26867), .C(n_2352), .Z(n_57378));
	notech_or4 i_25609(.A(n_59375), .B(n_62395), .C(n_60503), .D(\opcode[3] 
		), .Z(n_2352));
	notech_nand3 i_2191(.A(n_2042), .B(n_26867), .C(n_26243), .Z(n_57374));
	notech_or4 i_114932859(.A(n_62395), .B(n_62437), .C(n_28975), .D(n_60504
		), .Z(n_2192));
	notech_or4 i_157332863(.A(n_60507), .B(\opcode[3] ), .C(n_60558), .D(n_59375
		), .Z(n_2196));
	notech_nand3 i_162132835(.A(n_2042), .B(n_26785), .C(n_27081), .Z(n_2168
		));
	notech_nao3 i_21732922(.A(n_2340), .B(n_26785), .C(n_26663), .Z(n_2258)
		);
	notech_nand3 i_46363(.A(fsm[1]), .B(n_244056258), .C(n_27266), .Z(n_273688719
		));
	notech_nand3 i_124333054(.A(n_59183), .B(n_59889), .C(n_59771), .Z(n_55131
		));
	notech_or2 i_60433055(.A(n_26616), .B(n_206688847), .Z(n_55745));
	notech_nand2 i_1811(.A(n_59272), .B(n_59263), .Z(n_273588720));
	notech_or4 i_173133062(.A(n_2258), .B(n_59355), .C(n_59762), .D(n_60463)
		, .Z(n_54733));
	notech_or4 i_157533065(.A(n_2258), .B(n_206188852), .C(reps[2]), .D(n_60463
		), .Z(n_54862));
	notech_and4 i_46379(.A(fsm[1]), .B(n_244356261), .C(n_60748), .D(n_60735
		), .Z(n_273488721));
	notech_or4 i_158533099(.A(n_59762), .B(n_60490), .C(n_59967), .D(n_273288723
		), .Z(n_57414));
	notech_or4 i_2394(.A(n_2647), .B(n_272988726), .C(n_59762), .D(n_60463),
		 .Z(n_57372));
	notech_or4 i_71633104(.A(n_2258), .B(n_273288723), .C(n_59201), .D(n_60463
		), .Z(n_55634));
	notech_nand2 i_5375(.A(nZF), .B(n_1947), .Z(n_51738));
	notech_or4 i_8747(.A(n_212988815), .B(n_60579), .C(n_59817), .D(n_26862)
		, .Z(n_48496));
	notech_or4 i_1495(.A(n_59201), .B(n_60490), .C(n_59967), .D(n_272988726)
		, .Z(n_273388722));
	notech_or4 i_70833105(.A(n_59141), .B(n_60579), .C(n_59889), .D(n_273388722
		), .Z(n_55642));
	notech_or4 i_72533106(.A(n_2205), .B(n_26296), .C(n_276288695), .D(n_1990
		), .Z(n_55625));
	notech_nand2 i_72733107(.A(reps[2]), .B(n_26620), .Z(n_55623));
	notech_nao3 i_69333108(.A(n_190488901), .B(n_26374), .C(n_206688847), .Z
		(n_55657));
	notech_or4 i_168733064(.A(n_2831), .B(n_58904), .C(n_59364), .D(n_60463)
		, .Z(n_54769));
	notech_or2 i_11170(.A(n_54505), .B(n_55958), .Z(n_46073));
	notech_nao3 i_21232924(.A(n_2385), .B(n_2042), .C(n_2361), .Z(n_2260));
	notech_nao3 i_24833128(.A(n_27517), .B(n_27518), .C(opz[2]), .Z(n_56079)
		);
	notech_nand2 i_196(.A(\opcode[3] ), .B(n_62419), .Z(n_273288723));
	notech_or4 i_8944(.A(n_28975), .B(n_59762), .C(n_2588), .D(n_60507), .Z(n_48299
		));
	notech_nao3 i_20933051(.A(n_60558), .B(n_59375), .C(n_60490), .Z(n_56117
		));
	notech_nao3 i_427964(.A(n_2500), .B(n_224756218), .C(n_227488799), .Z(\opcode[3] 
		));
	notech_ao4 i_38933002(.A(n_2044), .B(n_54520), .C(n_56375), .D(n_26242),
		 .Z(n_55960));
	notech_ao4 i_39133118(.A(n_2044), .B(n_56547), .C(n_55858), .D(n_26242),
		 .Z(n_55958));
	notech_nand3 i_169333164(.A(n_59183), .B(n_59889), .C(n_26862), .Z(n_54764
		));
	notech_or2 i_177433158(.A(n_205788856), .B(n_26599), .Z(n_54698));
	notech_nand2 i_195(.A(n_62437), .B(n_60558), .Z(n_273188724));
	notech_or4 i_2187(.A(n_28975), .B(n_2260), .C(n_59201), .D(n_62419), .Z(n_57375
		));
	notech_ao4 i_144868818(.A(n_27341992), .B(n_27349), .C(n_56409), .D(n_26953
		), .Z(n_112984456));
	notech_ao4 i_144768819(.A(n_26595), .B(n_356476400), .C(n_28442003), .D(n_27316
		), .Z(n_113084457));
	notech_ao4 i_138268884(.A(n_151260594), .B(n_27335), .C(n_334862246), .D
		(n_26927), .Z(n_113184458));
	notech_ao4 i_138168885(.A(n_56153), .B(n_29709), .C(n_170860790), .D(n_27300
		), .Z(n_113284459));
	notech_ao4 i_138068886(.A(n_151260594), .B(n_27336), .C(n_334862246), .D
		(n_26929), .Z(n_113384460));
	notech_ao4 i_137968887(.A(n_56153), .B(n_29708), .C(n_170860790), .D(n_27301
		), .Z(n_113484461));
	notech_ao4 i_137868888(.A(n_151260594), .B(n_27337), .C(n_334862246), .D
		(n_26931), .Z(n_113584462));
	notech_ao4 i_137768889(.A(n_56153), .B(n_29707), .C(n_170860790), .D(n_27302
		), .Z(n_113684463));
	notech_ao4 i_137668890(.A(n_151260594), .B(n_27338), .C(n_334862246), .D
		(n_26933), .Z(n_113784464));
	notech_ao4 i_137568891(.A(n_56153), .B(n_29706), .C(n_170860790), .D(n_27304
		), .Z(n_113884465));
	notech_ao4 i_137468892(.A(n_151260594), .B(n_27339), .C(n_334862246), .D
		(n_26935), .Z(n_113984466));
	notech_ao4 i_137368893(.A(n_56153), .B(n_29705), .C(n_170860790), .D(n_27307
		), .Z(n_114084467));
	notech_ao4 i_137268894(.A(n_151260594), .B(n_27340), .C(n_334862246), .D
		(n_26937), .Z(n_114184468));
	notech_ao4 i_137168895(.A(n_56153), .B(n_29704), .C(n_170860790), .D(n_27308
		), .Z(n_114284469));
	notech_ao4 i_137068896(.A(n_151260594), .B(n_27341), .C(n_334862246), .D
		(n_26939), .Z(n_114384470));
	notech_ao4 i_136968897(.A(n_56153), .B(n_29703), .C(n_170860790), .D(n_27309
		), .Z(n_114484471));
	notech_ao4 i_136868898(.A(n_151260594), .B(n_27342), .C(n_334862246), .D
		(n_26941), .Z(n_114584472));
	notech_ao4 i_136768899(.A(n_56153), .B(n_29702), .C(n_170860790), .D(n_27310
		), .Z(n_114684473));
	notech_ao4 i_136668900(.A(n_151260594), .B(n_27343), .C(n_334862246), .D
		(n_26943), .Z(n_114784474));
	notech_ao4 i_136568901(.A(n_56153), .B(n_29701), .C(n_170860790), .D(n_27311
		), .Z(n_114884475));
	notech_ao4 i_136468902(.A(n_151260594), .B(n_27345), .C(n_334862246), .D
		(n_26945), .Z(n_114984476));
	notech_ao4 i_136368903(.A(n_56153), .B(n_29700), .C(n_170860790), .D(n_27312
		), .Z(n_115084477));
	notech_ao4 i_136268904(.A(n_151260594), .B(n_27346), .C(n_334862246), .D
		(n_26947), .Z(n_115184478));
	notech_ao4 i_136168905(.A(n_56153), .B(n_29699), .C(n_170860790), .D(n_27313
		), .Z(n_115284479));
	notech_ao4 i_135968906(.A(n_151260594), .B(n_27347), .C(n_334862246), .D
		(n_26949), .Z(n_115384480));
	notech_ao4 i_135868907(.A(n_56153), .B(n_29698), .C(n_170860790), .D(n_27314
		), .Z(n_115484481));
	notech_ao4 i_135768908(.A(n_151260594), .B(n_27348), .C(n_334862246), .D
		(n_26951), .Z(n_115584482));
	notech_ao4 i_135668909(.A(n_56153), .B(n_29697), .C(n_170860790), .D(n_27315
		), .Z(n_115684483));
	notech_ao4 i_135568910(.A(n_151260594), .B(n_27349), .C(n_334862246), .D
		(n_26953), .Z(n_115784484));
	notech_ao4 i_135468911(.A(n_56153), .B(n_29696), .C(n_170860790), .D(n_27316
		), .Z(n_115884485));
	notech_ao4 i_135368912(.A(n_27350), .B(n_151260594), .C(n_56336), .D(n_26955
		), .Z(n_115984486));
	notech_ao4 i_135268913(.A(n_56153), .B(n_29695), .C(n_170860790), .D(n_27317
		), .Z(n_116084487));
	notech_ao4 i_135168914(.A(n_53113), .B(n_27351), .C(n_56336), .D(n_26957
		), .Z(n_116184488));
	notech_ao4 i_135068915(.A(n_53234), .B(n_29694), .C(n_53964), .D(n_27318
		), .Z(n_116284489));
	notech_ao4 i_134968916(.A(n_53113), .B(n_27352), .C(n_56336), .D(n_26959
		), .Z(n_116384490));
	notech_ao4 i_134868917(.A(n_53234), .B(n_29693), .C(n_53964), .D(n_27319
		), .Z(n_116484491));
	notech_ao4 i_134768918(.A(n_53113), .B(n_27353), .C(n_56336), .D(n_26961
		), .Z(n_116584492));
	notech_ao4 i_134668919(.A(n_53234), .B(n_29691), .C(n_53964), .D(n_27320
		), .Z(n_116684493));
	notech_ao4 i_134568920(.A(n_53113), .B(n_27354), .C(n_56336), .D(n_26963
		), .Z(n_116784494));
	notech_ao4 i_134468921(.A(n_53234), .B(n_29690), .C(n_53964), .D(n_27321
		), .Z(n_116884495));
	notech_ao4 i_134368922(.A(n_53113), .B(n_27355), .C(n_56336), .D(n_26965
		), .Z(n_116984496));
	notech_ao4 i_134268923(.A(n_53234), .B(n_29689), .C(n_53964), .D(n_27322
		), .Z(n_117084497));
	notech_ao4 i_134168924(.A(n_53113), .B(n_27356), .C(n_56336), .D(n_26967
		), .Z(n_117184498));
	notech_ao4 i_134068925(.A(n_53234), .B(n_29688), .C(n_53964), .D(n_27323
		), .Z(n_117284499));
	notech_ao4 i_133968926(.A(n_53113), .B(n_27357), .C(n_56336), .D(n_26969
		), .Z(n_117384500));
	notech_ao4 i_133868927(.A(n_53234), .B(n_29687), .C(n_53964), .D(n_27324
		), .Z(n_117484501));
	notech_ao4 i_133768928(.A(n_53113), .B(n_27358), .C(n_56336), .D(n_26971
		), .Z(n_117584502));
	notech_ao4 i_133668929(.A(n_53234), .B(n_29686), .C(n_53964), .D(n_27325
		), .Z(n_117684503));
	notech_ao4 i_133568930(.A(n_53113), .B(n_27359), .C(n_56336), .D(n_26973
		), .Z(n_117784504));
	notech_ao4 i_133468931(.A(n_53234), .B(n_29685), .C(n_53964), .D(n_27326
		), .Z(n_117884505));
	notech_ao4 i_133368932(.A(n_53113), .B(n_27360), .C(n_56336), .D(n_26975
		), .Z(n_117984506));
	notech_ao4 i_133268933(.A(n_53234), .B(n_29684), .C(n_53964), .D(n_27327
		), .Z(n_118084507));
	notech_ao4 i_133168934(.A(n_53113), .B(n_27361), .C(n_56336), .D(n_26977
		), .Z(n_118184508));
	notech_ao4 i_133068935(.A(n_53234), .B(n_29683), .C(n_170860790), .D(n_27328
		), .Z(n_118284509));
	notech_ao4 i_132968936(.A(n_53113), .B(n_27362), .C(n_56336), .D(n_26979
		), .Z(n_118384510));
	notech_ao4 i_132868937(.A(n_53234), .B(n_29682), .C(n_53964), .D(n_27329
		), .Z(n_118484511));
	notech_ao4 i_132768938(.A(n_53113), .B(n_27363), .C(n_56336), .D(n_26983
		), .Z(n_118584512));
	notech_ao4 i_132668939(.A(n_53234), .B(n_29681), .C(n_53964), .D(n_27330
		), .Z(n_118684513));
	notech_ao4 i_132568940(.A(n_27364), .B(n_53113), .C(n_56336), .D(n_26985
		), .Z(n_118784514));
	notech_ao4 i_132468941(.A(n_53234), .B(n_29680), .C(n_53964), .D(n_27331
		), .Z(n_118884515));
	notech_ao4 i_132368942(.A(n_53964), .B(n_27332), .C(n_27365), .D(n_53113
		), .Z(n_118984516));
	notech_ao4 i_132268943(.A(n_53234), .B(n_29679), .C(n_56336), .D(n_26987
		), .Z(n_119084517));
	notech_ao4 i_125969006(.A(n_27333), .B(n_150960591), .C(n_334762245), .D
		(n_26923), .Z(n_119184518));
	notech_ao4 i_125869007(.A(n_56150), .B(n_29678), .C(n_27297), .D(n_171160793
		), .Z(n_119284519));
	notech_ao4 i_125769008(.A(n_27334), .B(n_150960591), .C(n_334762245), .D
		(n_26925), .Z(n_119384520));
	notech_ao4 i_125669009(.A(n_56150), .B(n_29677), .C(n_171160793), .D(n_27298
		), .Z(n_119484521));
	notech_ao4 i_125569010(.A(n_27335), .B(n_150960591), .C(n_334762245), .D
		(n_26927), .Z(n_119584522));
	notech_ao4 i_125469011(.A(n_56150), .B(n_29676), .C(n_171160793), .D(n_27300
		), .Z(n_119684523));
	notech_ao4 i_125369012(.A(n_27336), .B(n_150960591), .C(n_334762245), .D
		(n_26929), .Z(n_119784524));
	notech_ao4 i_125269013(.A(n_56150), .B(n_29675), .C(n_171160793), .D(n_27301
		), .Z(n_119884525));
	notech_ao4 i_125169014(.A(n_27337), .B(n_150960591), .C(n_334762245), .D
		(n_26931), .Z(n_119984526));
	notech_ao4 i_125069015(.A(n_56150), .B(n_29674), .C(n_171160793), .D(n_27302
		), .Z(n_120084527));
	notech_ao4 i_124969016(.A(n_27338), .B(n_150960591), .C(n_334762245), .D
		(n_26933), .Z(n_120184528));
	notech_ao4 i_124869017(.A(n_56150), .B(n_29673), .C(n_171160793), .D(n_27304
		), .Z(n_120284529));
	notech_ao4 i_124769018(.A(n_27339), .B(n_150960591), .C(n_334762245), .D
		(n_26935), .Z(n_120384530));
	notech_ao4 i_124669019(.A(n_56150), .B(n_29672), .C(n_171160793), .D(n_27307
		), .Z(n_120484531));
	notech_ao4 i_124569020(.A(n_27340), .B(n_150960591), .C(n_334762245), .D
		(n_26937), .Z(n_120584532));
	notech_ao4 i_124469021(.A(n_56150), .B(n_29671), .C(n_171160793), .D(n_27308
		), .Z(n_120684533));
	notech_ao4 i_124369022(.A(n_27341), .B(n_150960591), .C(n_334762245), .D
		(n_26939), .Z(n_120784534));
	notech_ao4 i_124269023(.A(n_56150), .B(n_29670), .C(n_171160793), .D(n_27309
		), .Z(n_120884535));
	notech_ao4 i_124169024(.A(n_27342), .B(n_150960591), .C(n_334762245), .D
		(n_26941), .Z(n_120984536));
	notech_ao4 i_124069025(.A(n_56150), .B(n_29669), .C(n_171160793), .D(n_27310
		), .Z(n_121084537));
	notech_ao4 i_123969026(.A(n_27343), .B(n_150960591), .C(n_334762245), .D
		(n_26943), .Z(n_121184538));
	notech_ao4 i_123869027(.A(n_56150), .B(n_29668), .C(n_171160793), .D(n_27311
		), .Z(n_121284539));
	notech_ao4 i_123769028(.A(n_27345), .B(n_150960591), .C(n_334762245), .D
		(n_26945), .Z(n_121384540));
	notech_ao4 i_123669029(.A(n_56150), .B(n_29667), .C(n_171160793), .D(n_27312
		), .Z(n_121484541));
	notech_ao4 i_123569030(.A(n_27346), .B(n_150960591), .C(n_334762245), .D
		(n_26947), .Z(n_121584542));
	notech_ao4 i_123469031(.A(n_56150), .B(n_29666), .C(n_171160793), .D(n_27313
		), .Z(n_121684543));
	notech_ao4 i_123369032(.A(n_27347), .B(n_150960591), .C(n_334762245), .D
		(n_26949), .Z(n_121784544));
	notech_ao4 i_123269033(.A(n_56150), .B(n_29665), .C(n_171160793), .D(n_27314
		), .Z(n_121884545));
	notech_ao4 i_123169034(.A(n_27348), .B(n_150960591), .C(n_56511), .D(n_26951
		), .Z(n_121984546));
	notech_ao4 i_123069035(.A(n_56150), .B(n_29664), .C(n_171160793), .D(n_27315
		), .Z(n_122084547));
	notech_ao4 i_122969036(.A(n_27349), .B(n_52811), .C(n_56511), .D(n_26953
		), .Z(n_122184548));
	notech_ao4 i_122869037(.A(n_52930), .B(n_29663), .C(n_53937), .D(n_27316
		), .Z(n_122284549));
	notech_ao4 i_122569040(.A(n_27351), .B(n_52811), .C(n_56511), .D(n_26957
		), .Z(n_122384550));
	notech_ao4 i_122469041(.A(n_52930), .B(n_29662), .C(n_53937), .D(n_27318
		), .Z(n_122484551));
	notech_ao4 i_122369042(.A(n_27352), .B(n_52811), .C(n_56511), .D(n_26959
		), .Z(n_122584552));
	notech_ao4 i_122269043(.A(n_52930), .B(n_29661), .C(n_53937), .D(n_27319
		), .Z(n_122684553));
	notech_ao4 i_122169044(.A(n_27353), .B(n_52811), .C(n_56511), .D(n_26961
		), .Z(n_122784554));
	notech_ao4 i_122069045(.A(n_52930), .B(n_29660), .C(n_53937), .D(n_27320
		), .Z(n_122884555));
	notech_ao4 i_121969046(.A(n_27354), .B(n_52811), .C(n_56511), .D(n_26963
		), .Z(n_122984556));
	notech_ao4 i_121869047(.A(n_52930), .B(n_29659), .C(n_53937), .D(n_27321
		), .Z(n_123084557));
	notech_ao4 i_121769048(.A(n_27355), .B(n_52811), .C(n_56511), .D(n_26965
		), .Z(n_123184558));
	notech_ao4 i_121669049(.A(n_52930), .B(n_29658), .C(n_53937), .D(n_27322
		), .Z(n_123284559));
	notech_ao4 i_121569050(.A(n_27356), .B(n_52811), .C(n_56511), .D(n_26967
		), .Z(n_123384560));
	notech_ao4 i_121469051(.A(n_52930), .B(n_29657), .C(n_53937), .D(n_27323
		), .Z(n_123484561));
	notech_ao4 i_121369052(.A(n_27357), .B(n_52811), .C(n_56511), .D(n_26969
		), .Z(n_123584562));
	notech_ao4 i_121269053(.A(n_52930), .B(n_29656), .C(n_53937), .D(n_27324
		), .Z(n_123684563));
	notech_ao4 i_121069054(.A(n_27358), .B(n_52811), .C(n_56511), .D(n_26971
		), .Z(n_123784564));
	notech_ao4 i_120969055(.A(n_52930), .B(n_29655), .C(n_53937), .D(n_27325
		), .Z(n_123884565));
	notech_ao4 i_120869056(.A(n_27359), .B(n_52811), .C(n_56511), .D(n_26973
		), .Z(n_123984566));
	notech_ao4 i_120769057(.A(n_52930), .B(n_29654), .C(n_53937), .D(n_27326
		), .Z(n_124084567));
	notech_ao4 i_120669058(.A(n_27360), .B(n_150960591), .C(n_56511), .D(n_26975
		), .Z(n_124184568));
	notech_ao4 i_120569059(.A(n_52930), .B(n_29653), .C(n_171160793), .D(n_27327
		), .Z(n_124284569));
	notech_ao4 i_120469060(.A(n_27361), .B(n_52811), .C(n_56511), .D(n_26977
		), .Z(n_124384570));
	notech_ao4 i_120369061(.A(n_52930), .B(n_29652), .C(n_53937), .D(n_27328
		), .Z(n_124484571));
	notech_ao4 i_120269062(.A(n_27362), .B(n_52811), .C(n_56511), .D(n_26979
		), .Z(n_124584572));
	notech_ao4 i_120169063(.A(n_52930), .B(n_29651), .C(n_53937), .D(n_27329
		), .Z(n_124684573));
	notech_ao4 i_120069064(.A(n_27363), .B(n_52811), .C(n_56511), .D(n_26983
		), .Z(n_124784574));
	notech_ao4 i_119969065(.A(n_52930), .B(n_29650), .C(n_53937), .D(n_27330
		), .Z(n_124884575));
	notech_ao4 i_119869066(.A(n_27364), .B(n_52811), .C(n_56511), .D(n_26985
		), .Z(n_124984576));
	notech_ao4 i_119769067(.A(n_52930), .B(n_29649), .C(n_53937), .D(n_27331
		), .Z(n_125084577));
	notech_and3 i_168273(.A(n_57380), .B(n_57423), .C(n_2781), .Z(n_125384580
		));
	notech_ao4 i_52383(.A(n_125384580), .B(n_60463), .C(n_55745), .D(n_321731604
		), .Z(\nbus_11334[0] ));
	notech_or4 i_2768247(.A(n_60602), .B(n_272988726), .C(n_58940), .D(n_60463
		), .Z(n_125484581));
	notech_nand2 i_47393(.A(n_125484581), .B(n_55657), .Z(n_9351));
	notech_or4 i_2968245(.A(n_60602), .B(n_272988726), .C(n_59364), .D(n_60463
		), .Z(n_125584582));
	notech_nand2 i_47316(.A(n_125584582), .B(n_55657), .Z(n_9257));
	notech_or4 i_3168243(.A(n_60602), .B(n_59201), .C(n_60463), .D(n_59210),
		 .Z(n_125684583));
	notech_nand2 i_48680(.A(n_125684583), .B(n_55657), .Z(n_11506));
	notech_or4 i_3368241(.A(n_60602), .B(n_2352), .C(n_60579), .D(n_59889), 
		.Z(n_125784584));
	notech_nand2 i_51299(.A(n_125784584), .B(n_55657), .Z(n_15204));
	notech_or4 i_3568239(.A(n_60602), .B(n_2196), .C(n_60577), .D(n_59889), 
		.Z(n_125884585));
	notech_nand2 i_47956(.A(n_125884585), .B(n_55657), .Z(n_10208));
	notech_or4 i_3868236(.A(n_60761), .B(n_60719), .C(n_126084587), .D(n_60577
		), .Z(n_125984586));
	notech_and4 i_268272(.A(n_57387), .B(n_54741), .C(n_57388), .D(n_57402),
		 .Z(n_126084587));
	notech_nand2 i_46218(.A(n_181485140), .B(n_125984586), .Z(n_7415));
	notech_ao4 i_46986(.A(n_35657), .B(n_60463), .C(n_56547), .D(n_54968), .Z
		(n_8785));
	notech_or4 i_4768227(.A(n_60761), .B(n_60719), .C(n_57387), .D(n_60577),
		 .Z(n_126284589));
	notech_nand2 i_51159(.A(n_300586325), .B(n_126284589), .Z(n_14930));
	notech_ao4 i_50990(.A(n_323688454), .B(n_60463), .C(n_206688847), .D(n_26616
		), .Z(n_14738));
	notech_or4 i_6468210(.A(n_28975), .B(n_2204), .C(n_2264), .D(n_62395), .Z
		(n_126384590));
	notech_or4 i_6268212(.A(n_60577), .B(n_59890), .C(n_26600), .D(n_276588692
		), .Z(n_126484591));
	notech_and4 i_6368211(.A(read_ack), .B(mask8b[2]), .C(n_26554), .D(n_26862
		), .Z(n_126584592));
	notech_nao3 i_48597(.A(n_126384590), .B(n_126484591), .C(n_126584592), .Z
		(\nbus_11302[0] ));
	notech_ao4 i_53371(.A(n_206688847), .B(n_26616), .C(n_54914), .D(n_60463
		), .Z(n_18841));
	notech_nand2 i_51019(.A(n_55745), .B(n_54896), .Z(n_14770));
	notech_or4 i_47350(.A(n_60577), .B(n_59817), .C(n_14770), .D(n_26601), .Z
		(\nbus_11283[0] ));
	notech_ao3 i_10868172(.A(n_26380), .B(read_ack), .C(n_107542794), .Z(n_126784594
		));
	notech_or2 i_51332(.A(n_126784594), .B(n_353288276), .Z(\nbus_11327[0] )
		);
	notech_nand3 i_52868(.A(n_55642), .B(n_55745), .C(n_182485150), .Z(\nbus_11341[0] 
		));
	notech_or4 i_11568165(.A(n_60540), .B(n_2204), .C(n_60558), .D(n_56260),
		 .Z(n_126984596));
	notech_nand2 i_52422(.A(n_55745), .B(n_126984596), .Z(n_17010));
	notech_and4 i_12668162(.A(n_2042), .B(n_26867), .C(n_26666), .D(n_26621)
		, .Z(n_127084597));
	notech_nao3 i_51189(.A(n_55745), .B(n_238685706), .C(n_127084597), .Z(n_14963
		));
	notech_or4 i_12968159(.A(n_2258), .B(n_60586), .C(n_59890), .D(n_55086),
		 .Z(n_127184598));
	notech_nand3 i_46422(.A(n_55808), .B(n_55745), .C(n_127184598), .Z(n_7558
		));
	notech_nand2 i_46353(.A(n_55625), .B(n_300286322), .Z(n_7511));
	notech_or4 i_21868073(.A(n_52251), .B(n_52370), .C(from_acu[3]), .D(n_27958
		), .Z(n_127384600));
	notech_or4 i_21368078(.A(from_acu[3]), .B(from_acu[2]), .C(n_52370), .D(n_27891
		), .Z(n_128084607));
	notech_nand2 i_611983(.A(n_184085166), .B(n_127384600), .Z(to_acu[5]));
	notech_or4 i_29467998(.A(n_52251), .B(n_52370), .C(from_acu[3]), .D(n_27963
		), .Z(n_128184608));
	notech_or4 i_28968003(.A(from_acu[3]), .B(from_acu[2]), .C(n_52370), .D(n_27897
		), .Z(n_128884615));
	notech_nand2 i_1111988(.A(n_184685172), .B(n_128184608), .Z(to_acu[10])
		);
	notech_or4 i_33967953(.A(n_52251), .B(n_52370), .C(from_acu[3]), .D(n_27966
		), .Z(n_128984616));
	notech_or4 i_33467958(.A(from_acu[3]), .B(from_acu[2]), .C(n_52370), .D(n_27900
		), .Z(n_129684623));
	notech_nand2 i_1411991(.A(n_185285178), .B(n_128984616), .Z(to_acu[13])
		);
	notech_or4 i_35467938(.A(n_52251), .B(n_52370), .C(from_acu[3]), .D(n_27967
		), .Z(n_129784624));
	notech_or4 i_34967943(.A(from_acu[3]), .B(from_acu[2]), .C(n_52370), .D(n_27901
		), .Z(n_130484631));
	notech_nand2 i_1511992(.A(n_185885184), .B(n_129784624), .Z(to_acu[14])
		);
	notech_or4 i_36967923(.A(n_52250), .B(n_52369), .C(from_acu[3]), .D(n_27968
		), .Z(n_130584632));
	notech_or4 i_36467928(.A(from_acu[3]), .B(from_acu[2]), .C(n_52369), .D(n_27902
		), .Z(n_131284639));
	notech_nand2 i_1611993(.A(n_130584632), .B(n_186485190), .Z(to_acu[15])
		);
	notech_or4 i_38467908(.A(n_52250), .B(n_52369), .C(from_acu[3]), .D(n_27969
		), .Z(n_131384640));
	notech_or4 i_37967913(.A(from_acu[3]), .B(from_acu[2]), .C(n_52369), .D(n_27903
		), .Z(n_132084647));
	notech_nand2 i_1711994(.A(n_187085196), .B(n_131384640), .Z(to_acu[16])
		);
	notech_or4 i_39967893(.A(n_52250), .B(n_52369), .C(from_acu[3]), .D(n_27970
		), .Z(n_132184648));
	notech_or4 i_39467898(.A(from_acu[3]), .B(from_acu[2]), .C(n_52369), .D(n_27904
		), .Z(n_132884655));
	notech_nand2 i_1811995(.A(n_187685202), .B(n_132184648), .Z(to_acu[17])
		);
	notech_or4 i_41467878(.A(n_52250), .B(n_52369), .C(from_acu[3]), .D(n_27971
		), .Z(n_132984656));
	notech_or4 i_40967883(.A(from_acu[3]), .B(from_acu[2]), .C(n_52369), .D(n_27905
		), .Z(n_133684663));
	notech_nand2 i_1911996(.A(n_188285208), .B(n_132984656), .Z(to_acu[18])
		);
	notech_or4 i_42967863(.A(n_52253), .B(n_52372), .C(from_acu[3]), .D(n_27972
		), .Z(n_133784664));
	notech_or4 i_42467868(.A(from_acu[3]), .B(from_acu[2]), .C(n_52372), .D(n_27906
		), .Z(n_134484671));
	notech_nand2 i_2011997(.A(n_188885214), .B(n_133784664), .Z(to_acu[19])
		);
	notech_or4 i_44467848(.A(n_52253), .B(n_52372), .C(from_acu[3]), .D(n_27973
		), .Z(n_134584672));
	notech_or4 i_43967853(.A(from_acu[3]), .B(from_acu[2]), .C(n_52372), .D(n_27907
		), .Z(n_135284679));
	notech_nand2 i_2111998(.A(n_189485220), .B(n_134584672), .Z(to_acu[20])
		);
	notech_or4 i_45967833(.A(n_52253), .B(n_52372), .C(from_acu[3]), .D(n_27974
		), .Z(n_135384680));
	notech_or4 i_45467838(.A(from_acu[3]), .B(from_acu[2]), .C(n_52372), .D(n_27908
		), .Z(n_136084687));
	notech_nand2 i_2211999(.A(n_190085226), .B(n_135384680), .Z(to_acu[21])
		);
	notech_or4 i_47467818(.A(n_52253), .B(n_52372), .C(from_acu[3]), .D(n_27975
		), .Z(n_136184688));
	notech_or4 i_46967823(.A(from_acu[3]), .B(from_acu[2]), .C(n_52372), .D(n_27909
		), .Z(n_136884695));
	notech_nand2 i_2312000(.A(n_190685232), .B(n_136184688), .Z(to_acu[22])
		);
	notech_or4 i_49067803(.A(n_52252), .B(n_52371), .C(from_acu[3]), .D(n_27976
		), .Z(n_136984696));
	notech_or4 i_48467808(.A(from_acu[3]), .B(from_acu[2]), .C(n_52371), .D(n_27910
		), .Z(n_137684703));
	notech_nand2 i_2412001(.A(n_191285238), .B(n_136984696), .Z(to_acu[23])
		);
	notech_or4 i_50567788(.A(from_acu[3]), .B(n_52252), .C(n_52371), .D(n_27977
		), .Z(n_137784704));
	notech_or4 i_50067793(.A(from_acu[3]), .B(from_acu[2]), .C(n_52371), .D(n_27911
		), .Z(n_138484711));
	notech_nand2 i_2512002(.A(n_191885244), .B(n_137784704), .Z(to_acu[24])
		);
	notech_or4 i_52067773(.A(n_52252), .B(n_52371), .C(from_acu[3]), .D(n_27978
		), .Z(n_138584712));
	notech_or4 i_51567778(.A(from_acu[3]), .B(from_acu[2]), .C(n_52371), .D(n_27912
		), .Z(n_139284719));
	notech_nand2 i_2612003(.A(n_192485250), .B(n_138584712), .Z(to_acu[25])
		);
	notech_or4 i_53567758(.A(n_52252), .B(n_52371), .C(from_acu[3]), .D(n_27979
		), .Z(n_139384720));
	notech_or4 i_53067763(.A(from_acu[3]), .B(from_acu[2]), .C(n_52371), .D(n_27913
		), .Z(n_140084727));
	notech_nand2 i_2712004(.A(n_193085256), .B(n_139384720), .Z(to_acu[26])
		);
	notech_or4 i_55067743(.A(n_52246), .B(n_52365), .C(from_acu[3]), .D(n_27980
		), .Z(n_140184728));
	notech_or4 i_54567748(.A(from_acu[3]), .B(from_acu[2]), .C(n_52365), .D(n_27914
		), .Z(n_140884735));
	notech_nand2 i_2812005(.A(n_193685262), .B(n_140184728), .Z(to_acu[27])
		);
	notech_or4 i_56567728(.A(n_52246), .B(n_52365), .C(from_acu[3]), .D(n_27981
		), .Z(n_140984736));
	notech_or4 i_56067733(.A(from_acu[3]), .B(from_acu[2]), .C(n_52365), .D(n_27915
		), .Z(n_141684743));
	notech_nand2 i_2912006(.A(n_194285268), .B(n_140984736), .Z(to_acu[28])
		);
	notech_or4 i_58067713(.A(n_52246), .B(n_52365), .C(from_acu[3]), .D(n_27982
		), .Z(n_141784744));
	notech_or4 i_57567718(.A(from_acu[3]), .B(from_acu[2]), .C(n_52365), .D(n_27916
		), .Z(n_142484751));
	notech_nand2 i_3012007(.A(n_194885274), .B(n_141784744), .Z(to_acu[29])
		);
	notech_or4 i_61067683(.A(n_52246), .B(n_52365), .C(from_acu[3]), .D(n_27984
		), .Z(n_142584752));
	notech_or4 i_60567688(.A(from_acu[3]), .B(from_acu[2]), .C(n_52365), .D(n_27918
		), .Z(n_143284759));
	notech_nand2 i_3212009(.A(n_195485280), .B(n_142584752), .Z(to_acu[31])
		);
	notech_or4 i_62767666(.A(n_52442), .B(n_52453), .C(from_acu[7]), .D(n_27953
		), .Z(n_143384760));
	notech_or4 i_62167672(.A(from_acu[7]), .B(from_acu[6]), .C(n_52453), .D(n_27885
		), .Z(n_144084767));
	notech_nand2 i_112234(.A(n_197585301), .B(n_143384760), .Z(to_acu[32])
		);
	notech_or4 i_64267651(.A(n_52442), .B(n_52453), .C(from_acu[7]), .D(n_27954
		), .Z(n_144184768));
	notech_or4 i_63667657(.A(from_acu[7]), .B(from_acu[6]), .C(n_52453), .D(n_27886
		), .Z(n_144884775));
	notech_nand2 i_212235(.A(n_198185307), .B(n_144184768), .Z(to_acu[33])
		);
	notech_or4 i_65767636(.A(n_52442), .B(n_52453), .C(from_acu[7]), .D(n_27955
		), .Z(n_144984776));
	notech_or4 i_65167642(.A(from_acu[7]), .B(from_acu[6]), .C(n_52453), .D(n_27887
		), .Z(n_145684783));
	notech_nand2 i_312236(.A(n_198785313), .B(n_144984776), .Z(to_acu[34])
		);
	notech_or4 i_67267621(.A(n_52442), .B(n_52453), .C(from_acu[7]), .D(n_27956
		), .Z(n_145784784));
	notech_or4 i_66667627(.A(from_acu[7]), .B(from_acu[6]), .C(n_52453), .D(n_27888
		), .Z(n_146484791));
	notech_nand2 i_412237(.A(n_199385319), .B(n_145784784), .Z(to_acu[35])
		);
	notech_or4 i_68767606(.A(n_52441), .B(n_52452), .C(from_acu[7]), .D(n_27957
		), .Z(n_146584792));
	notech_or4 i_68167612(.A(from_acu[7]), .B(from_acu[6]), .C(n_52452), .D(n_27889
		), .Z(n_147284799));
	notech_nand2 i_512238(.A(n_199985325), .B(n_146584792), .Z(to_acu[36])
		);
	notech_or4 i_70267591(.A(n_52441), .B(n_52452), .C(from_acu[7]), .D(n_27958
		), .Z(n_147384800));
	notech_or4 i_69667597(.A(from_acu[7]), .B(from_acu[6]), .C(n_52452), .D(n_27891
		), .Z(n_148084807));
	notech_nand2 i_612239(.A(n_200585331), .B(n_147384800), .Z(to_acu[37])
		);
	notech_or4 i_71767576(.A(n_52441), .B(n_52452), .C(from_acu[7]), .D(n_27959
		), .Z(n_148184808));
	notech_or4 i_71167582(.A(from_acu[7]), .B(from_acu[6]), .C(n_52452), .D(n_27893
		), .Z(n_148884815));
	notech_nand2 i_712240(.A(n_201185337), .B(n_148184808), .Z(to_acu[38])
		);
	notech_or4 i_73267561(.A(n_52441), .B(n_52452), .C(from_acu[7]), .D(n_27960
		), .Z(n_148984816));
	notech_or4 i_72667567(.A(from_acu[7]), .B(from_acu[6]), .C(n_52452), .D(n_27894
		), .Z(n_149684823));
	notech_nand2 i_812241(.A(n_201785343), .B(n_148984816), .Z(to_acu[39])
		);
	notech_or4 i_74767546(.A(n_52444), .B(n_52455), .C(from_acu[7]), .D(n_27961
		), .Z(n_149784824));
	notech_or4 i_74167552(.A(from_acu[7]), .B(from_acu[6]), .C(n_52455), .D(n_27895
		), .Z(n_150484831));
	notech_nand2 i_912242(.A(n_202385349), .B(n_149784824), .Z(to_acu[40])
		);
	notech_or4 i_76267531(.A(n_52444), .B(n_52455), .C(from_acu[7]), .D(n_27962
		), .Z(n_150584832));
	notech_or4 i_75667537(.A(from_acu[7]), .B(from_acu[6]), .C(n_52455), .D(n_27896
		), .Z(n_151284839));
	notech_nand2 i_1012243(.A(n_202985355), .B(n_150584832), .Z(to_acu[41])
		);
	notech_or4 i_77767516(.A(n_52444), .B(n_52455), .C(from_acu[7]), .D(n_27963
		), .Z(n_151384840));
	notech_or4 i_77167522(.A(from_acu[7]), .B(from_acu[6]), .C(n_52455), .D(n_27897
		), .Z(n_152084847));
	notech_nand2 i_1112244(.A(n_203585361), .B(n_151384840), .Z(to_acu[42])
		);
	notech_or4 i_79267501(.A(n_52444), .B(n_52455), .C(from_acu[7]), .D(n_27964
		), .Z(n_152184848));
	notech_or4 i_78667507(.A(from_acu[7]), .B(from_acu[6]), .C(n_52455), .D(n_27898
		), .Z(n_152884855));
	notech_nand2 i_1212245(.A(n_204185367), .B(n_152184848), .Z(to_acu[43])
		);
	notech_or4 i_80767486(.A(n_52443), .B(n_52454), .C(from_acu[7]), .D(n_27965
		), .Z(n_152984856));
	notech_or4 i_80167492(.A(from_acu[7]), .B(from_acu[6]), .C(n_52454), .D(n_27899
		), .Z(n_153684863));
	notech_nand2 i_1312246(.A(n_204785373), .B(n_152984856), .Z(to_acu[44])
		);
	notech_or4 i_82267471(.A(n_52443), .B(n_52454), .C(from_acu[7]), .D(n_27966
		), .Z(n_153784864));
	notech_or4 i_81667477(.A(from_acu[7]), .B(from_acu[6]), .C(n_52454), .D(n_27900
		), .Z(n_154484871));
	notech_nand2 i_1412247(.A(n_205385379), .B(n_153784864), .Z(to_acu[45])
		);
	notech_or4 i_83767456(.A(n_52443), .B(n_52454), .C(from_acu[7]), .D(n_27967
		), .Z(n_154584872));
	notech_or4 i_83167462(.A(from_acu[7]), .B(from_acu[6]), .C(n_52454), .D(n_27901
		), .Z(n_155284879));
	notech_nand2 i_1512248(.A(n_205985385), .B(n_154584872), .Z(to_acu[46])
		);
	notech_or4 i_85267441(.A(n_52443), .B(n_52454), .C(from_acu[7]), .D(n_27968
		), .Z(n_155384880));
	notech_or4 i_84667447(.A(from_acu[7]), .B(from_acu[6]), .C(n_52454), .D(n_27902
		), .Z(n_156084887));
	notech_nand2 i_1612249(.A(n_155384880), .B(n_206585391), .Z(to_acu[47])
		);
	notech_or4 i_86767426(.A(n_52437), .B(n_52448), .C(from_acu[7]), .D(n_27969
		), .Z(n_156184888));
	notech_or4 i_86167432(.A(from_acu[7]), .B(from_acu[6]), .C(n_52448), .D(n_27903
		), .Z(n_156884895));
	notech_nand2 i_1712250(.A(n_207185397), .B(n_156184888), .Z(to_acu[48])
		);
	notech_or4 i_88267411(.A(n_52437), .B(n_52448), .C(from_acu[7]), .D(n_27970
		), .Z(n_156984896));
	notech_or4 i_87667417(.A(from_acu[7]), .B(from_acu[6]), .C(n_52448), .D(n_27904
		), .Z(n_157684903));
	notech_nand2 i_1812251(.A(n_207785403), .B(n_156984896), .Z(to_acu[49])
		);
	notech_or4 i_89767396(.A(n_52437), .B(n_52448), .C(from_acu[7]), .D(n_27971
		), .Z(n_157784904));
	notech_or4 i_89167402(.A(from_acu[7]), .B(from_acu[6]), .C(n_52448), .D(n_27905
		), .Z(n_158484911));
	notech_nand2 i_1912252(.A(n_208385409), .B(n_157784904), .Z(to_acu[50])
		);
	notech_or4 i_91267381(.A(n_52437), .B(n_52448), .C(from_acu[7]), .D(n_27972
		), .Z(n_158584912));
	notech_or4 i_90667387(.A(from_acu[7]), .B(from_acu[6]), .C(n_52448), .D(n_27906
		), .Z(n_159284919));
	notech_nand2 i_2012253(.A(n_208985415), .B(n_158584912), .Z(to_acu[51])
		);
	notech_or4 i_92767366(.A(n_52436), .B(n_52447), .C(from_acu[7]), .D(n_27973
		), .Z(n_159384920));
	notech_or4 i_92167372(.A(from_acu[7]), .B(from_acu[6]), .C(n_52447), .D(n_27907
		), .Z(n_160084927));
	notech_nand2 i_2112254(.A(n_209585421), .B(n_159384920), .Z(to_acu[52])
		);
	notech_or4 i_94267351(.A(n_52436), .B(n_52447), .C(from_acu[7]), .D(n_27974
		), .Z(n_160184928));
	notech_or4 i_93667357(.A(from_acu[7]), .B(from_acu[6]), .C(n_52447), .D(n_27908
		), .Z(n_160884935));
	notech_nand2 i_2212255(.A(n_210185427), .B(n_160184928), .Z(to_acu[53])
		);
	notech_or4 i_95767336(.A(n_52436), .B(n_52447), .C(from_acu[7]), .D(n_27975
		), .Z(n_160984936));
	notech_or4 i_95167342(.A(from_acu[7]), .B(from_acu[6]), .C(n_52447), .D(n_27909
		), .Z(n_161684943));
	notech_nand2 i_2312256(.A(n_210785433), .B(n_160984936), .Z(to_acu[54])
		);
	notech_or4 i_97267321(.A(n_52436), .B(n_52447), .C(from_acu[7]), .D(n_27976
		), .Z(n_161784944));
	notech_or4 i_96667327(.A(from_acu[7]), .B(from_acu[6]), .C(n_52447), .D(n_27910
		), .Z(n_162484951));
	notech_nand2 i_2412257(.A(n_211385439), .B(n_161784944), .Z(to_acu[55])
		);
	notech_or4 i_98767306(.A(from_acu[7]), .B(n_52439), .C(n_52450), .D(n_27977
		), .Z(n_162584952));
	notech_or4 i_98167312(.A(from_acu[7]), .B(from_acu[6]), .C(n_52450), .D(n_27911
		), .Z(n_163284959));
	notech_nand2 i_2512258(.A(n_211985445), .B(n_162584952), .Z(to_acu[56])
		);
	notech_or4 i_100267291(.A(n_52439), .B(n_52450), .C(from_acu[7]), .D(n_27978
		), .Z(n_163384960));
	notech_or4 i_99667297(.A(from_acu[7]), .B(from_acu[6]), .C(n_52450), .D(n_27912
		), .Z(n_164084967));
	notech_nand2 i_2612259(.A(n_212585451), .B(n_163384960), .Z(to_acu[57])
		);
	notech_or4 i_101767276(.A(n_52439), .B(n_52450), .C(from_acu[7]), .D(n_27979
		), .Z(n_164184968));
	notech_or4 i_101167282(.A(from_acu[7]), .B(from_acu[6]), .C(n_52450), .D
		(n_27913), .Z(n_164884975));
	notech_nand2 i_2712260(.A(n_213185457), .B(n_164184968), .Z(to_acu[58])
		);
	notech_or4 i_103367261(.A(n_52439), .B(n_52450), .C(from_acu[7]), .D(n_27980
		), .Z(n_164984976));
	notech_or4 i_102667267(.A(from_acu[7]), .B(from_acu[6]), .C(n_52450), .D
		(n_27914), .Z(n_165684983));
	notech_nand2 i_2812261(.A(n_213785463), .B(n_164984976), .Z(to_acu[59])
		);
	notech_or4 i_104867246(.A(n_52438), .B(n_52449), .C(from_acu[7]), .D(n_27981
		), .Z(n_165784984));
	notech_or4 i_104267252(.A(from_acu[7]), .B(from_acu[6]), .C(n_52449), .D
		(n_27915), .Z(n_166484991));
	notech_nand2 i_2912262(.A(n_214385469), .B(n_165784984), .Z(to_acu[60])
		);
	notech_or4 i_106367231(.A(n_52438), .B(n_52449), .C(from_acu[7]), .D(n_27982
		), .Z(n_166584992));
	notech_or4 i_105767237(.A(from_acu[7]), .B(from_acu[6]), .C(n_52449), .D
		(n_27916), .Z(n_167284999));
	notech_nand2 i_3012263(.A(n_214985475), .B(n_166584992), .Z(to_acu[61])
		);
	notech_or4 i_107867216(.A(n_52438), .B(n_52449), .C(from_acu[7]), .D(n_27983
		), .Z(n_167385000));
	notech_or4 i_107267222(.A(from_acu[7]), .B(from_acu[6]), .C(n_52449), .D
		(n_27917), .Z(n_168085007));
	notech_nand2 i_3112264(.A(n_215585481), .B(n_167385000), .Z(to_acu[62])
		);
	notech_or4 i_109367201(.A(n_52438), .B(n_52449), .C(from_acu[7]), .D(n_27984
		), .Z(n_168185008));
	notech_or4 i_108767207(.A(from_acu[7]), .B(from_acu[6]), .C(n_52449), .D
		(n_27918), .Z(n_168885015));
	notech_nand2 i_3212265(.A(n_216185487), .B(n_168185008), .Z(to_acu[63])
		);
	notech_nand2 i_117803(.A(n_216385489), .B(n_216285488), .Z(write_data_26
		[0]));
	notech_nand2 i_317805(.A(n_216585491), .B(n_216485490), .Z(write_data_26
		[2]));
	notech_nand2 i_417806(.A(n_216785493), .B(n_216685492), .Z(write_data_26
		[3]));
	notech_nand2 i_517807(.A(n_216985495), .B(n_216885494), .Z(write_data_26
		[4]));
	notech_nand2 i_617808(.A(n_217185497), .B(n_217085496), .Z(write_data_26
		[5]));
	notech_nand2 i_817810(.A(n_217385499), .B(n_217285498), .Z(write_data_26
		[7]));
	notech_nand2 i_1817820(.A(n_217585501), .B(n_217485500), .Z(write_data_26
		[17]));
	notech_nand2 i_2517827(.A(n_217785503), .B(n_217685502), .Z(write_data_26
		[24]));
	notech_nand2 i_3017832(.A(n_217985505), .B(n_217885504), .Z(write_data_26
		[29]));
	notech_nand2 i_123667058(.A(opa[7]), .B(n_26592), .Z(n_172585052));
	notech_nand2 i_6486(.A(n_218485510), .B(n_172585052), .Z(n_18226));
	notech_or2 i_124167053(.A(n_55282), .B(n_56551), .Z(n_172885055));
	notech_and2 i_1168263(.A(n_218585511), .B(n_172885055), .Z(n_173285059)
		);
	notech_ao4 i_6497(.A(CFOF_mul), .B(n_57387), .C(n_57417), .D(n_173285059
		), .Z(n_14933));
	notech_nand2 i_323103(.A(n_54881), .B(n_218785513), .Z(n_11427));
	notech_ao4 i_223102(.A(n_218785513), .B(n_55331), .C(n_54881), .D(n_59753
		), .Z(n_11421));
	notech_ao4 i_123101(.A(n_218785513), .B(n_55342), .C(n_54881), .D(n_55356
		), .Z(n_11415));
	notech_nand2 i_134966945(.A(n_55758), .B(opb[21]), .Z(n_174385070));
	notech_nand3 i_2218624(.A(n_218985515), .B(n_218885514), .C(n_174385070)
		, .Z(n_18361));
	notech_nand2 i_135866936(.A(n_55758), .B(opb[20]), .Z(n_174885075));
	notech_nand3 i_2118623(.A(n_219285518), .B(n_219185517), .C(n_174885075)
		, .Z(n_18356));
	notech_nand2 i_136766927(.A(n_55758), .B(opb[19]), .Z(n_175385080));
	notech_nand3 i_2018622(.A(n_219585521), .B(n_219485520), .C(n_175385080)
		, .Z(n_18351));
	notech_nand2 i_137666918(.A(n_55758), .B(opb[18]), .Z(n_175885085));
	notech_nand3 i_1918621(.A(n_219985524), .B(n_219885523), .C(n_175885085)
		, .Z(n_18346));
	notech_nand2 i_138566909(.A(n_55758), .B(opb[17]), .Z(n_176385090));
	notech_nand3 i_1818620(.A(n_220285527), .B(n_220185526), .C(n_176385090)
		, .Z(n_18341));
	notech_nand2 i_139466900(.A(n_55758), .B(opb[16]), .Z(n_176885095));
	notech_nand3 i_1718619(.A(n_220685530), .B(n_220585529), .C(n_176885095)
		, .Z(n_18336));
	notech_nand2 i_140366891(.A(opb[14]), .B(n_264885968), .Z(n_177385100)
		);
	notech_nand3 i_1518617(.A(n_221085533), .B(n_220885532), .C(n_177385100)
		, .Z(n_18326));
	notech_nand2 i_141266882(.A(opb[13]), .B(n_264885968), .Z(n_177885105)
		);
	notech_nand3 i_1418616(.A(n_221385536), .B(n_221285535), .C(n_177885105)
		, .Z(n_18321));
	notech_nand2 i_142266873(.A(opb[12]), .B(n_264885968), .Z(n_178385110)
		);
	notech_nand3 i_1318615(.A(n_221685539), .B(n_221585538), .C(n_178385110)
		, .Z(n_18316));
	notech_nand2 i_143166864(.A(opb[11]), .B(n_264885968), .Z(n_178985115)
		);
	notech_nand3 i_1218614(.A(n_221985542), .B(n_221885541), .C(n_178985115)
		, .Z(n_18311));
	notech_nand2 i_144066855(.A(opb[10]), .B(n_264885968), .Z(n_179485120)
		);
	notech_nand3 i_1118613(.A(n_222285545), .B(n_222185544), .C(n_179485120)
		, .Z(n_18306));
	notech_nand2 i_144966846(.A(opb[9]), .B(n_264885968), .Z(n_179985125));
	notech_nand3 i_1018612(.A(n_222585548), .B(n_222485547), .C(n_179985125)
		, .Z(n_18301));
	notech_nand2 i_145866837(.A(opb[7]), .B(n_264885968), .Z(n_180485130));
	notech_nand3 i_818610(.A(n_222885551), .B(n_222785550), .C(n_180485130),
		 .Z(n_18291));
	notech_nand2 i_146766828(.A(opb[5]), .B(n_264885968), .Z(n_180985135));
	notech_nand3 i_618608(.A(n_223185554), .B(n_223085553), .C(n_180985135),
		 .Z(n_18281));
	notech_and4 i_4168233(.A(n_54811), .B(n_301586335), .C(n_54775), .D(n_55018
		), .Z(n_181485140));
	notech_ao4 i_11368167(.A(n_60463), .B(n_55210), .C(n_494), .D(n_353688272
		), .Z(n_182485150));
	notech_nand2 i_188768286(.A(n_28868), .B(n_28867), .Z(n_182885154));
	notech_and2 i_188968285(.A(n_28870), .B(n_28869), .Z(n_182985155));
	notech_or4 i_10368306(.A(n_28868), .B(n_28867), .C(from_acu[3]), .D(from_acu
		[2]), .Z(n_95342672));
	notech_or4 i_11768303(.A(n_28867), .B(from_acu[1]), .C(from_acu[3]), .D(from_acu
		[2]), .Z(n_95042669));
	notech_or4 i_10068307(.A(from_acu[0]), .B(from_acu[3]), .C(n_28869), .D(n_28868
		), .Z(n_94442663));
	notech_or4 i_11968302(.A(n_28868), .B(from_acu[0]), .C(from_acu[3]), .D(from_acu
		[2]), .Z(n_94242661));
	notech_or4 i_12168300(.A(n_28869), .B(from_acu[3]), .C(from_acu[1]), .D(n_28867
		), .Z(n_93942658));
	notech_and4 i_12568296(.A(from_acu[2]), .B(from_acu[1]), .C(from_acu[0])
		, .D(n_28870), .Z(n_93742656));
	notech_ao4 i_22168070(.A(n_27375), .B(n_52390), .C(n_27752), .D(n_52380)
		, .Z(n_183585161));
	notech_ao4 i_22268069(.A(n_52410), .B(n_27823), .C(n_52400), .D(n_27688)
		, .Z(n_183785163));
	notech_ao4 i_22368068(.A(n_28024), .B(n_52431), .C(n_52421), .D(n_27720)
		, .Z(n_183885164));
	notech_and4 i_22668065(.A(n_183885164), .B(n_183785163), .C(n_183585161)
		, .D(n_128084607), .Z(n_184085166));
	notech_ao4 i_29767995(.A(n_52390), .B(n_27380), .C(n_52380), .D(n_27757)
		, .Z(n_184185167));
	notech_ao4 i_29867994(.A(n_52410), .B(n_27828), .C(n_52400), .D(n_27693)
		, .Z(n_184385169));
	notech_ao4 i_29967993(.A(n_28029), .B(n_52431), .C(n_52421), .D(n_27725)
		, .Z(n_184485170));
	notech_and4 i_30267990(.A(n_184485170), .B(n_184385169), .C(n_184185167)
		, .D(n_128884615), .Z(n_184685172));
	notech_ao4 i_34267950(.A(n_52390), .B(n_27383), .C(n_52380), .D(n_27761)
		, .Z(n_184785173));
	notech_ao4 i_34367949(.A(n_52410), .B(n_27831), .C(n_52400), .D(n_27696)
		, .Z(n_184985175));
	notech_ao4 i_34467948(.A(n_28032), .B(n_52431), .C(n_52421), .D(n_27728)
		, .Z(n_185085176));
	notech_and4 i_34767945(.A(n_185085176), .B(n_184985175), .C(n_184785173)
		, .D(n_129684623), .Z(n_185285178));
	notech_ao4 i_35767935(.A(n_52390), .B(n_27384), .C(n_52380), .D(n_27763)
		, .Z(n_185385179));
	notech_ao4 i_35867934(.A(n_52410), .B(n_27832), .C(n_52400), .D(n_27697)
		, .Z(n_185585181));
	notech_ao4 i_35967933(.A(n_28033), .B(n_52431), .C(n_52421), .D(n_27729)
		, .Z(n_185685182));
	notech_and4 i_36267930(.A(n_185685182), .B(n_185585181), .C(n_185385179)
		, .D(n_130484631), .Z(n_185885184));
	notech_ao4 i_37267920(.A(n_52389), .B(n_27385), .C(n_52379), .D(n_27764)
		, .Z(n_185985185));
	notech_ao4 i_37367919(.A(n_52409), .B(n_27833), .C(n_52399), .D(n_27698)
		, .Z(n_186185187));
	notech_ao4 i_37467918(.A(n_28034), .B(n_52430), .C(n_52419), .D(n_27730)
		, .Z(n_186285188));
	notech_and4 i_37767915(.A(n_186285188), .B(n_186185187), .C(n_185985185)
		, .D(n_131284639), .Z(n_186485190));
	notech_ao4 i_38767905(.A(n_52389), .B(n_27386), .C(n_52379), .D(n_27766)
		, .Z(n_186585191));
	notech_ao4 i_38867904(.A(n_52409), .B(n_27834), .C(n_52399), .D(n_27699)
		, .Z(n_186785193));
	notech_ao4 i_38967903(.A(n_28035), .B(n_52430), .C(n_52419), .D(n_27731)
		, .Z(n_186885194));
	notech_and4 i_39267900(.A(n_186885194), .B(n_186785193), .C(n_186585191)
		, .D(n_132084647), .Z(n_187085196));
	notech_ao4 i_40267890(.A(n_52389), .B(n_27387), .C(n_52379), .D(n_27768)
		, .Z(n_187185197));
	notech_ao4 i_40367889(.A(n_52409), .B(n_27835), .C(n_52399), .D(n_27700)
		, .Z(n_187385199));
	notech_ao4 i_40467888(.A(n_28036), .B(n_52430), .C(n_52419), .D(n_27732)
		, .Z(n_187485200));
	notech_and4 i_40767885(.A(n_187485200), .B(n_187385199), .C(n_187185197)
		, .D(n_132884655), .Z(n_187685202));
	notech_ao4 i_41767875(.A(n_52389), .B(n_27388), .C(n_52379), .D(n_27769)
		, .Z(n_187785203));
	notech_ao4 i_41867874(.A(n_52409), .B(n_27836), .C(n_52399), .D(n_27701)
		, .Z(n_187985205));
	notech_ao4 i_41967873(.A(n_28037), .B(n_52430), .C(n_52419), .D(n_27733)
		, .Z(n_188085206));
	notech_and4 i_42267870(.A(n_188085206), .B(n_187985205), .C(n_187785203)
		, .D(n_133684663), .Z(n_188285208));
	notech_ao4 i_43267860(.A(n_52392), .B(n_27389), .C(n_52381), .D(n_27770)
		, .Z(n_188385209));
	notech_ao4 i_43367859(.A(n_52412), .B(n_27837), .C(n_52401), .D(n_27702)
		, .Z(n_188585211));
	notech_ao4 i_43467858(.A(n_28038), .B(n_52433), .C(n_52422), .D(n_27734)
		, .Z(n_188685212));
	notech_and4 i_43767855(.A(n_188685212), .B(n_188585211), .C(n_188385209)
		, .D(n_134484671), .Z(n_188885214));
	notech_ao4 i_44767845(.A(n_52392), .B(n_27390), .C(n_52381), .D(n_27772)
		, .Z(n_188985215));
	notech_ao4 i_44867844(.A(n_52412), .B(n_27838), .C(n_52401), .D(n_27703)
		, .Z(n_189185217));
	notech_ao4 i_44967843(.A(n_28039), .B(n_52433), .C(n_52422), .D(n_27735)
		, .Z(n_189285218));
	notech_and4 i_45267840(.A(n_189285218), .B(n_189185217), .C(n_188985215)
		, .D(n_135284679), .Z(n_189485220));
	notech_ao4 i_46267830(.A(n_52392), .B(n_27391), .C(n_52381), .D(n_27773)
		, .Z(n_189585221));
	notech_ao4 i_46367829(.A(n_52412), .B(n_27839), .C(n_52401), .D(n_27704)
		, .Z(n_189785223));
	notech_ao4 i_46467828(.A(n_28040), .B(n_52433), .C(n_52422), .D(n_27736)
		, .Z(n_189885224));
	notech_and4 i_46767825(.A(n_189885224), .B(n_189785223), .C(n_189585221)
		, .D(n_136084687), .Z(n_190085226));
	notech_ao4 i_47767815(.A(n_52392), .B(n_27392), .C(n_52381), .D(n_27774)
		, .Z(n_190185227));
	notech_ao4 i_47867814(.A(n_52412), .B(n_27840), .C(n_52401), .D(n_27705)
		, .Z(n_190385229));
	notech_ao4 i_47967813(.A(n_28041), .B(n_52433), .C(n_52422), .D(n_27737)
		, .Z(n_190485230));
	notech_and4 i_48267810(.A(n_190485230), .B(n_190385229), .C(n_190185227)
		, .D(n_136884695), .Z(n_190685232));
	notech_ao4 i_49367800(.A(n_52391), .B(n_27393), .C(n_52380), .D(n_27777)
		, .Z(n_190785233));
	notech_ao4 i_49467799(.A(n_52411), .B(n_27841), .C(n_52400), .D(n_27706)
		, .Z(n_190985235));
	notech_ao4 i_49567798(.A(n_28042), .B(n_52432), .C(n_52421), .D(n_27738)
		, .Z(n_191085236));
	notech_and4 i_49867795(.A(n_191085236), .B(n_190985235), .C(n_190785233)
		, .D(n_137684703), .Z(n_191285238));
	notech_ao4 i_50867785(.A(n_52391), .B(n_27394), .C(n_52380), .D(n_27778)
		, .Z(n_191385239));
	notech_ao4 i_50967784(.A(n_52411), .B(n_27842), .C(n_52400), .D(n_27707)
		, .Z(n_191585241));
	notech_ao4 i_51067783(.A(n_28043), .B(n_52432), .C(n_52421), .D(n_27739)
		, .Z(n_191685242));
	notech_and4 i_51367780(.A(n_191685242), .B(n_191585241), .C(n_191385239)
		, .D(n_138484711), .Z(n_191885244));
	notech_ao4 i_52367770(.A(n_52391), .B(n_27395), .C(n_52381), .D(n_27779)
		, .Z(n_191985245));
	notech_ao4 i_52467769(.A(n_52411), .B(n_27843), .C(n_52401), .D(n_27708)
		, .Z(n_192185247));
	notech_ao4 i_52567768(.A(n_28044), .B(n_52432), .C(n_52422), .D(n_27740)
		, .Z(n_192285248));
	notech_and4 i_52867765(.A(n_192285248), .B(n_192185247), .C(n_191985245)
		, .D(n_139284719), .Z(n_192485250));
	notech_ao4 i_53867755(.A(n_52391), .B(n_27396), .C(n_52381), .D(n_27780)
		, .Z(n_192585251));
	notech_ao4 i_53967754(.A(n_52411), .B(n_27844), .C(n_52401), .D(n_27709)
		, .Z(n_192785253));
	notech_ao4 i_54067753(.A(n_28045), .B(n_52432), .C(n_52422), .D(n_27741)
		, .Z(n_192885254));
	notech_and4 i_54367750(.A(n_192885254), .B(n_192785253), .C(n_192585251)
		, .D(n_140084727), .Z(n_193085256));
	notech_ao4 i_55367740(.A(n_52385), .B(n_27397), .C(n_52376), .D(n_27781)
		, .Z(n_193185257));
	notech_ao4 i_55467739(.A(n_52405), .B(n_27845), .C(n_52396), .D(n_27710)
		, .Z(n_193385259));
	notech_ao4 i_55567738(.A(n_28046), .B(n_52426), .C(n_52416), .D(n_27742)
		, .Z(n_193485260));
	notech_and4 i_55867735(.A(n_193485260), .B(n_193385259), .C(n_193185257)
		, .D(n_140884735), .Z(n_193685262));
	notech_ao4 i_56867725(.A(n_52385), .B(n_27398), .C(n_52375), .D(n_27782)
		, .Z(n_193785263));
	notech_ao4 i_56967724(.A(n_52405), .B(n_27846), .C(n_52395), .D(n_27711)
		, .Z(n_193985265));
	notech_ao4 i_57067723(.A(n_28047), .B(n_52426), .C(n_52415), .D(n_27743)
		, .Z(n_194085266));
	notech_and4 i_57367720(.A(n_194085266), .B(n_193985265), .C(n_193785263)
		, .D(n_141684743), .Z(n_194285268));
	notech_ao4 i_58367710(.A(n_52385), .B(n_27399), .C(n_52376), .D(n_27783)
		, .Z(n_194385269));
	notech_ao4 i_58467709(.A(n_52405), .B(n_27847), .C(n_52396), .D(n_27712)
		, .Z(n_194585271));
	notech_ao4 i_58567708(.A(n_28048), .B(n_52426), .C(n_52416), .D(n_27744)
		, .Z(n_194685272));
	notech_and4 i_58867705(.A(n_194685272), .B(n_194585271), .C(n_194385269)
		, .D(n_142484751), .Z(n_194885274));
	notech_ao4 i_61367680(.A(n_52385), .B(n_27401), .C(n_52376), .D(n_27785)
		, .Z(n_194985275));
	notech_ao4 i_61467679(.A(n_52405), .B(n_27849), .C(n_52396), .D(n_27714)
		, .Z(n_195185277));
	notech_ao4 i_61567678(.A(n_28050), .B(n_52426), .C(n_52416), .D(n_27746)
		, .Z(n_195285278));
	notech_and4 i_61867675(.A(n_195285278), .B(n_195185277), .C(n_194985275)
		, .D(n_143284759), .Z(n_195485280));
	notech_nand2 i_189168283(.A(n_28872), .B(n_28871), .Z(n_195585281));
	notech_nor2 i_189268282(.A(from_acu[7]), .B(from_acu[6]), .Z(n_195685282
		));
	notech_or4 i_12268299(.A(from_acu[7]), .B(n_28871), .C(from_acu[5]), .D(from_acu
		[6]), .Z(n_196185287));
	notech_or4 i_12368298(.A(from_acu[7]), .B(from_acu[6]), .C(n_28872), .D(from_acu
		[4]), .Z(n_196385289));
	notech_ao4 i_62967664(.A(n_52473), .B(n_27818), .C(n_52463), .D(n_27370)
		, .Z(n_196485290));
	notech_or4 i_9568309(.A(from_acu[7]), .B(n_28873), .C(from_acu[4]), .D(n_28872
		), .Z(n_196785293));
	notech_or4 i_12468297(.A(from_acu[7]), .B(n_28872), .C(n_28871), .D(from_acu
		[6]), .Z(n_196985295));
	notech_ao4 i_63067663(.A(n_52493), .B(n_27747), .C(n_52483), .D(n_27681)
		, .Z(n_197085296));
	notech_or4 i_9768308(.A(from_acu[7]), .B(n_28873), .C(n_28872), .D(n_28871
		), .Z(n_197185297));
	notech_or4 i_14168294(.A(from_acu[7]), .B(from_acu[5]), .C(n_28873), .D(n_28871
		), .Z(n_197285298));
	notech_ao4 i_63167662(.A(n_52513), .B(n_27715), .C(n_28019), .D(n_52503)
		, .Z(n_197385299));
	notech_and4 i_63467659(.A(n_197385299), .B(n_197085296), .C(n_196485290)
		, .D(n_144084767), .Z(n_197585301));
	notech_ao4 i_64467649(.A(n_52473), .B(n_27819), .C(n_52463), .D(n_27371)
		, .Z(n_197685302));
	notech_ao4 i_64567648(.A(n_52493), .B(n_27748), .C(n_52483), .D(n_27682)
		, .Z(n_197885304));
	notech_ao4 i_64667647(.A(n_52513), .B(n_27716), .C(n_28020), .D(n_52503)
		, .Z(n_197985305));
	notech_and4 i_64967644(.A(n_197985305), .B(n_197885304), .C(n_197685302)
		, .D(n_144884775), .Z(n_198185307));
	notech_ao4 i_65967634(.A(n_52473), .B(n_27820), .C(n_52463), .D(n_27372)
		, .Z(n_198285308));
	notech_ao4 i_66067633(.A(n_52493), .B(n_27749), .C(n_52483), .D(n_27685)
		, .Z(n_198485310));
	notech_ao4 i_66167632(.A(n_52513), .B(n_27717), .C(n_28021), .D(n_52503)
		, .Z(n_198585311));
	notech_and4 i_66467629(.A(n_198585311), .B(n_198485310), .C(n_198285308)
		, .D(n_145684783), .Z(n_198785313));
	notech_ao4 i_67467619(.A(n_52473), .B(n_27821), .C(n_52463), .D(n_27373)
		, .Z(n_198885314));
	notech_ao4 i_67567618(.A(n_52493), .B(n_27750), .C(n_52483), .D(n_27686)
		, .Z(n_199085316));
	notech_ao4 i_67667617(.A(n_52513), .B(n_27718), .C(n_52503), .D(n_28022)
		, .Z(n_199185317));
	notech_and4 i_67967614(.A(n_199185317), .B(n_199085316), .C(n_198885314)
		, .D(n_146484791), .Z(n_199385319));
	notech_ao4 i_68967604(.A(n_52472), .B(n_27822), .C(n_52462), .D(n_27374)
		, .Z(n_199485320));
	notech_ao4 i_69067603(.A(n_52492), .B(n_27751), .C(n_52482), .D(n_27687)
		, .Z(n_199685322));
	notech_ao4 i_69167602(.A(n_52512), .B(n_27719), .C(n_28023), .D(n_52502)
		, .Z(n_199785323));
	notech_and4 i_69467599(.A(n_199785323), .B(n_199685322), .C(n_199485320)
		, .D(n_147284799), .Z(n_199985325));
	notech_ao4 i_70467589(.A(n_52472), .B(n_27823), .C(n_52462), .D(n_27375)
		, .Z(n_200085326));
	notech_ao4 i_70567588(.A(n_52492), .B(n_27752), .C(n_52482), .D(n_27688)
		, .Z(n_200285328));
	notech_ao4 i_70667587(.A(n_52512), .B(n_27720), .C(n_52502), .D(n_28024)
		, .Z(n_200385329));
	notech_and4 i_70967584(.A(n_200385329), .B(n_200285328), .C(n_200085326)
		, .D(n_148084807), .Z(n_200585331));
	notech_ao4 i_71967574(.A(n_52472), .B(n_27824), .C(n_52462), .D(n_27376)
		, .Z(n_200685332));
	notech_ao4 i_72067573(.A(n_52492), .B(n_27753), .C(n_52482), .D(n_27689)
		, .Z(n_200885334));
	notech_ao4 i_72167572(.A(n_52512), .B(n_27721), .C(n_28025), .D(n_52502)
		, .Z(n_200985335));
	notech_and4 i_72467569(.A(n_200985335), .B(n_200885334), .C(n_200685332)
		, .D(n_148884815), .Z(n_201185337));
	notech_ao4 i_73467559(.A(n_52472), .B(n_27825), .C(n_52462), .D(n_27377)
		, .Z(n_201285338));
	notech_ao4 i_73567558(.A(n_52492), .B(n_27754), .C(n_52482), .D(n_27690)
		, .Z(n_201485340));
	notech_ao4 i_73667557(.A(n_52512), .B(n_27722), .C(n_28026), .D(n_52502)
		, .Z(n_201585341));
	notech_and4 i_73967554(.A(n_201585341), .B(n_201485340), .C(n_201285338)
		, .D(n_149684823), .Z(n_201785343));
	notech_ao4 i_74967544(.A(n_52475), .B(n_27826), .C(n_52464), .D(n_27378)
		, .Z(n_201885344));
	notech_ao4 i_75067543(.A(n_52495), .B(n_27755), .C(n_52484), .D(n_27691)
		, .Z(n_202085346));
	notech_ao4 i_75167542(.A(n_27723), .B(n_52515), .C(n_28027), .D(n_52504)
		, .Z(n_202185347));
	notech_and4 i_75467539(.A(n_202185347), .B(n_202085346), .C(n_201885344)
		, .D(n_150484831), .Z(n_202385349));
	notech_ao4 i_76467529(.A(n_52475), .B(n_27827), .C(n_52464), .D(n_27379)
		, .Z(n_202485350));
	notech_ao4 i_76567528(.A(n_52495), .B(n_27756), .C(n_52484), .D(n_27692)
		, .Z(n_202685352));
	notech_ao4 i_76667527(.A(n_52515), .B(n_27724), .C(n_28028), .D(n_52504)
		, .Z(n_202785353));
	notech_and4 i_76967524(.A(n_202785353), .B(n_202685352), .C(n_202485350)
		, .D(n_151284839), .Z(n_202985355));
	notech_ao4 i_77967514(.A(n_52475), .B(n_27828), .C(n_52464), .D(n_27380)
		, .Z(n_203085356));
	notech_ao4 i_78067513(.A(n_52495), .B(n_27757), .C(n_52484), .D(n_27693)
		, .Z(n_203285358));
	notech_ao4 i_78167512(.A(n_52515), .B(n_27725), .C(n_28029), .D(n_52504)
		, .Z(n_203385359));
	notech_and4 i_78467509(.A(n_203385359), .B(n_203285358), .C(n_203085356)
		, .D(n_152084847), .Z(n_203585361));
	notech_ao4 i_79467499(.A(n_52475), .B(n_27829), .C(n_52464), .D(n_27381)
		, .Z(n_203685362));
	notech_ao4 i_79567498(.A(n_52495), .B(n_27758), .C(n_52484), .D(n_27694)
		, .Z(n_203885364));
	notech_ao4 i_79667497(.A(n_52515), .B(n_27726), .C(n_28030), .D(n_52504)
		, .Z(n_203985365));
	notech_and4 i_79967494(.A(n_203985365), .B(n_203885364), .C(n_203685362)
		, .D(n_152884855), .Z(n_204185367));
	notech_ao4 i_80967484(.A(n_52474), .B(n_27830), .C(n_52463), .D(n_27382)
		, .Z(n_204285368));
	notech_ao4 i_81067483(.A(n_52494), .B(n_27760), .C(n_52483), .D(n_27695)
		, .Z(n_204485370));
	notech_ao4 i_81167482(.A(n_52514), .B(n_27727), .C(n_52503), .D(n_28031)
		, .Z(n_204585371));
	notech_and4 i_81467479(.A(n_204585371), .B(n_204485370), .C(n_204285368)
		, .D(n_153684863), .Z(n_204785373));
	notech_ao4 i_82467469(.A(n_52474), .B(n_27831), .C(n_52463), .D(n_27383)
		, .Z(n_204885374));
	notech_ao4 i_82567468(.A(n_52494), .B(n_27761), .C(n_52483), .D(n_27696)
		, .Z(n_205085376));
	notech_ao4 i_82667467(.A(n_52514), .B(n_27728), .C(n_28032), .D(n_52503)
		, .Z(n_205185377));
	notech_and4 i_82967464(.A(n_205185377), .B(n_205085376), .C(n_204885374)
		, .D(n_154484871), .Z(n_205385379));
	notech_ao4 i_83967454(.A(n_52474), .B(n_27832), .C(n_52464), .D(n_27384)
		, .Z(n_205485380));
	notech_ao4 i_84067453(.A(n_52494), .B(n_27763), .C(n_52484), .D(n_27697)
		, .Z(n_205685382));
	notech_ao4 i_84167452(.A(n_52514), .B(n_27729), .C(n_28033), .D(n_52504)
		, .Z(n_205785383));
	notech_and4 i_84467449(.A(n_205785383), .B(n_205685382), .C(n_205485380)
		, .D(n_155284879), .Z(n_205985385));
	notech_ao4 i_85467439(.A(n_52474), .B(n_27833), .C(n_52464), .D(n_27385)
		, .Z(n_206085386));
	notech_ao4 i_85567438(.A(n_52494), .B(n_27764), .C(n_52484), .D(n_27698)
		, .Z(n_206285388));
	notech_ao4 i_85667437(.A(n_52514), .B(n_27730), .C(n_28034), .D(n_52504)
		, .Z(n_206385389));
	notech_and4 i_85967434(.A(n_206385389), .B(n_206285388), .C(n_206085386)
		, .D(n_156084887), .Z(n_206585391));
	notech_ao4 i_86967424(.A(n_52468), .B(n_27834), .C(n_52459), .D(n_27386)
		, .Z(n_206685392));
	notech_ao4 i_87067423(.A(n_52488), .B(n_27766), .C(n_52479), .D(n_27699)
		, .Z(n_206885394));
	notech_ao4 i_87167422(.A(n_52508), .B(n_27731), .C(n_52499), .D(n_28035)
		, .Z(n_206985395));
	notech_and4 i_87467419(.A(n_206985395), .B(n_206885394), .C(n_206685392)
		, .D(n_156884895), .Z(n_207185397));
	notech_ao4 i_88467409(.A(n_52468), .B(n_27835), .C(n_52458), .D(n_27387)
		, .Z(n_207285398));
	notech_ao4 i_88567408(.A(n_52488), .B(n_27768), .C(n_52478), .D(n_27700)
		, .Z(n_207485400));
	notech_ao4 i_88667407(.A(n_52508), .B(n_27732), .C(n_28036), .D(n_52498)
		, .Z(n_207585401));
	notech_and4 i_88967404(.A(n_207585401), .B(n_207485400), .C(n_207285398)
		, .D(n_157684903), .Z(n_207785403));
	notech_ao4 i_89967394(.A(n_52468), .B(n_27836), .C(n_52459), .D(n_27388)
		, .Z(n_207885404));
	notech_ao4 i_90067393(.A(n_52488), .B(n_27769), .C(n_52479), .D(n_27701)
		, .Z(n_208085406));
	notech_ao4 i_90167392(.A(n_52508), .B(n_27733), .C(n_28037), .D(n_52499)
		, .Z(n_208185407));
	notech_and4 i_90467389(.A(n_208185407), .B(n_208085406), .C(n_207885404)
		, .D(n_158484911), .Z(n_208385409));
	notech_ao4 i_91467379(.A(n_52468), .B(n_27837), .C(n_52459), .D(n_27389)
		, .Z(n_208485410));
	notech_ao4 i_91567378(.A(n_52488), .B(n_27770), .C(n_52479), .D(n_27702)
		, .Z(n_208685412));
	notech_ao4 i_91667377(.A(n_52508), .B(n_27734), .C(n_28038), .D(n_52499)
		, .Z(n_208785413));
	notech_and4 i_91967374(.A(n_208785413), .B(n_208685412), .C(n_208485410)
		, .D(n_159284919), .Z(n_208985415));
	notech_ao4 i_92967364(.A(n_52467), .B(n_27838), .C(n_52458), .D(n_27390)
		, .Z(n_209085416));
	notech_ao4 i_93067363(.A(n_52487), .B(n_27772), .C(n_52478), .D(n_27703)
		, .Z(n_209285418));
	notech_ao4 i_93167362(.A(n_52507), .B(n_27735), .C(n_28039), .D(n_52498)
		, .Z(n_209385419));
	notech_and4 i_93467359(.A(n_209385419), .B(n_209285418), .C(n_209085416)
		, .D(n_160084927), .Z(n_209585421));
	notech_ao4 i_94467349(.A(n_52467), .B(n_27839), .C(n_52458), .D(n_27391)
		, .Z(n_209685422));
	notech_ao4 i_94567348(.A(n_52487), .B(n_27773), .C(n_52478), .D(n_27704)
		, .Z(n_209885424));
	notech_ao4 i_94667347(.A(n_52507), .B(n_27736), .C(n_28040), .D(n_52498)
		, .Z(n_209985425));
	notech_and4 i_94967344(.A(n_209985425), .B(n_209885424), .C(n_209685422)
		, .D(n_160884935), .Z(n_210185427));
	notech_ao4 i_95967334(.A(n_52467), .B(n_27840), .C(n_52458), .D(n_27392)
		, .Z(n_210285428));
	notech_ao4 i_96067333(.A(n_52487), .B(n_27774), .C(n_52478), .D(n_27705)
		, .Z(n_210485430));
	notech_ao4 i_96167332(.A(n_52507), .B(n_27737), .C(n_52498), .D(n_28041)
		, .Z(n_210585431));
	notech_and4 i_96467329(.A(n_210585431), .B(n_210485430), .C(n_210285428)
		, .D(n_161684943), .Z(n_210785433));
	notech_ao4 i_97467319(.A(n_52467), .B(n_27841), .C(n_52458), .D(n_27393)
		, .Z(n_210885434));
	notech_ao4 i_97567318(.A(n_52487), .B(n_27777), .C(n_52478), .D(n_27706)
		, .Z(n_211085436));
	notech_ao4 i_97667317(.A(n_52507), .B(n_27738), .C(n_28042), .D(n_52498)
		, .Z(n_211185437));
	notech_and4 i_97967314(.A(n_211185437), .B(n_211085436), .C(n_210885434)
		, .D(n_162484951), .Z(n_211385439));
	notech_ao4 i_98967304(.A(n_52470), .B(n_27842), .C(n_52460), .D(n_27394)
		, .Z(n_211485440));
	notech_ao4 i_99067303(.A(n_52490), .B(n_27778), .C(n_52480), .D(n_27707)
		, .Z(n_211685442));
	notech_ao4 i_99167302(.A(n_52510), .B(n_27739), .C(n_28043), .D(n_52500)
		, .Z(n_211785443));
	notech_and4 i_99467299(.A(n_211785443), .B(n_211685442), .C(n_211485440)
		, .D(n_163284959), .Z(n_211985445));
	notech_ao4 i_100467289(.A(n_52470), .B(n_27843), .C(n_52460), .D(n_27395
		), .Z(n_212085446));
	notech_ao4 i_100567288(.A(n_52490), .B(n_27779), .C(n_52480), .D(n_27708
		), .Z(n_212285448));
	notech_ao4 i_100667287(.A(n_52510), .B(n_27740), .C(n_28044), .D(n_52500
		), .Z(n_212385449));
	notech_and4 i_100967284(.A(n_212385449), .B(n_212285448), .C(n_212085446
		), .D(n_164084967), .Z(n_212585451));
	notech_ao4 i_101967274(.A(n_52470), .B(n_27844), .C(n_52462), .D(n_27396
		), .Z(n_212685452));
	notech_ao4 i_102067273(.A(n_52490), .B(n_27780), .C(n_52482), .D(n_27709
		), .Z(n_212885454));
	notech_ao4 i_102167272(.A(n_52510), .B(n_27741), .C(n_28045), .D(n_52502
		), .Z(n_212985455));
	notech_and4 i_102467269(.A(n_212985455), .B(n_212885454), .C(n_212685452
		), .D(n_164884975), .Z(n_213185457));
	notech_ao4 i_103567259(.A(n_52470), .B(n_27845), .C(n_52460), .D(n_27397
		), .Z(n_213285458));
	notech_ao4 i_103667258(.A(n_52490), .B(n_27781), .C(n_52480), .D(n_27710
		), .Z(n_213485460));
	notech_ao4 i_103767257(.A(n_52510), .B(n_27742), .C(n_28046), .D(n_52500
		), .Z(n_213585461));
	notech_and4 i_104067254(.A(n_213585461), .B(n_213485460), .C(n_213285458
		), .D(n_165684983), .Z(n_213785463));
	notech_ao4 i_105067244(.A(n_52469), .B(n_27846), .C(n_52459), .D(n_27398
		), .Z(n_213885464));
	notech_ao4 i_105167243(.A(n_52489), .B(n_27782), .C(n_52479), .D(n_27711
		), .Z(n_214085466));
	notech_ao4 i_105267242(.A(n_52509), .B(n_27743), .C(n_28047), .D(n_52499
		), .Z(n_214185467));
	notech_and4 i_105567239(.A(n_214185467), .B(n_214085466), .C(n_213885464
		), .D(n_166484991), .Z(n_214385469));
	notech_ao4 i_106567229(.A(n_52469), .B(n_27847), .C(n_52459), .D(n_27399
		), .Z(n_214485470));
	notech_ao4 i_106667228(.A(n_52489), .B(n_27783), .C(n_52479), .D(n_27712
		), .Z(n_214685472));
	notech_ao4 i_106767227(.A(n_52509), .B(n_27744), .C(n_28048), .D(n_52499
		), .Z(n_214785473));
	notech_and4 i_107067224(.A(n_214785473), .B(n_214685472), .C(n_214485470
		), .D(n_167284999), .Z(n_214985475));
	notech_ao4 i_108067214(.A(n_52469), .B(n_27848), .C(n_52460), .D(n_27400
		), .Z(n_215085476));
	notech_ao4 i_108167213(.A(n_52489), .B(n_27784), .C(n_52480), .D(n_27713
		), .Z(n_215285478));
	notech_ao4 i_108267212(.A(n_52509), .B(n_27745), .C(n_52500), .D(n_28049
		), .Z(n_215385479));
	notech_and4 i_108567209(.A(n_215385479), .B(n_215285478), .C(n_215085476
		), .D(n_168085007), .Z(n_215585481));
	notech_ao4 i_109567199(.A(n_52469), .B(n_27849), .C(n_52460), .D(n_27401
		), .Z(n_215685482));
	notech_ao4 i_109667198(.A(n_52489), .B(n_27785), .C(n_52480), .D(n_27714
		), .Z(n_215885484));
	notech_ao4 i_109767197(.A(n_52509), .B(n_27746), .C(n_52500), .D(n_28050
		), .Z(n_215985485));
	notech_and4 i_110067194(.A(n_215985485), .B(n_215885484), .C(n_215685482
		), .D(n_168885015), .Z(n_216185487));
	notech_ao4 i_111067184(.A(n_28442003), .B(n_27297), .C(n_56409), .D(n_26923
		), .Z(n_216285488));
	notech_ao4 i_111167183(.A(n_27341992), .B(n_27333), .C(n_26595), .D(n_2699
		), .Z(n_216385489));
	notech_ao4 i_112467170(.A(n_28442003), .B(n_27300), .C(n_56409), .D(n_26927
		), .Z(n_216485490));
	notech_ao4 i_112567169(.A(n_27341992), .B(n_27335), .C(n_26595), .D(n_322488466
		), .Z(n_216585491));
	notech_ao4 i_113167163(.A(n_28442003), .B(n_27301), .C(n_56409), .D(n_26929
		), .Z(n_216685492));
	notech_ao4 i_113267162(.A(n_27341992), .B(n_27336), .C(n_26595), .D(n_322688464
		), .Z(n_216785493));
	notech_ao4 i_113867156(.A(n_28442003), .B(n_27302), .C(n_56404), .D(n_26931
		), .Z(n_216885494));
	notech_ao4 i_113967155(.A(n_27341992), .B(n_27337), .C(n_26595), .D(n_321188478
		), .Z(n_216985495));
	notech_ao4 i_114567149(.A(n_28442003), .B(n_27304), .C(n_56404), .D(n_26933
		), .Z(n_217085496));
	notech_ao4 i_114667148(.A(n_27341992), .B(n_27338), .C(n_26595), .D(n_322788463
		), .Z(n_217185497));
	notech_ao4 i_115967135(.A(n_28442003), .B(n_27308), .C(n_56404), .D(n_26937
		), .Z(n_217285498));
	notech_ao4 i_116067134(.A(n_27341992), .B(n_27340), .C(n_26595), .D(n_57351
		), .Z(n_217385499));
	notech_ao4 i_120867086(.A(n_53296), .B(n_27318), .C(n_26957), .D(n_56404
		), .Z(n_217485500));
	notech_ao4 i_120967085(.A(n_53285), .B(n_27351), .C(n_53276), .D(n_2700)
		, .Z(n_217585501));
	notech_ao4 i_121567079(.A(n_53296), .B(n_27325), .C(n_56404), .D(n_26971
		), .Z(n_217685502));
	notech_ao4 i_121667078(.A(n_53285), .B(n_27358), .C(n_53276), .D(n_57334
		), .Z(n_217785503));
	notech_ao4 i_122267072(.A(n_53296), .B(n_27330), .C(n_56404), .D(n_26983
		), .Z(n_217885504));
	notech_ao4 i_122367071(.A(n_53285), .B(n_27363), .C(n_53276), .D(n_57329
		), .Z(n_217985505));
	notech_or4 i_164368289(.A(n_274588712), .B(n_60586), .C(n_59890), .D(n_106813462
		), .Z(n_218285508));
	notech_ao4 i_123767057(.A(n_26599), .B(n_56766), .C(n_57438), .D(n_58951
		), .Z(n_218485510));
	notech_ao4 i_124267052(.A(n_57438), .B(n_55252), .C(n_55253), .D(n_26599
		), .Z(n_218585511));
	notech_or4 i_124767047(.A(n_275488703), .B(n_59967), .C(n_59210), .D(n_54913
		), .Z(n_218685512));
	notech_ao4 i_48968292(.A(n_218685512), .B(n_59889), .C(n_48510), .D(n_2826
		), .Z(n_218785513));
	notech_ao4 i_135166943(.A(n_54762), .B(n_27391), .C(n_59817), .D(n_28898
		), .Z(n_218885514));
	notech_ao4 i_135066944(.A(n_55943), .B(n_58996), .C(n_54642), .D(n_27773
		), .Z(n_218985515));
	notech_ao4 i_136066934(.A(n_54762), .B(n_27390), .C(n_59817), .D(n_28897
		), .Z(n_219185517));
	notech_ao4 i_135966935(.A(n_55943), .B(n_59005), .C(n_54642), .D(n_27772
		), .Z(n_219285518));
	notech_ao4 i_136966925(.A(n_54762), .B(n_27389), .C(n_59817), .D(n_28894
		), .Z(n_219485520));
	notech_ao4 i_136866926(.A(n_55943), .B(n_59014), .C(n_54642), .D(n_27770
		), .Z(n_219585521));
	notech_ao4 i_137866916(.A(n_54762), .B(n_27388), .C(n_59817), .D(n_28893
		), .Z(n_219885523));
	notech_ao4 i_137766917(.A(n_55943), .B(n_58969), .C(n_54642), .D(n_27769
		), .Z(n_219985524));
	notech_ao4 i_138766907(.A(n_54762), .B(n_27387), .C(n_59817), .D(n_28892
		), .Z(n_220185526));
	notech_ao4 i_138666908(.A(n_55943), .B(n_58978), .C(n_54642), .D(n_27768
		), .Z(n_220285527));
	notech_ao4 i_139666898(.A(n_54762), .B(n_27386), .C(n_59817), .D(n_28891
		), .Z(n_220585529));
	notech_ao4 i_139566899(.A(n_55943), .B(n_58987), .C(n_54642), .D(n_27766
		), .Z(n_220685530));
	notech_ao4 i_140566889(.A(n_54762), .B(n_27384), .C(n_59817), .D(n_28889
		), .Z(n_220885532));
	notech_ao4 i_140466890(.A(n_55943), .B(nbus_11326[14]), .C(n_54642), .D(n_27763
		), .Z(n_221085533));
	notech_ao4 i_141466880(.A(n_54762), .B(n_27383), .C(n_59828), .D(n_28888
		), .Z(n_221285535));
	notech_ao4 i_141366881(.A(n_55943), .B(nbus_11326[13]), .C(n_54642), .D(n_27761
		), .Z(n_221385536));
	notech_ao4 i_142466871(.A(n_54762), .B(n_27382), .C(n_59828), .D(n_28887
		), .Z(n_221585538));
	notech_ao4 i_142366872(.A(n_55943), .B(nbus_11326[12]), .C(n_54642), .D(n_27760
		), .Z(n_221685539));
	notech_ao4 i_143366862(.A(n_54762), .B(n_27381), .C(n_59828), .D(n_28886
		), .Z(n_221885541));
	notech_ao4 i_143266863(.A(n_55943), .B(nbus_11326[11]), .C(n_54642), .D(n_27758
		), .Z(n_221985542));
	notech_ao4 i_144266853(.A(n_54762), .B(n_27380), .C(n_59828), .D(n_28885
		), .Z(n_222185544));
	notech_ao4 i_144166854(.A(n_55943), .B(nbus_11326[10]), .C(n_54642), .D(n_27757
		), .Z(n_222285545));
	notech_ao4 i_145166844(.A(n_54762), .B(n_27379), .C(n_59828), .D(n_28884
		), .Z(n_222485547));
	notech_ao4 i_145066845(.A(n_55943), .B(nbus_11326[9]), .C(n_54642), .D(n_27756
		), .Z(n_222585548));
	notech_ao4 i_146066835(.A(n_54762), .B(n_27377), .C(n_59826), .D(n_28882
		), .Z(n_222785550));
	notech_ao4 i_145966836(.A(n_55943), .B(nbus_11326[7]), .C(n_54642), .D(n_27754
		), .Z(n_222885551));
	notech_ao4 i_146966826(.A(n_54762), .B(n_27375), .C(n_59826), .D(n_28880
		), .Z(n_223085553));
	notech_ao4 i_146866827(.A(n_55943), .B(nbus_11326[5]), .C(n_27752), .D(n_54642
		), .Z(n_223185554));
	notech_nand2 i_7365685(.A(n_265185971), .B(n_59826), .Z(n_223485557));
	notech_xor2 i_3065638(.A(pipe_mul[1]), .B(pipe_mul[0]), .Z(n_223585558)
		);
	notech_and4 i_47265684(.A(n_61624), .B(n_55943), .C(n_238985709), .D(n_26610
		), .Z(n_223785560));
	notech_ao4 i_2465644(.A(n_260688757), .B(n_2605), .C(n_57448), .D(n_56067
		), .Z(n_223985562));
	notech_or2 i_13265538(.A(n_55115), .B(n_57417), .Z(n_224085563));
	notech_nand2 i_44465253(.A(divr_0[0]), .B(n_59889), .Z(n_224285565));
	notech_nand2 i_44765250(.A(divr_0[1]), .B(n_59880), .Z(n_224385566));
	notech_nand2 i_45065247(.A(divr_0[2]), .B(n_59880), .Z(n_224485567));
	notech_nand2 i_45365244(.A(divr_0[3]), .B(n_59876), .Z(n_224585568));
	notech_nand2 i_45665241(.A(divr_0[4]), .B(n_59876), .Z(n_224685569));
	notech_nand2 i_45965238(.A(divr_0[5]), .B(n_59876), .Z(n_224785570));
	notech_nand2 i_46265235(.A(divr_0[6]), .B(n_59880), .Z(n_224885571));
	notech_nand2 i_46565232(.A(divr_0[7]), .B(n_59880), .Z(n_224985572));
	notech_nand2 i_46865229(.A(divr_0[8]), .B(n_59880), .Z(n_225085573));
	notech_nand2 i_47165226(.A(divr_0[9]), .B(n_59880), .Z(n_225185574));
	notech_nand2 i_47565223(.A(divr_0[10]), .B(n_59880), .Z(n_225285575));
	notech_nand2 i_47865220(.A(divr_0[11]), .B(n_59876), .Z(n_225385576));
	notech_nand2 i_48165217(.A(divr_0[12]), .B(n_59876), .Z(n_225485577));
	notech_nand2 i_48465214(.A(divr_0[13]), .B(n_59876), .Z(n_225585578));
	notech_nand2 i_48765211(.A(divr_0[14]), .B(n_59876), .Z(n_225685579));
	notech_nand2 i_49065208(.A(divr_0[15]), .B(n_59876), .Z(n_225785580));
	notech_nand2 i_49365205(.A(divr_0[16]), .B(n_59876), .Z(n_225885581));
	notech_nand2 i_49665202(.A(divr_0[17]), .B(n_59876), .Z(n_225985582));
	notech_nand2 i_49965199(.A(divr_0[18]), .B(n_59876), .Z(n_226185583));
	notech_nand2 i_50265196(.A(divr_0[19]), .B(n_59876), .Z(n_226285584));
	notech_nand2 i_50565193(.A(divr_0[20]), .B(n_59876), .Z(n_226385585));
	notech_nand2 i_50865190(.A(divr_0[21]), .B(n_59876), .Z(n_226485586));
	notech_nand2 i_51165187(.A(divr_0[22]), .B(n_59881), .Z(n_226585587));
	notech_nand2 i_51465184(.A(divr_0[23]), .B(n_59881), .Z(n_226685588));
	notech_nand2 i_51765181(.A(divr_0[24]), .B(n_59881), .Z(n_226785589));
	notech_nand2 i_52065178(.A(divr_0[25]), .B(n_59881), .Z(n_226885590));
	notech_nand2 i_52365175(.A(divr_0[26]), .B(n_59881), .Z(n_226985591));
	notech_nand2 i_52665172(.A(divr_0[27]), .B(n_59881), .Z(n_227085592));
	notech_nand2 i_52965169(.A(divr_0[28]), .B(n_59881), .Z(n_227185593));
	notech_nand2 i_53265166(.A(divr_0[29]), .B(n_59881), .Z(n_227285594));
	notech_nand2 i_53565163(.A(divr_0[30]), .B(n_59881), .Z(n_227385595));
	notech_nand2 i_53865160(.A(divr_0[31]), .B(n_59881), .Z(n_227485596));
	notech_nand2 i_54165157(.A(divr_0[32]), .B(n_59881), .Z(n_227585597));
	notech_nand2 i_54465154(.A(divr_0[33]), .B(n_59880), .Z(n_227685598));
	notech_nand2 i_54765151(.A(divr_0[34]), .B(n_59880), .Z(n_227785599));
	notech_nand2 i_55065148(.A(divr_0[35]), .B(n_59880), .Z(n_227885600));
	notech_nand2 i_55365145(.A(divr_0[36]), .B(n_59880), .Z(n_227985601));
	notech_nand2 i_55665142(.A(divr_0[37]), .B(n_59880), .Z(n_228085602));
	notech_nand2 i_55965139(.A(divr_0[38]), .B(n_59881), .Z(n_228185603));
	notech_nand2 i_56265136(.A(divr_0[39]), .B(n_59881), .Z(n_228285604));
	notech_nand2 i_56565133(.A(divr_0[40]), .B(n_59881), .Z(n_228385605));
	notech_nand2 i_56865130(.A(divr_0[41]), .B(n_59880), .Z(n_228485606));
	notech_nand2 i_57165127(.A(divr_0[42]), .B(n_59880), .Z(n_228585607));
	notech_nand2 i_57465124(.A(divr_0[43]), .B(n_59907), .Z(n_228685608));
	notech_nand2 i_57765121(.A(divr_0[44]), .B(n_59907), .Z(n_228785609));
	notech_nand2 i_58065118(.A(divr_0[45]), .B(n_59903), .Z(n_228885610));
	notech_nand2 i_58365115(.A(divr_0[46]), .B(n_59903), .Z(n_228985611));
	notech_nand2 i_58665112(.A(divr_0[47]), .B(n_59903), .Z(n_229085612));
	notech_nand2 i_58965109(.A(divr_0[48]), .B(n_59907), .Z(n_229185613));
	notech_nand2 i_59265106(.A(divr_0[49]), .B(n_59907), .Z(n_229285614));
	notech_nand2 i_59565103(.A(divr_0[50]), .B(n_59907), .Z(n_229385615));
	notech_nand2 i_59865100(.A(divr_0[51]), .B(n_59907), .Z(n_229485616));
	notech_nand2 i_60165097(.A(divr_0[52]), .B(n_59907), .Z(n_229585617));
	notech_nand2 i_60465094(.A(divr_0[53]), .B(n_59903), .Z(n_229685618));
	notech_nand2 i_60765091(.A(divr_0[54]), .B(n_59903), .Z(n_229785619));
	notech_nand2 i_61065088(.A(divr_0[55]), .B(n_59903), .Z(n_229885620));
	notech_nand2 i_61365085(.A(divr_0[56]), .B(n_59903), .Z(n_229985621));
	notech_nand2 i_61665082(.A(divr_0[57]), .B(n_59903), .Z(n_230085622));
	notech_nand2 i_62065079(.A(divr_0[58]), .B(n_59903), .Z(n_230185623));
	notech_nand2 i_62365076(.A(divr_0[59]), .B(n_59903), .Z(n_230285624));
	notech_nand2 i_62665073(.A(divr_0[60]), .B(n_59903), .Z(n_230385625));
	notech_nand2 i_62965070(.A(divr_0[61]), .B(n_59903), .Z(n_230485626));
	notech_ao4 i_161365667(.A(n_2271), .B(n_59903), .C(n_172781715), .D(opc[
		31]), .Z(n_230585627));
	notech_nand2 i_63265067(.A(divr_0[62]), .B(n_59903), .Z(n_230685628));
	notech_nand2 i_63665063(.A(divr_0[63]), .B(n_59908), .Z(n_230885630));
	notech_and2 i_7165683(.A(n_265185971), .B(n_237685696), .Z(n_237585695)
		);
	notech_nand2 i_83764863(.A(n_275888699), .B(n_59908), .Z(n_237685696));
	notech_and2 i_84064860(.A(n_59826), .B(n_238085700), .Z(n_237985699));
	notech_nand3 i_2565643(.A(n_57415), .B(n_57417), .C(n_57387), .Z(n_238085700
		));
	notech_or4 i_85364847(.A(n_60536), .B(n_2258), .C(n_55149), .D(n_62419),
		 .Z(n_238285702));
	notech_or4 i_91464786(.A(n_60761), .B(n_60719), .C(n_60586), .D(n_238485704
		), .Z(n_238385703));
	notech_and3 i_065663(.A(n_57423), .B(n_57380), .C(n_238585705), .Z(n_238485704
		));
	notech_nand2 i_91564785(.A(n_2771), .B(n_55324), .Z(n_238585705));
	notech_or4 i_91664784(.A(n_56117), .B(n_59967), .C(n_59210), .D(n_60468)
		, .Z(n_238685706));
	notech_and4 i_16252(.A(n_26867), .B(n_2042), .C(n_26666), .D(n_59826), .Z
		(n_238785707));
	notech_ao3 i_16256(.A(calc_sz[1]), .B(n_56569), .C(n_223785560), .Z(n_238885708
		));
	notech_nand2 i_3365635(.A(n_26604), .B(n_59908), .Z(n_238985709));
	notech_nand2 i_3665632(.A(write_data_33[0]), .B(n_59908), .Z(n_239485714
		));
	notech_or2 i_4565623(.A(n_54754), .B(n_27371), .Z(n_239985719));
	notech_or2 i_5065618(.A(n_54754), .B(n_27372), .Z(n_240485724));
	notech_or2 i_5565613(.A(n_54754), .B(n_27373), .Z(n_240985729));
	notech_or2 i_6065608(.A(n_54754), .B(n_27374), .Z(n_241485734));
	notech_or2 i_6565603(.A(n_54754), .B(n_27376), .Z(n_241985739));
	notech_or2 i_7065598(.A(n_54754), .B(n_27378), .Z(n_242485744));
	notech_or2 i_7765593(.A(n_54754), .B(n_27385), .Z(n_242985749));
	notech_nand2 i_8265588(.A(write_data_33[22]), .B(n_59908), .Z(n_243485754
		));
	notech_nand2 i_8765583(.A(write_data_33[23]), .B(n_59908), .Z(n_243985759
		));
	notech_nand2 i_9265578(.A(write_data_33[24]), .B(n_59908), .Z(n_244485764
		));
	notech_nand2 i_9765573(.A(write_data_33[25]), .B(n_59908), .Z(n_244985769
		));
	notech_nand2 i_10265568(.A(write_data_33[26]), .B(n_59908), .Z(n_245485774
		));
	notech_nand2 i_10765563(.A(write_data_33[27]), .B(n_59908), .Z(n_245985779
		));
	notech_nand2 i_11265558(.A(write_data_33[28]), .B(n_59908), .Z(n_246485784
		));
	notech_nand2 i_11765553(.A(write_data_33[29]), .B(n_59907), .Z(n_246985789
		));
	notech_nand2 i_12265548(.A(write_data_33[30]), .B(n_59907), .Z(n_247485794
		));
	notech_nand2 i_12765543(.A(write_data_33[31]), .B(n_59907), .Z(n_247985799
		));
	notech_and2 i_16362(.A(n_223485557), .B(regs_10[0]), .Z(n_248085800));
	notech_and2 i_16364(.A(n_223485557), .B(regs_10[1]), .Z(n_248185801));
	notech_and2 i_16365(.A(n_223485557), .B(regs_10[2]), .Z(n_248285802));
	notech_and2 i_16366(.A(n_223485557), .B(regs_10[3]), .Z(n_248385803));
	notech_and2 i_16367(.A(n_223485557), .B(regs_10[4]), .Z(n_248485804));
	notech_and2 i_16368(.A(n_223485557), .B(regs_10[5]), .Z(n_248585805));
	notech_and2 i_16369(.A(n_223485557), .B(regs_10[6]), .Z(n_248685806));
	notech_and2 i_16370(.A(n_223485557), .B(regs_10[7]), .Z(n_248785807));
	notech_and2 i_16371(.A(n_223485557), .B(regs_10[8]), .Z(n_248885808));
	notech_and2 i_16372(.A(n_223485557), .B(regs_10[9]), .Z(n_248985809));
	notech_and2 i_16373(.A(n_223485557), .B(regs_10[10]), .Z(n_249085810));
	notech_and2 i_16374(.A(n_223485557), .B(regs_10[11]), .Z(n_249185811));
	notech_and2 i_16375(.A(n_223485557), .B(regs_10[12]), .Z(n_249285812));
	notech_and2 i_16376(.A(n_223485557), .B(regs_10[13]), .Z(n_249385813));
	notech_and2 i_16377(.A(n_223485557), .B(regs_10[14]), .Z(n_249485814));
	notech_and2 i_16378(.A(n_223485557), .B(regs_10[15]), .Z(n_249585815));
	notech_and2 i_16379(.A(n_52518), .B(regs_10[16]), .Z(n_249685816));
	notech_and2 i_16380(.A(n_52518), .B(regs_10[17]), .Z(n_249785817));
	notech_and2 i_16381(.A(n_52518), .B(regs_10[18]), .Z(n_249885818));
	notech_and2 i_16382(.A(n_52518), .B(regs_10[19]), .Z(n_249985819));
	notech_and2 i_16383(.A(n_52518), .B(regs_10[20]), .Z(n_250085820));
	notech_and2 i_16384(.A(n_52518), .B(regs_10[21]), .Z(n_250185821));
	notech_and2 i_16385(.A(n_52518), .B(regs_10[22]), .Z(n_250285822));
	notech_and2 i_16386(.A(n_52518), .B(regs_10[23]), .Z(n_250385823));
	notech_and2 i_16387(.A(regs_10[24]), .B(n_52518), .Z(n_250485824));
	notech_and2 i_16388(.A(n_52518), .B(regs_10[25]), .Z(n_250585825));
	notech_and2 i_16389(.A(n_52518), .B(regs_10[26]), .Z(n_250685826));
	notech_and2 i_16390(.A(n_52518), .B(regs_10[27]), .Z(n_250785827));
	notech_and2 i_16391(.A(n_52518), .B(regs_10[28]), .Z(n_250885828));
	notech_and2 i_16392(.A(n_52518), .B(regs_10[29]), .Z(n_250985829));
	notech_and2 i_16393(.A(n_52518), .B(regs_10[30]), .Z(n_251085830));
	notech_and2 i_16394(.A(n_52518), .B(regs_10[31]), .Z(n_251185831));
	notech_ao3 i_16895(.A(tcmp_arithbox), .B(n_59828), .C(n_57424), .Z(n_251285832
		));
	notech_or4 i_13065540(.A(n_1845), .B(n_326546823), .C(n_223985562), .D(n_207241703
		), .Z(n_251385833));
	notech_ao3 i_13165539(.A(n_620), .B(n_55040), .C(n_59364), .Z(n_251485834
		));
	notech_ao3 i_21758(.A(n_2771), .B(n_59828), .C(pipe_mul[0]), .Z(n_264385963
		));
	notech_and3 i_21760(.A(n_223585558), .B(n_2771), .C(n_59828), .Z(n_264485964
		));
	notech_nand3 i_42165716(.A(n_54727), .B(n_51840), .C(n_54967), .Z(n_264885968
		));
	notech_nao3 i_19365682(.A(n_244056258), .B(n_59907), .C(n_2582), .Z(n_265085970
		));
	notech_ao4 i_151065668(.A(n_58895), .B(n_1967), .C(n_2772), .D(n_59907),
		 .Z(n_265185971));
	notech_ao4 i_133664368(.A(n_54388), .B(n_29777), .C(n_207041701), .D(n_59095
		), .Z(n_265285972));
	notech_ao4 i_133564369(.A(n_54388), .B(n_29775), .C(n_54373), .D(n_59050
		), .Z(n_265385973));
	notech_ao4 i_133464370(.A(n_54388), .B(n_29774), .C(n_54373), .D(n_59104
		), .Z(n_265485974));
	notech_ao4 i_133364371(.A(n_54389), .B(n_29773), .C(n_54373), .D(nbus_11326
		[28]), .Z(n_265585975));
	notech_ao4 i_133264372(.A(n_54389), .B(n_29771), .C(n_54373), .D(nbus_11326
		[27]), .Z(n_265685976));
	notech_ao4 i_133164373(.A(n_54388), .B(n_29770), .C(n_54373), .D(n_59068
		), .Z(n_265785977));
	notech_ao4 i_133064374(.A(n_54388), .B(n_29769), .C(n_54373), .D(n_59023
		), .Z(n_265885978));
	notech_ao4 i_132964375(.A(n_54388), .B(n_29768), .C(n_54373), .D(n_59086
		), .Z(n_265985979));
	notech_ao4 i_132864376(.A(n_54388), .B(n_29767), .C(n_54373), .D(n_59041
		), .Z(n_266085980));
	notech_ao4 i_132764377(.A(n_54388), .B(n_29766), .C(n_54369), .D(n_59032
		), .Z(n_266185981));
	notech_ao4 i_132664378(.A(n_54388), .B(n_29765), .C(n_54369), .D(n_58996
		), .Z(n_266285982));
	notech_ao4 i_132564379(.A(n_54388), .B(n_29764), .C(n_54369), .D(n_59005
		), .Z(n_266385983));
	notech_ao4 i_132464380(.A(n_54388), .B(n_29763), .C(n_54373), .D(n_59014
		), .Z(n_266485984));
	notech_ao4 i_132364381(.A(n_54388), .B(n_29762), .C(n_54373), .D(n_58969
		), .Z(n_266585985));
	notech_ao4 i_132264382(.A(n_54388), .B(n_29759), .C(n_54373), .D(nbus_11326
		[17]), .Z(n_266685986));
	notech_ao4 i_132164383(.A(n_54389), .B(n_29758), .C(n_54373), .D(nbus_11326
		[16]), .Z(n_266785987));
	notech_ao4 i_132064384(.A(n_54389), .B(n_29757), .C(n_54373), .D(nbus_11326
		[15]), .Z(n_266885988));
	notech_ao4 i_131964385(.A(n_54389), .B(n_29756), .C(n_54374), .D(nbus_11326
		[14]), .Z(n_266985989));
	notech_ao4 i_131864386(.A(n_54389), .B(n_29755), .C(n_54374), .D(nbus_11326
		[13]), .Z(n_267085990));
	notech_ao4 i_131764387(.A(n_54389), .B(n_29754), .C(n_54374), .D(nbus_11326
		[12]), .Z(n_267185991));
	notech_ao4 i_131664388(.A(n_54389), .B(n_29753), .C(n_54374), .D(nbus_11326
		[11]), .Z(n_267285992));
	notech_ao4 i_131564389(.A(n_54389), .B(n_29752), .C(n_54374), .D(nbus_11326
		[10]), .Z(n_267385993));
	notech_ao4 i_131464390(.A(n_54389), .B(n_29751), .C(n_54374), .D(nbus_11326
		[9]), .Z(n_267485994));
	notech_ao4 i_131364391(.A(n_54389), .B(n_29750), .C(n_54374), .D(nbus_11326
		[8]), .Z(n_267585995));
	notech_ao4 i_131264392(.A(n_54389), .B(n_29749), .C(n_54374), .D(nbus_11326
		[7]), .Z(n_267685996));
	notech_ao4 i_131164393(.A(n_54389), .B(n_29748), .C(n_54374), .D(nbus_11326
		[6]), .Z(n_267785997));
	notech_ao4 i_131064394(.A(n_54389), .B(n_29747), .C(n_54374), .D(nbus_11326
		[5]), .Z(n_267885998));
	notech_ao4 i_130964395(.A(n_54389), .B(n_29746), .C(n_54373), .D(nbus_11326
		[4]), .Z(n_267985999));
	notech_ao4 i_130864396(.A(n_54389), .B(n_29745), .C(n_54374), .D(nbus_11326
		[3]), .Z(n_268086000));
	notech_ao4 i_130764397(.A(n_54389), .B(n_29744), .C(n_54374), .D(nbus_11326
		[2]), .Z(n_268186001));
	notech_ao4 i_130664398(.A(n_54389), .B(n_29743), .C(n_54374), .D(nbus_11326
		[1]), .Z(n_268286002));
	notech_ao4 i_130564399(.A(n_54388), .B(n_29742), .C(n_54374), .D(nbus_11326
		[0]), .Z(n_268386003));
	notech_ao4 i_130464400(.A(n_54383), .B(n_29741), .C(n_54369), .D(n_58951
		), .Z(n_268486004));
	notech_ao4 i_130364401(.A(n_54383), .B(n_29740), .C(n_54365), .D(n_56901
		), .Z(n_268586005));
	notech_ao4 i_130264402(.A(n_54378), .B(n_29739), .C(n_54365), .D(n_56892
		), .Z(n_268686006));
	notech_ao4 i_130164403(.A(n_54378), .B(n_29738), .C(n_54365), .D(n_56883
		), .Z(n_268786007));
	notech_ao4 i_130064404(.A(n_54383), .B(n_29737), .C(n_54365), .D(n_56874
		), .Z(n_268886008));
	notech_ao4 i_129964405(.A(n_54383), .B(n_29736), .C(n_54365), .D(n_56865
		), .Z(n_268986009));
	notech_ao4 i_129864406(.A(n_54383), .B(n_29735), .C(n_54365), .D(n_56856
		), .Z(n_269086010));
	notech_ao4 i_129764407(.A(n_54383), .B(n_29734), .C(n_54365), .D(n_56847
		), .Z(n_269186011));
	notech_ao4 i_129664408(.A(n_54378), .B(n_29733), .C(n_54365), .D(n_56838
		), .Z(n_269286012));
	notech_ao4 i_129564409(.A(n_54378), .B(n_29732), .C(n_54364), .D(n_56829
		), .Z(n_269386013));
	notech_ao4 i_129464410(.A(n_54378), .B(n_29731), .C(n_54364), .D(n_56820
		), .Z(n_269486014));
	notech_ao4 i_129364411(.A(n_54378), .B(n_29730), .C(n_54364), .D(n_56811
		), .Z(n_269586015));
	notech_ao4 i_129264412(.A(n_54378), .B(n_29729), .C(n_54364), .D(n_56802
		), .Z(n_269686016));
	notech_ao4 i_129164413(.A(n_54378), .B(n_29728), .C(n_54364), .D(n_56793
		), .Z(n_269786017));
	notech_ao4 i_129064414(.A(n_54378), .B(n_29727), .C(n_54364), .D(n_56784
		), .Z(n_269886018));
	notech_ao4 i_128964415(.A(n_54378), .B(n_29726), .C(n_54364), .D(n_56775
		), .Z(n_269986019));
	notech_ao4 i_128864416(.A(n_54383), .B(n_29725), .C(n_54365), .D(n_56766
		), .Z(n_270086020));
	notech_ao4 i_128764417(.A(n_54383), .B(n_29724), .C(n_54369), .D(nbus_11273
		[14]), .Z(n_270186021));
	notech_ao4 i_128664418(.A(n_54383), .B(n_29723), .C(n_54369), .D(n_56748
		), .Z(n_270286022));
	notech_ao4 i_128564419(.A(n_54383), .B(n_29722), .C(n_54369), .D(n_56739
		), .Z(n_270386023));
	notech_ao4 i_128464420(.A(n_54388), .B(n_29721), .C(n_54369), .D(n_56730
		), .Z(n_270486024));
	notech_ao4 i_128364421(.A(n_54388), .B(n_29720), .C(n_54369), .D(n_56721
		), .Z(n_270586025));
	notech_ao4 i_128264422(.A(n_54383), .B(n_29719), .C(n_54369), .D(n_56712
		), .Z(n_270686026));
	notech_ao4 i_128164423(.A(n_54383), .B(n_29718), .C(n_54369), .D(n_56703
		), .Z(n_270786027));
	notech_ao4 i_128064424(.A(n_54383), .B(n_29717), .C(n_54369), .D(n_57326
		), .Z(n_270886028));
	notech_ao4 i_127964425(.A(n_54383), .B(n_29716), .C(n_54365), .D(n_56694
		), .Z(n_270986029));
	notech_ao4 i_127864426(.A(n_54383), .B(n_29715), .C(n_54365), .D(nbus_11273
		[5]), .Z(n_271086030));
	notech_ao4 i_127764427(.A(n_54383), .B(n_29714), .C(n_54365), .D(n_56676
		), .Z(n_271186031));
	notech_ao4 i_127664428(.A(n_54383), .B(n_29713), .C(n_54365), .D(n_56667
		), .Z(n_271286032));
	notech_ao4 i_127564429(.A(n_54383), .B(n_29712), .C(n_54369), .D(n_56658
		), .Z(n_271386033));
	notech_ao4 i_127464430(.A(n_54383), .B(n_29711), .C(n_54369), .D(n_56649
		), .Z(n_271486034));
	notech_ao4 i_127364431(.A(n_54383), .B(n_29710), .C(n_54365), .D(n_58960
		), .Z(n_271586035));
	notech_ao4 i_99364707(.A(n_54754), .B(n_27401), .C(n_55943), .D(nbus_11326
		[31]), .Z(n_271986039));
	notech_ao4 i_99264708(.A(n_54637), .B(n_27785), .C(n_56943), .D(n_26608)
		, .Z(n_272186041));
	notech_ao4 i_99064710(.A(n_54754), .B(n_27400), .C(n_58505), .D(nbus_11326
		[30]), .Z(n_272286042));
	notech_ao4 i_98964711(.A(n_54637), .B(n_27784), .C(n_55234), .D(n_26608)
		, .Z(n_272486044));
	notech_ao4 i_98764713(.A(n_54754), .B(n_27399), .C(n_58505), .D(nbus_11326
		[29]), .Z(n_272586045));
	notech_ao4 i_98664714(.A(n_54637), .B(n_27783), .C(n_55249), .D(n_26608)
		, .Z(n_272786047));
	notech_ao4 i_98464716(.A(n_54754), .B(n_27398), .C(n_58505), .D(n_59077)
		, .Z(n_272886048));
	notech_ao4 i_98364717(.A(n_54637), .B(n_27782), .C(n_55261), .D(n_26608)
		, .Z(n_273086050));
	notech_ao4 i_98164719(.A(n_54754), .B(n_27397), .C(n_58505), .D(n_59059)
		, .Z(n_273186051));
	notech_ao4 i_98064720(.A(n_54637), .B(n_27781), .C(n_59328), .D(n_26608)
		, .Z(n_273386053));
	notech_ao4 i_97864722(.A(n_54762), .B(n_27396), .C(n_58505), .D(n_59068)
		, .Z(n_273486054));
	notech_ao4 i_97764723(.A(n_54637), .B(n_27780), .C(n_59337), .D(n_26608)
		, .Z(n_273686056));
	notech_ao4 i_97564725(.A(n_54754), .B(n_27395), .C(n_58505), .D(n_59023)
		, .Z(n_273786057));
	notech_ao4 i_97464726(.A(n_54637), .B(n_27779), .C(n_59346), .D(n_26608)
		, .Z(n_273986059));
	notech_ao4 i_97264728(.A(n_54754), .B(n_27394), .C(n_58505), .D(n_59086)
		, .Z(n_274086060));
	notech_ao4 i_97164729(.A(n_54637), .B(n_27778), .C(n_56207), .D(n_26608)
		, .Z(n_274286062));
	notech_ao4 i_96964731(.A(n_54754), .B(n_27393), .C(n_58505), .D(n_59041)
		, .Z(n_274386063));
	notech_ao4 i_96864732(.A(n_54637), .B(n_27777), .C(n_26608), .D(n_59319)
		, .Z(n_274586065));
	notech_ao4 i_96664734(.A(n_54754), .B(n_27392), .C(n_58505), .D(n_59032)
		, .Z(n_274686066));
	notech_ao4 i_96564735(.A(n_54637), .B(n_27774), .C(n_26608), .D(n_55647)
		, .Z(n_274886068));
	notech_ao4 i_96364737(.A(n_58505), .B(nbus_11326[15]), .C(n_55578), .D(n_26610
		), .Z(n_274986069));
	notech_ao4 i_96264738(.A(n_54637), .B(n_27764), .C(n_59828), .D(n_28890)
		, .Z(n_275186071));
	notech_ao4 i_96064740(.A(n_58505), .B(nbus_11326[8]), .C(n_55413), .D(n_26610
		), .Z(n_275286072));
	notech_ao4 i_95964741(.A(n_54637), .B(n_27755), .C(n_59828), .D(n_28883)
		, .Z(n_275486074));
	notech_ao4 i_95764743(.A(n_58505), .B(nbus_11326[6]), .C(n_55387), .D(n_26610
		), .Z(n_275586075));
	notech_ao4 i_95664744(.A(n_54642), .B(n_27753), .C(n_59828), .D(n_28881)
		, .Z(n_275786077));
	notech_ao4 i_95464746(.A(n_58505), .B(nbus_11326[4]), .C(n_55365), .D(n_26610
		), .Z(n_275886078));
	notech_ao4 i_95364747(.A(n_54637), .B(n_27751), .C(n_59828), .D(n_28879)
		, .Z(n_276086080));
	notech_ao4 i_95164749(.A(n_58505), .B(nbus_11326[3]), .C(n_55277), .D(n_26610
		), .Z(n_276186081));
	notech_ao4 i_95064750(.A(n_54637), .B(n_27750), .C(n_59828), .D(n_28878)
		, .Z(n_276386083));
	notech_ao4 i_94864752(.A(n_58505), .B(nbus_11326[2]), .C(n_55289), .D(n_26610
		), .Z(n_276486084));
	notech_ao4 i_94764753(.A(n_54637), .B(n_27749), .C(n_59828), .D(n_28876)
		, .Z(n_276686086));
	notech_ao4 i_94564755(.A(n_58505), .B(nbus_11326[1]), .C(n_26610), .D(n_59753
		), .Z(n_276786087));
	notech_ao4 i_94464756(.A(n_54637), .B(n_27748), .C(n_59828), .D(n_28875)
		, .Z(n_276986089));
	notech_ao4 i_92564775(.A(n_54754), .B(n_27370), .C(n_58505), .D(nbus_11326
		[0]), .Z(n_277086090));
	notech_ao4 i_92464776(.A(n_54637), .B(n_27747), .C(n_26608), .D(\nbus_11276[0] 
		), .Z(n_277286092));
	notech_nand2 i_92164779(.A(calc_sz[2]), .B(n_56569), .Z(n_277586095));
	notech_ao4 i_18763364(.A(n_2582), .B(n_2599), .C(n_278086100), .D(n_26612
		), .Z(n_277886098));
	notech_ao4 i_14063411(.A(n_57458), .B(n_57441), .C(n_278286102), .D(n_177260854
		), .Z(n_278086100));
	notech_ao4 i_11063438(.A(n_2585), .B(n_2582), .C(n_278486104), .D(n_26614
		), .Z(n_278286102));
	notech_and2 i_8363464(.A(n_2822), .B(n_275188706), .Z(n_278486104));
	notech_ao4 i_149262100(.A(n_53113), .B(n_27334), .C(n_53964), .D(n_27298
		), .Z(n_279386113));
	notech_ao4 i_149162101(.A(n_56336), .B(n_26925), .C(n_53234), .D(n_29779
		), .Z(n_279486114));
	notech_ao4 i_148462108(.A(n_27365), .B(n_52811), .C(n_53937), .D(n_27332
		), .Z(n_279586115));
	notech_ao4 i_148362109(.A(n_56511), .B(n_26987), .C(n_52930), .D(n_29778
		), .Z(n_279686116));
	notech_xor2 i_3255267(.A(vliw_pc[0]), .B(vliw_pc[1]), .Z(n_279786117));
	notech_xor2 i_3355266(.A(n_2789), .B(vliw_pc[2]), .Z(n_279886118));
	notech_xor2 i_3455265(.A(n_2790), .B(vliw_pc[3]), .Z(n_279986119));
	notech_ao4 i_3555264(.A(n_2832), .B(n_2790), .C(n_280786127), .D(n_27268
		), .Z(n_280086120));
	notech_ao4 i_54055317(.A(n_59150), .B(n_273488721), .C(n_60468), .D(n_281086130
		), .Z(n_280186121));
	notech_and4 i_2355275(.A(vliw_pc[1]), .B(vliw_pc[0]), .C(vliw_pc[2]), .D
		(vliw_pc[3]), .Z(n_280786127));
	notech_and4 i_3155268(.A(n_26785), .B(n_2042), .C(reps[2]), .D(n_27081),
		 .Z(n_281086130));
	notech_and2 i_16763(.A(n_279786117), .B(n_26617), .Z(n_281486134));
	notech_nor2 i_16764(.A(n_280186121), .B(n_279886118), .Z(n_281586135));
	notech_nor2 i_16765(.A(n_280186121), .B(n_279986119), .Z(n_281686136));
	notech_nor2 i_16766(.A(n_280186121), .B(n_280086120), .Z(n_281786137));
	notech_ao4 i_122354123(.A(n_54886), .B(n_59150), .C(vliw_pc[0]), .D(n_280186121
		), .Z(n_281886138));
	notech_or2 i_12949033(.A(n_53276), .B(n_271088745), .Z(n_281986139));
	notech_nand3 i_12849034(.A(n_60525), .B(n_26772), .C(temp_sp[31]), .Z(n_282286142
		));
	notech_nand3 i_3217834(.A(n_287786197), .B(n_281986139), .C(n_282286142)
		, .Z(write_data_26[31]));
	notech_or2 i_129647936(.A(n_54836), .B(n_28082), .Z(n_282386143));
	notech_nand3 i_3216841(.A(n_288086200), .B(n_287986199), .C(n_288686206)
		, .Z(n_9862));
	notech_or2 i_131547918(.A(n_54836), .B(n_28081), .Z(n_283286152));
	notech_nand3 i_3116840(.A(n_288886208), .B(n_288786207), .C(n_289486214)
		, .Z(n_9857));
	notech_or2 i_133547900(.A(n_54836), .B(n_28080), .Z(n_284186161));
	notech_nand3 i_3016839(.A(n_289686216), .B(n_289586215), .C(n_290286222)
		, .Z(n_9852));
	notech_or4 i_135347882(.A(n_244656264), .B(n_57404), .C(n_59908), .D(n_59077
		), .Z(n_285086170));
	notech_nand3 i_2916838(.A(n_290486224), .B(n_290386223), .C(n_291086230)
		, .Z(n_9847));
	notech_or4 i_137247864(.A(n_57383), .B(n_57404), .C(n_59908), .D(n_59059
		), .Z(n_285986179));
	notech_nand3 i_2816837(.A(n_291286232), .B(n_291186231), .C(n_291886238)
		, .Z(n_9842));
	notech_or4 i_157947666(.A(n_57383), .B(n_57404), .C(n_59908), .D(n_58987
		), .Z(n_286886188));
	notech_nand3 i_1716826(.A(n_292086240), .B(n_291986239), .C(n_292686246)
		, .Z(n_9787));
	notech_ao4 i_13049032(.A(n_53296), .B(n_27332), .C(n_53285), .D(n_27365)
		, .Z(n_287786197));
	notech_ao4 i_130847925(.A(n_54926), .B(nbus_11348[31]), .C(n_54908), .D(n_29780
		), .Z(n_287986199));
	notech_ao4 i_130947924(.A(n_54940), .B(n_29781), .C(n_56631), .D(n_29460
		), .Z(n_288086200));
	notech_ao4 i_131047923(.A(n_54863), .B(n_56943), .C(n_55122), .D(n_59095
		), .Z(n_288286202));
	notech_ao4 i_130747926(.A(n_54887), .B(n_28931), .C(n_54847), .D(nbus_11326
		[7]), .Z(n_288486204));
	notech_and4 i_131347920(.A(n_2312), .B(n_288486204), .C(n_288286202), .D
		(n_282386143), .Z(n_288686206));
	notech_ao4 i_132847907(.A(n_54926), .B(nbus_11348[30]), .C(n_54908), .D(n_29782
		), .Z(n_288786207));
	notech_ao4 i_132947906(.A(n_54940), .B(n_29783), .C(n_56631), .D(n_29458
		), .Z(n_288886208));
	notech_ao4 i_133047905(.A(n_54863), .B(\nbus_11276[30] ), .C(n_55122), .D
		(n_59050), .Z(n_289086210));
	notech_ao4 i_132747908(.A(n_54887), .B(n_28930), .C(n_54847), .D(nbus_11326
		[6]), .Z(n_289286212));
	notech_and4 i_133347902(.A(n_2312), .B(n_289286212), .C(n_289086210), .D
		(n_283286152), .Z(n_289486214));
	notech_ao4 i_134647889(.A(n_54926), .B(nbus_11348[29]), .C(n_54908), .D(n_29784
		), .Z(n_289586215));
	notech_ao4 i_134747888(.A(n_54940), .B(n_29785), .C(n_56631), .D(n_29462
		), .Z(n_289686216));
	notech_ao4 i_134847887(.A(n_54863), .B(\nbus_11276[29] ), .C(n_55122), .D
		(n_59104), .Z(n_289886218));
	notech_ao4 i_134547890(.A(n_54887), .B(n_28929), .C(n_54847), .D(nbus_11326
		[5]), .Z(n_290086220));
	notech_and4 i_135147884(.A(n_2312), .B(n_290086220), .C(n_289886218), .D
		(n_284186161), .Z(n_290286222));
	notech_ao4 i_136547871(.A(n_54887), .B(n_28928), .C(n_54863), .D(n_55261
		), .Z(n_290386223));
	notech_ao4 i_136647870(.A(n_54926), .B(nbus_11348[28]), .C(n_54908), .D(n_29786
		), .Z(n_290486224));
	notech_ao4 i_136747869(.A(n_2249), .B(n_29787), .C(n_56631), .D(n_29459)
		, .Z(n_290686226));
	notech_ao4 i_136447872(.A(n_54847), .B(nbus_11326[4]), .C(n_54836), .D(n_28079
		), .Z(n_290886228));
	notech_and4 i_137047866(.A(n_2312), .B(n_290886228), .C(n_290686226), .D
		(n_285086170), .Z(n_291086230));
	notech_ao4 i_138347853(.A(n_54887), .B(n_28927), .C(n_54863), .D(n_59328
		), .Z(n_291186231));
	notech_ao4 i_138447852(.A(n_54926), .B(nbus_11348[27]), .C(n_54908), .D(n_29788
		), .Z(n_291286232));
	notech_ao4 i_138547851(.A(n_54940), .B(n_29789), .C(n_56631), .D(n_29461
		), .Z(n_291486234));
	notech_ao4 i_138247854(.A(n_54847), .B(nbus_11326[3]), .C(n_54836), .D(n_28078
		), .Z(n_291686236));
	notech_and4 i_138847848(.A(n_2312), .B(n_291686236), .C(n_291486234), .D
		(n_285986179), .Z(n_291886238));
	notech_ao4 i_159047655(.A(n_54887), .B(n_28916), .C(n_54863), .D(n_55590
		), .Z(n_291986239));
	notech_ao4 i_159147654(.A(n_54926), .B(nbus_11348[16]), .C(n_54908), .D(n_29790
		), .Z(n_292086240));
	notech_ao4 i_159247653(.A(n_54940), .B(n_29791), .C(n_56631), .D(n_29463
		), .Z(n_292286242));
	notech_ao4 i_158947656(.A(n_54847), .B(nbus_11326[8]), .C(n_54836), .D(n_28067
		), .Z(n_292486244));
	notech_and4 i_159547650(.A(n_2312), .B(n_292486244), .C(n_292286242), .D
		(n_286886188), .Z(n_292686246));
	notech_ao4 i_209143342(.A(n_56404), .B(n_26969), .C(n_53276), .D(n_308921976
		), .Z(n_294786267));
	notech_ao4 i_209043343(.A(n_53285), .B(n_27357), .C(n_53296), .D(n_27324
		), .Z(n_294886268));
	notech_ao4 i_207543358(.A(n_56404), .B(n_26973), .C(n_308821975), .D(n_53276
		), .Z(n_294986269));
	notech_ao4 i_207443359(.A(n_53285), .B(n_27359), .C(n_53296), .D(n_27326
		), .Z(n_295086270));
	notech_ao4 i_205943374(.A(n_56409), .B(n_26975), .C(n_53276), .D(n_308721974
		), .Z(n_295186271));
	notech_ao4 i_205843375(.A(n_53285), .B(n_27360), .C(n_53296), .D(n_27327
		), .Z(n_295286272));
	notech_ao4 i_204343390(.A(n_56409), .B(n_26977), .C(n_308621973), .D(n_53276
		), .Z(n_295386273));
	notech_ao4 i_204243391(.A(n_53285), .B(n_27361), .C(n_53296), .D(n_27328
		), .Z(n_295486274));
	notech_ao4 i_202743406(.A(n_56409), .B(n_26979), .C(n_57330), .D(n_53276
		), .Z(n_295586275));
	notech_ao4 i_202643407(.A(n_53285), .B(n_27362), .C(n_53296), .D(n_27329
		), .Z(n_295686276));
	notech_ao4 i_207140221(.A(n_56409), .B(n_26959), .C(n_53276), .D(n_311318890
		), .Z(n_297786297));
	notech_ao4 i_207040222(.A(n_53285), .B(n_27352), .C(n_53296), .D(n_27319
		), .Z(n_297886298));
	notech_ao4 i_205540237(.A(n_56409), .B(n_26961), .C(n_26595), .D(n_311218889
		), .Z(n_297986299));
	notech_ao4 i_205440238(.A(n_53285), .B(n_27353), .C(n_53296), .D(n_27320
		), .Z(n_298086300));
	notech_ao4 i_203940253(.A(n_56414), .B(n_26963), .C(n_53276), .D(n_311118888
		), .Z(n_298186301));
	notech_ao4 i_203840254(.A(n_53285), .B(n_27354), .C(n_53296), .D(n_27321
		), .Z(n_298286302));
	notech_ao4 i_202340269(.A(n_56414), .B(n_26965), .C(n_53276), .D(n_311018887
		), .Z(n_298386303));
	notech_ao4 i_202240270(.A(n_53285), .B(n_27355), .C(n_53296), .D(n_27322
		), .Z(n_298486304));
	notech_ao4 i_200740285(.A(n_56409), .B(n_26967), .C(n_53276), .D(n_26618
		), .Z(n_298586305));
	notech_ao4 i_200640286(.A(n_53285), .B(n_27356), .C(n_53296), .D(n_27323
		), .Z(n_298686306));
	notech_or2 i_13038963(.A(n_53276), .B(n_271888737), .Z(n_298786307));
	notech_nand3 i_12938964(.A(n_60525), .B(n_26772), .C(temp_sp[14]), .Z(n_299086310
		));
	notech_nand3 i_1517817(.A(n_299586315), .B(n_298786307), .C(n_299086310)
		, .Z(write_data_26[14]));
	notech_or2 i_16738926(.A(n_53276), .B(n_271988736), .Z(n_299186311));
	notech_nand3 i_16638927(.A(n_60525), .B(n_26772), .C(temp_sp[16]), .Z(n_299486314
		));
	notech_nand3 i_1717819(.A(n_299786317), .B(n_299186311), .C(n_299486314)
		, .Z(write_data_26[16]));
	notech_ao4 i_13138962(.A(n_53296), .B(n_27315), .C(n_53285), .D(n_27348)
		, .Z(n_299586315));
	notech_ao4 i_16838925(.A(n_53296), .B(n_27317), .C(n_53285), .D(n_27350)
		, .Z(n_299786317));
	notech_or4 i_16745(.A(n_2831), .B(n_57404), .C(n_59364), .D(n_60468), .Z
		(n_299986319));
	notech_or4 i_48389(.A(n_274588712), .B(n_59967), .C(n_59958), .D(n_60468
		), .Z(n_300186321));
	notech_or4 i_117334576(.A(n_60761), .B(n_60719), .C(n_57418), .D(n_60586
		), .Z(n_300286322));
	notech_nand2 i_1617818(.A(n_113084457), .B(n_112984456), .Z(write_data_26
		[15]));
	notech_nand2 i_318061(.A(n_113284459), .B(n_113184458), .Z(write_data_28
		[2]));
	notech_nand2 i_418062(.A(n_113484461), .B(n_113384460), .Z(write_data_28
		[3]));
	notech_nand2 i_518063(.A(n_113684463), .B(n_113584462), .Z(write_data_28
		[4]));
	notech_nand2 i_618064(.A(n_113884465), .B(n_113784464), .Z(write_data_28
		[5]));
	notech_nand2 i_718065(.A(n_114084467), .B(n_113984466), .Z(write_data_28
		[6]));
	notech_nand2 i_818066(.A(n_114284469), .B(n_114184468), .Z(write_data_28
		[7]));
	notech_nand2 i_918067(.A(n_114484471), .B(n_114384470), .Z(write_data_28
		[8]));
	notech_nand2 i_1018068(.A(n_114684473), .B(n_114584472), .Z(write_data_28
		[9]));
	notech_nand2 i_1118069(.A(n_114884475), .B(n_114784474), .Z(write_data_28
		[10]));
	notech_nand2 i_1218070(.A(n_115084477), .B(n_114984476), .Z(write_data_28
		[11]));
	notech_nand2 i_1318071(.A(n_115284479), .B(n_115184478), .Z(write_data_28
		[12]));
	notech_nand2 i_1418072(.A(n_115484481), .B(n_115384480), .Z(write_data_28
		[13]));
	notech_nand2 i_1518073(.A(n_115684483), .B(n_115584482), .Z(write_data_28
		[14]));
	notech_nand2 i_1618074(.A(n_115884485), .B(n_115784484), .Z(write_data_28
		[15]));
	notech_nand2 i_1718075(.A(n_116084487), .B(n_115984486), .Z(write_data_28
		[16]));
	notech_nand2 i_1818076(.A(n_116284489), .B(n_116184488), .Z(write_data_28
		[17]));
	notech_nand2 i_1918077(.A(n_116484491), .B(n_116384490), .Z(write_data_28
		[18]));
	notech_nand2 i_2018078(.A(n_116684493), .B(n_116584492), .Z(write_data_28
		[19]));
	notech_nand2 i_2118079(.A(n_116884495), .B(n_116784494), .Z(write_data_28
		[20]));
	notech_nand2 i_2218080(.A(n_117084497), .B(n_116984496), .Z(write_data_28
		[21]));
	notech_nand2 i_2318081(.A(n_117284499), .B(n_117184498), .Z(write_data_28
		[22]));
	notech_nand2 i_2418082(.A(n_117484501), .B(n_117384500), .Z(write_data_28
		[23]));
	notech_nand2 i_2518083(.A(n_117684503), .B(n_117584502), .Z(write_data_28
		[24]));
	notech_nand2 i_2618084(.A(n_117884505), .B(n_117784504), .Z(write_data_28
		[25]));
	notech_nand2 i_2718085(.A(n_118084507), .B(n_117984506), .Z(write_data_28
		[26]));
	notech_nand2 i_2818086(.A(n_118284509), .B(n_118184508), .Z(write_data_28
		[27]));
	notech_nand2 i_2918087(.A(n_118484511), .B(n_118384510), .Z(write_data_28
		[28]));
	notech_nand2 i_3018088(.A(n_118684513), .B(n_118584512), .Z(write_data_28
		[29]));
	notech_nand2 i_3118089(.A(n_118884515), .B(n_118784514), .Z(write_data_28
		[30]));
	notech_nand2 i_3218090(.A(n_119084517), .B(n_118984516), .Z(write_data_28
		[31]));
	notech_nand2 i_118315(.A(n_119284519), .B(n_119184518), .Z(write_data_30
		[0]));
	notech_nand2 i_218316(.A(n_119484521), .B(n_119384520), .Z(write_data_30
		[1]));
	notech_nand2 i_318317(.A(n_119684523), .B(n_119584522), .Z(write_data_30
		[2]));
	notech_nand2 i_418318(.A(n_119884525), .B(n_119784524), .Z(write_data_30
		[3]));
	notech_nand2 i_518319(.A(n_120084527), .B(n_119984526), .Z(write_data_30
		[4]));
	notech_nand2 i_618320(.A(n_120284529), .B(n_120184528), .Z(write_data_30
		[5]));
	notech_nand2 i_718321(.A(n_120484531), .B(n_120384530), .Z(write_data_30
		[6]));
	notech_nand2 i_818322(.A(n_120684533), .B(n_120584532), .Z(write_data_30
		[7]));
	notech_nand2 i_918323(.A(n_120884535), .B(n_120784534), .Z(write_data_30
		[8]));
	notech_nand2 i_1018324(.A(n_121084537), .B(n_120984536), .Z(write_data_30
		[9]));
	notech_nand2 i_1118325(.A(n_121284539), .B(n_121184538), .Z(write_data_30
		[10]));
	notech_nand2 i_1218326(.A(n_121484541), .B(n_121384540), .Z(write_data_30
		[11]));
	notech_nand2 i_1318327(.A(n_121684543), .B(n_121584542), .Z(write_data_30
		[12]));
	notech_nand2 i_1418328(.A(n_121884545), .B(n_121784544), .Z(write_data_30
		[13]));
	notech_nand2 i_1518329(.A(n_122084547), .B(n_121984546), .Z(write_data_30
		[14]));
	notech_nand2 i_1618330(.A(n_122284549), .B(n_122184548), .Z(write_data_30
		[15]));
	notech_nand2 i_1818332(.A(n_122484551), .B(n_122384550), .Z(write_data_30
		[17]));
	notech_nand2 i_1918333(.A(n_122684553), .B(n_122584552), .Z(write_data_30
		[18]));
	notech_nand2 i_2018334(.A(n_122884555), .B(n_122784554), .Z(write_data_30
		[19]));
	notech_nand2 i_2118335(.A(n_123084557), .B(n_122984556), .Z(write_data_30
		[20]));
	notech_nand2 i_2218336(.A(n_123284559), .B(n_123184558), .Z(write_data_30
		[21]));
	notech_nand2 i_2318337(.A(n_123484561), .B(n_123384560), .Z(write_data_30
		[22]));
	notech_nand2 i_2418338(.A(n_123684563), .B(n_123584562), .Z(write_data_30
		[23]));
	notech_nand2 i_2518339(.A(n_123884565), .B(n_123784564), .Z(write_data_30
		[24]));
	notech_nand2 i_2618340(.A(n_124084567), .B(n_123984566), .Z(write_data_30
		[25]));
	notech_nand2 i_2718341(.A(n_124284569), .B(n_124184568), .Z(write_data_30
		[26]));
	notech_nand2 i_2818342(.A(n_124484571), .B(n_124384570), .Z(write_data_30
		[27]));
	notech_nand2 i_2918343(.A(n_124684573), .B(n_124584572), .Z(write_data_30
		[28]));
	notech_nand2 i_3018344(.A(n_124884575), .B(n_124784574), .Z(write_data_30
		[29]));
	notech_nand2 i_3118345(.A(n_125084577), .B(n_124984576), .Z(write_data_30
		[30]));
	notech_nao3 i_25268311(.A(n_253034156), .B(n_26621), .C(n_57417), .Z(n_300586325
		));
	notech_or4 i_16241(.A(n_2204), .B(n_60558), .C(n_60536), .D(n_2264), .Z(n_300686326
		));
	notech_or4 i_157133166(.A(n_2044), .B(n_35829), .C(n_26592), .D(n_60586)
		, .Z(n_54865));
	notech_or4 i_16742(.A(n_58913), .B(n_1844), .C(n_59762), .D(n_60468), .Z
		(n_300786327));
	notech_or4 i_16743(.A(n_58913), .B(n_57404), .C(n_59201), .D(n_60468), .Z
		(n_300886328));
	notech_or4 i_16744(.A(n_58913), .B(n_57404), .C(n_58940), .D(n_60468), .Z
		(n_300986329));
	notech_or4 i_183833182(.A(n_60536), .B(n_59364), .C(n_2588), .D(n_60507)
		, .Z(n_57391));
	notech_or4 i_17709(.A(n_57338), .B(n_218285508), .C(n_26315), .D(n_2796)
		, .Z(n_301086330));
	notech_or4 i_17712(.A(n_106813462), .B(n_274588712), .C(n_57371), .D(n_60468
		), .Z(n_301186331));
	notech_or4 i_18359(.A(n_60762), .B(n_60719), .C(n_55280), .D(n_60584), .Z
		(n_301286332));
	notech_or4 i_19672(.A(n_106813462), .B(n_274588712), .C(n_60479), .D(n_60468
		), .Z(n_301386333));
	notech_or4 i_20678(.A(n_59364), .B(n_59958), .C(n_60602), .D(n_60468), .Z
		(n_301486334));
	notech_or4 i_21673(.A(n_60762), .B(n_60719), .C(n_57424), .D(n_60584), .Z
		(n_301586335));
	notech_or4 i_50333186(.A(calc_sz[3]), .B(calc_sz[2]), .C(n_260688757), .D
		(n_204988864), .Z(n_55846));
	notech_nand3 i_46970(.A(n_55745), .B(n_238685706), .C(n_238385703), .Z(\nbus_11281[0] 
		));
	notech_and2 i_116265717(.A(n_51738), .B(n_2236), .Z(n_55210));
	notech_or4 i_4557(.A(n_60762), .B(n_60721), .C(n_55210), .D(n_60584), .Z
		(n_52420));
	notech_nand2 i_408365686(.A(n_54877), .B(n_238285702), .Z(n_10177));
	notech_nao3 i_7224(.A(n_251385833), .B(n_224085563), .C(n_251485834), .Z
		(n_7435));
	notech_ao4 i_3215337(.A(n_237585695), .B(n_27984), .C(n_265085970), .D(n_27554
		), .Z(n_15173));
	notech_ao4 i_3115336(.A(n_237585695), .B(n_27983), .C(n_265085970), .D(n_27553
		), .Z(n_15168));
	notech_ao4 i_3015335(.A(n_237585695), .B(n_27982), .C(n_265085970), .D(n_27552
		), .Z(n_15163));
	notech_ao4 i_2915334(.A(n_237585695), .B(n_27981), .C(n_265085970), .D(n_27551
		), .Z(n_15158));
	notech_ao4 i_2815333(.A(n_237585695), .B(n_27980), .C(n_265085970), .D(n_27550
		), .Z(n_15153));
	notech_ao4 i_2715332(.A(n_237585695), .B(n_27979), .C(n_265085970), .D(n_27549
		), .Z(n_15148));
	notech_ao4 i_2615331(.A(n_237585695), .B(n_27978), .C(n_265085970), .D(n_27548
		), .Z(n_15143));
	notech_ao4 i_2515330(.A(n_27977), .B(n_237585695), .C(n_265085970), .D(n_27546
		), .Z(n_15138));
	notech_ao4 i_2415329(.A(n_237585695), .B(n_27976), .C(n_265085970), .D(n_27545
		), .Z(n_15133));
	notech_ao4 i_2315328(.A(n_237585695), .B(n_27975), .C(n_265085970), .D(n_27542
		), .Z(n_15128));
	notech_ao4 i_2215327(.A(n_237585695), .B(n_27974), .C(n_265085970), .D(n_27541
		), .Z(n_15123));
	notech_ao4 i_2115326(.A(n_237585695), .B(n_27973), .C(n_265085970), .D(n_27540
		), .Z(n_15118));
	notech_ao4 i_2015325(.A(n_237585695), .B(n_27972), .C(n_265085970), .D(n_27539
		), .Z(n_15113));
	notech_ao4 i_1915324(.A(n_237585695), .B(n_27971), .C(n_265085970), .D(n_27538
		), .Z(n_15108));
	notech_ao4 i_1815323(.A(n_237585695), .B(n_27970), .C(n_265085970), .D(n_27537
		), .Z(n_15103));
	notech_ao4 i_1715322(.A(n_237585695), .B(n_27969), .C(n_265085970), .D(n_27535
		), .Z(n_15098));
	notech_ao4 i_1615321(.A(n_53650), .B(n_27968), .C(n_53641), .D(n_27534),
		 .Z(n_15093));
	notech_ao4 i_1515320(.A(n_53650), .B(n_27967), .C(n_53641), .D(n_27533),
		 .Z(n_15088));
	notech_ao4 i_1415319(.A(n_53650), .B(n_27966), .C(n_53641), .D(n_27532),
		 .Z(n_15083));
	notech_ao4 i_1315318(.A(n_53650), .B(n_27965), .C(n_53641), .D(n_27531),
		 .Z(n_15078));
	notech_ao4 i_1215317(.A(n_53650), .B(n_27964), .C(n_53641), .D(n_27530),
		 .Z(n_15073));
	notech_ao4 i_1115316(.A(n_53650), .B(n_27963), .C(n_53641), .D(n_27529),
		 .Z(n_15068));
	notech_ao4 i_1015315(.A(n_53650), .B(n_27962), .C(n_53641), .D(n_27528),
		 .Z(n_15063));
	notech_ao4 i_915314(.A(n_53650), .B(n_27961), .C(n_53641), .D(n_27527), 
		.Z(n_15058));
	notech_ao4 i_815313(.A(n_53650), .B(n_27960), .C(n_53641), .D(n_27526), 
		.Z(n_15053));
	notech_ao4 i_715312(.A(n_53650), .B(n_27959), .C(n_53641), .D(n_27525), 
		.Z(n_15048));
	notech_ao4 i_615311(.A(n_53650), .B(n_27958), .C(n_265085970), .D(n_27524
		), .Z(n_15043));
	notech_ao4 i_515310(.A(n_53650), .B(n_27957), .C(n_53641), .D(n_27523), 
		.Z(n_15038));
	notech_ao4 i_415309(.A(n_53650), .B(n_27956), .C(n_53641), .D(n_27522), 
		.Z(n_15033));
	notech_ao4 i_315308(.A(n_53650), .B(n_27955), .C(n_53641), .D(n_27521), 
		.Z(n_15028));
	notech_ao4 i_215307(.A(n_53650), .B(n_27954), .C(n_53641), .D(n_27520), 
		.Z(n_15023));
	notech_ao4 i_115306(.A(n_53650), .B(n_27953), .C(n_53641), .D(n_27519), 
		.Z(n_15018));
	notech_nand2 i_6427416(.A(n_265285972), .B(n_230885630), .Z(n_18012));
	notech_nand2 i_6327415(.A(n_265385973), .B(n_230685628), .Z(n_18007));
	notech_nand2 i_6227414(.A(n_265485974), .B(n_230485626), .Z(n_18002));
	notech_nand2 i_6127413(.A(n_265585975), .B(n_230385625), .Z(n_17997));
	notech_nand2 i_6027412(.A(n_265685976), .B(n_230285624), .Z(n_17992));
	notech_nand2 i_5927411(.A(n_265785977), .B(n_230185623), .Z(n_17987));
	notech_nand2 i_5827410(.A(n_265885978), .B(n_230085622), .Z(n_17982));
	notech_nand2 i_5727409(.A(n_265985979), .B(n_229985621), .Z(n_17977));
	notech_nand2 i_5627408(.A(n_266085980), .B(n_229885620), .Z(n_17972));
	notech_nand2 i_5527407(.A(n_266185981), .B(n_229785619), .Z(n_17967));
	notech_nand2 i_5427406(.A(n_266285982), .B(n_229685618), .Z(n_17962));
	notech_nand2 i_5327405(.A(n_266385983), .B(n_229585617), .Z(n_17957));
	notech_nand2 i_5227404(.A(n_266485984), .B(n_229485616), .Z(n_17952));
	notech_nand2 i_5127403(.A(n_266585985), .B(n_229385615), .Z(n_17947));
	notech_nand2 i_5027402(.A(n_266685986), .B(n_229285614), .Z(n_17942));
	notech_nand2 i_4927401(.A(n_266785987), .B(n_229185613), .Z(n_17937));
	notech_nand2 i_4827400(.A(n_266885988), .B(n_229085612), .Z(n_17932));
	notech_nand2 i_4727399(.A(n_266985989), .B(n_228985611), .Z(n_17927));
	notech_nand2 i_4627398(.A(n_267085990), .B(n_228885610), .Z(n_17922));
	notech_nand2 i_4527397(.A(n_267185991), .B(n_228785609), .Z(n_17917));
	notech_nand2 i_4427396(.A(n_267285992), .B(n_228685608), .Z(n_17912));
	notech_nand2 i_4327395(.A(n_267385993), .B(n_228585607), .Z(n_17907));
	notech_nand2 i_4227394(.A(n_267485994), .B(n_228485606), .Z(n_17902));
	notech_nand2 i_4127393(.A(n_267585995), .B(n_228385605), .Z(n_17897));
	notech_nand2 i_4027392(.A(n_267685996), .B(n_228285604), .Z(n_17892));
	notech_nand2 i_3927391(.A(n_267785997), .B(n_228185603), .Z(n_17887));
	notech_nand2 i_3827390(.A(n_267885998), .B(n_228085602), .Z(n_17882));
	notech_nand2 i_3727389(.A(n_267985999), .B(n_227985601), .Z(n_17877));
	notech_nand2 i_3627388(.A(n_268086000), .B(n_227885600), .Z(n_17872));
	notech_nand2 i_3527387(.A(n_268186001), .B(n_227785599), .Z(n_17867));
	notech_nand2 i_3427386(.A(n_268286002), .B(n_227685598), .Z(n_17862));
	notech_nand2 i_3327385(.A(n_268386003), .B(n_227585597), .Z(n_17857));
	notech_nand2 i_3227384(.A(n_268486004), .B(n_227485596), .Z(n_17852));
	notech_nand2 i_3127383(.A(n_268586005), .B(n_227385595), .Z(n_17847));
	notech_nand2 i_3027382(.A(n_268686006), .B(n_227285594), .Z(n_17842));
	notech_nand2 i_2927381(.A(n_268786007), .B(n_227185593), .Z(n_17837));
	notech_nand2 i_2827380(.A(n_268886008), .B(n_227085592), .Z(n_17832));
	notech_nand2 i_2727379(.A(n_268986009), .B(n_226985591), .Z(n_17827));
	notech_nand2 i_2627378(.A(n_269086010), .B(n_226885590), .Z(n_17822));
	notech_nand2 i_2527377(.A(n_269186011), .B(n_226785589), .Z(n_17817));
	notech_nand2 i_2427376(.A(n_269286012), .B(n_226685588), .Z(n_17812));
	notech_nand2 i_2327375(.A(n_269386013), .B(n_226585587), .Z(n_17807));
	notech_nand2 i_2227374(.A(n_269486014), .B(n_226485586), .Z(n_17802));
	notech_nand2 i_2127373(.A(n_269586015), .B(n_226385585), .Z(n_17797));
	notech_nand2 i_2027372(.A(n_269686016), .B(n_226285584), .Z(n_17792));
	notech_nand2 i_1927371(.A(n_269786017), .B(n_226185583), .Z(n_17787));
	notech_nand2 i_1827370(.A(n_269886018), .B(n_225985582), .Z(n_17782));
	notech_nand2 i_1727369(.A(n_269986019), .B(n_225885581), .Z(n_17777));
	notech_nand2 i_1627368(.A(n_270086020), .B(n_225785580), .Z(n_17772));
	notech_nand2 i_1527367(.A(n_270186021), .B(n_225685579), .Z(n_17767));
	notech_nand2 i_1427366(.A(n_270286022), .B(n_225585578), .Z(n_17762));
	notech_nand2 i_1327365(.A(n_270386023), .B(n_225485577), .Z(n_17757));
	notech_nand2 i_1227364(.A(n_270486024), .B(n_225385576), .Z(n_17752));
	notech_nand2 i_1127363(.A(n_270586025), .B(n_225285575), .Z(n_17747));
	notech_nand2 i_1027362(.A(n_270686026), .B(n_225185574), .Z(n_17742));
	notech_nand2 i_927361(.A(n_270786027), .B(n_225085573), .Z(n_17737));
	notech_nand2 i_827360(.A(n_270886028), .B(n_224985572), .Z(n_17732));
	notech_nand2 i_727359(.A(n_270986029), .B(n_224885571), .Z(n_17727));
	notech_nand2 i_627358(.A(n_271086030), .B(n_224785570), .Z(n_17722));
	notech_nand2 i_527357(.A(n_271186031), .B(n_224685569), .Z(n_17717));
	notech_nand2 i_427356(.A(n_271286032), .B(n_224585568), .Z(n_17712));
	notech_nand2 i_327355(.A(n_271386033), .B(n_224485567), .Z(n_17707));
	notech_nand2 i_227354(.A(n_271486034), .B(n_224385566), .Z(n_17702));
	notech_nand2 i_127353(.A(n_271586035), .B(n_224285565), .Z(n_17697));
	notech_nand3 i_3218634(.A(n_271986039), .B(n_272186041), .C(n_247985799)
		, .Z(n_18411));
	notech_nand3 i_3118633(.A(n_272286042), .B(n_272486044), .C(n_247485794)
		, .Z(n_18406));
	notech_nand3 i_3018632(.A(n_272586045), .B(n_272786047), .C(n_246985789)
		, .Z(n_18401));
	notech_nand3 i_2918631(.A(n_272886048), .B(n_273086050), .C(n_246485784)
		, .Z(n_18396));
	notech_nand3 i_2818630(.A(n_273186051), .B(n_273386053), .C(n_245985779)
		, .Z(n_18391));
	notech_nand3 i_2718629(.A(n_273486054), .B(n_273686056), .C(n_245485774)
		, .Z(n_18386));
	notech_nand3 i_2618628(.A(n_273786057), .B(n_273986059), .C(n_244985769)
		, .Z(n_18381));
	notech_nand3 i_2518627(.A(n_274086060), .B(n_274286062), .C(n_244485764)
		, .Z(n_18376));
	notech_nand3 i_2418626(.A(n_274386063), .B(n_274586065), .C(n_243985759)
		, .Z(n_18371));
	notech_nand3 i_2318625(.A(n_274686066), .B(n_274886068), .C(n_243485754)
		, .Z(n_18366));
	notech_nand3 i_1618618(.A(n_274986069), .B(n_275186071), .C(n_242985749)
		, .Z(n_18331));
	notech_nand3 i_918611(.A(n_242485744), .B(n_275286072), .C(n_275486074),
		 .Z(n_18296));
	notech_nand3 i_718609(.A(n_275586075), .B(n_275786077), .C(n_241985739),
		 .Z(n_18286));
	notech_nand3 i_518607(.A(n_275886078), .B(n_276086080), .C(n_241485734),
		 .Z(n_18276));
	notech_nand3 i_418606(.A(n_276186081), .B(n_276386083), .C(n_240985729),
		 .Z(n_18271));
	notech_nand3 i_318605(.A(n_276486084), .B(n_276686086), .C(n_240485724),
		 .Z(n_18266));
	notech_nand3 i_218604(.A(n_276786087), .B(n_276986089), .C(n_239985719),
		 .Z(n_18261));
	notech_nand3 i_118603(.A(n_277086090), .B(n_277286092), .C(n_239485714),
		 .Z(n_18256));
	notech_ao4 i_222678(.A(n_59807), .B(n_26604), .C(n_223785560), .D(n_277586095
		), .Z(n_17661));
	notech_or4 i_133765673(.A(n_60540), .B(n_2386), .C(n_62419), .D(n_59907)
		, .Z(n_207041701));
	notech_nao3 i_50233187(.A(n_59183), .B(n_26592), .C(n_2044), .Z(n_55847)
		);
	notech_or2 i_50433188(.A(n_56569), .B(n_204988864), .Z(n_55845));
	notech_nao3 i_830599(.A(calc_sz[1]), .B(n_27402), .C(n_2605), .Z(n_56112
		));
	notech_or4 i_2123(.A(n_60540), .B(n_59762), .C(n_60602), .D(n_62419), .Z
		(n_57384));
	notech_or4 i_148733194(.A(n_59364), .B(n_60490), .C(n_59967), .D(n_59210
		), .Z(n_57423));
	notech_nand3 i_51137(.A(n_211288830), .B(n_2188), .C(n_212788817), .Z(\nbus_11321[0] 
		));
	notech_nand3 i_2165(.A(n_2340), .B(n_26663), .C(n_26785), .Z(n_57380));
	notech_or4 i_4135657(.A(opa[1]), .B(opa[0]), .C(opa[2]), .D(opa[3]), .Z(n_326046828
		));
	notech_nand2 i_3935659(.A(n_56649), .B(nbus_11273[0]), .Z(n_326246826)
		);
	notech_ao3 i_29600(.A(n_2385), .B(n_2361), .C(n_274588712), .Z(n_273088725
		));
	notech_nand3 i_1735671(.A(n_26284), .B(n_56685), .C(n_56694), .Z(n_327446814
		));
	notech_nand3 i_1335673(.A(n_26283), .B(n_56676), .C(n_56685), .Z(n_327646812
		));
	notech_nand2 i_103635687(.A(n_26283), .B(n_56676), .Z(n_3290));
	notech_nand2 i_194(.A(n_60507), .B(n_60536), .Z(n_272988726));
	notech_or4 i_3035667(.A(n_59201), .B(n_60490), .C(n_59967), .D(n_59958),
		 .Z(n_327046818));
	notech_or2 i_1193(.A(n_2773), .B(n_58904), .Z(n_272888727));
	notech_nand3 i_3635662(.A(n_26285), .B(n_56694), .C(n_57326), .Z(n_326546823
		));
	notech_nand3 i_87235709(.A(n_56649), .B(nbus_11273[0]), .C(n_56658), .Z(n_55482
		));
	notech_or4 i_166935762(.A(n_60762), .B(n_60724), .C(n_57380), .D(n_60586
		), .Z(n_54784));
	notech_nand2 i_93(.A(n_62429), .B(n_60536), .Z(n_272788728));
	notech_or4 i_29100(.A(n_60490), .B(n_59967), .C(n_60558), .D(n_59375), .Z
		(n_272688729));
	notech_or4 i_153335766(.A(n_59762), .B(n_60490), .C(n_59967), .D(n_59958
		), .Z(n_57418));
	notech_or2 i_174133161(.A(n_2213), .B(n_1931), .Z(n_54725));
	notech_or4 i_107833180(.A(n_60767), .B(n_60724), .C(n_272588730), .D(n_59201
		), .Z(n_55292));
	notech_or4 i_174933098(.A(n_60770), .B(n_60724), .C(n_192288896), .D(n_55400
		), .Z(n_54719));
	notech_or4 i_103732991(.A(n_58940), .B(n_60490), .C(n_60770), .D(n_60724
		), .Z(n_55332));
	notech_or4 i_8733(.A(n_59201), .B(n_60490), .C(n_60770), .D(n_60724), .Z
		(n_48510));
	notech_nao3 i_32099(.A(n_60536), .B(n_62403), .C(n_2588), .Z(n_272588730
		));
	notech_and3 i_53833014(.A(n_55693), .B(n_2006), .C(n_55687), .Z(n_55811)
		);
	notech_ao3 i_75333036(.A(n_55236), .B(n_55263), .C(n_1897), .Z(n_55597)
		);
	notech_and3 i_76333024(.A(n_55216), .B(n_1898), .C(n_55264), .Z(n_55587)
		);
	notech_nao3 i_230(.A(n_2578), .B(n_60507), .C(n_60536), .Z(n_106813462)
		);
	notech_ao4 i_121833121(.A(n_55958), .B(n_54505), .C(n_2177), .D(eval_flag
		), .Z(n_55156));
	notech_ao4 i_73133130(.A(n_2591), .B(n_56041), .C(n_2213), .D(n_59219), 
		.Z(n_55619));
	notech_ao4 i_99833131(.A(n_57388), .B(n_59907), .C(n_2210), .D(n_26296),
		 .Z(n_55366));
	notech_ao4 i_112933132(.A(mask8b[2]), .B(n_1907), .C(n_222456215), .D(n_220856212
		), .Z(n_55243));
	notech_nand3 i_496(.A(n_59186), .B(n_59895), .C(n_59780), .Z(n_170914103
		));
	notech_or2 i_32071(.A(n_190688899), .B(instrc[107]), .Z(n_2320));
	notech_or4 i_32061(.A(n_58913), .B(n_59967), .C(n_59355), .D(n_55149), .Z
		(n_2323));
	notech_or4 i_32068(.A(n_58913), .B(n_2572), .C(n_2192), .D(n_59895), .Z(n_2322
		));
	notech_nand2 i_218060(.A(n_279486114), .B(n_279386113), .Z(write_data_28
		[1]));
	notech_nand2 i_3218346(.A(n_279686116), .B(n_279586115), .Z(write_data_30
		[31]));
	notech_ao4 i_7434(.A(n_60584), .B(n_59895), .C(n_277886098), .D(n_1910),
		 .Z(n_18925));
	notech_nao3 i_21603(.A(n_253034156), .B(n_273088725), .C(n_59355), .Z(n_35657
		));
	notech_nand2 i_126971(.A(n_58496), .B(n_281886138), .Z(n_9296));
	notech_or4 i_163732831(.A(n_60748), .B(n_60735), .C(n_60770), .D(n_192188897
		), .Z(n_2164));
	notech_or2 i_82732994(.A(n_2213), .B(n_56265), .Z(n_55526));
	notech_or4 i_32077(.A(n_58913), .B(n_59967), .C(n_59355), .D(n_1967), .Z
		(n_2319));
	notech_nand2 i_176132823(.A(n_2219), .B(n_274788710), .Z(n_2156));
	notech_nand2 i_2417826(.A(n_294886268), .B(n_294786267), .Z(write_data_26
		[23]));
	notech_nand2 i_2617828(.A(n_295086270), .B(n_294986269), .Z(write_data_26
		[25]));
	notech_nand2 i_2717829(.A(n_295286272), .B(n_295186271), .Z(write_data_26
		[26]));
	notech_nand2 i_2817830(.A(n_295486274), .B(n_295386273), .Z(write_data_26
		[27]));
	notech_nand2 i_2917831(.A(n_295686276), .B(n_295586275), .Z(write_data_26
		[28]));
	notech_nand2 i_1917821(.A(n_297886298), .B(n_297786297), .Z(write_data_26
		[18]));
	notech_nand2 i_2017822(.A(n_298086300), .B(n_297986299), .Z(write_data_26
		[19]));
	notech_nand2 i_2117823(.A(n_298286302), .B(n_298186301), .Z(write_data_26
		[20]));
	notech_nand2 i_2217824(.A(n_298486304), .B(n_298386303), .Z(write_data_26
		[21]));
	notech_nand2 i_2317825(.A(n_298686306), .B(n_298586305), .Z(write_data_26
		[22]));
	notech_nand3 i_55131(.A(n_300186321), .B(n_55745), .C(n_300286322), .Z(\nbus_11356[0] 
		));
	notech_nand2 i_52889(.A(n_300186321), .B(n_55625), .Z(n_17679));
	notech_or4 i_154932988(.A(n_59364), .B(n_60490), .C(n_57404), .D(n_59895
		), .Z(n_54884));
	notech_or4 i_172932989(.A(n_58940), .B(n_60494), .C(n_57404), .D(n_59895
		), .Z(n_54735));
	notech_or2 i_29977(.A(n_2255), .B(n_55958), .Z(n_2326));
	notech_nand2 i_114432860(.A(n_59780), .B(n_59895), .Z(n_2193));
	notech_or4 i_97232878(.A(n_56460), .B(n_55522), .C(n_1962), .D(n_56440),
		 .Z(n_2211));
	notech_or4 i_97132879(.A(n_55522), .B(n_2349), .C(n_55833), .D(n_60507),
		 .Z(n_2212));
	notech_nao3 i_25532917(.A(n_2578), .B(n_62419), .C(n_60536), .Z(n_2253)
		);
	notech_nand2 i_8539008(.A(read_data[17]), .B(n_59895), .Z(n_272488731)
		);
	notech_nand2 i_4039052(.A(n_55292), .B(n_272288733), .Z(n_272388732));
	notech_or4 i_110632865(.A(n_60768), .B(n_60724), .C(n_59762), .D(n_60494
		), .Z(n_2198));
	notech_or4 i_177539075(.A(n_59762), .B(n_60494), .C(n_59895), .D(n_106813462
		), .Z(n_89713291));
	notech_or4 i_165039076(.A(n_60768), .B(n_60724), .C(n_59762), .D(n_272588730
		), .Z(n_89513289));
	notech_ao4 i_116639078(.A(n_272888727), .B(n_59895), .C(n_2253), .D(n_1602
		), .Z(n_272288733));
	notech_or4 i_42839083(.A(calc_sz[3]), .B(calc_sz[0]), .C(n_260888755), .D
		(n_2318), .Z(n_88913283));
	notech_or4 i_32104(.A(n_59369), .B(n_60494), .C(n_274488713), .D(n_59895
		), .Z(n_2318));
	notech_or2 i_830596(.A(n_260988754), .B(n_260888755), .Z(n_56099));
	notech_nand3 i_42739084(.A(n_1969), .B(n_57438), .C(n_59807), .Z(n_88813282
		));
	notech_and4 i_143739090(.A(n_1780), .B(n_1779), .C(n_177588906), .D(n_1778
		), .Z(n_272188734));
	notech_and4 i_143939091(.A(n_175688923), .B(n_175588924), .C(n_1751), .D
		(n_1754), .Z(n_272088735));
	notech_and4 i_92729151(.A(n_171088929), .B(n_170988930), .C(n_170588934)
		, .D(n_170888931), .Z(n_271988736));
	notech_and4 i_92529149(.A(n_169688943), .B(n_169588944), .C(n_169188948)
		, .D(n_169488945), .Z(n_271888737));
	notech_or4 i_37039117(.A(n_60586), .B(n_59895), .C(n_1900), .D(n_26326),
		 .Z(n_55979));
	notech_or4 i_37139118(.A(n_60770), .B(n_60724), .C(n_54761), .D(n_60586)
		, .Z(n_55978));
	notech_mux2 i_1711674(.S(n_60138), .A(regs_14[16]), .B(add_len_pc32[16])
		, .Z(n_271788738));
	notech_or4 i_32739157(.A(n_60768), .B(n_60724), .C(n_54688), .D(n_60586)
		, .Z(n_56022));
	notech_nand3 i_8483(.A(opz[2]), .B(n_27517), .C(n_27518), .Z(n_48760));
	notech_nand2 i_117139161(.A(n_48760), .B(n_1562), .Z(n_57432));
	notech_or4 i_85942282(.A(n_1916), .B(n_1023), .C(n_60525), .D(n_1526), .Z
		(n_55495));
	notech_or2 i_85842284(.A(n_1526), .B(n_54527), .Z(n_55496));
	notech_nor2 i_3845339(.A(n_26443), .B(n_54151), .Z(n_303321920));
	notech_or2 i_5845319(.A(n_56063), .B(n_60586), .Z(n_301321900));
	notech_nand2 i_109345399(.A(n_56053), .B(n_301321900), .Z(n_55279));
	notech_nao3 i_155845400(.A(n_26592), .B(n_59186), .C(n_56502), .Z(n_54876
		));
	notech_nand2 i_242445406(.A(n_56053), .B(n_56052), .Z(n_54151));
	notech_or2 i_29645418(.A(n_55858), .B(n_60586), .Z(n_56053));
	notech_or4 i_158845422(.A(n_260688757), .B(n_2605), .C(n_56498), .D(n_60586
		), .Z(n_54851));
	notech_or2 i_153045425(.A(n_56058), .B(n_60586), .Z(n_54900));
	notech_or2 i_29745419(.A(n_55827), .B(n_60586), .Z(n_56052));
	notech_nor2 i_129145427(.A(n_55279), .B(n_26555), .Z(n_55088));
	notech_nand2 i_25491(.A(n_59186), .B(n_59894), .Z(n_123723224));
	notech_and2 i_105645407(.A(n_55978), .B(n_1491), .Z(n_55314));
	notech_ao4 i_105745408(.A(n_26326), .B(n_54874), .C(n_1492), .D(n_320788482
		), .Z(n_55313));
	notech_nao3 i_178733000(.A(n_55040), .B(n_59807), .C(n_59762), .Z(n_54687
		));
	notech_nao3 i_152933111(.A(n_55040), .B(n_59807), .C(n_59201), .Z(n_54901
		));
	notech_or4 i_930842(.A(instrc[123]), .B(instrc[121]), .C(n_28566), .D(n_60525
		), .Z(n_193714331));
	notech_or4 i_930751(.A(n_60549), .B(instrc[121]), .C(instrc[120]), .D(n_60525
		), .Z(n_165623643));
	notech_or4 i_4845329(.A(n_56460), .B(n_56469), .C(n_55522), .D(n_1492), 
		.Z(n_302321910));
	notech_or4 i_4345334(.A(n_59299), .B(n_59290), .C(n_55088), .D(n_59250),
		 .Z(n_302821915));
	notech_ao4 i_81339135(.A(n_60468), .B(n_55325), .C(n_317888511), .D(n_316888521
		), .Z(n_271688739));
	notech_ao4 i_81439136(.A(n_54688), .B(n_60468), .C(n_316888521), .D(n_320788482
		), .Z(n_271588740));
	notech_or4 i_140232847(.A(n_60540), .B(n_60507), .C(n_60563), .D(\opcode[1] 
		), .Z(n_2180));
	notech_or4 i_7633056(.A(n_60549), .B(n_59241), .C(n_28566), .D(n_59230),
		 .Z(n_56189));
	notech_or4 i_7733025(.A(n_60549), .B(n_59241), .C(instrc[120]), .D(n_59230
		), .Z(n_56188));
	notech_nao3 i_7933026(.A(instrc[121]), .B(n_59230), .C(n_1909), .Z(n_56186
		));
	notech_or2 i_8333029(.A(n_1913), .B(n_60525), .Z(n_56182));
	notech_or4 i_8533031(.A(n_60549), .B(instrc[121]), .C(instrc[120]), .D(n_59230
		), .Z(n_56180));
	notech_or4 i_8633032(.A(n_60549), .B(n_59241), .C(n_28566), .D(n_60527),
		 .Z(n_56179));
	notech_or2 i_8733033(.A(n_1916), .B(n_59235), .Z(n_56178));
	notech_nao3 i_8932926(.A(n_60527), .B(instrc[121]), .C(n_1909), .Z(n_2262
		));
	notech_or4 i_9033034(.A(n_60549), .B(n_60516), .C(n_28566), .D(n_59230),
		 .Z(n_56175));
	notech_or2 i_9132925(.A(n_1913), .B(n_59230), .Z(n_2261));
	notech_and2 i_187049160(.A(opc[1]), .B(n_59113), .Z(n_110723094));
	notech_or4 i_135549164(.A(n_56487), .B(n_56478), .C(n_2349), .D(n_1301),
		 .Z(n_123623223));
	notech_nao3 i_130449166(.A(n_62429), .B(n_26305), .C(n_263436789), .Z(n_123423221
		));
	notech_or4 i_103849172(.A(rep_en3), .B(rep_en2), .C(rep_en1), .D(n_26890
		), .Z(n_271488741));
	notech_nao3 i_77949176(.A(rep_en3), .B(n_26889), .C(rep_en2), .Z(n_271388742
		));
	notech_or4 i_39949186(.A(n_59263), .B(n_59272), .C(n_56177), .D(n_55798)
		, .Z(n_123223219));
	notech_nand2 i_24949189(.A(nbus_11326[0]), .B(nbus_11326[1]), .Z(n_149823485
		));
	notech_nand2 i_3149192(.A(opc_10[29]), .B(n_62405), .Z(n_110923096));
	notech_and4 i_145449194(.A(n_1443), .B(n_1442), .C(n_1438), .D(n_1441), 
		.Z(n_271288743));
	notech_and4 i_145349195(.A(n_145756185), .B(n_145656184), .C(n_145256180
		), .D(n_145556183), .Z(n_271188744));
	notech_and4 i_94229164(.A(n_1413), .B(n_1412), .C(n_1408), .D(n_1411), .Z
		(n_271088745));
	notech_and4 i_94149196(.A(n_1399), .B(n_1398), .C(n_1394), .D(n_1397), .Z
		(n_270988746));
	notech_nand3 i_29627(.A(opc[1]), .B(n_59113), .C(opc[2]), .Z(n_2708));
	notech_and4 i_145249211(.A(n_1428), .B(n_1427), .C(n_1423), .D(n_1426), 
		.Z(n_270688747));
	notech_or4 i_169049219(.A(rep_en3), .B(rep_en2), .C(rep_en1), .D(rep_en4
		), .Z(n_270588748));
	notech_nand2 i_164549220(.A(rep_en2), .B(n_26889), .Z(n_270488749));
	notech_ao3 i_112849225(.A(nbus_11326[0]), .B(nbus_11326[1]), .C(n_2770),
		 .Z(n_270388750));
	notech_nand3 i_1989(.A(n_56569), .B(n_56560), .C(n_56547), .Z(n_54520)
		);
	notech_and2 i_95749236(.A(n_55497), .B(n_54454), .Z(n_2702));
	notech_ao4 i_95649237(.A(n_26591), .B(n_29012), .C(n_318931576), .D(n_26277
		), .Z(n_2701));
	notech_and2 i_20306(.A(n_55827), .B(n_56063), .Z(n_36952));
	notech_and2 i_107232870(.A(n_26782), .B(n_59807), .Z(n_2203));
	notech_and4 i_67439079(.A(n_272488731), .B(n_174288925), .C(n_1600), .D(n_1597
		), .Z(n_43426147));
	notech_nand3 i_53033113(.A(n_205988854), .B(n_2215), .C(n_221888805), .Z
		(n_55819));
	notech_and4 i_91835755(.A(n_1874), .B(n_1873), .C(n_1869), .D(n_1872), .Z
		(n_57351));
	notech_ao4 i_93742285(.A(n_58895), .B(n_1041), .C(n_1529), .D(n_55995), 
		.Z(n_55424));
	notech_and2 i_95842283(.A(n_55496), .B(n_54459), .Z(n_55405));
	notech_and2 i_95942281(.A(n_55495), .B(n_54441), .Z(n_55404));
	notech_or4 i_36849188(.A(n_60770), .B(n_60724), .C(n_2180), .D(n_60602),
		 .Z(n_107626780));
	notech_or4 i_78233035(.A(n_55087), .B(n_1955), .C(n_55833), .D(n_59241),
		 .Z(n_55568));
	notech_or2 i_78333039(.A(n_55833), .B(n_190588900), .Z(n_55567));
	notech_or4 i_132142239(.A(n_56487), .B(n_56478), .C(n_56449), .D(n_1527)
		, .Z(n_308418861));
	notech_or4 i_40442251(.A(n_59263), .B(n_59272), .C(n_56196), .D(n_55798)
		, .Z(n_309618873));
	notech_or4 i_63042274(.A(n_59263), .B(n_59268), .C(n_56196), .D(n_56369)
		, .Z(n_55720));
	notech_and4 i_92829152(.A(n_1739), .B(n_1738), .C(n_1734), .D(n_1737), .Z
		(n_2700));
	notech_and4 i_91139147(.A(n_1725), .B(n_1724), .C(n_1720), .D(n_1723), .Z
		(n_2699));
	notech_or4 i_42933067(.A(n_60770), .B(n_60724), .C(n_56569), .D(n_1900),
		 .Z(n_55920));
	notech_or4 i_66333061(.A(n_56573), .B(n_56354), .C(n_56177), .D(n_59250)
		, .Z(n_55687));
	notech_or4 i_115633175(.A(n_55087), .B(n_1955), .C(n_205188862), .D(n_59241
		), .Z(n_55216));
	notech_or2 i_113633176(.A(n_205188862), .B(n_190588900), .Z(n_55236));
	notech_or4 i_54133013(.A(n_58945), .B(n_205588858), .C(n_60586), .D(n_59894
		), .Z(n_55808));
	notech_nand3 i_25798(.A(n_26625), .B(n_59780), .C(n_26554), .Z(n_2345)
		);
	notech_ao4 i_51533038(.A(n_204988864), .B(n_56547), .C(n_56345), .D(n_26228
		), .Z(n_55834));
	notech_ao4 i_51633181(.A(n_56059), .B(n_60586), .C(n_2250), .D(n_26228),
		 .Z(n_55833));
	notech_ao4 i_50733112(.A(n_2005), .B(n_59369), .C(n_2250), .D(n_55934), 
		.Z(n_55842));
	notech_or4 i_930845(.A(n_60549), .B(n_59241), .C(instrc[120]), .D(n_60527
		), .Z(n_197114365));
	notech_nand2 i_432927(.A(n_62429), .B(n_59375), .Z(n_2263));
	notech_nand2 i_132928(.A(n_62429), .B(\opcode[1] ), .Z(n_2264));
	notech_nao3 i_48332907(.A(n_59299), .B(n_58645), .C(n_59290), .Z(n_2242)
		);
	notech_nao3 i_47133057(.A(n_59259), .B(n_59268), .C(n_59277), .Z(n_55878
		));
	notech_nand3 i_47633015(.A(n_59299), .B(n_59290), .C(n_58645), .Z(n_55873
		));
	notech_nao3 i_47733016(.A(n_59299), .B(n_59290), .C(n_56158), .Z(n_55872
		));
	notech_or2 i_47833017(.A(n_56158), .B(n_56114), .Z(n_55871));
	notech_nao3 i_47933018(.A(n_59299), .B(n_59290), .C(n_56081), .Z(n_55870
		));
	notech_or4 i_48033019(.A(n_59259), .B(n_59268), .C(n_59299), .D(n_59290)
		, .Z(n_55869));
	notech_or2 i_48133020(.A(n_56177), .B(n_56074), .Z(n_55868));
	notech_or2 i_48433022(.A(n_56074), .B(n_59277), .Z(n_55865));
	notech_or2 i_48533023(.A(n_56158), .B(n_59277), .Z(n_55864));
	notech_or2 i_1970(.A(n_58660), .B(n_59281), .Z(n_54535));
	notech_nao3 i_2057(.A(n_59259), .B(n_59272), .C(n_56114), .Z(n_54465));
	notech_nand2 i_13187(.A(read_data[0]), .B(n_59894), .Z(n_2698));
	notech_or2 i_196951964(.A(n_1104), .B(n_2689), .Z(n_2697));
	notech_or4 i_130051970(.A(n_56460), .B(n_56431), .C(n_1085), .D(n_56440)
		, .Z(n_2694));
	notech_ao4 i_127351971(.A(n_55356), .B(n_55854), .C(n_1135), .D(n_28986)
		, .Z(n_2693));
	notech_ao3 i_25632916(.A(n_56487), .B(instrc[118]), .C(n_2349), .Z(n_2252
		));
	notech_nao3 i_97851977(.A(n_55567), .B(n_55263), .C(n_1897), .Z(n_2692)
		);
	notech_and3 i_97751978(.A(n_55568), .B(n_1898), .C(n_55264), .Z(n_2691)
		);
	notech_and3 i_61351986(.A(n_2006), .B(n_55842), .C(n_55693), .Z(n_2690)
		);
	notech_or2 i_24151994(.A(n_56460), .B(n_1189), .Z(n_2689));
	notech_nand2 i_1751996(.A(opc_10[17]), .B(n_62405), .Z(n_63826342));
	notech_and4 i_142351998(.A(n_1234), .B(n_1233), .C(n_1229), .D(n_1232), 
		.Z(n_2688));
	notech_or4 i_31960(.A(n_59299), .B(n_59290), .C(n_56074), .D(n_54089), .Z
		(n_2687));
	notech_or4 i_28433011(.A(n_60540), .B(n_56573), .C(n_59894), .D(n_2007),
		 .Z(n_56065));
	notech_or2 i_48233021(.A(n_56074), .B(n_56114), .Z(n_55867));
	notech_or4 i_31952(.A(n_59299), .B(n_59290), .C(n_56081), .D(n_55827), .Z
		(n_2686));
	notech_or2 i_188452007(.A(n_2660), .B(n_2689), .Z(n_54606));
	notech_ao4 i_32252010(.A(n_56498), .B(n_56560), .C(n_55807), .D(n_26227)
		, .Z(n_56027));
	notech_or4 i_27838(.A(n_56460), .B(n_56431), .C(n_56440), .D(n_2683), .Z
		(n_2685));
	notech_or4 i_27837(.A(n_56460), .B(n_56431), .C(n_2664), .D(n_56440), .Z
		(n_2684));
	notech_or2 i_205252019(.A(n_2683), .B(n_2650), .Z(n_54468));
	notech_and2 i_34551991(.A(n_56058), .B(n_1071), .Z(n_2683));
	notech_or4 i_210252020(.A(n_55087), .B(n_1069), .C(n_2683), .D(n_60516),
		 .Z(n_54428));
	notech_nao3 i_8433030(.A(n_60527), .B(n_59241), .C(n_1909), .Z(n_56181)
		);
	notech_nand2 i_25689(.A(n_56469), .B(n_28966), .Z(n_2349));
	notech_or2 i_22652026(.A(n_2349), .B(n_56431), .Z(n_56101));
	notech_nand2 i_26743(.A(opc[7]), .B(n_62405), .Z(n_2680));
	notech_nao3 i_327963(.A(n_2488), .B(n_2228), .C(n_224656217), .Z(opcode_289113
		));
	notech_nand2 i_26741(.A(opc_10[7]), .B(n_62405), .Z(n_2679));
	notech_or4 i_12998(.A(n_55087), .B(n_1069), .C(n_1188), .D(n_60516), .Z(n_2678
		));
	notech_or2 i_12999(.A(n_2650), .B(n_1188), .Z(n_2677));
	notech_or4 i_65733185(.A(n_56354), .B(n_56177), .C(n_56547), .D(n_59250)
		, .Z(n_55693));
	notech_or4 i_110833178(.A(n_55087), .B(n_1955), .C(n_55834), .D(n_28567)
		, .Z(n_55264));
	notech_or2 i_110933177(.A(n_55834), .B(n_190588900), .Z(n_55263));
	notech_mux2 i_811665(.S(n_60125), .A(n_563), .B(add_len_pc32[7]), .Z(n_2676
		));
	notech_and4 i_143052029(.A(n_1206), .B(n_1205), .C(n_1201), .D(n_1204), 
		.Z(n_2675));
	notech_and2 i_218249261(.A(n_55858), .B(n_36952), .Z(n_54367));
	notech_or2 i_2080(.A(n_56172), .B(n_56163), .Z(n_54446));
	notech_or2 i_27663(.A(n_55798), .B(n_56144), .Z(n_2674));
	notech_ao4 i_35151990(.A(n_56498), .B(n_56538), .C(n_56369), .D(n_26574)
		, .Z(n_2673));
	notech_or4 i_27648(.A(n_2349), .B(n_56431), .C(n_2673), .D(n_60507), .Z(n_2672
		));
	notech_or2 i_63352021(.A(n_56369), .B(n_56144), .Z(n_55717));
	notech_and2 i_59452037(.A(n_55717), .B(n_1084), .Z(n_2671));
	notech_or2 i_131152025(.A(n_2673), .B(n_2650), .Z(n_55068));
	notech_nand3 i_182152038(.A(n_2653), .B(n_55068), .C(n_2677), .Z(n_2670)
		);
	notech_or4 i_131052023(.A(n_55087), .B(n_1069), .C(n_2673), .D(n_60516),
		 .Z(n_55069));
	notech_and3 i_182352039(.A(n_2678), .B(n_2656), .C(n_55069), .Z(n_2669)
		);
	notech_and2 i_183452047(.A(n_55920), .B(n_2661), .Z(n_2668));
	notech_ao4 i_183552048(.A(n_2660), .B(n_2658), .C(n_1135), .D(n_59894), 
		.Z(n_2667));
	notech_and4 i_186552049(.A(n_2657), .B(n_2662), .C(n_55810), .D(n_1083),
		 .Z(n_2666));
	notech_and4 i_186752050(.A(n_61624), .B(n_56045), .C(n_2663), .D(n_1082)
		, .Z(n_2665));
	notech_and2 i_34249206(.A(n_54637), .B(n_54754), .Z(n_61624));
	notech_and4 i_252152055(.A(n_2673), .B(n_1188), .C(n_55667), .D(n_1073),
		 .Z(n_2664));
	notech_or4 i_209552059(.A(n_2740), .B(n_1076), .C(n_56025), .D(n_60527),
		 .Z(n_2663));
	notech_ao4 i_32452009(.A(n_56502), .B(n_56547), .C(n_55858), .D(n_26227)
		, .Z(n_56025));
	notech_or2 i_204452060(.A(n_56025), .B(n_2658), .Z(n_2662));
	notech_or4 i_178252061(.A(n_2740), .B(n_1076), .C(n_2660), .D(n_60527), 
		.Z(n_2661));
	notech_ao4 i_31852058(.A(n_56573), .B(n_56498), .C(n_55827), .D(n_26227)
		, .Z(n_2660));
	notech_or2 i_174052062(.A(n_2660), .B(n_2658), .Z(n_2659));
	notech_and3 i_148652046(.A(n_56260), .B(n_1077), .C(n_1075), .Z(n_2658)
		);
	notech_or2 i_124452068(.A(n_2658), .B(n_56029), .Z(n_2657));
	notech_or4 i_205652027(.A(n_55087), .B(n_1069), .C(n_55986), .D(n_60516)
		, .Z(n_2656));
	notech_and2 i_96552076(.A(n_2656), .B(n_2654), .Z(n_2655));
	notech_or4 i_86552077(.A(n_1069), .B(n_2651), .C(n_60516), .D(n_55087), 
		.Z(n_2654));
	notech_or2 i_205552028(.A(n_2650), .B(n_55986), .Z(n_2653));
	notech_nand2 i_96452078(.A(n_2653), .B(n_2649), .Z(n_2652));
	notech_and3 i_90651979(.A(n_56058), .B(n_1071), .C(n_1188), .Z(n_2651)
		);
	notech_and3 i_198452036(.A(n_56260), .B(n_1070), .C(n_1068), .Z(n_2650)
		);
	notech_or2 i_86452079(.A(n_2651), .B(n_2650), .Z(n_2649));
	notech_or4 i_156033165(.A(n_60770), .B(n_60724), .C(n_60583), .D(n_1900)
		, .Z(n_54874));
	notech_ao4 i_32052093(.A(n_56498), .B(n_56538), .C(n_56369), .D(n_26227)
		, .Z(n_56029));
	notech_and4 i_144052095(.A(n_1184), .B(n_1183), .C(n_1179), .D(n_1182), 
		.Z(n_2648));
	notech_ao3 i_5372(.A(n_60527), .B(instrc[107]), .C(n_1912), .Z(n_51741)
		);
	notech_nand3 i_1569(.A(n_2340), .B(n_26663), .C(n_2578), .Z(n_2647));
	notech_or4 i_31430(.A(n_273288723), .B(n_60602), .C(n_62395), .D(\opcode[1] 
		), .Z(n_323631623));
	notech_nao3 i_85755350(.A(n_318931576), .B(n_26320), .C(n_997), .Z(n_55497
		));
	notech_nand3 i_055294(.A(n_55658), .B(n_996), .C(n_56006), .Z(n_318931576
		));
	notech_or4 i_44855362(.A(n_60748), .B(n_60735), .C(n_60770), .D(n_1031),
		 .Z(n_55901));
	notech_or2 i_175033097(.A(n_55960), .B(n_54505), .Z(n_54718));
	notech_ao4 i_39033003(.A(n_56498), .B(n_56560), .C(n_55807), .D(n_26242)
		, .Z(n_55959));
	notech_nand2 i_21430(.A(n_56573), .B(n_56560), .Z(n_35829));
	notech_or2 i_146733169(.A(n_26570), .B(n_55836), .Z(n_54953));
	notech_or2 i_8233028(.A(n_1916), .B(n_60527), .Z(n_56183));
	notech_nao3 i_2088(.A(n_59299), .B(n_59290), .C(n_58656), .Z(n_54439));
	notech_or2 i_133857862(.A(n_2255), .B(n_1019), .Z(n_248534111));
	notech_or2 i_175833160(.A(n_55960), .B(n_54530), .Z(n_54711));
	notech_or4 i_22233044(.A(calc_sz[3]), .B(calc_sz[2]), .C(calc_sz[1]), .D
		(n_27402), .Z(n_56104));
	notech_nand2 i_77657878(.A(n_56560), .B(n_56547), .Z(n_250134127));
	notech_and2 i_82933009(.A(n_57374), .B(n_1900), .Z(n_55524));
	notech_or4 i_50833170(.A(n_58931), .B(n_59369), .C(n_60770), .D(n_60724)
		, .Z(n_55841));
	notech_or4 i_28235748(.A(n_1895), .B(n_1892), .C(n_1888), .D(n_1885), .Z
		(n_56067));
	notech_nor2 i_112735751(.A(n_1845), .B(n_326546823), .Z(n_55245));
	notech_nand2 i_211(.A(n_62395), .B(n_59375), .Z(n_2646));
	notech_ao4 i_36057901(.A(n_56498), .B(n_56560), .C(n_55807), .D(n_26805)
		, .Z(n_252434150));
	notech_or4 i_29233066(.A(n_60748), .B(n_60735), .C(n_60770), .D(n_54688)
		, .Z(n_56057));
	notech_and2 i_30457929(.A(n_56216), .B(n_1020), .Z(n_56045));
	notech_nand2 i_27357(.A(n_1016), .B(n_59807), .Z(n_254834174));
	notech_or4 i_28533041(.A(n_60540), .B(n_2007), .C(n_59895), .D(n_56538),
		 .Z(n_56064));
	notech_and2 i_249957941(.A(n_55580), .B(n_56369), .Z(n_54089));
	notech_or4 i_208657942(.A(n_1916), .B(n_1023), .C(n_55983), .D(n_60527),
		 .Z(n_54441));
	notech_ao4 i_36657922(.A(n_56498), .B(n_56547), .C(n_55858), .D(n_26805)
		, .Z(n_55983));
	notech_or2 i_206457945(.A(n_55983), .B(n_54527), .Z(n_54459));
	notech_or2 i_174557954(.A(n_54505), .B(n_55961), .Z(n_54722));
	notech_or4 i_157757955(.A(n_60770), .B(n_60721), .C(n_1031), .D(n_60583)
		, .Z(n_54860));
	notech_and2 i_1976(.A(n_56260), .B(n_2199), .Z(n_54530));
	notech_ao4 i_38833004(.A(n_56573), .B(n_56498), .C(n_55820), .D(n_26242)
		, .Z(n_55961));
	notech_or4 i_131757961(.A(n_1916), .B(n_1023), .C(n_55995), .D(n_60527),
		 .Z(n_55062));
	notech_and2 i_198057947(.A(n_1048), .B(n_56260), .Z(n_54527));
	notech_or2 i_131557962(.A(n_54527), .B(n_55995), .Z(n_55064));
	notech_and4 i_52833183(.A(n_56569), .B(n_56560), .C(n_56547), .D(n_54953
		), .Z(n_55821));
	notech_or4 i_110457966(.A(n_1046), .B(n_1035), .C(n_26191), .D(n_55821),
		 .Z(n_55268));
	notech_and3 i_106057969(.A(n_54718), .B(n_54722), .C(n_1044), .Z(n_55310
		));
	notech_ao3 i_51333171(.A(n_26887), .B(n_59807), .C(n_57378), .Z(n_55836)
		);
	notech_or2 i_169833163(.A(n_54530), .B(n_55958), .Z(n_54760));
	notech_ao3 i_101057971(.A(n_1039), .B(n_54760), .C(n_55831), .Z(n_55354)
		);
	notech_or4 i_28633010(.A(n_60540), .B(n_2007), .C(n_59895), .D(n_56560),
		 .Z(n_56063));
	notech_or4 i_28733012(.A(n_60540), .B(n_2007), .C(n_59895), .D(n_56551),
		 .Z(n_56062));
	notech_and2 i_77057975(.A(n_55807), .B(n_55858), .Z(n_55580));
	notech_or2 i_66557977(.A(n_55820), .B(n_55947), .Z(n_55685));
	notech_and3 i_62357978(.A(n_55685), .B(n_55776), .C(n_1040), .Z(n_55727)
		);
	notech_or2 i_57357986(.A(n_56369), .B(n_55952), .Z(n_55776));
	notech_nand2 i_53957988(.A(n_56056), .B(n_59807), .Z(n_55810));
	notech_nor2 i_101257970(.A(n_55836), .B(n_1027), .Z(n_55353));
	notech_nor2 i_51857989(.A(n_55353), .B(n_56551), .Z(n_55831));
	notech_nao3 i_178533008(.A(n_26599), .B(n_56551), .C(n_55524), .Z(n_54688
		));
	notech_and2 i_49557990(.A(n_54688), .B(n_1017), .Z(n_55854));
	notech_or2 i_254(.A(n_58913), .B(n_2825), .Z(n_2645));
	notech_or4 i_44657991(.A(n_60770), .B(n_60721), .C(n_59369), .D(n_58895)
		, .Z(n_55903));
	notech_or4 i_46316(.A(fsm[4]), .B(fsm[1]), .C(n_60721), .D(fsm[2]), .Z(n_159623583
		));
	notech_ao4 i_35457993(.A(n_56498), .B(n_56538), .C(n_56369), .D(n_26805)
		, .Z(n_55995));
	notech_ao4 i_34857995(.A(n_56569), .B(n_56502), .C(n_55820), .D(n_26805)
		, .Z(n_56001));
	notech_ao4 i_29357996(.A(n_26406), .B(n_26503), .C(n_26326), .D(n_250134127
		), .Z(n_56056));
	notech_or4 i_6730348(.A(n_327446814), .B(n_1845), .C(n_56067), .D(opa[7]
		), .Z(n_57433));
	notech_nao3 i_8033027(.A(n_60549), .B(n_28566), .C(n_2202), .Z(n_56185)
		);
	notech_or2 i_2074(.A(n_56172), .B(n_58656), .Z(n_54451));
	notech_or4 i_30749265(.A(n_60748), .B(n_60735), .C(n_60770), .D(n_54761)
		, .Z(n_101413408));
	notech_and4 i_94029163(.A(n_1523), .B(n_1522), .C(n_1518), .D(n_1521), .Z
		(n_57329));
	notech_or4 i_30349266(.A(n_60767), .B(n_60721), .C(n_1900), .D(n_26326),
		 .Z(n_101213406));
	notech_or4 i_29449267(.A(n_60748), .B(n_60735), .C(n_60767), .D(n_55325)
		, .Z(n_98113375));
	notech_nao3 i_118860578(.A(n_56460), .B(n_195658242), .C(n_995), .Z(n_260936764
		));
	notech_nao3 i_117960579(.A(n_56460), .B(n_195658242), .C(n_55825), .Z(n_261036765
		));
	notech_and3 i_44360596(.A(n_1012), .B(n_1014), .C(n_1006), .Z(n_262736782
		));
	notech_or2 i_43560598(.A(n_56369), .B(n_27597), .Z(n_262936784));
	notech_or4 i_28933190(.A(calc_sz[3]), .B(calc_sz[2]), .C(n_260688757), .D
		(n_56502), .Z(n_56060));
	notech_or4 i_23960603(.A(n_56460), .B(n_56487), .C(n_56478), .D(n_29010)
		, .Z(n_263436789));
	notech_ao4 i_35560600(.A(n_56502), .B(n_56560), .C(n_55807), .D(n_26582)
		, .Z(n_263136786));
	notech_or2 i_207160616(.A(n_54528), .B(n_55988), .Z(n_54453));
	notech_or4 i_207060617(.A(n_1909), .B(n_2202), .C(n_997), .D(n_55988), .Z
		(n_54454));
	notech_nand2 i_333155(.A(n_60504), .B(n_59375), .Z(n_56260));
	notech_or4 i_130760661(.A(n_1909), .B(n_2202), .C(n_997), .D(n_56000), .Z
		(n_55072));
	notech_and2 i_197960619(.A(n_56260), .B(n_1011), .Z(n_54528));
	notech_or2 i_130660662(.A(n_54528), .B(n_56000), .Z(n_55073));
	notech_and4 i_105260671(.A(n_55257), .B(n_318688503), .C(n_318288507), .D
		(n_55791), .Z(n_55317));
	notech_and4 i_105160672(.A(n_55265), .B(n_318788502), .C(n_318388506), .D
		(n_55790), .Z(n_55318));
	notech_ao4 i_93160683(.A(n_54874), .B(n_56551), .C(n_55825), .D(n_320888481
		), .Z(n_55430));
	notech_ao4 i_93060684(.A(n_1970), .B(n_60468), .C(n_55825), .D(n_54938),
		 .Z(n_55431));
	notech_and3 i_85460687(.A(n_55257), .B(n_318688503), .C(n_318288507), .Z
		(n_55500));
	notech_and3 i_85360688(.A(n_55265), .B(n_318788502), .C(n_318388506), .Z
		(n_55501));
	notech_and3 i_61160701(.A(n_131423301), .B(n_217058450), .C(n_55690), .Z
		(n_55739));
	notech_or4 i_56360705(.A(n_60583), .B(n_59894), .C(n_1900), .D(n_56551),
		 .Z(n_55786));
	notech_or4 i_56060706(.A(n_60768), .B(n_60721), .C(n_1970), .D(n_60584),
		 .Z(n_55789));
	notech_and2 i_138733173(.A(n_54698), .B(n_55325), .Z(n_55001));
	notech_or4 i_55960707(.A(n_60768), .B(n_60721), .C(n_60584), .D(n_55001)
		, .Z(n_55790));
	notech_nand3 i_55860708(.A(n_1016), .B(n_59186), .C(n_59807), .Z(n_55791
		));
	notech_or2 i_28833189(.A(n_56502), .B(n_56551), .Z(n_56061));
	notech_ao4 i_36160717(.A(n_56502), .B(n_56551), .C(n_55858), .D(n_26582)
		, .Z(n_55988));
	notech_nao3 i_29033042(.A(n_26599), .B(n_56551), .C(n_56502), .Z(n_56059
		));
	notech_ao4 i_34960718(.A(n_56502), .B(n_56538), .C(n_56369), .D(n_26582)
		, .Z(n_56000));
	notech_or2 i_29133191(.A(n_56569), .B(n_56502), .Z(n_56058));
	notech_ao4 i_34360719(.A(n_56573), .B(n_56502), .C(n_55827), .D(n_26582)
		, .Z(n_56006));
	notech_or2 i_27029(.A(n_56487), .B(n_28967), .Z(n_264436799));
	notech_or4 i_283(.A(n_60748), .B(n_60735), .C(n_60767), .D(n_60583), .Z(n_56066
		));
	notech_ao4 i_92570301(.A(n_2409), .B(n_56748), .C(n_2794), .D(n_29039), 
		.Z(n_2644));
	notech_and4 i_923(.A(n_264088752), .B(n_2631), .C(n_2636), .D(n_243556253
		), .Z(n_2642));
	notech_and4 i_920(.A(n_57312), .B(n_2637), .C(n_243456252), .D(n_243256250
		), .Z(n_264088752));
	notech_ao4 i_909(.A(n_2816), .B(n_28354), .C(n_2811), .D(n_28400), .Z(n_2637
		));
	notech_and3 i_919(.A(n_2634), .B(n_2633), .C(n_243156249), .Z(n_2636));
	notech_ao4 i_912(.A(n_2812), .B(n_56892), .C(n_280088689), .D(n_27578), 
		.Z(n_2634));
	notech_ao4 i_915(.A(n_2815), .B(n_28321), .C(n_55230), .D(n_55375), .Z(n_2633
		));
	notech_and4 i_918(.A(n_2628), .B(n_2627), .C(n_2626), .D(n_243356251), .Z
		(n_2631));
	notech_ao4 i_908(.A(n_56910), .B(n_27179), .C(n_56972), .D(n_27045), .Z(n_2628
		));
	notech_ao4 i_907(.A(n_57168), .B(n_27212), .C(n_2802), .D(n_28198), .Z(n_2627
		));
	notech_and4 i_910(.A(n_2623), .B(n_241956237), .C(n_2622), .D(n_242656244
		), .Z(n_2626));
	notech_ao4 i_903(.A(n_2813), .B(n_29038), .C(n_56640), .D(n_28096), .Z(n_2623
		));
	notech_and4 i_904(.A(n_241456232), .B(n_2619), .C(n_241556233), .D(n_241856236
		), .Z(n_2622));
	notech_and3 i_900(.A(n_2617), .B(n_241288763), .C(n_2413), .Z(n_2619));
	notech_ao4 i_896(.A(n_56932), .B(n_29036), .C(n_56921), .D(nbus_11326[13
		]), .Z(n_2617));
	notech_or4 i_514(.A(n_26663), .B(n_2340), .C(n_60558), .D(\opcode[1] ), 
		.Z(n_2616));
	notech_and3 i_117(.A(n_57371), .B(n_60479), .C(n_57358), .Z(n_2613));
	notech_or4 i_24(.A(n_59369), .B(n_60494), .C(n_106813462), .D(n_59894), 
		.Z(n_2612));
	notech_nao3 i_1754(.A(n_60540), .B(n_60504), .C(n_2588), .Z(n_2610));
	notech_nand2 i_489(.A(n_27404), .B(n_27402), .Z(n_260988754));
	notech_nand2 i_488(.A(calc_sz[2]), .B(n_27403), .Z(n_260888755));
	notech_nao3 i_485(.A(n_2042), .B(n_26867), .C(n_58940), .Z(n_260788756)
		);
	notech_nand2 i_481(.A(calc_sz[1]), .B(n_27402), .Z(n_260688757));
	notech_or2 i_25660(.A(calc_sz[2]), .B(calc_sz[3]), .Z(n_2605));
	notech_nao3 i_480(.A(n_2822), .B(n_275188706), .C(n_2603), .Z(n_2604));
	notech_nand3 i_1408(.A(n_2823), .B(n_275888699), .C(n_55641), .Z(n_2603)
		);
	notech_or4 i_512(.A(n_4737261), .B(n_26377), .C(n_26536), .D(n_26496), .Z
		(n_2601));
	notech_nand3 i_477(.A(n_27265), .B(n_27262), .C(n_27264), .Z(n_2599));
	notech_or4 i_471(.A(n_60748), .B(n_60735), .C(n_60767), .D(n_57326), .Z(n_2597
		));
	notech_nand2 i_1329(.A(n_276288695), .B(n_2593), .Z(n_2596));
	notech_nand2 i_25510(.A(n_276288695), .B(n_274788710), .Z(n_2594));
	notech_nao3 i_46362(.A(n_244056258), .B(n_27266), .C(fsm[1]), .Z(n_2593)
		);
	notech_nand2 i_25500(.A(n_222456215), .B(n_2225), .Z(n_2591));
	notech_nao3 i_200(.A(n_2385), .B(n_2361), .C(n_2831), .Z(n_2588));
	notech_or2 i_1111(.A(n_2361), .B(n_26869), .Z(n_2586));
	notech_nand3 i_2047(.A(n_60748), .B(n_60739), .C(n_27264), .Z(n_2585));
	notech_nand2 i_2010(.A(fsm[1]), .B(fsm[4]), .Z(n_2584));
	notech_or2 i_221(.A(fsm[1]), .B(n_27266), .Z(n_2582));
	notech_nao3 i_399(.A(n_27266), .B(n_27264), .C(fsm[1]), .Z(n_2580));
	notech_and2 i_1117(.A(n_2361), .B(n_26869), .Z(n_2578));
	notech_nor2 i_2046(.A(fsm[1]), .B(fsm[4]), .Z(n_2575));
	notech_nand2 i_73333184(.A(n_59210), .B(n_59958), .Z(n_2573));
	notech_nand2 i_1040(.A(n_2361), .B(n_2385), .Z(n_2572));
	notech_ao4 i_378(.A(n_245156269), .B(n_28521), .C(n_245756275), .D(n_28529
		), .Z(n_2569));
	notech_ao4 i_377(.A(n_245656274), .B(n_28537), .C(n_28545), .D(n_246156279
		), .Z(n_2568));
	notech_ao4 i_379(.A(n_245056268), .B(n_28505), .C(n_245256270), .D(n_28513
		), .Z(n_2567));
	notech_and2 i_727895(.A(n_2564), .B(n_2365), .Z(n_2565));
	notech_ao4 i_362(.A(n_247056288), .B(instrc[86]), .C(n_246956287), .D(instrc
		[78]), .Z(n_2564));
	notech_ao4 i_358(.A(instrc[94]), .B(n_247556293), .C(instrc[102]), .D(n_247456292
		), .Z(n_2563));
	notech_nao3 i_353(.A(n_235988764), .B(n_2560), .C(n_2360), .Z(n_2562));
	notech_and3 i_351(.A(n_2552), .B(n_2551), .C(n_2559), .Z(n_2560));
	notech_and4 i_350(.A(n_2557), .B(n_2556), .C(n_2554), .D(n_2358), .Z(n_2559
		));
	notech_ao4 i_344(.A(n_245156269), .B(n_28519), .C(n_245756275), .D(n_28527
		), .Z(n_2557));
	notech_ao4 i_343(.A(n_245656274), .B(n_28535), .C(n_246156279), .D(n_28543
		), .Z(n_2556));
	notech_ao4 i_342(.A(n_246056278), .B(n_28551), .C(n_247456292), .D(n_29033
		), .Z(n_2554));
	notech_ao4 i_346(.A(n_246956287), .B(n_28558), .C(n_247556293), .D(n_29034
		), .Z(n_2552));
	notech_ao4 i_345(.A(n_245056268), .B(n_28503), .C(n_245256270), .D(n_28511
		), .Z(n_2551));
	notech_or2 i_1455(.A(n_2340), .B(n_231756227), .Z(n_2550));
	notech_and4 i_323(.A(n_253988758), .B(n_253888759), .C(n_2546), .D(n_2338
		), .Z(n_2548));
	notech_and4 i_321(.A(n_2544), .B(n_2543), .C(n_2541), .D(n_2337), .Z(n_2546
		));
	notech_ao4 i_315(.A(n_245156269), .B(n_28522), .C(n_245756275), .D(n_28530
		), .Z(n_2544));
	notech_ao4 i_314(.A(n_245656274), .B(n_28538), .C(n_246156279), .D(n_28546
		), .Z(n_2543));
	notech_and2 i_16361(.A(pt_fault), .B(n_29792), .Z(n_67587010));
	notech_and2 i_25199(.A(had_lgjmp), .B(\nbus_14523[31] ), .Z(pg_en));
	notech_ao4 i_151068756(.A(n_21051), .B(n_27333), .C(n_56583), .D(n_26923
		), .Z(n_134587616));
	notech_ao4 i_150968757(.A(n_152160603), .B(n_28986), .C(n_135360435), .D
		(n_27297), .Z(n_134687617));
	notech_ao4 i_150668760(.A(n_21051), .B(n_27335), .C(n_56583), .D(n_26927
		), .Z(n_134787618));
	notech_ao4 i_150568761(.A(n_152160603), .B(n_29050), .C(n_135360435), .D
		(n_27300), .Z(n_134887619));
	notech_ao4 i_150468762(.A(n_21051), .B(n_27336), .C(n_56583), .D(n_26929
		), .Z(n_134987620));
	notech_ao4 i_150368763(.A(n_152160603), .B(n_29043), .C(n_135360435), .D
		(n_27301), .Z(n_135087621));
	notech_ao4 i_150268764(.A(n_21051), .B(n_27337), .C(n_56583), .D(n_26931
		), .Z(n_135187622));
	notech_ao4 i_150168765(.A(n_152160603), .B(n_29063), .C(n_135360435), .D
		(n_27302), .Z(n_135287623));
	notech_ao4 i_150068766(.A(n_21051), .B(n_27338), .C(n_56583), .D(n_26933
		), .Z(n_135387624));
	notech_ao4 i_149968767(.A(n_152160603), .B(n_29065), .C(n_135360435), .D
		(n_27304), .Z(n_135487625));
	notech_ao4 i_149868768(.A(n_21051), .B(n_27339), .C(n_56583), .D(n_26935
		), .Z(n_135587626));
	notech_ao4 i_149768769(.A(n_152160603), .B(n_29068), .C(n_135360435), .D
		(n_27307), .Z(n_135687627));
	notech_ao4 i_149668770(.A(n_21051), .B(n_27340), .C(n_56583), .D(n_26937
		), .Z(n_135787628));
	notech_ao4 i_149568771(.A(n_152160603), .B(n_28983), .C(n_135360435), .D
		(n_27308), .Z(n_135887629));
	notech_ao4 i_149468772(.A(n_21051), .B(n_27341), .C(n_56583), .D(n_26939
		), .Z(n_135987630));
	notech_ao4 i_149368773(.A(n_152160603), .B(n_29045), .C(n_135360435), .D
		(n_27309), .Z(n_136087631));
	notech_ao4 i_149268774(.A(n_21051), .B(n_27342), .C(n_56583), .D(n_26941
		), .Z(n_136187632));
	notech_ao4 i_149168775(.A(n_152160603), .B(n_29048), .C(n_135360435), .D
		(n_27310), .Z(n_136287633));
	notech_ao4 i_149068776(.A(n_21051), .B(n_27343), .C(n_56583), .D(n_26943
		), .Z(n_136387634));
	notech_ao4 i_148968777(.A(n_152160603), .B(n_29077), .C(n_135360435), .D
		(n_27311), .Z(n_136487635));
	notech_ao4 i_148868778(.A(n_21051), .B(n_27345), .C(n_56583), .D(n_26945
		), .Z(n_136587636));
	notech_ao4 i_148768779(.A(n_152160603), .B(n_29080), .C(n_135360435), .D
		(n_27312), .Z(n_136687637));
	notech_ao4 i_148668780(.A(n_21051), .B(n_27346), .C(n_56583), .D(n_26947
		), .Z(n_136787638));
	notech_ao4 i_148568781(.A(n_152160603), .B(n_29084), .C(n_135360435), .D
		(n_27313), .Z(n_136887639));
	notech_ao4 i_148468782(.A(n_21051), .B(n_27347), .C(n_56583), .D(n_26949
		), .Z(n_136987640));
	notech_ao4 i_148368783(.A(n_152160603), .B(n_29037), .C(n_135360435), .D
		(n_27314), .Z(n_137087641));
	notech_ao4 i_148268784(.A(n_21051), .B(n_27348), .C(n_56583), .D(n_26951
		), .Z(n_137187642));
	notech_ao4 i_148168785(.A(n_152160603), .B(n_29006), .C(n_135360435), .D
		(n_27315), .Z(n_137287643));
	notech_ao4 i_148068786(.A(n_21051), .B(n_27349), .C(n_56578), .D(n_26953
		), .Z(n_137387644));
	notech_ao4 i_147968787(.A(n_152160603), .B(n_29087), .C(n_53973), .D(n_27316
		), .Z(n_137487645));
	notech_ao4 i_147868788(.A(n_53307), .B(n_27350), .C(n_56578), .D(n_26955
		), .Z(n_137587646));
	notech_ao4 i_147768789(.A(n_53318), .B(n_29004), .C(n_53973), .D(n_27317
		), .Z(n_137687647));
	notech_ao4 i_147668790(.A(n_53307), .B(n_27351), .C(n_56578), .D(n_26957
		), .Z(n_137787648));
	notech_ao4 i_147568791(.A(n_53318), .B(n_28987), .C(n_53973), .D(n_27318
		), .Z(n_137887649));
	notech_ao4 i_147468792(.A(n_53307), .B(n_27352), .C(n_56578), .D(n_26959
		), .Z(n_137987650));
	notech_ao4 i_147368793(.A(n_53318), .B(n_29165), .C(n_53973), .D(n_27319
		), .Z(n_138087651));
	notech_ao4 i_147268794(.A(n_53307), .B(n_27353), .C(n_56578), .D(n_26961
		), .Z(n_138187652));
	notech_ao4 i_147168795(.A(n_53318), .B(n_29167), .C(n_53973), .D(n_27320
		), .Z(n_138287653));
	notech_ao4 i_147068796(.A(n_53307), .B(n_27354), .C(n_56578), .D(n_26963
		), .Z(n_138387654));
	notech_ao4 i_146968797(.A(n_53318), .B(n_29169), .C(n_53973), .D(n_27321
		), .Z(n_138487655));
	notech_ao4 i_146868798(.A(n_53307), .B(n_27355), .C(n_56578), .D(n_26965
		), .Z(n_138587656));
	notech_ao4 i_146768799(.A(n_53318), .B(n_29172), .C(n_53973), .D(n_27322
		), .Z(n_138687657));
	notech_ao4 i_146668800(.A(n_53307), .B(n_27356), .C(n_56578), .D(n_26967
		), .Z(n_138787658));
	notech_ao4 i_146568801(.A(n_53318), .B(n_29174), .C(n_53973), .D(n_27323
		), .Z(n_138887659));
	notech_ao4 i_146468802(.A(n_53307), .B(n_27357), .C(n_56578), .D(n_26969
		), .Z(n_138987660));
	notech_ao4 i_146368803(.A(n_53318), .B(n_29152), .C(n_53973), .D(n_27324
		), .Z(n_139087661));
	notech_ao4 i_146268804(.A(n_53307), .B(n_27358), .C(n_56578), .D(n_26971
		), .Z(n_139187662));
	notech_ao4 i_146168805(.A(n_53318), .B(n_29137), .C(n_53973), .D(n_27325
		), .Z(n_139287663));
	notech_ao4 i_146068806(.A(n_53307), .B(n_27359), .C(n_56578), .D(n_26973
		), .Z(n_139387664));
	notech_ao4 i_145968807(.A(n_53318), .B(n_29215), .C(n_53973), .D(n_27326
		), .Z(n_139487665));
	notech_ao4 i_145868808(.A(n_53307), .B(n_27360), .C(n_56583), .D(n_26975
		), .Z(n_139587666));
	notech_ao4 i_145768809(.A(n_53318), .B(n_29156), .C(n_135360435), .D(n_27327
		), .Z(n_139687667));
	notech_ao4 i_145668810(.A(n_53307), .B(n_27361), .C(n_56578), .D(n_26977
		), .Z(n_139787668));
	notech_ao4 i_145568811(.A(n_53318), .B(n_29154), .C(n_53973), .D(n_27328
		), .Z(n_139887669));
	notech_ao4 i_145468812(.A(n_53307), .B(n_27362), .C(n_56578), .D(n_26979
		), .Z(n_139987670));
	notech_ao4 i_145368813(.A(n_53318), .B(n_29219), .C(n_53973), .D(n_27329
		), .Z(n_140087671));
	notech_ao4 i_145268814(.A(n_53307), .B(n_27363), .C(n_56578), .D(n_26983
		), .Z(n_140187672));
	notech_ao4 i_145168815(.A(n_53318), .B(n_28977), .C(n_53973), .D(n_27330
		), .Z(n_140287673));
	notech_ao4 i_145068816(.A(n_53307), .B(n_27364), .C(n_56578), .D(n_26985
		), .Z(n_140387674));
	notech_ao4 i_144968817(.A(n_53318), .B(n_28997), .C(n_53973), .D(n_27331
		), .Z(n_140487675));
	notech_ao4 i_144668820(.A(n_152060602), .B(n_27333), .C(n_56425), .D(n_26923
		), .Z(n_140587676));
	notech_ao4 i_144568821(.A(n_151760599), .B(n_28051), .C(n_151960601), .D
		(n_27297), .Z(n_140687677));
	notech_ao4 i_144468822(.A(n_152060602), .B(n_27335), .C(n_56425), .D(n_26927
		), .Z(n_140787678));
	notech_ao4 i_144368823(.A(n_151760599), .B(n_28053), .C(n_151960601), .D
		(n_27300), .Z(n_140887679));
	notech_ao4 i_144268824(.A(n_152060602), .B(n_27336), .C(n_56425), .D(n_26929
		), .Z(n_140987680));
	notech_ao4 i_144168825(.A(n_151760599), .B(n_28054), .C(n_151960601), .D
		(n_27301), .Z(n_141087681));
	notech_ao4 i_144068826(.A(n_152060602), .B(n_27337), .C(n_56425), .D(n_26931
		), .Z(n_141187682));
	notech_ao4 i_143968827(.A(n_151760599), .B(n_28055), .C(n_151960601), .D
		(n_27302), .Z(n_141287683));
	notech_ao4 i_143868828(.A(n_152060602), .B(n_27338), .C(n_56425), .D(n_26933
		), .Z(n_141387684));
	notech_ao4 i_143768829(.A(n_151760599), .B(n_28056), .C(n_151960601), .D
		(n_27304), .Z(n_141487685));
	notech_ao4 i_143668830(.A(n_152060602), .B(n_27339), .C(n_56425), .D(n_26935
		), .Z(n_141587686));
	notech_ao4 i_143568831(.A(n_151760599), .B(n_28057), .C(n_151960601), .D
		(n_27307), .Z(n_141687687));
	notech_ao4 i_143468832(.A(n_152060602), .B(n_27340), .C(n_56425), .D(n_26937
		), .Z(n_141787688));
	notech_ao4 i_143368833(.A(n_151760599), .B(n_28058), .C(n_151960601), .D
		(n_27308), .Z(n_141887689));
	notech_ao4 i_143268834(.A(n_152060602), .B(n_27341), .C(n_56425), .D(n_26939
		), .Z(n_141987690));
	notech_ao4 i_143168835(.A(n_151760599), .B(n_28059), .C(n_151960601), .D
		(n_27309), .Z(n_142087691));
	notech_ao4 i_143068836(.A(n_152060602), .B(n_27342), .C(n_56425), .D(n_26941
		), .Z(n_142187692));
	notech_ao4 i_142968837(.A(n_151760599), .B(n_28060), .C(n_151960601), .D
		(n_27310), .Z(n_142287693));
	notech_ao4 i_142868838(.A(n_152060602), .B(n_27343), .C(n_56425), .D(n_26943
		), .Z(n_142387694));
	notech_ao4 i_142768839(.A(n_151760599), .B(n_28061), .C(n_151960601), .D
		(n_27311), .Z(n_142487695));
	notech_ao4 i_142668840(.A(n_152060602), .B(n_27345), .C(n_56425), .D(n_26945
		), .Z(n_142587696));
	notech_ao4 i_142568841(.A(n_151760599), .B(n_28062), .C(n_151960601), .D
		(n_27312), .Z(n_142687697));
	notech_ao4 i_142468842(.A(n_152060602), .B(n_27346), .C(n_56425), .D(n_26947
		), .Z(n_142787698));
	notech_ao4 i_142368843(.A(n_151760599), .B(n_28063), .C(n_151960601), .D
		(n_27313), .Z(n_142887699));
	notech_ao4 i_142268844(.A(n_152060602), .B(n_27347), .C(n_56425), .D(n_26949
		), .Z(n_142987700));
	notech_ao4 i_142168845(.A(n_151760599), .B(n_28064), .C(n_151960601), .D
		(n_27314), .Z(n_143087701));
	notech_ao4 i_142068846(.A(n_152060602), .B(n_27348), .C(n_56425), .D(n_26951
		), .Z(n_143187702));
	notech_ao4 i_141968847(.A(n_151760599), .B(n_28065), .C(n_151960601), .D
		(n_27315), .Z(n_143287703));
	notech_ao4 i_141868848(.A(n_152060602), .B(n_27349), .C(n_56420), .D(n_26953
		), .Z(n_143387704));
	notech_ao4 i_141768849(.A(n_151760599), .B(n_28066), .C(n_151960601), .D
		(n_27316), .Z(n_143487705));
	notech_ao4 i_141668850(.A(n_53245), .B(n_27350), .C(n_56420), .D(n_26955
		), .Z(n_143587706));
	notech_ao4 i_141568851(.A(n_53265), .B(n_28067), .C(n_53256), .D(n_27317
		), .Z(n_143687707));
	notech_ao4 i_141468852(.A(n_53245), .B(n_27351), .C(n_56420), .D(n_26957
		), .Z(n_143787708));
	notech_ao4 i_141368853(.A(n_53265), .B(n_28068), .C(n_53256), .D(n_27318
		), .Z(n_143887709));
	notech_ao4 i_141268854(.A(n_53245), .B(n_27352), .C(n_56420), .D(n_26959
		), .Z(n_143987710));
	notech_ao4 i_141168855(.A(n_53265), .B(n_28069), .C(n_53256), .D(n_27319
		), .Z(n_144087711));
	notech_ao4 i_141068856(.A(n_53245), .B(n_27353), .C(n_56420), .D(n_26961
		), .Z(n_144187712));
	notech_ao4 i_140968857(.A(n_53265), .B(n_28070), .C(n_53256), .D(n_27320
		), .Z(n_144287713));
	notech_ao4 i_140868858(.A(n_53245), .B(n_27354), .C(n_56420), .D(n_26963
		), .Z(n_144387714));
	notech_ao4 i_140768859(.A(n_53265), .B(n_28071), .C(n_53256), .D(n_27321
		), .Z(n_144487715));
	notech_ao4 i_140668860(.A(n_53245), .B(n_27355), .C(n_56420), .D(n_26965
		), .Z(n_147787716));
	notech_ao4 i_140568861(.A(n_53265), .B(n_28072), .C(n_53256), .D(n_27322
		), .Z(n_147887717));
	notech_ao4 i_140468862(.A(n_53245), .B(n_27356), .C(n_56420), .D(n_26967
		), .Z(n_147987718));
	notech_ao4 i_140368863(.A(n_53265), .B(n_28073), .C(n_53256), .D(n_27323
		), .Z(n_148087719));
	notech_ao4 i_140268864(.A(n_53245), .B(n_27357), .C(n_56420), .D(n_26969
		), .Z(n_148187720));
	notech_ao4 i_140168865(.A(n_53265), .B(n_28074), .C(n_53256), .D(n_27324
		), .Z(n_148287721));
	notech_ao4 i_140068866(.A(n_53245), .B(n_27358), .C(n_56420), .D(n_26971
		), .Z(n_148387722));
	notech_ao4 i_139968867(.A(n_53265), .B(n_28075), .C(n_53256), .D(n_27325
		), .Z(n_148487723));
	notech_ao4 i_139868868(.A(n_53245), .B(n_27359), .C(n_56420), .D(n_26973
		), .Z(n_148587724));
	notech_ao4 i_139768869(.A(n_53265), .B(n_28076), .C(n_53256), .D(n_27326
		), .Z(n_148687725));
	notech_ao4 i_139668870(.A(n_53245), .B(n_27360), .C(n_56425), .D(n_26975
		), .Z(n_148787726));
	notech_ao4 i_139568871(.A(n_53265), .B(n_28077), .C(n_151960601), .D(n_27327
		), .Z(n_148887727));
	notech_ao4 i_139468872(.A(n_53245), .B(n_27361), .C(n_56420), .D(n_26977
		), .Z(n_148987728));
	notech_ao4 i_139368873(.A(n_53265), .B(n_28078), .C(n_53256), .D(n_27328
		), .Z(n_149087729));
	notech_ao4 i_139268874(.A(n_53245), .B(n_27362), .C(n_56420), .D(n_26979
		), .Z(n_149187730));
	notech_ao4 i_139168875(.A(n_53265), .B(n_28079), .C(n_53256), .D(n_27329
		), .Z(n_149287731));
	notech_ao4 i_139068876(.A(n_53245), .B(n_27363), .C(n_56420), .D(n_26983
		), .Z(n_149387732));
	notech_ao4 i_138968877(.A(n_53265), .B(n_28080), .C(n_53256), .D(n_27330
		), .Z(n_149487733));
	notech_ao4 i_138868878(.A(n_53245), .B(n_27364), .C(n_56420), .D(n_26985
		), .Z(n_149587734));
	notech_ao4 i_138768879(.A(n_53265), .B(n_28081), .C(n_53256), .D(n_27331
		), .Z(n_149687735));
	notech_ao4 i_138668880(.A(n_53256), .B(n_27332), .C(n_53245), .D(n_27365
		), .Z(n_149787736));
	notech_ao4 i_138568881(.A(n_56420), .B(n_26987), .C(n_53265), .D(n_28082
		), .Z(n_149887737));
	notech_ao4 i_132168944(.A(n_176260844), .B(n_27333), .C(n_341962313), .D
		(n_26923), .Z(n_149987738));
	notech_ao4 i_132068945(.A(n_151060592), .B(n_29898), .C(n_171060792), .D
		(n_27297), .Z(n_150087739));
	notech_ao4 i_131968946(.A(n_176260844), .B(n_27334), .C(n_341962313), .D
		(n_26925), .Z(n_150187740));
	notech_ao4 i_131868947(.A(n_151060592), .B(n_29897), .C(n_171060792), .D
		(n_27298), .Z(n_150287741));
	notech_ao4 i_131768948(.A(n_176260844), .B(n_27335), .C(n_341962313), .D
		(n_26927), .Z(n_150387742));
	notech_ao4 i_131668949(.A(n_151060592), .B(n_29896), .C(n_171060792), .D
		(n_27300), .Z(n_150487743));
	notech_ao4 i_131568950(.A(n_176260844), .B(n_27336), .C(n_341962313), .D
		(n_26929), .Z(n_150587744));
	notech_ao4 i_131468951(.A(n_151060592), .B(n_29895), .C(n_171060792), .D
		(n_27301), .Z(n_150687745));
	notech_ao4 i_131368952(.A(n_176260844), .B(n_27337), .C(n_341962313), .D
		(n_26931), .Z(n_150787746));
	notech_ao4 i_131268953(.A(n_151060592), .B(n_29894), .C(n_171060792), .D
		(n_27302), .Z(n_150887747));
	notech_ao4 i_131168954(.A(n_176260844), .B(n_27338), .C(n_341962313), .D
		(n_26933), .Z(n_150987748));
	notech_ao4 i_131068955(.A(n_151060592), .B(n_29893), .C(n_171060792), .D
		(n_27304), .Z(n_151087749));
	notech_ao4 i_130968956(.A(n_176260844), .B(n_27339), .C(n_341962313), .D
		(n_26935), .Z(n_151187750));
	notech_ao4 i_130868957(.A(n_151060592), .B(n_29892), .C(n_171060792), .D
		(n_27307), .Z(n_151287751));
	notech_ao4 i_130768958(.A(n_176260844), .B(n_27340), .C(n_341962313), .D
		(n_26937), .Z(n_151387752));
	notech_ao4 i_130668959(.A(n_151060592), .B(n_29891), .C(n_171060792), .D
		(n_27308), .Z(n_151487753));
	notech_ao4 i_130568960(.A(n_176260844), .B(n_27341), .C(n_341962313), .D
		(n_26939), .Z(n_151587754));
	notech_ao4 i_130468961(.A(n_151060592), .B(n_29890), .C(n_171060792), .D
		(n_27309), .Z(n_151687755));
	notech_ao4 i_130368962(.A(n_176260844), .B(n_27342), .C(n_341962313), .D
		(n_26941), .Z(n_151787756));
	notech_ao4 i_130268963(.A(n_151060592), .B(n_29889), .C(n_171060792), .D
		(n_27310), .Z(n_151887757));
	notech_ao4 i_130168964(.A(n_176260844), .B(n_27343), .C(n_341962313), .D
		(n_26943), .Z(n_151987758));
	notech_ao4 i_130068965(.A(n_151060592), .B(n_29888), .C(n_171060792), .D
		(n_27311), .Z(n_152087759));
	notech_ao4 i_129968966(.A(n_176260844), .B(n_27345), .C(n_341962313), .D
		(n_26945), .Z(n_152187760));
	notech_ao4 i_129868967(.A(n_151060592), .B(n_29887), .C(n_171060792), .D
		(n_27312), .Z(n_152287761));
	notech_ao4 i_129768968(.A(n_176260844), .B(n_27346), .C(n_341962313), .D
		(n_26947), .Z(n_152387762));
	notech_ao4 i_129668969(.A(n_151060592), .B(n_29886), .C(n_171060792), .D
		(n_27313), .Z(n_152487763));
	notech_ao4 i_129568970(.A(n_176260844), .B(n_27347), .C(n_341962313), .D
		(n_26949), .Z(n_152587764));
	notech_ao4 i_129468971(.A(n_151060592), .B(n_29885), .C(n_171060792), .D
		(n_27314), .Z(n_152687765));
	notech_ao4 i_129368972(.A(n_53906), .B(n_27348), .C(n_56520), .D(n_26951
		), .Z(n_152787766));
	notech_ao4 i_129268973(.A(n_151060592), .B(n_29884), .C(n_171060792), .D
		(n_27315), .Z(n_152887767));
	notech_ao4 i_128968976(.A(n_53906), .B(n_27350), .C(n_56520), .D(n_26955
		), .Z(n_152987768));
	notech_ao4 i_128868977(.A(n_53051), .B(n_29883), .C(n_53946), .D(n_27317
		), .Z(n_153087769));
	notech_ao4 i_128768978(.A(n_53906), .B(n_27351), .C(n_56520), .D(n_26957
		), .Z(n_153187770));
	notech_ao4 i_128668979(.A(n_53051), .B(n_29882), .C(n_53946), .D(n_27318
		), .Z(n_153287771));
	notech_ao4 i_128568980(.A(n_53906), .B(n_27352), .C(n_56520), .D(n_26959
		), .Z(n_153387772));
	notech_ao4 i_128468981(.A(n_53051), .B(n_29881), .C(n_53946), .D(n_27319
		), .Z(n_153487773));
	notech_ao4 i_128368982(.A(n_53906), .B(n_27353), .C(n_56520), .D(n_26961
		), .Z(n_153587774));
	notech_ao4 i_128268983(.A(n_53051), .B(n_29880), .C(n_53946), .D(n_27320
		), .Z(n_153687775));
	notech_ao4 i_128168984(.A(n_53906), .B(n_27354), .C(n_56520), .D(n_26963
		), .Z(n_153787776));
	notech_ao4 i_128068985(.A(n_53051), .B(n_29879), .C(n_53946), .D(n_27321
		), .Z(n_153887777));
	notech_ao4 i_127968986(.A(n_53906), .B(n_27355), .C(n_56520), .D(n_26965
		), .Z(n_153987778));
	notech_ao4 i_127868987(.A(n_53051), .B(n_29878), .C(n_53946), .D(n_27322
		), .Z(n_154087779));
	notech_ao4 i_127768988(.A(n_53906), .B(n_27356), .C(n_56520), .D(n_26967
		), .Z(n_154187780));
	notech_ao4 i_127668989(.A(n_53051), .B(n_29877), .C(n_53946), .D(n_27323
		), .Z(n_154287781));
	notech_ao4 i_127568990(.A(n_53906), .B(n_27357), .C(n_56520), .D(n_26969
		), .Z(n_154387782));
	notech_ao4 i_127468991(.A(n_53051), .B(n_29876), .C(n_53946), .D(n_27324
		), .Z(n_154487783));
	notech_ao4 i_127368992(.A(n_53906), .B(n_27358), .C(n_56520), .D(n_26971
		), .Z(n_154587784));
	notech_ao4 i_127268993(.A(n_53051), .B(n_29875), .C(n_53946), .D(n_27325
		), .Z(n_154687785));
	notech_ao4 i_127168994(.A(n_53906), .B(n_27359), .C(n_56520), .D(n_26973
		), .Z(n_154787786));
	notech_ao4 i_127068995(.A(n_53051), .B(n_29874), .C(n_53946), .D(n_27326
		), .Z(n_154887787));
	notech_ao4 i_126968996(.A(n_176260844), .B(n_27360), .C(n_56520), .D(n_26975
		), .Z(n_154987788));
	notech_ao4 i_126868997(.A(n_53051), .B(n_29873), .C(n_171060792), .D(n_27327
		), .Z(n_155087789));
	notech_ao4 i_126768998(.A(n_53906), .B(n_27361), .C(n_56520), .D(n_26977
		), .Z(n_155187790));
	notech_ao4 i_126668999(.A(n_53051), .B(n_29872), .C(n_53946), .D(n_27328
		), .Z(n_155287791));
	notech_ao4 i_126569000(.A(n_53906), .B(n_27362), .C(n_56520), .D(n_26979
		), .Z(n_155387792));
	notech_ao4 i_126469001(.A(n_53051), .B(n_29871), .C(n_53946), .D(n_27329
		), .Z(n_155487793));
	notech_ao4 i_126369002(.A(n_53906), .B(n_27363), .C(n_56520), .D(n_26983
		), .Z(n_155587794));
	notech_ao4 i_126269003(.A(n_53051), .B(n_29870), .C(n_53946), .D(n_27330
		), .Z(n_155687795));
	notech_ao4 i_126169004(.A(n_53906), .B(n_27364), .C(n_56520), .D(n_26985
		), .Z(n_155787796));
	notech_ao4 i_126069005(.A(n_53051), .B(n_29868), .C(n_53946), .D(n_27331
		), .Z(n_155887797));
	notech_ao4 i_119669068(.A(n_150760589), .B(n_27333), .C(n_334662244), .D
		(n_26923), .Z(n_155987798));
	notech_ao4 i_119569069(.A(n_56147), .B(n_29867), .C(n_27297), .D(n_150660588
		), .Z(n_156087799));
	notech_ao4 i_119469070(.A(n_150760589), .B(n_27334), .C(n_334662244), .D
		(n_26925), .Z(n_156187800));
	notech_ao4 i_119369071(.A(n_56147), .B(n_29864), .C(n_150660588), .D(n_27298
		), .Z(n_156287801));
	notech_ao4 i_119269072(.A(n_150760589), .B(n_27335), .C(n_334662244), .D
		(n_26927), .Z(n_156387802));
	notech_ao4 i_119169073(.A(n_56147), .B(n_29863), .C(n_150660588), .D(n_27300
		), .Z(n_156487803));
	notech_ao4 i_119069074(.A(n_150760589), .B(n_27336), .C(n_334662244), .D
		(n_26929), .Z(n_156587804));
	notech_ao4 i_118969075(.A(n_56147), .B(n_29860), .C(n_150660588), .D(n_27301
		), .Z(n_156687805));
	notech_ao4 i_118869076(.A(n_150760589), .B(n_27337), .C(n_334662244), .D
		(n_26931), .Z(n_156787806));
	notech_ao4 i_118769077(.A(n_56147), .B(n_29859), .C(n_150660588), .D(n_27302
		), .Z(n_156887807));
	notech_ao4 i_118669078(.A(n_150760589), .B(n_27338), .C(n_334662244), .D
		(n_26933), .Z(n_156987808));
	notech_ao4 i_118569079(.A(n_56147), .B(n_29858), .C(n_150660588), .D(n_27304
		), .Z(n_157087809));
	notech_ao4 i_118469080(.A(n_150760589), .B(n_27339), .C(n_334662244), .D
		(n_26935), .Z(n_157187810));
	notech_ao4 i_118369081(.A(n_56147), .B(n_29856), .C(n_150660588), .D(n_27307
		), .Z(n_157287811));
	notech_ao4 i_118269082(.A(n_150760589), .B(n_27340), .C(n_334662244), .D
		(n_26937), .Z(n_157387812));
	notech_ao4 i_118169083(.A(n_56147), .B(n_29855), .C(n_150660588), .D(n_27308
		), .Z(n_157487813));
	notech_ao4 i_118069084(.A(n_150760589), .B(n_27341), .C(n_334662244), .D
		(n_26939), .Z(n_157587814));
	notech_ao4 i_117969085(.A(n_56147), .B(n_29854), .C(n_150660588), .D(n_27309
		), .Z(n_157687815));
	notech_ao4 i_117669088(.A(n_150760589), .B(n_27343), .C(n_334662244), .D
		(n_26943), .Z(n_157787816));
	notech_ao4 i_117569089(.A(n_56147), .B(n_29853), .C(n_150660588), .D(n_27311
		), .Z(n_157887817));
	notech_ao4 i_117469090(.A(n_150760589), .B(n_27345), .C(n_334662244), .D
		(n_26945), .Z(n_157987818));
	notech_ao4 i_117369091(.A(n_56147), .B(n_29852), .C(n_150660588), .D(n_27312
		), .Z(n_158087819));
	notech_ao4 i_117269092(.A(n_150760589), .B(n_27346), .C(n_334662244), .D
		(n_26947), .Z(n_158187820));
	notech_ao4 i_117169093(.A(n_56147), .B(n_29851), .C(n_150660588), .D(n_27313
		), .Z(n_158287821));
	notech_ao4 i_117069094(.A(n_150760589), .B(n_27347), .C(n_334662244), .D
		(n_26949), .Z(n_158387822));
	notech_ao4 i_116969095(.A(n_56147), .B(n_29850), .C(n_150660588), .D(n_27314
		), .Z(n_158487823));
	notech_ao4 i_116869096(.A(n_150760589), .B(n_27348), .C(n_334662244), .D
		(n_26951), .Z(n_158587824));
	notech_ao4 i_116769097(.A(n_56147), .B(n_29849), .C(n_150660588), .D(n_27315
		), .Z(n_158687825));
	notech_ao4 i_116669098(.A(n_150760589), .B(n_27349), .C(n_334662244), .D
		(n_26953), .Z(n_158787826));
	notech_ao4 i_116569099(.A(n_56147), .B(n_29848), .C(n_150660588), .D(n_27316
		), .Z(n_158887827));
	notech_ao4 i_116469100(.A(n_52670), .B(n_27350), .C(n_56529), .D(n_26955
		), .Z(n_158987828));
	notech_ao4 i_116369101(.A(n_52800), .B(n_29847), .C(n_52681), .D(n_27317
		), .Z(n_159087829));
	notech_ao4 i_116269102(.A(n_52670), .B(n_27351), .C(n_56529), .D(n_26957
		), .Z(n_159187830));
	notech_ao4 i_116169103(.A(n_52800), .B(n_29846), .C(n_52681), .D(n_27318
		), .Z(n_159287831));
	notech_ao4 i_116069104(.A(n_52670), .B(n_27352), .C(n_56529), .D(n_26959
		), .Z(n_159387832));
	notech_ao4 i_115969105(.A(n_52800), .B(n_29845), .C(n_52681), .D(n_27319
		), .Z(n_159487833));
	notech_ao4 i_115869106(.A(n_52670), .B(n_27353), .C(n_56529), .D(n_26961
		), .Z(n_159587834));
	notech_ao4 i_115769107(.A(n_52800), .B(n_29844), .C(n_52681), .D(n_27320
		), .Z(n_159687835));
	notech_ao4 i_115669108(.A(n_52670), .B(n_27354), .C(n_56529), .D(n_26963
		), .Z(n_159787836));
	notech_ao4 i_115569109(.A(n_52800), .B(n_29843), .C(n_52681), .D(n_27321
		), .Z(n_159887837));
	notech_ao4 i_115469110(.A(n_52670), .B(n_27355), .C(n_56529), .D(n_26965
		), .Z(n_159987838));
	notech_ao4 i_115369111(.A(n_52800), .B(n_29842), .C(n_52681), .D(n_27322
		), .Z(n_160087839));
	notech_ao4 i_115269112(.A(n_52670), .B(n_27356), .C(n_56529), .D(n_26967
		), .Z(n_160187840));
	notech_ao4 i_115169113(.A(n_52800), .B(n_29841), .C(n_52681), .D(n_27323
		), .Z(n_160287841));
	notech_ao4 i_115069114(.A(n_52670), .B(n_27357), .C(n_56529), .D(n_26969
		), .Z(n_160387842));
	notech_ao4 i_114969115(.A(n_52800), .B(n_29840), .C(n_52681), .D(n_27324
		), .Z(n_160487843));
	notech_ao4 i_114869116(.A(n_52670), .B(n_27358), .C(n_56529), .D(n_26971
		), .Z(n_160587844));
	notech_ao4 i_114769117(.A(n_52800), .B(n_29839), .C(n_52681), .D(n_27325
		), .Z(n_160687845));
	notech_ao4 i_114669118(.A(n_52670), .B(n_27359), .C(n_56529), .D(n_26973
		), .Z(n_160787846));
	notech_ao4 i_114569119(.A(n_52800), .B(n_29838), .C(n_52681), .D(n_27326
		), .Z(n_160887847));
	notech_ao4 i_114469120(.A(n_52670), .B(n_27360), .C(n_56529), .D(n_26975
		), .Z(n_160987848));
	notech_ao4 i_114369121(.A(n_52800), .B(n_29837), .C(n_150660588), .D(n_27327
		), .Z(n_161087849));
	notech_ao4 i_114269122(.A(n_52670), .B(n_27361), .C(n_56529), .D(n_26977
		), .Z(n_161187850));
	notech_ao4 i_114169123(.A(n_52800), .B(n_29836), .C(n_52681), .D(n_27328
		), .Z(n_161287851));
	notech_ao4 i_114069124(.A(n_52670), .B(n_27362), .C(n_56529), .D(n_26979
		), .Z(n_161387852));
	notech_ao4 i_113969125(.A(n_52800), .B(n_29835), .C(n_52681), .D(n_27329
		), .Z(n_161487853));
	notech_ao4 i_113869126(.A(n_52670), .B(n_27363), .C(n_56529), .D(n_26983
		), .Z(n_161587854));
	notech_ao4 i_113769127(.A(n_52800), .B(n_29833), .C(n_52681), .D(n_27330
		), .Z(n_161687855));
	notech_ao4 i_113669128(.A(n_52681), .B(n_27332), .C(n_52670), .D(n_27365
		), .Z(n_161787856));
	notech_ao4 i_113569129(.A(n_52800), .B(n_29832), .C(n_56529), .D(n_26987
		), .Z(n_161887857));
	notech_ao4 i_113469130(.A(n_27334), .B(n_150460586), .C(n_334962247), .D
		(n_26925), .Z(n_161987858));
	notech_ao4 i_113369131(.A(n_56160), .B(n_29831), .C(n_170960791), .D(n_27298
		), .Z(n_162087859));
	notech_ao4 i_113269132(.A(n_27335), .B(n_150460586), .C(n_334962247), .D
		(n_26927), .Z(n_162187860));
	notech_ao4 i_113169133(.A(n_56160), .B(n_29830), .C(n_170960791), .D(n_27300
		), .Z(n_162287861));
	notech_ao4 i_113069134(.A(n_27336), .B(n_150460586), .C(n_334962247), .D
		(n_26929), .Z(n_162387862));
	notech_ao4 i_112969135(.A(n_56160), .B(n_29829), .C(n_170960791), .D(n_27301
		), .Z(n_162487863));
	notech_ao4 i_112869136(.A(n_27337), .B(n_150460586), .C(n_334962247), .D
		(n_26931), .Z(n_162587864));
	notech_ao4 i_112769137(.A(n_56160), .B(n_29828), .C(n_170960791), .D(n_27302
		), .Z(n_162687865));
	notech_ao4 i_112669138(.A(n_27338), .B(n_150460586), .C(n_334962247), .D
		(n_26933), .Z(n_162787866));
	notech_ao4 i_112569139(.A(n_56160), .B(n_29827), .C(n_170960791), .D(n_27304
		), .Z(n_162887867));
	notech_ao4 i_112469140(.A(n_27339), .B(n_150460586), .C(n_334962247), .D
		(n_26935), .Z(n_162987868));
	notech_ao4 i_112369141(.A(n_56160), .B(n_29825), .C(n_170960791), .D(n_27307
		), .Z(n_163087869));
	notech_ao4 i_112269142(.A(n_27340), .B(n_150460586), .C(n_334962247), .D
		(n_26937), .Z(n_163187870));
	notech_ao4 i_112169143(.A(n_56160), .B(n_29824), .C(n_170960791), .D(n_27308
		), .Z(n_163287871));
	notech_ao4 i_112069144(.A(n_27341), .B(n_150460586), .C(n_334962247), .D
		(n_26939), .Z(n_163387872));
	notech_ao4 i_111969145(.A(n_56160), .B(n_29822), .C(n_170960791), .D(n_27309
		), .Z(n_163487873));
	notech_ao4 i_111869146(.A(n_27342), .B(n_150460586), .C(n_334962247), .D
		(n_26941), .Z(n_163587874));
	notech_ao4 i_111769147(.A(n_56160), .B(n_29821), .C(n_170960791), .D(n_27310
		), .Z(n_163687875));
	notech_ao4 i_111669148(.A(n_27343), .B(n_150460586), .C(n_334962247), .D
		(n_26943), .Z(n_163787876));
	notech_ao4 i_111569149(.A(n_56160), .B(n_29820), .C(n_170960791), .D(n_27311
		), .Z(n_163887877));
	notech_ao4 i_111469150(.A(n_27345), .B(n_150460586), .C(n_334962247), .D
		(n_26945), .Z(n_163987878));
	notech_ao4 i_111369151(.A(n_56160), .B(n_29819), .C(n_170960791), .D(n_27312
		), .Z(n_164087879));
	notech_ao4 i_111269152(.A(n_27346), .B(n_150460586), .C(n_334962247), .D
		(n_26947), .Z(n_164187880));
	notech_ao4 i_111169153(.A(n_56160), .B(n_29817), .C(n_170960791), .D(n_27313
		), .Z(n_164287881));
	notech_ao4 i_111069154(.A(n_27347), .B(n_150460586), .C(n_334962247), .D
		(n_26949), .Z(n_164387882));
	notech_ao4 i_110969155(.A(n_56160), .B(n_29815), .C(n_170960791), .D(n_27314
		), .Z(n_164487883));
	notech_ao4 i_110869156(.A(n_27348), .B(n_150460586), .C(n_334962247), .D
		(n_26951), .Z(n_164587884));
	notech_ao4 i_110769157(.A(n_56160), .B(n_29812), .C(n_170960791), .D(n_27315
		), .Z(n_164687885));
	notech_ao4 i_110669158(.A(n_27349), .B(n_150460586), .C(n_56327), .D(n_26953
		), .Z(n_164787886));
	notech_ao4 i_110569159(.A(n_56160), .B(n_29811), .C(n_170960791), .D(n_27316
		), .Z(n_164887887));
	notech_ao4 i_110469160(.A(n_27350), .B(n_52540), .C(n_56327), .D(n_26955
		), .Z(n_164987888));
	notech_ao4 i_110369161(.A(n_52659), .B(n_29809), .C(n_53955), .D(n_27317
		), .Z(n_165087889));
	notech_ao4 i_110269162(.A(n_27351), .B(n_52540), .C(n_56327), .D(n_26957
		), .Z(n_165187890));
	notech_ao4 i_110169163(.A(n_52659), .B(n_29808), .C(n_53955), .D(n_27318
		), .Z(n_165287891));
	notech_ao4 i_110069164(.A(n_27352), .B(n_52540), .C(n_56327), .D(n_26959
		), .Z(n_165387892));
	notech_ao4 i_109969165(.A(n_52659), .B(n_29807), .C(n_53955), .D(n_27319
		), .Z(n_165487893));
	notech_ao4 i_109869166(.A(n_27353), .B(n_52540), .C(n_56327), .D(n_26961
		), .Z(n_165587894));
	notech_ao4 i_109769167(.A(n_52659), .B(n_29806), .C(n_53955), .D(n_27320
		), .Z(n_165687895));
	notech_ao4 i_109669168(.A(n_27354), .B(n_52540), .C(n_56327), .D(n_26963
		), .Z(n_165787896));
	notech_ao4 i_109569169(.A(n_52659), .B(n_29805), .C(n_53955), .D(n_27321
		), .Z(n_165887897));
	notech_ao4 i_109469170(.A(n_27355), .B(n_52540), .C(n_56327), .D(n_26965
		), .Z(n_165987898));
	notech_ao4 i_109369171(.A(n_52659), .B(n_29804), .C(n_53955), .D(n_27322
		), .Z(n_166087899));
	notech_ao4 i_109169172(.A(n_27356), .B(n_52540), .C(n_56327), .D(n_26967
		), .Z(n_166187900));
	notech_ao4 i_109069173(.A(n_52659), .B(n_29803), .C(n_53955), .D(n_27323
		), .Z(n_166287901));
	notech_ao4 i_108969174(.A(n_27357), .B(n_52540), .C(n_56327), .D(n_26969
		), .Z(n_166387902));
	notech_ao4 i_108869175(.A(n_52659), .B(n_29801), .C(n_53955), .D(n_27324
		), .Z(n_166487903));
	notech_ao4 i_108769176(.A(n_27358), .B(n_52540), .C(n_56327), .D(n_26971
		), .Z(n_166587904));
	notech_ao4 i_108669177(.A(n_52659), .B(n_29800), .C(n_53955), .D(n_27325
		), .Z(n_166687905));
	notech_ao4 i_108569178(.A(n_27359), .B(n_52540), .C(n_56327), .D(n_26973
		), .Z(n_166787906));
	notech_ao4 i_108469179(.A(n_52659), .B(n_29799), .C(n_53955), .D(n_27326
		), .Z(n_166887907));
	notech_ao4 i_108369180(.A(n_27360), .B(n_150460586), .C(n_56327), .D(n_26975
		), .Z(n_166987908));
	notech_ao4 i_108269181(.A(n_52659), .B(n_29797), .C(n_170960791), .D(n_27327
		), .Z(n_167087909));
	notech_ao4 i_108169182(.A(n_27361), .B(n_52540), .C(n_56327), .D(n_26977
		), .Z(n_167187910));
	notech_ao4 i_108069183(.A(n_52659), .B(n_29796), .C(n_53955), .D(n_27328
		), .Z(n_167287911));
	notech_ao4 i_107769186(.A(n_27363), .B(n_52540), .C(n_56327), .D(n_26983
		), .Z(n_167387912));
	notech_ao4 i_107669187(.A(n_52659), .B(n_29795), .C(n_53955), .D(n_27330
		), .Z(n_167487913));
	notech_ao4 i_107569188(.A(n_27364), .B(n_52540), .C(n_56327), .D(n_26985
		), .Z(n_167587914));
	notech_ao4 i_107469189(.A(n_52659), .B(n_29794), .C(n_53955), .D(n_27331
		), .Z(n_167687915));
	notech_ao4 i_107369190(.A(n_53955), .B(n_27332), .C(n_27365), .D(n_52540
		), .Z(n_167787916));
	notech_ao4 i_107269191(.A(n_52659), .B(n_29793), .C(n_56327), .D(n_26987
		), .Z(n_167887917));
	notech_xor2 i_1368261(.A(all_cnt[2]), .B(n_55323), .Z(n_167987918));
	notech_xor2 i_1468260(.A(all_cnt[3]), .B(n_26624), .Z(n_168087919));
	notech_or4 i_14268148(.A(n_52245), .B(n_52364), .C(from_acu[3]), .D(n_27953
		), .Z(n_168187920));
	notech_or4 i_13668153(.A(from_acu[3]), .B(from_acu[2]), .C(n_52364), .D(n_27885
		), .Z(n_168887927));
	notech_nand2 i_111978(.A(n_178788026), .B(n_168187920), .Z(to_acu[0]));
	notech_or4 i_15768133(.A(n_52245), .B(n_52364), .C(from_acu[3]), .D(n_27954
		), .Z(n_168987928));
	notech_or4 i_15268138(.A(from_acu[3]), .B(from_acu[2]), .C(n_52364), .D(n_27886
		), .Z(n_169687935));
	notech_nand2 i_211979(.A(n_179388032), .B(n_168987928), .Z(to_acu[1]));
	notech_or4 i_17268118(.A(n_52245), .B(n_52364), .C(from_acu[3]), .D(n_27955
		), .Z(n_169787936));
	notech_or4 i_16768123(.A(from_acu[3]), .B(from_acu[2]), .C(n_52364), .D(n_27887
		), .Z(n_170487943));
	notech_nand2 i_311980(.A(n_179988038), .B(n_169787936), .Z(to_acu[2]));
	notech_or4 i_18768103(.A(n_52245), .B(n_52364), .C(from_acu[3]), .D(n_27956
		), .Z(n_170587944));
	notech_or4 i_18268108(.A(from_acu[3]), .B(from_acu[2]), .C(n_52364), .D(n_27888
		), .Z(n_171287951));
	notech_nand2 i_411981(.A(n_180588044), .B(n_170587944), .Z(to_acu[3]));
	notech_or4 i_20368088(.A(n_52248), .B(n_52367), .C(from_acu[3]), .D(n_27957
		), .Z(n_171387952));
	notech_or4 i_19868093(.A(from_acu[3]), .B(from_acu[2]), .C(n_52367), .D(n_27889
		), .Z(n_172087959));
	notech_nand2 i_511982(.A(n_181188050), .B(n_171387952), .Z(to_acu[4]));
	notech_or4 i_23368058(.A(n_52248), .B(n_52367), .C(from_acu[3]), .D(n_27959
		), .Z(n_172187960));
	notech_or4 i_22868063(.A(from_acu[3]), .B(from_acu[2]), .C(n_52367), .D(n_27893
		), .Z(n_172887967));
	notech_nand2 i_711984(.A(n_181788056), .B(n_172187960), .Z(to_acu[6]));
	notech_or4 i_24868043(.A(n_52248), .B(n_52367), .C(from_acu[3]), .D(n_27960
		), .Z(n_172987968));
	notech_or4 i_24368048(.A(from_acu[3]), .B(from_acu[2]), .C(n_52367), .D(n_27894
		), .Z(n_173687975));
	notech_nand2 i_811985(.A(n_182388062), .B(n_172987968), .Z(to_acu[7]));
	notech_or4 i_26468028(.A(n_52248), .B(n_52367), .C(from_acu[3]), .D(n_27961
		), .Z(n_173787976));
	notech_or4 i_25968033(.A(from_acu[3]), .B(from_acu[2]), .C(n_52367), .D(n_27895
		), .Z(n_174487983));
	notech_nand2 i_911986(.A(n_182988068), .B(n_173787976), .Z(to_acu[8]));
	notech_or4 i_27968013(.A(n_52247), .B(n_52366), .C(from_acu[3]), .D(n_27962
		), .Z(n_174587984));
	notech_or4 i_27468018(.A(from_acu[3]), .B(from_acu[2]), .C(n_52366), .D(n_27896
		), .Z(n_175287991));
	notech_nand2 i_1011987(.A(n_183588074), .B(n_174587984), .Z(to_acu[9])
		);
	notech_or4 i_30967983(.A(n_52247), .B(n_52366), .C(from_acu[3]), .D(n_27964
		), .Z(n_175387992));
	notech_or4 i_30467988(.A(from_acu[3]), .B(from_acu[2]), .C(n_52366), .D(n_27898
		), .Z(n_176087999));
	notech_nand2 i_1211989(.A(n_184188080), .B(n_175387992), .Z(to_acu[11])
		);
	notech_or4 i_32467968(.A(n_52247), .B(n_52366), .C(from_acu[3]), .D(n_27965
		), .Z(n_176188000));
	notech_or4 i_31967973(.A(from_acu[3]), .B(from_acu[2]), .C(n_52366), .D(n_27899
		), .Z(n_176888007));
	notech_nand2 i_1311990(.A(n_184788086), .B(n_176188000), .Z(to_acu[12])
		);
	notech_or4 i_59567698(.A(n_52247), .B(n_52366), .C(from_acu[3]), .D(n_27983
		), .Z(n_176988008));
	notech_or4 i_59067703(.A(from_acu[3]), .B(from_acu[2]), .C(n_52366), .D(n_27917
		), .Z(n_177688015));
	notech_nand2 i_3112008(.A(n_185388092), .B(n_176988008), .Z(to_acu[30])
		);
	notech_ao4 i_222479(.A(n_27556), .B(n_189388132), .C(n_59807), .D(n_2351
		), .Z(n_7831));
	notech_ao4 i_14568145(.A(n_52384), .B(n_27370), .C(n_52375), .D(n_27747)
		, .Z(n_178288021));
	notech_ao4 i_14668144(.A(n_52404), .B(n_27818), .C(n_52395), .D(n_27681)
		, .Z(n_178488023));
	notech_ao4 i_14768143(.A(n_52425), .B(n_28019), .C(n_52415), .D(n_27715)
		, .Z(n_178588024));
	notech_and4 i_15068140(.A(n_178588024), .B(n_178488023), .C(n_178288021)
		, .D(n_168887927), .Z(n_178788026));
	notech_ao4 i_16068130(.A(n_52384), .B(n_27371), .C(n_52375), .D(n_27748)
		, .Z(n_178888027));
	notech_ao4 i_16168129(.A(n_52404), .B(n_27819), .C(n_52395), .D(n_27682)
		, .Z(n_179088029));
	notech_ao4 i_16268128(.A(n_52425), .B(n_28020), .C(n_52415), .D(n_27716)
		, .Z(n_179188030));
	notech_and4 i_16568125(.A(n_179188030), .B(n_179088029), .C(n_178888027)
		, .D(n_169687935), .Z(n_179388032));
	notech_ao4 i_17568115(.A(n_52384), .B(n_27372), .C(n_52375), .D(n_27749)
		, .Z(n_179488033));
	notech_ao4 i_17668114(.A(n_52404), .B(n_27820), .C(n_52395), .D(n_27685)
		, .Z(n_179688035));
	notech_ao4 i_17768113(.A(n_52425), .B(n_28021), .C(n_52415), .D(n_27717)
		, .Z(n_179788036));
	notech_and4 i_18068110(.A(n_179788036), .B(n_179688035), .C(n_179488033)
		, .D(n_170487943), .Z(n_179988038));
	notech_ao4 i_19068100(.A(n_52384), .B(n_27373), .C(n_52375), .D(n_27750)
		, .Z(n_180088039));
	notech_ao4 i_19168099(.A(n_52404), .B(n_27821), .C(n_52395), .D(n_27686)
		, .Z(n_180288041));
	notech_ao4 i_19368098(.A(n_28022), .B(n_52425), .C(n_52415), .D(n_27718)
		, .Z(n_180388042));
	notech_and4 i_19668095(.A(n_180388042), .B(n_180288041), .C(n_180088039)
		, .D(n_171287951), .Z(n_180588044));
	notech_ao4 i_20668085(.A(n_52387), .B(n_27374), .C(n_52377), .D(n_27751)
		, .Z(n_180688045));
	notech_ao4 i_20768084(.A(n_52407), .B(n_27822), .C(n_52397), .D(n_27687)
		, .Z(n_180888047));
	notech_ao4 i_20868083(.A(n_52428), .B(n_28023), .C(n_52417), .D(n_27719)
		, .Z(n_180988048));
	notech_and4 i_21168080(.A(n_180988048), .B(n_180888047), .C(n_180688045)
		, .D(n_172087959), .Z(n_181188050));
	notech_ao4 i_23668055(.A(n_52387), .B(n_27376), .C(n_52377), .D(n_27753)
		, .Z(n_181288051));
	notech_ao4 i_23768054(.A(n_52407), .B(n_27824), .C(n_52397), .D(n_27689)
		, .Z(n_181488053));
	notech_ao4 i_23868053(.A(n_52428), .B(n_28025), .C(n_52417), .D(n_27721)
		, .Z(n_181588054));
	notech_and4 i_24168050(.A(n_181588054), .B(n_181488053), .C(n_181288051)
		, .D(n_172887967), .Z(n_181788056));
	notech_ao4 i_25168040(.A(n_52387), .B(n_27377), .C(n_52379), .D(n_27754)
		, .Z(n_181888057));
	notech_ao4 i_25368039(.A(n_52407), .B(n_27825), .C(n_52399), .D(n_27690)
		, .Z(n_182088059));
	notech_ao4 i_25468038(.A(n_52428), .B(n_28026), .C(n_52419), .D(n_27722)
		, .Z(n_182188060));
	notech_and4 i_25768035(.A(n_182188060), .B(n_182088059), .C(n_181888057)
		, .D(n_173687975), .Z(n_182388062));
	notech_ao4 i_26768025(.A(n_52387), .B(n_27378), .C(n_52377), .D(n_27755)
		, .Z(n_182488063));
	notech_ao4 i_26868024(.A(n_52407), .B(n_27826), .C(n_52397), .D(n_27691)
		, .Z(n_182688065));
	notech_ao4 i_26968023(.A(n_28027), .B(n_52428), .C(n_52417), .D(n_27723)
		, .Z(n_182788066));
	notech_and4 i_27268020(.A(n_182788066), .B(n_182688065), .C(n_182488063)
		, .D(n_174487983), .Z(n_182988068));
	notech_ao4 i_28268010(.A(n_52386), .B(n_27379), .C(n_52376), .D(n_27756)
		, .Z(n_183088069));
	notech_ao4 i_28368009(.A(n_52406), .B(n_27827), .C(n_52396), .D(n_27692)
		, .Z(n_183288071));
	notech_ao4 i_28468008(.A(n_52427), .B(n_28028), .C(n_52416), .D(n_27724)
		, .Z(n_183388072));
	notech_and4 i_28768005(.A(n_183388072), .B(n_183288071), .C(n_183088069)
		, .D(n_175287991), .Z(n_183588074));
	notech_ao4 i_31267980(.A(n_52386), .B(n_27381), .C(n_52376), .D(n_27758)
		, .Z(n_183688075));
	notech_ao4 i_31367979(.A(n_52406), .B(n_27829), .C(n_52396), .D(n_27694)
		, .Z(n_183888077));
	notech_ao4 i_31467978(.A(n_52427), .B(n_28030), .C(n_52416), .D(n_27726)
		, .Z(n_183988078));
	notech_and4 i_31767975(.A(n_183988078), .B(n_183888077), .C(n_183688075)
		, .D(n_176087999), .Z(n_184188080));
	notech_ao4 i_32767965(.A(n_52386), .B(n_27382), .C(n_52377), .D(n_27760)
		, .Z(n_184288081));
	notech_ao4 i_32867964(.A(n_52406), .B(n_27830), .C(n_52397), .D(n_27695)
		, .Z(n_184488083));
	notech_ao4 i_32967963(.A(n_28031), .B(n_52427), .C(n_52417), .D(n_27727)
		, .Z(n_184588084));
	notech_and4 i_33267960(.A(n_184588084), .B(n_184488083), .C(n_184288081)
		, .D(n_176888007), .Z(n_184788086));
	notech_ao4 i_59867695(.A(n_52386), .B(n_27400), .C(n_52377), .D(n_27784)
		, .Z(n_184888087));
	notech_ao4 i_59967694(.A(n_52406), .B(n_27848), .C(n_52397), .D(n_27713)
		, .Z(n_185088089));
	notech_ao4 i_60067693(.A(n_28049), .B(n_52427), .C(n_52417), .D(n_27745)
		, .Z(n_185188090));
	notech_and4 i_60367690(.A(n_185188090), .B(n_185088089), .C(n_184888087)
		, .D(n_177688015), .Z(n_185388092));
	notech_and2 i_16747(.A(opb[2]), .B(n_59807), .Z(n_185488093));
	notech_and2 i_16748(.A(opb[3]), .B(n_59807), .Z(n_185588094));
	notech_and2 i_16749(.A(opb[5]), .B(n_59809), .Z(n_185688095));
	notech_and2 i_16750(.A(opb[6]), .B(n_59807), .Z(n_185788096));
	notech_and2 i_16751(.A(opb[7]), .B(n_59807), .Z(n_185888097));
	notech_and2 i_16752(.A(opb[8]), .B(n_59807), .Z(n_185988098));
	notech_and2 i_16753(.A(opb[9]), .B(n_59807), .Z(n_186088099));
	notech_and2 i_16754(.A(opb[10]), .B(n_59807), .Z(n_186188100));
	notech_and2 i_16755(.A(opb[11]), .B(n_59807), .Z(n_186288101));
	notech_and2 i_16756(.A(opb[12]), .B(n_59819), .Z(n_186388102));
	notech_and2 i_16757(.A(opb[13]), .B(n_59819), .Z(n_186488103));
	notech_and2 i_16758(.A(opb[14]), .B(n_59819), .Z(n_186588104));
	notech_and2 i_16759(.A(opb[15]), .B(n_59819), .Z(n_186688105));
	notech_ao3 i_72362849(.A(temp_ss[31]), .B(n_56578), .C(n_53973), .Z(n_188188120
		));
	notech_or2 i_72462848(.A(n_53307), .B(n_27365), .Z(n_188288121));
	notech_ao4 i_150262090(.A(n_56578), .B(n_26987), .C(n_53318), .D(n_28996
		), .Z(n_188588124));
	notech_ao4 i_148962103(.A(n_53906), .B(n_27365), .C(n_53946), .D(n_27332
		), .Z(n_188688125));
	notech_ao4 i_148862104(.A(n_56520), .B(n_26987), .C(n_53051), .D(n_29901
		), .Z(n_188788126));
	notech_ao4 i_147862114(.A(n_52681), .B(n_27331), .C(n_52670), .D(n_27364
		), .Z(n_188888127));
	notech_ao4 i_147762115(.A(n_56529), .B(n_26985), .C(n_52800), .D(n_29900
		), .Z(n_188988128));
	notech_ao4 i_147362119(.A(n_27333), .B(n_52540), .C(n_27297), .D(n_53955
		), .Z(n_189088129));
	notech_ao4 i_147262120(.A(n_56327), .B(n_26923), .C(n_52659), .D(n_29899
		), .Z(n_189188130));
	notech_ao4 i_313(.A(n_246056278), .B(n_28553), .C(n_247456292), .D(n_29029
		), .Z(n_2541));
	notech_ao4 i_317(.A(n_246956287), .B(n_28561), .C(n_247556293), .D(n_29030
		), .Z(n_253988758));
	notech_ao4 i_316(.A(n_245056268), .B(n_28506), .C(n_245256270), .D(n_28514
		), .Z(n_253888759));
	notech_and4 i_295(.A(n_2527), .B(n_2526), .C(n_2534), .D(n_231588765), .Z
		(n_2536));
	notech_and4 i_293(.A(n_2532), .B(n_2531), .C(n_2529), .D(n_231456226), .Z
		(n_2534));
	notech_ao4 i_287(.A(n_245156269), .B(n_28520), .C(n_245756275), .D(n_28528
		), .Z(n_2532));
	notech_ao4 i_286(.A(n_245656274), .B(n_28536), .C(n_246156279), .D(n_28544
		), .Z(n_2531));
	notech_ao4 i_285(.A(n_246056278), .B(n_28552), .C(n_247456292), .D(n_29025
		), .Z(n_2529));
	notech_ao4 i_289(.A(n_246956287), .B(n_28559), .C(n_247556293), .D(n_29026
		), .Z(n_2527));
	notech_ao4 i_288(.A(n_245056268), .B(n_28504), .C(n_245256270), .D(n_28512
		), .Z(n_2526));
	notech_and4 i_266(.A(n_2515), .B(n_2514), .C(n_2522), .D(n_230188772), .Z
		(n_2524));
	notech_and4 i_264(.A(n_2520), .B(n_2519), .C(n_2517), .D(n_230088773), .Z
		(n_2522));
	notech_ao4 i_257(.A(n_245156269), .B(n_28516), .C(n_245756275), .D(n_28524
		), .Z(n_2520));
	notech_ao4 i_256(.A(n_245656274), .B(n_28532), .C(n_246156279), .D(n_28540
		), .Z(n_2519));
	notech_ao4 i_255(.A(n_246056278), .B(n_28548), .C(n_247456292), .D(n_29022
		), .Z(n_2517));
	notech_ao4 i_260(.A(n_246956287), .B(n_28555), .C(n_247556293), .D(n_29023
		), .Z(n_2515));
	notech_ao4 i_259(.A(n_245056268), .B(n_28500), .C(n_245256270), .D(n_28508
		), .Z(n_2514));
	notech_and4 i_236(.A(n_2503), .B(n_250288762), .C(n_2510), .D(n_228788786
		), .Z(n_2512));
	notech_and4 i_234(.A(n_2508), .B(n_2507), .C(n_2505), .D(n_228688787), .Z
		(n_2510));
	notech_mux2 i_112266(.S(n_60125), .A(n_1445), .B(regs_14[0]), .Z(pc_out[
		0]));
	notech_mux2 i_212267(.S(n_60125), .A(n_1446), .B(regs_14[1]), .Z(pc_out[
		1]));
	notech_mux2 i_312268(.S(n_60125), .A(n_1447), .B(regs_14[2]), .Z(pc_out[
		2]));
	notech_mux2 i_412269(.S(n_60125), .A(n_1448), .B(regs_14[3]), .Z(pc_out[
		3]));
	notech_mux2 i_512270(.S(n_60130), .A(n_1449), .B(regs_14[4]), .Z(pc_out[
		4]));
	notech_mux2 i_612271(.S(n_60130), .A(n_1450), .B(regs_14[5]), .Z(pc_out[
		5]));
	notech_mux2 i_712272(.S(n_60125), .A(n_1451), .B(regs_14[6]), .Z(pc_out[
		6]));
	notech_mux2 i_812273(.S(n_60130), .A(n_1452), .B(regs_14[7]), .Z(pc_out[
		7]));
	notech_mux2 i_912274(.S(n_60125), .A(n_1453), .B(regs_14[8]), .Z(pc_out[
		8]));
	notech_mux2 i_1012275(.S(n_60125), .A(n_1454), .B(regs_14[9]), .Z(pc_out
		[9]));
	notech_mux2 i_1112276(.S(n_60125), .A(n_1455), .B(regs_14[10]), .Z(pc_out
		[10]));
	notech_mux2 i_1212277(.S(n_60125), .A(n_1456), .B(regs_14[11]), .Z(pc_out
		[11]));
	notech_mux2 i_1312278(.S(n_60125), .A(n_1457), .B(regs_14[12]), .Z(pc_out
		[12]));
	notech_mux2 i_1412279(.S(n_60125), .A(n_1458), .B(regs_14[13]), .Z(pc_out
		[13]));
	notech_mux2 i_1512280(.S(n_60125), .A(n_1459), .B(regs_14[14]), .Z(pc_out
		[14]));
	notech_mux2 i_1612281(.S(n_60125), .A(n_1460), .B(regs_14[15]), .Z(pc_out
		[15]));
	notech_mux2 i_1712282(.S(n_60125), .A(n_1461), .B(regs_14[16]), .Z(pc_out
		[16]));
	notech_mux2 i_1812283(.S(n_60130), .A(n_1462), .B(regs_14[17]), .Z(pc_out
		[17]));
	notech_mux2 i_1912284(.S(n_60130), .A(n_1463), .B(regs_14[18]), .Z(pc_out
		[18]));
	notech_mux2 i_2012285(.S(n_60130), .A(n_1464), .B(regs_14[19]), .Z(pc_out
		[19]));
	notech_mux2 i_2112286(.S(n_60130), .A(n_1465), .B(regs_14[20]), .Z(pc_out
		[20]));
	notech_mux2 i_2212287(.S(n_60130), .A(n_1466), .B(regs_14[21]), .Z(pc_out
		[21]));
	notech_mux2 i_2312288(.S(n_60130), .A(n_1467), .B(regs_14[22]), .Z(pc_out
		[22]));
	notech_mux2 i_2412289(.S(n_60136), .A(n_1468), .B(regs_14[23]), .Z(pc_out
		[23]));
	notech_mux2 i_2512290(.S(n_60130), .A(n_1469), .B(regs_14[24]), .Z(pc_out
		[24]));
	notech_mux2 i_2612291(.S(n_60130), .A(n_1470), .B(regs_14[25]), .Z(pc_out
		[25]));
	notech_mux2 i_2712292(.S(n_60130), .A(n_1471), .B(regs_14[26]), .Z(pc_out
		[26]));
	notech_mux2 i_2812293(.S(n_60130), .A(n_1472), .B(regs_14[27]), .Z(pc_out
		[27]));
	notech_mux2 i_2912294(.S(n_60130), .A(n_1473), .B(regs_14[28]), .Z(pc_out
		[28]));
	notech_mux2 i_3012295(.S(n_60130), .A(n_1474), .B(regs_14[29]), .Z(pc_out
		[29]));
	notech_mux2 i_3112296(.S(n_60130), .A(n_1475), .B(regs_14[30]), .Z(pc_out
		[30]));
	notech_mux2 i_3212297(.S(n_60130), .A(n_1476), .B(regs_14[31]), .Z(pc_out
		[31]));
	notech_nand2 i_117675(.A(n_134687617), .B(n_134587616), .Z(write_data_25
		[0]));
	notech_nand2 i_317677(.A(n_134887619), .B(n_134787618), .Z(write_data_25
		[2]));
	notech_nand2 i_417678(.A(n_135087621), .B(n_134987620), .Z(write_data_25
		[3]));
	notech_nand2 i_517679(.A(n_135287623), .B(n_135187622), .Z(write_data_25
		[4]));
	notech_nand2 i_617680(.A(n_135487625), .B(n_135387624), .Z(write_data_25
		[5]));
	notech_nand2 i_717681(.A(n_135687627), .B(n_135587626), .Z(write_data_25
		[6]));
	notech_nand2 i_817682(.A(n_135887629), .B(n_135787628), .Z(write_data_25
		[7]));
	notech_nand2 i_917683(.A(n_136087631), .B(n_135987630), .Z(write_data_25
		[8]));
	notech_nand2 i_1017684(.A(n_136287633), .B(n_136187632), .Z(write_data_25
		[9]));
	notech_nand2 i_1117685(.A(n_136487635), .B(n_136387634), .Z(write_data_25
		[10]));
	notech_nand2 i_1217686(.A(n_136687637), .B(n_136587636), .Z(write_data_25
		[11]));
	notech_nand2 i_1317687(.A(n_136887639), .B(n_136787638), .Z(write_data_25
		[12]));
	notech_nand2 i_1417688(.A(n_137087641), .B(n_136987640), .Z(write_data_25
		[13]));
	notech_nand2 i_1517689(.A(n_137287643), .B(n_137187642), .Z(write_data_25
		[14]));
	notech_nand2 i_1617690(.A(n_137487645), .B(n_137387644), .Z(write_data_25
		[15]));
	notech_nand2 i_1717691(.A(n_137687647), .B(n_137587646), .Z(write_data_25
		[16]));
	notech_nand2 i_1817692(.A(n_137887649), .B(n_137787648), .Z(write_data_25
		[17]));
	notech_nand2 i_1917693(.A(n_138087651), .B(n_137987650), .Z(write_data_25
		[18]));
	notech_nand2 i_2017694(.A(n_138287653), .B(n_138187652), .Z(write_data_25
		[19]));
	notech_nand2 i_2117695(.A(n_138487655), .B(n_138387654), .Z(write_data_25
		[20]));
	notech_nand2 i_2217696(.A(n_138687657), .B(n_138587656), .Z(write_data_25
		[21]));
	notech_nand2 i_2317697(.A(n_138887659), .B(n_138787658), .Z(write_data_25
		[22]));
	notech_nand2 i_2417698(.A(n_139087661), .B(n_138987660), .Z(write_data_25
		[23]));
	notech_nand2 i_2517699(.A(n_139287663), .B(n_139187662), .Z(write_data_25
		[24]));
	notech_nand2 i_2617700(.A(n_139487665), .B(n_139387664), .Z(write_data_25
		[25]));
	notech_nand2 i_2717701(.A(n_139687667), .B(n_139587666), .Z(write_data_25
		[26]));
	notech_nand2 i_2817702(.A(n_139887669), .B(n_139787668), .Z(write_data_25
		[27]));
	notech_nand2 i_2917703(.A(n_140087671), .B(n_139987670), .Z(write_data_25
		[28]));
	notech_nand2 i_3017704(.A(n_140287673), .B(n_140187672), .Z(write_data_25
		[29]));
	notech_nand2 i_3117705(.A(n_140487675), .B(n_140387674), .Z(write_data_25
		[30]));
	notech_nand2 i_117931(.A(n_140687677), .B(n_140587676), .Z(write_data_27
		[0]));
	notech_nand2 i_317933(.A(n_140887679), .B(n_140787678), .Z(write_data_27
		[2]));
	notech_nand2 i_417934(.A(n_141087681), .B(n_140987680), .Z(write_data_27
		[3]));
	notech_nand2 i_517935(.A(n_141287683), .B(n_141187682), .Z(write_data_27
		[4]));
	notech_nand2 i_617936(.A(n_141487685), .B(n_141387684), .Z(write_data_27
		[5]));
	notech_nand2 i_717937(.A(n_141687687), .B(n_141587686), .Z(write_data_27
		[6]));
	notech_nand2 i_817938(.A(n_141887689), .B(n_141787688), .Z(write_data_27
		[7]));
	notech_nand2 i_917939(.A(n_142087691), .B(n_141987690), .Z(write_data_27
		[8]));
	notech_nand2 i_1017940(.A(n_142287693), .B(n_142187692), .Z(write_data_27
		[9]));
	notech_nand2 i_1117941(.A(n_142487695), .B(n_142387694), .Z(write_data_27
		[10]));
	notech_nand2 i_1217942(.A(n_142687697), .B(n_142587696), .Z(write_data_27
		[11]));
	notech_nand2 i_1317943(.A(n_142887699), .B(n_142787698), .Z(write_data_27
		[12]));
	notech_nand2 i_1417944(.A(n_143087701), .B(n_142987700), .Z(write_data_27
		[13]));
	notech_nand2 i_1517945(.A(n_143287703), .B(n_143187702), .Z(write_data_27
		[14]));
	notech_nand2 i_1617946(.A(n_143487705), .B(n_143387704), .Z(write_data_27
		[15]));
	notech_nand2 i_1717947(.A(n_143687707), .B(n_143587706), .Z(write_data_27
		[16]));
	notech_nand2 i_1817948(.A(n_143887709), .B(n_143787708), .Z(write_data_27
		[17]));
	notech_nand2 i_1917949(.A(n_144087711), .B(n_143987710), .Z(write_data_27
		[18]));
	notech_nand2 i_2017950(.A(n_144287713), .B(n_144187712), .Z(write_data_27
		[19]));
	notech_nand2 i_2117951(.A(n_144487715), .B(n_144387714), .Z(write_data_27
		[20]));
	notech_nand2 i_2217952(.A(n_147887717), .B(n_147787716), .Z(write_data_27
		[21]));
	notech_nand2 i_2317953(.A(n_148087719), .B(n_147987718), .Z(write_data_27
		[22]));
	notech_nand2 i_2417954(.A(n_148287721), .B(n_148187720), .Z(write_data_27
		[23]));
	notech_nand2 i_2517955(.A(n_148487723), .B(n_148387722), .Z(write_data_27
		[24]));
	notech_nand2 i_2617956(.A(n_148687725), .B(n_148587724), .Z(write_data_27
		[25]));
	notech_nand2 i_2717957(.A(n_148887727), .B(n_148787726), .Z(write_data_27
		[26]));
	notech_nand2 i_2817958(.A(n_149087729), .B(n_148987728), .Z(write_data_27
		[27]));
	notech_nand2 i_2917959(.A(n_149287731), .B(n_149187730), .Z(write_data_27
		[28]));
	notech_nand2 i_3017960(.A(n_149487733), .B(n_149387732), .Z(write_data_27
		[29]));
	notech_nand2 i_3117961(.A(n_149687735), .B(n_149587734), .Z(write_data_27
		[30]));
	notech_nand2 i_3217962(.A(n_149887737), .B(n_149787736), .Z(write_data_27
		[31]));
	notech_nand2 i_118187(.A(n_150087739), .B(n_149987738), .Z(write_data_29
		[0]));
	notech_nand2 i_218188(.A(n_150287741), .B(n_150187740), .Z(write_data_29
		[1]));
	notech_nand2 i_318189(.A(n_150487743), .B(n_150387742), .Z(write_data_29
		[2]));
	notech_nand2 i_418190(.A(n_150687745), .B(n_150587744), .Z(write_data_29
		[3]));
	notech_nand2 i_518191(.A(n_150887747), .B(n_150787746), .Z(write_data_29
		[4]));
	notech_nand2 i_618192(.A(n_151087749), .B(n_150987748), .Z(write_data_29
		[5]));
	notech_nand2 i_718193(.A(n_151287751), .B(n_151187750), .Z(write_data_29
		[6]));
	notech_nand2 i_818194(.A(n_151487753), .B(n_151387752), .Z(write_data_29
		[7]));
	notech_nand2 i_918195(.A(n_151687755), .B(n_151587754), .Z(write_data_29
		[8]));
	notech_nand2 i_1018196(.A(n_151887757), .B(n_151787756), .Z(write_data_29
		[9]));
	notech_nand2 i_1118197(.A(n_152087759), .B(n_151987758), .Z(write_data_29
		[10]));
	notech_nand2 i_1218198(.A(n_152287761), .B(n_152187760), .Z(write_data_29
		[11]));
	notech_nand2 i_1318199(.A(n_152487763), .B(n_152387762), .Z(write_data_29
		[12]));
	notech_nand2 i_1418200(.A(n_152687765), .B(n_152587764), .Z(write_data_29
		[13]));
	notech_nand2 i_1518201(.A(n_152887767), .B(n_152787766), .Z(write_data_29
		[14]));
	notech_nand2 i_1718203(.A(n_153087769), .B(n_152987768), .Z(write_data_29
		[16]));
	notech_nand2 i_1818204(.A(n_153287771), .B(n_153187770), .Z(write_data_29
		[17]));
	notech_nand2 i_1918205(.A(n_153487773), .B(n_153387772), .Z(write_data_29
		[18]));
	notech_nand2 i_2018206(.A(n_153687775), .B(n_153587774), .Z(write_data_29
		[19]));
	notech_nand2 i_2118207(.A(n_153887777), .B(n_153787776), .Z(write_data_29
		[20]));
	notech_nand2 i_2218208(.A(n_154087779), .B(n_153987778), .Z(write_data_29
		[21]));
	notech_nand2 i_2318209(.A(n_154287781), .B(n_154187780), .Z(write_data_29
		[22]));
	notech_nand2 i_2418210(.A(n_154487783), .B(n_154387782), .Z(write_data_29
		[23]));
	notech_nand2 i_2518211(.A(n_154687785), .B(n_154587784), .Z(write_data_29
		[24]));
	notech_nand2 i_2618212(.A(n_154887787), .B(n_154787786), .Z(write_data_29
		[25]));
	notech_nand2 i_2718213(.A(n_155087789), .B(n_154987788), .Z(write_data_29
		[26]));
	notech_nand2 i_2818214(.A(n_155287791), .B(n_155187790), .Z(write_data_29
		[27]));
	notech_nand2 i_2918215(.A(n_155487793), .B(n_155387792), .Z(write_data_29
		[28]));
	notech_nand2 i_3018216(.A(n_155687795), .B(n_155587794), .Z(write_data_29
		[29]));
	notech_nand2 i_3118217(.A(n_155887797), .B(n_155787796), .Z(write_data_29
		[30]));
	notech_nand2 i_118443(.A(n_156087799), .B(n_155987798), .Z(write_data_31
		[0]));
	notech_nand2 i_218444(.A(n_156287801), .B(n_156187800), .Z(write_data_31
		[1]));
	notech_nand2 i_318445(.A(n_156487803), .B(n_156387802), .Z(write_data_31
		[2]));
	notech_nand2 i_418446(.A(n_156687805), .B(n_156587804), .Z(write_data_31
		[3]));
	notech_nand2 i_518447(.A(n_156887807), .B(n_156787806), .Z(write_data_31
		[4]));
	notech_nand2 i_618448(.A(n_157087809), .B(n_156987808), .Z(write_data_31
		[5]));
	notech_nand2 i_718449(.A(n_157287811), .B(n_157187810), .Z(write_data_31
		[6]));
	notech_nand2 i_818450(.A(n_157487813), .B(n_157387812), .Z(write_data_31
		[7]));
	notech_nand2 i_918451(.A(n_157687815), .B(n_157587814), .Z(write_data_31
		[8]));
	notech_nand2 i_1118453(.A(n_157887817), .B(n_157787816), .Z(write_data_31
		[10]));
	notech_nand2 i_1218454(.A(n_158087819), .B(n_157987818), .Z(write_data_31
		[11]));
	notech_nand2 i_1318455(.A(n_158287821), .B(n_158187820), .Z(write_data_31
		[12]));
	notech_nand2 i_1418456(.A(n_158487823), .B(n_158387822), .Z(write_data_31
		[13]));
	notech_nand2 i_1518457(.A(n_158687825), .B(n_158587824), .Z(write_data_31
		[14]));
	notech_nand2 i_1618458(.A(n_158887827), .B(n_158787826), .Z(write_data_31
		[15]));
	notech_nand2 i_1718459(.A(n_159087829), .B(n_158987828), .Z(write_data_31
		[16]));
	notech_nand2 i_1818460(.A(n_159287831), .B(n_159187830), .Z(write_data_31
		[17]));
	notech_nand2 i_1918461(.A(n_159487833), .B(n_159387832), .Z(write_data_31
		[18]));
	notech_nand2 i_2018462(.A(n_159687835), .B(n_159587834), .Z(write_data_31
		[19]));
	notech_nand2 i_2118463(.A(n_159887837), .B(n_159787836), .Z(write_data_31
		[20]));
	notech_nand2 i_2218464(.A(n_160087839), .B(n_159987838), .Z(write_data_31
		[21]));
	notech_nand2 i_2318465(.A(n_160287841), .B(n_160187840), .Z(write_data_31
		[22]));
	notech_nand2 i_2418466(.A(n_160487843), .B(n_160387842), .Z(write_data_31
		[23]));
	notech_nand2 i_2518467(.A(n_160687845), .B(n_160587844), .Z(write_data_31
		[24]));
	notech_nand2 i_2618468(.A(n_160887847), .B(n_160787846), .Z(write_data_31
		[25]));
	notech_nand2 i_2718469(.A(n_161087849), .B(n_160987848), .Z(write_data_31
		[26]));
	notech_nand2 i_2818470(.A(n_161287851), .B(n_161187850), .Z(write_data_31
		[27]));
	notech_nand2 i_2918471(.A(n_161487853), .B(n_161387852), .Z(write_data_31
		[28]));
	notech_nand2 i_3018472(.A(n_161687855), .B(n_161587854), .Z(write_data_31
		[29]));
	notech_nand2 i_3218474(.A(n_161887857), .B(n_161787856), .Z(write_data_31
		[31]));
	notech_nand2 i_218572(.A(n_162087859), .B(n_161987858), .Z(write_data_32
		[1]));
	notech_nand2 i_318573(.A(n_162287861), .B(n_162187860), .Z(write_data_32
		[2]));
	notech_nand2 i_418574(.A(n_162487863), .B(n_162387862), .Z(write_data_32
		[3]));
	notech_nand2 i_518575(.A(n_162687865), .B(n_162587864), .Z(write_data_32
		[4]));
	notech_nand2 i_618576(.A(n_162887867), .B(n_162787866), .Z(write_data_32
		[5]));
	notech_nand2 i_718577(.A(n_163087869), .B(n_162987868), .Z(write_data_32
		[6]));
	notech_nand2 i_818578(.A(n_163287871), .B(n_163187870), .Z(write_data_32
		[7]));
	notech_nand2 i_918579(.A(n_163487873), .B(n_163387872), .Z(write_data_32
		[8]));
	notech_nand2 i_1018580(.A(n_163687875), .B(n_163587874), .Z(write_data_32
		[9]));
	notech_nand2 i_1118581(.A(n_163887877), .B(n_163787876), .Z(write_data_32
		[10]));
	notech_nand2 i_1218582(.A(n_164087879), .B(n_163987878), .Z(write_data_32
		[11]));
	notech_nand2 i_1318583(.A(n_164287881), .B(n_164187880), .Z(write_data_32
		[12]));
	notech_nand2 i_1418584(.A(n_164487883), .B(n_164387882), .Z(write_data_32
		[13]));
	notech_nand2 i_1518585(.A(n_164687885), .B(n_164587884), .Z(write_data_32
		[14]));
	notech_nand2 i_1618586(.A(n_164887887), .B(n_164787886), .Z(write_data_32
		[15]));
	notech_nand2 i_1718587(.A(n_165087889), .B(n_164987888), .Z(write_data_32
		[16]));
	notech_nand2 i_1818588(.A(n_165287891), .B(n_165187890), .Z(write_data_32
		[17]));
	notech_nand2 i_1918589(.A(n_165487893), .B(n_165387892), .Z(write_data_32
		[18]));
	notech_nand2 i_2018590(.A(n_165687895), .B(n_165587894), .Z(write_data_32
		[19]));
	notech_nand2 i_2118591(.A(n_165887897), .B(n_165787896), .Z(write_data_32
		[20]));
	notech_nand2 i_2218592(.A(n_166087899), .B(n_165987898), .Z(write_data_32
		[21]));
	notech_nand2 i_2318593(.A(n_166287901), .B(n_166187900), .Z(write_data_32
		[22]));
	notech_nand2 i_2418594(.A(n_166487903), .B(n_166387902), .Z(write_data_32
		[23]));
	notech_nand2 i_2518595(.A(n_166687905), .B(n_166587904), .Z(write_data_32
		[24]));
	notech_nand2 i_2618596(.A(n_166887907), .B(n_166787906), .Z(write_data_32
		[25]));
	notech_nand2 i_2718597(.A(n_167087909), .B(n_166987908), .Z(write_data_32
		[26]));
	notech_nand2 i_2818598(.A(n_167287911), .B(n_167187910), .Z(write_data_32
		[27]));
	notech_nand2 i_3018600(.A(n_167487913), .B(n_167387912), .Z(write_data_32
		[29]));
	notech_nand2 i_3118601(.A(n_167687915), .B(n_167587914), .Z(write_data_32
		[30]));
	notech_nand2 i_3218602(.A(n_167887917), .B(n_167787916), .Z(write_data_32
		[31]));
	notech_xor2 i_22370263(.A(\eflags[7] ), .B(\eflags[11] ), .Z(\cond[12] )
		);
	notech_nand2 i_6770264(.A(n_29792), .B(n_59186), .Z(\nbus_11274[0] ));
	notech_or2 i_121170262(.A(\eflags[6] ), .B(\cond[12] ), .Z(\cond[14] )
		);
	notech_or2 i_98770261(.A(\eflags[0] ), .B(\eflags[6] ), .Z(\cond[6] ));
	notech_mux2 i_3211721(.S(n_60423), .A(cr2[31]), .B(icr2[31]), .Z(n_7797)
		);
	notech_mux2 i_3111720(.S(n_60423), .A(cr2[30]), .B(icr2[30]), .Z(n_7791)
		);
	notech_mux2 i_3011719(.S(n_60423), .A(cr2[29]), .B(icr2[29]), .Z(n_7785)
		);
	notech_mux2 i_2911718(.S(n_60423), .A(cr2[28]), .B(icr2[28]), .Z(n_7779)
		);
	notech_mux2 i_2811717(.S(n_60423), .A(cr2[27]), .B(icr2[27]), .Z(n_7773)
		);
	notech_mux2 i_2711716(.S(n_60423), .A(cr2[26]), .B(icr2[26]), .Z(n_7767)
		);
	notech_mux2 i_2611715(.S(n_60423), .A(cr2[25]), .B(icr2[25]), .Z(n_7761)
		);
	notech_mux2 i_2511714(.S(n_60423), .A(cr2[24]), .B(icr2[24]), .Z(n_7755)
		);
	notech_mux2 i_2411713(.S(n_60419), .A(cr2[23]), .B(icr2[23]), .Z(n_7749)
		);
	notech_mux2 i_2311712(.S(n_60419), .A(cr2[22]), .B(icr2[22]), .Z(n_7743)
		);
	notech_mux2 i_2211711(.S(n_60419), .A(cr2[21]), .B(icr2[21]), .Z(n_7737)
		);
	notech_mux2 i_2111710(.S(n_60423), .A(cr2[20]), .B(icr2[20]), .Z(n_7731)
		);
	notech_mux2 i_2011709(.S(n_60423), .A(cr2[19]), .B(icr2[19]), .Z(n_7725)
		);
	notech_mux2 i_1911708(.S(n_60423), .A(cr2[18]), .B(icr2[18]), .Z(n_7719)
		);
	notech_mux2 i_1811707(.S(n_60423), .A(cr2[17]), .B(icr2[17]), .Z(n_7713)
		);
	notech_mux2 i_1711706(.S(n_60423), .A(cr2[16]), .B(icr2[16]), .Z(n_7707)
		);
	notech_mux2 i_1611705(.S(n_60424), .A(cr2[15]), .B(icr2[15]), .Z(n_7701)
		);
	notech_mux2 i_1511704(.S(n_60424), .A(cr2[14]), .B(icr2[14]), .Z(n_7695)
		);
	notech_mux2 i_1411703(.S(n_60424), .A(cr2[13]), .B(icr2[13]), .Z(n_7689)
		);
	notech_mux2 i_1311702(.S(n_60424), .A(cr2[12]), .B(icr2[12]), .Z(n_7683)
		);
	notech_mux2 i_1211701(.S(n_60424), .A(cr2[11]), .B(icr2[11]), .Z(n_7677)
		);
	notech_mux2 i_1111700(.S(n_60424), .A(cr2[10]), .B(icr2[10]), .Z(n_7671)
		);
	notech_mux2 i_1011699(.S(n_60424), .A(cr2[9]), .B(icr2[9]), .Z(n_7665)
		);
	notech_mux2 i_911698(.S(n_60424), .A(cr2[8]), .B(icr2[8]), .Z(n_7659));
	notech_mux2 i_811697(.S(n_60424), .A(cr2[7]), .B(icr2[7]), .Z(n_7653));
	notech_mux2 i_711696(.S(n_60424), .A(cr2[6]), .B(icr2[6]), .Z(n_7647));
	notech_mux2 i_611695(.S(n_60423), .A(cr2[5]), .B(icr2[5]), .Z(n_7641));
	notech_mux2 i_511694(.S(n_60424), .A(cr2[4]), .B(icr2[4]), .Z(n_7635));
	notech_mux2 i_411693(.S(n_60424), .A(cr2[3]), .B(icr2[3]), .Z(n_7629));
	notech_mux2 i_311692(.S(n_60424), .A(cr2[2]), .B(icr2[2]), .Z(n_7623));
	notech_mux2 i_211691(.S(n_60424), .A(cr2[1]), .B(icr2[1]), .Z(n_7617));
	notech_mux2 i_111690(.S(n_60415), .A(cr2[0]), .B(icr2[0]), .Z(n_7611));
	notech_mux2 i_3211753(.S(n_55326), .A(n_852), .B(n_851), .Z(n_16184));
	notech_mux2 i_3111752(.S(n_55322), .A(n_850), .B(n_849), .Z(n_16177));
	notech_mux2 i_3011751(.S(n_55326), .A(n_848), .B(n_847), .Z(n_16170));
	notech_mux2 i_2911750(.S(n_55326), .A(n_846), .B(n_845), .Z(n_16163));
	notech_mux2 i_2811749(.S(n_55326), .A(n_844), .B(n_843), .Z(n_16156));
	notech_mux2 i_2711748(.S(n_55322), .A(n_842), .B(n_841), .Z(n_16149));
	notech_mux2 i_2611747(.S(n_55322), .A(n_840), .B(n_839), .Z(n_16142));
	notech_mux2 i_2511746(.S(n_55322), .A(n_838), .B(n_837), .Z(n_16135));
	notech_mux2 i_2411745(.S(n_55322), .A(n_836), .B(n_835), .Z(n_16128));
	notech_mux2 i_2311744(.S(n_55322), .A(n_834), .B(n_833), .Z(n_16121));
	notech_mux2 i_2211743(.S(n_55326), .A(n_832), .B(n_831), .Z(n_16114));
	notech_mux2 i_2111742(.S(n_55326), .A(n_830), .B(n_829), .Z(n_16107));
	notech_mux2 i_2011741(.S(n_55326), .A(n_828), .B(n_827), .Z(n_16100));
	notech_mux2 i_1911740(.S(n_55326), .A(n_826), .B(n_825), .Z(n_16093));
	notech_mux2 i_1811739(.S(n_55326), .A(n_824), .B(n_823), .Z(n_16086));
	notech_mux2 i_1711738(.S(n_55326), .A(n_822), .B(n_821), .Z(n_16079));
	notech_mux2 i_1611737(.S(n_55326), .A(n_820), .B(n_819), .Z(n_16072));
	notech_mux2 i_1511736(.S(n_55326), .A(n_818), .B(n_817), .Z(n_16065));
	notech_mux2 i_1411735(.S(n_55326), .A(n_816), .B(n_815), .Z(n_16058));
	notech_mux2 i_1311734(.S(n_55326), .A(n_814), .B(n_813), .Z(n_16051));
	notech_mux2 i_1211733(.S(n_55322), .A(n_812), .B(n_811), .Z(n_16044));
	notech_mux2 i_1111732(.S(n_55326), .A(n_810), .B(n_809), .Z(n_16037));
	notech_mux2 i_1011731(.S(n_55326), .A(n_808), .B(n_807), .Z(n_16030));
	notech_mux2 i_911730(.S(n_55326), .A(n_806), .B(n_805), .Z(n_16023));
	notech_mux2 i_811729(.S(n_55326), .A(n_804), .B(n_803), .Z(n_16016));
	notech_mux2 i_711728(.S(n_55326), .A(n_802), .B(n_801), .Z(n_16009));
	notech_mux2 i_611727(.S(n_55326), .A(n_800), .B(n_799), .Z(n_16002));
	notech_mux2 i_511726(.S(n_55322), .A(n_798), .B(n_797), .Z(n_15995));
	notech_mux2 i_411725(.S(n_55322), .A(n_796), .B(n_795), .Z(n_15988));
	notech_mux2 i_311724(.S(n_55322), .A(n_794), .B(n_793), .Z(n_15981));
	notech_mux2 i_211723(.S(n_55322), .A(n_792), .B(n_791), .Z(n_15974));
	notech_mux2 i_111722(.S(n_55322), .A(n_790), .B(n_789), .Z(n_15967));
	notech_ao4 i_225(.A(n_245156269), .B(n_28515), .C(n_245756275), .D(n_28523
		), .Z(n_2508));
	notech_ao4 i_224(.A(n_245656274), .B(n_28531), .C(n_246156279), .D(n_28539
		), .Z(n_2507));
	notech_or2 i_25029(.A(all_cnt[0]), .B(n_59819), .Z(n_189388132));
	notech_and2 i_25032(.A(n_167987918), .B(n_59899), .Z(n_189488133));
	notech_and2 i_25033(.A(n_168087919), .B(n_59899), .Z(n_189588134));
	notech_ao4 i_223(.A(n_246056278), .B(n_28547), .C(n_247456292), .D(n_29019
		), .Z(n_2505));
	notech_ao4 i_227(.A(n_246956287), .B(n_28554), .C(n_247556293), .D(n_29020
		), .Z(n_2503));
	notech_ao4 i_226(.A(n_245056268), .B(n_28499), .C(n_245256270), .D(n_28507
		), .Z(n_250288762));
	notech_and4 i_193(.A(n_2491), .B(n_2490), .C(n_2498), .D(n_227388800), .Z
		(n_2500));
	notech_and4 i_191(.A(n_2496), .B(n_2495), .C(n_2493), .D(n_227288801), .Z
		(n_2498));
	notech_ao4 i_185(.A(n_245156269), .B(n_28518), .C(n_245756275), .D(n_28526
		), .Z(n_2496));
	notech_ao4 i_184(.A(n_245656274), .B(n_28534), .C(n_246156279), .D(n_28542
		), .Z(n_2495));
	notech_nao3 i_3217706(.A(n_188588124), .B(n_188288121), .C(n_188188120),
		 .Z(write_data_25[31]));
	notech_nand2 i_3218218(.A(n_188788126), .B(n_188688125), .Z(write_data_29
		[31]));
	notech_nand2 i_3118473(.A(n_188988128), .B(n_188888127), .Z(write_data_31
		[30]));
	notech_nand2 i_118571(.A(n_189188130), .B(n_189088129), .Z(write_data_32
		[0]));
	notech_nand3 i_8221(.A(n_26625), .B(n_273688719), .C(n_59899), .Z(n_11475
		));
	notech_ao4 i_183(.A(n_246056278), .B(n_28550), .C(n_247456292), .D(n_29016
		), .Z(n_2493));
	notech_reg_set fsmf_reg_0(.CP(n_62061), .D(n_60739), .SD(n_61176), .Q(fsmf
		[0]));
	notech_reg_set fsmf_reg_1(.CP(n_62061), .D(fsm[1]), .SD(n_61176), .Q(fsmf
		[1]));
	notech_reg_set fsmf_reg_2(.CP(n_62061), .D(fsm[2]), .SD(n_61176), .Q(fsmf
		[2]));
	notech_reg_set fsmf_reg_3(.CP(n_62061), .D(n_60752), .SD(n_61176), .Q(fsmf
		[3]));
	notech_reg fsmf_reg_4(.CP(n_62061), .D(fsm[4]), .CD(n_61176), .Q(fsmf[4]
		));
	notech_reg calc_sz_reg_0(.CP(n_62061), .D(n_16591), .CD(n_61175), .Q(calc_sz
		[0]));
	notech_mux2 i_71(.S(n_26628), .A(calc_sz[0]), .B(instrc[108]), .Z(n_16591
		));
	notech_reg calc_sz_reg_1(.CP(n_62061), .D(n_16597), .CD(n_61175), .Q(calc_sz
		[1]));
	notech_mux2 i_86(.S(n_26628), .A(calc_sz[1]), .B(instrc[109]), .Z(n_16597
		));
	notech_ao4 i_187(.A(n_246956287), .B(n_28557), .C(n_247556293), .D(n_29017
		), .Z(n_2491));
	notech_reg calc_sz_reg_2(.CP(n_62061), .D(n_16603), .CD(n_61175), .Q(calc_sz
		[2]));
	notech_mux2 i_110(.S(n_26628), .A(calc_sz[2]), .B(instrc[110]), .Z(n_16603
		));
	notech_ao4 i_186(.A(n_245056268), .B(n_28502), .C(n_245256270), .D(n_28510
		), .Z(n_2490));
	notech_reg calc_sz_reg_3(.CP(n_62061), .D(n_16609), .CD(n_61175), .Q(calc_sz
		[3]));
	notech_mux2 i_451(.S(n_26628), .A(calc_sz[3]), .B(instrc[111]), .Z(n_16609
		));
	notech_reg tsc_reg_0(.CP(n_62061), .D(n_363), .CD(n_61175), .Q(tsc[0])
		);
	notech_reg tsc_reg_1(.CP(n_62061), .D(n_365), .CD(n_61175), .Q(tsc[1])
		);
	notech_reg tsc_reg_2(.CP(n_62061), .D(n_367), .CD(n_61175), .Q(tsc[2])
		);
	notech_reg tsc_reg_3(.CP(n_62163), .D(n_369), .CD(n_61175), .Q(tsc[3])
		);
	notech_reg tsc_reg_4(.CP(n_62163), .D(n_371), .CD(n_61175), .Q(tsc[4])
		);
	notech_reg tsc_reg_5(.CP(n_62163), .D(n_373), .CD(n_61176), .Q(tsc[5])
		);
	notech_reg tsc_reg_6(.CP(n_62163), .D(n_375), .CD(n_61177), .Q(tsc[6])
		);
	notech_reg tsc_reg_7(.CP(n_62163), .D(n_377), .CD(n_61177), .Q(tsc[7])
		);
	notech_reg tsc_reg_8(.CP(n_62163), .D(n_379), .CD(n_61177), .Q(tsc[8])
		);
	notech_reg tsc_reg_9(.CP(n_62163), .D(n_381), .CD(n_61177), .Q(tsc[9])
		);
	notech_reg tsc_reg_10(.CP(n_62163), .D(n_383), .CD(n_61177), .Q(tsc[10])
		);
	notech_reg tsc_reg_11(.CP(n_62163), .D(n_385), .CD(n_61177), .Q(tsc[11])
		);
	notech_reg tsc_reg_12(.CP(n_62163), .D(n_387), .CD(n_61178), .Q(tsc[12])
		);
	notech_reg tsc_reg_13(.CP(n_62163), .D(n_389), .CD(n_61177), .Q(tsc[13])
		);
	notech_reg tsc_reg_14(.CP(n_62163), .D(n_391), .CD(n_61177), .Q(tsc[14])
		);
	notech_reg tsc_reg_15(.CP(n_62163), .D(n_393), .CD(n_61176), .Q(tsc[15])
		);
	notech_reg tsc_reg_16(.CP(n_62163), .D(n_395), .CD(n_61176), .Q(tsc[16])
		);
	notech_reg tsc_reg_17(.CP(n_62163), .D(n_397), .CD(n_61176), .Q(tsc[17])
		);
	notech_reg tsc_reg_18(.CP(n_62163), .D(n_399), .CD(n_61176), .Q(tsc[18])
		);
	notech_reg tsc_reg_19(.CP(n_62163), .D(n_401), .CD(n_61177), .Q(tsc[19])
		);
	notech_reg tsc_reg_20(.CP(n_62163), .D(n_403), .CD(n_61177), .Q(tsc[20])
		);
	notech_reg tsc_reg_21(.CP(n_62163), .D(n_405), .CD(n_61177), .Q(tsc[21])
		);
	notech_reg tsc_reg_22(.CP(n_62161), .D(n_407), .CD(n_61177), .Q(tsc[22])
		);
	notech_reg tsc_reg_23(.CP(n_62161), .D(n_409), .CD(n_61177), .Q(tsc[23])
		);
	notech_reg tsc_reg_24(.CP(n_62223), .D(n_411), .CD(n_61171), .Q(tsc[24])
		);
	notech_reg tsc_reg_25(.CP(n_62223), .D(n_413), .CD(n_61169), .Q(tsc[25])
		);
	notech_reg tsc_reg_26(.CP(n_62223), .D(n_415), .CD(n_61170), .Q(tsc[26])
		);
	notech_reg tsc_reg_27(.CP(n_62223), .D(n_417), .CD(n_61169), .Q(tsc[27])
		);
	notech_reg tsc_reg_28(.CP(n_62223), .D(n_419), .CD(n_61169), .Q(tsc[28])
		);
	notech_reg tsc_reg_29(.CP(n_62223), .D(n_421), .CD(n_61170), .Q(tsc[29])
		);
	notech_reg tsc_reg_30(.CP(n_62223), .D(n_423), .CD(n_61170), .Q(tsc[30])
		);
	notech_reg tsc_reg_31(.CP(n_62223), .D(n_425), .CD(n_61170), .Q(tsc[31])
		);
	notech_reg tsc_reg_32(.CP(n_62223), .D(n_427), .CD(n_61170), .Q(tsc[32])
		);
	notech_reg tsc_reg_33(.CP(n_62223), .D(n_429), .CD(n_61170), .Q(tsc[33])
		);
	notech_reg tsc_reg_34(.CP(n_62223), .D(n_431), .CD(n_61169), .Q(tsc[34])
		);
	notech_reg tsc_reg_35(.CP(n_62223), .D(n_433), .CD(n_61169), .Q(tsc[35])
		);
	notech_reg tsc_reg_36(.CP(n_62223), .D(n_435), .CD(n_61169), .Q(tsc[36])
		);
	notech_reg tsc_reg_37(.CP(n_62223), .D(n_437), .CD(n_61169), .Q(tsc[37])
		);
	notech_reg tsc_reg_38(.CP(n_62223), .D(n_439), .CD(n_61169), .Q(tsc[38])
		);
	notech_reg tsc_reg_39(.CP(n_62223), .D(n_441), .CD(n_61169), .Q(tsc[39])
		);
	notech_reg tsc_reg_40(.CP(n_62223), .D(n_443), .CD(n_61169), .Q(tsc[40])
		);
	notech_reg tsc_reg_41(.CP(n_62223), .D(n_445), .CD(n_61169), .Q(tsc[41])
		);
	notech_reg tsc_reg_42(.CP(n_62161), .D(n_447), .CD(n_61169), .Q(tsc[42])
		);
	notech_reg tsc_reg_43(.CP(n_62161), .D(n_449), .CD(n_61170), .Q(tsc[43])
		);
	notech_reg tsc_reg_44(.CP(n_62161), .D(n_451), .CD(n_61171), .Q(tsc[44])
		);
	notech_reg tsc_reg_45(.CP(n_62161), .D(n_453), .CD(n_61171), .Q(tsc[45])
		);
	notech_reg tsc_reg_46(.CP(n_62161), .D(n_455), .CD(n_61171), .Q(tsc[46])
		);
	notech_reg tsc_reg_47(.CP(n_62161), .D(n_457), .CD(n_61171), .Q(tsc[47])
		);
	notech_reg tsc_reg_48(.CP(n_62161), .D(n_459), .CD(n_61171), .Q(tsc[48])
		);
	notech_reg tsc_reg_49(.CP(n_62161), .D(n_461), .CD(n_61171), .Q(tsc[49])
		);
	notech_reg tsc_reg_50(.CP(n_62161), .D(n_463), .CD(n_61171), .Q(tsc[50])
		);
	notech_reg tsc_reg_51(.CP(n_62161), .D(n_465), .CD(n_61171), .Q(tsc[51])
		);
	notech_reg tsc_reg_52(.CP(n_62223), .D(n_467), .CD(n_61171), .Q(tsc[52])
		);
	notech_reg tsc_reg_53(.CP(n_62159), .D(n_469), .CD(n_61170), .Q(tsc[53])
		);
	notech_reg tsc_reg_54(.CP(n_62159), .D(n_471), .CD(n_61170), .Q(tsc[54])
		);
	notech_reg tsc_reg_55(.CP(n_62219), .D(n_473), .CD(n_61170), .Q(tsc[55])
		);
	notech_reg tsc_reg_56(.CP(n_62219), .D(n_475), .CD(n_61170), .Q(tsc[56])
		);
	notech_reg tsc_reg_57(.CP(n_62219), .D(n_477), .CD(n_61170), .Q(tsc[57])
		);
	notech_reg tsc_reg_58(.CP(n_62219), .D(n_479), .CD(n_61171), .Q(tsc[58])
		);
	notech_reg tsc_reg_59(.CP(n_62219), .D(n_481), .CD(n_61171), .Q(tsc[59])
		);
	notech_reg tsc_reg_60(.CP(n_62219), .D(n_483), .CD(n_61170), .Q(tsc[60])
		);
	notech_reg tsc_reg_61(.CP(n_62219), .D(n_485), .CD(n_61171), .Q(tsc[61])
		);
	notech_reg tsc_reg_62(.CP(n_62219), .D(n_487), .CD(n_61178), .Q(tsc[62])
		);
	notech_reg tsc_reg_63(.CP(n_62219), .D(n_489), .CD(n_61182), .Q(tsc[63])
		);
	notech_reg_set first_rep_reg(.CP(n_62219), .D(n_16752), .SD(n_61183), .Q
		(first_rep));
	notech_mux2 i_1885(.S(n_14770), .A(first_rep), .B(n_59780), .Z(n_16752)
		);
	notech_and4 i_166(.A(n_2479), .B(n_2478), .C(n_2486), .D(n_2245), .Z(n_2488
		));
	notech_reg_set fecx_reg(.CP(n_62303), .D(n_16760), .SD(1'b1), .Q(fecx)
		);
	notech_mux2 i_1894(.S(n_26631), .A(fecx), .B(n_26620), .Z(n_16760));
	notech_reg sav_ecx_reg_0(.CP(n_62303), .D(n_16767), .CD(n_61182), .Q(sav_ecx
		[0]));
	notech_mux2 i_1902(.S(n_59134), .A(ecx[0]), .B(sav_ecx[0]), .Z(n_16767)
		);
	notech_and4 i_164(.A(n_2484), .B(n_2483), .C(n_2481), .D(n_224488804), .Z
		(n_2486));
	notech_reg sav_ecx_reg_1(.CP(n_62303), .D(n_16774), .CD(n_61182), .Q(sav_ecx
		[1]));
	notech_mux2 i_1911(.S(n_59134), .A(ecx[1]), .B(sav_ecx[1]), .Z(n_16774)
		);
	notech_reg sav_ecx_reg_2(.CP(n_62303), .D(n_16781), .CD(n_61183), .Q(sav_ecx
		[2]));
	notech_mux2 i_1920(.S(n_59134), .A(ecx[2]), .B(sav_ecx[2]), .Z(n_16781)
		);
	notech_ao4 i_155(.A(n_245156269), .B(n_28517), .C(n_245756275), .D(n_28525
		), .Z(n_2484));
	notech_reg sav_ecx_reg_3(.CP(n_62303), .D(n_16788), .CD(n_61183), .Q(sav_ecx
		[3]));
	notech_mux2 i_1928(.S(n_59134), .A(ecx[3]), .B(sav_ecx[3]), .Z(n_16788)
		);
	notech_ao4 i_154(.A(n_245656274), .B(n_28533), .C(n_246156279), .D(n_28541
		), .Z(n_2483));
	notech_reg sav_ecx_reg_4(.CP(n_62303), .D(n_16796), .CD(n_61183), .Q(sav_ecx
		[4]));
	notech_mux2 i_1936(.S(n_59134), .A(ecx[4]), .B(sav_ecx[4]), .Z(n_16796)
		);
	notech_reg sav_ecx_reg_5(.CP(n_62303), .D(n_16803), .CD(n_61183), .Q(sav_ecx
		[5]));
	notech_mux2 i_1944(.S(n_59134), .A(ecx[5]), .B(sav_ecx[5]), .Z(n_16803)
		);
	notech_ao4 i_153(.A(n_246056278), .B(n_28549), .C(n_247456292), .D(n_29013
		), .Z(n_2481));
	notech_reg sav_ecx_reg_6(.CP(n_62303), .D(n_16810), .CD(n_61183), .Q(sav_ecx
		[6]));
	notech_mux2 i_1952(.S(n_59135), .A(ecx[6]), .B(sav_ecx[6]), .Z(n_16810)
		);
	notech_reg sav_ecx_reg_7(.CP(n_62303), .D(n_16817), .CD(n_61182), .Q(sav_ecx
		[7]));
	notech_mux2 i_1960(.S(n_59135), .A(ecx[7]), .B(sav_ecx[7]), .Z(n_16817)
		);
	notech_ao4 i_157(.A(n_246956287), .B(n_28556), .C(n_247556293), .D(n_29014
		), .Z(n_2479));
	notech_reg sav_ecx_reg_8(.CP(n_62303), .D(n_16824), .CD(n_61182), .Q(sav_ecx
		[8]));
	notech_mux2 i_1969(.S(n_59135), .A(ecx[8]), .B(sav_ecx[8]), .Z(n_16824)
		);
	notech_ao4 i_156(.A(n_245056268), .B(n_28501), .C(n_245256270), .D(n_28509
		), .Z(n_2478));
	notech_reg sav_ecx_reg_9(.CP(n_62303), .D(n_16832), .CD(n_61182), .Q(sav_ecx
		[9]));
	notech_mux2 i_1980(.S(n_59134), .A(ecx[9]), .B(sav_ecx[9]), .Z(n_16832)
		);
	notech_reg sav_ecx_reg_10(.CP(n_62303), .D(n_16839), .CD(n_61182), .Q(sav_ecx
		[10]));
	notech_mux2 i_1991(.S(n_59134), .A(ecx[10]), .B(sav_ecx[10]), .Z(n_16839
		));
	notech_and2 i_1179596(.A(n_247556293), .B(n_247456292), .Z(n_247656294)
		);
	notech_reg sav_ecx_reg_11(.CP(n_62303), .D(n_16846), .CD(n_61182), .Q(sav_ecx
		[11]));
	notech_mux2 i_1999(.S(n_59135), .A(ecx[11]), .B(sav_ecx[11]), .Z(n_16846
		));
	notech_nand3 i_46318(.A(vliw_pc[1]), .B(vliw_pc[0]), .C(n_246556283), .Z
		(n_247556293));
	notech_reg sav_ecx_reg_12(.CP(n_62303), .D(n_16853), .CD(n_61182), .Q(sav_ecx
		[12]));
	notech_mux2 i_2012(.S(n_59129), .A(ecx[12]), .B(sav_ecx[12]), .Z(n_16853
		));
	notech_nao3 i_46317(.A(vliw_pc[2]), .B(n_244756265), .C(n_2832), .Z(n_247456292
		));
	notech_reg sav_ecx_reg_13(.CP(n_62303), .D(n_16860), .CD(n_61182), .Q(sav_ecx
		[13]));
	notech_mux2 i_2025(.S(n_59129), .A(ecx[13]), .B(sav_ecx[13]), .Z(n_16860
		));
	notech_reg sav_ecx_reg_14(.CP(n_62303), .D(n_16868), .CD(n_61182), .Q(sav_ecx
		[14]));
	notech_mux2 i_2034(.S(n_59129), .A(ecx[14]), .B(sav_ecx[14]), .Z(n_16868
		));
	notech_and2 i_2084(.A(n_247156289), .B(n_246856286), .Z(n_247256290));
	notech_reg sav_ecx_reg_15(.CP(n_62303), .D(n_16875), .CD(n_61182), .Q(sav_ecx
		[15]));
	notech_mux2 i_2042(.S(n_59129), .A(ecx[15]), .B(sav_ecx[15]), .Z(n_16875
		));
	notech_and2 i_1479595(.A(n_247056288), .B(n_246956287), .Z(n_247156289)
		);
	notech_reg sav_ecx_reg_16(.CP(n_62303), .D(n_16882), .CD(n_61183), .Q(sav_ecx
		[16]));
	notech_mux2 i_2053(.S(n_59129), .A(ecx[16]), .B(sav_ecx[16]), .Z(n_16882
		));
	notech_nao3 i_1279594(.A(vliw_pc[1]), .B(n_246556283), .C(vliw_pc[0]), .Z
		(n_247056288));
	notech_reg sav_ecx_reg_17(.CP(n_62219), .D(n_16889), .CD(n_61186), .Q(sav_ecx
		[17]));
	notech_mux2 i_2064(.S(n_59129), .A(ecx[17]), .B(sav_ecx[17]), .Z(n_16889
		));
	notech_nao3 i_46320(.A(vliw_pc[0]), .B(n_246556283), .C(vliw_pc[1]), .Z(n_246956287
		));
	notech_reg sav_ecx_reg_18(.CP(n_62303), .D(n_16895), .CD(n_61186), .Q(sav_ecx
		[18]));
	notech_mux2 i_2072(.S(n_59134), .A(ecx[18]), .B(sav_ecx[18]), .Z(n_16895
		));
	notech_and3 i_328(.A(n_246656284), .B(n_246456282), .C(n_246356281), .Z(n_246856286
		));
	notech_reg sav_ecx_reg_19(.CP(n_62221), .D(n_16901), .CD(n_61186), .Q(sav_ecx
		[19]));
	notech_mux2 i_2085(.S(n_59134), .A(ecx[19]), .B(sav_ecx[19]), .Z(n_16901
		));
	notech_reg sav_ecx_reg_20(.CP(n_62221), .D(n_16907), .CD(n_61186), .Q(sav_ecx
		[20]));
	notech_mux2 i_2095(.S(n_59134), .A(ecx[20]), .B(sav_ecx[20]), .Z(n_16907
		));
	notech_or4 i_46321(.A(vliw_pc[0]), .B(vliw_pc[1]), .C(vliw_pc[2]), .D(n_2832
		), .Z(n_246656284));
	notech_reg sav_ecx_reg_21(.CP(n_62221), .D(n_16913), .CD(n_61186), .Q(sav_ecx
		[21]));
	notech_mux2 i_2105(.S(n_59134), .A(ecx[21]), .B(sav_ecx[21]), .Z(n_16913
		));
	notech_ao3 i_2015(.A(vliw_pc[3]), .B(n_27268), .C(vliw_pc[2]), .Z(n_246556283
		));
	notech_reg sav_ecx_reg_22(.CP(n_62221), .D(n_16919), .CD(n_61186), .Q(sav_ecx
		[22]));
	notech_mux2 i_2113(.S(n_59134), .A(ecx[22]), .B(sav_ecx[22]), .Z(n_16919
		));
	notech_nao3 i_1130932(.A(vliw_pc[2]), .B(n_244856266), .C(n_2789), .Z(n_246456282
		));
	notech_reg sav_ecx_reg_23(.CP(n_62221), .D(n_16925), .CD(n_61186), .Q(sav_ecx
		[23]));
	notech_mux2 i_2122(.S(n_59134), .A(ecx[23]), .B(sav_ecx[23]), .Z(n_16925
		));
	notech_ao3 i_2058(.A(n_246056278), .B(n_245956277), .C(n_26877), .Z(n_246356281
		));
	notech_reg sav_ecx_reg_24(.CP(n_62221), .D(n_16931), .CD(n_61186), .Q(sav_ecx
		[24]));
	notech_mux2 i_2131(.S(n_59137), .A(ecx[24]), .B(sav_ecx[24]), .Z(n_16931
		));
	notech_reg sav_ecx_reg_25(.CP(n_62221), .D(n_16937), .CD(n_61186), .Q(sav_ecx
		[25]));
	notech_mux2 i_2139(.S(n_59137), .A(ecx[25]), .B(sav_ecx[25]), .Z(n_16937
		));
	notech_nao3 i_46324(.A(vliw_pc[2]), .B(n_244856266), .C(n_54510), .Z(n_246156279
		));
	notech_reg sav_ecx_reg_26(.CP(n_62221), .D(n_16943), .CD(n_61183), .Q(sav_ecx
		[26]));
	notech_mux2 i_2148(.S(n_59137), .A(ecx[26]), .B(sav_ecx[26]), .Z(n_16943
		));
	notech_nao3 i_46323(.A(vliw_pc[2]), .B(n_244856266), .C(n_54500), .Z(n_246056278
		));
	notech_reg sav_ecx_reg_27(.CP(n_62221), .D(n_16949), .CD(n_61183), .Q(sav_ecx
		[27]));
	notech_mux2 i_2157(.S(n_59137), .A(ecx[27]), .B(sav_ecx[27]), .Z(n_16949
		));
	notech_and4 i_301(.A(n_245256270), .B(n_245156269), .C(n_245056268), .D(n_245856276
		), .Z(n_245956277));
	notech_reg sav_ecx_reg_28(.CP(n_62221), .D(n_16955), .CD(n_61183), .Q(sav_ecx
		[28]));
	notech_mux2 i_2166(.S(n_59137), .A(ecx[28]), .B(sav_ecx[28]), .Z(n_16955
		));
	notech_and2 i_20(.A(n_245756275), .B(n_245656274), .Z(n_245856276));
	notech_reg sav_ecx_reg_29(.CP(n_62221), .D(n_16961), .CD(n_61183), .Q(sav_ecx
		[29]));
	notech_mux2 i_2176(.S(n_59137), .A(ecx[29]), .B(sav_ecx[29]), .Z(n_16961
		));
	notech_or4 i_46326(.A(vliw_pc[3]), .B(vliw_pc[2]), .C(vliw_pc[4]), .D(n_2789
		), .Z(n_245756275));
	notech_reg sav_ecx_reg_30(.CP(n_62221), .D(n_16967), .CD(n_61183), .Q(sav_ecx
		[30]));
	notech_mux2 i_2185(.S(n_59137), .A(ecx[30]), .B(sav_ecx[30]), .Z(n_16967
		));
	notech_nand3 i_46325(.A(vliw_pc[2]), .B(n_244856266), .C(n_244756265), .Z
		(n_245656274));
	notech_reg sav_ecx_reg_31(.CP(n_62221), .D(n_16973), .CD(n_61186), .Q(sav_ecx
		[31]));
	notech_mux2 i_2195(.S(n_59137), .A(ecx[31]), .B(sav_ecx[31]), .Z(n_16973
		));
	notech_reg fesp_reg(.CP(n_62221), .D(n_16984), .CD(n_61186), .Q(fesp));
	notech_or4 i_2204(.A(n_60767), .B(n_60721), .C(n_55248), .D(n_9223), .Z(n_16981
		));
	notech_and4 i_2205(.A(n_54862), .B(n_42082), .C(n_206482046), .D(fesp), 
		.Z(n_16982));
	notech_nao3 i_2208(.A(n_16981), .B(1'b1), .C(n_16982), .Z(n_16984));
	notech_reg_set sav_esp_reg_0(.CP(n_62221), .D(n_16985), .SD(1'b1), .Q(sav_esp
		[0]));
	notech_mux2 i_2211(.S(n_335083325), .A(regs_4[0]), .B(sav_esp[0]), .Z(n_16985
		));
	notech_reg_set sav_esp_reg_1(.CP(n_62221), .D(n_16991), .SD(1'b1), .Q(sav_esp
		[1]));
	notech_mux2 i_2219(.S(n_335083325), .A(regs_4[1]), .B(sav_esp[1]), .Z(n_16991
		));
	notech_or4 i_46328(.A(vliw_pc[3]), .B(vliw_pc[2]), .C(vliw_pc[4]), .D(n_54510
		), .Z(n_245256270));
	notech_reg_set sav_esp_reg_2(.CP(n_62221), .D(n_16997), .SD(1'b1), .Q(sav_esp
		[2]));
	notech_mux2 i_2227(.S(n_335083325), .A(regs_4[2]), .B(sav_esp[2]), .Z(n_16997
		));
	notech_or4 i_46327(.A(vliw_pc[3]), .B(vliw_pc[2]), .C(vliw_pc[4]), .D(n_54500
		), .Z(n_245156269));
	notech_reg_set sav_esp_reg_3(.CP(n_62221), .D(n_17003), .SD(1'b1), .Q(sav_esp
		[3]));
	notech_mux2 i_2236(.S(n_335083325), .A(regs_4[3]), .B(sav_esp[3]), .Z(n_17003
		));
	notech_nao3 i_46329(.A(n_244856266), .B(n_244756265), .C(vliw_pc[2]), .Z
		(n_245056268));
	notech_reg_set sav_esp_reg_4(.CP(n_62221), .D(n_17009), .SD(1'b1), .Q(sav_esp
		[4]));
	notech_mux2 i_2244(.S(n_335083325), .A(regs_4[4]), .B(sav_esp[4]), .Z(n_17009
		));
	notech_reg_set sav_esp_reg_5(.CP(n_62159), .D(n_17016), .SD(1'b1), .Q(sav_esp
		[5]));
	notech_mux2 i_2252(.S(n_335083325), .A(regs_4[5]), .B(sav_esp[5]), .Z(n_17016
		));
	notech_nor2 i_1877(.A(vliw_pc[3]), .B(vliw_pc[4]), .Z(n_244856266));
	notech_reg_set sav_esp_reg_6(.CP(n_62159), .D(n_17022), .SD(1'b1), .Q(sav_esp
		[6]));
	notech_mux2 i_2260(.S(n_335083325), .A(regs_4[6]), .B(sav_esp[6]), .Z(n_17022
		));
	notech_nor2 i_1990(.A(vliw_pc[0]), .B(vliw_pc[1]), .Z(n_244756265));
	notech_reg_set sav_esp_reg_7(.CP(n_62159), .D(n_17028), .SD(1'b1), .Q(sav_esp
		[7]));
	notech_mux2 i_2268(.S(n_335083325), .A(regs_4[7]), .B(sav_esp[7]), .Z(n_17028
		));
	notech_nao3 i_21033193(.A(n_62395), .B(n_59375), .C(n_60494), .Z(n_244656264
		));
	notech_reg_set sav_esp_reg_8(.CP(n_62159), .D(n_17034), .SD(1'b1), .Q(sav_esp
		[8]));
	notech_mux2 i_2276(.S(n_335083325), .A(regs_4[8]), .B(sav_esp[8]), .Z(n_17034
		));
	notech_and2 i_2077(.A(n_60739), .B(n_27265), .Z(n_244556263));
	notech_reg_set sav_esp_reg_9(.CP(n_62159), .D(n_17040), .SD(1'b1), .Q(sav_esp
		[9]));
	notech_mux2 i_2284(.S(n_335083325), .A(regs_4[9]), .B(sav_esp[9]), .Z(n_17040
		));
	notech_reg_set sav_esp_reg_10(.CP(n_62159), .D(n_17046), .SD(1'b1), .Q(sav_esp
		[10]));
	notech_mux2 i_2292(.S(n_335083325), .A(regs_4[10]), .B(sav_esp[10]), .Z(n_17046
		));
	notech_and2 i_16844(.A(fsm[2]), .B(n_27266), .Z(n_244356261));
	notech_reg_set sav_esp_reg_11(.CP(n_62159), .D(n_17052), .SD(1'b1), .Q(sav_esp
		[11]));
	notech_mux2 i_2300(.S(n_335083325), .A(regs_4[11]), .B(sav_esp[11]), .Z(n_17052
		));
	notech_nand2 i_1919(.A(n_27265), .B(n_27262), .Z(n_244256260));
	notech_reg_set sav_esp_reg_12(.CP(n_62159), .D(n_17058), .SD(1'b1), .Q(sav_esp
		[12]));
	notech_mux2 i_2308(.S(n_335083325), .A(regs_4[12]), .B(sav_esp[12]), .Z(n_17058
		));
	notech_reg_set sav_esp_reg_13(.CP(n_62159), .D(n_17064), .SD(1'b1), .Q(sav_esp
		[13]));
	notech_mux2 i_2316(.S(n_335083325), .A(regs_4[13]), .B(sav_esp[13]), .Z(n_17064
		));
	notech_and3 i_2021(.A(n_60752), .B(n_27262), .C(n_27264), .Z(n_244056258
		));
	notech_reg_set sav_esp_reg_14(.CP(n_62159), .D(n_17070), .SD(1'b1), .Q(sav_esp
		[14]));
	notech_mux2 i_2324(.S(n_335083325), .A(regs_4[14]), .B(sav_esp[14]), .Z(n_17070
		));
	notech_reg_set sav_esp_reg_15(.CP(n_62219), .D(n_17076), .SD(1'b1), .Q(sav_esp
		[15]));
	notech_mux2 i_2332(.S(n_335083325), .A(regs_4[15]), .B(sav_esp[15]), .Z(n_17076
		));
	notech_nand3 i_1417400(.A(n_2644), .B(n_243656254), .C(n_2642), .Z(n_17274
		));
	notech_reg_set sav_esp_reg_16(.CP(n_62213), .D(n_17082), .SD(1'b1), .Q(sav_esp
		[16]));
	notech_mux2 i_2340(.S(n_53630), .A(regs_4[16]), .B(sav_esp[16]), .Z(n_17082
		));
	notech_reg_set sav_esp_reg_17(.CP(n_62157), .D(n_17088), .SD(1'b1), .Q(sav_esp
		[17]));
	notech_mux2 i_2348(.S(n_53630), .A(regs_4[17]), .B(sav_esp[17]), .Z(n_17088
		));
	notech_reg_set sav_esp_reg_18(.CP(n_62213), .D(n_17094), .SD(1'b1), .Q(sav_esp
		[18]));
	notech_mux2 i_2356(.S(n_53630), .A(regs_4[18]), .B(sav_esp[18]), .Z(n_17094
		));
	notech_nand2 i_866(.A(resa_shiftbox[13]), .B(n_26288), .Z(n_243656254)
		);
	notech_reg_set sav_esp_reg_19(.CP(n_62213), .D(n_17100), .SD(1'b1), .Q(sav_esp
		[19]));
	notech_mux2 i_2364(.S(n_53630), .A(regs_4[19]), .B(sav_esp[19]), .Z(n_17100
		));
	notech_or2 i_879(.A(n_56952), .B(n_55552), .Z(n_243556253));
	notech_reg_set sav_esp_reg_20(.CP(n_62213), .D(n_17106), .SD(1'b1), .Q(sav_esp
		[20]));
	notech_mux2 i_2372(.S(n_53630), .A(regs_4[20]), .B(sav_esp[20]), .Z(n_17106
		));
	notech_or4 i_871(.A(n_2610), .B(n_273188724), .C(n_59899), .D(n_27566), 
		.Z(n_243456252));
	notech_reg_set sav_esp_reg_21(.CP(n_62213), .D(n_17112), .SD(1'b1), .Q(sav_esp
		[21]));
	notech_mux2 i_2380(.S(n_53630), .A(regs_4[21]), .B(sav_esp[21]), .Z(n_17112
		));
	notech_nao3 i_893(.A(n_57438), .B(nbus_140[13]), .C(n_2833), .Z(n_243356251
		));
	notech_reg_set sav_esp_reg_22(.CP(n_62213), .D(n_17118), .SD(1'b1), .Q(sav_esp
		[22]));
	notech_mux2 i_2388(.S(n_53630), .A(regs_4[22]), .B(sav_esp[22]), .Z(n_17118
		));
	notech_or4 i_892(.A(n_260988754), .B(n_260888755), .C(n_2833), .D(n_28281
		), .Z(n_243256250));
	notech_reg_set sav_esp_reg_23(.CP(n_62213), .D(n_17124), .SD(1'b1), .Q(sav_esp
		[23]));
	notech_mux2 i_2397(.S(n_53630), .A(regs_4[23]), .B(sav_esp[23]), .Z(n_17124
		));
	notech_nao3 i_891(.A(n_57438), .B(nbus_142[13]), .C(n_2834), .Z(n_243156249
		));
	notech_reg_set sav_esp_reg_24(.CP(n_62213), .D(n_17130), .SD(1'b1), .Q(sav_esp
		[24]));
	notech_mux2 i_2405(.S(n_53630), .A(regs_4[24]), .B(sav_esp[24]), .Z(n_17130
		));
	notech_reg_set sav_esp_reg_25(.CP(n_62213), .D(n_17136), .SD(1'b1), .Q(sav_esp
		[25]));
	notech_mux2 i_2413(.S(n_53630), .A(regs_4[25]), .B(sav_esp[25]), .Z(n_17136
		));
	notech_reg_set sav_esp_reg_26(.CP(n_62213), .D(n_17142), .SD(1'b1), .Q(sav_esp
		[26]));
	notech_mux2 i_2421(.S(n_53630), .A(regs_4[26]), .B(sav_esp[26]), .Z(n_17142
		));
	notech_reg_set sav_esp_reg_27(.CP(n_62213), .D(n_17148), .SD(1'b1), .Q(sav_esp
		[27]));
	notech_mux2 i_2429(.S(n_53630), .A(regs_4[27]), .B(sav_esp[27]), .Z(n_17148
		));
	notech_reg_set sav_esp_reg_28(.CP(n_62299), .D(n_17154), .SD(1'b1), .Q(sav_esp
		[28]));
	notech_mux2 i_2437(.S(n_53630), .A(regs_4[28]), .B(sav_esp[28]), .Z(n_17154
		));
	notech_or4 i_873(.A(n_60767), .B(n_60724), .C(n_57390), .D(n_56685), .Z(n_242656244
		));
	notech_reg_set sav_esp_reg_29(.CP(n_62299), .D(n_17160), .SD(1'b1), .Q(sav_esp
		[29]));
	notech_mux2 i_2445(.S(n_53630), .A(regs_4[29]), .B(sav_esp[29]), .Z(n_17160
		));
	notech_reg_set sav_esp_reg_30(.CP(n_62299), .D(n_17166), .SD(1'b1), .Q(sav_esp
		[30]));
	notech_mux2 i_2453(.S(n_53630), .A(regs_4[30]), .B(sav_esp[30]), .Z(n_17166
		));
	notech_reg_set sav_esp_reg_31(.CP(n_62299), .D(n_17172), .SD(1'b1), .Q(sav_esp
		[31]));
	notech_mux2 i_2461(.S(n_53630), .A(regs_4[31]), .B(sav_esp[31]), .Z(n_17172
		));
	notech_reg sav_esi_reg_0(.CP(n_62299), .D(n_17178), .CD(n_61183), .Q(sav_esi
		[0]));
	notech_mux2 i_2470(.S(n_59137), .A(regs_6[0]), .B(sav_esi[0]), .Z(n_17178
		));
	notech_reg sav_esi_reg_1(.CP(n_62299), .D(n_17184), .CD(n_61186), .Q(sav_esi
		[1]));
	notech_mux2 i_2478(.S(n_59137), .A(regs_6[1]), .B(sav_esi[1]), .Z(n_17184
		));
	notech_reg sav_esi_reg_2(.CP(n_62299), .D(n_17190), .CD(n_61182), .Q(sav_esi
		[2]));
	notech_mux2 i_2486(.S(n_59137), .A(regs_6[2]), .B(sav_esi[2]), .Z(n_17190
		));
	notech_reg sav_esi_reg_3(.CP(n_62299), .D(n_17197), .CD(n_61180), .Q(sav_esi
		[3]));
	notech_mux2 i_2494(.S(n_59137), .A(regs_6[3]), .B(sav_esi[3]), .Z(n_17197
		));
	notech_or2 i_894(.A(n_2820), .B(n_55249), .Z(n_241956237));
	notech_reg sav_esi_reg_4(.CP(n_62299), .D(n_17204), .CD(n_61180), .Q(sav_esi
		[4]));
	notech_mux2 i_2503(.S(n_59135), .A(regs_6[4]), .B(sav_esi[4]), .Z(n_17204
		));
	notech_nao3 i_888(.A(n_26650), .B(opa_0[13]), .C(n_57438), .Z(n_241856236
		));
	notech_reg sav_esi_reg_5(.CP(n_62299), .D(n_17211), .CD(n_61178), .Q(sav_esi
		[5]));
	notech_mux2 i_2511(.S(n_59135), .A(regs_6[5]), .B(sav_esi[5]), .Z(n_17211
		));
	notech_reg sav_esi_reg_6(.CP(n_62299), .D(n_17218), .CD(n_61178), .Q(sav_esi
		[6]));
	notech_mux2 i_2519(.S(n_59135), .A(regs_6[6]), .B(sav_esi[6]), .Z(n_17218
		));
	notech_reg sav_esi_reg_7(.CP(n_62299), .D(n_17225), .CD(n_61180), .Q(sav_esi
		[7]));
	notech_mux2 i_2527(.S(n_59135), .A(regs_6[7]), .B(sav_esi[7]), .Z(n_17225
		));
	notech_nao3 i_870(.A(resa_arithbox[13]), .B(n_59819), .C(n_57424), .Z(n_241556233
		));
	notech_reg sav_esi_reg_8(.CP(n_62299), .D(n_17233), .CD(n_61180), .Q(sav_esi
		[8]));
	notech_mux2 i_2535(.S(n_59135), .A(regs_6[8]), .B(sav_esi[8]), .Z(n_17233
		));
	notech_nao3 i_883(.A(resa_shift4box[13]), .B(n_26856), .C(n_275988698), 
		.Z(n_241456232));
	notech_reg sav_esi_reg_9(.CP(n_62299), .D(n_17240), .CD(n_61180), .Q(sav_esi
		[9]));
	notech_mux2 i_2543(.S(n_59135), .A(regs_6[9]), .B(sav_esi[9]), .Z(n_17240
		));
	notech_or2 i_867(.A(n_57298), .B(n_29037), .Z(n_2413));
	notech_reg sav_esi_reg_10(.CP(n_62299), .D(n_17247), .CD(n_61180), .Q(sav_esi
		[10]));
	notech_mux2 i_2551(.S(n_59135), .A(regs_6[10]), .B(sav_esi[10]), .Z(n_17247
		));
	notech_nand2 i_868(.A(readio_data[13]), .B(n_26287), .Z(n_241288763));
	notech_reg sav_esi_reg_11(.CP(n_62299), .D(n_17254), .CD(n_61180), .Q(sav_esi
		[11]));
	notech_mux2 i_2559(.S(n_59137), .A(regs_6[11]), .B(sav_esi[11]), .Z(n_17254
		));
	notech_reg sav_esi_reg_12(.CP(n_62299), .D(n_17261), .CD(n_61178), .Q(sav_esi
		[12]));
	notech_mux2 i_2567(.S(n_59137), .A(regs_6[12]), .B(sav_esi[12]), .Z(n_17261
		));
	notech_reg sav_esi_reg_13(.CP(n_62299), .D(n_17269), .CD(n_61178), .Q(sav_esi
		[13]));
	notech_mux2 i_2575(.S(n_59135), .A(regs_6[13]), .B(sav_esi[13]), .Z(n_17269
		));
	notech_ao4 i_127(.A(n_2390), .B(n_59899), .C(n_2799), .D(nbus_11279[13])
		, .Z(n_2409));
	notech_reg sav_esi_reg_14(.CP(n_62299), .D(n_17276), .CD(n_61178), .Q(sav_esi
		[14]));
	notech_mux2 i_2583(.S(n_59135), .A(regs_6[14]), .B(sav_esi[14]), .Z(n_17276
		));
	notech_reg sav_esi_reg_15(.CP(n_62363), .D(n_17283), .CD(n_61178), .Q(sav_esi
		[15]));
	notech_mux2 i_2591(.S(n_59135), .A(regs_6[15]), .B(sav_esi[15]), .Z(n_17283
		));
	notech_and3 i_130(.A(n_2822), .B(n_2823), .C(n_2824), .Z(n_2407));
	notech_reg sav_esi_reg_16(.CP(n_62297), .D(n_17290), .CD(n_61178), .Q(sav_esi
		[16]));
	notech_mux2 i_2599(.S(n_59129), .A(regs_6[16]), .B(sav_esi[16]), .Z(n_17290
		));
	notech_or4 i_523(.A(n_2793), .B(n_59771), .C(n_59159), .D(n_2407), .Z(n_2406
		));
	notech_reg sav_esi_reg_17(.CP(n_62363), .D(n_17297), .CD(n_61178), .Q(sav_esi
		[17]));
	notech_mux2 i_2607(.S(n_59122), .A(regs_6[17]), .B(sav_esi[17]), .Z(n_17297
		));
	notech_ao4 i_586(.A(n_494), .B(n_55641), .C(n_57445), .D(n_59150), .Z(n_55763
		));
	notech_reg sav_esi_reg_18(.CP(n_62363), .D(n_17305), .CD(n_61178), .Q(sav_esi
		[18]));
	notech_mux2 i_2615(.S(n_59122), .A(regs_6[18]), .B(sav_esi[18]), .Z(n_17305
		));
	notech_reg sav_esi_reg_19(.CP(n_62363), .D(n_17312), .CD(n_61178), .Q(sav_esi
		[19]));
	notech_mux2 i_2623(.S(n_59122), .A(regs_6[19]), .B(sav_esi[19]), .Z(n_17312
		));
	notech_reg sav_esi_reg_20(.CP(n_62363), .D(n_17319), .CD(n_61178), .Q(sav_esi
		[20]));
	notech_mux2 i_2631(.S(n_59122), .A(regs_6[20]), .B(sav_esi[20]), .Z(n_17319
		));
	notech_reg sav_esi_reg_21(.CP(n_62363), .D(n_17326), .CD(n_61180), .Q(sav_esi
		[21]));
	notech_mux2 i_2639(.S(n_59122), .A(regs_6[21]), .B(sav_esi[21]), .Z(n_17326
		));
	notech_reg sav_esi_reg_22(.CP(n_62363), .D(n_17333), .CD(n_61181), .Q(sav_esi
		[22]));
	notech_mux2 i_2647(.S(n_59122), .A(regs_6[22]), .B(sav_esi[22]), .Z(n_17333
		));
	notech_or4 i_1686(.A(n_2793), .B(n_59771), .C(n_59159), .D(n_57441), .Z(n_54770
		));
	notech_reg sav_esi_reg_23(.CP(n_62363), .D(n_17341), .CD(n_61181), .Q(sav_esi
		[23]));
	notech_mux2 i_2655(.S(n_59135), .A(regs_6[23]), .B(sav_esi[23]), .Z(n_17341
		));
	notech_ao4 i_511(.A(n_106813462), .B(n_2616), .C(n_58895), .D(n_58940), 
		.Z(n_55838));
	notech_reg sav_esi_reg_24(.CP(n_62363), .D(n_17348), .CD(n_61181), .Q(sav_esi
		[24]));
	notech_mux2 i_2663(.S(n_59135), .A(regs_6[24]), .B(sav_esi[24]), .Z(n_17348
		));
	notech_reg sav_esi_reg_25(.CP(n_62363), .D(n_17355), .CD(n_61181), .Q(sav_esi
		[25]));
	notech_mux2 i_2671(.S(n_59135), .A(regs_6[25]), .B(sav_esi[25]), .Z(n_17355
		));
	notech_reg sav_esi_reg_26(.CP(n_62363), .D(n_17362), .CD(n_61181), .Q(sav_esi
		[26]));
	notech_mux2 i_2679(.S(n_59135), .A(regs_6[26]), .B(sav_esi[26]), .Z(n_17362
		));
	notech_or4 i_1810(.A(n_58913), .B(n_59967), .C(n_58940), .D(n_59355), .Z
		(n_57392));
	notech_reg sav_esi_reg_27(.CP(n_62363), .D(n_17369), .CD(n_61181), .Q(sav_esi
		[27]));
	notech_mux2 i_2687(.S(n_59135), .A(regs_6[27]), .B(sav_esi[27]), .Z(n_17369
		));
	notech_or4 i_1766(.A(n_59210), .B(n_2588), .C(n_60558), .D(\opcode[1] ),
		 .Z(n_57397));
	notech_reg sav_esi_reg_28(.CP(n_62363), .D(n_17377), .CD(n_61181), .Q(sav_esi
		[28]));
	notech_mux2 i_2695(.S(n_59135), .A(regs_6[28]), .B(sav_esi[28]), .Z(n_17377
		));
	notech_nand2 i_1220(.A(n_2776), .B(n_57384), .Z(n_55154));
	notech_reg sav_esi_reg_29(.CP(n_62363), .D(n_17384), .CD(n_61181), .Q(sav_esi
		[29]));
	notech_mux2 i_2703(.S(n_59122), .A(regs_6[29]), .B(sav_esi[29]), .Z(n_17384
		));
	notech_or4 i_1759(.A(n_59210), .B(n_2588), .C(\opcode[0] ), .D(\opcode[1] 
		), .Z(n_57398));
	notech_reg sav_esi_reg_30(.CP(n_62363), .D(n_17390), .CD(n_61181), .Q(sav_esi
		[30]));
	notech_mux2 i_2711(.S(n_59122), .A(regs_6[30]), .B(sav_esi[30]), .Z(n_17390
		));
	notech_or2 i_92232881(.A(n_2361), .B(n_2385), .Z(n_2399));
	notech_reg sav_esi_reg_31(.CP(n_62363), .D(n_17396), .CD(n_61180), .Q(sav_esi
		[31]));
	notech_mux2 i_2719(.S(n_59122), .A(regs_6[31]), .B(sav_esi[31]), .Z(n_17396
		));
	notech_reg sav_edi_reg_0(.CP(n_62363), .D(n_17402), .CD(n_61180), .Q(sav_edi
		[0]));
	notech_mux2 i_2727(.S(n_59122), .A(regs_7[0]), .B(sav_edi[0]), .Z(n_17402
		));
	notech_or4 i_1843(.A(n_58913), .B(n_59967), .C(n_273288723), .D(n_59201)
		, .Z(n_57390));
	notech_reg sav_edi_reg_1(.CP(n_62363), .D(n_17408), .CD(n_61180), .Q(sav_edi
		[1]));
	notech_mux2 i_2735(.S(n_59122), .A(regs_7[1]), .B(sav_edi[1]), .Z(n_17408
		));
	notech_reg sav_edi_reg_2(.CP(n_62363), .D(n_17414), .CD(n_61180), .Q(sav_edi
		[2]));
	notech_mux2 i_2743(.S(n_59122), .A(regs_7[2]), .B(sav_edi[2]), .Z(n_17414
		));
	notech_or4 i_1678(.A(n_60494), .B(n_58904), .C(n_60558), .D(n_59375), .Z
		(n_54777));
	notech_reg sav_edi_reg_3(.CP(n_62297), .D(n_17420), .CD(n_61180), .Q(sav_edi
		[3]));
	notech_mux2 i_2751(.S(n_59122), .A(regs_7[3]), .B(sav_edi[3]), .Z(n_17420
		));
	notech_or4 i_1531(.A(n_60490), .B(n_58904), .C(\opcode[0] ), .D(\opcode[1] 
		), .Z(n_54899));
	notech_reg sav_edi_reg_4(.CP(n_62297), .D(n_17426), .CD(n_61181), .Q(sav_edi
		[4]));
	notech_mux2 i_2759(.S(n_59122), .A(regs_7[4]), .B(sav_edi[4]), .Z(n_17426
		));
	notech_reg sav_edi_reg_5(.CP(n_62297), .D(n_17432), .CD(n_61181), .Q(sav_edi
		[5]));
	notech_mux2 i_2767(.S(n_59122), .A(regs_7[5]), .B(sav_edi[5]), .Z(n_17432
		));
	notech_reg sav_edi_reg_6(.CP(n_62297), .D(n_17438), .CD(n_61181), .Q(sav_edi
		[6]));
	notech_mux2 i_2775(.S(n_59122), .A(regs_7[6]), .B(sav_edi[6]), .Z(n_17438
		));
	notech_reg sav_edi_reg_7(.CP(n_62297), .D(n_17444), .CD(n_61181), .Q(sav_edi
		[7]));
	notech_mux2 i_2783(.S(n_59122), .A(regs_7[7]), .B(sav_edi[7]), .Z(n_17444
		));
	notech_or4 i_459(.A(n_59355), .B(n_2647), .C(\opcode[0] ), .D(\opcode[1] 
		), .Z(n_2395));
	notech_reg sav_edi_reg_8(.CP(n_62297), .D(n_17450), .CD(n_61169), .Q(sav_edi
		[8]));
	notech_mux2 i_2791(.S(n_59122), .A(regs_7[8]), .B(sav_edi[8]), .Z(n_17450
		));
	notech_or4 i_1784(.A(n_62395), .B(\opcode[1] ), .C(n_60540), .D(n_62405)
		, .Z(n_54689));
	notech_reg sav_edi_reg_9(.CP(n_62297), .D(n_17456), .CD(n_61158), .Q(sav_edi
		[9]));
	notech_mux2 i_2799(.S(n_59129), .A(regs_7[9]), .B(sav_edi[9]), .Z(n_17456
		));
	notech_or4 i_454(.A(n_60540), .B(n_275488703), .C(n_60504), .D(n_2586), 
		.Z(n_2394));
	notech_reg sav_edi_reg_10(.CP(n_62297), .D(n_17462), .CD(n_61158), .Q(sav_edi
		[10]));
	notech_mux2 i_2807(.S(n_59129), .A(regs_7[10]), .B(sav_edi[10]), .Z(n_17462
		));
	notech_ao4 i_828(.A(n_272688729), .B(n_59210), .C(n_274588712), .D(n_2826
		), .Z(n_55525));
	notech_reg sav_edi_reg_11(.CP(n_62297), .D(n_17468), .CD(n_61158), .Q(sav_edi
		[11]));
	notech_mux2 i_2815(.S(n_59129), .A(regs_7[11]), .B(sav_edi[11]), .Z(n_17468
		));
	notech_reg sav_edi_reg_12(.CP(n_62297), .D(n_17474), .CD(n_61158), .Q(sav_edi
		[12]));
	notech_mux2 i_2823(.S(n_59129), .A(regs_7[12]), .B(sav_edi[12]), .Z(n_17474
		));
	notech_reg sav_edi_reg_13(.CP(n_62297), .D(n_17480), .CD(n_61158), .Q(sav_edi
		[13]));
	notech_mux2 i_2831(.S(n_59129), .A(regs_7[13]), .B(sav_edi[13]), .Z(n_17480
		));
	notech_reg sav_edi_reg_14(.CP(n_62213), .D(n_17486), .CD(n_61158), .Q(sav_edi
		[14]));
	notech_mux2 i_2839(.S(n_59129), .A(regs_7[14]), .B(sav_edi[14]), .Z(n_17486
		));
	notech_or2 i_1742(.A(n_2386), .B(n_273288723), .Z(n_57400));
	notech_reg sav_edi_reg_15(.CP(n_62157), .D(n_17492), .CD(n_61158), .Q(sav_edi
		[15]));
	notech_mux2 i_2847(.S(n_59129), .A(regs_7[15]), .B(sav_edi[15]), .Z(n_17492
		));
	notech_and3 i_426(.A(n_57400), .B(n_272888727), .C(n_2787), .Z(n_2390)
		);
	notech_reg sav_edi_reg_16(.CP(n_62301), .D(n_17498), .CD(n_61158), .Q(sav_edi
		[16]));
	notech_mux2 i_2855(.S(n_59129), .A(regs_7[16]), .B(sav_edi[16]), .Z(n_17498
		));
	notech_reg sav_edi_reg_17(.CP(n_62215), .D(n_17504), .CD(n_61158), .Q(sav_edi
		[17]));
	notech_mux2 i_2863(.S(n_59129), .A(regs_7[17]), .B(sav_edi[17]), .Z(n_17504
		));
	notech_ao4 i_416(.A(n_26865), .B(n_2586), .C(n_274488713), .D(\opcode[1] 
		), .Z(n_2388));
	notech_reg sav_edi_reg_18(.CP(n_62215), .D(n_17510), .CD(n_61157), .Q(sav_edi
		[18]));
	notech_mux2 i_2871(.S(n_59129), .A(regs_7[18]), .B(sav_edi[18]), .Z(n_17510
		));
	notech_or4 i_1178(.A(n_60752), .B(n_60739), .C(n_60768), .D(n_57423), .Z
		(n_55195));
	notech_reg sav_edi_reg_19(.CP(n_62215), .D(n_17516), .CD(n_61157), .Q(sav_edi
		[19]));
	notech_mux2 i_2879(.S(n_59129), .A(regs_7[19]), .B(sav_edi[19]), .Z(n_17516
		));
	notech_or2 i_394(.A(n_2386), .B(n_26865), .Z(n_2387));
	notech_reg sav_edi_reg_20(.CP(n_62215), .D(n_17522), .CD(n_61157), .Q(sav_edi
		[20]));
	notech_mux2 i_2887(.S(n_59129), .A(regs_7[20]), .B(sav_edi[20]), .Z(n_17522
		));
	notech_or4 i_29516(.A(n_60490), .B(\opcode[0] ), .C(\opcode[1] ), .D(n_2399
		), .Z(n_2386));
	notech_reg sav_edi_reg_21(.CP(n_62215), .D(n_17528), .CD(n_61157), .Q(sav_edi
		[21]));
	notech_mux2 i_2895(.S(n_59134), .A(regs_7[21]), .B(sav_edi[21]), .Z(n_17528
		));
	notech_nand2 i_1215(.A(n_2775), .B(n_2774), .Z(n_55159));
	notech_reg sav_edi_reg_22(.CP(n_62215), .D(n_17534), .CD(n_61157), .Q(sav_edi
		[22]));
	notech_mux2 i_2903(.S(n_59134), .A(regs_7[22]), .B(sav_edi[22]), .Z(n_17534
		));
	notech_and2 i_97470268(.A(n_2768), .B(n_2769), .Z(n_55389));
	notech_reg sav_edi_reg_23(.CP(n_62215), .D(n_17540), .CD(n_61157), .Q(sav_edi
		[23]));
	notech_mux2 i_2911(.S(n_59134), .A(regs_7[23]), .B(sav_edi[23]), .Z(n_17540
		));
	notech_and4 i_727967(.A(n_2569), .B(n_2568), .C(n_2567), .D(n_2377), .Z(n_2385
		));
	notech_reg sav_edi_reg_24(.CP(n_62215), .D(n_17546), .CD(n_61157), .Q(sav_edi
		[24]));
	notech_mux2 i_2919(.S(n_59134), .A(regs_7[24]), .B(sav_edi[24]), .Z(n_17546
		));
	notech_reg sav_edi_reg_25(.CP(n_62215), .D(n_17552), .CD(n_61157), .Q(sav_edi
		[25]));
	notech_mux2 i_2927(.S(n_59134), .A(regs_7[25]), .B(sav_edi[25]), .Z(n_17552
		));
	notech_reg sav_edi_reg_26(.CP(n_62215), .D(n_17558), .CD(n_61157), .Q(sav_edi
		[26]));
	notech_mux2 i_2935(.S(n_59134), .A(regs_7[26]), .B(sav_edi[26]), .Z(n_17558
		));
	notech_reg sav_edi_reg_27(.CP(n_62301), .D(n_17564), .CD(n_61158), .Q(sav_edi
		[27]));
	notech_mux2 i_2943(.S(n_59137), .A(regs_7[27]), .B(sav_edi[27]), .Z(n_17564
		));
	notech_reg sav_edi_reg_28(.CP(n_62301), .D(n_17570), .CD(n_61159), .Q(sav_edi
		[28]));
	notech_mux2 i_2951(.S(n_59137), .A(regs_7[28]), .B(sav_edi[28]), .Z(n_17570
		));
	notech_reg sav_edi_reg_29(.CP(n_62301), .D(n_17576), .CD(n_61159), .Q(sav_edi
		[29]));
	notech_mux2 i_2959(.S(n_59137), .A(regs_7[29]), .B(sav_edi[29]), .Z(n_17576
		));
	notech_reg sav_edi_reg_30(.CP(n_62301), .D(n_17582), .CD(n_61159), .Q(sav_edi
		[30]));
	notech_mux2 i_2967(.S(n_59137), .A(regs_7[30]), .B(sav_edi[30]), .Z(n_17582
		));
	notech_mux2 i_113(.S(n_246056278), .A(instrc[54]), .B(n_2376), .Z(n_2378
		));
	notech_reg sav_edi_reg_31(.CP(n_62301), .D(n_17588), .CD(n_61159), .Q(sav_edi
		[31]));
	notech_mux2 i_2975(.S(n_59137), .A(regs_7[31]), .B(sav_edi[31]), .Z(n_17588
		));
	notech_nao3 i_375(.A(n_245956277), .B(n_2378), .C(n_26877), .Z(n_2377)
		);
	notech_reg fepc_reg(.CP(n_62301), .D(n_17594), .CD(n_61159), .Q(fepc));
	notech_mux2 i_2983(.S(n_10174), .A(fepc), .B(n_10177), .Z(n_17594));
	notech_mux2 i_104(.S(n_246456282), .A(instrc[62]), .B(n_2373), .Z(n_2376
		));
	notech_reg_set sav_epc_reg_0(.CP(n_62301), .D(n_17600), .SD(1'b1), .Q(sav_epc
		[0]));
	notech_mux2 i_2991(.S(n_26800), .A(sav_epc[0]), .B(regs_14[0]), .Z(n_17600
		));
	notech_reg_set sav_epc_reg_1(.CP(n_62301), .D(n_17606), .SD(1'b1), .Q(sav_epc
		[1]));
	notech_mux2 i_2999(.S(n_26800), .A(sav_epc[1]), .B(regs_14[1]), .Z(n_17606
		));
	notech_reg_set sav_epc_reg_2(.CP(n_62301), .D(n_17612), .SD(1'b1), .Q(sav_epc
		[2]));
	notech_mux2 i_3007(.S(n_26800), .A(sav_epc[2]), .B(regs_14[2]), .Z(n_17612
		));
	notech_mux2 i_95(.S(n_246656284), .A(instrc[70]), .B(n_2565), .Z(n_2373)
		);
	notech_reg_set sav_epc_reg_3(.CP(n_62301), .D(n_17618), .SD(1'b1), .Q(sav_epc
		[3]));
	notech_mux2 i_3015(.S(n_26800), .A(sav_epc[3]), .B(regs_14[3]), .Z(n_17618
		));
	notech_reg_set sav_epc_reg_4(.CP(n_62301), .D(n_17624), .SD(1'b1), .Q(sav_epc
		[4]));
	notech_mux2 i_3023(.S(n_26800), .A(sav_epc[4]), .B(regs_14[4]), .Z(n_17624
		));
	notech_reg_set sav_epc_reg_5(.CP(n_62301), .D(n_17630), .SD(1'b1), .Q(sav_epc
		[5]));
	notech_mux2 i_3031(.S(n_26800), .A(sav_epc[5]), .B(regs_14[5]), .Z(n_17630
		));
	notech_reg_set sav_epc_reg_6(.CP(n_62301), .D(n_17636), .SD(1'b1), .Q(sav_epc
		[6]));
	notech_mux2 i_3039(.S(n_26800), .A(sav_epc[6]), .B(regs_14[6]), .Z(n_17636
		));
	notech_reg_set sav_epc_reg_7(.CP(n_62301), .D(n_17642), .SD(1'b1), .Q(sav_epc
		[7]));
	notech_mux2 i_3047(.S(n_26800), .A(sav_epc[7]), .B(regs_14[7]), .Z(n_17642
		));
	notech_reg_set sav_epc_reg_8(.CP(n_62301), .D(n_17648), .SD(1'b1), .Q(sav_epc
		[8]));
	notech_mux2 i_3055(.S(n_26800), .A(sav_epc[8]), .B(regs_14[8]), .Z(n_17648
		));
	notech_reg_set sav_epc_reg_9(.CP(n_62301), .D(n_17654), .SD(1'b1), .Q(sav_epc
		[9]));
	notech_mux2 i_3063(.S(n_26800), .A(sav_epc[9]), .B(regs_14[9]), .Z(n_17654
		));
	notech_nand2 i_131(.A(n_2563), .B(n_2362), .Z(n_2366));
	notech_reg_set sav_epc_reg_10(.CP(n_62301), .D(n_17662), .SD(1'b1), .Q(sav_epc
		[10]));
	notech_mux2 i_3071(.S(n_26800), .A(sav_epc[10]), .B(regs_14[10]), .Z(n_17662
		));
	notech_nand2 i_361(.A(n_247156289), .B(n_2366), .Z(n_2365));
	notech_reg_set sav_epc_reg_11(.CP(n_62301), .D(n_17668), .SD(1'b1), .Q(sav_epc
		[11]));
	notech_mux2 i_3079(.S(n_26800), .A(sav_epc[11]), .B(regs_14[11]), .Z(n_17668
		));
	notech_reg_set sav_epc_reg_12(.CP(n_62215), .D(n_17674), .SD(1'b1), .Q(sav_epc
		[12]));
	notech_mux2 i_3087(.S(n_26800), .A(sav_epc[12]), .B(regs_14[12]), .Z(n_17674
		));
	notech_reg_set sav_epc_reg_13(.CP(n_62215), .D(n_17681), .SD(1'b1), .Q(sav_epc
		[13]));
	notech_mux2 i_3095(.S(n_26800), .A(sav_epc[13]), .B(regs_14[13]), .Z(n_17681
		));
	notech_nand2 i_357(.A(n_247656294), .B(n_28970), .Z(n_2362));
	notech_reg_set sav_epc_reg_14(.CP(n_62217), .D(n_17687), .SD(1'b1), .Q(sav_epc
		[14]));
	notech_mux2 i_3103(.S(n_26800), .A(sav_epc[14]), .B(regs_14[14]), .Z(n_17687
		));
	notech_nor2 i_527965(.A(n_2341), .B(n_2562), .Z(n_2361));
	notech_reg_set sav_epc_reg_15(.CP(n_62217), .D(n_17693), .SD(1'b1), .Q(sav_epc
		[15]));
	notech_mux2 i_3111(.S(n_26800), .A(sav_epc[15]), .B(regs_14[15]), .Z(n_17693
		));
	notech_ao3 i_326(.A(n_244856266), .B(instrc[60]), .C(n_2790), .Z(n_2360)
		);
	notech_reg_set sav_epc_reg_16(.CP(n_62217), .D(n_17700), .SD(1'b1), .Q(sav_epc
		[16]));
	notech_mux2 i_3119(.S(n_53833), .A(sav_epc[16]), .B(regs_14[16]), .Z(n_17700
		));
	notech_or2 i_341(.A(n_247056288), .B(n_29035), .Z(n_235988764));
	notech_reg_set sav_epc_reg_17(.CP(n_62217), .D(n_17708), .SD(1'b1), .Q(sav_epc
		[17]));
	notech_mux2 i_3127(.S(n_53833), .A(sav_epc[17]), .B(regs_14[17]), .Z(n_17708
		));
	notech_nand3 i_333(.A(n_244756265), .B(n_246556283), .C(instrc[68]), .Z(n_2358
		));
	notech_reg_set sav_epc_reg_18(.CP(n_62217), .D(n_17715), .SD(1'b1), .Q(sav_epc
		[18]));
	notech_mux2 i_3135(.S(n_53833), .A(sav_epc[18]), .B(regs_14[18]), .Z(n_17715
		));
	notech_reg_set sav_epc_reg_19(.CP(n_62217), .D(n_17723), .SD(1'b1), .Q(sav_epc
		[19]));
	notech_mux2 i_3143(.S(n_53833), .A(sav_epc[19]), .B(regs_14[19]), .Z(n_17723
		));
	notech_reg_set sav_epc_reg_20(.CP(n_62217), .D(n_17730), .SD(1'b1), .Q(sav_epc
		[20]));
	notech_mux2 i_3151(.S(n_53833), .A(sav_epc[20]), .B(regs_14[20]), .Z(n_17730
		));
	notech_reg_set sav_epc_reg_21(.CP(n_62217), .D(n_17738), .SD(1'b1), .Q(sav_epc
		[21]));
	notech_mux2 i_3159(.S(n_53833), .A(sav_epc[21]), .B(regs_14[21]), .Z(n_17738
		));
	notech_reg_set sav_epc_reg_22(.CP(n_62217), .D(n_17745), .SD(1'b1), .Q(sav_epc
		[22]));
	notech_mux2 i_3167(.S(n_53833), .A(sav_epc[22]), .B(regs_14[22]), .Z(n_17745
		));
	notech_reg_set sav_epc_reg_23(.CP(n_62217), .D(n_17753), .SD(1'b1), .Q(sav_epc
		[23]));
	notech_mux2 i_3175(.S(n_53833), .A(sav_epc[23]), .B(regs_14[23]), .Z(n_17753
		));
	notech_reg_set sav_epc_reg_24(.CP(n_62217), .D(n_17760), .SD(1'b1), .Q(sav_epc
		[24]));
	notech_mux2 i_3183(.S(n_53833), .A(sav_epc[24]), .B(regs_14[24]), .Z(n_17760
		));
	notech_reg_set sav_epc_reg_25(.CP(n_62217), .D(n_17768), .SD(1'b1), .Q(sav_epc
		[25]));
	notech_mux2 i_3191(.S(n_53833), .A(sav_epc[25]), .B(regs_14[25]), .Z(n_17768
		));
	notech_reg_set sav_epc_reg_26(.CP(n_62217), .D(n_17775), .SD(1'b1), .Q(sav_epc
		[26]));
	notech_mux2 i_3199(.S(n_53833), .A(sav_epc[26]), .B(regs_14[26]), .Z(n_17775
		));
	notech_reg_set sav_epc_reg_27(.CP(n_62217), .D(n_17783), .SD(1'b1), .Q(sav_epc
		[27]));
	notech_mux2 i_3207(.S(n_53833), .A(sav_epc[27]), .B(regs_14[27]), .Z(n_17783
		));
	notech_reg_set sav_epc_reg_28(.CP(n_62217), .D(n_17790), .SD(1'b1), .Q(sav_epc
		[28]));
	notech_mux2 i_3215(.S(n_53833), .A(sav_epc[28]), .B(regs_14[28]), .Z(n_17790
		));
	notech_and4 i_327(.A(n_247656294), .B(n_247156289), .C(n_246856286), .D(instrc
		[124]), .Z(n_2341));
	notech_reg_set sav_epc_reg_29(.CP(n_62217), .D(n_17798), .SD(1'b1), .Q(sav_epc
		[29]));
	notech_mux2 i_3223(.S(n_53833), .A(sav_epc[29]), .B(regs_14[29]), .Z(n_17798
		));
	notech_nao3 i_827968(.A(n_2548), .B(n_2321), .C(n_2339), .Z(n_2340));
	notech_reg_set sav_epc_reg_30(.CP(n_62217), .D(n_17805), .SD(1'b1), .Q(sav_epc
		[30]));
	notech_mux2 i_3231(.S(n_53833), .A(sav_epc[30]), .B(regs_14[30]), .Z(n_17805
		));
	notech_ao3 i_298(.A(n_244856266), .B(instrc[63]), .C(n_2790), .Z(n_2339)
		);
	notech_reg_set sav_epc_reg_31(.CP(n_62217), .D(n_17813), .SD(1'b1), .Q(sav_epc
		[31]));
	notech_mux2 i_3239(.S(n_53833), .A(sav_epc[31]), .B(regs_14[31]), .Z(n_17813
		));
	notech_or2 i_312(.A(n_247056288), .B(n_29031), .Z(n_2338));
	notech_reg_set all_cnt_reg_0(.CP(n_62217), .D(n_17820), .SD(1'b1), .Q(all_cnt
		[0]));
	notech_mux2 i_3247(.S(n_26803), .A(all_cnt[0]), .B(n_26626), .Z(n_17820)
		);
	notech_nand3 i_304(.A(n_244756265), .B(n_246556283), .C(instrc[71]), .Z(n_2337
		));
	notech_reg_set all_cnt_reg_1(.CP(n_62157), .D(n_17828), .SD(1'b1), .Q(all_cnt
		[1]));
	notech_mux2 i_3255(.S(n_26803), .A(all_cnt[1]), .B(n_26801), .Z(n_17828)
		);
	notech_reg_set all_cnt_reg_2(.CP(n_62157), .D(n_17835), .SD(1'b1), .Q(all_cnt
		[2]));
	notech_mux2 i_3263(.S(n_26803), .A(all_cnt[2]), .B(n_189488133), .Z(n_17835
		));
	notech_reg_set all_cnt_reg_3(.CP(n_62157), .D(n_17843), .SD(1'b1), .Q(all_cnt
		[3]));
	notech_mux2 i_3271(.S(n_26803), .A(all_cnt[3]), .B(n_189588134), .Z(n_17843
		));
	notech_reg regs_reg_14_0(.CP(n_62157), .D(n_17850), .CD(n_61160), .Q(regs_14
		[0]));
	notech_mux2 i_3279(.S(n_26808), .A(regs_14[0]), .B(n_20111), .Z(n_17850)
		);
	notech_reg regs_reg_14_1(.CP(n_62157), .D(n_17858), .CD(n_61160), .Q(regs_14
		[1]));
	notech_mux2 i_3287(.S(n_26808), .A(regs_14[1]), .B(n_20117), .Z(n_17858)
		);
	notech_reg regs_reg_14_2(.CP(n_62157), .D(n_17865), .CD(n_61159), .Q(regs_14
		[2]));
	notech_mux2 i_3295(.S(n_26808), .A(regs_14[2]), .B(n_20123), .Z(n_17865)
		);
	notech_reg regs_reg_14_3(.CP(n_62157), .D(n_17873), .CD(n_61159), .Q(regs_14
		[3]));
	notech_mux2 i_3303(.S(n_26808), .A(regs_14[3]), .B(n_20129), .Z(n_17873)
		);
	notech_reg regs_reg_14_4(.CP(n_62157), .D(n_17880), .CD(n_61158), .Q(regs_14
		[4]));
	notech_mux2 i_3311(.S(n_26808), .A(regs_14[4]), .B(n_20135), .Z(n_17880)
		);
	notech_reg regs_reg_14_5(.CP(n_62157), .D(n_17888), .CD(n_61159), .Q(regs_14
		[5]));
	notech_mux2 i_3319(.S(n_26808), .A(regs_14[5]), .B(n_20141), .Z(n_17888)
		);
	notech_reg regs_reg_14_6(.CP(n_62157), .D(n_17895), .CD(n_61158), .Q(regs_14
		[6]));
	notech_mux2 i_3327(.S(n_26808), .A(regs_14[6]), .B(n_20147), .Z(n_17895)
		);
	notech_reg regs_reg_14_7(.CP(n_62297), .D(n_17903), .CD(n_61158), .Q(regs_14
		[7]));
	notech_mux2 i_3335(.S(n_26808), .A(regs_14[7]), .B(n_20153), .Z(n_17903)
		);
	notech_nand3 i_299(.A(n_247656294), .B(n_247256290), .C(instrc[127]), .Z
		(n_2321));
	notech_reg regs_reg_14_8(.CP(n_62155), .D(n_17910), .CD(n_61159), .Q(regs_14
		[8]));
	notech_mux2 i_3343(.S(n_26808), .A(regs_14[8]), .B(n_20159), .Z(n_17910)
		);
	notech_nao3 i_627966(.A(n_2536), .B(n_230388770), .C(n_2316), .Z(n_231756227
		));
	notech_reg regs_reg_14_9(.CP(n_62155), .D(n_17918), .CD(n_61159), .Q(regs_14
		[9]));
	notech_mux2 i_3351(.S(n_26808), .A(regs_14[9]), .B(n_20165), .Z(n_17918)
		);
	notech_ao3 i_270(.A(n_244856266), .B(instrc[61]), .C(n_2790), .Z(n_2316)
		);
	notech_reg_set regs_reg_14_10(.CP(n_62205), .D(n_17925), .SD(n_61159), .Q
		(regs_14[10]));
	notech_mux2 i_3359(.S(n_26808), .A(regs_14[10]), .B(n_20171), .Z(n_17925
		));
	notech_or2 i_284(.A(n_247056288), .B(n_29027), .Z(n_231588765));
	notech_reg_set regs_reg_14_11(.CP(n_62205), .D(n_17933), .SD(n_61159), .Q
		(regs_14[11]));
	notech_mux2 i_3367(.S(n_26808), .A(regs_14[11]), .B(n_20177), .Z(n_17933
		));
	notech_nand3 i_275(.A(n_244756265), .B(n_246556283), .C(instrc[69]), .Z(n_231456226
		));
	notech_reg_set regs_reg_14_12(.CP(n_62205), .D(n_17940), .SD(n_61159), .Q
		(regs_14[12]));
	notech_mux2 i_3375(.S(n_26808), .A(regs_14[12]), .B(n_20183), .Z(n_17940
		));
	notech_reg_set regs_reg_14_13(.CP(n_62205), .D(n_17948), .SD(n_61157), .Q
		(regs_14[13]));
	notech_mux2 i_3383(.S(n_26808), .A(regs_14[13]), .B(n_20189), .Z(n_17948
		));
	notech_reg_set regs_reg_14_14(.CP(n_62205), .D(n_17955), .SD(n_61154), .Q
		(regs_14[14]));
	notech_mux2 i_3391(.S(n_26808), .A(regs_14[14]), .B(n_20195), .Z(n_17955
		));
	notech_reg_set regs_reg_14_15(.CP(n_62205), .D(n_17963), .SD(n_61154), .Q
		(regs_14[15]));
	notech_mux2 i_3399(.S(n_26808), .A(regs_14[15]), .B(n_20201), .Z(n_17963
		));
	notech_reg_set regs_reg_14_16(.CP(n_62205), .D(n_17970), .SD(n_61154), .Q
		(regs_14[16]));
	notech_mux2 i_3407(.S(n_55508), .A(regs_14[16]), .B(n_20207), .Z(n_17970
		));
	notech_reg_set regs_reg_14_17(.CP(n_62205), .D(n_17978), .SD(n_61154), .Q
		(regs_14[17]));
	notech_mux2 i_3415(.S(n_55508), .A(regs_14[17]), .B(n_20213), .Z(n_17978
		));
	notech_reg_set regs_reg_14_18(.CP(n_62205), .D(n_17985), .SD(n_61154), .Q
		(regs_14[18]));
	notech_mux2 i_3423(.S(n_55508), .A(regs_14[18]), .B(n_20219), .Z(n_17985
		));
	notech_reg_set regs_reg_14_19(.CP(n_62205), .D(n_17993), .SD(n_61154), .Q
		(regs_14[19]));
	notech_mux2 i_3431(.S(n_55508), .A(regs_14[19]), .B(n_20225), .Z(n_17993
		));
	notech_reg regs_reg_14_20(.CP(n_62289), .D(n_18000), .CD(n_61154), .Q(regs_14
		[20]));
	notech_mux2 i_3439(.S(n_55508), .A(regs_14[20]), .B(n_20231), .Z(n_18000
		));
	notech_reg regs_reg_14_21(.CP(n_62289), .D(n_18008), .CD(n_61154), .Q(regs_14
		[21]));
	notech_mux2 i_3447(.S(n_55508), .A(regs_14[21]), .B(n_20237), .Z(n_18008
		));
	notech_reg regs_reg_14_22(.CP(n_62289), .D(n_18015), .CD(n_61154), .Q(regs_14
		[22]));
	notech_mux2 i_3455(.S(n_55508), .A(regs_14[22]), .B(n_20243), .Z(n_18015
		));
	notech_nand3 i_271(.A(n_247656294), .B(n_247256290), .C(instrc[125]), .Z
		(n_230388770));
	notech_reg regs_reg_14_23(.CP(n_62289), .D(n_18021), .CD(n_61153), .Q(regs_14
		[23]));
	notech_mux2 i_3463(.S(n_55508), .A(regs_14[23]), .B(n_20249), .Z(n_18021
		));
	notech_nao3 i_227962(.A(n_2524), .B(n_228988784), .C(n_230288771), .Z(\opcode[1] 
		));
	notech_reg regs_reg_14_24(.CP(n_62289), .D(n_18027), .CD(n_61153), .Q(regs_14
		[24]));
	notech_mux2 i_3471(.S(n_55508), .A(regs_14[24]), .B(n_20255), .Z(n_18027
		));
	notech_ao3 i_239(.A(n_244856266), .B(instrc[57]), .C(n_2790), .Z(n_230288771
		));
	notech_reg regs_reg_14_25(.CP(n_62289), .D(n_18033), .CD(n_61153), .Q(regs_14
		[25]));
	notech_mux2 i_3479(.S(n_55508), .A(regs_14[25]), .B(n_20261), .Z(n_18033
		));
	notech_or2 i_253(.A(n_247056288), .B(n_29024), .Z(n_230188772));
	notech_reg regs_reg_14_26(.CP(n_62289), .D(n_18039), .CD(n_61153), .Q(regs_14
		[26]));
	notech_mux2 i_3487(.S(n_55508), .A(regs_14[26]), .B(n_20267), .Z(n_18039
		));
	notech_nand3 i_244(.A(n_244756265), .B(n_246556283), .C(instrc[65]), .Z(n_230088773
		));
	notech_reg regs_reg_14_27(.CP(n_62289), .D(n_18045), .CD(n_61153), .Q(regs_14
		[27]));
	notech_mux2 i_3495(.S(n_55508), .A(regs_14[27]), .B(n_20273), .Z(n_18045
		));
	notech_reg regs_reg_14_28(.CP(n_62289), .D(n_18051), .CD(n_61153), .Q(regs_14
		[28]));
	notech_mux2 i_3503(.S(n_55508), .A(regs_14[28]), .B(n_20279), .Z(n_18051
		));
	notech_reg regs_reg_14_29(.CP(n_62289), .D(n_18057), .CD(n_61154), .Q(regs_14
		[29]));
	notech_mux2 i_3511(.S(n_55508), .A(regs_14[29]), .B(n_20285), .Z(n_18057
		));
	notech_reg regs_reg_14_30(.CP(n_62289), .D(n_18063), .CD(n_61153), .Q(regs_14
		[30]));
	notech_mux2 i_3519(.S(n_55508), .A(regs_14[30]), .B(n_20291), .Z(n_18063
		));
	notech_reg regs_reg_14_31(.CP(n_62289), .D(n_18069), .CD(n_61153), .Q(regs_14
		[31]));
	notech_mux2 i_3527(.S(n_55508), .A(regs_14[31]), .B(n_20297), .Z(n_18069
		));
	notech_reg regs_reg_13_0(.CP(n_62289), .D(n_18075), .CD(n_61154), .Q(gs[
		0]));
	notech_mux2 i_3535(.S(\nbus_11351[0] ), .A(gs[0]), .B(n_26809), .Z(n_18075
		));
	notech_reg regs_reg_13_1(.CP(n_62289), .D(n_18081), .CD(n_61155), .Q(gs[
		1]));
	notech_mux2 i_3543(.S(\nbus_11351[0] ), .A(gs[1]), .B(n_26810), .Z(n_18081
		));
	notech_reg regs_reg_13_2(.CP(n_62289), .D(n_18087), .CD(n_61155), .Q(gs[
		2]));
	notech_mux2 i_3551(.S(\nbus_11351[0] ), .A(n_55322), .B(n_26811), .Z(n_18087
		));
	notech_reg regs_reg_13_3(.CP(n_62289), .D(n_18093), .CD(n_61155), .Q(gs[
		3]));
	notech_mux2 i_3559(.S(\nbus_11351[0] ), .A(gs[3]), .B(n_19803), .Z(n_18093
		));
	notech_reg regs_reg_13_4(.CP(n_62289), .D(n_18099), .CD(n_61155), .Q(gs[
		4]));
	notech_mux2 i_3567(.S(\nbus_11351[0] ), .A(gs[4]), .B(n_26812), .Z(n_18099
		));
	notech_reg regs_reg_13_5(.CP(n_62289), .D(n_18105), .CD(n_61155), .Q(gs[
		5]));
	notech_mux2 i_3575(.S(\nbus_11351[0] ), .A(gs[5]), .B(n_19815), .Z(n_18105
		));
	notech_nand3 i_240(.A(n_247656294), .B(n_247256290), .C(n_60516), .Z(n_228988784
		));
	notech_reg regs_reg_13_6(.CP(n_62289), .D(n_18111), .CD(n_61157), .Q(gs[
		6]));
	notech_mux2 i_3583(.S(\nbus_11351[0] ), .A(gs[6]), .B(n_26813), .Z(n_18111
		));
	notech_ao3 i_203(.A(n_244856266), .B(instrc[56]), .C(n_2790), .Z(n_228888785
		));
	notech_reg regs_reg_13_7(.CP(n_62287), .D(n_18117), .CD(n_61157), .Q(gs[
		7]));
	notech_mux2 i_3591(.S(\nbus_11351[0] ), .A(gs[7]), .B(n_26814), .Z(n_18117
		));
	notech_or2 i_222(.A(n_247056288), .B(n_29021), .Z(n_228788786));
	notech_reg regs_reg_13_8(.CP(n_62287), .D(n_18123), .CD(n_61155), .Q(gs[
		8]));
	notech_mux2 i_3599(.S(\nbus_11351[0] ), .A(gs[8]), .B(n_19833), .Z(n_18123
		));
	notech_nand3 i_208(.A(n_244756265), .B(n_246556283), .C(instrc[64]), .Z(n_228688787
		));
	notech_reg regs_reg_13_9(.CP(n_62359), .D(n_18129), .CD(n_61157), .Q(gs[
		9]));
	notech_mux2 i_3607(.S(\nbus_11351[0] ), .A(gs[9]), .B(n_19839), .Z(n_18129
		));
	notech_reg regs_reg_13_10(.CP(n_62359), .D(n_18135), .CD(n_61155), .Q(gs
		[10]));
	notech_mux2 i_3615(.S(\nbus_11351[0] ), .A(gs[10]), .B(n_26815), .Z(n_18135
		));
	notech_reg regs_reg_13_11(.CP(n_62359), .D(n_18141), .CD(n_61155), .Q(gs
		[11]));
	notech_mux2 i_3623(.S(\nbus_11351[0] ), .A(gs[11]), .B(n_19851), .Z(n_18141
		));
	notech_reg regs_reg_13_12(.CP(n_62359), .D(n_18147), .CD(n_61154), .Q(gs
		[12]));
	notech_mux2 i_3631(.S(\nbus_11351[0] ), .A(gs[12]), .B(n_19857), .Z(n_18147
		));
	notech_reg regs_reg_13_13(.CP(n_62359), .D(n_18153), .CD(n_61154), .Q(gs
		[13]));
	notech_mux2 i_3639(.S(\nbus_11351[0] ), .A(gs[13]), .B(n_19863), .Z(n_18153
		));
	notech_reg regs_reg_13_14(.CP(n_62359), .D(n_18159), .CD(n_61155), .Q(gs
		[14]));
	notech_mux2 i_3647(.S(\nbus_11351[0] ), .A(gs[14]), .B(n_19869), .Z(n_18159
		));
	notech_reg regs_reg_13_15(.CP(n_62359), .D(n_18165), .CD(n_61155), .Q(gs
		[15]));
	notech_mux2 i_3655(.S(\nbus_11351[0] ), .A(gs[15]), .B(n_26816), .Z(n_18165
		));
	notech_reg regs_reg_13_16(.CP(n_62359), .D(n_18171), .CD(n_61155), .Q(gs
		[16]));
	notech_mux2 i_3663(.S(n_53884), .A(gs[16]), .B(n_19881), .Z(n_18171));
	notech_reg regs_reg_13_17(.CP(n_62359), .D(n_18177), .CD(n_61155), .Q(gs
		[17]));
	notech_mux2 i_3671(.S(n_53884), .A(gs[17]), .B(n_19887), .Z(n_18177));
	notech_reg regs_reg_13_18(.CP(n_62359), .D(n_18183), .CD(n_61155), .Q(gs
		[18]));
	notech_mux2 i_3679(.S(n_53884), .A(gs[18]), .B(n_19893), .Z(n_18183));
	notech_reg regs_reg_13_19(.CP(n_62359), .D(n_18189), .CD(n_61160), .Q(gs
		[19]));
	notech_mux2 i_3687(.S(n_53884), .A(gs[19]), .B(n_19899), .Z(n_18189));
	notech_nand3 i_204(.A(n_247656294), .B(n_247256290), .C(instrc[120]), .Z
		(n_227588798));
	notech_reg regs_reg_13_20(.CP(n_62359), .D(n_18195), .CD(n_61166), .Q(gs
		[20]));
	notech_mux2 i_3695(.S(n_53884), .A(gs[20]), .B(n_19905), .Z(n_18195));
	notech_ao3 i_169(.A(n_244856266), .B(instrc[59]), .C(n_2790), .Z(n_227488799
		));
	notech_reg regs_reg_13_21(.CP(n_62359), .D(n_18201), .CD(n_61166), .Q(gs
		[21]));
	notech_mux2 i_3703(.S(n_53884), .A(gs[21]), .B(n_19911), .Z(n_18201));
	notech_or2 i_182(.A(n_247056288), .B(n_29018), .Z(n_227388800));
	notech_reg regs_reg_13_22(.CP(n_62359), .D(n_18207), .CD(n_61165), .Q(gs
		[22]));
	notech_mux2 i_3711(.S(n_53884), .A(gs[22]), .B(n_26817), .Z(n_18207));
	notech_nand3 i_174(.A(n_244756265), .B(n_246556283), .C(instrc[67]), .Z(n_227288801
		));
	notech_reg regs_reg_13_23(.CP(n_62359), .D(n_18213), .CD(n_61165), .Q(gs
		[23]));
	notech_mux2 i_3719(.S(n_53884), .A(gs[23]), .B(n_19923), .Z(n_18213));
	notech_reg regs_reg_13_24(.CP(n_62359), .D(n_18219), .CD(n_61166), .Q(gs
		[24]));
	notech_mux2 i_3727(.S(n_53884), .A(gs[24]), .B(n_19929), .Z(n_18219));
	notech_reg regs_reg_13_25(.CP(n_62359), .D(n_18227), .CD(n_61166), .Q(gs
		[25]));
	notech_mux2 i_3735(.S(n_53884), .A(gs[25]), .B(n_19935), .Z(n_18227));
	notech_reg regs_reg_13_26(.CP(n_62359), .D(n_18233), .CD(n_61166), .Q(gs
		[26]));
	notech_mux2 i_3743(.S(n_53884), .A(gs[26]), .B(n_19941), .Z(n_18233));
	notech_reg regs_reg_13_27(.CP(n_62287), .D(n_18239), .CD(n_61166), .Q(gs
		[27]));
	notech_mux2 i_3751(.S(n_53884), .A(gs[27]), .B(n_19947), .Z(n_18239));
	notech_reg regs_reg_13_28(.CP(n_62287), .D(n_18245), .CD(n_61166), .Q(gs
		[28]));
	notech_mux2 i_3759(.S(n_53884), .A(gs[28]), .B(n_19953), .Z(n_18245));
	notech_reg regs_reg_13_29(.CP(n_62287), .D(n_18251), .CD(n_61165), .Q(gs
		[29]));
	notech_mux2 i_3767(.S(n_53884), .A(gs[29]), .B(n_26818), .Z(n_18251));
	notech_reg regs_reg_13_30(.CP(n_62287), .D(n_18258), .CD(n_61165), .Q(gs
		[30]));
	notech_mux2 i_3775(.S(n_53884), .A(gs[30]), .B(n_26819), .Z(n_18258));
	notech_reg regs_reg_13_31(.CP(n_62287), .D(n_18265), .CD(n_61165), .Q(gs
		[31]));
	notech_mux2 i_3783(.S(n_53884), .A(gs[31]), .B(n_19971), .Z(n_18265));
	notech_reg regs_reg_12_0(.CP(n_62287), .D(n_18273), .CD(n_61165), .Q(regs_12
		[0]));
	notech_mux2 i_3791(.S(\nbus_11350[0] ), .A(regs_12[0]), .B(n_19437), .Z(n_18273
		));
	notech_reg regs_reg_12_1(.CP(n_62287), .D(n_18280), .CD(n_61165), .Q(regs_12
		[1]));
	notech_mux2 i_3799(.S(\nbus_11350[0] ), .A(regs_12[1]), .B(n_26820), .Z(n_18280
		));
	notech_nand3 i_170(.A(n_247656294), .B(n_247256290), .C(n_60549), .Z(n_224756218
		));
	notech_reg regs_reg_12_2(.CP(n_62287), .D(n_18288), .CD(n_61165), .Q(regs_12
		[2]));
	notech_mux2 i_3807(.S(\nbus_11350[0] ), .A(regs_12[2]), .B(n_26822), .Z(n_18288
		));
	notech_ao3 i_139(.A(instrc[58]), .B(n_244856266), .C(n_2790), .Z(n_224656217
		));
	notech_reg regs_reg_12_3(.CP(n_62287), .D(n_18295), .CD(n_61165), .Q(regs_12
		[3]));
	notech_mux2 i_3815(.S(\nbus_11350[0] ), .A(regs_12[3]), .B(n_19455), .Z(n_18295
		));
	notech_or2 i_152(.A(n_247056288), .B(n_29015), .Z(n_2245));
	notech_reg regs_reg_12_4(.CP(n_62287), .D(n_18303), .CD(n_61165), .Q(regs_12
		[4]));
	notech_mux2 i_3823(.S(\nbus_11350[0] ), .A(regs_12[4]), .B(n_26823), .Z(n_18303
		));
	notech_nand3 i_144(.A(instrc[66]), .B(n_244756265), .C(n_246556283), .Z(n_224488804
		));
	notech_reg regs_reg_12_5(.CP(n_62359), .D(n_18310), .CD(n_61165), .Q(regs_12
		[5]));
	notech_mux2 i_3831(.S(\nbus_11350[0] ), .A(regs_12[5]), .B(n_19467), .Z(n_18310
		));
	notech_reg regs_reg_12_6(.CP(n_62355), .D(n_18318), .CD(n_61166), .Q(regs_12
		[6]));
	notech_mux2 i_3839(.S(\nbus_11350[0] ), .A(regs_12[6]), .B(n_26824), .Z(n_18318
		));
	notech_reg regs_reg_12_7(.CP(n_62285), .D(n_18325), .CD(n_61168), .Q(regs_12
		[7]));
	notech_mux2 i_3847(.S(\nbus_11350[0] ), .A(regs_12[7]), .B(n_26825), .Z(n_18325
		));
	notech_reg regs_reg_12_8(.CP(n_62355), .D(n_18333), .CD(n_61168), .Q(regs_12
		[8]));
	notech_mux2 i_3855(.S(\nbus_11350[0] ), .A(regs_12[8]), .B(n_26827), .Z(n_18333
		));
	notech_reg regs_reg_12_9(.CP(n_62355), .D(n_18340), .CD(n_61168), .Q(regs_12
		[9]));
	notech_mux2 i_3863(.S(\nbus_11350[0] ), .A(regs_12[9]), .B(n_19491), .Z(n_18340
		));
	notech_reg regs_reg_12_10(.CP(n_62355), .D(n_18348), .CD(n_61168), .Q(regs_12
		[10]));
	notech_mux2 i_3871(.S(\nbus_11350[0] ), .A(regs_12[10]), .B(n_19497), .Z
		(n_18348));
	notech_reg regs_reg_12_11(.CP(n_62355), .D(n_18355), .CD(n_61168), .Q(regs_12
		[11]));
	notech_mux2 i_3879(.S(\nbus_11350[0] ), .A(regs_12[11]), .B(n_19503), .Z
		(n_18355));
	notech_reg regs_reg_12_12(.CP(n_62355), .D(n_18363), .CD(n_61168), .Q(regs_12
		[12]));
	notech_mux2 i_3887(.S(\nbus_11350[0] ), .A(regs_12[12]), .B(n_19509), .Z
		(n_18363));
	notech_reg regs_reg_12_13(.CP(n_62355), .D(n_18370), .CD(n_61168), .Q(regs_12
		[13]));
	notech_mux2 i_3895(.S(\nbus_11350[0] ), .A(regs_12[13]), .B(n_19515), .Z
		(n_18370));
	notech_reg regs_reg_12_14(.CP(n_62355), .D(n_18378), .CD(n_61168), .Q(regs_12
		[14]));
	notech_mux2 i_3903(.S(\nbus_11350[0] ), .A(regs_12[14]), .B(n_19521), .Z
		(n_18378));
	notech_reg regs_reg_12_15(.CP(n_62355), .D(n_18385), .CD(n_61168), .Q(regs_12
		[15]));
	notech_mux2 i_3911(.S(\nbus_11350[0] ), .A(regs_12[15]), .B(n_26828), .Z
		(n_18385));
	notech_nand3 i_140(.A(n_247656294), .B(n_247256290), .C(n_60527), .Z(n_2228
		));
	notech_reg regs_reg_12_16(.CP(n_62355), .D(n_18393), .CD(n_61166), .Q(regs_12
		[16]));
	notech_mux2 i_3919(.S(n_53895), .A(regs_12[16]), .B(n_19533), .Z(n_18393
		));
	notech_nand2 i_2001(.A(vliw_pc[0]), .B(n_27267), .Z(n_54510));
	notech_reg regs_reg_12_17(.CP(n_62355), .D(n_18400), .CD(n_61166), .Q(regs_12
		[17]));
	notech_mux2 i_3927(.S(n_53895), .A(regs_12[17]), .B(n_19539), .Z(n_18400
		));
	notech_or2 i_2013(.A(vliw_pc[0]), .B(n_27267), .Z(n_54500));
	notech_reg regs_reg_12_18(.CP(n_62355), .D(n_18408), .CD(n_61166), .Q(regs_12
		[18]));
	notech_mux2 i_3935(.S(n_53895), .A(regs_12[18]), .B(n_19545), .Z(n_18408
		));
	notech_and4 i_100(.A(n_54777), .B(n_2788), .C(n_57380), .D(n_26291), .Z(n_2227
		));
	notech_reg regs_reg_12_19(.CP(n_62387), .D(n_18415), .CD(n_61166), .Q(regs_12
		[19]));
	notech_mux2 i_3943(.S(n_53895), .A(regs_12[19]), .B(n_19551), .Z(n_18415
		));
	notech_and4 i_46366(.A(fsm[1]), .B(n_244356261), .C(n_60752), .D(n_27262
		), .Z(n_57446));
	notech_reg regs_reg_12_20(.CP(n_62387), .D(n_18421), .CD(n_61166), .Q(regs_12
		[20]));
	notech_mux2 i_3951(.S(n_53895), .A(regs_12[20]), .B(n_19557), .Z(n_18421
		));
	notech_nand3 i_46357(.A(n_244556263), .B(n_2575), .C(n_27264), .Z(n_2225
		));
	notech_reg regs_reg_12_21(.CP(n_62387), .D(n_18427), .CD(n_61168), .Q(regs_12
		[21]));
	notech_mux2 i_3959(.S(n_53895), .A(regs_12[21]), .B(n_19563), .Z(n_18427
		));
	notech_nand3 i_46359(.A(n_206788846), .B(n_27265), .C(n_27262), .Z(n_222456215
		));
	notech_reg regs_reg_12_22(.CP(n_62387), .D(n_18433), .CD(n_61168), .Q(regs_12
		[22]));
	notech_mux2 i_3967(.S(n_53895), .A(regs_12[22]), .B(n_26829), .Z(n_18433
		));
	notech_or4 i_113932861(.A(n_62427), .B(\opcode[3] ), .C(n_60558), .D(n_59375
		), .Z(n_222356214));
	notech_reg regs_reg_12_23(.CP(n_62387), .D(n_18439), .CD(n_61168), .Q(regs_12
		[23]));
	notech_mux2 i_3975(.S(n_53895), .A(regs_12[23]), .B(n_19575), .Z(n_18439
		));
	notech_or4 i_159332840(.A(n_2385), .B(n_2361), .C(n_59369), .D(n_60490),
		 .Z(n_2221));
	notech_reg regs_reg_12_24(.CP(n_62387), .D(n_18445), .CD(n_61168), .Q(regs_12
		[24]));
	notech_mux2 i_3983(.S(n_53895), .A(regs_12[24]), .B(n_19581), .Z(n_18445
		));
	notech_reg regs_reg_12_25(.CP(n_62387), .D(n_18451), .CD(n_61165), .Q(regs_12
		[25]));
	notech_mux2 i_3991(.S(n_53895), .A(regs_12[25]), .B(n_19587), .Z(n_18451
		));
	notech_ao3 i_121631868(.A(n_2225), .B(n_222456215), .C(n_275988698), .Z(n_2219
		));
	notech_reg regs_reg_12_26(.CP(n_62387), .D(n_18457), .CD(n_61163), .Q(regs_12
		[26]));
	notech_mux2 i_3999(.S(n_53895), .A(regs_12[26]), .B(n_19593), .Z(n_18457
		));
	notech_and3 i_124131846(.A(n_58496), .B(n_54733), .C(n_54784), .Z(n_221888805
		));
	notech_reg regs_reg_12_27(.CP(n_62387), .D(n_18463), .CD(n_61163), .Q(regs_12
		[27]));
	notech_mux2 i_4007(.S(n_53895), .A(regs_12[27]), .B(n_19599), .Z(n_18463
		));
	notech_reg regs_reg_12_28(.CP(n_62387), .D(n_18469), .CD(n_61160), .Q(regs_12
		[28]));
	notech_mux2 i_4015(.S(n_53895), .A(regs_12[28]), .B(n_19605), .Z(n_18469
		));
	notech_reg regs_reg_12_29(.CP(n_62387), .D(n_18475), .CD(n_61163), .Q(regs_12
		[29]));
	notech_mux2 i_4023(.S(n_53895), .A(regs_12[29]), .B(n_26830), .Z(n_18475
		));
	notech_ao4 i_124231845(.A(n_2168), .B(n_60468), .C(n_59150), .D(n_26625)
		, .Z(n_2215));
	notech_reg regs_reg_12_30(.CP(n_62387), .D(n_18481), .CD(n_61163), .Q(regs_12
		[30]));
	notech_mux2 i_4031(.S(n_53895), .A(regs_12[30]), .B(n_26831), .Z(n_18481
		));
	notech_reg regs_reg_12_31(.CP(n_62387), .D(n_18487), .CD(n_61163), .Q(regs_12
		[31]));
	notech_mux2 i_4039(.S(n_53895), .A(regs_12[31]), .B(n_19623), .Z(n_18487
		));
	notech_nao3 i_127031825(.A(n_2225), .B(n_222456215), .C(n_276088697), .Z
		(n_2210));
	notech_reg regs_reg_11_0(.CP(n_62387), .D(n_18493), .CD(n_61163), .Q(regs_11
		[0]));
	notech_mux2 i_4047(.S(n_26844), .A(regs_11[0]), .B(n_26832), .Z(n_18493)
		);
	notech_nand2 i_127131824(.A(n_59899), .B(n_2225), .Z(n_220856212));
	notech_reg regs_reg_11_1(.CP(n_62387), .D(n_18499), .CD(n_61163), .Q(regs_11
		[1]));
	notech_mux2 i_4055(.S(n_26844), .A(regs_11[1]), .B(n_26833), .Z(n_18499)
		);
	notech_reg regs_reg_11_2(.CP(n_62387), .D(n_18505), .CD(n_61163), .Q(regs_11
		[2]));
	notech_mux2 i_4063(.S(n_26844), .A(regs_11[2]), .B(n_26834), .Z(n_18505)
		);
	notech_reg regs_reg_11_3(.CP(n_62387), .D(n_18511), .CD(n_61160), .Q(regs_11
		[3]));
	notech_mux2 i_4071(.S(n_26844), .A(regs_11[3]), .B(n_19107), .Z(n_18511)
		);
	notech_nand2 i_130931792(.A(n_59241), .B(n_59230), .Z(n_2202));
	notech_reg regs_reg_11_4(.CP(n_62387), .D(n_18517), .CD(n_61160), .Q(regs_11
		[4]));
	notech_mux2 i_4079(.S(n_26844), .A(regs_11[4]), .B(n_26835), .Z(n_18517)
		);
	notech_reg regs_reg_11_5(.CP(n_62355), .D(n_18523), .CD(n_61160), .Q(regs_11
		[5]));
	notech_mux2 i_4087(.S(n_26844), .A(regs_11[5]), .B(n_19119), .Z(n_18523)
		);
	notech_nand3 i_130631795(.A(n_222456215), .B(n_2225), .C(n_273488721), .Z
		(n_2200));
	notech_reg regs_reg_11_6(.CP(n_62387), .D(n_18529), .CD(n_61160), .Q(regs_11
		[6]));
	notech_mux2 i_4095(.S(n_26844), .A(regs_11[6]), .B(n_26836), .Z(n_18529)
		);
	notech_ao4 i_131131790(.A(n_2263), .B(n_26229), .C(n_1936), .D(n_26313),
		 .Z(n_2199));
	notech_reg regs_reg_11_7(.CP(n_62357), .D(n_18535), .CD(n_61160), .Q(regs_11
		[7]));
	notech_mux2 i_4103(.S(n_26844), .A(regs_11[7]), .B(n_26837), .Z(n_18535)
		);
	notech_nand2 i_185232818(.A(n_59299), .B(n_59290), .Z(n_2197));
	notech_reg regs_reg_11_8(.CP(n_62357), .D(n_18541), .CD(n_61160), .Q(regs_11
		[8]));
	notech_mux2 i_4111(.S(n_26844), .A(regs_11[8]), .B(n_26838), .Z(n_18541)
		);
	notech_reg regs_reg_11_9(.CP(n_62357), .D(n_18547), .CD(n_61160), .Q(regs_11
		[9]));
	notech_mux2 i_4119(.S(n_26844), .A(regs_11[9]), .B(n_19143), .Z(n_18547)
		);
	notech_or2 i_187432816(.A(n_59299), .B(n_59290), .Z(n_2189));
	notech_reg regs_reg_11_10(.CP(n_62357), .D(n_18553), .CD(n_61160), .Q(regs_11
		[10]));
	notech_mux2 i_4127(.S(n_26844), .A(regs_11[10]), .B(n_26839), .Z(n_18553
		));
	notech_and4 i_132531776(.A(n_276188696), .B(n_213488810), .C(n_59186), .D
		(n_2185), .Z(n_2188));
	notech_reg regs_reg_11_11(.CP(n_62357), .D(n_18559), .CD(n_61160), .Q(regs_11
		[11]));
	notech_mux2 i_4135(.S(n_26844), .A(regs_11[11]), .B(n_19155), .Z(n_18559
		));
	notech_reg regs_reg_11_12(.CP(n_62357), .D(n_18565), .CD(n_61163), .Q(regs_11
		[12]));
	notech_mux2 i_4143(.S(n_26844), .A(regs_11[12]), .B(n_19161), .Z(n_18565
		));
	notech_reg regs_reg_11_13(.CP(n_62357), .D(n_18571), .CD(n_61164), .Q(regs_11
		[13]));
	notech_mux2 i_4151(.S(n_26844), .A(regs_11[13]), .B(n_19167), .Z(n_18571
		));
	notech_ao3 i_131931782(.A(n_59137), .B(n_55657), .C(n_26622), .Z(n_2185)
		);
	notech_reg regs_reg_11_14(.CP(n_62357), .D(n_18577), .CD(n_61164), .Q(regs_11
		[14]));
	notech_mux2 i_4159(.S(n_26844), .A(regs_11[14]), .B(n_19173), .Z(n_18577
		));
	notech_reg regs_reg_11_15(.CP(n_62357), .D(n_18583), .CD(n_61164), .Q(regs_11
		[15]));
	notech_mux2 i_4167(.S(n_26844), .A(regs_11[15]), .B(n_26840), .Z(n_18583
		));
	notech_reg regs_reg_11_16(.CP(n_62357), .D(n_18589), .CD(n_61164), .Q(regs_11
		[16]));
	notech_mux2 i_4175(.S(n_53915), .A(regs_11[16]), .B(n_19185), .Z(n_18589
		));
	notech_reg regs_reg_11_17(.CP(n_62357), .D(n_18595), .CD(n_61164), .Q(regs_11
		[17]));
	notech_mux2 i_4183(.S(n_53915), .A(regs_11[17]), .B(n_19191), .Z(n_18595
		));
	notech_reg regs_reg_11_18(.CP(n_62357), .D(n_18601), .CD(n_61164), .Q(regs_11
		[18]));
	notech_mux2 i_4191(.S(n_53915), .A(regs_11[18]), .B(n_19197), .Z(n_18601
		));
	notech_ao4 i_133931763(.A(n_2169), .B(n_26889), .C(n_271388742), .D(n_1954
		), .Z(n_2174));
	notech_reg regs_reg_11_19(.CP(n_62357), .D(n_18607), .CD(n_61165), .Q(regs_11
		[19]));
	notech_mux2 i_4199(.S(n_53915), .A(regs_11[19]), .B(n_19203), .Z(n_18607
		));
	notech_reg regs_reg_11_20(.CP(n_62357), .D(n_18613), .CD(n_61164), .Q(regs_11
		[20]));
	notech_mux2 i_4207(.S(n_53915), .A(regs_11[20]), .B(n_19209), .Z(n_18613
		));
	notech_and4 i_134831757(.A(n_59104), .B(n_59095), .C(n_59086), .D(n_2171
		), .Z(n_2172));
	notech_reg regs_reg_11_21(.CP(n_62357), .D(n_18619), .CD(n_61164), .Q(regs_11
		[21]));
	notech_mux2 i_4215(.S(n_53915), .A(regs_11[21]), .B(n_19215), .Z(n_18619
		));
	notech_ao3 i_134431760(.A(n_2169), .B(n_59077), .C(opc[15]), .Z(n_2171)
		);
	notech_reg regs_reg_11_22(.CP(n_62357), .D(n_18625), .CD(n_61163), .Q(regs_11
		[22]));
	notech_mux2 i_4223(.S(n_53915), .A(regs_11[22]), .B(n_26841), .Z(n_18625
		));
	notech_reg regs_reg_11_23(.CP(n_62357), .D(n_18631), .CD(n_61163), .Q(regs_11
		[23]));
	notech_mux2 i_4231(.S(n_53915), .A(regs_11[23]), .B(n_19227), .Z(n_18631
		));
	notech_and4 i_7832789(.A(n_270388750), .B(nbus_11326[5]), .C(nbus_11326[
		7]), .D(nbus_11326[6]), .Z(n_2169));
	notech_reg regs_reg_11_24(.CP(n_62357), .D(n_18637), .CD(n_61163), .Q(regs_11
		[24]));
	notech_mux2 i_4239(.S(n_53915), .A(regs_11[24]), .B(n_19233), .Z(n_18637
		));
	notech_reg regs_reg_11_25(.CP(n_62357), .D(n_18643), .CD(n_61163), .Q(regs_11
		[25]));
	notech_mux2 i_4247(.S(n_53915), .A(regs_11[25]), .B(n_19239), .Z(n_18643
		));
	notech_reg regs_reg_11_26(.CP(n_62285), .D(n_18649), .CD(n_61164), .Q(regs_11
		[26]));
	notech_mux2 i_4255(.S(n_53915), .A(regs_11[26]), .B(n_19245), .Z(n_18649
		));
	notech_reg regs_reg_11_27(.CP(n_62285), .D(n_18655), .CD(n_61164), .Q(regs_11
		[27]));
	notech_mux2 i_4263(.S(n_53915), .A(regs_11[27]), .B(n_19251), .Z(n_18655
		));
	notech_reg regs_reg_11_28(.CP(n_62285), .D(n_18661), .CD(n_61164), .Q(regs_11
		[28]));
	notech_mux2 i_4271(.S(n_53915), .A(regs_11[28]), .B(n_19257), .Z(n_18661
		));
	notech_and4 i_135331752(.A(n_59068), .B(n_59059), .C(n_59050), .D(n_2158
		), .Z(n_2162));
	notech_reg regs_reg_11_29(.CP(n_62285), .D(n_18667), .CD(n_61164), .Q(regs_11
		[29]));
	notech_mux2 i_4279(.S(n_53915), .A(regs_11[29]), .B(n_26842), .Z(n_18667
		));
	notech_reg regs_reg_11_30(.CP(n_62285), .D(n_18673), .CD(n_61164), .Q(regs_11
		[30]));
	notech_mux2 i_4287(.S(n_53915), .A(regs_11[30]), .B(n_26843), .Z(n_18673
		));
	notech_reg regs_reg_11_31(.CP(n_62285), .D(n_18679), .CD(n_61208), .Q(regs_11
		[31]));
	notech_mux2 i_4295(.S(n_53915), .A(regs_11[31]), .B(n_19275), .Z(n_18679
		));
	notech_and3 i_135231753(.A(n_59041), .B(n_59032), .C(n_59023), .Z(n_2158
		));
	notech_reg regs_reg_10_0(.CP(n_62285), .D(n_18685), .CD(n_61208), .Q(regs_10
		[0]));
	notech_mux2 i_4303(.S(n_26852), .A(regs_10[0]), .B(n_26845), .Z(n_18685)
		);
	notech_reg regs_reg_10_1(.CP(n_62285), .D(n_18691), .CD(n_61208), .Q(regs_10
		[1]));
	notech_mux2 i_4311(.S(n_26852), .A(regs_10[1]), .B(n_26846), .Z(n_18691)
		);
	notech_reg regs_reg_10_2(.CP(n_62285), .D(n_18697), .CD(n_61208), .Q(regs_10
		[2]));
	notech_mux2 i_4319(.S(n_26852), .A(regs_10[2]), .B(n_26847), .Z(n_18697)
		);
	notech_and4 i_135931746(.A(n_59014), .B(n_59005), .C(n_58996), .D(n_2150
		), .Z(n_2153));
	notech_reg regs_reg_10_3(.CP(n_62285), .D(n_18703), .CD(n_61208), .Q(regs_10
		[3]));
	notech_mux2 i_4327(.S(n_26852), .A(regs_10[3]), .B(n_8997), .Z(n_18703)
		);
	notech_reg regs_reg_10_4(.CP(n_62205), .D(n_18709), .CD(n_61208), .Q(regs_10
		[4]));
	notech_mux2 i_4335(.S(n_26852), .A(regs_10[4]), .B(n_26848), .Z(n_18709)
		);
	notech_reg regs_reg_10_5(.CP(n_62285), .D(n_18715), .CD(n_61208), .Q(regs_10
		[5]));
	notech_mux2 i_4343(.S(n_26852), .A(regs_10[5]), .B(n_9009), .Z(n_18715)
		);
	notech_and3 i_135831747(.A(n_58987), .B(n_58978), .C(n_58969), .Z(n_2150
		));
	notech_reg regs_reg_10_6(.CP(n_62291), .D(n_18721), .CD(n_61208), .Q(regs_10
		[6]));
	notech_mux2 i_4351(.S(n_26852), .A(regs_10[6]), .B(n_26849), .Z(n_18721)
		);
	notech_reg regs_reg_10_7(.CP(n_62207), .D(n_18727), .CD(n_61208), .Q(regs_10
		[7]));
	notech_mux2 i_4359(.S(n_26852), .A(regs_10[7]), .B(n_26850), .Z(n_18727)
		);
	notech_and4 i_136531740(.A(nbus_11326[12]), .B(nbus_11326[13]), .C(n_2144
		), .D(nbus_11326[14]), .Z(n_214888806));
	notech_reg regs_reg_10_8(.CP(n_62207), .D(n_18733), .CD(n_61205), .Q(regs_10
		[8]));
	notech_mux2 i_4367(.S(n_26852), .A(regs_10[8]), .B(n_9027), .Z(n_18733)
		);
	notech_reg regs_reg_10_9(.CP(n_62207), .D(n_18739), .CD(n_61205), .Q(regs_10
		[9]));
	notech_mux2 i_4375(.S(n_26852), .A(regs_10[9]), .B(n_9033), .Z(n_18739)
		);
	notech_reg regs_reg_10_10(.CP(n_62207), .D(n_18745), .CD(n_61205), .Q(regs_10
		[10]));
	notech_mux2 i_4383(.S(n_26852), .A(regs_10[10]), .B(n_9039), .Z(n_18745)
		);
	notech_and4 i_136431741(.A(nbus_11326[10]), .B(nbus_11326[11]), .C(nbus_11326
		[9]), .D(nbus_11326[8]), .Z(n_2144));
	notech_reg regs_reg_10_11(.CP(n_62207), .D(n_18751), .CD(n_61205), .Q(regs_10
		[11]));
	notech_mux2 i_4391(.S(n_26852), .A(regs_10[11]), .B(n_9045), .Z(n_18751)
		);
	notech_reg regs_reg_10_12(.CP(n_62207), .D(n_18757), .CD(n_61205), .Q(regs_10
		[12]));
	notech_mux2 i_4399(.S(n_26852), .A(regs_10[12]), .B(n_9051), .Z(n_18757)
		);
	notech_reg regs_reg_10_13(.CP(n_62207), .D(n_18763), .CD(n_61208), .Q(regs_10
		[13]));
	notech_mux2 i_4407(.S(n_26852), .A(regs_10[13]), .B(n_9057), .Z(n_18763)
		);
	notech_reg regs_reg_10_14(.CP(n_62207), .D(n_18769), .CD(n_61208), .Q(regs_10
		[14]));
	notech_mux2 i_4415(.S(n_26852), .A(regs_10[14]), .B(n_9063), .Z(n_18769)
		);
	notech_reg regs_reg_10_15(.CP(n_62207), .D(n_18775), .CD(n_61205), .Q(regs_10
		[15]));
	notech_mux2 i_4423(.S(n_26852), .A(regs_10[15]), .B(n_26851), .Z(n_18775
		));
	notech_reg regs_reg_10_16(.CP(n_62207), .D(n_18781), .CD(n_61208), .Q(regs_10
		[16]));
	notech_mux2 i_4431(.S(n_53926), .A(regs_10[16]), .B(n_9075), .Z(n_18781)
		);
	notech_reg regs_reg_10_17(.CP(n_62293), .D(n_18787), .CD(n_61208), .Q(regs_10
		[17]));
	notech_mux2 i_4439(.S(n_53926), .A(regs_10[17]), .B(n_9081), .Z(n_18787)
		);
	notech_reg regs_reg_10_18(.CP(n_62293), .D(n_18793), .CD(n_61209), .Q(regs_10
		[18]));
	notech_mux2 i_4447(.S(n_53926), .A(regs_10[18]), .B(n_9087), .Z(n_18793)
		);
	notech_xor2 i_137331733(.A(nbus_11326[4]), .B(n_48760), .Z(n_213688808)
		);
	notech_reg regs_reg_10_19(.CP(n_62293), .D(n_18799), .CD(n_61209), .Q(regs_10
		[19]));
	notech_mux2 i_4455(.S(n_53926), .A(regs_10[19]), .B(n_9093), .Z(n_18799)
		);
	notech_reg regs_reg_10_20(.CP(n_62293), .D(n_18805), .CD(n_61209), .Q(regs_10
		[20]));
	notech_mux2 i_4463(.S(n_53926), .A(regs_10[20]), .B(n_9099), .Z(n_18805)
		);
	notech_and4 i_132431777(.A(n_54862), .B(n_54818), .C(n_48496), .D(n_213388811
		), .Z(n_213488810));
	notech_reg regs_reg_10_21(.CP(n_62293), .D(n_18811), .CD(n_61209), .Q(regs_10
		[21]));
	notech_mux2 i_4471(.S(n_53926), .A(regs_10[21]), .B(n_9105), .Z(n_18811)
		);
	notech_ao4 i_132131780(.A(n_2190), .B(n_190388902), .C(n_994), .D(n_273388722
		), .Z(n_213388811));
	notech_reg regs_reg_10_22(.CP(n_62293), .D(n_18817), .CD(n_61210), .Q(regs_10
		[22]));
	notech_mux2 i_4479(.S(n_53926), .A(regs_10[22]), .B(n_9111), .Z(n_18817)
		);
	notech_reg regs_reg_10_23(.CP(n_62293), .D(n_18823), .CD(n_61210), .Q(regs_10
		[23]));
	notech_mux2 i_4487(.S(n_53926), .A(regs_10[23]), .B(n_9117), .Z(n_18823)
		);
	notech_reg regs_reg_10_24(.CP(n_62293), .D(n_18829), .CD(n_61210), .Q(regs_10
		[24]));
	notech_mux2 i_4495(.S(n_53926), .A(regs_10[24]), .B(n_9123), .Z(n_18829)
		);
	notech_reg regs_reg_10_25(.CP(n_62293), .D(n_18835), .CD(n_61210), .Q(regs_10
		[25]));
	notech_mux2 i_4503(.S(n_53926), .A(regs_10[25]), .B(n_9129), .Z(n_18835)
		);
	notech_nao3 i_137831729(.A(n_206788846), .B(n_26497), .C(n_60724), .Z(n_212988815
		));
	notech_reg regs_reg_10_26(.CP(n_62293), .D(n_18842), .CD(n_61210), .Q(regs_10
		[26]));
	notech_mux2 i_4511(.S(n_53926), .A(regs_10[26]), .B(n_9135), .Z(n_18842)
		);
	notech_reg regs_reg_10_27(.CP(n_62293), .D(n_18849), .CD(n_61209), .Q(regs_10
		[27]));
	notech_mux2 i_4519(.S(n_53926), .A(regs_10[27]), .B(n_9141), .Z(n_18849)
		);
	notech_and4 i_132931772(.A(n_2175), .B(n_2191), .C(n_1914), .D(n_212488820
		), .Z(n_212788817));
	notech_reg regs_reg_10_28(.CP(n_62293), .D(n_18855), .CD(n_61209), .Q(regs_10
		[28]));
	notech_mux2 i_4527(.S(n_53926), .A(regs_10[28]), .B(n_9147), .Z(n_18855)
		);
	notech_reg regs_reg_10_29(.CP(n_62293), .D(n_18862), .CD(n_61209), .Q(regs_10
		[29]));
	notech_mux2 i_4535(.S(n_53926), .A(regs_10[29]), .B(n_9153), .Z(n_18862)
		);
	notech_reg regs_reg_10_30(.CP(n_62293), .D(n_18868), .CD(n_61209), .Q(regs_10
		[30]));
	notech_mux2 i_4543(.S(n_53926), .A(regs_10[30]), .B(n_9159), .Z(n_18868)
		);
	notech_and2 i_132731774(.A(n_1918), .B(n_26745), .Z(n_212488820));
	notech_reg regs_reg_10_31(.CP(n_62293), .D(n_18874), .CD(n_61209), .Q(regs_10
		[31]));
	notech_mux2 i_4551(.S(n_53926), .A(regs_10[31]), .B(n_9165), .Z(n_18874)
		);
	notech_reg regs_reg_9_0(.CP(n_62293), .D(n_18880), .CD(n_61209), .Q(cs[0
		]));
	notech_mux2 i_4560(.S(\nbus_11332[0] ), .A(cs[0]), .B(n_26853), .Z(n_18880
		));
	notech_reg regs_reg_9_1(.CP(n_62293), .D(n_18886), .CD(n_61209), .Q(cs[1
		]));
	notech_mux2 i_4568(.S(\nbus_11332[0] ), .A(cs[1]), .B(n_26854), .Z(n_18886
		));
	notech_ao4 i_138831722(.A(n_275788700), .B(n_494), .C(n_1945), .D(n_60468
		), .Z(n_212188823));
	notech_reg regs_reg_9_2(.CP(n_62293), .D(n_18892), .CD(n_61209), .Q(\nbus_14524[2] 
		));
	notech_mux2 i_4576(.S(\nbus_11332[0] ), .A(\nbus_14524[2] ), .B(n_26855)
		, .Z(n_18892));
	notech_reg regs_reg_9_3(.CP(n_62293), .D(n_18898), .CD(n_61209), .Q(\nbus_14524[3] 
		));
	notech_mux2 i_4584(.S(\nbus_11332[0] ), .A(\nbus_14524[3] ), .B(n_26857)
		, .Z(n_18898));
	notech_reg regs_reg_9_4(.CP(n_62361), .D(n_18904), .CD(n_61205), .Q(\nbus_14524[4] 
		));
	notech_mux2 i_4592(.S(\nbus_11332[0] ), .A(\nbus_14524[4] ), .B(n_26858)
		, .Z(n_18904));
	notech_and3 i_162432834(.A(n_57419), .B(n_276588692), .C(n_2105), .Z(n_211888826
		));
	notech_reg regs_reg_9_5(.CP(n_62291), .D(n_18910), .CD(n_61203), .Q(\nbus_14524[5] 
		));
	notech_mux2 i_4600(.S(\nbus_11332[0] ), .A(\nbus_14524[5] ), .B(n_16729)
		, .Z(n_18910));
	notech_reg regs_reg_9_6(.CP(n_62361), .D(n_18916), .CD(n_61203), .Q(\nbus_14524[6] 
		));
	notech_mux2 i_4608(.S(\nbus_11332[0] ), .A(\nbus_14524[6] ), .B(n_26859)
		, .Z(n_18916));
	notech_reg regs_reg_9_7(.CP(n_62361), .D(n_18923), .CD(n_61203), .Q(\nbus_14524[7] 
		));
	notech_mux2 i_4616(.S(\nbus_11332[0] ), .A(\nbus_14524[7] ), .B(n_26860)
		, .Z(n_18923));
	notech_ao4 i_138531724(.A(n_2209), .B(n_2192), .C(n_2161), .D(n_2205), .Z
		(n_211588829));
	notech_reg regs_reg_9_8(.CP(n_62361), .D(n_18930), .CD(n_61203), .Q(\nbus_14524[8] 
		));
	notech_mux2 i_4624(.S(\nbus_11332[0] ), .A(\nbus_14524[8] ), .B(n_26861)
		, .Z(n_18930));
	notech_reg regs_reg_9_9(.CP(n_62361), .D(n_18936), .CD(n_61203), .Q(\nbus_14524[9] 
		));
	notech_mux2 i_4632(.S(\nbus_11332[0] ), .A(\nbus_14524[9] ), .B(n_26863)
		, .Z(n_18936));
	notech_and4 i_133531767(.A(n_2155), .B(n_211088832), .C(n_2073), .D(n_1981
		), .Z(n_211288830));
	notech_reg regs_reg_9_10(.CP(n_62361), .D(n_18942), .CD(n_61203), .Q(\nbus_14524[10] 
		));
	notech_mux2 i_4640(.S(\nbus_11332[0] ), .A(\nbus_14524[10] ), .B(n_26864
		), .Z(n_18942));
	notech_reg regs_reg_9_11(.CP(n_62361), .D(n_18948), .CD(n_61203), .Q(\nbus_14524[11] 
		));
	notech_mux2 i_4648(.S(\nbus_11332[0] ), .A(\nbus_14524[11] ), .B(n_16765
		), .Z(n_18948));
	notech_ao4 i_133131771(.A(n_274788710), .B(n_2205), .C(n_192088898), .D(n_60468
		), .Z(n_211088832));
	notech_reg regs_reg_9_12(.CP(n_62361), .D(n_18954), .CD(n_61203), .Q(\nbus_14524[12] 
		));
	notech_mux2 i_4656(.S(\nbus_11332[0] ), .A(\nbus_14524[12] ), .B(n_16771
		), .Z(n_18954));
	notech_reg regs_reg_9_13(.CP(n_62361), .D(n_18960), .CD(n_61203), .Q(\nbus_14524[13] 
		));
	notech_mux2 i_4664(.S(\nbus_11332[0] ), .A(\nbus_14524[13] ), .B(n_16777
		), .Z(n_18960));
	notech_reg regs_reg_9_14(.CP(n_62361), .D(n_18966), .CD(n_61202), .Q(\nbus_14524[14] 
		));
	notech_mux2 i_4672(.S(\nbus_11332[0] ), .A(\nbus_14524[14] ), .B(n_16783
		), .Z(n_18966));
	notech_ao4 i_139631716(.A(n_2271), .B(n_27112), .C(n_1943), .D(n_57423),
		 .Z(n_2106));
	notech_reg regs_reg_9_15(.CP(n_62361), .D(n_18972), .CD(n_61202), .Q(\nbus_14524[15] 
		));
	notech_mux2 i_4680(.S(\nbus_11332[0] ), .A(\nbus_14524[15] ), .B(n_26866
		), .Z(n_18972));
	notech_reg regs_reg_9_16(.CP(n_62361), .D(n_18978), .CD(n_61202), .Q(\nbus_14524[16] 
		));
	notech_mux2 i_4688(.S(n_56316), .A(\nbus_14524[16] ), .B(n_16795), .Z(n_18978
		));
	notech_or4 i_140331710(.A(n_210288837), .B(opb[24]), .C(opb[13]), .D(opb
		[9]), .Z(n_210388836));
	notech_reg regs_reg_9_17(.CP(n_62361), .D(n_18984), .CD(n_61202), .Q(\nbus_14524[17] 
		));
	notech_mux2 i_4696(.S(n_56316), .A(\nbus_14524[17] ), .B(n_16801), .Z(n_18984
		));
	notech_or4 i_139931713(.A(opb[15]), .B(opb[28]), .C(n_2096), .D(n_209988840
		), .Z(n_210288837));
	notech_reg regs_reg_9_18(.CP(n_62361), .D(n_18990), .CD(n_61202), .Q(\nbus_14524[18] 
		));
	notech_mux2 i_4704(.S(n_56316), .A(\nbus_14524[18] ), .B(n_16807), .Z(n_18990
		));
	notech_reg regs_reg_9_19(.CP(n_62361), .D(n_18996), .CD(n_61203), .Q(\nbus_14524[19] 
		));
	notech_mux2 i_4712(.S(n_56316), .A(\nbus_14524[19] ), .B(n_16813), .Z(n_18996
		));
	notech_reg regs_reg_9_20(.CP(n_62361), .D(n_19002), .CD(n_61203), .Q(\nbus_14524[20] 
		));
	notech_mux2 i_4720(.S(n_56316), .A(\nbus_14524[20] ), .B(n_16819), .Z(n_19002
		));
	notech_or4 i_142631689(.A(opb[7]), .B(opb[5]), .C(opb[4]), .D(opb[6]), .Z
		(n_209988840));
	notech_reg regs_reg_9_21(.CP(n_62361), .D(n_19008), .CD(n_61203), .Q(\nbus_14524[21] 
		));
	notech_mux2 i_4728(.S(n_56316), .A(\nbus_14524[21] ), .B(n_16825), .Z(n_19008
		));
	notech_reg regs_reg_9_22(.CP(n_62361), .D(n_19014), .CD(n_61203), .Q(\nbus_14524[22] 
		));
	notech_mux2 i_4736(.S(n_56316), .A(\nbus_14524[22] ), .B(n_26868), .Z(n_19014
		));
	notech_reg regs_reg_9_23(.CP(n_62361), .D(n_19020), .CD(n_61204), .Q(\nbus_14524[23] 
		));
	notech_mux2 i_4744(.S(n_56316), .A(\nbus_14524[23] ), .B(n_16837), .Z(n_19020
		));
	notech_or4 i_142931686(.A(opb[0]), .B(opb[1]), .C(opb[2]), .D(opb[3]), .Z
		(n_2096));
	notech_reg regs_reg_9_24(.CP(n_62291), .D(n_19026), .CD(n_61204), .Q(\nbus_14524[24] 
		));
	notech_mux2 i_4752(.S(n_56316), .A(\nbus_14524[24] ), .B(n_16843), .Z(n_19026
		));
	notech_reg regs_reg_9_25(.CP(n_62291), .D(n_19032), .CD(n_61205), .Q(\nbus_14524[25] 
		));
	notech_mux2 i_4760(.S(n_56316), .A(\nbus_14524[25] ), .B(n_16849), .Z(n_19032
		));
	notech_reg regs_reg_9_26(.CP(n_62291), .D(n_19038), .CD(n_61204), .Q(\nbus_14524[26] 
		));
	notech_mux2 i_4768(.S(n_56316), .A(\nbus_14524[26] ), .B(n_16855), .Z(n_19038
		));
	notech_reg regs_reg_9_27(.CP(n_62291), .D(n_19044), .CD(n_61204), .Q(\nbus_14524[27] 
		));
	notech_mux2 i_4776(.S(n_56316), .A(\nbus_14524[27] ), .B(n_16861), .Z(n_19044
		));
	notech_reg regs_reg_9_28(.CP(n_62291), .D(n_19050), .CD(n_61205), .Q(\nbus_14524[28] 
		));
	notech_mux2 i_4784(.S(n_56316), .A(\nbus_14524[28] ), .B(n_16867), .Z(n_19050
		));
	notech_or4 i_140831705(.A(opb[30]), .B(opb[29]), .C(opb[31]), .D(n_2088)
		, .Z(n_2091));
	notech_reg regs_reg_9_29(.CP(n_62291), .D(n_19056), .CD(n_61205), .Q(\nbus_14524[29] 
		));
	notech_mux2 i_4792(.S(n_56316), .A(\nbus_14524[29] ), .B(n_16873), .Z(n_19056
		));
	notech_reg regs_reg_9_30(.CP(n_62291), .D(n_19062), .CD(n_61205), .Q(\nbus_14524[30] 
		));
	notech_mux2 i_4800(.S(n_56316), .A(\nbus_14524[30] ), .B(n_26870), .Z(n_19062
		));
	notech_reg regs_reg_9_31(.CP(n_62291), .D(n_19068), .CD(n_61205), .Q(\nbus_14524[31] 
		));
	notech_mux2 i_4808(.S(n_56316), .A(\nbus_14524[31] ), .B(n_16885), .Z(n_19068
		));
	notech_nand3 i_140731706(.A(n_59346), .B(n_59337), .C(n_59328), .Z(n_2088
		));
	notech_reg regs_reg_8_0(.CP(n_62291), .D(n_19074), .CD(n_61205), .Q(regs_8
		[0]));
	notech_mux2 i_4816(.S(n_26881), .A(regs_8[0]), .B(n_26871), .Z(n_19074)
		);
	notech_reg regs_reg_8_1(.CP(n_62291), .D(n_19080), .CD(n_61204), .Q(regs_8
		[1]));
	notech_mux2 i_4824(.S(n_26881), .A(regs_8[1]), .B(n_26872), .Z(n_19080)
		);
	notech_reg regs_reg_8_2(.CP(n_62207), .D(n_19086), .CD(n_61204), .Q(regs_8
		[2]));
	notech_mux2 i_4832(.S(n_26881), .A(regs_8[2]), .B(n_26873), .Z(n_19086)
		);
	notech_or4 i_141431699(.A(opb[18]), .B(opb[19]), .C(opb[20]), .D(n_2084)
		, .Z(n_2085));
	notech_reg regs_reg_8_3(.CP(n_62207), .D(n_19093), .CD(n_61204), .Q(regs_8
		[3]));
	notech_mux2 i_4840(.S(n_26881), .A(regs_8[3]), .B(n_13833), .Z(n_19093)
		);
	notech_nao3 i_141131702(.A(n_59319), .B(n_59310), .C(opb[22]), .Z(n_2084
		));
	notech_reg regs_reg_8_4(.CP(n_62295), .D(n_19100), .CD(n_61204), .Q(regs_8
		[4]));
	notech_mux2 i_4848(.S(n_26881), .A(regs_8[4]), .B(n_26874), .Z(n_19100)
		);
	notech_reg regs_reg_8_5(.CP(n_62209), .D(n_19108), .CD(n_61204), .Q(regs_8
		[5]));
	notech_mux2 i_4856(.S(n_26881), .A(regs_8[5]), .B(n_13845), .Z(n_19108)
		);
	notech_reg regs_reg_8_6(.CP(n_62209), .D(n_19115), .CD(n_61204), .Q(regs_8
		[6]));
	notech_mux2 i_4864(.S(n_26881), .A(regs_8[6]), .B(n_26875), .Z(n_19115)
		);
	notech_reg regs_reg_8_7(.CP(n_62209), .D(n_19122), .CD(n_61204), .Q(regs_8
		[7]));
	notech_mux2 i_4872(.S(n_26881), .A(regs_8[7]), .B(n_26876), .Z(n_19122)
		);
	notech_or4 i_142031693(.A(opb[14]), .B(opb[16]), .C(opb[17]), .D(n_2077)
		, .Z(n_2080));
	notech_reg regs_reg_8_8(.CP(n_62209), .D(n_19129), .CD(n_61204), .Q(regs_8
		[8]));
	notech_mux2 i_4880(.S(n_26881), .A(regs_8[8]), .B(n_13863), .Z(n_19129)
		);
	notech_reg regs_reg_8_9(.CP(n_62209), .D(n_19136), .CD(n_61204), .Q(regs_8
		[9]));
	notech_mux2 i_4888(.S(n_26881), .A(regs_8[9]), .B(n_13869), .Z(n_19136)
		);
	notech_reg regs_reg_8_10(.CP(n_62209), .D(n_19144), .CD(n_61210), .Q(regs_8
		[10]));
	notech_mux2 i_4896(.S(n_26881), .A(regs_8[10]), .B(n_13875), .Z(n_19144)
		);
	notech_or4 i_141931694(.A(opb[11]), .B(opb[12]), .C(opb[8]), .D(opb[10])
		, .Z(n_2077));
	notech_reg regs_reg_8_11(.CP(n_62209), .D(n_19151), .CD(n_61215), .Q(regs_8
		[11]));
	notech_mux2 i_4904(.S(n_26881), .A(regs_8[11]), .B(n_13881), .Z(n_19151)
		);
	notech_reg regs_reg_8_12(.CP(n_62209), .D(n_19158), .CD(n_61215), .Q(regs_8
		[12]));
	notech_mux2 i_4912(.S(n_26881), .A(regs_8[12]), .B(n_13887), .Z(n_19158)
		);
	notech_reg regs_reg_8_13(.CP(n_62209), .D(n_19165), .CD(n_61215), .Q(regs_8
		[13]));
	notech_mux2 i_4920(.S(n_26881), .A(regs_8[13]), .B(n_13893), .Z(n_19165)
		);
	notech_reg regs_reg_8_14(.CP(n_62209), .D(n_19172), .CD(n_61215), .Q(regs_8
		[14]));
	notech_mux2 i_4928(.S(n_26881), .A(regs_8[14]), .B(n_13899), .Z(n_19172)
		);
	notech_ao4 i_133331769(.A(n_1941), .B(n_2209), .C(n_1940), .D(n_206988844
		), .Z(n_2073));
	notech_reg regs_reg_8_15(.CP(n_62295), .D(n_19180), .CD(n_61215), .Q(regs_8
		[15]));
	notech_mux2 i_4936(.S(n_26881), .A(regs_8[15]), .B(n_26878), .Z(n_19180)
		);
	notech_ao4 i_143031685(.A(n_2352), .B(nZF), .C(n_54689), .D(n_26403), .Z
		(n_2072));
	notech_reg regs_reg_8_16(.CP(n_62295), .D(n_19187), .CD(n_61215), .Q(regs_8
		[16]));
	notech_mux2 i_4944(.S(n_53982), .A(regs_8[16]), .B(n_13911), .Z(n_19187)
		);
	notech_ao4 i_143131684(.A(n_27146), .B(n_2196), .C(n_2107), .D(n_22579221
		), .Z(n_207188842));
	notech_reg regs_reg_8_17(.CP(n_62295), .D(n_19194), .CD(n_61215), .Q(regs_8
		[17]));
	notech_mux2 i_4952(.S(n_53982), .A(regs_8[17]), .B(n_13917), .Z(n_19194)
		);
	notech_reg regs_reg_8_18(.CP(n_62295), .D(n_19201), .CD(n_61215), .Q(regs_8
		[18]));
	notech_mux2 i_4960(.S(n_53982), .A(regs_8[18]), .B(n_13923), .Z(n_19201)
		);
	notech_nand2 i_143331682(.A(n_26616), .B(n_26773), .Z(n_206988844));
	notech_reg regs_reg_8_19(.CP(n_62295), .D(n_19208), .CD(n_61215), .Q(regs_8
		[19]));
	notech_mux2 i_4968(.S(n_53982), .A(regs_8[19]), .B(n_13929), .Z(n_19208)
		);
	notech_reg regs_reg_8_20(.CP(n_62295), .D(n_19216), .CD(n_61214), .Q(regs_8
		[20]));
	notech_mux2 i_4976(.S(n_53982), .A(regs_8[20]), .B(n_13935), .Z(n_19216)
		);
	notech_ao3 i_143531680(.A(fsm[2]), .B(n_27266), .C(fsm[1]), .Z(n_206788846
		));
	notech_reg regs_reg_8_21(.CP(n_62295), .D(n_19223), .CD(n_61214), .Q(regs_8
		[21]));
	notech_mux2 i_4984(.S(n_53982), .A(regs_8[21]), .B(n_13941), .Z(n_19223)
		);
	notech_or4 i_54332900(.A(n_2601), .B(n_494), .C(n_26380), .D(n_2604), .Z
		(n_206688847));
	notech_reg regs_reg_8_22(.CP(n_62295), .D(n_19230), .CD(n_61214), .Q(regs_8
		[22]));
	notech_mux2 i_4992(.S(n_53982), .A(regs_8[22]), .B(n_26879), .Z(n_19230)
		);
	notech_reg regs_reg_8_23(.CP(n_62295), .D(n_19237), .CD(n_61214), .Q(regs_8
		[23]));
	notech_mux2 i_5000(.S(n_53982), .A(regs_8[23]), .B(n_13953), .Z(n_19237)
		);
	notech_ao4 i_144831667(.A(n_59210), .B(n_59369), .C(n_59201), .D(n_26865
		), .Z(n_206488849));
	notech_reg regs_reg_8_24(.CP(n_62295), .D(n_19244), .CD(n_61214), .Q(regs_8
		[24]));
	notech_mux2 i_5008(.S(n_53982), .A(regs_8[24]), .B(n_13959), .Z(n_19244)
		);
	notech_reg regs_reg_8_25(.CP(n_62295), .D(n_19252), .CD(n_61214), .Q(regs_8
		[25]));
	notech_mux2 i_5016(.S(n_53982), .A(regs_8[25]), .B(n_13965), .Z(n_19252)
		);
	notech_or2 i_185832817(.A(n_59299), .B(n_28564), .Z(n_206288851));
	notech_reg regs_reg_8_26(.CP(n_62295), .D(n_19259), .CD(n_61214), .Q(regs_8
		[26]));
	notech_mux2 i_5024(.S(n_53982), .A(regs_8[26]), .B(n_13971), .Z(n_19259)
		);
	notech_or4 i_148431634(.A(n_60540), .B(n_60504), .C(n_60558), .D(n_59375
		), .Z(n_206188852));
	notech_reg regs_reg_8_27(.CP(n_62295), .D(n_19266), .CD(n_61214), .Q(regs_8
		[27]));
	notech_mux2 i_5032(.S(n_53982), .A(regs_8[27]), .B(n_13977), .Z(n_19266)
		);
	notech_reg regs_reg_8_28(.CP(n_62295), .D(n_19273), .CD(n_61214), .Q(regs_8
		[28]));
	notech_mux2 i_5040(.S(n_53982), .A(regs_8[28]), .B(n_13983), .Z(n_19273)
		);
	notech_and3 i_51032903(.A(n_1960), .B(n_54874), .C(n_195988889), .Z(n_205988854
		));
	notech_reg regs_reg_8_29(.CP(n_62295), .D(n_19280), .CD(n_61215), .Q(regs_8
		[29]));
	notech_mux2 i_5048(.S(n_53982), .A(regs_8[29]), .B(n_26880), .Z(n_19280)
		);
	notech_nao3 i_80133052(.A(n_57378), .B(n_57374), .C(n_26406), .Z(n_205888855
		));
	notech_reg regs_reg_8_30(.CP(n_62295), .D(n_19286), .CD(n_61216), .Q(regs_8
		[30]));
	notech_mux2 i_5056(.S(n_53982), .A(regs_8[30]), .B(n_13995), .Z(n_19286)
		);
	notech_ao4 i_73933053(.A(n_58931), .B(n_59369), .C(n_2260), .D(n_2352), 
		.Z(n_205788856));
	notech_reg regs_reg_8_31(.CP(n_62295), .D(n_19292), .CD(n_61216), .Q(regs_8
		[31]));
	notech_mux2 i_5064(.S(n_53982), .A(regs_8[31]), .B(n_14001), .Z(n_19292)
		);
	notech_ao3 i_148631632(.A(n_59183), .B(n_59817), .C(n_58940), .Z(n_205688857
		));
	notech_reg regs_reg_7_0(.CP(n_62295), .D(n_19298), .CD(n_61216), .Q(regs_7
		[0]));
	notech_mux2 i_5072(.S(\nbus_11310[0] ), .A(regs_7[0]), .B(n_13467), .Z(n_19298
		));
	notech_nao3 i_120932856(.A(n_2042), .B(n_26867), .C(n_59355), .Z(n_205588858
		));
	notech_reg regs_reg_7_1(.CP(n_62209), .D(n_19304), .CD(n_61216), .Q(regs_7
		[1]));
	notech_mux2 i_5080(.S(\nbus_11310[0] ), .A(regs_7[1]), .B(n_13473), .Z(n_19304
		));
	notech_reg regs_reg_7_2(.CP(n_62209), .D(n_19310), .CD(n_61216), .Q(regs_7
		[2]));
	notech_mux2 i_5088(.S(\nbus_11310[0] ), .A(regs_7[2]), .B(n_13479), .Z(n_19310
		));
	notech_reg regs_reg_7_3(.CP(n_62211), .D(n_19316), .CD(n_61216), .Q(regs_7
		[3]));
	notech_mux2 i_5096(.S(\nbus_11310[0] ), .A(regs_7[3]), .B(n_13485), .Z(n_19316
		));
	notech_reg regs_reg_7_4(.CP(n_62211), .D(n_19322), .CD(n_61216), .Q(regs_7
		[4]));
	notech_mux2 i_5104(.S(\nbus_11310[0] ), .A(regs_7[4]), .B(n_13491), .Z(n_19322
		));
	notech_ao4 i_51433037(.A(n_56573), .B(n_204988864), .C(n_2241), .D(n_26228
		), .Z(n_205188862));
	notech_reg regs_reg_7_5(.CP(n_62211), .D(n_19328), .CD(n_61216), .Q(regs_7
		[5]));
	notech_mux2 i_5112(.S(\nbus_11310[0] ), .A(regs_7[5]), .B(n_13497), .Z(n_19328
		));
	notech_or4 i_164132830(.A(n_60540), .B(n_2007), .C(n_59899), .D(n_60583)
		, .Z(n_205088863));
	notech_reg regs_reg_7_6(.CP(n_62211), .D(n_19334), .CD(n_61216), .Q(regs_7
		[6]));
	notech_mux2 i_5120(.S(\nbus_11310[0] ), .A(regs_7[6]), .B(n_26882), .Z(n_19334
		));
	notech_or2 i_164232829(.A(n_56502), .B(n_60583), .Z(n_204988864));
	notech_reg regs_reg_7_7(.CP(n_62211), .D(n_19340), .CD(n_61215), .Q(regs_7
		[7]));
	notech_mux2 i_5128(.S(\nbus_11310[0] ), .A(regs_7[7]), .B(n_26883), .Z(n_19340
		));
	notech_ao4 i_153431594(.A(n_2252), .B(n_2263), .C(n_1955), .D(n_26322), 
		.Z(n_204888865));
	notech_reg regs_reg_7_8(.CP(n_62211), .D(n_19346), .CD(n_61215), .Q(regs_7
		[8]));
	notech_mux2 i_5136(.S(\nbus_11310[0] ), .A(regs_7[8]), .B(n_13515), .Z(n_19346
		));
	notech_nand2 i_182632819(.A(n_59299), .B(n_28564), .Z(n_204788866));
	notech_reg regs_reg_7_9(.CP(n_62211), .D(n_19352), .CD(n_61215), .Q(regs_7
		[9]));
	notech_mux2 i_5144(.S(\nbus_11310[0] ), .A(regs_7[9]), .B(n_26884), .Z(n_19352
		));
	notech_reg regs_reg_7_10(.CP(n_62211), .D(n_19358), .CD(n_61215), .Q(regs_7
		[10]));
	notech_mux2 i_5152(.S(\nbus_11310[0] ), .A(regs_7[10]), .B(n_26885), .Z(n_19358
		));
	notech_reg regs_reg_7_11(.CP(n_62211), .D(n_19364), .CD(n_61216), .Q(regs_7
		[11]));
	notech_mux2 i_5160(.S(\nbus_11310[0] ), .A(regs_7[11]), .B(n_13533), .Z(n_19364
		));
	notech_nao3 i_1968(.A(n_60540), .B(n_59817), .C(n_2007), .Z(n_2044));
	notech_reg regs_reg_7_12(.CP(n_62211), .D(n_19370), .CD(n_61216), .Q(regs_7
		[12]));
	notech_mux2 i_5168(.S(\nbus_11310[0] ), .A(regs_7[12]), .B(n_13539), .Z(n_19370
		));
	notech_reg regs_reg_7_13(.CP(n_62211), .D(n_19376), .CD(n_61216), .Q(regs_7
		[13]));
	notech_mux2 i_5176(.S(\nbus_11310[0] ), .A(regs_7[13]), .B(n_13545), .Z(n_19376
		));
	notech_and2 i_173632825(.A(n_2340), .B(n_231756227), .Z(n_2042));
	notech_reg regs_reg_7_14(.CP(n_62211), .D(n_19382), .CD(n_61216), .Q(regs_7
		[14]));
	notech_mux2 i_5184(.S(\nbus_11310[0] ), .A(regs_7[14]), .B(n_13551), .Z(n_19382
		));
	notech_ao3 i_153231596(.A(calc_sz[1]), .B(n_27404), .C(calc_sz[2]), .Z(n_2041
		));
	notech_reg regs_reg_7_15(.CP(n_62211), .D(n_19388), .CD(n_61216), .Q(regs_7
		[15]));
	notech_mux2 i_5192(.S(\nbus_11310[0] ), .A(regs_7[15]), .B(n_13557), .Z(n_19388
		));
	notech_reg regs_reg_7_16(.CP(n_62211), .D(n_19394), .CD(n_61214), .Q(regs_7
		[16]));
	notech_mux2 i_5200(.S(n_54004), .A(regs_7[16]), .B(n_13563), .Z(n_19394)
		);
	notech_reg regs_reg_7_17(.CP(n_62211), .D(n_19400), .CD(n_61211), .Q(regs_7
		[17]));
	notech_mux2 i_5208(.S(n_54004), .A(regs_7[17]), .B(n_13569), .Z(n_19400)
		);
	notech_or4 i_154631584(.A(ecx[1]), .B(ecx[0]), .C(ecx[2]), .D(ecx[3]), .Z
		(n_2038));
	notech_reg regs_reg_7_18(.CP(n_62211), .D(n_19406), .CD(n_61211), .Q(regs_7
		[18]));
	notech_mux2 i_5216(.S(n_54004), .A(regs_7[18]), .B(n_13575), .Z(n_19406)
		);
	notech_reg regs_reg_7_19(.CP(n_62211), .D(n_19412), .CD(n_61211), .Q(regs_7
		[19]));
	notech_mux2 i_5224(.S(n_54004), .A(regs_7[19]), .B(n_13581), .Z(n_19412)
		);
	notech_reg regs_reg_7_20(.CP(n_62211), .D(n_19418), .CD(n_61211), .Q(regs_7
		[20]));
	notech_mux2 i_5232(.S(n_54004), .A(regs_7[20]), .B(n_13587), .Z(n_19418)
		);
	notech_or4 i_155031581(.A(ecx[4]), .B(ecx[5]), .C(ecx[6]), .D(ecx[7]), .Z
		(n_2035));
	notech_reg regs_reg_7_21(.CP(n_62211), .D(n_19424), .CD(n_61211), .Q(regs_7
		[21]));
	notech_mux2 i_5240(.S(n_54004), .A(regs_7[21]), .B(n_13593), .Z(n_19424)
		);
	notech_reg regs_reg_7_22(.CP(n_62155), .D(n_19430), .CD(n_61211), .Q(regs_7
		[22]));
	notech_mux2 i_5248(.S(n_54004), .A(regs_7[22]), .B(n_13599), .Z(n_19430)
		);
	notech_reg regs_reg_7_23(.CP(n_62155), .D(n_19436), .CD(n_61211), .Q(regs_7
		[23]));
	notech_mux2 i_5257(.S(n_54004), .A(regs_7[23]), .B(n_13605), .Z(n_19436)
		);
	notech_reg regs_reg_7_24(.CP(n_62155), .D(n_19444), .CD(n_61211), .Q(regs_7
		[24]));
	notech_mux2 i_5265(.S(n_54004), .A(regs_7[24]), .B(n_13611), .Z(n_19444)
		);
	notech_or4 i_155531577(.A(ecx[10]), .B(ecx[8]), .C(ecx[9]), .D(ecx[11]),
		 .Z(n_2031));
	notech_reg regs_reg_7_25(.CP(n_62155), .D(n_19451), .CD(n_61211), .Q(regs_7
		[25]));
	notech_mux2 i_5273(.S(n_54004), .A(regs_7[25]), .B(n_13617), .Z(n_19451)
		);
	notech_reg regs_reg_7_26(.CP(n_62155), .D(n_19458), .CD(n_61210), .Q(regs_7
		[26]));
	notech_mux2 i_5281(.S(n_54004), .A(regs_7[26]), .B(n_13623), .Z(n_19458)
		);
	notech_reg regs_reg_7_27(.CP(n_62155), .D(n_19465), .CD(n_61210), .Q(regs_7
		[27]));
	notech_mux2 i_5289(.S(n_54004), .A(regs_7[27]), .B(n_13629), .Z(n_19465)
		);
	notech_or4 i_156231573(.A(ecx[15]), .B(ecx[12]), .C(ecx[13]), .D(n_2025)
		, .Z(n_2028));
	notech_reg regs_reg_7_28(.CP(n_62155), .D(n_19472), .CD(n_61210), .Q(regs_7
		[28]));
	notech_mux2 i_5297(.S(n_54004), .A(regs_7[28]), .B(n_13635), .Z(n_19472)
		);
	notech_reg regs_reg_7_29(.CP(n_62155), .D(n_19480), .CD(n_61210), .Q(regs_7
		[29]));
	notech_mux2 i_5305(.S(n_54004), .A(regs_7[29]), .B(n_13641), .Z(n_19480)
		);
	notech_reg regs_reg_7_30(.CP(n_62155), .D(n_19487), .CD(n_61210), .Q(regs_7
		[30]));
	notech_mux2 i_5313(.S(n_54004), .A(regs_7[30]), .B(n_13647), .Z(n_19487)
		);
	notech_or2 i_155831575(.A(ecx[14]), .B(n_2010), .Z(n_2025));
	notech_reg regs_reg_7_31(.CP(n_62155), .D(n_19494), .CD(n_61211), .Q(regs_7
		[31]));
	notech_mux2 i_5321(.S(n_54004), .A(regs_7[31]), .B(n_13653), .Z(n_19494)
		);
	notech_reg pipe_mul_reg_0(.CP(n_62205), .D(n_19501), .CD(n_61211), .Q(pipe_mul
		[0]));
	notech_mux2 i_5329(.S(\nbus_11281[0] ), .A(pipe_mul[0]), .B(n_264385963)
		, .Z(n_19501));
	notech_or4 i_156631569(.A(ecx[31]), .B(ecx[30]), .C(ecx[29]), .D(ecx[28]
		), .Z(n_202388868));
	notech_reg pipe_mul_reg_1(.CP(n_62195), .D(n_19508), .CD(n_61210), .Q(pipe_mul
		[1]));
	notech_mux2 i_5337(.S(\nbus_11281[0] ), .A(pipe_mul[1]), .B(n_264485964)
		, .Z(n_19508));
	notech_reg CFOF_mul_reg(.CP(n_62195), .D(n_19516), .CD(n_61210), .Q(CFOF_mul
		));
	notech_mux2 i_5345(.S(n_208741718), .A(n_8721), .B(CFOF_mul), .Z(n_19516
		));
	notech_reg eval_flag_reg(.CP(n_62195), .D(n_19523), .CD(n_61211), .Q(eval_flag
		));
	notech_or2 i_5353(.A(n_19525), .B(n_19526), .Z(n_19523));
	notech_ao4 i_5354(.A(n_55569), .B(n_237985699), .C(n_26589), .D(n_26507)
		, .Z(n_19525));
	notech_and3 i_5355(.A(n_166781655), .B(eval_flag), .C(n_54968), .Z(n_19526
		));
	notech_or4 i_156931566(.A(ecx[26]), .B(ecx[27]), .C(ecx[24]), .D(ecx[25]
		), .Z(n_202088871));
	notech_reg rep_en1_reg(.CP(n_62195), .D(n_19530), .CD(n_61213), .Q(rep_en1
		));
	notech_mux2 i_5361(.S(n_9351), .A(rep_en1), .B(n_59819), .Z(n_19530));
	notech_reg rep_en2_reg(.CP(n_62195), .D(n_19537), .CD(n_61213), .Q(rep_en2
		));
	notech_mux2 i_5369(.S(n_9257), .A(rep_en2), .B(n_59819), .Z(n_19537));
	notech_reg rep_en3_reg(.CP(n_62195), .D(n_19544), .CD(n_61213), .Q(rep_en3
		));
	notech_mux2 i_5379(.S(n_11506), .A(rep_en3), .B(n_59819), .Z(n_19544));
	notech_reg rep_en4_reg(.CP(n_62195), .D(n_19552), .CD(n_61213), .Q(rep_en4
		));
	notech_mux2 i_5388(.S(n_15204), .A(rep_en4), .B(n_59819), .Z(n_19552));
	notech_or4 i_157931562(.A(ecx[23]), .B(ecx[20]), .C(ecx[22]), .D(ecx[21]
		), .Z(n_201688875));
	notech_reg rep_en5_reg(.CP(n_62195), .D(n_19559), .CD(n_61213), .Q(rep_en5
		));
	notech_mux2 i_5397(.S(n_10208), .A(rep_en5), .B(n_59819), .Z(n_19559));
	notech_reg nCF_reg(.CP(n_62195), .D(n_19566), .CD(n_61214), .Q(nCF));
	notech_mux2 i_5407(.S(n_7415), .A(nCF), .B(n_7418), .Z(n_19566));
	notech_reg nPF_reg(.CP(n_62195), .D(n_19574), .CD(n_61214), .Q(nPF));
	notech_mux2 i_5415(.S(n_26893), .A(nPF), .B(n_156774435), .Z(n_19574));
	notech_or4 i_158231559(.A(ecx[18]), .B(ecx[19]), .C(ecx[17]), .D(ecx[16]
		), .Z(n_201388878));
	notech_reg nAF_reg(.CP(n_62195), .D(n_19583), .CD(n_61214), .Q(nAF));
	notech_mux2 i_5423(.S(n_301586335), .A(nAF_arithbox), .B(nAF), .Z(n_19583
		));
	notech_reg nSF_reg(.CP(n_62195), .D(n_19591), .CD(n_61214), .Q(nSF));
	notech_mux2 i_5431(.S(n_300586325), .A(n_18226), .B(nSF), .Z(n_19591));
	notech_reg opas_reg(.CP(n_62271), .D(n_19600), .CD(n_61213), .Q(opas));
	notech_mux2 i_5439(.S(n_301586335), .A(opas_arithbox), .B(opas), .Z(n_19600
		));
	notech_and2 i_73232286(.A(n_1966), .B(n_60130), .Z(n_2010));
	notech_reg opbs_reg(.CP(n_62271), .D(n_19608), .CD(n_61213), .Q(opbs));
	notech_mux2 i_5447(.S(n_301586335), .A(opbs_arithbox), .B(opbs), .Z(n_19608
		));
	notech_reg nOF_reg(.CP(n_62271), .D(n_19616), .CD(n_61211), .Q(nOF));
	notech_mux2 i_5455(.S(n_14930), .A(nOF), .B(n_26895), .Z(n_19616));
	notech_reg regs_reg_15_0(.CP(n_62271), .D(n_19625), .CD(n_61213), .Q(\eflags[0] 
		));
	notech_mux2 i_5463(.S(\nbus_11353[0] ), .A(\eflags[0] ), .B(n_20601), .Z
		(n_19625));
	notech_nao3 i_25655(.A(n_2042), .B(n_2361), .C(n_2385), .Z(n_2007));
	notech_reg regs_reg_15_1(.CP(n_62271), .D(n_19632), .CD(n_61213), .Q(\eflags[1] 
		));
	notech_mux2 i_5471(.S(\nbus_11353[1] ), .A(\eflags[1] ), .B(n_20607), .Z
		(n_19632));
	notech_or4 i_15108(.A(n_260688757), .B(n_2605), .C(n_56354), .D(n_55934)
		, .Z(n_2006));
	notech_reg regs_reg_15_2(.CP(n_62271), .D(n_19639), .CD(n_61213), .Q(\eflags[2] 
		));
	notech_mux2 i_5479(.S(\nbus_11353[2] ), .A(\eflags[2] ), .B(n_20613), .Z
		(n_19639));
	notech_or4 i_25813(.A(n_58913), .B(n_58904), .C(n_60583), .D(n_59899), .Z
		(n_2005));
	notech_reg regs_reg_15_3(.CP(n_62271), .D(n_19646), .CD(n_61213), .Q(\eflags[3] 
		));
	notech_mux2 i_5487(.S(\nbus_11353[1] ), .A(\eflags[3] ), .B(n_20619), .Z
		(n_19646));
	notech_reg regs_reg_15_4(.CP(n_62271), .D(n_19653), .CD(n_61213), .Q(\eflags[4] 
		));
	notech_mux2 i_5495(.S(\nbus_11353[0] ), .A(\eflags[4] ), .B(n_26896), .Z
		(n_19653));
	notech_reg regs_reg_15_5(.CP(n_62271), .D(n_19660), .CD(n_61213), .Q(\eflags[5] 
		));
	notech_mux2 i_5503(.S(\nbus_11353[1] ), .A(\eflags[5] ), .B(n_20631), .Z
		(n_19660));
	notech_reg regs_reg_15_6(.CP(n_62271), .D(n_19667), .CD(n_61202), .Q(\eflags[6] 
		));
	notech_mux2 i_5511(.S(\nbus_11353[6] ), .A(\eflags[6] ), .B(n_20637), .Z
		(n_19667));
	notech_reg regs_reg_15_7(.CP(n_62271), .D(n_19673), .CD(n_61191), .Q(\eflags[7] 
		));
	notech_mux2 i_5519(.S(\nbus_11353[6] ), .A(\eflags[7] ), .B(n_20643), .Z
		(n_19673));
	notech_reg regs_reg_15_8(.CP(n_62271), .D(n_19680), .CD(n_61191), .Q(\eflags[8] 
		));
	notech_mux2 i_5527(.S(\nbus_11353[8] ), .A(\eflags[8] ), .B(n_26897), .Z
		(n_19680));
	notech_reg regs_reg_15_9(.CP(n_62271), .D(n_19687), .CD(n_61191), .Q(ie)
		);
	notech_mux2 i_5535(.S(\nbus_11353[9] ), .A(ie), .B(n_20655), .Z(n_19687)
		);
	notech_reg regs_reg_15_10(.CP(n_62271), .D(n_19694), .CD(n_61191), .Q(\eflags[10] 
		));
	notech_mux2 i_5543(.S(n_26898), .A(n_55460), .B(n_20661), .Z(n_19694));
	notech_reg regs_reg_15_11(.CP(n_62271), .D(n_19700), .CD(n_61191), .Q(\eflags[11] 
		));
	notech_mux2 i_5551(.S(\nbus_11353[6] ), .A(\eflags[11] ), .B(n_20667), .Z
		(n_19700));
	notech_or4 i_63332365(.A(n_58940), .B(n_60494), .C(n_59967), .D(n_59355)
		, .Z(n_199688883));
	notech_reg regs_reg_15_12(.CP(n_62271), .D(n_19706), .CD(n_61192), .Q(\eflags[12] 
		));
	notech_mux2 i_5559(.S(\nbus_11353[12] ), .A(\eflags[12] ), .B(n_20673), 
		.Z(n_19706));
	notech_reg regs_reg_15_13(.CP(n_62271), .D(n_19713), .CD(n_61192), .Q(\eflags[13] 
		));
	notech_mux2 i_5567(.S(\nbus_11353[12] ), .A(\eflags[13] ), .B(n_20679), 
		.Z(n_19713));
	notech_reg regs_reg_15_14(.CP(n_62271), .D(n_19720), .CD(n_61191), .Q(\eflags[14] 
		));
	notech_mux2 i_5575(.S(\nbus_11353[12] ), .A(\eflags[14] ), .B(n_26899), 
		.Z(n_19720));
	notech_reg regs_reg_15_15(.CP(n_62271), .D(n_19726), .CD(n_61192), .Q(\eflags[15] 
		));
	notech_mux2 i_5583(.S(\nbus_11353[1] ), .A(\eflags[15] ), .B(n_20691), .Z
		(n_19726));
	notech_reg regs_reg_15_16(.CP(n_62269), .D(n_19733), .CD(n_61191), .Q(\eflags[16] 
		));
	notech_mux2 i_5591(.S(\nbus_11353[12] ), .A(\eflags[16] ), .B(n_20697), 
		.Z(n_19733));
	notech_nao3 i_63732361(.A(n_244056258), .B(n_26590), .C(n_2582), .Z(n_199188888
		));
	notech_reg regs_reg_15_17(.CP(n_62269), .D(n_19739), .CD(n_61191), .Q(\eflags[17] 
		));
	notech_mux2 i_5599(.S(\nbus_11353[12] ), .A(\eflags[17] ), .B(n_20703), 
		.Z(n_19739));
	notech_nor2 i_64132357(.A(writeio_ack), .B(readio_ack), .Z(n_1990));
	notech_reg regs_reg_15_18(.CP(n_62345), .D(n_19745), .CD(n_61189), .Q(\eflags[18] 
		));
	notech_mux2 i_5607(.S(\nbus_11353[12] ), .A(\eflags[18] ), .B(n_20709), 
		.Z(n_19745));
	notech_and2 i_64832350(.A(nbus_11326[3]), .B(n_57432), .Z(n_1989));
	notech_reg regs_reg_15_19(.CP(n_62345), .D(n_19751), .CD(n_61189), .Q(\eflags[19] 
		));
	notech_mux2 i_5615(.S(\nbus_11353[12] ), .A(\eflags[19] ), .B(n_20715), 
		.Z(n_19751));
	notech_reg regs_reg_15_20(.CP(n_62345), .D(n_19757), .CD(n_61191), .Q(\eflags[20] 
		));
	notech_mux2 i_5623(.S(\nbus_11353[12] ), .A(\eflags[20] ), .B(n_20721), 
		.Z(n_19757));
	notech_reg regs_reg_15_21(.CP(n_62345), .D(n_19763), .CD(n_61191), .Q(\eflags[21] 
		));
	notech_mux2 i_5631(.S(\nbus_11353[12] ), .A(\eflags[21] ), .B(n_20727), 
		.Z(n_19763));
	notech_and3 i_65032349(.A(n_48760), .B(n_1562), .C(opc[3]), .Z(n_1986)
		);
	notech_reg regs_reg_15_22(.CP(n_62345), .D(n_19769), .CD(n_61191), .Q(\eflags[22] 
		));
	notech_mux2 i_5639(.S(\nbus_11353[12] ), .A(\eflags[22] ), .B(n_20733), 
		.Z(n_19769));
	notech_ao4 i_64332355(.A(n_149823485), .B(n_2770), .C(n_26553), .D(n_1953
		), .Z(n_1985));
	notech_reg regs_reg_15_23(.CP(n_62345), .D(n_19775), .CD(n_61191), .Q(\eflags[23] 
		));
	notech_mux2 i_5647(.S(\nbus_11353[12] ), .A(\eflags[23] ), .B(n_20739), 
		.Z(n_19775));
	notech_nao3 i_64232356(.A(n_1951), .B(nbus_11273[0]), .C(n_271488741), .Z
		(n_1984));
	notech_reg regs_reg_15_24(.CP(n_62345), .D(n_19781), .CD(n_61191), .Q(\eflags[24] 
		));
	notech_mux2 i_5655(.S(\nbus_11353[12] ), .A(\eflags[24] ), .B(n_20745), 
		.Z(n_19781));
	notech_reg regs_reg_15_25(.CP(n_62345), .D(n_19788), .CD(n_61192), .Q(\eflags[25] 
		));
	notech_mux2 i_5663(.S(\nbus_11353[12] ), .A(\eflags[25] ), .B(n_26900), 
		.Z(n_19788));
	notech_reg regs_reg_15_26(.CP(n_62345), .D(n_19795), .CD(n_61193), .Q(\eflags[26] 
		));
	notech_mux2 i_5671(.S(\nbus_11353[12] ), .A(\eflags[26] ), .B(n_26901), 
		.Z(n_19795));
	notech_or4 i_62132377(.A(n_60602), .B(n_60583), .C(n_59899), .D(n_2226),
		 .Z(n_1981));
	notech_reg regs_reg_15_27(.CP(n_62345), .D(n_19802), .CD(n_61193), .Q(\eflags[27] 
		));
	notech_mux2 i_5679(.S(\nbus_11353[12] ), .A(\eflags[27] ), .B(n_26902), 
		.Z(n_19802));
	notech_reg regs_reg_15_28(.CP(n_62345), .D(n_19810), .CD(n_61193), .Q(\eflags[28] 
		));
	notech_mux2 i_5687(.S(\nbus_11353[12] ), .A(\eflags[28] ), .B(n_26903), 
		.Z(n_19810));
	notech_reg regs_reg_15_29(.CP(n_62345), .D(n_19817), .CD(n_61193), .Q(\eflags[29] 
		));
	notech_mux2 i_5695(.S(\nbus_11353[12] ), .A(\eflags[29] ), .B(n_20775), 
		.Z(n_19817));
	notech_reg regs_reg_15_30(.CP(n_62345), .D(n_19824), .CD(n_61193), .Q(\eflags[30] 
		));
	notech_mux2 i_5703(.S(\nbus_11353[12] ), .A(\eflags[30] ), .B(n_20781), 
		.Z(n_19824));
	notech_reg regs_reg_15_31(.CP(n_62345), .D(n_19831), .CD(n_61193), .Q(\eflags[31] 
		));
	notech_mux2 i_5711(.S(\nbus_11353[12] ), .A(\eflags[31] ), .B(n_20787), 
		.Z(n_19831));
	notech_nand2 i_27130(.A(n_56469), .B(n_56460), .Z(n_1976));
	notech_reg regs_reg_6_0(.CP(n_62345), .D(n_19838), .CD(n_61193), .Q(regs_6
		[0]));
	notech_mux2 i_5719(.S(\nbus_11331[0] ), .A(regs_6[0]), .B(n_16350), .Z(n_19838
		));
	notech_reg regs_reg_6_1(.CP(n_62345), .D(n_19846), .CD(n_61193), .Q(regs_6
		[1]));
	notech_mux2 i_5727(.S(\nbus_11331[0] ), .A(regs_6[1]), .B(n_16356), .Z(n_19846
		));
	notech_reg regs_reg_6_2(.CP(n_62345), .D(n_19853), .CD(n_61193), .Q(regs_6
		[2]));
	notech_mux2 i_5735(.S(\nbus_11331[0] ), .A(regs_6[2]), .B(n_16362), .Z(n_19853
		));
	notech_or4 i_11332766(.A(n_1909), .B(n_60516), .C(n_60527), .D(n_28571),
		 .Z(n_1973));
	notech_reg regs_reg_6_3(.CP(n_62345), .D(n_19860), .CD(n_61192), .Q(regs_6
		[3]));
	notech_mux2 i_5743(.S(\nbus_11331[0] ), .A(regs_6[3]), .B(n_26904), .Z(n_19860
		));
	notech_nand2 i_32069(.A(n_274788710), .B(n_59899), .Z(n_1972));
	notech_reg regs_reg_6_4(.CP(n_62269), .D(n_19867), .CD(n_61192), .Q(regs_6
		[4]));
	notech_mux2 i_5751(.S(\nbus_11331[0] ), .A(regs_6[4]), .B(n_16374), .Z(n_19867
		));
	notech_reg regs_reg_6_5(.CP(n_62269), .D(n_19874), .CD(n_61192), .Q(regs_6
		[5]));
	notech_mux2 i_5759(.S(\nbus_11331[0] ), .A(regs_6[5]), .B(n_26905), .Z(n_19874
		));
	notech_nand2 i_27360(.A(n_205888855), .B(n_26592), .Z(n_1970));
	notech_reg regs_reg_6_6(.CP(n_62269), .D(n_19882), .CD(n_61192), .Q(regs_6
		[6]));
	notech_mux2 i_5767(.S(\nbus_11331[0] ), .A(regs_6[6]), .B(n_26906), .Z(n_19882
		));
	notech_nor2 i_29683(.A(n_57383), .B(n_274488713), .Z(n_1969));
	notech_reg regs_reg_6_7(.CP(n_62269), .D(n_19889), .CD(n_61192), .Q(regs_6
		[7]));
	notech_mux2 i_5775(.S(\nbus_11331[0] ), .A(regs_6[7]), .B(n_26907), .Z(n_19889
		));
	notech_or4 i_29739(.A(n_59369), .B(n_60494), .C(n_60768), .D(n_60724), .Z
		(n_1968));
	notech_reg regs_reg_6_8(.CP(n_62269), .D(n_19896), .CD(n_61192), .Q(regs_6
		[8]));
	notech_mux2 i_5783(.S(\nbus_11331[0] ), .A(regs_6[8]), .B(n_16398), .Z(n_19896
		));
	notech_or4 i_30881(.A(n_60752), .B(n_60739), .C(n_60768), .D(n_59201), .Z
		(n_1967));
	notech_reg regs_reg_6_9(.CP(n_62269), .D(n_19903), .CD(n_61192), .Q(regs_6
		[9]));
	notech_mux2 i_5791(.S(\nbus_11331[0] ), .A(regs_6[9]), .B(n_26908), .Z(n_19903
		));
	notech_or4 i_15832721(.A(n_202388868), .B(n_202088871), .C(n_201688875),
		 .D(n_201388878), .Z(n_1966));
	notech_reg regs_reg_6_10(.CP(n_62269), .D(n_19910), .CD(n_61192), .Q(regs_6
		[10]));
	notech_mux2 i_5799(.S(\nbus_11331[0] ), .A(regs_6[10]), .B(n_26909), .Z(n_19910
		));
	notech_reg regs_reg_6_11(.CP(n_62269), .D(n_19918), .CD(n_61192), .Q(regs_6
		[11]));
	notech_mux2 i_5807(.S(\nbus_11331[0] ), .A(regs_6[11]), .B(n_16416), .Z(n_19918
		));
	notech_reg regs_reg_6_12(.CP(n_62269), .D(n_19925), .CD(n_61189), .Q(regs_6
		[12]));
	notech_mux2 i_5815(.S(\nbus_11331[0] ), .A(regs_6[12]), .B(n_16422), .Z(n_19925
		));
	notech_or4 i_71832294(.A(n_260688757), .B(n_2605), .C(n_56354), .D(n_26228
		), .Z(n_1963));
	notech_reg regs_reg_6_13(.CP(n_62269), .D(n_19932), .CD(n_61187), .Q(regs_6
		[13]));
	notech_mux2 i_5823(.S(\nbus_11331[0] ), .A(regs_6[13]), .B(n_16428), .Z(n_19932
		));
	notech_and4 i_71732295(.A(n_55846), .B(n_1963), .C(n_205188862), .D(n_55834
		), .Z(n_1962));
	notech_reg regs_reg_6_14(.CP(n_62345), .D(n_19939), .CD(n_61187), .Q(regs_6
		[14]));
	notech_mux2 i_5831(.S(\nbus_11331[0] ), .A(regs_6[14]), .B(n_26910), .Z(n_19939
		));
	notech_and3 i_16132718(.A(n_205788856), .B(n_57375), .C(n_57374), .Z(n_1961
		));
	notech_reg regs_reg_6_15(.CP(n_62267), .D(n_19946), .CD(n_61187), .Q(regs_6
		[15]));
	notech_mux2 i_5839(.S(\nbus_11331[0] ), .A(regs_6[15]), .B(n_16440), .Z(n_19946
		));
	notech_or4 i_71532296(.A(n_60768), .B(n_60721), .C(n_60584), .D(n_1961),
		 .Z(n_1960));
	notech_reg regs_reg_6_16(.CP(n_62267), .D(n_19954), .CD(n_61187), .Q(regs_6
		[16]));
	notech_mux2 i_5847(.S(n_54035), .A(regs_6[16]), .B(n_16446), .Z(n_19954)
		);
	notech_or4 i_71232297(.A(n_2258), .B(n_2180), .C(n_60584), .D(n_59899), 
		.Z(n_195988889));
	notech_reg regs_reg_6_17(.CP(n_62341), .D(n_19961), .CD(n_61187), .Q(regs_6
		[17]));
	notech_mux2 i_5855(.S(n_54035), .A(regs_6[17]), .B(n_16452), .Z(n_19961)
		);
	notech_or4 i_71132298(.A(n_57380), .B(cond_1), .C(n_60584), .D(n_59898),
		 .Z(n_1958));
	notech_reg regs_reg_6_18(.CP(n_62341), .D(n_19968), .CD(n_61188), .Q(regs_6
		[18]));
	notech_mux2 i_5863(.S(n_54035), .A(regs_6[18]), .B(n_16458), .Z(n_19968)
		);
	notech_reg regs_reg_6_19(.CP(n_62341), .D(n_19975), .CD(n_61188), .Q(regs_6
		[19]));
	notech_mux2 i_5871(.S(n_54035), .A(regs_6[19]), .B(n_16464), .Z(n_19975)
		);
	notech_reg regs_reg_6_20(.CP(n_62341), .D(n_19981), .CD(n_61188), .Q(regs_6
		[20]));
	notech_mux2 i_5879(.S(n_54035), .A(regs_6[20]), .B(n_16470), .Z(n_19981)
		);
	notech_ao4 i_180732820(.A(n_59375), .B(n_62405), .C(n_2252), .D(n_2264),
		 .Z(n_1955));
	notech_reg regs_reg_6_21(.CP(n_62341), .D(n_19987), .CD(n_61188), .Q(regs_6
		[21]));
	notech_mux2 i_5887(.S(n_54035), .A(regs_6[21]), .B(n_16476), .Z(n_19987)
		);
	notech_and4 i_65132348(.A(n_2172), .B(n_2162), .C(n_2153), .D(n_214888806
		), .Z(n_1954));
	notech_reg regs_reg_6_22(.CP(n_62341), .D(n_19993), .CD(n_61187), .Q(regs_6
		[22]));
	notech_mux2 i_5895(.S(n_54035), .A(regs_6[22]), .B(n_16482), .Z(n_19993)
		);
	notech_ao3 i_64532353(.A(rep_en5), .B(n_58951), .C(n_270588748), .Z(n_1953
		));
	notech_reg regs_reg_6_23(.CP(n_62341), .D(n_19999), .CD(n_61187), .Q(regs_6
		[23]));
	notech_mux2 i_5903(.S(n_54035), .A(regs_6[23]), .B(n_16488), .Z(n_19999)
		);
	notech_reg regs_reg_6_24(.CP(n_62341), .D(n_20005), .CD(n_61186), .Q(regs_6
		[24]));
	notech_mux2 i_5911(.S(n_54035), .A(regs_6[24]), .B(n_16494), .Z(n_20005)
		);
	notech_or4 i_12332756(.A(n_2708), .B(n_1986), .C(n_1989), .D(n_213688808
		), .Z(n_1951));
	notech_reg regs_reg_6_25(.CP(n_62341), .D(n_20011), .CD(n_61187), .Q(regs_6
		[25]));
	notech_mux2 i_5919(.S(n_54035), .A(regs_6[25]), .B(n_16500), .Z(n_20011)
		);
	notech_or4 i_64032358(.A(n_62427), .B(\opcode[3] ), .C(\opcode[0] ), .D(\opcode[1] 
		), .Z(n_1950));
	notech_reg regs_reg_6_26(.CP(n_62341), .D(n_20017), .CD(n_61187), .Q(regs_6
		[26]));
	notech_mux2 i_5927(.S(n_54035), .A(regs_6[26]), .B(n_16506), .Z(n_20017)
		);
	notech_nao3 i_63632362(.A(start_up), .B(n_26773), .C(n_26616), .Z(n_1949
		));
	notech_reg regs_reg_6_27(.CP(n_62383), .D(n_20023), .CD(n_61187), .Q(regs_6
		[27]));
	notech_mux2 i_5935(.S(n_54035), .A(regs_6[27]), .B(n_16512), .Z(n_20023)
		);
	notech_reg regs_reg_6_28(.CP(n_62383), .D(n_20029), .CD(n_61187), .Q(regs_6
		[28]));
	notech_mux2 i_5943(.S(n_54035), .A(regs_6[28]), .B(n_16518), .Z(n_20029)
		);
	notech_nand2 i_63432364(.A(n_55843), .B(n_57384), .Z(n_1947));
	notech_reg regs_reg_6_29(.CP(n_62383), .D(n_20035), .CD(n_61187), .Q(regs_6
		[29]));
	notech_mux2 i_5951(.S(n_54035), .A(regs_6[29]), .B(n_16524), .Z(n_20035)
		);
	notech_reg regs_reg_6_30(.CP(n_62383), .D(n_20041), .CD(n_61187), .Q(regs_6
		[30]));
	notech_mux2 i_5959(.S(n_54035), .A(regs_6[30]), .B(n_26911), .Z(n_20041)
		);
	notech_and3 i_16232717(.A(n_55644), .B(n_2236), .C(n_51738), .Z(n_1945)
		);
	notech_reg regs_reg_6_31(.CP(n_62383), .D(n_20047), .CD(n_61188), .Q(regs_6
		[31]));
	notech_mux2 i_5967(.S(n_54035), .A(regs_6[31]), .B(n_16536), .Z(n_20047)
		);
	notech_or4 i_19632710(.A(n_210388836), .B(n_2091), .C(n_2085), .D(n_2080
		), .Z(n_1944));
	notech_reg regs_reg_5_0(.CP(n_62383), .D(n_20053), .CD(n_61189), .Q(regs_5
		[0]));
	notech_mux2 i_5975(.S(\nbus_11309[0] ), .A(regs_5[0]), .B(n_26912), .Z(n_20053
		));
	notech_ao4 i_19532711(.A(n_59281), .B(n_59250), .C(n_29040), .D(n_59219)
		, .Z(n_1943));
	notech_reg regs_reg_5_1(.CP(n_62383), .D(n_20059), .CD(n_61189), .Q(regs_5
		[1]));
	notech_mux2 i_5983(.S(\nbus_11309[0] ), .A(regs_5[1]), .B(n_26913), .Z(n_20059
		));
	notech_nand3 i_62732371(.A(n_59762), .B(n_59369), .C(n_59201), .Z(n_1942
		));
	notech_reg regs_reg_5_2(.CP(n_62383), .D(n_20065), .CD(n_61189), .Q(regs_5
		[2]));
	notech_mux2 i_5991(.S(\nbus_11309[0] ), .A(regs_5[2]), .B(n_26914), .Z(n_20065
		));
	notech_and2 i_11232767(.A(n_2072), .B(n_207188842), .Z(n_1941));
	notech_reg regs_reg_5_3(.CP(n_62383), .D(n_20071), .CD(n_61189), .Q(regs_5
		[3]));
	notech_mux2 i_5999(.S(\nbus_11309[0] ), .A(regs_5[3]), .B(n_13133), .Z(n_20071
		));
	notech_and3 i_11132768(.A(n_206788846), .B(n_60752), .C(n_60739), .Z(n_1940
		));
	notech_reg regs_reg_5_4(.CP(n_62383), .D(n_20077), .CD(n_61189), .Q(regs_5
		[4]));
	notech_mux2 i_6007(.S(\nbus_11309[0] ), .A(regs_5[4]), .B(n_26915), .Z(n_20077
		));
	notech_reg regs_reg_5_5(.CP(n_62383), .D(n_20083), .CD(n_61189), .Q(regs_5
		[5]));
	notech_mux2 i_6015(.S(\nbus_11309[0] ), .A(regs_5[5]), .B(n_13145), .Z(n_20083
		));
	notech_reg regs_reg_5_6(.CP(n_62383), .D(n_20089), .CD(n_61189), .Q(regs_5
		[6]));
	notech_mux2 i_6023(.S(\nbus_11309[0] ), .A(regs_5[6]), .B(n_26916), .Z(n_20089
		));
	notech_reg regs_reg_5_7(.CP(n_62383), .D(n_20095), .CD(n_61189), .Q(regs_5
		[7]));
	notech_mux2 i_6031(.S(\nbus_11309[0] ), .A(regs_5[7]), .B(n_26917), .Z(n_20095
		));
	notech_ao4 i_179732821(.A(n_59375), .B(n_62405), .C(n_2264), .D(n_26229)
		, .Z(n_1936));
	notech_reg regs_reg_5_8(.CP(n_62383), .D(n_20101), .CD(n_61189), .Q(regs_5
		[8]));
	notech_mux2 i_6039(.S(\nbus_11309[0] ), .A(regs_5[8]), .B(n_13163), .Z(n_20101
		));
	notech_reg regs_reg_5_9(.CP(n_62383), .D(n_20107), .CD(n_61188), .Q(regs_5
		[9]));
	notech_mux2 i_6047(.S(\nbus_11309[0] ), .A(regs_5[9]), .B(n_13169), .Z(n_20107
		));
	notech_nao3 i_61132386(.A(n_59230), .B(n_57162), .C(n_1916), .Z(n_1934)
		);
	notech_reg regs_reg_5_10(.CP(n_62383), .D(n_20114), .CD(n_61188), .Q(regs_5
		[10]));
	notech_mux2 i_6055(.S(\nbus_11309[0] ), .A(regs_5[10]), .B(n_13175), .Z(n_20114
		));
	notech_reg regs_reg_5_11(.CP(n_62383), .D(n_20121), .CD(n_61188), .Q(regs_5
		[11]));
	notech_mux2 i_6064(.S(\nbus_11309[0] ), .A(regs_5[11]), .B(n_13181), .Z(n_20121
		));
	notech_nao3 i_11432765(.A(n_59230), .B(n_56079), .C(n_273888717), .Z(n_1932
		));
	notech_reg regs_reg_5_12(.CP(n_62383), .D(n_20128), .CD(n_61188), .Q(regs_5
		[12]));
	notech_mux2 i_6072(.S(\nbus_11309[0] ), .A(regs_5[12]), .B(n_13187), .Z(n_20128
		));
	notech_and4 i_60932388(.A(n_56305), .B(n_1934), .C(n_1973), .D(n_1932), 
		.Z(n_1931));
	notech_reg regs_reg_5_13(.CP(n_62341), .D(n_20136), .CD(n_61188), .Q(regs_5
		[13]));
	notech_mux2 i_6080(.S(\nbus_11309[0] ), .A(regs_5[13]), .B(n_13193), .Z(n_20136
		));
	notech_reg regs_reg_5_14(.CP(n_62383), .D(n_20143), .CD(n_61188), .Q(regs_5
		[14]));
	notech_mux2 i_6088(.S(\nbus_11309[0] ), .A(regs_5[14]), .B(n_13199), .Z(n_20143
		));
	notech_reg regs_reg_5_15(.CP(n_62343), .D(n_20150), .CD(n_61189), .Q(regs_5
		[15]));
	notech_mux2 i_6096(.S(\nbus_11309[0] ), .A(regs_5[15]), .B(n_26918), .Z(n_20150
		));
	notech_reg regs_reg_5_16(.CP(n_62343), .D(n_20157), .CD(n_61188), .Q(regs_5
		[16]));
	notech_mux2 i_6104(.S(n_54055), .A(regs_5[16]), .B(n_13211), .Z(n_20157)
		);
	notech_reg regs_reg_5_17(.CP(n_62343), .D(n_20164), .CD(n_61188), .Q(regs_5
		[17]));
	notech_mux2 i_6112(.S(n_54055), .A(regs_5[17]), .B(n_13217), .Z(n_20164)
		);
	notech_reg regs_reg_5_18(.CP(n_62343), .D(n_20172), .CD(n_61193), .Q(regs_5
		[18]));
	notech_mux2 i_6120(.S(n_54055), .A(regs_5[18]), .B(n_13223), .Z(n_20172)
		);
	notech_reg regs_reg_5_19(.CP(n_62343), .D(n_20179), .CD(n_61199), .Q(regs_5
		[19]));
	notech_mux2 i_6128(.S(n_54055), .A(regs_5[19]), .B(n_13229), .Z(n_20179)
		);
	notech_reg regs_reg_5_20(.CP(n_62343), .D(n_20186), .CD(n_61199), .Q(regs_5
		[20]));
	notech_mux2 i_6136(.S(n_54055), .A(regs_5[20]), .B(n_13235), .Z(n_20186)
		);
	notech_reg regs_reg_5_21(.CP(n_62343), .D(n_20193), .CD(n_61199), .Q(regs_5
		[21]));
	notech_mux2 i_6144(.S(n_54055), .A(regs_5[21]), .B(n_13241), .Z(n_20193)
		);
	notech_and2 i_49932463(.A(n_48299), .B(n_54899), .Z(n_192288896));
	notech_reg regs_reg_5_22(.CP(n_62343), .D(n_20200), .CD(n_61199), .Q(regs_5
		[22]));
	notech_mux2 i_6152(.S(n_54055), .A(regs_5[22]), .B(n_26919), .Z(n_20200)
		);
	notech_and3 i_49032469(.A(n_2776), .B(n_54777), .C(n_57391), .Z(n_192188897
		));
	notech_reg regs_reg_5_23(.CP(n_62343), .D(n_20208), .CD(n_61199), .Q(regs_5
		[23]));
	notech_mux2 i_6160(.S(n_54055), .A(regs_5[23]), .B(n_13253), .Z(n_20208)
		);
	notech_and4 i_19432712(.A(n_57414), .B(n_2269), .C(n_2106), .D(n_1862), 
		.Z(n_192088898));
	notech_reg regs_reg_5_24(.CP(n_62343), .D(n_20215), .CD(n_61199), .Q(regs_5
		[24]));
	notech_mux2 i_6168(.S(n_54055), .A(regs_5[24]), .B(n_13259), .Z(n_20215)
		);
	notech_nand2 i_16867(.A(n_58922), .B(n_211588829), .Z(n_1919));
	notech_reg regs_reg_5_25(.CP(n_62343), .D(n_20222), .CD(n_61200), .Q(regs_5
		[25]));
	notech_mux2 i_6176(.S(n_54055), .A(regs_5[25]), .B(n_13265), .Z(n_20222)
		);
	notech_ao3 i_162632833(.A(n_212188823), .B(n_2176), .C(n_26510), .Z(n_1918
		));
	notech_reg regs_reg_5_26(.CP(n_62343), .D(n_20229), .CD(n_61199), .Q(regs_5
		[26]));
	notech_mux2 i_6184(.S(n_54055), .A(regs_5[26]), .B(n_13271), .Z(n_20229)
		);
	notech_reg regs_reg_5_27(.CP(n_62343), .D(n_20236), .CD(n_61199), .Q(regs_5
		[27]));
	notech_mux2 i_6192(.S(n_54055), .A(regs_5[27]), .B(n_13277), .Z(n_20236)
		);
	notech_nand3 i_161532837(.A(instrc[123]), .B(n_59241), .C(instrc[120]), 
		.Z(n_1916));
	notech_reg regs_reg_5_28(.CP(n_62343), .D(n_20244), .CD(n_61198), .Q(regs_5
		[28]));
	notech_mux2 i_6200(.S(n_54055), .A(regs_5[28]), .B(n_13283), .Z(n_20244)
		);
	notech_nand3 i_161432838(.A(n_205988854), .B(n_1958), .C(n_1949), .Z(n_1915
		));
	notech_reg regs_reg_5_29(.CP(n_62343), .D(n_20251), .CD(n_61198), .Q(regs_5
		[29]));
	notech_mux2 i_6208(.S(n_54055), .A(regs_5[29]), .B(n_13289), .Z(n_20251)
		);
	notech_and4 i_159832839(.A(n_2113), .B(n_55634), .C(n_199188888), .D(n_26751
		), .Z(n_1914));
	notech_reg regs_reg_5_30(.CP(n_62343), .D(n_20258), .CD(n_61198), .Q(regs_5
		[30]));
	notech_mux2 i_6216(.S(n_54055), .A(regs_5[30]), .B(n_26920), .Z(n_20258)
		);
	notech_nand3 i_157832841(.A(n_60549), .B(n_60516), .C(instrc[120]), .Z(n_1913
		));
	notech_reg regs_reg_5_31(.CP(n_62343), .D(n_20265), .CD(n_61198), .Q(regs_5
		[31]));
	notech_mux2 i_6224(.S(n_54055), .A(regs_5[31]), .B(n_13301), .Z(n_20265)
		);
	notech_nao3 i_149332845(.A(n_60516), .B(instrc[120]), .C(n_60549), .Z(n_1912
		));
	notech_reg sav_cs_reg_0(.CP(n_62343), .D(n_20272), .CD(n_61199), .Q(sav_cs
		[0]));
	notech_mux2 i_6232(.S(n_301486334), .A(cs[0]), .B(sav_cs[0]), .Z(n_20272
		));
	notech_nao3 i_125032852(.A(n_2042), .B(n_26867), .C(n_59210), .Z(n_1911)
		);
	notech_reg sav_cs_reg_1(.CP(n_62343), .D(n_20280), .CD(n_61199), .Q(sav_cs
		[1]));
	notech_mux2 i_6240(.S(n_301486334), .A(cs[1]), .B(sav_cs[1]), .Z(n_20280
		));
	notech_nand3 i_111232864(.A(n_59183), .B(n_59898), .C(n_2225), .Z(n_1910
		));
	notech_reg tss_esp0_reg(.CP(n_62267), .D(n_20287), .CD(n_61199), .Q(tss_esp0
		));
	notech_mux2 i_6248(.S(n_26921), .A(tss_esp0), .B(n_59819), .Z(n_20287)
		);
	notech_nand2 i_110132866(.A(n_60549), .B(n_28566), .Z(n_1909));
	notech_reg_set temp_sp_reg_0(.CP(n_62267), .D(n_20294), .SD(1'b1), .Q(temp_sp
		[0]));
	notech_mux2 i_6256(.S(\nbus_11323[0] ), .A(temp_sp[0]), .B(n_26922), .Z(n_20294
		));
	notech_or4 i_102832873(.A(n_60752), .B(n_60739), .C(n_60768), .D(n_59762
		), .Z(n_1908));
	notech_reg_set temp_sp_reg_1(.CP(n_62267), .D(n_20301), .SD(1'b1), .Q(temp_sp
		[1]));
	notech_mux2 i_6264(.S(\nbus_11323[0] ), .A(temp_sp[1]), .B(n_26924), .Z(n_20301
		));
	notech_nand2 i_100032874(.A(n_59898), .B(n_26862), .Z(n_1907));
	notech_reg_set temp_sp_reg_2(.CP(n_62267), .D(n_20307), .SD(1'b1), .Q(temp_sp
		[2]));
	notech_mux2 i_6272(.S(\nbus_11323[0] ), .A(temp_sp[2]), .B(n_26926), .Z(n_20307
		));
	notech_ao4 i_72832886(.A(n_57423), .B(n_59898), .C(n_1972), .D(n_2200), 
		.Z(n_190688899));
	notech_reg_set temp_sp_reg_3(.CP(n_62267), .D(n_20313), .SD(1'b1), .Q(temp_sp
		[3]));
	notech_mux2 i_6280(.S(\nbus_11323[0] ), .A(temp_sp[3]), .B(n_26928), .Z(n_20313
		));
	notech_and2 i_1986(.A(n_204888865), .B(n_56260), .Z(n_190588900));
	notech_reg_set temp_sp_reg_4(.CP(n_62267), .D(n_20319), .SD(1'b1), .Q(temp_sp
		[4]));
	notech_mux2 i_6288(.S(\nbus_11323[0] ), .A(temp_sp[4]), .B(n_26930), .Z(n_20319
		));
	notech_and4 i_60532893(.A(n_60748), .B(n_60735), .C(n_26616), .D(n_206788846
		), .Z(n_190488901));
	notech_reg_set temp_sp_reg_5(.CP(n_62267), .D(n_20325), .SD(1'b1), .Q(temp_sp
		[5]));
	notech_mux2 i_6296(.S(\nbus_11323[0] ), .A(temp_sp[5]), .B(n_26932), .Z(n_20325
		));
	notech_nao3 i_56532894(.A(n_59183), .B(n_59898), .C(n_275088707), .Z(n_190388902
		));
	notech_reg_set temp_sp_reg_6(.CP(n_62267), .D(n_20331), .SD(1'b1), .Q(temp_sp
		[6]));
	notech_mux2 i_6304(.S(\nbus_11323[0] ), .A(temp_sp[6]), .B(n_26934), .Z(n_20331
		));
	notech_and2 i_51732902(.A(n_55846), .B(n_1963), .Z(n_190288903));
	notech_reg_set temp_sp_reg_7(.CP(n_62267), .D(n_20337), .SD(1'b1), .Q(temp_sp
		[7]));
	notech_mux2 i_6312(.S(\nbus_11323[0] ), .A(temp_sp[7]), .B(n_26936), .Z(n_20337
		));
	notech_or4 i_25332918(.A(n_60490), .B(n_59967), .C(n_60558), .D(\opcode[1] 
		), .Z(n_1901));
	notech_reg_set temp_sp_reg_8(.CP(n_62267), .D(n_20343), .SD(1'b1), .Q(temp_sp
		[8]));
	notech_mux2 i_6320(.S(\nbus_11323[0] ), .A(temp_sp[8]), .B(n_26938), .Z(n_20343
		));
	notech_nao3 i_2174(.A(n_2042), .B(n_26867), .C(n_2196), .Z(n_1900));
	notech_reg_set temp_sp_reg_9(.CP(n_62341), .D(n_20349), .SD(1'b1), .Q(temp_sp
		[9]));
	notech_mux2 i_6328(.S(\nbus_11323[0] ), .A(temp_sp[9]), .B(n_26940), .Z(n_20349
		));
	notech_and2 i_188033007(.A(n_27517), .B(n_27518), .Z(n_1899));
	notech_reg_set temp_sp_reg_10(.CP(n_62335), .D(n_20355), .SD(1'b1), .Q(temp_sp
		[10]));
	notech_mux2 i_6336(.S(\nbus_11323[0] ), .A(temp_sp[10]), .B(n_26942), .Z
		(n_20355));
	notech_or4 i_15100(.A(n_55087), .B(n_1955), .C(n_59241), .D(n_190288903)
		, .Z(n_1898));
	notech_reg_set temp_sp_reg_11(.CP(n_62335), .D(n_20361), .SD(1'b1), .Q(temp_sp
		[11]));
	notech_mux2 i_6344(.S(\nbus_11323[0] ), .A(temp_sp[11]), .B(n_26944), .Z
		(n_20361));
	notech_nor2 i_15102(.A(n_190288903), .B(n_190588900), .Z(n_1897));
	notech_reg_set temp_sp_reg_12(.CP(n_62335), .D(n_20367), .SD(1'b1), .Q(temp_sp
		[12]));
	notech_mux2 i_6352(.S(\nbus_11323[0] ), .A(temp_sp[12]), .B(n_26946), .Z
		(n_20367));
	notech_reg_set temp_sp_reg_13(.CP(n_62335), .D(n_20373), .SD(1'b1), .Q(temp_sp
		[13]));
	notech_mux2 i_6360(.S(\nbus_11323[0] ), .A(temp_sp[13]), .B(n_26948), .Z
		(n_20373));
	notech_or4 i_215633613(.A(opa[16]), .B(opa[17]), .C(opa[18]), .D(opa[19]
		), .Z(n_1895));
	notech_reg_set temp_sp_reg_14(.CP(n_62335), .D(n_20379), .SD(1'b1), .Q(temp_sp
		[14]));
	notech_mux2 i_6368(.S(\nbus_11323[0] ), .A(temp_sp[14]), .B(n_26950), .Z
		(n_20379));
	notech_reg_set temp_sp_reg_15(.CP(n_62335), .D(n_20385), .SD(1'b1), .Q(temp_sp
		[15]));
	notech_mux2 i_6377(.S(\nbus_11323[0] ), .A(temp_sp[15]), .B(n_26952), .Z
		(n_20385));
	notech_reg_set temp_sp_reg_16(.CP(n_62335), .D(n_20391), .SD(1'b1), .Q(temp_sp
		[16]));
	notech_mux2 i_6385(.S(n_53661), .A(temp_sp[16]), .B(n_26954), .Z(n_20391
		));
	notech_or4 i_215933610(.A(opa[20]), .B(opa[21]), .C(opa[22]), .D(opa[23]
		), .Z(n_1892));
	notech_reg_set temp_sp_reg_17(.CP(n_62335), .D(n_20397), .SD(1'b1), .Q(temp_sp
		[17]));
	notech_mux2 i_6393(.S(n_53661), .A(temp_sp[17]), .B(n_26956), .Z(n_20397
		));
	notech_reg_set temp_sp_reg_18(.CP(n_62335), .D(n_20403), .SD(1'b1), .Q(temp_sp
		[18]));
	notech_mux2 i_6402(.S(n_53661), .A(temp_sp[18]), .B(n_26958), .Z(n_20403
		));
	notech_reg_set temp_sp_reg_19(.CP(n_62335), .D(n_20409), .SD(1'b1), .Q(temp_sp
		[19]));
	notech_mux2 i_6410(.S(n_53661), .A(temp_sp[19]), .B(n_26960), .Z(n_20409
		));
	notech_reg_set temp_sp_reg_20(.CP(n_62335), .D(n_20415), .SD(1'b1), .Q(temp_sp
		[20]));
	notech_mux2 i_6418(.S(n_53661), .A(temp_sp[20]), .B(n_26962), .Z(n_20415
		));
	notech_or4 i_216333606(.A(opa[24]), .B(opa[25]), .C(opa[26]), .D(opa[27]
		), .Z(n_1888));
	notech_reg_set temp_sp_reg_21(.CP(n_62335), .D(n_20421), .SD(1'b1), .Q(temp_sp
		[21]));
	notech_mux2 i_6426(.S(n_53661), .A(temp_sp[21]), .B(n_26964), .Z(n_20421
		));
	notech_reg_set temp_sp_reg_22(.CP(n_62379), .D(n_20427), .SD(1'b1), .Q(temp_sp
		[22]));
	notech_mux2 i_6434(.S(n_53661), .A(temp_sp[22]), .B(n_26966), .Z(n_20427
		));
	notech_reg_set temp_sp_reg_23(.CP(n_62379), .D(n_20433), .SD(1'b1), .Q(temp_sp
		[23]));
	notech_mux2 i_6443(.S(n_53661), .A(temp_sp[23]), .B(n_26968), .Z(n_20433
		));
	notech_or4 i_216633603(.A(opa[28]), .B(opa[29]), .C(opa[30]), .D(opa[31]
		), .Z(n_1885));
	notech_reg_set temp_sp_reg_24(.CP(n_62379), .D(n_20439), .SD(1'b1), .Q(temp_sp
		[24]));
	notech_mux2 i_6451(.S(n_53661), .A(temp_sp[24]), .B(n_26970), .Z(n_20439
		));
	notech_reg_set temp_sp_reg_25(.CP(n_62379), .D(n_20445), .SD(1'b1), .Q(temp_sp
		[25]));
	notech_mux2 i_6459(.S(n_53661), .A(temp_sp[25]), .B(n_26972), .Z(n_20445
		));
	notech_reg_set temp_sp_reg_26(.CP(n_62379), .D(n_20451), .SD(1'b1), .Q(temp_sp
		[26]));
	notech_mux2 i_6467(.S(n_53661), .A(temp_sp[26]), .B(n_26974), .Z(n_20451
		));
	notech_reg_set temp_sp_reg_27(.CP(n_62379), .D(n_20457), .SD(1'b1), .Q(temp_sp
		[27]));
	notech_mux2 i_6475(.S(n_53661), .A(temp_sp[27]), .B(n_26976), .Z(n_20457
		));
	notech_reg_set temp_sp_reg_28(.CP(n_62379), .D(n_20463), .SD(1'b1), .Q(temp_sp
		[28]));
	notech_mux2 i_6483(.S(n_53661), .A(temp_sp[28]), .B(n_26978), .Z(n_20463
		));
	notech_nand2 i_217133598(.A(n_56721), .B(n_56730), .Z(n_1880));
	notech_reg_set temp_sp_reg_29(.CP(n_62379), .D(n_20469), .SD(1'b1), .Q(temp_sp
		[29]));
	notech_mux2 i_6492(.S(n_53661), .A(temp_sp[29]), .B(n_26980), .Z(n_20469
		));
	notech_or4 i_217533594(.A(opa[14]), .B(opa[15]), .C(opa[12]), .D(opa[13]
		), .Z(n_1879));
	notech_reg_set temp_sp_reg_30(.CP(n_62379), .D(n_20475), .SD(1'b1), .Q(temp_sp
		[30]));
	notech_mux2 i_6501(.S(n_53661), .A(temp_sp[30]), .B(n_26984), .Z(n_20475
		));
	notech_reg_set temp_sp_reg_31(.CP(n_62379), .D(n_20481), .SD(1'b1), .Q(temp_sp
		[31]));
	notech_mux2 i_6509(.S(n_53661), .A(temp_sp[31]), .B(n_26986), .Z(n_20481
		));
	notech_reg regs_reg_4_0(.CP(n_62379), .D(n_20487), .CD(n_61199), .Q(regs_4
		[0]));
	notech_mux2 i_6517(.S(n_27000), .A(regs_4[0]), .B(n_12767), .Z(n_20487)
		);
	notech_reg regs_reg_4_1(.CP(n_62379), .D(n_20493), .CD(n_61199), .Q(regs_4
		[1]));
	notech_mux2 i_6525(.S(n_27000), .A(regs_4[1]), .B(n_26988), .Z(n_20493)
		);
	notech_reg regs_reg_4_2(.CP(n_62379), .D(n_20500), .CD(n_61200), .Q(regs_4
		[2]));
	notech_mux2 i_6533(.S(n_27000), .A(regs_4[2]), .B(n_26989), .Z(n_20500)
		);
	notech_ao4 i_217933590(.A(n_28981), .B(n_56246), .C(n_56235), .D(n_27722
		), .Z(n_1874));
	notech_reg regs_reg_4_3(.CP(n_62379), .D(n_20507), .CD(n_61202), .Q(regs_4
		[3]));
	notech_mux2 i_6541(.S(n_27000), .A(regs_4[3]), .B(n_26992), .Z(n_20507)
		);
	notech_ao4 i_218033589(.A(n_56255), .B(n_27793), .C(n_27825), .D(n_57358
		), .Z(n_1873));
	notech_reg regs_reg_4_4(.CP(n_62379), .D(n_20513), .CD(n_61202), .Q(regs_4
		[4]));
	notech_mux2 i_6549(.S(n_27000), .A(regs_4[4]), .B(n_26993), .Z(n_20513)
		);
	notech_and2 i_218433585(.A(n_1871), .B(n_1870), .Z(n_1872));
	notech_reg regs_reg_4_5(.CP(n_62379), .D(n_20519), .CD(n_61200), .Q(regs_4
		[5]));
	notech_mux2 i_6557(.S(n_27000), .A(regs_4[5]), .B(n_26996), .Z(n_20519)
		);
	notech_ao4 i_218233587(.A(n_56226), .B(n_27992), .C(n_56414), .D(n_27960
		), .Z(n_1871));
	notech_reg regs_reg_4_6(.CP(n_62379), .D(n_20525), .CD(n_61200), .Q(regs_4
		[6]));
	notech_mux2 i_6565(.S(n_27000), .A(regs_4[6]), .B(n_26997), .Z(n_20525)
		);
	notech_ao4 i_218333586(.A(n_56305), .B(n_27613), .C(n_27926), .D(n_56296
		), .Z(n_1870));
	notech_reg regs_reg_4_7(.CP(n_62379), .D(n_20531), .CD(n_61202), .Q(regs_4
		[7]));
	notech_mux2 i_6573(.S(n_27000), .A(regs_4[7]), .B(n_26998), .Z(n_20531)
		);
	notech_and4 i_219233577(.A(n_1867), .B(n_1866), .C(n_1864), .D(n_1863), 
		.Z(n_1869));
	notech_reg regs_reg_4_8(.CP(n_62379), .D(n_20537), .CD(n_61202), .Q(regs_4
		[8]));
	notech_mux2 i_6581(.S(n_27000), .A(regs_4[8]), .B(n_12815), .Z(n_20537)
		);
	notech_reg regs_reg_4_9(.CP(n_62391), .D(n_20543), .CD(n_61202), .Q(regs_4
		[9]));
	notech_mux2 i_6589(.S(n_27000), .A(regs_4[9]), .B(n_12821), .Z(n_20543)
		);
	notech_ao4 i_218633583(.A(n_56395), .B(n_28980), .C(n_60479), .D(n_27894
		), .Z(n_1867));
	notech_reg regs_reg_4_10(.CP(n_62391), .D(n_20549), .CD(n_61202), .Q(regs_4
		[10]));
	notech_mux2 i_6597(.S(n_27000), .A(regs_4[10]), .B(n_12827), .Z(n_20549)
		);
	notech_ao4 i_218733582(.A(n_56285), .B(n_27647), .C(n_56276), .D(n_27857
		), .Z(n_1866));
	notech_reg regs_reg_4_11(.CP(n_62391), .D(n_20555), .CD(n_61202), .Q(regs_4
		[11]));
	notech_mux2 i_6606(.S(n_27000), .A(regs_4[11]), .B(n_12833), .Z(n_20555)
		);
	notech_reg regs_reg_4_12(.CP(n_62391), .D(n_20561), .CD(n_61200), .Q(regs_4
		[12]));
	notech_mux2 i_6614(.S(n_27000), .A(regs_4[12]), .B(n_12839), .Z(n_20561)
		);
	notech_ao4 i_218933580(.A(n_56265), .B(n_27690), .C(n_57371), .D(n_27377
		), .Z(n_1864));
	notech_reg regs_reg_4_13(.CP(n_62391), .D(n_20568), .CD(n_61200), .Q(regs_4
		[13]));
	notech_mux2 i_6622(.S(n_27000), .A(regs_4[13]), .B(n_12845), .Z(n_20568)
		);
	notech_ao4 i_219033579(.A(n_57338), .B(n_27754), .C(n_28026), .D(n_59219
		), .Z(n_1863));
	notech_reg regs_reg_4_14(.CP(n_62391), .D(n_20575), .CD(n_61200), .Q(regs_4
		[14]));
	notech_mux2 i_6630(.S(n_27000), .A(regs_4[14]), .B(n_12851), .Z(n_20575)
		);
	notech_and2 i_35125(.A(n_57418), .B(n_327046818), .Z(n_1862));
	notech_reg regs_reg_4_15(.CP(n_62391), .D(n_20581), .CD(n_61200), .Q(regs_4
		[15]));
	notech_mux2 i_6638(.S(n_27000), .A(regs_4[15]), .B(n_12857), .Z(n_20581)
		);
	notech_reg regs_reg_4_16(.CP(n_62391), .D(n_20587), .CD(n_61200), .Q(regs_4
		[16]));
	notech_mux2 i_6646(.S(n_54101), .A(regs_4[16]), .B(n_12863), .Z(n_20587)
		);
	notech_reg regs_reg_4_17(.CP(n_62391), .D(n_20593), .CD(n_61200), .Q(regs_4
		[17]));
	notech_mux2 i_6654(.S(n_54101), .A(regs_4[17]), .B(n_12869), .Z(n_20593)
		);
	notech_reg regs_reg_4_18(.CP(n_62391), .D(n_20599), .CD(n_61200), .Q(regs_4
		[18]));
	notech_mux2 i_6662(.S(n_54101), .A(regs_4[18]), .B(n_12875), .Z(n_20599)
		);
	notech_reg regs_reg_4_19(.CP(n_62391), .D(n_20606), .CD(n_61200), .Q(regs_4
		[19]));
	notech_mux2 i_6670(.S(n_54101), .A(regs_4[19]), .B(n_12881), .Z(n_20606)
		);
	notech_reg regs_reg_4_20(.CP(n_62391), .D(n_20614), .CD(n_61200), .Q(regs_4
		[20]));
	notech_mux2 i_6678(.S(n_54101), .A(regs_4[20]), .B(n_12887), .Z(n_20614)
		);
	notech_reg regs_reg_4_21(.CP(n_62391), .D(n_20621), .CD(n_61198), .Q(regs_4
		[21]));
	notech_mux2 i_6686(.S(n_54101), .A(regs_4[21]), .B(n_12893), .Z(n_20621)
		);
	notech_reg regs_reg_4_22(.CP(n_62391), .D(n_20628), .CD(n_61194), .Q(regs_4
		[22]));
	notech_mux2 i_6694(.S(n_54101), .A(regs_4[22]), .B(n_12899), .Z(n_20628)
		);
	notech_reg regs_reg_4_23(.CP(n_62391), .D(n_20635), .CD(n_61194), .Q(regs_4
		[23]));
	notech_mux2 i_6702(.S(n_54101), .A(regs_4[23]), .B(n_12905), .Z(n_20635)
		);
	notech_reg regs_reg_4_24(.CP(n_62391), .D(n_20644), .CD(n_61194), .Q(regs_4
		[24]));
	notech_mux2 i_6710(.S(n_54101), .A(regs_4[24]), .B(n_12911), .Z(n_20644)
		);
	notech_reg regs_reg_4_25(.CP(n_62391), .D(n_20652), .CD(n_61194), .Q(regs_4
		[25]));
	notech_mux2 i_6718(.S(n_54101), .A(regs_4[25]), .B(n_12917), .Z(n_20652)
		);
	notech_reg regs_reg_4_26(.CP(n_62391), .D(n_20659), .CD(n_61194), .Q(regs_4
		[26]));
	notech_mux2 i_6726(.S(n_54101), .A(regs_4[26]), .B(n_12923), .Z(n_20659)
		);
	notech_reg regs_reg_4_27(.CP(n_62391), .D(n_20666), .CD(n_61197), .Q(regs_4
		[27]));
	notech_mux2 i_6734(.S(n_54101), .A(regs_4[27]), .B(n_12929), .Z(n_20666)
		);
	notech_reg regs_reg_4_28(.CP(n_62391), .D(n_20674), .CD(n_61197), .Q(regs_4
		[28]));
	notech_mux2 i_6742(.S(n_54101), .A(regs_4[28]), .B(n_12935), .Z(n_20674)
		);
	notech_reg regs_reg_4_29(.CP(n_62377), .D(n_20681), .CD(n_61194), .Q(regs_4
		[29]));
	notech_mux2 i_6750(.S(n_54101), .A(regs_4[29]), .B(n_12941), .Z(n_20681)
		);
	notech_reg regs_reg_4_30(.CP(n_62377), .D(n_20688), .CD(n_61194), .Q(regs_4
		[30]));
	notech_mux2 i_6758(.S(n_54101), .A(regs_4[30]), .B(n_12947), .Z(n_20688)
		);
	notech_reg regs_reg_4_31(.CP(n_62377), .D(n_20695), .CD(n_61193), .Q(regs_4
		[31]));
	notech_mux2 i_6766(.S(n_54101), .A(regs_4[31]), .B(n_12953), .Z(n_20695)
		);
	notech_or4 i_29703(.A(n_1879), .B(opa[8]), .C(opa[9]), .D(n_1880), .Z(n_1845
		));
	notech_reg regs_reg_3_0(.CP(n_62377), .D(n_20702), .CD(n_61194), .Q(regs_3
		[0]));
	notech_mux2 i_6774(.S(n_27022), .A(regs_3[0]), .B(n_27002), .Z(n_20702)
		);
	notech_or4 i_25735693(.A(n_2341), .B(n_2562), .C(n_2385), .D(n_59210), .Z
		(n_1844));
	notech_reg regs_reg_3_1(.CP(n_62377), .D(n_20710), .CD(n_61193), .Q(regs_3
		[1]));
	notech_mux2 i_6782(.S(n_27022), .A(regs_3[1]), .B(n_27004), .Z(n_20710)
		);
	notech_reg regs_reg_3_2(.CP(n_62377), .D(n_20717), .CD(n_61193), .Q(regs_3
		[2]));
	notech_mux2 i_6790(.S(n_27022), .A(regs_3[2]), .B(n_27005), .Z(n_20717)
		);
	notech_ao4 i_219936963(.A(n_261036765), .B(n_82713221), .C(n_260936764),
		 .D(n_82813222), .Z(n_1842));
	notech_reg regs_reg_3_3(.CP(n_62377), .D(n_20724), .CD(n_61194), .Q(regs_3
		[3]));
	notech_mux2 i_6798(.S(n_27022), .A(regs_3[3]), .B(n_12419), .Z(n_20724)
		);
	notech_and4 i_219836964(.A(n_1834), .B(n_1833), .C(n_1839), .D(n_1682), 
		.Z(n_1841));
	notech_reg regs_reg_3_4(.CP(n_62377), .D(n_20735), .CD(n_61194), .Q(regs_3
		[4]));
	notech_mux2 i_6806(.S(n_27022), .A(regs_3[4]), .B(n_27006), .Z(n_20735)
		);
	notech_reg regs_reg_3_5(.CP(n_62377), .D(n_20742), .CD(n_61194), .Q(regs_3
		[5]));
	notech_mux2 i_6814(.S(n_27022), .A(regs_3[5]), .B(n_12431), .Z(n_20742)
		);
	notech_and4 i_219636966(.A(n_54860), .B(n_1836), .C(n_167488959), .D(n_1681
		), .Z(n_1839));
	notech_reg regs_reg_3_6(.CP(n_62377), .D(n_20749), .CD(n_61194), .Q(regs_3
		[6]));
	notech_mux2 i_6822(.S(n_27022), .A(regs_3[6]), .B(n_27007), .Z(n_20749)
		);
	notech_reg regs_reg_3_7(.CP(n_62377), .D(n_20756), .CD(n_61194), .Q(regs_3
		[7]));
	notech_mux2 i_6830(.S(n_27022), .A(regs_3[7]), .B(n_27008), .Z(n_20756)
		);
	notech_reg regs_reg_3_8(.CP(n_62377), .D(n_20764), .CD(n_61197), .Q(regs_3
		[8]));
	notech_mux2 i_6838(.S(n_27022), .A(regs_3[8]), .B(n_27009), .Z(n_20764)
		);
	notech_ao4 i_219336969(.A(n_59150), .B(n_27533), .C(n_55739), .D(n_27579
		), .Z(n_1836));
	notech_reg regs_reg_3_9(.CP(n_62377), .D(n_20771), .CD(n_61198), .Q(regs_3
		[9]));
	notech_mux2 i_6846(.S(n_27022), .A(regs_3[9]), .B(n_12455), .Z(n_20771)
		);
	notech_reg regs_reg_3_10(.CP(n_62381), .D(n_20778), .CD(n_61198), .Q(regs_3
		[10]));
	notech_mux2 i_6854(.S(n_27022), .A(regs_3[10]), .B(n_27010), .Z(n_20778)
		);
	notech_ao4 i_219236970(.A(n_55318), .B(n_56757), .C(n_55317), .D(n_55566
		), .Z(n_1834));
	notech_reg regs_reg_3_11(.CP(n_62337), .D(n_20785), .CD(n_61197), .Q(regs_3
		[11]));
	notech_mux2 i_6862(.S(n_27022), .A(regs_3[11]), .B(n_12467), .Z(n_20785)
		);
	notech_ao4 i_219136971(.A(n_55431), .B(n_29006), .C(n_318588504), .D(n_29007
		), .Z(n_1833));
	notech_reg regs_reg_3_12(.CP(n_62337), .D(n_20792), .CD(n_61198), .Q(regs_3
		[12]));
	notech_mux2 i_6870(.S(n_27022), .A(regs_3[12]), .B(n_12473), .Z(n_20792)
		);
	notech_reg regs_reg_3_13(.CP(n_62337), .D(n_20798), .CD(n_61198), .Q(regs_3
		[13]));
	notech_mux2 i_6878(.S(n_27022), .A(regs_3[13]), .B(n_27011), .Z(n_20798)
		);
	notech_and4 i_167937477(.A(n_1828), .B(n_1671), .C(n_1791), .D(n_166888964
		), .Z(n_1831));
	notech_reg regs_reg_3_14(.CP(n_62337), .D(n_20804), .CD(n_61198), .Q(regs_3
		[14]));
	notech_mux2 i_6886(.S(n_27022), .A(regs_3[14]), .B(n_12485), .Z(n_20804)
		);
	notech_reg regs_reg_3_15(.CP(n_62337), .D(n_20811), .CD(n_61198), .Q(regs_3
		[15]));
	notech_mux2 i_6894(.S(n_27022), .A(regs_3[15]), .B(n_27012), .Z(n_20811)
		);
	notech_reg regs_reg_3_16(.CP(n_62337), .D(n_20818), .CD(n_61198), .Q(regs_3
		[16]));
	notech_mux2 i_6902(.S(n_54112), .A(regs_3[16]), .B(n_12497), .Z(n_20818)
		);
	notech_and4 i_167537481(.A(n_1793), .B(n_1792), .C(n_1820), .D(n_36812763
		), .Z(n_1828));
	notech_reg regs_reg_3_17(.CP(n_62337), .D(n_20824), .CD(n_61198), .Q(regs_3
		[17]));
	notech_mux2 i_6910(.S(n_54112), .A(regs_3[17]), .B(n_12503), .Z(n_20824)
		);
	notech_reg regs_reg_3_18(.CP(n_62337), .D(n_20830), .CD(n_61197), .Q(regs_3
		[18]));
	notech_mux2 i_6918(.S(n_54112), .A(regs_3[18]), .B(n_27013), .Z(n_20830)
		);
	notech_and4 i_167337483(.A(n_180756206), .B(n_180656205), .C(n_1796), .D
		(n_166788965), .Z(n_1820));
	notech_reg regs_reg_3_19(.CP(n_62337), .D(n_20836), .CD(n_61197), .Q(regs_3
		[19]));
	notech_mux2 i_6926(.S(n_54112), .A(regs_3[19]), .B(n_27014), .Z(n_20836)
		);
	notech_reg regs_reg_3_20(.CP(n_62337), .D(n_20842), .CD(n_61197), .Q(regs_3
		[20]));
	notech_mux2 i_6934(.S(n_54112), .A(regs_3[20]), .B(n_12521), .Z(n_20842)
		);
	notech_ao4 i_166737489(.A(n_55526), .B(n_28570), .C(n_55102), .D(n_28788
		), .Z(n_180756206));
	notech_reg regs_reg_3_21(.CP(n_62381), .D(n_20850), .CD(n_61197), .Q(regs_3
		[21]));
	notech_mux2 i_6942(.S(n_54112), .A(regs_3[21]), .B(n_27015), .Z(n_20850)
		);
	notech_ao4 i_166637490(.A(n_55181), .B(n_28973), .C(n_55161), .D(n_28815
		), .Z(n_180656205));
	notech_reg regs_reg_3_22(.CP(n_62381), .D(n_20857), .CD(n_61197), .Q(regs_3
		[22]));
	notech_mux2 i_6950(.S(n_54112), .A(regs_3[22]), .B(n_27016), .Z(n_20857)
		);
	notech_reg regs_reg_3_23(.CP(n_62381), .D(n_20864), .CD(n_61197), .Q(regs_3
		[23]));
	notech_mux2 i_6958(.S(n_54112), .A(regs_3[23]), .B(n_12539), .Z(n_20864)
		);
	notech_ao4 i_166537491(.A(n_55122), .B(n_55234), .C(n_55111), .D(nbus_11326
		[6]), .Z(n_1796));
	notech_reg regs_reg_3_24(.CP(n_62381), .D(n_20871), .CD(n_61197), .Q(regs_3
		[24]));
	notech_mux2 i_6966(.S(n_54112), .A(regs_3[24]), .B(n_27017), .Z(n_20871)
		);
	notech_reg regs_reg_3_25(.CP(n_62381), .D(n_20878), .CD(n_61197), .Q(regs_3
		[25]));
	notech_mux2 i_6975(.S(n_54112), .A(regs_3[25]), .B(n_12551), .Z(n_20878)
		);
	notech_ao4 i_166937487(.A(n_55136), .B(n_27579), .C(n_55170), .D(n_56757
		), .Z(n_1793));
	notech_reg regs_reg_3_26(.CP(n_62381), .D(n_20886), .CD(n_61197), .Q(regs_3
		[26]));
	notech_mux2 i_6983(.S(n_54112), .A(regs_3[26]), .B(n_27018), .Z(n_20886)
		);
	notech_ao4 i_166837488(.A(n_55192), .B(nbus_11326[14]), .C(n_55091), .D(n_28625
		), .Z(n_1792));
	notech_reg regs_reg_3_27(.CP(n_62381), .D(n_20896), .CD(n_61153), .Q(regs_3
		[27]));
	notech_mux2 i_6991(.S(n_54112), .A(regs_3[27]), .B(n_12563), .Z(n_20896)
		);
	notech_and2 i_4739045(.A(n_54725), .B(n_54719), .Z(n_36812763));
	notech_reg regs_reg_3_28(.CP(n_62381), .D(n_20904), .CD(n_61107), .Q(regs_3
		[28]));
	notech_mux2 i_6999(.S(n_54112), .A(regs_3[28]), .B(n_27020), .Z(n_20904)
		);
	notech_ao4 i_167737479(.A(n_89513289), .B(n_27599), .C(n_88913283), .D(n_28844
		), .Z(n_1791));
	notech_reg regs_reg_3_29(.CP(n_62381), .D(n_20911), .CD(n_61107), .Q(regs_3
		[29]));
	notech_mux2 i_7007(.S(n_54112), .A(regs_3[29]), .B(n_12575), .Z(n_20911)
		);
	notech_reg regs_reg_3_30(.CP(n_62381), .D(n_20918), .CD(n_61107), .Q(regs_3
		[30]));
	notech_mux2 i_7015(.S(n_54112), .A(regs_3[30]), .B(n_27021), .Z(n_20918)
		);
	notech_reg regs_reg_3_31(.CP(n_62381), .D(n_20925), .CD(n_61107), .Q(regs_3
		[31]));
	notech_mux2 i_7023(.S(n_54112), .A(regs_3[31]), .B(n_12587), .Z(n_20925)
		);
	notech_and4 i_128437867(.A(n_1784), .B(n_1783), .C(n_165288976), .D(n_1653
		), .Z(n_1788));
	notech_reg regs_reg_2_0(.CP(n_62381), .D(n_20932), .CD(n_61107), .Q(regs_2
		[0]));
	notech_mux2 i_7031(.S(n_27035), .A(regs_2[0]), .B(n_12049), .Z(n_20932)
		);
	notech_reg regs_reg_2_1(.CP(n_62381), .D(n_20940), .CD(n_61108), .Q(regs_2
		[1]));
	notech_mux2 i_7039(.S(n_27035), .A(regs_2[1]), .B(n_27023), .Z(n_20940)
		);
	notech_reg regs_reg_2_2(.CP(n_62381), .D(n_20947), .CD(n_61108), .Q(regs_2
		[2]));
	notech_mux2 i_7047(.S(n_27035), .A(regs_2[2]), .B(n_27024), .Z(n_20947)
		);
	notech_ao4 i_128037871(.A(n_55310), .B(n_55566), .C(n_55354), .D(n_29006
		), .Z(n_1784));
	notech_reg regs_reg_2_3(.CP(n_62381), .D(n_20954), .CD(n_61108), .Q(regs_2
		[3]));
	notech_mux2 i_7055(.S(n_27035), .A(regs_2[3]), .B(n_12067), .Z(n_20954)
		);
	notech_ao4 i_128137870(.A(n_55727), .B(n_27579), .C(n_56757), .D(n_26548
		), .Z(n_1783));
	notech_reg regs_reg_2_4(.CP(n_62381), .D(n_20961), .CD(n_61108), .Q(regs_2
		[4]));
	notech_mux2 i_7063(.S(n_27035), .A(regs_2[4]), .B(n_27025), .Z(n_20961)
		);
	notech_or2 i_63539082(.A(n_272188734), .B(n_55858), .Z(n_80913203));
	notech_reg regs_reg_2_5(.CP(n_62381), .D(n_20968), .CD(n_61107), .Q(regs_2
		[5]));
	notech_mux2 i_7072(.S(n_27035), .A(regs_2[5]), .B(n_12079), .Z(n_20968)
		);
	notech_nand2 i_5139087(.A(opc_10[14]), .B(n_62405), .Z(n_82713221));
	notech_reg regs_reg_2_6(.CP(n_62381), .D(n_20979), .CD(n_61107), .Q(regs_2
		[6]));
	notech_mux2 i_7080(.S(n_27035), .A(regs_2[6]), .B(n_12085), .Z(n_20979)
		);
	notech_nand2 i_1139088(.A(n_62427), .B(opc[14]), .Z(n_82813222));
	notech_reg regs_reg_2_7(.CP(n_62337), .D(n_20986), .CD(n_61104), .Q(regs_2
		[7]));
	notech_mux2 i_7088(.S(n_27035), .A(regs_2[7]), .B(n_27026), .Z(n_20986)
		);
	notech_reg regs_reg_2_8(.CP(n_62337), .D(n_20994), .CD(n_61104), .Q(regs_2
		[8]));
	notech_mux2 i_7096(.S(n_27035), .A(regs_2[8]), .B(n_27027), .Z(n_20994)
		);
	notech_reg regs_reg_2_9(.CP(n_62339), .D(n_21001), .CD(n_61107), .Q(regs_2
		[9]));
	notech_mux2 i_7104(.S(n_27035), .A(regs_2[9]), .B(n_27028), .Z(n_21001)
		);
	notech_ao4 i_80138315(.A(n_58487), .B(n_28033), .C(n_55952), .D(n_29000)
		, .Z(n_1780));
	notech_reg regs_reg_2_10(.CP(n_62339), .D(n_21008), .CD(n_61107), .Q(regs_2
		[10]));
	notech_mux2 i_7112(.S(n_27035), .A(regs_2[10]), .B(n_27029), .Z(n_21008)
		);
	notech_ao4 i_80038316(.A(n_55972), .B(n_27999), .C(n_55992), .D(n_27967)
		, .Z(n_1779));
	notech_reg regs_reg_2_11(.CP(n_62339), .D(n_21015), .CD(n_61107), .Q(regs_2
		[11]));
	notech_mux2 i_7120(.S(n_27035), .A(regs_2[11]), .B(n_12115), .Z(n_21015)
		);
	notech_and2 i_80638312(.A(n_177788904), .B(n_177688905), .Z(n_1778));
	notech_reg regs_reg_2_12(.CP(n_62339), .D(n_21022), .CD(n_61107), .Q(regs_2
		[12]));
	notech_mux2 i_7128(.S(n_27035), .A(regs_2[12]), .B(n_27030), .Z(n_21022)
		);
	notech_ao4 i_79938317(.A(n_56013), .B(n_27933), .C(n_56033), .D(n_27901)
		, .Z(n_177788904));
	notech_reg regs_reg_2_13(.CP(n_62339), .D(n_21030), .CD(n_61107), .Q(regs_2
		[13]));
	notech_mux2 i_7136(.S(n_27035), .A(regs_2[13]), .B(n_12127), .Z(n_21030)
		);
	notech_ao4 i_79838318(.A(n_56049), .B(n_27864), .C(n_55879), .D(n_27832)
		, .Z(n_177688905));
	notech_reg regs_reg_2_14(.CP(n_62339), .D(n_21036), .CD(n_61108), .Q(regs_2
		[14]));
	notech_mux2 i_7144(.S(n_27035), .A(regs_2[14]), .B(n_12133), .Z(n_21036)
		);
	notech_and4 i_80838310(.A(n_1773), .B(n_177288907), .C(n_177088909), .D(n_176988910
		), .Z(n_177588906));
	notech_reg regs_reg_2_15(.CP(n_62339), .D(n_21042), .CD(n_61109), .Q(regs_2
		[15]));
	notech_mux2 i_7152(.S(n_27035), .A(regs_2[15]), .B(n_12139), .Z(n_21042)
		);
	notech_reg regs_reg_2_16(.CP(n_62339), .D(n_21048), .CD(n_61109), .Q(regs_2
		[16]));
	notech_mux2 i_7160(.S(n_54137), .A(regs_2[16]), .B(n_12145), .Z(n_21048)
		);
	notech_ao4 i_79738319(.A(n_55934), .B(n_27800), .C(n_55893), .D(n_27763)
		, .Z(n_1773));
	notech_reg regs_reg_2_17(.CP(n_62339), .D(n_21057), .CD(n_61109), .Q(regs_2
		[17]));
	notech_mux2 i_7168(.S(n_54137), .A(regs_2[17]), .B(n_12151), .Z(n_21057)
		);
	notech_ao4 i_79638320(.A(n_55910), .B(n_27729), .C(n_55924), .D(n_27384)
		, .Z(n_177288907));
	notech_reg regs_reg_2_18(.CP(n_62339), .D(n_21063), .CD(n_61109), .Q(regs_2
		[18]));
	notech_mux2 i_7176(.S(n_54137), .A(regs_2[18]), .B(n_12157), .Z(n_21063)
		);
	notech_reg regs_reg_2_19(.CP(n_62339), .D(n_21069), .CD(n_61109), .Q(regs_2
		[19]));
	notech_mux2 i_7184(.S(n_54137), .A(regs_2[19]), .B(n_27031), .Z(n_21069)
		);
	notech_ao4 i_79538321(.A(n_56092), .B(n_27697), .C(n_56130), .D(n_27657)
		, .Z(n_177088909));
	notech_reg regs_reg_2_20(.CP(n_62339), .D(n_21075), .CD(n_61109), .Q(regs_2
		[20]));
	notech_mux2 i_7192(.S(n_54137), .A(regs_2[20]), .B(n_27032), .Z(n_21075)
		);
	notech_ao4 i_79438322(.A(n_56144), .B(n_27620), .C(n_56386), .D(n_29001)
		, .Z(n_176988910));
	notech_reg regs_reg_2_21(.CP(n_62339), .D(n_21081), .CD(n_61109), .Q(regs_2
		[21]));
	notech_mux2 i_7200(.S(n_54137), .A(regs_2[21]), .B(n_12175), .Z(n_21081)
		);
	notech_reg regs_reg_2_22(.CP(n_62339), .D(n_21087), .CD(n_61109), .Q(regs_2
		[22]));
	notech_mux2 i_7208(.S(n_54137), .A(regs_2[22]), .B(n_12181), .Z(n_21087)
		);
	notech_reg regs_reg_2_23(.CP(n_62339), .D(n_21093), .CD(n_61109), .Q(regs_2
		[23]));
	notech_mux2 i_7216(.S(n_54137), .A(regs_2[23]), .B(n_27033), .Z(n_21093)
		);
	notech_nand2 i_77238342(.A(n_176588914), .B(n_1628), .Z(n_176688913));
	notech_reg regs_reg_2_24(.CP(n_62339), .D(n_21099), .CD(n_61108), .Q(regs_2
		[24]));
	notech_mux2 i_7225(.S(n_54137), .A(regs_2[24]), .B(n_12193), .Z(n_21099)
		);
	notech_and4 i_77138343(.A(n_176388916), .B(n_176288917), .C(n_176088919)
		, .D(n_175988920), .Z(n_176588914));
	notech_reg regs_reg_2_25(.CP(n_62339), .D(n_21105), .CD(n_61108), .Q(regs_2
		[25]));
	notech_mux2 i_7233(.S(n_54137), .A(regs_2[25]), .B(n_12199), .Z(n_21105)
		);
	notech_reg regs_reg_2_26(.CP(n_62339), .D(n_21111), .CD(n_61108), .Q(regs_2
		[26]));
	notech_mux2 i_7241(.S(n_54137), .A(regs_2[26]), .B(n_12205), .Z(n_21111)
		);
	notech_ao4 i_76838346(.A(n_59183), .B(n_26781), .C(n_55842), .D(n_27582)
		, .Z(n_176388916));
	notech_reg regs_reg_2_27(.CP(n_62339), .D(n_21117), .CD(n_61108), .Q(regs_2
		[27]));
	notech_mux2 i_7249(.S(n_54137), .A(regs_2[27]), .B(n_27034), .Z(n_21117)
		);
	notech_ao4 i_76738347(.A(n_58922), .B(n_29005), .C(n_55492), .D(n_27535)
		, .Z(n_176288917));
	notech_reg regs_reg_2_28(.CP(n_62265), .D(n_21124), .CD(n_61108), .Q(regs_2
		[28]));
	notech_mux2 i_7257(.S(n_54137), .A(regs_2[28]), .B(n_12217), .Z(n_21124)
		);
	notech_reg regs_reg_2_29(.CP(n_62265), .D(n_21131), .CD(n_61109), .Q(regs_2
		[29]));
	notech_mux2 i_7265(.S(n_54137), .A(regs_2[29]), .B(n_12223), .Z(n_21131)
		);
	notech_ao4 i_76638348(.A(n_29004), .B(n_55597), .C(n_55568), .D(n_55590)
		, .Z(n_176088919));
	notech_reg regs_reg_2_30(.CP(n_62265), .D(n_21139), .CD(n_61109), .Q(regs_2
		[30]));
	notech_mux2 i_7273(.S(n_54137), .A(regs_2[30]), .B(n_12229), .Z(n_21139)
		);
	notech_ao4 i_76538349(.A(n_55567), .B(n_56775), .C(n_2212), .D(n_58987),
		 .Z(n_175988920));
	notech_reg regs_reg_2_31(.CP(n_62265), .D(n_21146), .CD(n_61108), .Q(regs_2
		[31]));
	notech_mux2 i_7281(.S(n_54137), .A(regs_2[31]), .B(n_12235), .Z(n_21146)
		);
	notech_reg_set cr0_reg_0(.CP(n_62265), .D(n_21154), .SD(n_61108), .Q(\nbus_14527[0] 
		));
	notech_mux2 i_7289(.S(n_301386333), .A(opa[0]), .B(n_60130), .Z(n_21154)
		);
	notech_reg cr0_reg_1(.CP(n_62265), .D(n_21161), .CD(n_61104), .Q(\nbus_14523[1] 
		));
	notech_mux2 i_7297(.S(n_301386333), .A(opa[1]), .B(\nbus_14523[1] ), .Z(n_21161
		));
	notech_reg cr0_reg_2(.CP(n_62265), .D(n_21169), .CD(n_61102), .Q(cr0[2])
		);
	notech_mux2 i_7305(.S(n_301386333), .A(opa[2]), .B(cr0[2]), .Z(n_21169)
		);
	notech_ao4 i_74638368(.A(n_55934), .B(n_27802), .C(n_55924), .D(n_27386)
		, .Z(n_175688923));
	notech_reg cr0_reg_3(.CP(n_62265), .D(n_21176), .CD(n_61102), .Q(\nbus_14523[3] 
		));
	notech_mux2 i_7313(.S(n_301386333), .A(opa[3]), .B(\nbus_14523[3] ), .Z(n_21176
		));
	notech_ao4 i_74538369(.A(n_58487), .B(n_28035), .C(n_56092), .D(n_27699)
		, .Z(n_175588924));
	notech_reg cr0_reg_4(.CP(n_62265), .D(n_21184), .CD(n_61102), .Q(\nbus_14523[4] 
		));
	notech_mux2 i_7321(.S(n_301386333), .A(opa[4]), .B(\nbus_14523[4] ), .Z(n_21184
		));
	notech_and2 i_74938365(.A(n_1753), .B(n_1752), .Z(n_1754));
	notech_reg cr0_reg_5(.CP(n_62265), .D(n_21191), .CD(n_61102), .Q(\nbus_14523[5] 
		));
	notech_mux2 i_7329(.S(n_301386333), .A(opa[5]), .B(\nbus_14523[5] ), .Z(n_21191
		));
	notech_ao4 i_74438370(.A(n_56049), .B(n_27867), .C(n_56130), .D(n_27659)
		, .Z(n_1753));
	notech_reg cr0_reg_6(.CP(n_62265), .D(n_21199), .CD(n_61102), .Q(\nbus_14523[6] 
		));
	notech_mux2 i_7337(.S(n_301386333), .A(opa[6]), .B(\nbus_14523[6] ), .Z(n_21199
		));
	notech_ao4 i_74338371(.A(n_56033), .B(n_27903), .C(n_56386), .D(n_29003)
		, .Z(n_1752));
	notech_reg cr0_reg_7(.CP(n_62265), .D(n_21206), .CD(n_61103), .Q(\nbus_14523[7] 
		));
	notech_mux2 i_7345(.S(n_301386333), .A(opa[7]), .B(\nbus_14523[7] ), .Z(n_21206
		));
	notech_and4 i_75138363(.A(n_1749), .B(n_1748), .C(n_1746), .D(n_1745), .Z
		(n_1751));
	notech_reg cr0_reg_8(.CP(n_62347), .D(n_21214), .CD(n_61103), .Q(\nbus_14523[8] 
		));
	notech_mux2 i_7353(.S(n_301386333), .A(opa[8]), .B(\nbus_14523[8] ), .Z(n_21214
		));
	notech_reg cr0_reg_9(.CP(n_62197), .D(n_21221), .CD(n_61102), .Q(\nbus_14523[9] 
		));
	notech_mux2 i_7361(.S(n_301386333), .A(opa[9]), .B(\nbus_14523[9] ), .Z(n_21221
		));
	notech_ao4 i_74238372(.A(n_56013), .B(n_27935), .C(n_56144), .D(n_27622)
		, .Z(n_1749));
	notech_reg cr0_reg_10(.CP(n_62197), .D(n_21229), .CD(n_61102), .Q(\nbus_14523[10] 
		));
	notech_mux2 i_7369(.S(n_301386333), .A(opa[10]), .B(\nbus_14523[10] ), .Z
		(n_21229));
	notech_ao4 i_74138373(.A(n_55992), .B(n_27969), .C(n_55893), .D(n_27766)
		, .Z(n_1748));
	notech_reg cr0_reg_11(.CP(n_62197), .D(n_21236), .CD(n_61101), .Q(\nbus_14523[11] 
		));
	notech_mux2 i_7377(.S(n_301386333), .A(opa[11]), .B(\nbus_14523[11] ), .Z
		(n_21236));
	notech_reg cr0_reg_12(.CP(n_62197), .D(n_21244), .CD(n_61101), .Q(\nbus_14523[12] 
		));
	notech_mux2 i_7385(.S(n_301386333), .A(opa[12]), .B(\nbus_14523[12] ), .Z
		(n_21244));
	notech_ao4 i_74038374(.A(n_55972), .B(n_28001), .C(n_55879), .D(n_27834)
		, .Z(n_1746));
	notech_reg cr0_reg_13(.CP(n_62197), .D(n_21251), .CD(n_61101), .Q(\nbus_14523[13] 
		));
	notech_mux2 i_7393(.S(n_301386333), .A(opa[13]), .B(\nbus_14523[13] ), .Z
		(n_21251));
	notech_ao4 i_73938375(.A(n_55910), .B(n_27731), .C(n_55952), .D(n_29002)
		, .Z(n_1745));
	notech_reg cr0_reg_14(.CP(n_62197), .D(n_21259), .CD(n_61101), .Q(\nbus_14523[14] 
		));
	notech_mux2 i_7401(.S(n_301386333), .A(opa[14]), .B(\nbus_14523[14] ), .Z
		(n_21259));
	notech_reg cr0_reg_15(.CP(n_62197), .D(n_21266), .CD(n_61102), .Q(\nbus_14523[15] 
		));
	notech_mux2 i_7409(.S(n_301386333), .A(opa[15]), .B(\nbus_14523[15] ), .Z
		(n_21266));
	notech_reg cr0_reg_16(.CP(n_62197), .D(n_21274), .CD(n_61102), .Q(cr0[16
		]));
	notech_mux2 i_7417(.S(n_60452), .A(opa[16]), .B(cr0[16]), .Z(n_21274));
	notech_ao4 i_71438400(.A(n_98113375), .B(n_56784), .C(n_101413408), .D(n_28987
		), .Z(n_174288925));
	notech_reg cr0_reg_17(.CP(n_62197), .D(n_21281), .CD(n_61102), .Q(\nbus_14523[17] 
		));
	notech_mux2 i_7425(.S(n_60452), .A(opa[17]), .B(\nbus_14523[17] ), .Z(n_21281
		));
	notech_reg cr0_reg_18(.CP(n_62197), .D(n_21287), .CD(n_61102), .Q(\nbus_14523[18] 
		));
	notech_mux2 i_7433(.S(n_60452), .A(opa[18]), .B(\nbus_14523[18] ), .Z(n_21287
		));
	notech_reg cr0_reg_19(.CP(n_62277), .D(n_21293), .CD(n_61102), .Q(\nbus_14523[19] 
		));
	notech_mux2 i_7442(.S(n_60452), .A(opa[19]), .B(\nbus_14523[19] ), .Z(n_21293
		));
	notech_ao4 i_69538419(.A(n_56255), .B(n_27803), .C(n_57371), .D(n_27387)
		, .Z(n_1739));
	notech_reg cr0_reg_20(.CP(n_62277), .D(n_21299), .CD(n_61103), .Q(\nbus_14523[20] 
		));
	notech_mux2 i_7450(.S(n_60452), .A(opa[20]), .B(\nbus_14523[20] ), .Z(n_21299
		));
	notech_ao4 i_69438420(.A(n_59219), .B(n_28036), .C(n_56265), .D(n_27700)
		, .Z(n_1738));
	notech_reg cr0_reg_21(.CP(n_62277), .D(n_21305), .CD(n_61104), .Q(\nbus_14523[21] 
		));
	notech_mux2 i_7458(.S(n_60452), .A(opa[21]), .B(\nbus_14523[21] ), .Z(n_21305
		));
	notech_and2 i_69838416(.A(n_1736), .B(n_1735), .Z(n_1737));
	notech_reg cr0_reg_22(.CP(n_62277), .D(n_21312), .CD(n_61104), .Q(\nbus_14523[22] 
		));
	notech_mux2 i_7466(.S(n_60452), .A(opa[22]), .B(\nbus_14523[22] ), .Z(n_21312
		));
	notech_ao4 i_69338421(.A(n_56276), .B(n_27868), .C(n_56285), .D(n_27660)
		, .Z(n_1736));
	notech_reg cr0_reg_23(.CP(n_62277), .D(n_21319), .CD(n_61104), .Q(\nbus_14523[23] 
		));
	notech_mux2 i_7474(.S(n_60452), .A(opa[23]), .B(\nbus_14523[23] ), .Z(n_21319
		));
	notech_ao4 i_69238422(.A(n_60479), .B(n_27904), .C(n_56395), .D(n_28978)
		, .Z(n_1735));
	notech_reg cr0_reg_24(.CP(n_62277), .D(n_21326), .CD(n_61104), .Q(\nbus_14523[24] 
		));
	notech_mux2 i_7482(.S(n_60452), .A(opa[24]), .B(\nbus_14523[24] ), .Z(n_21326
		));
	notech_and4 i_70038414(.A(n_1732), .B(n_1731), .C(n_1729), .D(n_1728), .Z
		(n_1734));
	notech_reg cr0_reg_25(.CP(n_62277), .D(n_21334), .CD(n_61104), .Q(\nbus_14523[25] 
		));
	notech_mux2 i_7490(.S(n_60452), .A(opa[25]), .B(\nbus_14523[25] ), .Z(n_21334
		));
	notech_reg cr0_reg_26(.CP(n_62277), .D(n_21341), .CD(n_61104), .Q(\nbus_14523[26] 
		));
	notech_mux2 i_7498(.S(n_60452), .A(opa[26]), .B(\nbus_14523[26] ), .Z(n_21341
		));
	notech_ao4 i_69138423(.A(n_56296), .B(n_27937), .C(n_56305), .D(n_27623)
		, .Z(n_1732));
	notech_reg cr0_reg_27(.CP(n_62277), .D(n_21348), .CD(n_61104), .Q(\nbus_14523[27] 
		));
	notech_mux2 i_7506(.S(n_60452), .A(opa[27]), .B(\nbus_14523[27] ), .Z(n_21348
		));
	notech_ao4 i_69038424(.A(n_56409), .B(n_27970), .C(n_57338), .D(n_27768)
		, .Z(n_1731));
	notech_reg cr0_reg_28(.CP(n_62277), .D(n_21355), .CD(n_61104), .Q(\nbus_14523[28] 
		));
	notech_mux2 i_7514(.S(n_60452), .A(opa[28]), .B(\nbus_14523[28] ), .Z(n_21355
		));
	notech_reg cr0_reg_29(.CP(n_62277), .D(n_21362), .CD(n_61104), .Q(\nbus_14523[29] 
		));
	notech_mux2 i_7522(.S(n_60452), .A(opa[29]), .B(\nbus_14523[29] ), .Z(n_21362
		));
	notech_ao4 i_68938425(.A(n_56226), .B(n_28002), .C(n_27835), .D(n_57358)
		, .Z(n_1729));
	notech_reg cr0_reg_30(.CP(n_62277), .D(n_21370), .CD(n_61103), .Q(\nbus_14523[30] 
		));
	notech_mux2 i_7530(.S(n_60452), .A(opa[30]), .B(\nbus_14523[30] ), .Z(n_21370
		));
	notech_ao4 i_68838426(.A(n_56235), .B(n_27732), .C(n_56246), .D(n_28979)
		, .Z(n_1728));
	notech_reg cr0_reg_31(.CP(n_62277), .D(n_21377), .CD(n_61103), .Q(\nbus_14523[31] 
		));
	notech_mux2 i_7541(.S(n_60452), .A(opa[31]), .B(\nbus_14523[31] ), .Z(n_21377
		));
	notech_reg mask8b_reg_0(.CP(n_62277), .D(n_21384), .CD(n_61103), .Q(mask8b
		[0]));
	notech_mux2 i_7549(.S(\nbus_11302[0] ), .A(mask8b[0]), .B(n_27062), .Z(n_21384
		));
	notech_reg mask8b_reg_1(.CP(n_62277), .D(n_21391), .CD(n_61103), .Q(mask8b
		[1]));
	notech_mux2 i_7557(.S(\nbus_11302[0] ), .A(mask8b[1]), .B(n_27063), .Z(n_21391
		));
	notech_ao4 i_28138813(.A(n_56255), .B(n_27786), .C(n_57371), .D(n_27370)
		, .Z(n_1725));
	notech_reg mask8b_reg_2(.CP(n_62277), .D(n_21398), .CD(n_61103), .Q(mask8b
		[2]));
	notech_mux2 i_7565(.S(\nbus_11302[0] ), .A(mask8b[2]), .B(n_11427), .Z(n_21398
		));
	notech_ao4 i_28038814(.A(n_59224), .B(n_28019), .C(n_56265), .D(n_27681)
		, .Z(n_1724));
	notech_reg opb_reg_0(.CP(n_62277), .D(n_21405), .CD(n_61103), .Q(opb[0])
		);
	notech_mux2 i_7573(.S(n_27069), .A(opb[0]), .B(n_27065), .Z(n_21405));
	notech_and2 i_28438810(.A(n_1722), .B(n_172188926), .Z(n_1723));
	notech_reg opb_reg_1(.CP(n_62277), .D(n_21411), .CD(n_61103), .Q(opb[1])
		);
	notech_mux2 i_7581(.S(n_27069), .A(opb[1]), .B(n_14098), .Z(n_21411));
	notech_ao4 i_27938815(.A(n_56276), .B(n_27850), .C(n_56290), .D(n_27639)
		, .Z(n_1722));
	notech_reg opb_reg_2(.CP(n_62277), .D(n_21417), .CD(n_61103), .Q(opb[2])
		);
	notech_mux2 i_7589(.S(n_27069), .A(opb[2]), .B(n_27066), .Z(n_21417));
	notech_ao4 i_27838816(.A(n_60479), .B(n_27885), .C(n_56395), .D(n_27559)
		, .Z(n_172188926));
	notech_reg opb_reg_3(.CP(n_62275), .D(n_21423), .CD(n_61103), .Q(opb[3])
		);
	notech_mux2 i_7597(.S(n_27069), .A(opb[3]), .B(n_27067), .Z(n_21423));
	notech_and4 i_28638808(.A(n_1718), .B(n_1717), .C(n_1715), .D(n_1714), .Z
		(n_1720));
	notech_reg opb_reg_4(.CP(n_62275), .D(n_21429), .CD(n_61109), .Q(opb[4])
		);
	notech_mux2 i_7605(.S(n_27069), .A(opb[4]), .B(n_14116), .Z(n_21429));
	notech_reg opb_reg_5(.CP(n_62351), .D(n_21435), .CD(n_61115), .Q(opb[5])
		);
	notech_mux2 i_7613(.S(n_27069), .A(opb[5]), .B(n_14122), .Z(n_21435));
	notech_ao4 i_27738817(.A(n_56296), .B(n_27919), .C(n_56310), .D(n_27602)
		, .Z(n_1718));
	notech_reg opb_reg_6(.CP(n_62351), .D(n_21441), .CD(n_61115), .Q(opb[6])
		);
	notech_mux2 i_7621(.S(n_27069), .A(opb[6]), .B(n_14128), .Z(n_21441));
	notech_ao4 i_27638818(.A(n_56409), .B(n_27953), .C(n_57343), .D(n_27747)
		, .Z(n_1717));
	notech_reg opb_reg_7(.CP(n_62351), .D(n_21447), .CD(n_61114), .Q(opb[7])
		);
	notech_mux2 i_7629(.S(n_27069), .A(opb[7]), .B(n_14134), .Z(n_21447));
	notech_reg opb_reg_8(.CP(n_62351), .D(n_21453), .CD(n_61115), .Q(opb[8])
		);
	notech_mux2 i_7637(.S(n_27069), .A(opb[8]), .B(n_14140), .Z(n_21453));
	notech_ao4 i_27538819(.A(n_56226), .B(n_27985), .C(n_27818), .D(n_57358)
		, .Z(n_1715));
	notech_reg opb_reg_9(.CP(n_62351), .D(n_21459), .CD(n_61115), .Q(opb[9])
		);
	notech_mux2 i_7645(.S(n_27069), .A(opb[9]), .B(n_27068), .Z(n_21459));
	notech_ao4 i_27438820(.A(n_56240), .B(n_27715), .C(n_56246), .D(n_28985)
		, .Z(n_1714));
	notech_reg opb_reg_10(.CP(n_62351), .D(n_21465), .CD(n_61115), .Q(opb[10
		]));
	notech_mux2 i_7653(.S(n_27069), .A(opb[10]), .B(n_14152), .Z(n_21465));
	notech_nand2 i_169749210(.A(n_56538), .B(n_205888855), .Z(n_54761));
	notech_reg opb_reg_11(.CP(n_62351), .D(n_21471), .CD(n_61115), .Q(opb[11
		]));
	notech_mux2 i_7661(.S(n_27069), .A(opb[11]), .B(n_14158), .Z(n_21471));
	notech_nao3 i_104449228(.A(n_26599), .B(n_56551), .C(n_205788856), .Z(n_55325
		));
	notech_reg opb_reg_12(.CP(n_62351), .D(n_21477), .CD(n_61115), .Q(opb[12
		]));
	notech_mux2 i_7669(.S(n_27069), .A(opb[12]), .B(n_14164), .Z(n_21477));
	notech_reg opb_reg_13(.CP(n_62351), .D(n_21483), .CD(n_61115), .Q(opb[13
		]));
	notech_mux2 i_7677(.S(n_27069), .A(opb[13]), .B(n_14170), .Z(n_21483));
	notech_reg opb_reg_14(.CP(n_62351), .D(n_21489), .CD(n_61114), .Q(opb[14
		]));
	notech_mux2 i_7685(.S(n_27069), .A(opb[14]), .B(n_14176), .Z(n_21489));
	notech_reg opb_reg_15(.CP(n_62351), .D(n_21495), .CD(n_61114), .Q(opb[15
		]));
	notech_mux2 i_7693(.S(n_27069), .A(opb[15]), .B(n_14182), .Z(n_21495));
	notech_ao4 i_15738936(.A(n_2262), .B(n_27802), .C(n_57367), .D(n_27386),
		 .Z(n_171088929));
	notech_reg opb_reg_16(.CP(n_62351), .D(n_21501), .CD(n_61114), .Q(opb[16
		]));
	notech_mux2 i_7701(.S(\nbus_11314[16] ), .A(opb[16]), .B(n_27070), .Z(n_21501
		));
	notech_ao4 i_15638937(.A(n_59219), .B(n_28035), .C(n_56265), .D(n_27699)
		, .Z(n_170988930));
	notech_reg opb_reg_17(.CP(n_62351), .D(n_21507), .CD(n_61114), .Q(opb[17
		]));
	notech_mux2 i_7709(.S(\nbus_11314[16] ), .A(opb[17]), .B(n_27071), .Z(n_21507
		));
	notech_and2 i_16038933(.A(n_170788932), .B(n_170688933), .Z(n_170888931)
		);
	notech_reg opb_reg_18(.CP(n_62351), .D(n_21513), .CD(n_61114), .Q(opb[18
		]));
	notech_mux2 i_7717(.S(\nbus_11314[16] ), .A(opb[18]), .B(n_14200), .Z(n_21513
		));
	notech_ao4 i_15538938(.A(n_56276), .B(n_27867), .C(n_56285), .D(n_27659)
		, .Z(n_170788932));
	notech_reg opb_reg_19(.CP(n_62351), .D(n_21519), .CD(n_61114), .Q(opb[19
		]));
	notech_mux2 i_7726(.S(\nbus_11314[16] ), .A(opb[19]), .B(n_14206), .Z(n_21519
		));
	notech_ao4 i_15438939(.A(n_60479), .B(n_27903), .C(n_56395), .D(n_29003)
		, .Z(n_170688933));
	notech_reg opb_reg_20(.CP(n_62351), .D(n_21525), .CD(n_61114), .Q(opb[20
		]));
	notech_mux2 i_7734(.S(\nbus_11314[16] ), .A(opb[20]), .B(n_14212), .Z(n_21525
		));
	notech_and4 i_16238931(.A(n_170388936), .B(n_170288937), .C(n_170088939)
		, .D(n_169988940), .Z(n_170588934));
	notech_reg opb_reg_21(.CP(n_62351), .D(n_21531), .CD(n_61114), .Q(opb[21
		]));
	notech_mux2 i_7742(.S(\nbus_11314[16] ), .A(opb[21]), .B(n_14218), .Z(n_21531
		));
	notech_reg opb_reg_22(.CP(n_62351), .D(n_21537), .CD(n_61114), .Q(opb[22
		]));
	notech_mux2 i_7750(.S(\nbus_11314[16] ), .A(opb[22]), .B(n_14224), .Z(n_21537
		));
	notech_ao4 i_15338940(.A(n_27935), .B(n_56296), .C(n_56305), .D(n_27622)
		, .Z(n_170388936));
	notech_reg opb_reg_23(.CP(n_62275), .D(n_21543), .CD(n_61115), .Q(opb[23
		]));
	notech_mux2 i_7758(.S(\nbus_11314[16] ), .A(opb[23]), .B(n_14230), .Z(n_21543
		));
	notech_ao4 i_15238941(.A(n_56409), .B(n_27969), .C(n_57338), .D(n_27766)
		, .Z(n_170288937));
	notech_reg opb_reg_24(.CP(n_62275), .D(n_21549), .CD(n_61118), .Q(opb[24
		]));
	notech_mux2 i_7766(.S(\nbus_11314[16] ), .A(opb[24]), .B(n_14236), .Z(n_21549
		));
	notech_reg opb_reg_25(.CP(n_62275), .D(n_21555), .CD(n_61118), .Q(opb[25
		]));
	notech_mux2 i_7774(.S(\nbus_11314[16] ), .A(opb[25]), .B(n_14242), .Z(n_21555
		));
	notech_ao4 i_15138942(.A(n_28001), .B(n_56226), .C(n_27834), .D(n_57358)
		, .Z(n_170088939));
	notech_reg opb_reg_26(.CP(n_62275), .D(n_21561), .CD(n_61118), .Q(opb[26
		]));
	notech_mux2 i_7782(.S(\nbus_11314[16] ), .A(opb[26]), .B(n_14248), .Z(n_21561
		));
	notech_ao4 i_15038943(.A(n_56235), .B(n_27731), .C(n_29002), .D(n_56246)
		, .Z(n_169988940));
	notech_reg opb_reg_27(.CP(n_62275), .D(n_21567), .CD(n_61118), .Q(opb[27
		]));
	notech_mux2 i_7790(.S(\nbus_11314[16] ), .A(opb[27]), .B(n_14254), .Z(n_21567
		));
	notech_reg opb_reg_28(.CP(n_62275), .D(n_21573), .CD(n_61118), .Q(opb[28
		]));
	notech_mux2 i_7798(.S(\nbus_11314[16] ), .A(opb[28]), .B(n_14260), .Z(n_21573
		));
	notech_reg opb_reg_29(.CP(n_62275), .D(n_21579), .CD(n_61119), .Q(opb[29
		]));
	notech_mux2 i_7806(.S(\nbus_11314[16] ), .A(opb[29]), .B(n_14266), .Z(n_21579
		));
	notech_ao4 i_12038973(.A(n_56255), .B(n_27800), .C(n_57367), .D(n_27384)
		, .Z(n_169688943));
	notech_reg opb_reg_30(.CP(n_62275), .D(n_21585), .CD(n_61119), .Q(opb[30
		]));
	notech_mux2 i_7814(.S(\nbus_11314[16] ), .A(opb[30]), .B(n_27072), .Z(n_21585
		));
	notech_ao4 i_11938974(.A(n_59219), .B(n_28033), .C(n_56265), .D(n_27697)
		, .Z(n_169588944));
	notech_reg opb_reg_31(.CP(n_62275), .D(n_21591), .CD(n_61118), .Q(opb[31
		]));
	notech_mux2 i_7822(.S(\nbus_11314[16] ), .A(opb[31]), .B(n_27073), .Z(n_21591
		));
	notech_and2 i_12338970(.A(n_169388946), .B(n_169288947), .Z(n_169488945)
		);
	notech_reg_set divq_reg_0(.CP(n_62275), .D(n_21597), .SD(1'b1), .Q(divq[
		0]));
	notech_mux2 i_7830(.S(n_54358), .A(divq[0]), .B(n_8312), .Z(n_21597));
	notech_ao4 i_11838975(.A(n_56276), .B(n_27864), .C(n_56285), .D(n_27657)
		, .Z(n_169388946));
	notech_reg_set divq_reg_1(.CP(n_62351), .D(n_21603), .SD(1'b1), .Q(divq[
		1]));
	notech_mux2 i_7838(.S(n_54358), .A(divq[1]), .B(n_8317), .Z(n_21603));
	notech_ao4 i_11738976(.A(n_60479), .B(n_27901), .C(n_56395), .D(n_29001)
		, .Z(n_169288947));
	notech_reg_set divq_reg_2(.CP(n_62197), .D(n_21609), .SD(1'b1), .Q(divq[
		2]));
	notech_mux2 i_7846(.S(n_54358), .A(divq[2]), .B(n_8322), .Z(n_21609));
	notech_and4 i_12538968(.A(n_168988950), .B(n_168888951), .C(n_168688953)
		, .D(n_168588954), .Z(n_169188948));
	notech_reg_set divq_reg_3(.CP(n_62273), .D(n_21615), .SD(1'b1), .Q(divq[
		3]));
	notech_mux2 i_7854(.S(n_54358), .A(divq[3]), .B(n_8327), .Z(n_21615));
	notech_reg_set divq_reg_4(.CP(n_62347), .D(n_21621), .SD(1'b1), .Q(divq[
		4]));
	notech_mux2 i_7862(.S(n_54358), .A(divq[4]), .B(n_8332), .Z(n_21621));
	notech_ao4 i_11638977(.A(n_56296), .B(n_27933), .C(n_56305), .D(n_27620)
		, .Z(n_168988950));
	notech_reg_set divq_reg_5(.CP(n_62347), .D(n_21627), .SD(1'b1), .Q(divq[
		5]));
	notech_mux2 i_7870(.S(n_54358), .A(divq[5]), .B(n_8337), .Z(n_21627));
	notech_ao4 i_11538978(.A(n_56409), .B(n_27967), .C(n_57338), .D(n_27763)
		, .Z(n_168888951));
	notech_reg_set divq_reg_6(.CP(n_62347), .D(n_21633), .SD(1'b1), .Q(divq[
		6]));
	notech_mux2 i_7878(.S(n_54358), .A(divq[6]), .B(n_8342), .Z(n_21633));
	notech_reg_set divq_reg_7(.CP(n_62347), .D(n_21639), .SD(1'b1), .Q(divq[
		7]));
	notech_mux2 i_7886(.S(n_54358), .A(divq[7]), .B(n_8347), .Z(n_21639));
	notech_ao4 i_11438979(.A(n_56226), .B(n_27999), .C(n_27832), .D(n_57358)
		, .Z(n_168688953));
	notech_reg_set divq_reg_8(.CP(n_62347), .D(n_21645), .SD(1'b1), .Q(divq[
		8]));
	notech_mux2 i_7894(.S(n_54358), .A(divq[8]), .B(n_8352), .Z(n_21645));
	notech_ao4 i_11338980(.A(n_56235), .B(n_27729), .C(n_29000), .D(n_56246)
		, .Z(n_168588954));
	notech_reg_set divq_reg_9(.CP(n_62347), .D(n_21651), .SD(1'b1), .Q(divq[
		9]));
	notech_mux2 i_7902(.S(n_54358), .A(divq[9]), .B(n_8357), .Z(n_21651));
	notech_nand3 i_1516664(.A(n_1842), .B(n_1841), .C(n_167388960), .Z(n_11776
		));
	notech_reg_set divq_reg_10(.CP(n_62347), .D(n_21657), .SD(1'b1), .Q(divq
		[10]));
	notech_mux2 i_7910(.S(n_54358), .A(divq[10]), .B(n_8362), .Z(n_21657));
	notech_reg_set divq_reg_11(.CP(n_62347), .D(n_21663), .SD(1'b1), .Q(divq
		[11]));
	notech_mux2 i_7918(.S(n_54358), .A(divq[11]), .B(n_8367), .Z(n_21663));
	notech_reg_set divq_reg_12(.CP(n_62347), .D(n_21669), .SD(1'b1), .Q(divq
		[12]));
	notech_mux2 i_7926(.S(n_54358), .A(divq[12]), .B(n_8372), .Z(n_21669));
	notech_or4 i_218736975(.A(n_58656), .B(n_59277), .C(n_56345), .D(n_272188734
		), .Z(n_1682));
	notech_reg_set divq_reg_13(.CP(n_62347), .D(n_21675), .SD(1'b1), .Q(divq
		[13]));
	notech_mux2 i_7934(.S(n_54358), .A(divq[13]), .B(n_8377), .Z(n_21675));
	notech_nand2 i_218536977(.A(sav_ecx[14]), .B(n_60584), .Z(n_1681));
	notech_reg_set divq_reg_14(.CP(n_62347), .D(n_21681), .SD(1'b1), .Q(divq
		[14]));
	notech_mux2 i_7942(.S(n_54358), .A(divq[14]), .B(n_8382), .Z(n_21681));
	notech_reg_set divq_reg_15(.CP(n_62385), .D(n_21687), .SD(1'b1), .Q(divq
		[15]));
	notech_mux2 i_7950(.S(n_54358), .A(divq[15]), .B(n_8387), .Z(n_21687));
	notech_reg_set divq_reg_16(.CP(n_62385), .D(n_21693), .SD(1'b1), .Q(divq
		[16]));
	notech_mux2 i_7958(.S(n_54360), .A(divq[16]), .B(n_8392), .Z(n_21693));
	notech_reg_set divq_reg_17(.CP(n_62385), .D(n_21699), .SD(1'b1), .Q(divq
		[17]));
	notech_mux2 i_7966(.S(n_54360), .A(divq[17]), .B(n_8397), .Z(n_21699));
	notech_reg_set divq_reg_18(.CP(n_62385), .D(n_21705), .SD(1'b1), .Q(divq
		[18]));
	notech_mux2 i_7974(.S(n_54360), .A(divq[18]), .B(n_8402), .Z(n_21705));
	notech_reg_set divq_reg_19(.CP(n_62385), .D(n_21711), .SD(1'b1), .Q(divq
		[19]));
	notech_mux2 i_7982(.S(n_54360), .A(divq[19]), .B(n_8407), .Z(n_21711));
	notech_reg_set divq_reg_20(.CP(n_62385), .D(n_21717), .SD(1'b1), .Q(divq
		[20]));
	notech_mux2 i_7990(.S(n_54360), .A(divq[20]), .B(n_8412), .Z(n_21717));
	notech_nao3 i_217836984(.A(\regs_1[14] ), .B(n_28140), .C(n_58496), .Z(n_167488959
		));
	notech_reg_set divq_reg_21(.CP(n_62385), .D(n_21723), .SD(1'b1), .Q(divq
		[21]));
	notech_mux2 i_7998(.S(n_54360), .A(divq[21]), .B(n_8417), .Z(n_21723));
	notech_or2 i_218636976(.A(n_271888737), .B(n_55430), .Z(n_167388960));
	notech_reg_set divq_reg_22(.CP(n_62385), .D(n_21729), .SD(1'b1), .Q(divq
		[22]));
	notech_mux2 i_8006(.S(n_54360), .A(divq[22]), .B(n_8422), .Z(n_21729));
	notech_nand3 i_1516184(.A(n_1831), .B(n_167288961), .C(n_165688973), .Z(n_14176
		));
	notech_reg_set divq_reg_23(.CP(n_62385), .D(n_21735), .SD(1'b1), .Q(divq
		[23]));
	notech_mux2 i_8014(.S(n_54360), .A(divq[23]), .B(n_8427), .Z(n_21735));
	notech_nand2 i_166437492(.A(n_272388732), .B(opb[14]), .Z(n_167288961)
		);
	notech_reg_set divq_reg_24(.CP(n_62385), .D(n_21741), .SD(1'b1), .Q(divq
		[24]));
	notech_mux2 i_8023(.S(n_54360), .A(divq[24]), .B(n_8432), .Z(n_21741));
	notech_nao3 i_166337493(.A(imm[46]), .B(n_26795), .C(n_2198), .Z(n_1671)
		);
	notech_reg_set divq_reg_25(.CP(n_62385), .D(n_21747), .SD(1'b1), .Q(divq
		[25]));
	notech_mux2 i_8031(.S(n_54360), .A(divq[25]), .B(n_8437), .Z(n_21747));
	notech_reg_set divq_reg_26(.CP(n_62385), .D(n_21753), .SD(1'b1), .Q(divq
		[26]));
	notech_mux2 i_8039(.S(n_54360), .A(divq[26]), .B(n_8442), .Z(n_21753));
	notech_reg_set divq_reg_27(.CP(n_62385), .D(n_21759), .SD(1'b1), .Q(divq
		[27]));
	notech_mux2 i_8047(.S(n_54360), .A(divq[27]), .B(n_8447), .Z(n_21759));
	notech_nao3 i_166037496(.A(n_57438), .B(nbus_138[14]), .C(n_2318), .Z(n_166888964
		));
	notech_reg_set divq_reg_28(.CP(n_62385), .D(n_21765), .SD(1'b1), .Q(divq
		[28]));
	notech_mux2 i_8055(.S(n_54360), .A(divq[28]), .B(n_8452), .Z(n_21765));
	notech_or2 i_165837498(.A(n_55204), .B(n_27533), .Z(n_166788965));
	notech_reg_set divq_reg_29(.CP(n_62385), .D(n_21771), .SD(1'b1), .Q(divq
		[29]));
	notech_mux2 i_8063(.S(n_54360), .A(divq[29]), .B(n_8457), .Z(n_21771));
	notech_reg_set divq_reg_30(.CP(n_62385), .D(n_21777), .SD(1'b1), .Q(divq
		[30]));
	notech_mux2 i_8071(.S(n_54360), .A(divq[30]), .B(n_8462), .Z(n_21777));
	notech_reg_set divq_reg_31(.CP(n_62385), .D(n_21783), .SD(1'b1), .Q(divq
		[31]));
	notech_mux2 i_8079(.S(n_54360), .A(divq[31]), .B(n_8467), .Z(n_21783));
	notech_reg_set divq_reg_32(.CP(n_62385), .D(n_21789), .SD(1'b1), .Q(divq
		[32]));
	notech_mux2 i_8087(.S(n_54353), .A(divq[32]), .B(n_8472), .Z(n_21789));
	notech_reg_set divq_reg_33(.CP(n_62347), .D(n_21795), .SD(1'b1), .Q(divq
		[33]));
	notech_mux2 i_8095(.S(n_54353), .A(divq[33]), .B(n_27075), .Z(n_21795)
		);
	notech_reg_set divq_reg_34(.CP(n_62385), .D(n_21801), .SD(1'b1), .Q(divq
		[34]));
	notech_mux2 i_8103(.S(n_54353), .A(divq[34]), .B(n_27077), .Z(n_21801)
		);
	notech_reg_set divq_reg_35(.CP(n_62349), .D(n_21807), .SD(1'b1), .Q(divq
		[35]));
	notech_mux2 i_8111(.S(n_54353), .A(divq[35]), .B(n_27078), .Z(n_21807)
		);
	notech_reg_set divq_reg_36(.CP(n_62349), .D(n_21813), .SD(1'b1), .Q(divq
		[36]));
	notech_mux2 i_8119(.S(n_54353), .A(divq[36]), .B(n_27079), .Z(n_21813)
		);
	notech_reg_set divq_reg_37(.CP(n_62349), .D(n_21819), .SD(1'b1), .Q(divq
		[37]));
	notech_mux2 i_8127(.S(n_54353), .A(divq[37]), .B(n_27080), .Z(n_21819)
		);
	notech_reg_set divq_reg_38(.CP(n_62349), .D(n_21825), .SD(1'b1), .Q(divq
		[38]));
	notech_mux2 i_8135(.S(n_54353), .A(divq[38]), .B(n_27082), .Z(n_21825)
		);
	notech_reg_set divq_reg_39(.CP(n_62349), .D(n_21831), .SD(1'b1), .Q(divq
		[39]));
	notech_mux2 i_8143(.S(n_54353), .A(divq[39]), .B(n_27083), .Z(n_21831)
		);
	notech_or2 i_165937497(.A(n_271888737), .B(n_55075), .Z(n_165688973));
	notech_reg_set divq_reg_40(.CP(n_62349), .D(n_21837), .SD(1'b1), .Q(divq
		[40]));
	notech_mux2 i_8151(.S(n_54353), .A(divq[40]), .B(n_27084), .Z(n_21837)
		);
	notech_and4 i_1521306(.A(n_1788), .B(n_164788981), .C(n_165488975), .D(n_165588974
		), .Z(n_20685));
	notech_reg_set divq_reg_41(.CP(n_62349), .D(n_21843), .SD(1'b1), .Q(divq
		[41]));
	notech_mux2 i_8159(.S(n_54353), .A(divq[41]), .B(n_27086), .Z(n_21843)
		);
	notech_or2 i_127637875(.A(n_55156), .B(n_271888737), .Z(n_165588974));
	notech_reg_set divq_reg_42(.CP(n_62349), .D(n_21849), .SD(1'b1), .Q(divq
		[42]));
	notech_mux2 i_8167(.S(n_54353), .A(divq[42]), .B(n_27087), .Z(n_21849)
		);
	notech_or4 i_127837873(.A(n_55958), .B(n_2255), .C(n_28065), .D(n_60507)
		, .Z(n_165488975));
	notech_reg_set divq_reg_43(.CP(n_62349), .D(n_21855), .SD(1'b1), .Q(divq
		[43]));
	notech_mux2 i_8175(.S(n_54353), .A(divq[43]), .B(n_27088), .Z(n_21855)
		);
	notech_nao3 i_127737874(.A(n_62427), .B(opc[14]), .C(n_248534111), .Z(n_1653
		));
	notech_reg_set divq_reg_44(.CP(n_62349), .D(n_21861), .SD(1'b1), .Q(divq
		[44]));
	notech_mux2 i_8183(.S(n_54353), .A(divq[44]), .B(n_27089), .Z(n_21861)
		);
	notech_nand3 i_127537876(.A(n_59780), .B(n_59899), .C(read_data[14]), .Z
		(n_165288976));
	notech_reg_set divq_reg_45(.CP(n_62349), .D(n_21867), .SD(1'b1), .Q(divq
		[45]));
	notech_mux2 i_8191(.S(n_54353), .A(divq[45]), .B(n_27090), .Z(n_21867)
		);
	notech_reg_set divq_reg_46(.CP(n_62349), .D(n_21873), .SD(1'b1), .Q(divq
		[46]));
	notech_mux2 i_8199(.S(n_54353), .A(divq[46]), .B(n_27091), .Z(n_21873)
		);
	notech_reg_set divq_reg_47(.CP(n_62349), .D(n_21879), .SD(1'b1), .Q(divq
		[47]));
	notech_mux2 i_8207(.S(n_54353), .A(divq[47]), .B(n_27092), .Z(n_21879)
		);
	notech_reg_set divq_reg_48(.CP(n_62349), .D(n_21885), .SD(1'b1), .Q(divq
		[48]));
	notech_mux2 i_8215(.S(n_54355), .A(divq[48]), .B(n_27094), .Z(n_21885)
		);
	notech_reg_set divq_reg_49(.CP(n_62349), .D(n_21891), .SD(1'b1), .Q(divq
		[49]));
	notech_mux2 i_8225(.S(n_54355), .A(divq[49]), .B(n_27097), .Z(n_21891)
		);
	notech_or2 i_127937872(.A(n_55952), .B(n_80913203), .Z(n_164788981));
	notech_reg_set divq_reg_50(.CP(n_62349), .D(n_21897), .SD(1'b1), .Q(divq
		[50]));
	notech_mux2 i_8234(.S(n_54355), .A(divq[50]), .B(n_27098), .Z(n_21897)
		);
	notech_reg_set divq_reg_51(.CP(n_62349), .D(n_21903), .SD(1'b1), .Q(divq
		[51]));
	notech_mux2 i_8242(.S(n_54355), .A(divq[51]), .B(n_27099), .Z(n_21903)
		);
	notech_reg_set divq_reg_52(.CP(n_62349), .D(n_21909), .SD(1'b1), .Q(divq
		[52]));
	notech_mux2 i_8250(.S(n_54355), .A(divq[52]), .B(n_27100), .Z(n_21909)
		);
	notech_reg_set divq_reg_53(.CP(n_62349), .D(n_21915), .SD(1'b1), .Q(divq
		[53]));
	notech_mux2 i_8258(.S(n_54355), .A(divq[53]), .B(n_27101), .Z(n_21915)
		);
	notech_reg_set divq_reg_54(.CP(n_62273), .D(n_21921), .SD(1'b1), .Q(divq
		[54]));
	notech_mux2 i_8266(.S(n_54355), .A(divq[54]), .B(n_27102), .Z(n_21921)
		);
	notech_reg_set divq_reg_55(.CP(n_62273), .D(n_21927), .SD(1'b1), .Q(divq
		[55]));
	notech_mux2 i_8274(.S(n_54355), .A(divq[55]), .B(n_27103), .Z(n_21927)
		);
	notech_reg_set divq_reg_56(.CP(n_62273), .D(n_21933), .SD(1'b1), .Q(divq
		[56]));
	notech_mux2 i_8282(.S(n_54355), .A(divq[56]), .B(n_27104), .Z(n_21933)
		);
	notech_reg_set divq_reg_57(.CP(n_62273), .D(n_21939), .SD(1'b1), .Q(divq
		[57]));
	notech_mux2 i_8290(.S(n_54355), .A(divq[57]), .B(n_27105), .Z(n_21939)
		);
	notech_reg_set divq_reg_58(.CP(n_62273), .D(n_21945), .SD(1'b1), .Q(divq
		[58]));
	notech_mux2 i_8298(.S(n_54355), .A(divq[58]), .B(n_27106), .Z(n_21945)
		);
	notech_reg_set divq_reg_59(.CP(n_62273), .D(n_21951), .SD(1'b1), .Q(divq
		[59]));
	notech_mux2 i_8306(.S(n_54355), .A(divq[59]), .B(n_27107), .Z(n_21951)
		);
	notech_reg_set divq_reg_60(.CP(n_62273), .D(n_21957), .SD(1'b1), .Q(divq
		[60]));
	notech_mux2 i_8314(.S(n_54355), .A(divq[60]), .B(n_27108), .Z(n_21957)
		);
	notech_reg_set divq_reg_61(.CP(n_62273), .D(n_21963), .SD(1'b1), .Q(divq
		[61]));
	notech_mux2 i_8322(.S(n_54355), .A(divq[61]), .B(n_27109), .Z(n_21963)
		);
	notech_reg_set divq_reg_62(.CP(n_62273), .D(n_21969), .SD(1'b1), .Q(divq
		[62]));
	notech_mux2 i_8330(.S(n_54355), .A(divq[62]), .B(n_27110), .Z(n_21969)
		);
	notech_reg_set divq_reg_63(.CP(n_62273), .D(n_21975), .SD(1'b1), .Q(divq
		[63]));
	notech_mux2 i_8338(.S(n_54355), .A(divq[63]), .B(n_335283327), .Z(n_21975
		));
	notech_reg_set divr_reg_0(.CP(n_62197), .D(n_21981), .SD(1'b1), .Q(divr[
		0]));
	notech_mux2 i_8346(.S(n_54399), .A(divr[0]), .B(n_17697), .Z(n_21981));
	notech_reg_set divr_reg_1(.CP(n_62273), .D(n_21987), .SD(1'b1), .Q(divr[
		1]));
	notech_mux2 i_8354(.S(n_54399), .A(divr[1]), .B(n_17702), .Z(n_21987));
	notech_reg_set divr_reg_2(.CP(n_62279), .D(n_21993), .SD(1'b1), .Q(divr[
		2]));
	notech_mux2 i_8362(.S(n_54399), .A(divr[2]), .B(n_17707), .Z(n_21993));
	notech_or4 i_1720636(.A(n_162988996), .B(n_176688913), .C(n_163088995), 
		.D(n_161989005), .Z(n_20207));
	notech_reg_set divr_reg_3(.CP(n_62199), .D(n_21999), .SD(1'b1), .Q(divr[
		3]));
	notech_mux2 i_8370(.S(n_54399), .A(divr[3]), .B(n_17712), .Z(n_21999));
	notech_nor2 i_76338351(.A(n_55811), .B(n_272088735), .Z(n_163088995));
	notech_reg_set divr_reg_4(.CP(n_62199), .D(n_22007), .SD(1'b1), .Q(divr[
		4]));
	notech_mux2 i_8378(.S(n_54399), .A(divr[4]), .B(n_17717), .Z(n_22007));
	notech_ao3 i_76438350(.A(opc_10[16]), .B(n_62405), .C(n_2211), .Z(n_162988996
		));
	notech_reg_set divr_reg_5(.CP(n_62199), .D(n_22015), .SD(1'b1), .Q(divr[
		5]));
	notech_mux2 i_8386(.S(n_54399), .A(divr[5]), .B(n_17722), .Z(n_22015));
	notech_nand2 i_76138353(.A(n_271788738), .B(n_55819), .Z(n_1628));
	notech_reg_set divr_reg_6(.CP(n_62199), .D(n_22021), .SD(1'b1), .Q(divr[
		6]));
	notech_mux2 i_8394(.S(n_54399), .A(divr[6]), .B(n_17727), .Z(n_22021));
	notech_reg_set divr_reg_7(.CP(n_62199), .D(n_22027), .SD(1'b1), .Q(divr[
		7]));
	notech_mux2 i_8402(.S(n_54399), .A(divr[7]), .B(n_17732), .Z(n_22027));
	notech_reg_set divr_reg_8(.CP(n_62199), .D(n_22033), .SD(1'b1), .Q(divr[
		8]));
	notech_mux2 i_8410(.S(n_54399), .A(divr[8]), .B(n_17737), .Z(n_22033));
	notech_reg_set divr_reg_9(.CP(n_62199), .D(n_22039), .SD(1'b1), .Q(divr[
		9]));
	notech_mux2 i_8418(.S(n_54399), .A(divr[9]), .B(n_17742), .Z(n_22039));
	notech_reg_set divr_reg_10(.CP(n_62199), .D(n_22045), .SD(1'b1), .Q(divr
		[10]));
	notech_mux2 i_8426(.S(n_54399), .A(divr[10]), .B(n_17747), .Z(n_22045)
		);
	notech_reg_set divr_reg_11(.CP(n_62199), .D(n_22052), .SD(1'b1), .Q(divr
		[11]));
	notech_mux2 i_8434(.S(n_54399), .A(divr[11]), .B(n_17752), .Z(n_22052)
		);
	notech_reg_set divr_reg_12(.CP(n_62199), .D(n_22059), .SD(1'b1), .Q(divr
		[12]));
	notech_mux2 i_8442(.S(n_54399), .A(divr[12]), .B(n_17757), .Z(n_22059)
		);
	notech_reg_set divr_reg_13(.CP(n_62281), .D(n_22065), .SD(1'b1), .Q(divr
		[13]));
	notech_mux2 i_8450(.S(n_54399), .A(divr[13]), .B(n_17762), .Z(n_22065)
		);
	notech_reg_set divr_reg_14(.CP(n_62281), .D(n_22071), .SD(1'b1), .Q(divr
		[14]));
	notech_mux2 i_8458(.S(n_54399), .A(divr[14]), .B(n_17767), .Z(n_22071)
		);
	notech_nor2 i_76238352(.A(n_55587), .B(n_271988736), .Z(n_161989005));
	notech_reg_set divr_reg_15(.CP(n_62281), .D(n_22077), .SD(1'b1), .Q(divr
		[15]));
	notech_mux2 i_8466(.S(n_54399), .A(divr[15]), .B(n_17772), .Z(n_22077)
		);
	notech_reg_set divr_reg_16(.CP(n_62281), .D(n_22083), .SD(1'b1), .Q(divr
		[16]));
	notech_mux2 i_8474(.S(n_54401), .A(divr[16]), .B(n_17777), .Z(n_22083)
		);
	notech_reg_set divr_reg_17(.CP(n_62281), .D(n_22089), .SD(1'b1), .Q(divr
		[17]));
	notech_mux2 i_8482(.S(n_54401), .A(divr[17]), .B(n_17782), .Z(n_22089)
		);
	notech_reg_set divr_reg_18(.CP(n_62281), .D(n_22095), .SD(1'b1), .Q(divr
		[18]));
	notech_mux2 i_8492(.S(n_54401), .A(divr[18]), .B(n_17787), .Z(n_22095)
		);
	notech_reg_set divr_reg_19(.CP(n_62281), .D(n_22101), .SD(1'b1), .Q(divr
		[19]));
	notech_mux2 i_8500(.S(n_54401), .A(divr[19]), .B(n_17792), .Z(n_22101)
		);
	notech_reg_set divr_reg_20(.CP(n_62281), .D(n_22107), .SD(1'b1), .Q(divr
		[20]));
	notech_mux2 i_8508(.S(n_54401), .A(divr[20]), .B(n_17797), .Z(n_22107)
		);
	notech_reg_set divr_reg_21(.CP(n_62281), .D(n_22113), .SD(1'b1), .Q(divr
		[21]));
	notech_mux2 i_8516(.S(n_54401), .A(divr[21]), .B(n_17802), .Z(n_22113)
		);
	notech_reg_set divr_reg_22(.CP(n_62281), .D(n_22120), .SD(1'b1), .Q(divr
		[22]));
	notech_mux2 i_8524(.S(n_54401), .A(divr[22]), .B(n_17807), .Z(n_22120)
		);
	notech_reg_set divr_reg_23(.CP(n_62281), .D(n_22129), .SD(1'b1), .Q(divr
		[23]));
	notech_mux2 i_8532(.S(n_54401), .A(divr[23]), .B(n_17812), .Z(n_22129)
		);
	notech_reg_set divr_reg_24(.CP(n_62281), .D(n_22138), .SD(1'b1), .Q(divr
		[24]));
	notech_mux2 i_8540(.S(n_54401), .A(divr[24]), .B(n_17817), .Z(n_22138)
		);
	notech_reg_set divr_reg_25(.CP(n_62281), .D(n_22145), .SD(1'b1), .Q(divr
		[25]));
	notech_mux2 i_8548(.S(n_54401), .A(divr[25]), .B(n_17822), .Z(n_22145)
		);
	notech_reg_set divr_reg_26(.CP(n_62281), .D(n_22152), .SD(1'b1), .Q(divr
		[26]));
	notech_mux2 i_8556(.S(n_54401), .A(divr[26]), .B(n_17827), .Z(n_22152)
		);
	notech_reg_set divr_reg_27(.CP(n_62281), .D(n_22159), .SD(1'b1), .Q(divr
		[27]));
	notech_mux2 i_8564(.S(n_54401), .A(divr[27]), .B(n_17832), .Z(n_22159)
		);
	notech_reg_set divr_reg_28(.CP(n_62281), .D(n_22165), .SD(1'b1), .Q(divr
		[28]));
	notech_mux2 i_8572(.S(n_54401), .A(divr[28]), .B(n_17837), .Z(n_22165)
		);
	notech_reg_set divr_reg_29(.CP(n_62281), .D(n_22173), .SD(1'b1), .Q(divr
		[29]));
	notech_mux2 i_8580(.S(n_54401), .A(divr[29]), .B(n_17842), .Z(n_22173)
		);
	notech_reg_set divr_reg_30(.CP(n_62281), .D(n_22180), .SD(1'b1), .Q(divr
		[30]));
	notech_mux2 i_8588(.S(n_54401), .A(divr[30]), .B(n_17847), .Z(n_22180)
		);
	notech_reg_set divr_reg_31(.CP(n_62281), .D(n_22187), .SD(1'b1), .Q(divr
		[31]));
	notech_mux2 i_8596(.S(n_54401), .A(divr[31]), .B(n_17852), .Z(n_22187)
		);
	notech_and2 i_9538998(.A(n_55332), .B(n_48510), .Z(n_1602));
	notech_reg_set divr_reg_32(.CP(n_62353), .D(n_22193), .SD(1'b1), .Q(divr
		[32]));
	notech_mux2 i_8604(.S(n_54394), .A(divr[32]), .B(n_17857), .Z(n_22193)
		);
	notech_reg_set divr_reg_33(.CP(n_62279), .D(n_22199), .SD(1'b1), .Q(divr
		[33]));
	notech_mux2 i_8612(.S(n_54394), .A(divr[33]), .B(n_17862), .Z(n_22199)
		);
	notech_or2 i_71238402(.A(n_56216), .B(n_55600), .Z(n_1600));
	notech_reg_set divr_reg_34(.CP(n_62353), .D(n_22205), .SD(1'b1), .Q(divr
		[34]));
	notech_mux2 i_8620(.S(n_54394), .A(divr[34]), .B(n_17867), .Z(n_22205)
		);
	notech_reg_set divr_reg_35(.CP(n_62353), .D(n_22211), .SD(1'b1), .Q(divr
		[35]));
	notech_mux2 i_8628(.S(n_54394), .A(divr[35]), .B(n_17872), .Z(n_22211)
		);
	notech_reg_set divr_reg_36(.CP(n_62353), .D(n_22217), .SD(1'b1), .Q(divr
		[36]));
	notech_mux2 i_8636(.S(n_54394), .A(divr[36]), .B(n_17877), .Z(n_22217)
		);
	notech_nao3 i_71338401(.A(n_2203), .B(n_56538), .C(n_2700), .Z(n_1597)
		);
	notech_reg_set divr_reg_37(.CP(n_62353), .D(n_22223), .SD(1'b1), .Q(divr
		[37]));
	notech_mux2 i_8644(.S(n_54394), .A(divr[37]), .B(n_17882), .Z(n_22223)
		);
	notech_reg_set divr_reg_38(.CP(n_62353), .D(n_22229), .SD(1'b1), .Q(divr
		[38]));
	notech_mux2 i_8652(.S(n_54394), .A(divr[38]), .B(n_17887), .Z(n_22229)
		);
	notech_reg_set divr_reg_39(.CP(n_62353), .D(n_22235), .SD(1'b1), .Q(divr
		[39]));
	notech_mux2 i_8660(.S(n_54394), .A(divr[39]), .B(n_17892), .Z(n_22235)
		);
	notech_reg_set divr_reg_40(.CP(n_62353), .D(n_22241), .SD(1'b1), .Q(divr
		[40]));
	notech_mux2 i_8668(.S(n_54394), .A(divr[40]), .B(n_17897), .Z(n_22241)
		);
	notech_reg_set divr_reg_41(.CP(n_62353), .D(n_22247), .SD(1'b1), .Q(divr
		[41]));
	notech_mux2 i_8676(.S(n_54394), .A(divr[41]), .B(n_17902), .Z(n_22247)
		);
	notech_reg_set divr_reg_42(.CP(n_62353), .D(n_22253), .SD(1'b1), .Q(divr
		[42]));
	notech_mux2 i_8684(.S(n_54394), .A(divr[42]), .B(n_17907), .Z(n_22253)
		);
	notech_reg_set divr_reg_43(.CP(n_62353), .D(n_22259), .SD(1'b1), .Q(divr
		[43]));
	notech_mux2 i_8692(.S(n_54394), .A(divr[43]), .B(n_17912), .Z(n_22259)
		);
	notech_reg_set divr_reg_44(.CP(n_62353), .D(n_22265), .SD(1'b1), .Q(divr
		[44]));
	notech_mux2 i_8700(.S(n_54394), .A(divr[44]), .B(n_17917), .Z(n_22265)
		);
	notech_reg_set divr_reg_45(.CP(n_62353), .D(n_22271), .SD(1'b1), .Q(divr
		[45]));
	notech_mux2 i_8708(.S(n_54394), .A(divr[45]), .B(n_17922), .Z(n_22271)
		);
	notech_reg_set divr_reg_46(.CP(n_62353), .D(n_22277), .SD(1'b1), .Q(divr
		[46]));
	notech_mux2 i_8716(.S(n_54394), .A(divr[46]), .B(n_17927), .Z(n_22277)
		);
	notech_reg_set divr_reg_47(.CP(n_62353), .D(n_22283), .SD(1'b1), .Q(divr
		[47]));
	notech_mux2 i_8724(.S(n_54394), .A(divr[47]), .B(n_17932), .Z(n_22283)
		);
	notech_reg_set divr_reg_48(.CP(n_62353), .D(n_22289), .SD(1'b1), .Q(divr
		[48]));
	notech_mux2 i_8734(.S(n_54396), .A(divr[48]), .B(n_17937), .Z(n_22289)
		);
	notech_reg_set divr_reg_49(.CP(n_62353), .D(n_22295), .SD(1'b1), .Q(divr
		[49]));
	notech_mux2 i_8742(.S(n_54396), .A(divr[49]), .B(n_17942), .Z(n_22295)
		);
	notech_reg_set divr_reg_50(.CP(n_62353), .D(n_22301), .SD(1'b1), .Q(divr
		[50]));
	notech_mux2 i_8751(.S(n_54396), .A(divr[50]), .B(n_17947), .Z(n_22301)
		);
	notech_reg_set divr_reg_51(.CP(n_62353), .D(n_22307), .SD(1'b1), .Q(divr
		[51]));
	notech_mux2 i_8759(.S(n_54396), .A(divr[51]), .B(n_17952), .Z(n_22307)
		);
	notech_reg_set divr_reg_52(.CP(n_62279), .D(n_22313), .SD(1'b1), .Q(divr
		[52]));
	notech_mux2 i_8767(.S(n_54396), .A(divr[52]), .B(n_17957), .Z(n_22313)
		);
	notech_reg_set divr_reg_53(.CP(n_62279), .D(n_22319), .SD(1'b1), .Q(divr
		[53]));
	notech_mux2 i_8775(.S(n_54396), .A(divr[53]), .B(n_17962), .Z(n_22319)
		);
	notech_reg_set divr_reg_54(.CP(n_62279), .D(n_22325), .SD(1'b1), .Q(divr
		[54]));
	notech_mux2 i_8783(.S(n_54396), .A(divr[54]), .B(n_17967), .Z(n_22325)
		);
	notech_reg_set divr_reg_55(.CP(n_62279), .D(n_22331), .SD(1'b1), .Q(divr
		[55]));
	notech_mux2 i_8791(.S(n_54396), .A(divr[55]), .B(n_17972), .Z(n_22331)
		);
	notech_reg_set divr_reg_56(.CP(n_62279), .D(n_22337), .SD(1'b1), .Q(divr
		[56]));
	notech_mux2 i_8799(.S(n_54396), .A(divr[56]), .B(n_17977), .Z(n_22337)
		);
	notech_reg_set divr_reg_57(.CP(n_62279), .D(n_22343), .SD(1'b1), .Q(divr
		[57]));
	notech_mux2 i_8807(.S(n_54396), .A(divr[57]), .B(n_17982), .Z(n_22343)
		);
	notech_reg_set divr_reg_58(.CP(n_62279), .D(n_22349), .SD(1'b1), .Q(divr
		[58]));
	notech_mux2 i_8815(.S(n_54396), .A(divr[58]), .B(n_17987), .Z(n_22349)
		);
	notech_reg_set divr_reg_59(.CP(n_62279), .D(n_22355), .SD(1'b1), .Q(divr
		[59]));
	notech_mux2 i_8823(.S(n_54396), .A(divr[59]), .B(n_17992), .Z(n_22355)
		);
	notech_reg_set divr_reg_60(.CP(n_62279), .D(n_22361), .SD(1'b1), .Q(divr
		[60]));
	notech_mux2 i_8831(.S(n_54396), .A(divr[60]), .B(n_17997), .Z(n_22361)
		);
	notech_reg_set divr_reg_61(.CP(n_62279), .D(n_22367), .SD(1'b1), .Q(divr
		[61]));
	notech_mux2 i_8839(.S(n_54396), .A(divr[61]), .B(n_18002), .Z(n_22367)
		);
	notech_reg_set divr_reg_62(.CP(n_62199), .D(n_22373), .SD(1'b1), .Q(divr
		[62]));
	notech_mux2 i_8847(.S(n_54396), .A(divr[62]), .B(n_18007), .Z(n_22373)
		);
	notech_reg_set divr_reg_63(.CP(n_62199), .D(n_22379), .SD(1'b1), .Q(divr
		[63]));
	notech_mux2 i_8855(.S(n_54396), .A(divr[63]), .B(n_18012), .Z(n_22379)
		);
	notech_reg_set opd_reg_0(.CP(n_62283), .D(n_22385), .SD(1'b1), .Q(opd[0]
		));
	notech_mux2 i_8863(.S(\nbus_11355[0] ), .A(opd[0]), .B(n_21122), .Z(n_22385
		));
	notech_reg_set opd_reg_1(.CP(n_62201), .D(n_22391), .SD(1'b1), .Q(opd[1]
		));
	notech_mux2 i_8871(.S(\nbus_11355[0] ), .A(opd[1]), .B(n_27114), .Z(n_22391
		));
	notech_reg_set opd_reg_2(.CP(n_62201), .D(n_22397), .SD(1'b1), .Q(opd[2]
		));
	notech_mux2 i_8879(.S(\nbus_11355[0] ), .A(opd[2]), .B(n_21132), .Z(n_22397
		));
	notech_reg_set opd_reg_3(.CP(n_62201), .D(n_22403), .SD(1'b1), .Q(opd[3]
		));
	notech_mux2 i_8887(.S(\nbus_11355[0] ), .A(opd[3]), .B(n_21137), .Z(n_22403
		));
	notech_reg_set opd_reg_4(.CP(n_62201), .D(n_22409), .SD(1'b1), .Q(opd[4]
		));
	notech_mux2 i_8895(.S(\nbus_11355[0] ), .A(opd[4]), .B(n_21142), .Z(n_22409
		));
	notech_reg_set opd_reg_5(.CP(n_62201), .D(n_22415), .SD(1'b1), .Q(opd[5]
		));
	notech_mux2 i_8903(.S(\nbus_11355[0] ), .A(opd[5]), .B(n_21147), .Z(n_22415
		));
	notech_reg_set opd_reg_6(.CP(n_62201), .D(n_22421), .SD(1'b1), .Q(opd[6]
		));
	notech_mux2 i_8911(.S(n_57470), .A(n_27115), .B(opd[6]), .Z(n_22421));
	notech_reg_set opd_reg_7(.CP(n_62201), .D(n_22427), .SD(1'b1), .Q(opd[7]
		));
	notech_mux2 i_8919(.S(n_57470), .A(n_27116), .B(opd[7]), .Z(n_22427));
	notech_nao3 i_17238921(.A(n_27517), .B(opz[1]), .C(opz[2]), .Z(n_1562)
		);
	notech_reg_set opd_reg_8(.CP(n_62201), .D(n_22433), .SD(1'b1), .Q(opd[8]
		));
	notech_mux2 i_8927(.S(n_57470), .A(n_27117), .B(opd[8]), .Z(n_22433));
	notech_reg_set opd_reg_9(.CP(n_62201), .D(n_22439), .SD(1'b1), .Q(opd[9]
		));
	notech_mux2 i_8935(.S(n_57470), .A(n_27118), .B(opd[9]), .Z(n_22439));
	notech_reg_set opd_reg_10(.CP(n_62201), .D(n_22445), .SD(1'b1), .Q(opd[
		10]));
	notech_mux2 i_8943(.S(n_57470), .A(n_27119), .B(opd[10]), .Z(n_22445));
	notech_reg_set opd_reg_11(.CP(n_62283), .D(n_22451), .SD(1'b1), .Q(opd[
		11]));
	notech_mux2 i_8952(.S(n_57470), .A(n_27120), .B(opd[11]), .Z(n_22451));
	notech_reg_set opd_reg_12(.CP(n_62283), .D(n_22457), .SD(1'b1), .Q(opd[
		12]));
	notech_mux2 i_8960(.S(n_57470), .A(n_27121), .B(opd[12]), .Z(n_22457));
	notech_reg_set opd_reg_13(.CP(n_62283), .D(n_22463), .SD(1'b1), .Q(opd[
		13]));
	notech_mux2 i_8968(.S(n_57470), .A(n_27122), .B(opd[13]), .Z(n_22463));
	notech_reg_set opd_reg_14(.CP(n_62283), .D(n_22469), .SD(1'b1), .Q(opd[
		14]));
	notech_mux2 i_8976(.S(n_57470), .A(n_27123), .B(opd[14]), .Z(n_22469));
	notech_reg_set opd_reg_15(.CP(n_62283), .D(n_22475), .SD(1'b1), .Q(opd[
		15]));
	notech_mux2 i_8984(.S(n_57470), .A(n_27124), .B(opd[15]), .Z(n_22475));
	notech_reg_set opd_reg_16(.CP(n_62283), .D(n_22481), .SD(1'b1), .Q(opd[
		16]));
	notech_mux2 i_8992(.S(\nbus_11355[16] ), .A(opd[16]), .B(n_21202), .Z(n_22481
		));
	notech_reg_set opd_reg_17(.CP(n_62283), .D(n_22487), .SD(1'b1), .Q(opd[
		17]));
	notech_mux2 i_9000(.S(\nbus_11355[16] ), .A(opd[17]), .B(n_21207), .Z(n_22487
		));
	notech_reg_set opd_reg_18(.CP(n_62283), .D(n_22493), .SD(1'b1), .Q(opd[
		18]));
	notech_mux2 i_9008(.S(\nbus_11355[16] ), .A(opd[18]), .B(n_21212), .Z(n_22493
		));
	notech_reg_set opd_reg_19(.CP(n_62283), .D(n_22499), .SD(1'b1), .Q(opd[
		19]));
	notech_mux2 i_9016(.S(\nbus_11355[16] ), .A(opd[19]), .B(n_21217), .Z(n_22499
		));
	notech_reg_set opd_reg_20(.CP(n_62283), .D(n_22505), .SD(1'b1), .Q(opd[
		20]));
	notech_mux2 i_9024(.S(\nbus_11355[16] ), .A(opd[20]), .B(n_21222), .Z(n_22505
		));
	notech_reg_set opd_reg_21(.CP(n_62283), .D(n_22511), .SD(1'b1), .Q(opd[
		21]));
	notech_mux2 i_9032(.S(\nbus_11355[16] ), .A(opd[21]), .B(n_21227), .Z(n_22511
		));
	notech_reg_set opd_reg_22(.CP(n_62283), .D(n_22517), .SD(1'b1), .Q(opd[
		22]));
	notech_mux2 i_9040(.S(\nbus_11355[16] ), .A(opd[22]), .B(n_21232), .Z(n_22517
		));
	notech_reg_set opd_reg_23(.CP(n_62283), .D(n_22523), .SD(1'b1), .Q(opd[
		23]));
	notech_mux2 i_9048(.S(\nbus_11355[16] ), .A(opd[23]), .B(n_21237), .Z(n_22523
		));
	notech_reg_set opd_reg_24(.CP(n_62283), .D(n_22529), .SD(1'b1), .Q(opd[
		24]));
	notech_mux2 i_9056(.S(\nbus_11355[16] ), .A(opd[24]), .B(n_21242), .Z(n_22529
		));
	notech_reg_set opd_reg_25(.CP(n_62283), .D(n_22535), .SD(1'b1), .Q(opd[
		25]));
	notech_mux2 i_9064(.S(\nbus_11355[16] ), .A(opd[25]), .B(n_21247), .Z(n_22535
		));
	notech_reg_set opd_reg_26(.CP(n_62283), .D(n_22541), .SD(1'b1), .Q(opd[
		26]));
	notech_mux2 i_9072(.S(\nbus_11355[16] ), .A(opd[26]), .B(n_21252), .Z(n_22541
		));
	notech_reg_set opd_reg_27(.CP(n_62283), .D(n_22547), .SD(1'b1), .Q(opd[
		27]));
	notech_mux2 i_9080(.S(\nbus_11355[16] ), .A(opd[27]), .B(n_21257), .Z(n_22547
		));
	notech_reg_set opd_reg_28(.CP(n_62283), .D(n_22553), .SD(1'b1), .Q(opd[
		28]));
	notech_mux2 i_9089(.S(\nbus_11355[16] ), .A(opd[28]), .B(n_21262), .Z(n_22553
		));
	notech_reg_set opd_reg_29(.CP(n_62201), .D(n_22559), .SD(1'b1), .Q(opd[
		29]));
	notech_mux2 i_9097(.S(\nbus_11355[16] ), .A(opd[29]), .B(n_21267), .Z(n_22559
		));
	notech_reg_set opd_reg_30(.CP(n_62201), .D(n_22565), .SD(1'b1), .Q(opd[
		30]));
	notech_mux2 i_9105(.S(\nbus_11355[16] ), .A(opd[30]), .B(n_21272), .Z(n_22565
		));
	notech_reg_set opd_reg_31(.CP(n_62203), .D(n_22571), .SD(1'b1), .Q(opd[
		31]));
	notech_mux2 i_9113(.S(\nbus_11355[16] ), .A(opd[31]), .B(n_27125), .Z(n_22571
		));
	notech_reg regs_reg_1_0(.CP(n_62203), .D(n_22577), .CD(n_61119), .Q(ecx[
		0]));
	notech_mux2 i_9121(.S(\nbus_11305[0] ), .A(ecx[0]), .B(n_11692), .Z(n_22577
		));
	notech_reg regs_reg_1_1(.CP(n_62203), .D(n_22583), .CD(n_61115), .Q(ecx[
		1]));
	notech_mux2 i_9129(.S(\nbus_11305[0] ), .A(ecx[1]), .B(n_27126), .Z(n_22583
		));
	notech_reg regs_reg_1_2(.CP(n_62203), .D(n_22589), .CD(n_61118), .Q(ecx[
		2]));
	notech_mux2 i_9137(.S(\nbus_11305[0] ), .A(ecx[2]), .B(n_27127), .Z(n_22589
		));
	notech_reg regs_reg_1_3(.CP(n_62203), .D(n_22595), .CD(n_61115), .Q(ecx[
		3]));
	notech_mux2 i_9145(.S(\nbus_11305[0] ), .A(ecx[3]), .B(n_27128), .Z(n_22595
		));
	notech_reg regs_reg_1_4(.CP(n_62203), .D(n_22601), .CD(n_61115), .Q(ecx[
		4]));
	notech_mux2 i_9153(.S(\nbus_11305[0] ), .A(ecx[4]), .B(n_27129), .Z(n_22601
		));
	notech_reg regs_reg_1_5(.CP(n_62203), .D(n_22607), .CD(n_61118), .Q(ecx[
		5]));
	notech_mux2 i_9161(.S(\nbus_11305[0] ), .A(ecx[5]), .B(n_27130), .Z(n_22607
		));
	notech_reg regs_reg_1_6(.CP(n_62203), .D(n_22613), .CD(n_61118), .Q(ecx[
		6]));
	notech_mux2 i_9169(.S(\nbus_11305[0] ), .A(ecx[6]), .B(n_27131), .Z(n_22613
		));
	notech_reg regs_reg_1_7(.CP(n_62203), .D(n_22619), .CD(n_61118), .Q(ecx[
		7]));
	notech_mux2 i_9177(.S(\nbus_11305[0] ), .A(ecx[7]), .B(n_27132), .Z(n_22619
		));
	notech_reg regs_reg_1_8(.CP(n_62203), .D(n_22625), .CD(n_61118), .Q(ecx[
		8]));
	notech_mux2 i_9185(.S(\nbus_11305[0] ), .A(ecx[8]), .B(n_11740), .Z(n_22625
		));
	notech_or4 i_28524(.A(n_56487), .B(n_56478), .C(n_56449), .D(n_60507), .Z
		(n_1529));
	notech_reg regs_reg_1_9(.CP(n_62203), .D(n_22631), .CD(n_61118), .Q(ecx[
		9]));
	notech_mux2 i_9193(.S(\nbus_11305[0] ), .A(ecx[9]), .B(n_27133), .Z(n_22631
		));
	notech_reg regs_reg_1_10(.CP(n_62203), .D(n_22638), .CD(n_61114), .Q(ecx
		[10]));
	notech_mux2 i_9201(.S(\nbus_11305[0] ), .A(ecx[10]), .B(n_27134), .Z(n_22638
		));
	notech_and3 i_99441276(.A(n_55667), .B(n_1526), .C(n_1022), .Z(n_1527)
		);
	notech_reg regs_reg_1_11(.CP(n_62203), .D(n_22647), .CD(n_61110), .Q(ecx
		[11]));
	notech_mux2 i_9209(.S(\nbus_11305[0] ), .A(ecx[11]), .B(n_11758), .Z(n_22647
		));
	notech_and3 i_90342243(.A(n_55658), .B(n_1021), .C(n_56001), .Z(n_1526)
		);
	notech_reg regs_reg_1_12(.CP(n_62203), .D(n_22657), .CD(n_61112), .Q(ecx
		[12]));
	notech_mux2 i_9217(.S(\nbus_11305[0] ), .A(ecx[12]), .B(n_11764), .Z(n_22657
		));
	notech_reg regs_reg_1_13(.CP(n_62203), .D(n_22665), .CD(n_61110), .Q(ecx
		[13]));
	notech_mux2 i_9225(.S(\nbus_11305[0] ), .A(ecx[13]), .B(n_11770), .Z(n_22665
		));
	notech_reg regs_reg_1_14(.CP(n_62203), .D(n_22671), .CD(n_61110), .Q(ecx
		[14]));
	notech_mux2 i_9233(.S(\nbus_11305[0] ), .A(ecx[14]), .B(n_11776), .Z(n_22671
		));
	notech_ao4 i_200443429(.A(n_56246), .B(n_28993), .C(n_56235), .D(n_27744
		), .Z(n_1523));
	notech_reg regs_reg_1_15(.CP(n_62203), .D(n_22677), .CD(n_61112), .Q(ecx
		[15]));
	notech_mux2 i_9241(.S(\nbus_11305[0] ), .A(ecx[15]), .B(n_11782), .Z(n_22677
		));
	notech_ao4 i_200543428(.A(n_56255), .B(n_27815), .C(n_27847), .D(n_57358
		), .Z(n_1522));
	notech_reg regs_reg_1_16(.CP(n_62203), .D(n_22683), .CD(n_61112), .Q(ecx
		[16]));
	notech_mux2 i_9249(.S(\nbus_11305[16] ), .A(ecx[16]), .B(n_11788), .Z(n_22683
		));
	notech_and2 i_200943424(.A(n_1520), .B(n_1519), .Z(n_1521));
	notech_reg regs_reg_1_17(.CP(n_62203), .D(n_22689), .CD(n_61112), .Q(ecx
		[17]));
	notech_mux2 i_9257(.S(\nbus_11305[16] ), .A(ecx[17]), .B(n_11794), .Z(n_22689
		));
	notech_ao4 i_200743426(.A(n_56226), .B(n_28016), .C(n_57338), .D(n_27783
		), .Z(n_1520));
	notech_reg regs_reg_1_18(.CP(n_62153), .D(n_22695), .CD(n_61112), .Q(ecx
		[18]));
	notech_mux2 i_9265(.S(\nbus_11305[16] ), .A(ecx[18]), .B(n_11800), .Z(n_22695
		));
	notech_ao4 i_200843425(.A(n_56409), .B(n_27982), .C(n_56305), .D(n_27635
		), .Z(n_1519));
	notech_reg regs_reg_1_19(.CP(n_62153), .D(n_22701), .CD(n_61112), .Q(ecx
		[19]));
	notech_mux2 i_9273(.S(\nbus_11305[16] ), .A(ecx[19]), .B(n_27135), .Z(n_22701
		));
	notech_and4 i_201743416(.A(n_1516), .B(n_1515), .C(n_1513), .D(n_1512), 
		.Z(n_1518));
	notech_reg regs_reg_1_20(.CP(n_62153), .D(n_22708), .CD(n_61110), .Q(ecx
		[20]));
	notech_mux2 i_9282(.S(\nbus_11305[16] ), .A(ecx[20]), .B(n_27136), .Z(n_22708
		));
	notech_reg regs_reg_1_21(.CP(n_62153), .D(n_22714), .CD(n_61110), .Q(ecx
		[21]));
	notech_mux2 i_9290(.S(\nbus_11305[16] ), .A(ecx[21]), .B(n_11818), .Z(n_22714
		));
	notech_ao4 i_201143422(.A(n_56296), .B(n_27950), .C(n_56395), .D(n_28992
		), .Z(n_1516));
	notech_reg regs_reg_1_22(.CP(n_62153), .D(n_22720), .CD(n_61110), .Q(ecx
		[22]));
	notech_mux2 i_9298(.S(\nbus_11305[16] ), .A(ecx[22]), .B(n_11824), .Z(n_22720
		));
	notech_ao4 i_201243421(.A(n_60479), .B(n_27916), .C(n_56285), .D(n_27677
		), .Z(n_1515));
	notech_reg regs_reg_1_23(.CP(n_62153), .D(n_22726), .CD(n_61110), .Q(ecx
		[23]));
	notech_mux2 i_9306(.S(\nbus_11305[16] ), .A(ecx[23]), .B(n_27137), .Z(n_22726
		));
	notech_reg regs_reg_1_24(.CP(n_62153), .D(n_22732), .CD(n_61110), .Q(ecx
		[24]));
	notech_mux2 i_9315(.S(\nbus_11305[16] ), .A(ecx[24]), .B(n_27138), .Z(n_22732
		));
	notech_ao4 i_201443419(.A(n_56276), .B(n_27882), .C(n_56265), .D(n_27712
		), .Z(n_1513));
	notech_reg regs_reg_1_25(.CP(n_62153), .D(n_22738), .CD(n_61110), .Q(ecx
		[25]));
	notech_mux2 i_9323(.S(\nbus_11305[16] ), .A(ecx[25]), .B(n_27139), .Z(n_22738
		));
	notech_ao4 i_201543418(.A(n_59219), .B(n_28048), .C(n_57367), .D(n_27399
		), .Z(n_1512));
	notech_reg regs_reg_1_26(.CP(n_62153), .D(n_22744), .CD(n_61110), .Q(ecx
		[26]));
	notech_mux2 i_9331(.S(\nbus_11305[16] ), .A(ecx[26]), .B(n_11848), .Z(n_22744
		));
	notech_reg regs_reg_1_27(.CP(n_62153), .D(n_22750), .CD(n_61110), .Q(ecx
		[27]));
	notech_mux2 i_9339(.S(\nbus_11305[16] ), .A(ecx[27]), .B(n_11854), .Z(n_22750
		));
	notech_ao4 i_202343410(.A(n_55667), .B(n_60584), .C(n_303321920), .D(n_26581
		), .Z(n_1510));
	notech_reg regs_reg_1_28(.CP(n_62153), .D(n_22756), .CD(n_61110), .Q(ecx
		[28]));
	notech_mux2 i_9347(.S(\nbus_11305[16] ), .A(ecx[28]), .B(n_27140), .Z(n_22756
		));
	notech_reg regs_reg_1_29(.CP(n_62153), .D(n_22762), .CD(n_61112), .Q(ecx
		[29]));
	notech_mux2 i_9355(.S(\nbus_11305[16] ), .A(ecx[29]), .B(n_11866), .Z(n_22762
		));
	notech_reg regs_reg_1_30(.CP(n_62369), .D(n_22768), .CD(n_61113), .Q(ecx
		[30]));
	notech_mux2 i_9363(.S(\nbus_11305[16] ), .A(ecx[30]), .B(n_27141), .Z(n_22768
		));
	notech_reg regs_reg_1_31(.CP(n_62077), .D(n_22774), .CD(n_61113), .Q(ecx
		[31]));
	notech_mux2 i_9371(.S(\nbus_11305[16] ), .A(ecx[31]), .B(n_11878), .Z(n_22774
		));
	notech_reg sign_div_reg(.CP(n_62077), .D(n_22780), .CD(n_61113), .Q(sign_div
		));
	notech_mux2 i_9379(.S(n_301286332), .A(n_26586), .B(sign_div), .Z(n_22780
		));
	notech_reg_set opc_reg_0(.CP(n_62077), .D(n_22786), .SD(1'b1), .Q(opc[0]
		));
	notech_mux2 i_9387(.S(n_27142), .A(opc[0]), .B(n_9707), .Z(n_22786));
	notech_reg_set opc_reg_1(.CP(n_62077), .D(n_22792), .SD(1'b1), .Q(opc[1]
		));
	notech_mux2 i_9395(.S(n_27142), .A(opc[1]), .B(n_9712), .Z(n_22792));
	notech_reg_set opc_reg_2(.CP(n_62077), .D(n_22798), .SD(1'b1), .Q(opc[2]
		));
	notech_mux2 i_9403(.S(n_27142), .A(opc[2]), .B(n_9717), .Z(n_22798));
	notech_reg_set opc_reg_3(.CP(n_62077), .D(n_22804), .SD(1'b1), .Q(opc[3]
		));
	notech_mux2 i_9411(.S(n_27142), .A(opc[3]), .B(n_9722), .Z(n_22804));
	notech_reg_set opc_reg_4(.CP(n_62077), .D(n_22810), .SD(1'b1), .Q(opc[4]
		));
	notech_mux2 i_9419(.S(n_27142), .A(opc[4]), .B(n_9727), .Z(n_22810));
	notech_reg_set opc_reg_5(.CP(n_62077), .D(n_22816), .SD(1'b1), .Q(opc[5]
		));
	notech_mux2 i_9427(.S(n_27143), .A(opc[5]), .B(n_9732), .Z(n_22816));
	notech_reg_set opc_reg_6(.CP(n_62077), .D(n_22822), .SD(1'b1), .Q(opc[6]
		));
	notech_mux2 i_9435(.S(n_27143), .A(opc[6]), .B(n_9737), .Z(n_22822));
	notech_reg_set opc_reg_7(.CP(n_62173), .D(n_22828), .SD(1'b1), .Q(opc[7]
		));
	notech_mux2 i_9443(.S(n_27143), .A(opc[7]), .B(n_9742), .Z(n_22828));
	notech_reg_set opc_reg_8(.CP(n_62173), .D(n_22834), .SD(1'b1), .Q(opc[8]
		));
	notech_mux2 i_9451(.S(n_27144), .A(opc[8]), .B(n_9747), .Z(n_22834));
	notech_reg_set opc_reg_9(.CP(n_62173), .D(n_22840), .SD(1'b1), .Q(opc[9]
		));
	notech_mux2 i_9459(.S(n_27144), .A(opc[9]), .B(n_9752), .Z(n_22840));
	notech_reg_set opc_reg_10(.CP(n_62173), .D(n_22846), .SD(1'b1), .Q(opc[
		10]));
	notech_mux2 i_9467(.S(n_27144), .A(opc[10]), .B(n_9757), .Z(n_22846));
	notech_reg_set opc_reg_11(.CP(n_62173), .D(n_22852), .SD(1'b1), .Q(opc[
		11]));
	notech_mux2 i_9475(.S(n_27144), .A(opc[11]), .B(n_9762), .Z(n_22852));
	notech_reg_set opc_reg_12(.CP(n_62173), .D(n_22858), .SD(1'b1), .Q(opc[
		12]));
	notech_mux2 i_9483(.S(n_27144), .A(opc[12]), .B(n_9767), .Z(n_22858));
	notech_and3 i_246545372(.A(n_54851), .B(n_54900), .C(n_1510), .Z(n_1492)
		);
	notech_reg_set opc_reg_13(.CP(n_62173), .D(n_22864), .SD(1'b1), .Q(opc[
		13]));
	notech_mux2 i_9491(.S(n_27144), .A(opc[13]), .B(n_9772), .Z(n_22864));
	notech_or2 i_89345431(.A(n_1492), .B(n_317888511), .Z(n_1491));
	notech_reg_set opc_reg_14(.CP(n_62173), .D(n_22870), .SD(1'b1), .Q(opc[
		14]));
	notech_mux2 i_9499(.S(n_27144), .A(opc[14]), .B(n_9777), .Z(n_22870));
	notech_reg_set opc_reg_15(.CP(n_62173), .D(n_22876), .SD(1'b1), .Q(opc[
		15]));
	notech_mux2 i_9507(.S(n_27144), .A(opc[15]), .B(n_9782), .Z(n_22876));
	notech_reg_set opc_reg_16(.CP(n_62173), .D(n_22882), .SD(1'b1), .Q(opc[
		16]));
	notech_mux2 i_9515(.S(n_27145), .A(opc[16]), .B(n_9787), .Z(n_22882));
	notech_reg_set opc_reg_17(.CP(n_62173), .D(n_22888), .SD(1'b1), .Q(opc[
		17]));
	notech_mux2 i_9523(.S(n_27145), .A(opc[17]), .B(n_9792), .Z(n_22888));
	notech_and4 i_88348326(.A(n_1480), .B(n_1479), .C(n_1485), .D(n_1383), .Z
		(n_1487));
	notech_reg_set opc_reg_18(.CP(n_62173), .D(n_22894), .SD(1'b1), .Q(opc[
		18]));
	notech_mux2 i_9531(.S(n_27145), .A(opc[18]), .B(n_9797), .Z(n_22894));
	notech_reg_set opc_reg_19(.CP(n_62173), .D(n_22900), .SD(1'b1), .Q(opc[
		19]));
	notech_mux2 i_9539(.S(n_27145), .A(opc[19]), .B(n_9802), .Z(n_22900));
	notech_and3 i_88148328(.A(n_1483), .B(n_148289037), .C(n_1382), .Z(n_1485
		));
	notech_reg_set opc_reg_20(.CP(n_62173), .D(n_22906), .SD(1'b1), .Q(opc[
		20]));
	notech_mux2 i_9547(.S(n_27145), .A(opc[20]), .B(n_9807), .Z(n_22906));
	notech_reg_set opc_reg_21(.CP(n_62173), .D(n_22912), .SD(1'b1), .Q(opc[
		21]));
	notech_mux2 i_9555(.S(n_27145), .A(opc[21]), .B(n_9812), .Z(n_22912));
	notech_ao4 i_87448334(.A(n_54024), .B(n_28999), .C(n_321688474), .D(n_28998
		), .Z(n_1483));
	notech_reg_set opc_reg_22(.CP(n_62173), .D(n_22918), .SD(1'b1), .Q(opc[
		22]));
	notech_mux2 i_9565(.S(n_27145), .A(opc[22]), .B(n_9817), .Z(n_22918));
	notech_ao4 i_87848331(.A(n_56901), .B(n_317288517), .C(n_28997), .D(n_1491
		), .Z(n_148289037));
	notech_reg_set opc_reg_23(.CP(n_62173), .D(n_22924), .SD(1'b1), .Q(opc[
		23]));
	notech_mux2 i_9573(.S(n_27145), .A(opc[23]), .B(n_9822), .Z(n_22924));
	notech_reg_set opc_reg_24(.CP(n_62173), .D(n_22930), .SD(1'b1), .Q(opc[
		24]));
	notech_mux2 i_9581(.S(n_27145), .A(opc[24]), .B(n_9827), .Z(n_22930));
	notech_ao4 i_87648332(.A(n_317488515), .B(n_55234), .C(n_320088489), .D(n_27599
		), .Z(n_1480));
	notech_reg_set opc_reg_25(.CP(n_62173), .D(n_22936), .SD(1'b1), .Q(opc[
		25]));
	notech_mux2 i_9589(.S(n_27145), .A(opc[25]), .B(n_9832), .Z(n_22936));
	notech_ao4 i_87548333(.A(n_59163), .B(n_27553), .C(n_55133), .D(n_59050)
		, .Z(n_1479));
	notech_reg_set opc_reg_26(.CP(n_62171), .D(n_22942), .SD(1'b1), .Q(opc[
		26]));
	notech_mux2 i_9597(.S(n_27145), .A(opc[26]), .B(n_9837), .Z(n_22942));
	notech_and3 i_48849180(.A(n_1373), .B(n_1477), .C(n_1370), .Z(n_82622813
		));
	notech_reg_set opc_reg_27(.CP(n_62171), .D(n_22948), .SD(1'b1), .Q(opc[
		27]));
	notech_mux2 i_9605(.S(n_27145), .A(opc[27]), .B(n_9842), .Z(n_22948));
	notech_reg_set opc_reg_28(.CP(n_62243), .D(n_22954), .SD(1'b1), .Q(opc[
		28]));
	notech_mux2 i_9613(.S(n_27145), .A(opc[28]), .B(n_9847), .Z(n_22954));
	notech_ao4 i_85848348(.A(n_55234), .B(n_56022), .C(n_28997), .D(n_55978)
		, .Z(n_1477));
	notech_reg_set opc_reg_29(.CP(n_62243), .D(n_22960), .SD(1'b1), .Q(opc[
		29]));
	notech_mux2 i_9621(.S(n_27145), .A(opc[29]), .B(n_9852), .Z(n_22960));
	notech_reg_set opc_reg_30(.CP(n_62243), .D(n_22966), .SD(1'b1), .Q(opc[
		30]));
	notech_mux2 i_9629(.S(n_27145), .A(opc[30]), .B(n_9857), .Z(n_22966));
	notech_reg_set opc_reg_31(.CP(n_62243), .D(n_22972), .SD(1'b1), .Q(opc[
		31]));
	notech_mux2 i_9637(.S(n_27145), .A(opc[31]), .B(n_9862), .Z(n_22972));
	notech_nand3 i_85048356(.A(n_146856196), .B(n_146756195), .C(n_147356201
		), .Z(n_147456202));
	notech_reg nZF_reg(.CP(n_62243), .D(n_22978), .CD(n_61113), .Q(nZF));
	notech_mux2 i_9645(.S(n_7432), .A(nZF), .B(n_7435), .Z(n_22978));
	notech_and3 i_84948357(.A(n_147156199), .B(n_147056198), .C(n_1367), .Z(n_147356201
		));
	notech_reg regs_reg_0_0(.CP(n_62243), .D(n_22984), .CD(n_61113), .Q(regs_0
		[0]));
	notech_mux2 i_9653(.S(n_27163), .A(regs_0[0]), .B(n_27147), .Z(n_22984)
		);
	notech_reg regs_reg_0_1(.CP(n_62243), .D(n_22990), .CD(n_61113), .Q(regs_0
		[1]));
	notech_mux2 i_9661(.S(n_27163), .A(regs_0[1]), .B(n_15780), .Z(n_22990)
		);
	notech_ao4 i_84348363(.A(n_54024), .B(n_28995), .C(n_321688474), .D(n_28994
		), .Z(n_147156199));
	notech_reg regs_reg_0_2(.CP(n_62243), .D(n_22999), .CD(n_61114), .Q(regs_0
		[2]));
	notech_mux2 i_9669(.S(n_27163), .A(regs_0[2]), .B(n_15786), .Z(n_22999)
		);
	notech_ao4 i_84648360(.A(n_271688739), .B(n_58951), .C(n_320088489), .D(n_27601
		), .Z(n_147056198));
	notech_reg regs_reg_0_3(.CP(n_62243), .D(n_23008), .CD(n_61113), .Q(regs_0
		[3]));
	notech_mux2 i_9677(.S(n_27163), .A(regs_0[3]), .B(n_15792), .Z(n_23008)
		);
	notech_reg regs_reg_0_4(.CP(n_62243), .D(n_23016), .CD(n_61113), .Q(regs_0
		[4]));
	notech_mux2 i_9685(.S(n_27163), .A(regs_0[4]), .B(n_27148), .Z(n_23016)
		);
	notech_ao4 i_84548361(.A(n_27554), .B(n_59163), .C(n_55314), .D(n_28996)
		, .Z(n_146856196));
	notech_reg regs_reg_0_5(.CP(n_62243), .D(n_23024), .CD(n_61112), .Q(regs_0
		[5]));
	notech_mux2 i_9693(.S(n_27163), .A(regs_0[5]), .B(n_27149), .Z(n_23024)
		);
	notech_ao4 i_84448362(.A(n_271588740), .B(n_56943), .C(n_59095), .D(n_55133
		), .Z(n_146756195));
	notech_reg regs_reg_0_6(.CP(n_62243), .D(n_23032), .CD(n_61112), .Q(regs_0
		[6]));
	notech_mux2 i_9701(.S(n_27163), .A(regs_0[6]), .B(n_27150), .Z(n_23032)
		);
	notech_reg regs_reg_0_7(.CP(n_62243), .D(n_23041), .CD(n_61112), .Q(regs_0
		[7]));
	notech_mux2 i_9709(.S(n_27163), .A(regs_0[7]), .B(n_15816), .Z(n_23041)
		);
	notech_reg regs_reg_0_8(.CP(n_62243), .D(n_23050), .CD(n_61112), .Q(regs_0
		[8]));
	notech_mux2 i_9717(.S(n_27163), .A(regs_0[8]), .B(n_15822), .Z(n_23050)
		);
	notech_ao4 i_68748506(.A(n_2702), .B(n_57329), .C(n_28977), .D(n_26450),
		 .Z(n_146456192));
	notech_reg regs_reg_0_9(.CP(n_62243), .D(n_23057), .CD(n_61112), .Q(regs_0
		[9]));
	notech_mux2 i_9725(.S(n_27163), .A(regs_0[9]), .B(n_15828), .Z(n_23057)
		);
	notech_and4 i_68648507(.A(n_146156189), .B(n_1351), .C(n_262736782), .D(n_1354
		), .Z(n_146356191));
	notech_reg regs_reg_0_10(.CP(n_62243), .D(n_23064), .CD(n_61113), .Q(regs_0
		[10]));
	notech_mux2 i_9733(.S(n_27163), .A(regs_0[10]), .B(n_15834), .Z(n_23064)
		);
	notech_reg regs_reg_0_11(.CP(n_62243), .D(n_23070), .CD(n_61113), .Q(regs_0
		[11]));
	notech_mux2 i_9741(.S(n_27163), .A(regs_0[11]), .B(n_15840), .Z(n_23070)
		);
	notech_ao4 i_68448509(.A(n_55073), .B(n_56892), .C(n_55072), .D(n_55249)
		, .Z(n_146156189));
	notech_reg regs_reg_0_12(.CP(n_62243), .D(n_23076), .CD(n_61113), .Q(regs_0
		[12]));
	notech_mux2 i_9749(.S(n_27163), .A(regs_0[12]), .B(n_15846), .Z(n_23076)
		);
	notech_reg regs_reg_0_13(.CP(n_62171), .D(n_23082), .CD(n_61113), .Q(regs_0
		[13]));
	notech_mux2 i_9757(.S(n_27163), .A(regs_0[13]), .B(n_15852), .Z(n_23082)
		);
	notech_reg regs_reg_0_14(.CP(n_62171), .D(n_23088), .CD(n_61101), .Q(regs_0
		[14]));
	notech_mux2 i_9765(.S(n_27163), .A(regs_0[14]), .B(n_15858), .Z(n_23088)
		);
	notech_reg regs_reg_0_15(.CP(n_62171), .D(n_23094), .CD(n_61090), .Q(regs_0
		[15]));
	notech_mux2 i_9773(.S(n_27163), .A(regs_0[15]), .B(n_15864), .Z(n_23094)
		);
	notech_reg regs_reg_0_16(.CP(n_62171), .D(n_23100), .CD(n_61090), .Q(regs_0
		[16]));
	notech_mux2 i_9781(.S(n_54158), .A(regs_0[16]), .B(n_15870), .Z(n_23100)
		);
	notech_ao4 i_36448810(.A(n_58487), .B(n_28049), .C(n_55952), .D(n_28988)
		, .Z(n_145756185));
	notech_reg regs_reg_0_17(.CP(n_62171), .D(n_23106), .CD(n_61088), .Q(regs_0
		[17]));
	notech_mux2 i_9789(.S(n_54158), .A(regs_0[17]), .B(n_15876), .Z(n_23106)
		);
	notech_ao4 i_36348811(.A(n_55972), .B(n_28017), .C(n_55992), .D(n_27983)
		, .Z(n_145656184));
	notech_reg regs_reg_0_18(.CP(n_62171), .D(n_23112), .CD(n_61090), .Q(regs_0
		[18]));
	notech_mux2 i_9797(.S(n_54158), .A(regs_0[18]), .B(n_27151), .Z(n_23112)
		);
	notech_and2 i_36748807(.A(n_145456182), .B(n_145356181), .Z(n_145556183)
		);
	notech_reg regs_reg_0_19(.CP(n_62171), .D(n_23118), .CD(n_61090), .Q(regs_0
		[19]));
	notech_mux2 i_9805(.S(n_54158), .A(regs_0[19]), .B(n_27152), .Z(n_23118)
		);
	notech_ao4 i_36248812(.A(n_56013), .B(n_27951), .C(n_56033), .D(n_27917)
		, .Z(n_145456182));
	notech_reg regs_reg_0_20(.CP(n_62171), .D(n_23124), .CD(n_61090), .Q(regs_0
		[20]));
	notech_mux2 i_9813(.S(n_54158), .A(regs_0[20]), .B(n_27153), .Z(n_23124)
		);
	notech_ao4 i_36148813(.A(n_56043), .B(n_27883), .C(n_55879), .D(n_27848)
		, .Z(n_145356181));
	notech_reg regs_reg_0_21(.CP(n_62171), .D(n_23130), .CD(n_61090), .Q(regs_0
		[21]));
	notech_mux2 i_9821(.S(n_54158), .A(regs_0[21]), .B(n_27154), .Z(n_23130)
		);
	notech_and4 i_37048805(.A(n_145056178), .B(n_144956177), .C(n_144756175)
		, .D(n_144656174), .Z(n_145256180));
	notech_reg regs_reg_0_22(.CP(n_62243), .D(n_23136), .CD(n_61090), .Q(regs_0
		[22]));
	notech_mux2 i_9829(.S(n_54158), .A(regs_0[22]), .B(n_27155), .Z(n_23136)
		);
	notech_reg regs_reg_0_23(.CP(n_62169), .D(n_23143), .CD(n_61090), .Q(regs_0
		[23]));
	notech_mux2 i_9837(.S(n_54158), .A(regs_0[23]), .B(n_27156), .Z(n_23143)
		);
	notech_ao4 i_36048814(.A(n_55940), .B(n_27816), .C(n_55888), .D(n_27784)
		, .Z(n_145056178));
	notech_reg regs_reg_0_24(.CP(n_62169), .D(n_23149), .CD(n_61088), .Q(regs_0
		[24]));
	notech_mux2 i_9845(.S(n_54158), .A(regs_0[24]), .B(n_27157), .Z(n_23149)
		);
	notech_ao4 i_35948815(.A(n_55910), .B(n_27745), .C(n_55924), .D(n_27400)
		, .Z(n_144956177));
	notech_reg regs_reg_0_25(.CP(n_62239), .D(n_23155), .CD(n_61088), .Q(regs_0
		[25]));
	notech_mux2 i_9853(.S(n_54158), .A(regs_0[25]), .B(n_27158), .Z(n_23155)
		);
	notech_reg regs_reg_0_26(.CP(n_62239), .D(n_23161), .CD(n_61088), .Q(regs_0
		[26]));
	notech_mux2 i_9861(.S(n_54158), .A(regs_0[26]), .B(n_27159), .Z(n_23161)
		);
	notech_ao4 i_35848816(.A(n_56092), .B(n_27713), .C(n_56130), .D(n_27679)
		, .Z(n_144756175));
	notech_reg regs_reg_0_27(.CP(n_62239), .D(n_23167), .CD(n_61088), .Q(regs_0
		[27]));
	notech_mux2 i_9869(.S(n_54158), .A(regs_0[27]), .B(n_27160), .Z(n_23167)
		);
	notech_ao4 i_35748817(.A(n_56144), .B(n_27636), .C(n_56386), .D(n_28989)
		, .Z(n_144656174));
	notech_reg regs_reg_0_28(.CP(n_62239), .D(n_23173), .CD(n_61088), .Q(regs_0
		[28]));
	notech_mux2 i_9877(.S(n_54158), .A(regs_0[28]), .B(n_27161), .Z(n_23173)
		);
	notech_reg regs_reg_0_29(.CP(n_62239), .D(n_23179), .CD(n_61088), .Q(regs_0
		[29]));
	notech_mux2 i_9885(.S(n_54158), .A(regs_0[29]), .B(n_27162), .Z(n_23179)
		);
	notech_reg regs_reg_0_30(.CP(n_62239), .D(n_23187), .CD(n_61088), .Q(regs_0
		[30]));
	notech_mux2 i_9893(.S(n_54158), .A(regs_0[30]), .B(n_15954), .Z(n_23187)
		);
	notech_reg regs_reg_0_31(.CP(n_62239), .D(n_23194), .CD(n_61088), .Q(regs_0
		[31]));
	notech_mux2 i_9901(.S(n_54158), .A(regs_0[31]), .B(n_15960), .Z(n_23194)
		);
	notech_ao4 i_30548863(.A(n_55934), .B(n_27817), .C(n_55924), .D(n_27401)
		, .Z(n_1443));
	notech_reg cr1_reg_0(.CP(n_62239), .D(n_23200), .CD(n_61088), .Q(nbus_14522
		[0]));
	notech_mux2 i_9909(.S(n_301186331), .A(opa[0]), .B(nbus_14522[0]), .Z(n_23200
		));
	notech_ao4 i_30448864(.A(n_58483), .B(n_28050), .C(n_56092), .D(n_27714)
		, .Z(n_1442));
	notech_reg cr1_reg_1(.CP(n_62239), .D(n_23206), .CD(n_61090), .Q(nbus_14522
		[1]));
	notech_mux2 i_9917(.S(n_301186331), .A(opa[1]), .B(nbus_14522[1]), .Z(n_23206
		));
	notech_and2 i_30948860(.A(n_1440), .B(n_1439), .Z(n_1441));
	notech_reg cr1_reg_2(.CP(n_62323), .D(n_23212), .CD(n_61091), .Q(nbus_14522
		[2]));
	notech_mux2 i_9926(.S(n_301186331), .A(opa[2]), .B(nbus_14522[2]), .Z(n_23212
		));
	notech_ao4 i_30248865(.A(n_56043), .B(n_27884), .C(n_56126), .D(n_27680)
		, .Z(n_1440));
	notech_reg cr1_reg_3(.CP(n_62323), .D(n_23218), .CD(n_61091), .Q(nbus_14522
		[3]));
	notech_mux2 i_9934(.S(n_301186331), .A(opa[3]), .B(nbus_14522[3]), .Z(n_23218
		));
	notech_ao4 i_30148866(.A(n_56033), .B(n_27918), .C(n_56382), .D(n_28991)
		, .Z(n_1439));
	notech_reg cr1_reg_4(.CP(n_62323), .D(n_23224), .CD(n_61091), .Q(nbus_14522
		[4]));
	notech_mux2 i_9942(.S(n_301186331), .A(opa[4]), .B(nbus_14522[4]), .Z(n_23224
		));
	notech_and4 i_31148858(.A(n_1436), .B(n_1435), .C(n_1433), .D(n_1432), .Z
		(n_1438));
	notech_reg cr1_reg_5(.CP(n_62323), .D(n_23230), .CD(n_61091), .Q(nbus_14522
		[5]));
	notech_mux2 i_9950(.S(n_301186331), .A(opa[5]), .B(nbus_14522[5]), .Z(n_23230
		));
	notech_reg cr1_reg_6(.CP(n_62323), .D(n_23237), .CD(n_61091), .Q(nbus_14522
		[6]));
	notech_mux2 i_9958(.S(n_301186331), .A(opa[6]), .B(nbus_14522[6]), .Z(n_23237
		));
	notech_ao4 i_30048867(.A(n_56009), .B(n_27952), .C(n_56139), .D(n_27638)
		, .Z(n_1436));
	notech_reg cr1_reg_7(.CP(n_62323), .D(n_23243), .CD(n_61092), .Q(nbus_14522
		[7]));
	notech_mux2 i_9966(.S(n_301186331), .A(opa[7]), .B(nbus_14522[7]), .Z(n_23243
		));
	notech_ao4 i_29948868(.A(n_55992), .B(n_27984), .C(n_55888), .D(n_27785)
		, .Z(n_1435));
	notech_reg cr1_reg_8(.CP(n_62323), .D(n_23249), .CD(n_61092), .Q(nbus_14522
		[8]));
	notech_mux2 i_9974(.S(n_301186331), .A(opa[8]), .B(nbus_14522[8]), .Z(n_23249
		));
	notech_reg cr1_reg_9(.CP(n_62323), .D(n_23255), .CD(n_61091), .Q(nbus_14522
		[9]));
	notech_mux2 i_9982(.S(n_301186331), .A(opa[9]), .B(nbus_14522[9]), .Z(n_23255
		));
	notech_ao4 i_29848869(.A(n_55972), .B(n_28018), .C(n_55879), .D(n_27849)
		, .Z(n_1433));
	notech_reg cr1_reg_10(.CP(n_62323), .D(n_23261), .CD(n_61092), .Q(nbus_14522
		[10]));
	notech_mux2 i_9990(.S(n_301186331), .A(opa[10]), .B(nbus_14522[10]), .Z(n_23261
		));
	notech_ao4 i_29748870(.A(n_55906), .B(n_27746), .C(n_55952), .D(n_28990)
		, .Z(n_1432));
	notech_reg cr1_reg_11(.CP(n_62323), .D(n_23267), .CD(n_61090), .Q(nbus_14522
		[11]));
	notech_mux2 i_9998(.S(n_301186331), .A(opa[11]), .B(nbus_14522[11]), .Z(n_23267
		));
	notech_reg cr1_reg_12(.CP(n_62323), .D(n_23273), .CD(n_61091), .Q(nbus_14522
		[12]));
	notech_mux2 i_10006(.S(n_301186331), .A(opa[12]), .B(nbus_14522[12]), .Z
		(n_23273));
	notech_reg cr1_reg_13(.CP(n_62323), .D(n_23279), .CD(n_61090), .Q(nbus_14522
		[13]));
	notech_mux2 i_10014(.S(n_301186331), .A(opa[13]), .B(nbus_14522[13]), .Z
		(n_23279));
	notech_reg cr1_reg_14(.CP(n_62323), .D(n_23285), .CD(n_61090), .Q(nbus_14522
		[14]));
	notech_mux2 i_10022(.S(n_301186331), .A(opa[14]), .B(nbus_14522[14]), .Z
		(n_23285));
	notech_ao4 i_26148905(.A(n_58483), .B(n_28048), .C(n_55952), .D(n_28993)
		, .Z(n_1428));
	notech_reg cr1_reg_15(.CP(n_62323), .D(n_23291), .CD(n_61091), .Q(nbus_14522
		[15]));
	notech_mux2 i_10030(.S(n_301186331), .A(opa[15]), .B(nbus_14522[15]), .Z
		(n_23291));
	notech_ao4 i_26048906(.A(n_55965), .B(n_28016), .C(n_55992), .D(n_27982)
		, .Z(n_1427));
	notech_reg cr1_reg_16(.CP(n_62323), .D(n_23297), .CD(n_61091), .Q(nbus_14522
		[16]));
	notech_mux2 i_10038(.S(n_53853), .A(opa[16]), .B(nbus_14522[16]), .Z(n_23297
		));
	notech_and2 i_26448902(.A(n_1425), .B(n_1424), .Z(n_1426));
	notech_reg cr1_reg_17(.CP(n_62323), .D(n_23303), .CD(n_61091), .Q(nbus_14522
		[17]));
	notech_mux2 i_10047(.S(n_53853), .A(opa[17]), .B(nbus_14522[17]), .Z(n_23303
		));
	notech_ao4 i_25948907(.A(n_56009), .B(n_27950), .C(n_56033), .D(n_27916)
		, .Z(n_1425));
	notech_reg cr1_reg_18(.CP(n_62323), .D(n_23309), .CD(n_61091), .Q(nbus_14522
		[18]));
	notech_mux2 i_10055(.S(n_53853), .A(opa[18]), .B(nbus_14522[18]), .Z(n_23309
		));
	notech_ao4 i_25848908(.A(n_56043), .B(n_27882), .C(n_55879), .D(n_27847)
		, .Z(n_1424));
	notech_reg cr1_reg_19(.CP(n_62323), .D(n_23315), .CD(n_61091), .Q(nbus_14522
		[19]));
	notech_mux2 i_10063(.S(n_53853), .A(opa[19]), .B(nbus_14522[19]), .Z(n_23315
		));
	notech_and4 i_26648900(.A(n_1421), .B(n_1420), .C(n_1418), .D(n_1417), .Z
		(n_1423));
	notech_reg cr1_reg_20(.CP(n_62239), .D(n_23321), .CD(n_61088), .Q(nbus_14522
		[20]));
	notech_mux2 i_10071(.S(n_53853), .A(opa[20]), .B(nbus_14522[20]), .Z(n_23321
		));
	notech_reg cr1_reg_21(.CP(n_62323), .D(n_23327), .CD(n_61085), .Q(nbus_14522
		[21]));
	notech_mux2 i_10079(.S(n_53853), .A(opa[21]), .B(nbus_14522[21]), .Z(n_23327
		));
	notech_ao4 i_25748909(.A(n_55934), .B(n_27815), .C(n_55888), .D(n_27783)
		, .Z(n_1421));
	notech_reg cr1_reg_22(.CP(n_62241), .D(n_23333), .CD(n_61086), .Q(nbus_14522
		[22]));
	notech_mux2 i_10087(.S(n_53853), .A(opa[22]), .B(nbus_14522[22]), .Z(n_23333
		));
	notech_ao4 i_25648910(.A(n_55906), .B(n_27744), .C(n_55924), .D(n_27399)
		, .Z(n_1420));
	notech_reg cr1_reg_23(.CP(n_62241), .D(n_23339), .CD(n_61085), .Q(nbus_14522
		[23]));
	notech_mux2 i_10095(.S(n_53853), .A(opa[23]), .B(nbus_14522[23]), .Z(n_23339
		));
	notech_reg cr1_reg_24(.CP(n_62241), .D(n_23345), .CD(n_61085), .Q(nbus_14522
		[24]));
	notech_mux2 i_10103(.S(n_53853), .A(opa[24]), .B(nbus_14522[24]), .Z(n_23345
		));
	notech_ao4 i_25548911(.A(n_56092), .B(n_27712), .C(n_56126), .D(n_27677)
		, .Z(n_1418));
	notech_reg cr1_reg_25(.CP(n_62241), .D(n_23351), .CD(n_61086), .Q(nbus_14522
		[25]));
	notech_mux2 i_10111(.S(n_53853), .A(opa[25]), .B(nbus_14522[25]), .Z(n_23351
		));
	notech_ao4 i_25448912(.A(n_56139), .B(n_27635), .C(n_56382), .D(n_28992)
		, .Z(n_1417));
	notech_reg cr1_reg_26(.CP(n_62241), .D(n_23359), .CD(n_61086), .Q(nbus_14522
		[26]));
	notech_mux2 i_10119(.S(n_53853), .A(opa[26]), .B(nbus_14522[26]), .Z(n_23359
		));
	notech_nor2 i_22948935(.A(n_2180), .B(n_60602), .Z(n_1416));
	notech_reg cr1_reg_27(.CP(n_62241), .D(n_23366), .CD(n_61086), .Q(nbus_14522
		[27]));
	notech_mux2 i_10127(.S(n_53853), .A(opa[27]), .B(nbus_14522[27]), .Z(n_23366
		));
	notech_reg cr1_reg_28(.CP(n_62241), .D(n_23374), .CD(n_61086), .Q(nbus_14522
		[28]));
	notech_mux2 i_10135(.S(n_53853), .A(opa[28]), .B(nbus_14522[28]), .Z(n_23374
		));
	notech_reg cr1_reg_29(.CP(n_62241), .D(n_23387), .CD(n_61086), .Q(nbus_14522
		[29]));
	notech_mux2 i_10143(.S(n_53853), .A(opa[29]), .B(nbus_14522[29]), .Z(n_23387
		));
	notech_ao4 i_11949043(.A(n_56255), .B(n_27817), .C(n_57371), .D(n_27401)
		, .Z(n_1413));
	notech_reg cr1_reg_30(.CP(n_62241), .D(n_23393), .CD(n_61085), .Q(nbus_14522
		[30]));
	notech_mux2 i_10151(.S(n_53853), .A(opa[30]), .B(nbus_14522[30]), .Z(n_23393
		));
	notech_ao4 i_11849044(.A(n_59219), .B(n_28050), .C(n_56265), .D(n_27714)
		, .Z(n_1412));
	notech_reg cr1_reg_31(.CP(n_62241), .D(n_23399), .CD(n_61085), .Q(nbus_14522
		[31]));
	notech_mux2 i_10159(.S(n_53853), .A(opa[31]), .B(nbus_14522[31]), .Z(n_23399
		));
	notech_and2 i_12249040(.A(n_1410), .B(n_1409), .Z(n_1411));
	notech_reg cr2_reg_reg_0(.CP(n_62241), .D(n_23405), .CD(n_61085), .Q(cr2_reg
		[0]));
	notech_mux2 i_10167(.S(\nbus_11274[0] ), .A(cr2_reg[0]), .B(n_7611), .Z(n_23405
		));
	notech_ao4 i_11749045(.A(n_56276), .B(n_27884), .C(n_56285), .D(n_27680)
		, .Z(n_1410));
	notech_reg cr2_reg_reg_1(.CP(n_62241), .D(n_23411), .CD(n_61085), .Q(cr2_reg
		[1]));
	notech_mux2 i_10175(.S(\nbus_11274[0] ), .A(cr2_reg[1]), .B(n_7617), .Z(n_23411
		));
	notech_ao4 i_11649046(.A(n_60479), .B(n_27918), .C(n_56395), .D(n_28991)
		, .Z(n_1409));
	notech_reg cr2_reg_reg_2(.CP(n_62241), .D(n_23417), .CD(n_61085), .Q(cr2_reg
		[2]));
	notech_mux2 i_10183(.S(\nbus_11274[0] ), .A(cr2_reg[2]), .B(n_7623), .Z(n_23417
		));
	notech_and4 i_12449038(.A(n_1406), .B(n_1405), .C(n_1403), .D(n_1402), .Z
		(n_1408));
	notech_reg cr2_reg_reg_3(.CP(n_62241), .D(n_23423), .CD(n_61085), .Q(cr2_reg
		[3]));
	notech_mux2 i_10191(.S(\nbus_11274[0] ), .A(cr2_reg[3]), .B(n_7629), .Z(n_23423
		));
	notech_reg cr2_reg_reg_4(.CP(n_62241), .D(n_23429), .CD(n_61085), .Q(cr2_reg
		[4]));
	notech_mux2 i_10199(.S(\nbus_11274[0] ), .A(cr2_reg[4]), .B(n_7635), .Z(n_23429
		));
	notech_ao4 i_11549047(.A(n_27952), .B(n_56296), .C(n_56305), .D(n_27638)
		, .Z(n_1406));
	notech_reg cr2_reg_reg_5(.CP(n_62241), .D(n_23435), .CD(n_61085), .Q(cr2_reg
		[5]));
	notech_mux2 i_10207(.S(\nbus_11274[0] ), .A(cr2_reg[5]), .B(n_7641), .Z(n_23435
		));
	notech_ao4 i_11449048(.A(n_56409), .B(n_27984), .C(n_57338), .D(n_27785)
		, .Z(n_1405));
	notech_reg cr2_reg_reg_6(.CP(n_62241), .D(n_23441), .CD(n_61085), .Q(cr2_reg
		[6]));
	notech_mux2 i_10215(.S(\nbus_11274[0] ), .A(cr2_reg[6]), .B(n_7647), .Z(n_23441
		));
	notech_reg cr2_reg_reg_7(.CP(n_62241), .D(n_23447), .CD(n_61086), .Q(cr2_reg
		[7]));
	notech_mux2 i_10223(.S(\nbus_11274[0] ), .A(cr2_reg[7]), .B(n_7653), .Z(n_23447
		));
	notech_ao4 i_11349049(.A(n_28018), .B(n_56226), .C(n_27849), .D(n_57358)
		, .Z(n_1403));
	notech_reg cr2_reg_reg_8(.CP(n_62241), .D(n_23453), .CD(n_61087), .Q(cr2_reg
		[8]));
	notech_mux2 i_10231(.S(\nbus_11274[0] ), .A(cr2_reg[8]), .B(n_7659), .Z(n_23453
		));
	notech_ao4 i_11249050(.A(n_56235), .B(n_27746), .C(n_28990), .D(n_56246)
		, .Z(n_1402));
	notech_reg cr2_reg_reg_9(.CP(n_62169), .D(n_23459), .CD(n_61087), .Q(cr2_reg
		[9]));
	notech_mux2 i_10239(.S(\nbus_11274[0] ), .A(cr2_reg[9]), .B(n_7665), .Z(n_23459
		));
	notech_reg cr2_reg_reg_10(.CP(n_62169), .D(n_23465), .CD(n_61087), .Q(cr2_reg
		[10]));
	notech_mux2 i_10247(.S(\nbus_11274[0] ), .A(cr2_reg[10]), .B(n_7671), .Z
		(n_23465));
	notech_reg cr2_reg_reg_11(.CP(n_62169), .D(n_23471), .CD(n_61087), .Q(cr2_reg
		[11]));
	notech_mux2 i_10255(.S(\nbus_11274[0] ), .A(cr2_reg[11]), .B(n_7677), .Z
		(n_23471));
	notech_ao4 i_8249080(.A(n_57371), .B(n_27400), .C(n_59219), .D(n_28049),
		 .Z(n_1399));
	notech_reg cr2_reg_reg_12(.CP(n_62169), .D(n_23477), .CD(n_61087), .Q(cr2_reg
		[12]));
	notech_mux2 i_10263(.S(\nbus_11274[0] ), .A(cr2_reg[12]), .B(n_7683), .Z
		(n_23477));
	notech_ao4 i_8149081(.A(n_56265), .B(n_27713), .C(n_56276), .D(n_27883),
		 .Z(n_1398));
	notech_reg cr2_reg_reg_13(.CP(n_62169), .D(n_23483), .CD(n_61087), .Q(cr2_reg
		[13]));
	notech_mux2 i_10271(.S(\nbus_11274[0] ), .A(cr2_reg[13]), .B(n_7689), .Z
		(n_23483));
	notech_and2 i_8549077(.A(n_1396), .B(n_1395), .Z(n_1397));
	notech_reg cr2_reg_reg_14(.CP(n_62169), .D(n_23489), .CD(n_61088), .Q(cr2_reg
		[14]));
	notech_mux2 i_10279(.S(\nbus_11274[0] ), .A(cr2_reg[14]), .B(n_7695), .Z
		(n_23489));
	notech_ao4 i_8049082(.A(n_56285), .B(n_27679), .C(n_60479), .D(n_27917),
		 .Z(n_1396));
	notech_reg cr2_reg_reg_15(.CP(n_62169), .D(n_23495), .CD(n_61087), .Q(cr2_reg
		[15]));
	notech_mux2 i_10287(.S(\nbus_11274[0] ), .A(cr2_reg[15]), .B(n_7701), .Z
		(n_23495));
	notech_ao4 i_7949083(.A(n_56395), .B(n_28989), .C(n_27951), .D(n_56296),
		 .Z(n_1395));
	notech_reg cr2_reg_reg_16(.CP(n_62169), .D(n_23501), .CD(n_61087), .Q(cr2_reg
		[16]));
	notech_mux2 i_10295(.S(\nbus_11274[0] ), .A(cr2_reg[16]), .B(n_7707), .Z
		(n_23501));
	notech_and4 i_8749075(.A(n_1392), .B(n_1391), .C(n_1389), .D(n_1388), .Z
		(n_1394));
	notech_reg cr2_reg_reg_17(.CP(n_62169), .D(n_23507), .CD(n_61086), .Q(cr2_reg
		[17]));
	notech_mux2 i_10303(.S(\nbus_11274[0] ), .A(cr2_reg[17]), .B(n_7713), .Z
		(n_23507));
	notech_reg cr2_reg_reg_18(.CP(n_62239), .D(n_23513), .CD(n_61086), .Q(cr2_reg
		[18]));
	notech_mux2 i_10311(.S(n_53864), .A(cr2_reg[18]), .B(n_7719), .Z(n_23513
		));
	notech_ao4 i_7849084(.A(n_56305), .B(n_27636), .C(n_56409), .D(n_27983),
		 .Z(n_1392));
	notech_reg cr2_reg_reg_19(.CP(n_62233), .D(n_23519), .CD(n_61086), .Q(cr2_reg
		[19]));
	notech_mux2 i_10319(.S(n_53864), .A(cr2_reg[19]), .B(n_7725), .Z(n_23519
		));
	notech_ao4 i_7749085(.A(n_57338), .B(n_27784), .C(n_28017), .D(n_56226),
		 .Z(n_1391));
	notech_reg cr2_reg_reg_20(.CP(n_62167), .D(n_23525), .CD(n_61086), .Q(cr2_reg
		[20]));
	notech_mux2 i_10327(.S(n_53864), .A(cr2_reg[20]), .B(n_7731), .Z(n_23525
		));
	notech_reg cr2_reg_reg_21(.CP(n_62233), .D(n_23531), .CD(n_61086), .Q(cr2_reg
		[21]));
	notech_mux2 i_10335(.S(n_53864), .A(cr2_reg[21]), .B(n_7737), .Z(n_23531
		));
	notech_ao4 i_7649086(.A(n_57358), .B(n_27848), .C(n_56255), .D(n_27816),
		 .Z(n_1389));
	notech_reg cr2_reg_reg_22(.CP(n_62233), .D(n_23537), .CD(n_61087), .Q(cr2_reg
		[22]));
	notech_mux2 i_10343(.S(n_53864), .A(cr2_reg[22]), .B(n_7743), .Z(n_23537
		));
	notech_ao4 i_7549087(.A(n_56235), .B(n_27745), .C(n_28988), .D(n_56246),
		 .Z(n_1388));
	notech_reg cr2_reg_reg_23(.CP(n_62233), .D(n_23543), .CD(n_61087), .Q(cr2_reg
		[23]));
	notech_mux2 i_10351(.S(n_53864), .A(cr2_reg[23]), .B(n_7749), .Z(n_23543
		));
	notech_reg cr2_reg_reg_24(.CP(n_62233), .D(n_23549), .CD(n_61087), .Q(cr2_reg
		[24]));
	notech_mux2 i_10359(.S(n_53864), .A(cr2_reg[24]), .B(n_7755), .Z(n_23549
		));
	notech_reg cr2_reg_reg_25(.CP(n_62233), .D(n_23555), .CD(n_61087), .Q(cr2_reg
		[25]));
	notech_mux2 i_10367(.S(n_53864), .A(cr2_reg[25]), .B(n_7761), .Z(n_23555
		));
	notech_and4 i_3121578(.A(n_1487), .B(n_1385), .C(n_82622813), .D(n_1384)
		, .Z(n_16530));
	notech_reg cr2_reg_reg_26(.CP(n_62233), .D(n_23561), .CD(n_61092), .Q(cr2_reg
		[26]));
	notech_mux2 i_10375(.S(n_53864), .A(cr2_reg[26]), .B(n_7767), .Z(n_23561
		));
	notech_or4 i_86948337(.A(n_182758113), .B(n_56265), .C(n_270988746), .D(n_1492
		), .Z(n_1385));
	notech_reg cr2_reg_reg_27(.CP(n_62233), .D(n_23567), .CD(n_61098), .Q(cr2_reg
		[27]));
	notech_mux2 i_10383(.S(n_53864), .A(cr2_reg[27]), .B(n_7773), .Z(n_23567
		));
	notech_or2 i_87248336(.A(n_271188744), .B(n_302821915), .Z(n_1384));
	notech_reg cr2_reg_reg_28(.CP(n_62233), .D(n_23573), .CD(n_61098), .Q(cr2_reg
		[28]));
	notech_mux2 i_10391(.S(n_53864), .A(cr2_reg[28]), .B(n_7779), .Z(n_23573
		));
	notech_or4 i_87348335(.A(n_320988480), .B(n_1492), .C(n_28081), .D(n_60504
		), .Z(n_1383));
	notech_reg cr2_reg_reg_29(.CP(n_62233), .D(n_23579), .CD(n_61098), .Q(cr2_reg
		[29]));
	notech_mux2 i_10400(.S(n_53864), .A(cr2_reg[29]), .B(n_7785), .Z(n_23579
		));
	notech_nand2 i_86848338(.A(sav_esi[30]), .B(n_60584), .Z(n_1382));
	notech_reg cr2_reg_reg_30(.CP(n_62319), .D(n_23585), .CD(n_61098), .Q(cr2_reg
		[30]));
	notech_mux2 i_10409(.S(n_53864), .A(cr2_reg[30]), .B(n_7791), .Z(n_23585
		));
	notech_reg cr2_reg_reg_31(.CP(n_62319), .D(n_23591), .CD(n_61098), .Q(cr2_reg
		[31]));
	notech_mux2 i_10417(.S(n_53864), .A(cr2_reg[31]), .B(n_7797), .Z(n_23591
		));
	notech_reg cr3_reg_0(.CP(n_62319), .D(n_23597), .CD(n_61098), .Q(\nbus_14521[0] 
		));
	notech_mux2 i_10425(.S(n_301086330), .A(opa[0]), .B(\nbus_14521[0] ), .Z
		(n_23597));
	notech_reg cr3_reg_1(.CP(n_62319), .D(n_23603), .CD(n_61098), .Q(\nbus_14521[1] 
		));
	notech_mux2 i_10433(.S(n_301086330), .A(opa[1]), .B(\nbus_14521[1] ), .Z
		(n_23603));
	notech_reg cr3_reg_2(.CP(n_62319), .D(n_23609), .CD(n_61098), .Q(\nbus_14521[2] 
		));
	notech_mux2 i_10441(.S(n_301086330), .A(opa[2]), .B(\nbus_14521[2] ), .Z
		(n_23609));
	notech_reg cr3_reg_3(.CP(n_62319), .D(n_23615), .CD(n_61098), .Q(\nbus_14521[3] 
		));
	notech_mux2 i_10449(.S(n_301086330), .A(opa[3]), .B(\nbus_14521[3] ), .Z
		(n_23615));
	notech_reg cr3_reg_4(.CP(n_62319), .D(n_23621), .CD(n_61097), .Q(\nbus_14521[4] 
		));
	notech_mux2 i_10457(.S(n_301086330), .A(opa[4]), .B(\nbus_14521[4] ), .Z
		(n_23621));
	notech_reg cr3_reg_5(.CP(n_62319), .D(n_23627), .CD(n_61097), .Q(\nbus_14521[5] 
		));
	notech_mux2 i_10465(.S(n_301086330), .A(opa[5]), .B(\nbus_14521[5] ), .Z
		(n_23627));
	notech_reg cr3_reg_6(.CP(n_62319), .D(n_23633), .CD(n_61097), .Q(\nbus_14521[6] 
		));
	notech_mux2 i_10473(.S(n_301086330), .A(opa[6]), .B(\nbus_14521[6] ), .Z
		(n_23633));
	notech_or4 i_85648350(.A(n_54520), .B(n_205788856), .C(n_60468), .D(n_56901
		), .Z(n_1373));
	notech_reg cr3_reg_7(.CP(n_62319), .D(n_23639), .CD(n_61097), .Q(\nbus_14521[7] 
		));
	notech_mux2 i_10481(.S(n_301086330), .A(opa[7]), .B(\nbus_14521[7] ), .Z
		(n_23639));
	notech_reg cr3_reg_8(.CP(n_62319), .D(n_23645), .CD(n_61097), .Q(\nbus_14521[8] 
		));
	notech_mux2 i_10489(.S(n_301086330), .A(opa[8]), .B(\nbus_14521[8] ), .Z
		(n_23645));
	notech_reg cr3_reg_9(.CP(n_62319), .D(n_23651), .CD(n_61098), .Q(\nbus_14521[9] 
		));
	notech_mux2 i_10497(.S(n_301086330), .A(opa[9]), .B(\nbus_14521[9] ), .Z
		(n_23651));
	notech_nao3 i_85748349(.A(n_26506), .B(n_56538), .C(n_270988746), .Z(n_1370
		));
	notech_reg cr3_reg_10(.CP(n_62319), .D(n_23657), .CD(n_61098), .Q(\nbus_14521[10] 
		));
	notech_mux2 i_10505(.S(n_301086330), .A(opa[10]), .B(\nbus_14521[10] ), 
		.Z(n_23657));
	notech_or4 i_3221579(.A(n_1368), .B(n_147456202), .C(n_1369), .D(n_1358)
		, .Z(n_16536));
	notech_reg cr3_reg_11(.CP(n_62319), .D(n_23663), .CD(n_61097), .Q(\nbus_14521[11] 
		));
	notech_mux2 i_10513(.S(n_301086330), .A(opa[11]), .B(\nbus_14521[11] ), 
		.Z(n_23663));
	notech_nor2 i_84148365(.A(n_271288743), .B(n_302821915), .Z(n_1369));
	notech_reg cr3_reg_12(.CP(n_62319), .D(n_23669), .CD(n_61098), .Q(cr3[12
		]));
	notech_mux2 i_10521(.S(n_301086330), .A(opa[12]), .B(cr3[12]), .Z(n_23669
		));
	notech_ao3 i_84248364(.A(opc_10[31]), .B(n_62405), .C(n_302321910), .Z(n_1368
		));
	notech_reg cr3_reg_13(.CP(n_62319), .D(n_23675), .CD(n_61099), .Q(cr3[13
		]));
	notech_mux2 i_10529(.S(n_301086330), .A(opa[13]), .B(cr3[13]), .Z(n_23675
		));
	notech_nand2 i_83948367(.A(sav_esi[31]), .B(n_60584), .Z(n_1367));
	notech_reg cr3_reg_14(.CP(n_62319), .D(n_23681), .CD(n_61101), .Q(cr3[14
		]));
	notech_mux2 i_10537(.S(n_301086330), .A(opa[14]), .B(cr3[14]), .Z(n_23681
		));
	notech_reg cr3_reg_15(.CP(n_62319), .D(n_23687), .CD(n_61101), .Q(cr3[15
		]));
	notech_mux2 i_10545(.S(n_301086330), .A(opa[15]), .B(cr3[15]), .Z(n_23687
		));
	notech_reg cr3_reg_16(.CP(n_62319), .D(n_23693), .CD(n_61099), .Q(cr3[16
		]));
	notech_mux2 i_10553(.S(n_55214), .A(opa[16]), .B(cr3[16]), .Z(n_23693)
		);
	notech_reg cr3_reg_17(.CP(n_62373), .D(n_23699), .CD(n_61099), .Q(cr3[17
		]));
	notech_mux2 i_10561(.S(n_55214), .A(opa[17]), .B(cr3[17]), .Z(n_23699)
		);
	notech_reg cr3_reg_18(.CP(n_62317), .D(n_23705), .CD(n_61101), .Q(cr3[18
		]));
	notech_mux2 i_10569(.S(n_55214), .A(opa[18]), .B(cr3[18]), .Z(n_23705)
		);
	notech_reg cr3_reg_19(.CP(n_62373), .D(n_23711), .CD(n_61101), .Q(cr3[19
		]));
	notech_mux2 i_10577(.S(n_55214), .A(opa[19]), .B(cr3[19]), .Z(n_23711)
		);
	notech_reg cr3_reg_20(.CP(n_62373), .D(n_23717), .CD(n_61101), .Q(cr3[20
		]));
	notech_mux2 i_10585(.S(n_55214), .A(opa[20]), .B(cr3[20]), .Z(n_23717)
		);
	notech_reg cr3_reg_21(.CP(n_62373), .D(n_23723), .CD(n_61101), .Q(cr3[21
		]));
	notech_mux2 i_10593(.S(n_55214), .A(opa[21]), .B(cr3[21]), .Z(n_23723)
		);
	notech_reg cr3_reg_22(.CP(n_62373), .D(n_23729), .CD(n_61101), .Q(cr3[22
		]));
	notech_mux2 i_10601(.S(n_55214), .A(opa[22]), .B(cr3[22]), .Z(n_23729)
		);
	notech_nor2 i_84048366(.A(n_55313), .B(n_271088745), .Z(n_1358));
	notech_reg cr3_reg_23(.CP(n_62373), .D(n_23735), .CD(n_61099), .Q(cr3[23
		]));
	notech_mux2 i_10609(.S(n_55214), .A(opa[23]), .B(cr3[23]), .Z(n_23735)
		);
	notech_and4 i_3021065(.A(n_146456192), .B(n_146356191), .C(n_1357), .D(n_1350
		), .Z(n_13989));
	notech_reg cr3_reg_24(.CP(n_62373), .D(n_23741), .CD(n_61099), .Q(cr3[24
		]));
	notech_mux2 i_10617(.S(n_55214), .A(opa[24]), .B(cr3[24]), .Z(n_23741)
		);
	notech_nao3 i_68148511(.A(opc_10[29]), .B(n_62405), .C(n_123623223), .Z(n_1357
		));
	notech_reg cr3_reg_25(.CP(n_62373), .D(n_23747), .CD(n_61099), .Q(cr3[25
		]));
	notech_mux2 i_10625(.S(n_55214), .A(opa[25]), .B(cr3[25]), .Z(n_23747)
		);
	notech_reg cr3_reg_26(.CP(n_62373), .D(n_23753), .CD(n_61099), .Q(cr3[26
		]));
	notech_mux2 i_10633(.S(n_55214), .A(opa[26]), .B(cr3[26]), .Z(n_23753)
		);
	notech_reg cr3_reg_27(.CP(n_62373), .D(n_23761), .CD(n_61099), .Q(cr3[27
		]));
	notech_mux2 i_10641(.S(n_55214), .A(opa[27]), .B(cr3[27]), .Z(n_23761)
		);
	notech_or2 i_68048512(.A(n_123423221), .B(n_59104), .Z(n_1354));
	notech_reg cr3_reg_28(.CP(n_62373), .D(n_23767), .CD(n_61099), .Q(cr3[28
		]));
	notech_mux2 i_10649(.S(n_55214), .A(opa[28]), .B(cr3[28]), .Z(n_23767)
		);
	notech_reg cr3_reg_29(.CP(n_62373), .D(n_23773), .CD(n_61099), .Q(cr3[29
		]));
	notech_mux2 i_10657(.S(n_55214), .A(opa[29]), .B(cr3[29]), .Z(n_23773)
		);
	notech_reg cr3_reg_30(.CP(n_62373), .D(n_23779), .CD(n_61099), .Q(cr3[30
		]));
	notech_mux2 i_10665(.S(n_55214), .A(opa[30]), .B(cr3[30]), .Z(n_23779)
		);
	notech_or4 i_67448518(.A(n_59263), .B(n_59272), .C(n_56172), .D(n_262936784
		), .Z(n_1351));
	notech_reg cr3_reg_31(.CP(n_62373), .D(n_23785), .CD(n_61099), .Q(cr3[31
		]));
	notech_mux2 i_10673(.S(n_55214), .A(opa[31]), .B(cr3[31]), .Z(n_23785)
		);
	notech_or4 i_67948513(.A(n_56177), .B(n_58660), .C(n_55798), .D(n_270688747
		), .Z(n_1350));
	notech_reg opa_reg_0(.CP(n_62373), .D(n_23791), .CD(n_61097), .Q(opa[0])
		);
	notech_mux2 i_10681(.S(n_27249), .A(opa[0]), .B(n_27239), .Z(n_23791));
	notech_reg opa_reg_1(.CP(n_62373), .D(n_23797), .CD(n_61093), .Q(opa[1])
		);
	notech_mux2 i_10689(.S(n_27249), .A(opa[1]), .B(n_27240), .Z(n_23797));
	notech_reg opa_reg_2(.CP(n_62373), .D(n_23803), .CD(n_61093), .Q(opa[2])
		);
	notech_mux2 i_10697(.S(n_27249), .A(opa[2]), .B(n_27241), .Z(n_23803));
	notech_reg opa_reg_3(.CP(n_62373), .D(n_23809), .CD(n_61093), .Q(opa[3])
		);
	notech_mux2 i_10705(.S(n_27249), .A(opa[3]), .B(n_27242), .Z(n_23809));
	notech_reg opa_reg_4(.CP(n_62373), .D(n_23815), .CD(n_61093), .Q(opa[4])
		);
	notech_mux2 i_10713(.S(n_27249), .A(opa[4]), .B(n_27243), .Z(n_23815));
	notech_reg opa_reg_5(.CP(n_62317), .D(n_23821), .CD(n_61093), .Q(opa[5])
		);
	notech_mux2 i_10721(.S(n_27249), .A(opa[5]), .B(n_27244), .Z(n_23821));
	notech_reg opa_reg_6(.CP(n_62317), .D(n_23827), .CD(n_61093), .Q(opa[6])
		);
	notech_mux2 i_10732(.S(n_27249), .A(opa[6]), .B(n_27245), .Z(n_23827));
	notech_reg opa_reg_7(.CP(n_62317), .D(n_23833), .CD(n_61093), .Q(opa[7])
		);
	notech_mux2 i_10740(.S(n_27249), .A(opa[7]), .B(n_27248), .Z(n_23833));
	notech_reg opa_reg_8(.CP(n_62317), .D(n_23839), .CD(n_61093), .Q(opa[8])
		);
	notech_mux2 i_10748(.S(n_27257), .A(opa[8]), .B(n_27250), .Z(n_23839));
	notech_reg opa_reg_9(.CP(n_62317), .D(n_23845), .CD(n_61093), .Q(opa[9])
		);
	notech_mux2 i_10756(.S(n_27257), .A(opa[9]), .B(n_27251), .Z(n_23845));
	notech_reg opa_reg_10(.CP(n_62317), .D(n_23851), .CD(n_61092), .Q(opa[10
		]));
	notech_mux2 i_10764(.S(n_27257), .A(opa[10]), .B(n_27252), .Z(n_23851)
		);
	notech_reg opa_reg_11(.CP(n_62317), .D(n_23857), .CD(n_61092), .Q(opa[11
		]));
	notech_mux2 i_10772(.S(n_27257), .A(opa[11]), .B(n_27253), .Z(n_23857)
		);
	notech_reg opa_reg_12(.CP(n_62317), .D(n_23863), .CD(n_61092), .Q(opa[12
		]));
	notech_mux2 i_10780(.S(n_27257), .A(opa[12]), .B(n_27254), .Z(n_23863)
		);
	notech_reg opa_reg_13(.CP(n_62317), .D(n_23869), .CD(n_61092), .Q(opa[13
		]));
	notech_mux2 i_10788(.S(n_27257), .A(opa[13]), .B(n_17274), .Z(n_23869)
		);
	notech_reg opa_reg_14(.CP(n_62317), .D(n_23875), .CD(n_61092), .Q(opa[14
		]));
	notech_mux2 i_10796(.S(n_27257), .A(opa[14]), .B(n_27255), .Z(n_23875)
		);
	notech_reg opa_reg_15(.CP(n_62233), .D(n_23881), .CD(n_61092), .Q(opa[15
		]));
	notech_mux2 i_10804(.S(n_27257), .A(opa[15]), .B(n_27256), .Z(n_23881)
		);
	notech_reg opa_reg_16(.CP(n_62167), .D(n_23887), .CD(n_61093), .Q(opa[16
		]));
	notech_mux2 i_10812(.S(n_27258), .A(opa[16]), .B(n_17292), .Z(n_23887)
		);
	notech_reg opa_reg_17(.CP(n_62321), .D(n_23893), .CD(n_61092), .Q(opa[17
		]));
	notech_mux2 i_10820(.S(n_27258), .A(opa[17]), .B(n_17298), .Z(n_23893)
		);
	notech_reg opa_reg_18(.CP(n_62235), .D(n_23899), .CD(n_61092), .Q(opa[18
		]));
	notech_mux2 i_10828(.S(n_27258), .A(opa[18]), .B(n_17304), .Z(n_23899)
		);
	notech_reg opa_reg_19(.CP(n_62235), .D(n_23905), .CD(n_61093), .Q(opa[19
		]));
	notech_mux2 i_10836(.S(n_27258), .A(opa[19]), .B(n_17310), .Z(n_23905)
		);
	notech_reg opa_reg_20(.CP(n_62235), .D(n_23911), .CD(n_61096), .Q(opa[20
		]));
	notech_mux2 i_10844(.S(n_27258), .A(opa[20]), .B(n_17316), .Z(n_23911)
		);
	notech_reg opa_reg_21(.CP(n_62235), .D(n_23917), .CD(n_61096), .Q(opa[21
		]));
	notech_mux2 i_10852(.S(n_27258), .A(opa[21]), .B(n_17322), .Z(n_23917)
		);
	notech_reg opa_reg_22(.CP(n_62235), .D(n_23923), .CD(n_61096), .Q(opa[22
		]));
	notech_mux2 i_10860(.S(n_27258), .A(opa[22]), .B(n_17328), .Z(n_23923)
		);
	notech_reg opa_reg_23(.CP(n_62235), .D(n_23929), .CD(n_61096), .Q(opa[23
		]));
	notech_mux2 i_10868(.S(n_27258), .A(opa[23]), .B(n_17334), .Z(n_23929)
		);
	notech_reg opa_reg_24(.CP(n_62235), .D(n_23935), .CD(n_61097), .Q(opa[24
		]));
	notech_mux2 i_10876(.S(n_27258), .A(opa[24]), .B(n_17340), .Z(n_23935)
		);
	notech_reg opa_reg_25(.CP(n_62235), .D(n_23941), .CD(n_61097), .Q(opa[25
		]));
	notech_mux2 i_10884(.S(n_27258), .A(opa[25]), .B(n_17346), .Z(n_23941)
		);
	notech_reg opa_reg_26(.CP(n_62235), .D(n_23949), .CD(n_61097), .Q(opa[26
		]));
	notech_mux2 i_10892(.S(n_27258), .A(opa[26]), .B(n_17352), .Z(n_23949)
		);
	notech_reg opa_reg_27(.CP(n_62321), .D(n_23955), .CD(n_61097), .Q(opa[27
		]));
	notech_mux2 i_10900(.S(n_27258), .A(opa[27]), .B(n_17358), .Z(n_23955)
		);
	notech_reg opa_reg_28(.CP(n_62321), .D(n_23961), .CD(n_61097), .Q(opa[28
		]));
	notech_mux2 i_10908(.S(n_27258), .A(opa[28]), .B(n_17364), .Z(n_23961)
		);
	notech_reg opa_reg_29(.CP(n_62321), .D(n_23967), .CD(n_61096), .Q(opa[29
		]));
	notech_mux2 i_10916(.S(n_27258), .A(opa[29]), .B(n_17370), .Z(n_23967)
		);
	notech_reg opa_reg_30(.CP(n_62321), .D(n_23974), .CD(n_61096), .Q(opa[30
		]));
	notech_mux2 i_10924(.S(n_27258), .A(opa[30]), .B(n_17376), .Z(n_23974)
		);
	notech_reg opa_reg_31(.CP(n_62321), .D(n_23980), .CD(n_61093), .Q(opa[31
		]));
	notech_mux2 i_10932(.S(n_27258), .A(opa[31]), .B(n_17382), .Z(n_23980)
		);
	notech_reg tcmp_reg(.CP(n_62321), .D(n_23986), .CD(n_61096), .Q(tcmp));
	notech_mux2 i_10940(.S(n_27259), .A(n_59141), .B(n_251285832), .Z(n_23986
		));
	notech_reg sema_rw_reg(.CP(n_62321), .D(n_23992), .CD(n_61096), .Q(sema_rw
		));
	notech_mux2 i_10948(.S(n_27261), .A(sema_rw), .B(n_26473), .Z(n_23992)
		);
	notech_reg_set fsm_reg_0(.CP(n_62321), .D(n_23998), .SD(n_61096), .Q(fsm
		[0]));
	notech_mux2 i_10956(.S(\nbus_11321[0] ), .A(n_60735), .B(n_14896), .Z(n_23998
		));
	notech_reg_set fsm_reg_1(.CP(n_62321), .D(n_24004), .SD(n_61096), .Q(fsm
		[1]));
	notech_mux2 i_10965(.S(\nbus_11321[0] ), .A(fsm[1]), .B(n_14902), .Z(n_24004
		));
	notech_reg_set fsm_reg_2(.CP(n_62321), .D(n_24010), .SD(n_61096), .Q(fsm
		[2]));
	notech_mux2 i_10973(.S(\nbus_11321[0] ), .A(fsm[2]), .B(n_27263), .Z(n_24010
		));
	notech_reg_set fsm_reg_3(.CP(n_62321), .D(n_24016), .SD(n_61096), .Q(fsm
		[3]));
	notech_mux2 i_10981(.S(\nbus_11321[0] ), .A(n_60748), .B(n_14914), .Z(n_24016
		));
	notech_reg fsm_reg_4(.CP(n_62321), .D(n_24022), .CD(n_61142), .Q(fsm[4])
		);
	notech_mux2 i_10989(.S(\nbus_11321[0] ), .A(fsm[4]), .B(n_14920), .Z(n_24022
		));
	notech_reg vliw_pc_reg_0(.CP(n_62321), .D(n_24028), .CD(n_61142), .Q(vliw_pc
		[0]));
	notech_mux2 i_10998(.S(\nbus_11283[0] ), .A(vliw_pc[0]), .B(n_9296), .Z(n_24028
		));
	notech_reg vliw_pc_reg_1(.CP(n_62321), .D(n_24034), .CD(n_61142), .Q(vliw_pc
		[1]));
	notech_mux2 i_11008(.S(\nbus_11283[0] ), .A(vliw_pc[1]), .B(n_281486134)
		, .Z(n_24034));
	notech_reg vliw_pc_reg_2(.CP(n_62321), .D(n_24040), .CD(n_61142), .Q(vliw_pc
		[2]));
	notech_mux2 i_11016(.S(\nbus_11283[0] ), .A(vliw_pc[2]), .B(n_281586135)
		, .Z(n_24040));
	notech_reg vliw_pc_reg_3(.CP(n_62321), .D(n_24046), .CD(n_61142), .Q(vliw_pc
		[3]));
	notech_mux2 i_11024(.S(\nbus_11283[0] ), .A(vliw_pc[3]), .B(n_281686136)
		, .Z(n_24046));
	notech_reg vliw_pc_reg_4(.CP(n_62321), .D(n_24052), .CD(n_61142), .Q(vliw_pc
		[4]));
	notech_mux2 i_11032(.S(\nbus_11283[0] ), .A(vliw_pc[4]), .B(n_281786137)
		, .Z(n_24052));
	notech_reg io_add_reg_0(.CP(n_62321), .D(n_24058), .CD(n_61142), .Q(io_add
		[0]));
	notech_mux2 i_11040(.S(\nbus_11356[0] ), .A(io_add[0]), .B(n_322388467),
		 .Z(n_24058));
	notech_reg io_add_reg_1(.CP(n_62235), .D(n_24064), .CD(n_61142), .Q(io_add
		[1]));
	notech_mux2 i_11048(.S(\nbus_11356[0] ), .A(io_add[1]), .B(n_26493), .Z(n_24064
		));
	notech_reg io_add_reg_2(.CP(n_62235), .D(n_24070), .CD(n_61142), .Q(io_add
		[2]));
	notech_mux2 i_11056(.S(\nbus_11356[0] ), .A(io_add[2]), .B(n_185488093),
		 .Z(n_24070));
	notech_reg io_add_reg_3(.CP(n_62237), .D(n_24076), .CD(n_61141), .Q(io_add
		[3]));
	notech_mux2 i_11064(.S(\nbus_11356[0] ), .A(io_add[3]), .B(n_185588094),
		 .Z(n_24076));
	notech_reg io_add_reg_4(.CP(n_62237), .D(n_24084), .CD(n_61141), .Q(io_add
		[4]));
	notech_mux2 i_11072(.S(\nbus_11356[0] ), .A(io_add[4]), .B(n_365988136),
		 .Z(n_24084));
	notech_nor2 i_23548929(.A(n_318931576), .B(n_26277), .Z(n_1301));
	notech_reg io_add_reg_5(.CP(n_62237), .D(n_24090), .CD(n_61141), .Q(io_add
		[5]));
	notech_mux2 i_11080(.S(\nbus_11356[0] ), .A(io_add[5]), .B(n_185688095),
		 .Z(n_24090));
	notech_reg io_add_reg_6(.CP(n_62237), .D(n_24096), .CD(n_61141), .Q(io_add
		[6]));
	notech_mux2 i_11088(.S(\nbus_11356[0] ), .A(io_add[6]), .B(n_185788096),
		 .Z(n_24096));
	notech_reg io_add_reg_7(.CP(n_62237), .D(n_24102), .CD(n_61141), .Q(io_add
		[7]));
	notech_mux2 i_11096(.S(\nbus_11356[0] ), .A(io_add[7]), .B(n_185888097),
		 .Z(n_24102));
	notech_reg io_add_reg_8(.CP(n_62237), .D(n_24108), .CD(n_61142), .Q(io_add
		[8]));
	notech_mux2 i_11104(.S(\nbus_11356[0] ), .A(io_add[8]), .B(n_185988098),
		 .Z(n_24108));
	notech_reg io_add_reg_9(.CP(n_62237), .D(n_24114), .CD(n_61142), .Q(io_add
		[9]));
	notech_mux2 i_11112(.S(\nbus_11356[0] ), .A(io_add[9]), .B(n_186088099),
		 .Z(n_24114));
	notech_reg io_add_reg_10(.CP(n_62237), .D(n_24120), .CD(n_61142), .Q(io_add
		[10]));
	notech_mux2 i_11120(.S(\nbus_11356[0] ), .A(io_add[10]), .B(n_186188100)
		, .Z(n_24120));
	notech_reg io_add_reg_11(.CP(n_62237), .D(n_24126), .CD(n_61142), .Q(io_add
		[11]));
	notech_mux2 i_11128(.S(\nbus_11356[0] ), .A(io_add[11]), .B(n_186288101)
		, .Z(n_24126));
	notech_reg io_add_reg_12(.CP(n_62237), .D(n_24132), .CD(n_61143), .Q(io_add
		[12]));
	notech_mux2 i_11136(.S(\nbus_11356[0] ), .A(io_add[12]), .B(n_186388102)
		, .Z(n_24132));
	notech_reg io_add_reg_13(.CP(n_62237), .D(n_24138), .CD(n_61143), .Q(io_add
		[13]));
	notech_mux2 i_11144(.S(\nbus_11356[0] ), .A(io_add[13]), .B(n_186488103)
		, .Z(n_24138));
	notech_reg io_add_reg_14(.CP(n_62237), .D(n_24144), .CD(n_61144), .Q(io_add
		[14]));
	notech_mux2 i_11152(.S(\nbus_11356[0] ), .A(io_add[14]), .B(n_186588104)
		, .Z(n_24144));
	notech_reg io_add_reg_15(.CP(n_62237), .D(n_24150), .CD(n_61143), .Q(io_add
		[15]));
	notech_mux2 i_11160(.S(\nbus_11356[0] ), .A(io_add[15]), .B(n_186688105)
		, .Z(n_24150));
	notech_reg ldtr_reg_0(.CP(n_62237), .D(n_24156), .CD(n_61143), .Q(ldtr[0
		]));
	notech_mux2 i_11168(.S(n_299986319), .A(opb[0]), .B(ldtr[0]), .Z(n_24156
		));
	notech_reg ldtr_reg_1(.CP(n_62237), .D(n_24166), .CD(n_61144), .Q(ldtr[1
		]));
	notech_mux2 i_11177(.S(n_299986319), .A(opb[1]), .B(ldtr[1]), .Z(n_24166
		));
	notech_reg ldtr_reg_2(.CP(n_62237), .D(n_24173), .CD(n_61144), .Q(ldtr[2
		]));
	notech_mux2 i_11185(.S(n_299986319), .A(opb[2]), .B(ldtr[2]), .Z(n_24173
		));
	notech_reg ldtr_reg_3(.CP(n_62237), .D(n_24179), .CD(n_61144), .Q(ldtr[3
		]));
	notech_mux2 i_11193(.S(n_299986319), .A(opb[3]), .B(ldtr[3]), .Z(n_24179
		));
	notech_reg ldtr_reg_4(.CP(n_62237), .D(n_24185), .CD(n_61144), .Q(ldtr[4
		]));
	notech_mux2 i_11201(.S(n_299986319), .A(opb[4]), .B(ldtr[4]), .Z(n_24185
		));
	notech_reg ldtr_reg_5(.CP(n_62237), .D(n_24191), .CD(n_61144), .Q(ldtr[5
		]));
	notech_mux2 i_11210(.S(n_299986319), .A(opb[5]), .B(ldtr[5]), .Z(n_24191
		));
	notech_reg ldtr_reg_6(.CP(n_62167), .D(n_24197), .CD(n_61143), .Q(ldtr[6
		]));
	notech_mux2 i_11218(.S(n_299986319), .A(opb[6]), .B(ldtr[6]), .Z(n_24197
		));
	notech_reg ldtr_reg_7(.CP(n_62167), .D(n_24203), .CD(n_61143), .Q(ldtr[7
		]));
	notech_mux2 i_11226(.S(n_299986319), .A(opb[7]), .B(ldtr[7]), .Z(n_24203
		));
	notech_reg ldtr_reg_8(.CP(n_62167), .D(n_24209), .CD(n_61143), .Q(ldtr[8
		]));
	notech_mux2 i_11234(.S(n_299986319), .A(opb[8]), .B(ldtr[8]), .Z(n_24209
		));
	notech_reg ldtr_reg_9(.CP(n_62167), .D(n_24215), .CD(n_61143), .Q(ldtr[9
		]));
	notech_mux2 i_11243(.S(n_299986319), .A(opb[9]), .B(ldtr[9]), .Z(n_24215
		));
	notech_reg ldtr_reg_10(.CP(n_62167), .D(n_24221), .CD(n_61143), .Q(ldtr[
		10]));
	notech_mux2 i_11251(.S(n_299986319), .A(opb[10]), .B(ldtr[10]), .Z(n_24221
		));
	notech_reg ldtr_reg_11(.CP(n_62167), .D(n_24227), .CD(n_61143), .Q(ldtr[
		11]));
	notech_mux2 i_11259(.S(n_299986319), .A(opb[11]), .B(ldtr[11]), .Z(n_24227
		));
	notech_reg ldtr_reg_12(.CP(n_62167), .D(n_24233), .CD(n_61143), .Q(ldtr[
		12]));
	notech_mux2 i_11267(.S(n_299986319), .A(opb[12]), .B(ldtr[12]), .Z(n_24233
		));
	notech_reg ldtr_reg_13(.CP(n_62167), .D(n_24239), .CD(n_61143), .Q(ldtr[
		13]));
	notech_mux2 i_11275(.S(n_299986319), .A(opb[13]), .B(ldtr[13]), .Z(n_24239
		));
	notech_reg ldtr_reg_14(.CP(n_62167), .D(n_24245), .CD(n_61143), .Q(ldtr[
		14]));
	notech_mux2 i_11283(.S(n_299986319), .A(opb[14]), .B(ldtr[14]), .Z(n_24245
		));
	notech_reg ldtr_reg_15(.CP(n_62317), .D(n_24251), .CD(n_61141), .Q(ldtr[
		15]));
	notech_mux2 i_11291(.S(n_299986319), .A(opb[15]), .B(ldtr[15]), .Z(n_24251
		));
	notech_reg ldtr_reg_16(.CP(n_62225), .D(n_24257), .CD(n_61137), .Q(ldtr[
		16]));
	notech_mux2 i_11300(.S(n_53557), .A(opb[16]), .B(ldtr[16]), .Z(n_24257)
		);
	notech_reg ldtr_reg_17(.CP(n_62165), .D(n_24263), .CD(n_61137), .Q(ldtr[
		17]));
	notech_mux2 i_11308(.S(n_53557), .A(opb[17]), .B(ldtr[17]), .Z(n_24263)
		);
	notech_reg ldtr_reg_18(.CP(n_62225), .D(n_24269), .CD(n_61137), .Q(ldtr[
		18]));
	notech_mux2 i_11316(.S(n_53557), .A(opb[18]), .B(ldtr[18]), .Z(n_24269)
		);
	notech_reg ldtr_reg_19(.CP(n_62225), .D(n_24275), .CD(n_61137), .Q(ldtr[
		19]));
	notech_mux2 i_11324(.S(n_53557), .A(opb[19]), .B(ldtr[19]), .Z(n_24275)
		);
	notech_reg ldtr_reg_20(.CP(n_62225), .D(n_24281), .CD(n_61137), .Q(ldtr[
		20]));
	notech_mux2 i_11332(.S(n_53557), .A(opb[20]), .B(ldtr[20]), .Z(n_24281)
		);
	notech_reg ldtr_reg_21(.CP(n_62225), .D(n_24287), .CD(n_61137), .Q(ldtr[
		21]));
	notech_mux2 i_11340(.S(n_53557), .A(opb[21]), .B(ldtr[21]), .Z(n_24287)
		);
	notech_reg ldtr_reg_22(.CP(n_62225), .D(n_24295), .CD(n_61138), .Q(ldtr[
		22]));
	notech_mux2 i_11348(.S(n_53557), .A(opb[22]), .B(ldtr[22]), .Z(n_24295)
		);
	notech_reg ldtr_reg_23(.CP(n_62225), .D(n_24301), .CD(n_61137), .Q(ldtr[
		23]));
	notech_mux2 i_11356(.S(n_53557), .A(opb[23]), .B(ldtr[23]), .Z(n_24301)
		);
	notech_and4 i_137350668(.A(n_1168), .B(n_1263), .C(n_1169), .D(n_1170), 
		.Z(n_1266));
	notech_reg ldtr_reg_24(.CP(n_62225), .D(n_24307), .CD(n_61137), .Q(ldtr[
		24]));
	notech_mux2 i_11364(.S(n_53557), .A(opb[24]), .B(ldtr[24]), .Z(n_24307)
		);
	notech_reg ldtr_reg_25(.CP(n_62225), .D(n_24313), .CD(n_61136), .Q(ldtr[
		25]));
	notech_mux2 i_11372(.S(n_53557), .A(opb[25]), .B(ldtr[25]), .Z(n_24313)
		);
	notech_reg ldtr_reg_26(.CP(n_62225), .D(n_24319), .CD(n_61136), .Q(ldtr[
		26]));
	notech_mux2 i_11380(.S(n_53557), .A(opb[26]), .B(ldtr[26]), .Z(n_24319)
		);
	notech_and4 i_137050671(.A(n_1260), .B(n_1166), .C(n_2698), .D(n_1167), 
		.Z(n_1263));
	notech_reg ldtr_reg_27(.CP(n_62309), .D(n_24325), .CD(n_61136), .Q(ldtr[
		27]));
	notech_mux2 i_11389(.S(n_53557), .A(opb[27]), .B(ldtr[27]), .Z(n_24325)
		);
	notech_reg ldtr_reg_28(.CP(n_62309), .D(n_24331), .CD(n_61136), .Q(ldtr[
		28]));
	notech_mux2 i_11397(.S(n_53557), .A(opb[28]), .B(ldtr[28]), .Z(n_24331)
		);
	notech_reg ldtr_reg_29(.CP(n_62309), .D(n_24337), .CD(n_61137), .Q(ldtr[
		29]));
	notech_mux2 i_11405(.S(n_53557), .A(opb[29]), .B(ldtr[29]), .Z(n_24337)
		);
	notech_ao4 i_136750674(.A(n_1031), .B(n_59899), .C(n_107626780), .D(n_28714
		), .Z(n_1260));
	notech_reg ldtr_reg_30(.CP(n_62309), .D(n_24343), .CD(n_61137), .Q(ldtr[
		30]));
	notech_mux2 i_11413(.S(n_53557), .A(opb[30]), .B(ldtr[30]), .Z(n_24343)
		);
	notech_reg ldtr_reg_31(.CP(n_62309), .D(n_24349), .CD(n_61137), .Q(ldtr[
		31]));
	notech_mux2 i_11421(.S(n_53557), .A(opb[31]), .B(ldtr[31]), .Z(n_24349)
		);
	notech_reg gdtr_reg_0(.CP(n_62309), .D(n_24355), .CD(n_61137), .Q(gdtr[0
		]));
	notech_mux2 i_11429(.S(n_300986329), .A(opb[0]), .B(gdtr[0]), .Z(n_24355
		));
	notech_nand2 i_107150954(.A(n_1256), .B(n_1255), .Z(n_1257));
	notech_reg gdtr_reg_1(.CP(n_62309), .D(n_24361), .CD(n_61137), .Q(gdtr[1
		]));
	notech_mux2 i_11437(.S(n_300986329), .A(opb[1]), .B(gdtr[1]), .Z(n_24361
		));
	notech_ao4 i_106950956(.A(n_28987), .B(n_55405), .C(n_55404), .D(n_2700)
		, .Z(n_1256));
	notech_reg gdtr_reg_2(.CP(n_62309), .D(n_24368), .CD(n_61138), .Q(gdtr[2
		]));
	notech_mux2 i_11445(.S(n_300986329), .A(opb[2]), .B(gdtr[2]), .Z(n_24368
		));
	notech_ao4 i_106850957(.A(n_55062), .B(n_55600), .C(n_55064), .D(n_56784
		), .Z(n_1255));
	notech_reg gdtr_reg_3(.CP(n_62309), .D(n_24375), .CD(n_61141), .Q(gdtr[3
		]));
	notech_mux2 i_11453(.S(n_300986329), .A(opb[3]), .B(gdtr[3]), .Z(n_24375
		));
	notech_nand3 i_107050955(.A(n_43426147), .B(n_1157), .C(n_1162), .Z(n_1254
		));
	notech_reg gdtr_reg_4(.CP(n_62309), .D(n_24381), .CD(n_61141), .Q(gdtr[4
		]));
	notech_mux2 i_11461(.S(n_300986329), .A(opb[4]), .B(gdtr[4]), .Z(n_24381
		));
	notech_reg gdtr_reg_5(.CP(n_62309), .D(n_24387), .CD(n_61138), .Q(gdtr[5
		]));
	notech_mux2 i_11469(.S(n_300986329), .A(opb[5]), .B(gdtr[5]), .Z(n_24387
		));
	notech_reg gdtr_reg_6(.CP(n_62309), .D(n_24393), .CD(n_61138), .Q(gdtr[6
		]));
	notech_mux2 i_11477(.S(n_300986329), .A(opb[6]), .B(gdtr[6]), .Z(n_24393
		));
	notech_reg gdtr_reg_7(.CP(n_62309), .D(n_24399), .CD(n_61141), .Q(gdtr[7
		]));
	notech_mux2 i_11485(.S(n_300986329), .A(opb[7]), .B(gdtr[7]), .Z(n_24399
		));
	notech_nand3 i_100751018(.A(n_1152), .B(n_1248), .C(n_1153), .Z(n_1250)
		);
	notech_reg gdtr_reg_8(.CP(n_62309), .D(n_24405), .CD(n_61141), .Q(gdtr[8
		]));
	notech_mux2 i_11493(.S(n_300986329), .A(opb[8]), .B(gdtr[8]), .Z(n_24405
		));
	notech_reg gdtr_reg_9(.CP(n_62309), .D(n_24411), .CD(n_61141), .Q(gdtr[9
		]));
	notech_mux2 i_11501(.S(n_300986329), .A(opb[9]), .B(gdtr[9]), .Z(n_24411
		));
	notech_and3 i_100551020(.A(n_1246), .B(n_41726130), .C(n_1151), .Z(n_1248
		));
	notech_reg gdtr_reg_10(.CP(n_62309), .D(n_24417), .CD(n_61141), .Q(gdtr[
		10]));
	notech_mux2 i_11509(.S(n_300986329), .A(opb[10]), .B(gdtr[10]), .Z(n_24417
		));
	notech_reg gdtr_reg_11(.CP(n_62309), .D(n_24423), .CD(n_61141), .Q(gdtr[
		11]));
	notech_mux2 i_11517(.S(n_300986329), .A(opb[11]), .B(gdtr[11]), .Z(n_24423
		));
	notech_ao4 i_100351022(.A(n_2685), .B(n_43626149), .C(n_2671), .D(n_55342
		), .Z(n_1246));
	notech_reg gdtr_reg_12(.CP(n_62309), .D(n_24429), .CD(n_61138), .Q(gdtr[
		12]));
	notech_mux2 i_11525(.S(n_300986329), .A(opb[12]), .B(gdtr[12]), .Z(n_24429
		));
	notech_reg gdtr_reg_13(.CP(n_62309), .D(n_24435), .CD(n_61138), .Q(gdtr[
		13]));
	notech_mux2 i_11533(.S(n_300986329), .A(opb[13]), .B(gdtr[13]), .Z(n_24435
		));
	notech_reg gdtr_reg_14(.CP(n_62307), .D(n_24441), .CD(n_61138), .Q(gdtr[
		14]));
	notech_mux2 i_11541(.S(n_300986329), .A(opb[14]), .B(gdtr[14]), .Z(n_24441
		));
	notech_or4 i_89451124(.A(n_1143), .B(n_1240), .C(n_1144), .D(n_1145), .Z
		(n_1243));
	notech_reg gdtr_reg_15(.CP(n_62307), .D(n_24447), .CD(n_61138), .Q(gdtr[
		15]));
	notech_mux2 i_11549(.S(n_300986329), .A(opb[15]), .B(gdtr[15]), .Z(n_24447
		));
	notech_reg gdtr_reg_16(.CP(n_62369), .D(n_24453), .CD(n_61138), .Q(gdtr[
		16]));
	notech_mux2 i_11557(.S(n_53705), .A(opb[16]), .B(gdtr[16]), .Z(n_24453)
		);
	notech_reg gdtr_reg_17(.CP(n_62369), .D(n_24459), .CD(n_61138), .Q(gdtr[
		17]));
	notech_mux2 i_11565(.S(n_53705), .A(opb[17]), .B(gdtr[17]), .Z(n_24459)
		);
	notech_nand3 i_89151127(.A(n_43426147), .B(n_1141), .C(n_1142), .Z(n_1240
		));
	notech_reg gdtr_reg_18(.CP(n_62369), .D(n_24465), .CD(n_61138), .Q(gdtr[
		18]));
	notech_mux2 i_11574(.S(n_53705), .A(opb[18]), .B(gdtr[18]), .Z(n_24465)
		);
	notech_reg gdtr_reg_19(.CP(n_62369), .D(n_24471), .CD(n_61138), .Q(gdtr[
		19]));
	notech_mux2 i_11582(.S(n_53705), .A(opb[19]), .B(gdtr[19]), .Z(n_24471)
		);
	notech_and3 i_66951985(.A(n_2698), .B(n_1237), .C(n_1137), .Z(n_41726130
		));
	notech_reg gdtr_reg_20(.CP(n_62369), .D(n_24477), .CD(n_61138), .Q(gdtr[
		20]));
	notech_mux2 i_11590(.S(n_53705), .A(opb[20]), .B(gdtr[20]), .Z(n_24477)
		);
	notech_reg gdtr_reg_21(.CP(n_62369), .D(n_24483), .CD(n_61144), .Q(gdtr[
		21]));
	notech_mux2 i_11598(.S(n_53705), .A(opb[21]), .B(gdtr[21]), .Z(n_24483)
		);
	notech_ao4 i_86251154(.A(n_55810), .B(n_58960), .C(n_2699), .D(n_55920),
		 .Z(n_1237));
	notech_reg gdtr_reg_22(.CP(n_62369), .D(n_24489), .CD(n_61149), .Q(gdtr[
		22]));
	notech_mux2 i_11606(.S(n_53705), .A(opb[22]), .B(gdtr[22]), .Z(n_24489)
		);
	notech_reg gdtr_reg_23(.CP(n_62369), .D(n_24495), .CD(n_61149), .Q(gdtr[
		23]));
	notech_mux2 i_11614(.S(n_53705), .A(opb[23]), .B(gdtr[23]), .Z(n_24495)
		);
	notech_nand2 i_6551995(.A(opc_10[0]), .B(n_62405), .Z(n_43626149));
	notech_reg gdtr_reg_24(.CP(n_62369), .D(n_24503), .CD(n_61149), .Q(gdtr[
		24]));
	notech_mux2 i_11622(.S(n_53705), .A(opb[24]), .B(gdtr[24]), .Z(n_24503)
		);
	notech_reg gdtr_reg_25(.CP(n_62369), .D(n_24512), .CD(n_61149), .Q(gdtr[
		25]));
	notech_mux2 i_11630(.S(n_53705), .A(opb[25]), .B(gdtr[25]), .Z(n_24512)
		);
	notech_reg gdtr_reg_26(.CP(n_62369), .D(n_24520), .CD(n_61149), .Q(gdtr[
		26]));
	notech_mux2 i_11638(.S(n_53705), .A(opb[26]), .B(gdtr[26]), .Z(n_24520)
		);
	notech_ao4 i_80451205(.A(n_58483), .B(n_28019), .C(n_55947), .D(n_28985)
		, .Z(n_1234));
	notech_reg gdtr_reg_27(.CP(n_62077), .D(n_24526), .CD(n_61149), .Q(gdtr[
		27]));
	notech_mux2 i_11646(.S(n_53705), .A(opb[27]), .B(gdtr[27]), .Z(n_24526)
		);
	notech_ao4 i_80351206(.A(n_55965), .B(n_27985), .C(n_55992), .D(n_27953)
		, .Z(n_1233));
	notech_reg gdtr_reg_28(.CP(n_62369), .D(n_24532), .CD(n_61149), .Q(gdtr[
		28]));
	notech_mux2 i_11654(.S(n_53705), .A(opb[28]), .B(gdtr[28]), .Z(n_24532)
		);
	notech_and2 i_80751202(.A(n_1231), .B(n_1230), .Z(n_1232));
	notech_reg gdtr_reg_29(.CP(n_62369), .D(n_24538), .CD(n_61149), .Q(gdtr[
		29]));
	notech_mux2 i_11662(.S(n_53705), .A(opb[29]), .B(gdtr[29]), .Z(n_24538)
		);
	notech_ao4 i_80251207(.A(n_56009), .B(n_27919), .C(n_56033), .D(n_27885)
		, .Z(n_1231));
	notech_reg gdtr_reg_30(.CP(n_62369), .D(n_24544), .CD(n_61149), .Q(gdtr[
		30]));
	notech_mux2 i_11670(.S(n_53705), .A(opb[30]), .B(gdtr[30]), .Z(n_24544)
		);
	notech_ao4 i_80151208(.A(n_56043), .B(n_27850), .C(n_55879), .D(n_27818)
		, .Z(n_1230));
	notech_reg gdtr_reg_31(.CP(n_62369), .D(n_24550), .CD(n_61148), .Q(gdtr[
		31]));
	notech_mux2 i_11678(.S(n_53705), .A(opb[31]), .B(gdtr[31]), .Z(n_24550)
		);
	notech_and4 i_80951200(.A(n_1227), .B(n_1226), .C(n_1224), .D(n_1223), .Z
		(n_1229));
	notech_reg Daddrgs_reg_0(.CP(n_62369), .D(n_15967), .CD(n_61148), .Q(Daddrgs
		[0]));
	notech_reg Daddrgs_reg_1(.CP(n_62369), .D(n_15974), .CD(n_61148), .Q(Daddrgs
		[1]));
	notech_reg Daddrgs_reg_2(.CP(n_62307), .D(n_15981), .CD(n_61148), .Q(Daddrgs
		[2]));
	notech_reg Daddrgs_reg_3(.CP(n_62307), .D(n_15988), .CD(n_61148), .Q(Daddrgs
		[3]));
	notech_reg Daddrgs_reg_4(.CP(n_62307), .D(n_15995), .CD(n_61149), .Q(Daddrgs
		[4]));
	notech_reg Daddrgs_reg_5(.CP(n_62307), .D(n_16002), .CD(n_61149), .Q(Daddrgs
		[5]));
	notech_reg Daddrgs_reg_6(.CP(n_62307), .D(n_16009), .CD(n_61148), .Q(Daddrgs
		[6]));
	notech_reg Daddrgs_reg_7(.CP(n_62307), .D(n_16016), .CD(n_61148), .Q(Daddrgs
		[7]));
	notech_reg Daddrgs_reg_8(.CP(n_62307), .D(n_16023), .CD(n_61149), .Q(Daddrgs
		[8]));
	notech_reg Daddrgs_reg_9(.CP(n_62307), .D(n_16030), .CD(n_61152), .Q(Daddrgs
		[9]));
	notech_reg Daddrgs_reg_10(.CP(n_62307), .D(n_16037), .CD(n_61152), .Q(Daddrgs
		[10]));
	notech_reg Daddrgs_reg_11(.CP(n_62369), .D(n_16044), .CD(n_61152), .Q(Daddrgs
		[11]));
	notech_reg Daddrgs_reg_12(.CP(n_62365), .D(n_16051), .CD(n_61152), .Q(Daddrgs
		[12]));
	notech_reg Daddrgs_reg_13(.CP(n_62305), .D(n_16058), .CD(n_61152), .Q(Daddrgs
		[13]));
	notech_reg Daddrgs_reg_14(.CP(n_62365), .D(n_16065), .CD(n_61153), .Q(Daddrgs
		[14]));
	notech_reg Daddrgs_reg_15(.CP(n_62365), .D(n_16072), .CD(n_61153), .Q(Daddrgs
		[15]));
	notech_reg Daddrgs_reg_16(.CP(n_62365), .D(n_16079), .CD(n_61153), .Q(Daddrgs
		[16]));
	notech_reg Daddrgs_reg_17(.CP(n_62365), .D(n_16086), .CD(n_61153), .Q(Daddrgs
		[17]));
	notech_reg Daddrgs_reg_18(.CP(n_62365), .D(n_16093), .CD(n_61152), .Q(Daddrgs
		[18]));
	notech_reg Daddrgs_reg_19(.CP(n_62365), .D(n_16100), .CD(n_61152), .Q(Daddrgs
		[19]));
	notech_reg Daddrgs_reg_20(.CP(n_62365), .D(n_16107), .CD(n_61149), .Q(Daddrgs
		[20]));
	notech_reg Daddrgs_reg_21(.CP(n_62365), .D(n_16114), .CD(n_61152), .Q(Daddrgs
		[21]));
	notech_reg Daddrgs_reg_22(.CP(n_62365), .D(n_16121), .CD(n_61152), .Q(Daddrgs
		[22]));
	notech_reg Daddrgs_reg_23(.CP(n_62365), .D(n_16128), .CD(n_61152), .Q(Daddrgs
		[23]));
	notech_reg Daddrgs_reg_24(.CP(n_62389), .D(n_16135), .CD(n_61152), .Q(Daddrgs
		[24]));
	notech_reg Daddrgs_reg_25(.CP(n_62389), .D(n_16142), .CD(n_61152), .Q(Daddrgs
		[25]));
	notech_reg Daddrgs_reg_26(.CP(n_62389), .D(n_16149), .CD(n_61152), .Q(Daddrgs
		[26]));
	notech_reg Daddrgs_reg_27(.CP(n_62389), .D(n_16156), .CD(n_61148), .Q(Daddrgs
		[27]));
	notech_reg Daddrgs_reg_28(.CP(n_62389), .D(n_16163), .CD(n_61146), .Q(Daddrgs
		[28]));
	notech_reg Daddrgs_reg_29(.CP(n_62389), .D(n_16170), .CD(n_61146), .Q(Daddrgs
		[29]));
	notech_reg Daddrgs_reg_30(.CP(n_62389), .D(n_16177), .CD(n_61146), .Q(Daddrgs
		[30]));
	notech_reg Daddrgs_reg_31(.CP(n_62389), .D(n_16184), .CD(n_61146), .Q(Daddrgs
		[31]));
	notech_reg idtr_reg_0(.CP(n_62389), .D(n_24621), .CD(n_61146), .Q(idtr[0
		]));
	notech_mux2 i_11819(.S(n_300886328), .A(opb[0]), .B(idtr[0]), .Z(n_24621
		));
	notech_reg idtr_reg_1(.CP(n_62389), .D(n_24627), .CD(n_61146), .Q(idtr[1
		]));
	notech_mux2 i_11827(.S(n_300886328), .A(opb[1]), .B(idtr[1]), .Z(n_24627
		));
	notech_ao4 i_80051209(.A(n_55934), .B(n_27786), .C(n_55893), .D(n_27747)
		, .Z(n_1227));
	notech_reg idtr_reg_2(.CP(n_62389), .D(n_24633), .CD(n_61146), .Q(idtr[2
		]));
	notech_mux2 i_11835(.S(n_300886328), .A(opb[2]), .B(idtr[2]), .Z(n_24633
		));
	notech_ao4 i_79951210(.A(n_55906), .B(n_27715), .C(n_55924), .D(n_27370)
		, .Z(n_1226));
	notech_reg idtr_reg_3(.CP(n_62389), .D(n_24639), .CD(n_61146), .Q(idtr[3
		]));
	notech_mux2 i_11843(.S(n_300886328), .A(opb[3]), .B(idtr[3]), .Z(n_24639
		));
	notech_reg idtr_reg_4(.CP(n_62389), .D(n_24645), .CD(n_61146), .Q(idtr[4
		]));
	notech_mux2 i_11851(.S(n_300886328), .A(opb[4]), .B(idtr[4]), .Z(n_24645
		));
	notech_ao4 i_79851211(.A(n_56092), .B(n_27681), .C(n_56126), .D(n_27639)
		, .Z(n_1224));
	notech_reg idtr_reg_5(.CP(n_62389), .D(n_24651), .CD(n_61144), .Q(idtr[5
		]));
	notech_mux2 i_11861(.S(n_300886328), .A(opb[5]), .B(idtr[5]), .Z(n_24651
		));
	notech_ao4 i_79751212(.A(n_56139), .B(n_27602), .C(n_56382), .D(n_27559)
		, .Z(n_1223));
	notech_reg idtr_reg_6(.CP(n_62389), .D(n_24657), .CD(n_61144), .Q(idtr[6
		]));
	notech_mux2 i_11869(.S(n_300886328), .A(opb[6]), .B(idtr[6]), .Z(n_24657
		));
	notech_nand2 i_1251997(.A(n_62427), .B(opc[0]), .Z(n_46226175));
	notech_reg idtr_reg_7(.CP(n_62389), .D(n_24664), .CD(n_61144), .Q(idtr[7
		]));
	notech_mux2 i_11877(.S(n_300886328), .A(opb[7]), .B(idtr[7]), .Z(n_24664
		));
	notech_reg idtr_reg_8(.CP(n_62389), .D(n_24670), .CD(n_61144), .Q(idtr[8
		]));
	notech_mux2 i_11885(.S(n_300886328), .A(opb[8]), .B(idtr[8]), .Z(n_24670
		));
	notech_and4 i_63151370(.A(n_1112), .B(n_1111), .C(n_1218), .D(n_1115), .Z
		(n_1221));
	notech_reg idtr_reg_9(.CP(n_62389), .D(n_24676), .CD(n_61144), .Q(idtr[9
		]));
	notech_mux2 i_11893(.S(n_300886328), .A(opb[9]), .B(idtr[9]), .Z(n_24676
		));
	notech_reg idtr_reg_10(.CP(n_62365), .D(n_24682), .CD(n_61146), .Q(idtr[
		10]));
	notech_mux2 i_11901(.S(n_300886328), .A(opb[10]), .B(idtr[10]), .Z(n_24682
		));
	notech_reg idtr_reg_11(.CP(n_62389), .D(n_24689), .CD(n_61146), .Q(idtr[
		11]));
	notech_mux2 i_11909(.S(n_300886328), .A(opb[11]), .B(idtr[11]), .Z(n_24689
		));
	notech_and3 i_62751374(.A(n_1216), .B(n_1215), .C(n_1110), .Z(n_1218));
	notech_reg idtr_reg_12(.CP(n_62367), .D(n_24695), .CD(n_61144), .Q(idtr[
		12]));
	notech_mux2 i_11917(.S(n_300886328), .A(opb[12]), .B(idtr[12]), .Z(n_24695
		));
	notech_reg idtr_reg_13(.CP(n_62367), .D(n_24701), .CD(n_61146), .Q(idtr[
		13]));
	notech_mux2 i_11925(.S(n_300886328), .A(opb[13]), .B(idtr[13]), .Z(n_24701
		));
	notech_ao4 i_62451377(.A(n_58922), .B(n_28982), .C(n_55492), .D(n_27526)
		, .Z(n_1216));
	notech_reg idtr_reg_14(.CP(n_62367), .D(n_24707), .CD(n_61146), .Q(idtr[
		14]));
	notech_mux2 i_11933(.S(n_300886328), .A(opb[14]), .B(idtr[14]), .Z(n_24707
		));
	notech_ao4 i_62551376(.A(n_57351), .B(n_55216), .C(n_28983), .D(n_55236)
		, .Z(n_1215));
	notech_reg idtr_reg_15(.CP(n_62367), .D(n_24713), .CD(n_61147), .Q(idtr[
		15]));
	notech_mux2 i_11941(.S(n_300886328), .A(opb[15]), .B(idtr[15]), .Z(n_24713
		));
	notech_or4 i_120351973(.A(n_56460), .B(n_55522), .C(n_205188862), .D(n_56440
		), .Z(n_54526258));
	notech_reg idtr_reg_16(.CP(n_62367), .D(n_24719), .CD(n_61147), .Q(idtr[
		16]));
	notech_mux2 i_11949(.S(n_53716), .A(opb[16]), .B(idtr[16]), .Z(n_24719)
		);
	notech_reg idtr_reg_17(.CP(n_62367), .D(n_24725), .CD(n_61147), .Q(idtr[
		17]));
	notech_mux2 i_11957(.S(n_53716), .A(opb[17]), .B(idtr[17]), .Z(n_24725)
		);
	notech_ao4 i_63051371(.A(n_2691), .B(n_55400), .C(n_2690), .D(n_27570), 
		.Z(n_1213));
	notech_reg idtr_reg_18(.CP(n_62367), .D(n_24731), .CD(n_61147), .Q(idtr[
		18]));
	notech_mux2 i_11965(.S(n_53716), .A(opb[18]), .B(idtr[18]), .Z(n_24731)
		);
	notech_reg idtr_reg_19(.CP(n_62367), .D(n_24737), .CD(n_61148), .Q(idtr[
		19]));
	notech_mux2 i_11973(.S(n_53716), .A(opb[19]), .B(idtr[19]), .Z(n_24737)
		);
	notech_reg idtr_reg_20(.CP(n_62367), .D(n_24743), .CD(n_61148), .Q(idtr[
		20]));
	notech_mux2 i_11981(.S(n_53716), .A(opb[20]), .B(idtr[20]), .Z(n_24743)
		);
	notech_ao4 i_63251369(.A(n_2680), .B(n_55426267), .C(n_2675), .D(n_55687
		), .Z(n_1210));
	notech_reg idtr_reg_21(.CP(n_62367), .D(n_24749), .CD(n_61148), .Q(idtr[
		21]));
	notech_mux2 i_11989(.S(n_53716), .A(opb[21]), .B(idtr[21]), .Z(n_24749)
		);
	notech_or4 i_118951976(.A(n_56460), .B(n_55522), .C(n_1105), .D(n_56440)
		, .Z(n_55426267));
	notech_reg idtr_reg_22(.CP(n_62367), .D(n_24755), .CD(n_61148), .Q(idtr[
		22]));
	notech_mux2 i_11997(.S(n_53716), .A(opb[22]), .B(idtr[22]), .Z(n_24755)
		);
	notech_reg idtr_reg_23(.CP(n_62367), .D(n_24761), .CD(n_61148), .Q(idtr[
		23]));
	notech_mux2 i_12005(.S(n_53716), .A(opb[23]), .B(idtr[23]), .Z(n_24761)
		);
	notech_reg idtr_reg_24(.CP(n_62367), .D(n_24767), .CD(n_61147), .Q(idtr[
		24]));
	notech_mux2 i_12013(.S(n_53716), .A(opb[24]), .B(idtr[24]), .Z(n_24767)
		);
	notech_reg idtr_reg_25(.CP(n_62367), .D(n_24773), .CD(n_61147), .Q(idtr[
		25]));
	notech_mux2 i_12021(.S(n_53716), .A(opb[25]), .B(idtr[25]), .Z(n_24773)
		);
	notech_ao4 i_51751471(.A(n_58487), .B(n_28026), .C(n_55947), .D(n_28981)
		, .Z(n_1206));
	notech_reg idtr_reg_26(.CP(n_62367), .D(n_24779), .CD(n_61147), .Q(idtr[
		26]));
	notech_mux2 i_12029(.S(n_53716), .A(opb[26]), .B(idtr[26]), .Z(n_24779)
		);
	notech_ao4 i_51651472(.A(n_55972), .B(n_27992), .C(n_55992), .D(n_27960)
		, .Z(n_1205));
	notech_reg idtr_reg_27(.CP(n_62367), .D(n_24785), .CD(n_61147), .Q(idtr[
		27]));
	notech_mux2 i_12037(.S(n_53716), .A(opb[27]), .B(idtr[27]), .Z(n_24785)
		);
	notech_and2 i_52551468(.A(n_1203), .B(n_1202), .Z(n_1204));
	notech_reg idtr_reg_28(.CP(n_62367), .D(n_24791), .CD(n_61147), .Q(idtr[
		28]));
	notech_mux2 i_12045(.S(n_53716), .A(opb[28]), .B(idtr[28]), .Z(n_24791)
		);
	notech_ao4 i_51551473(.A(n_56013), .B(n_27926), .C(n_56033), .D(n_27894)
		, .Z(n_1203));
	notech_reg idtr_reg_29(.CP(n_62367), .D(n_24797), .CD(n_61147), .Q(idtr[
		29]));
	notech_mux2 i_12053(.S(n_53716), .A(opb[29]), .B(idtr[29]), .Z(n_24797)
		);
	notech_ao4 i_51451474(.A(n_56049), .B(n_27857), .C(n_55879), .D(n_27825)
		, .Z(n_1202));
	notech_reg idtr_reg_30(.CP(n_62367), .D(n_24803), .CD(n_61147), .Q(idtr[
		30]));
	notech_mux2 i_12061(.S(n_53716), .A(opb[30]), .B(idtr[30]), .Z(n_24803)
		);
	notech_and4 i_52851466(.A(n_1199), .B(n_1198), .C(n_1196), .D(n_1195), .Z
		(n_1201));
	notech_reg idtr_reg_31(.CP(n_62305), .D(n_24809), .CD(n_61147), .Q(idtr[
		31]));
	notech_mux2 i_12069(.S(n_53716), .A(opb[31]), .B(idtr[31]), .Z(n_24809)
		);
	notech_reg tr_reg_3(.CP(n_62305), .D(n_24815), .CD(n_61147), .Q(\tr[3] )
		);
	notech_mux2 i_12077(.S(n_300786327), .A(opb[3]), .B(\tr[3] ), .Z(n_24815
		));
	notech_ao4 i_51351475(.A(n_55934), .B(n_27793), .C(n_55893), .D(n_27754)
		, .Z(n_1199));
	notech_reg tr_reg_4(.CP(n_62305), .D(n_24821), .CD(n_61136), .Q(\tr[4] )
		);
	notech_mux2 i_12085(.S(n_300786327), .A(opb[4]), .B(\tr[4] ), .Z(n_24821
		));
	notech_ao4 i_51251476(.A(n_55910), .B(n_27722), .C(n_55924), .D(n_27377)
		, .Z(n_1198));
	notech_reg tr_reg_5(.CP(n_62305), .D(n_24827), .CD(n_61124), .Q(\tr[5] )
		);
	notech_mux2 i_12093(.S(n_300786327), .A(opb[5]), .B(\tr[5] ), .Z(n_24827
		));
	notech_reg tr_reg_6(.CP(n_62305), .D(n_24833), .CD(n_61124), .Q(\tr[6] )
		);
	notech_mux2 i_12101(.S(n_300786327), .A(opb[6]), .B(\tr[6] ), .Z(n_24833
		));
	notech_ao4 i_51151477(.A(n_56092), .B(n_27690), .C(n_56130), .D(n_27647)
		, .Z(n_1196));
	notech_reg tr_reg_7(.CP(n_62305), .D(n_24839), .CD(n_61124), .Q(\tr[7] )
		);
	notech_mux2 i_12109(.S(n_300786327), .A(opb[7]), .B(\tr[7] ), .Z(n_24839
		));
	notech_ao4 i_51051478(.A(n_56144), .B(n_27613), .C(n_56386), .D(n_28980)
		, .Z(n_1195));
	notech_reg tr_reg_8(.CP(n_62305), .D(n_24845), .CD(n_61124), .Q(\tr[8] )
		);
	notech_mux2 i_12117(.S(n_300786327), .A(opb[8]), .B(\tr[8] ), .Z(n_24845
		));
	notech_reg tr_reg_9(.CP(n_62305), .D(n_24851), .CD(n_61124), .Q(\tr[9] )
		);
	notech_mux2 i_12125(.S(n_300786327), .A(opb[9]), .B(\tr[9] ), .Z(n_24851
		));
	notech_reg tr_reg_10(.CP(n_62305), .D(n_24857), .CD(n_61124), .Q(\tr[10] 
		));
	notech_mux2 i_12133(.S(n_300786327), .A(opb[10]), .B(\tr[10] ), .Z(n_24857
		));
	notech_reg tr_reg_11(.CP(n_62225), .D(n_24863), .CD(n_61124), .Q(\tr[11] 
		));
	notech_mux2 i_12141(.S(n_300786327), .A(opb[11]), .B(\tr[11] ), .Z(n_24863
		));
	notech_reg tr_reg_12(.CP(n_62305), .D(n_24869), .CD(n_61124), .Q(\tr[12] 
		));
	notech_mux2 i_12149(.S(n_300786327), .A(opb[12]), .B(\tr[12] ), .Z(n_24869
		));
	notech_reg tr_reg_13(.CP(n_62311), .D(n_24875), .CD(n_61124), .Q(\tr[13] 
		));
	notech_mux2 i_12157(.S(n_300786327), .A(opb[13]), .B(\tr[13] ), .Z(n_24875
		));
	notech_nao3 i_19951774(.A(n_56487), .B(n_56440), .C(n_56478), .Z(n_1189)
		);
	notech_reg tr_reg_14(.CP(n_62227), .D(n_24881), .CD(n_61123), .Q(\tr[14] 
		));
	notech_mux2 i_12165(.S(n_300786327), .A(opb[14]), .B(\tr[14] ), .Z(n_24881
		));
	notech_ao4 i_35751989(.A(n_56502), .B(n_56560), .C(n_55807), .D(n_26574)
		, .Z(n_1188));
	notech_reg tr_reg_15(.CP(n_62227), .D(n_24887), .CD(n_61123), .Q(\tr[15] 
		));
	notech_mux2 i_12173(.S(n_300786327), .A(opb[15]), .B(\tr[15] ), .Z(n_24887
		));
	notech_reg desc_reg_0(.CP(n_62227), .D(n_24893), .CD(n_61123), .Q(desc[0
		]));
	notech_mux2 i_12181(.S(n_57461), .A(read_data[0]), .B(desc[0]), .Z(n_24893
		));
	notech_reg desc_reg_1(.CP(n_62227), .D(n_24899), .CD(n_61123), .Q(desc[1
		]));
	notech_mux2 i_12189(.S(n_57461), .A(read_data[1]), .B(desc[1]), .Z(n_24899
		));
	notech_reg desc_reg_2(.CP(n_62227), .D(n_24905), .CD(n_61123), .Q(desc[2
		]));
	notech_mux2 i_12197(.S(n_57461), .A(read_data[2]), .B(desc[2]), .Z(n_24905
		));
	notech_ao4 i_10351870(.A(n_55934), .B(n_27803), .C(n_58487), .D(n_28036)
		, .Z(n_1184));
	notech_reg desc_reg_3(.CP(n_62227), .D(n_24911), .CD(n_61124), .Q(desc[3
		]));
	notech_mux2 i_12205(.S(n_57461), .A(read_data[3]), .B(desc[3]), .Z(n_24911
		));
	notech_ao4 i_10251871(.A(n_55952), .B(n_28979), .C(n_55972), .D(n_28002)
		, .Z(n_1183));
	notech_reg desc_reg_4(.CP(n_62227), .D(n_24917), .CD(n_61124), .Q(desc[4
		]));
	notech_mux2 i_12213(.S(n_57461), .A(read_data[4]), .B(desc[4]), .Z(n_24917
		));
	notech_and2 i_10651867(.A(n_1181), .B(n_1180), .Z(n_1182));
	notech_reg desc_reg_5(.CP(n_62227), .D(n_24923), .CD(n_61123), .Q(desc[5
		]));
	notech_mux2 i_12221(.S(n_57461), .A(read_data[5]), .B(desc[5]), .Z(n_24923
		));
	notech_ao4 i_10151872(.A(n_55992), .B(n_27970), .C(n_56013), .D(n_27937)
		, .Z(n_1181));
	notech_reg desc_reg_6(.CP(n_62227), .D(n_24929), .CD(n_61123), .Q(desc[6
		]));
	notech_mux2 i_12229(.S(n_57461), .A(read_data[6]), .B(desc[6]), .Z(n_24929
		));
	notech_ao4 i_10051873(.A(n_56033), .B(n_27904), .C(n_56049), .D(n_27868)
		, .Z(n_1180));
	notech_reg desc_reg_7(.CP(n_62313), .D(n_24935), .CD(n_61124), .Q(desc[7
		]));
	notech_mux2 i_12237(.S(n_57461), .A(read_data[7]), .B(desc[7]), .Z(n_24935
		));
	notech_and4 i_10851865(.A(n_1177), .B(n_1176), .C(n_1174), .D(n_1173), .Z
		(n_1179));
	notech_reg desc_reg_8(.CP(n_62313), .D(n_24941), .CD(n_61125), .Q(desc[8
		]));
	notech_mux2 i_12245(.S(n_57461), .A(read_data[8]), .B(desc[8]), .Z(n_24941
		));
	notech_reg desc_reg_9(.CP(n_62313), .D(n_24947), .CD(n_61126), .Q(desc[9
		]));
	notech_mux2 i_12253(.S(n_57461), .A(read_data[9]), .B(desc[9]), .Z(n_24947
		));
	notech_ao4 i_9951874(.A(n_55879), .B(n_27835), .C(n_55893), .D(n_27768),
		 .Z(n_1177));
	notech_reg desc_reg_10(.CP(n_62313), .D(n_24953), .CD(n_61125), .Q(desc[
		10]));
	notech_mux2 i_12261(.S(n_57461), .A(read_data[10]), .B(desc[10]), .Z(n_24953
		));
	notech_ao4 i_9851875(.A(n_55910), .B(n_27732), .C(n_55924), .D(n_27387),
		 .Z(n_1176));
	notech_reg desc_reg_11(.CP(n_62313), .D(n_24959), .CD(n_61125), .Q(desc[
		11]));
	notech_mux2 i_12269(.S(n_57461), .A(read_data[11]), .B(desc[11]), .Z(n_24959
		));
	notech_reg desc_reg_12(.CP(n_62313), .D(n_24967), .CD(n_61126), .Q(desc[
		12]));
	notech_mux2 i_12277(.S(n_57461), .A(read_data[12]), .B(desc[12]), .Z(n_24967
		));
	notech_ao4 i_9751876(.A(n_56092), .B(n_27700), .C(n_56130), .D(n_27660),
		 .Z(n_1174));
	notech_reg desc_reg_13(.CP(n_62313), .D(n_24974), .CD(n_61126), .Q(desc[
		13]));
	notech_mux2 i_12285(.S(n_58532), .A(read_data[13]), .B(desc[13]), .Z(n_24974
		));
	notech_ao4 i_9651877(.A(n_56144), .B(n_27623), .C(n_56386), .D(n_28978),
		 .Z(n_1173));
	notech_reg desc_reg_14(.CP(n_62313), .D(n_24981), .CD(n_61126), .Q(desc[
		14]));
	notech_mux2 i_12293(.S(n_58532), .A(read_data[14]), .B(desc[14]), .Z(n_24981
		));
	notech_or4 i_121900(.A(n_1171), .B(n_1172), .C(n_1164), .D(n_27344), .Z(n_12049
		));
	notech_reg desc_reg_15(.CP(n_62313), .D(n_24988), .CD(n_61126), .Q(desc[
		15]));
	notech_mux2 i_12301(.S(n_58532), .A(read_data[15]), .B(desc[15]), .Z(n_24988
		));
	notech_nor2 i_136150680(.A(n_2667), .B(n_28986), .Z(n_1172));
	notech_reg desc_reg_16(.CP(n_62313), .D(n_24994), .CD(n_61126), .Q(desc[
		16]));
	notech_mux2 i_12309(.S(n_58532), .A(read_data[16]), .B(desc[16]), .Z(n_24994
		));
	notech_nor2 i_135950682(.A(n_2665), .B(n_55356), .Z(n_1171));
	notech_reg desc_reg_17(.CP(n_62313), .D(n_25001), .CD(n_61125), .Q(desc[
		17]));
	notech_mux2 i_12317(.S(n_58532), .A(read_data[17]), .B(desc[17]), .Z(n_25001
		));
	notech_or2 i_136250679(.A(n_2699), .B(n_2668), .Z(n_1170));
	notech_reg desc_reg_18(.CP(n_62313), .D(n_25007), .CD(n_61125), .Q(desc[
		18]));
	notech_mux2 i_12325(.S(n_58532), .A(read_data[18]), .B(desc[18]), .Z(n_25007
		));
	notech_nao3 i_136650675(.A(n_62427), .B(opc[0]), .C(n_2697), .Z(n_1169)
		);
	notech_reg desc_reg_19(.CP(n_62313), .D(n_25015), .CD(n_61125), .Q(desc[
		19]));
	notech_mux2 i_12333(.S(n_58532), .A(read_data[19]), .B(desc[19]), .Z(n_25015
		));
	notech_or4 i_136450677(.A(n_56081), .B(n_56114), .C(n_55827), .D(n_2688)
		, .Z(n_1168));
	notech_reg desc_reg_20(.CP(n_62313), .D(n_25022), .CD(n_61125), .Q(desc[
		20]));
	notech_mux2 i_12341(.S(n_58532), .A(read_data[20]), .B(desc[20]), .Z(n_25022
		));
	notech_nao3 i_136550676(.A(opc_10[0]), .B(opcode_289113), .C(n_54606), .Z
		(n_1167));
	notech_reg desc_reg_21(.CP(n_62313), .D(n_25028), .CD(n_61125), .Q(desc[
		21]));
	notech_mux2 i_12350(.S(n_58532), .A(read_data[21]), .B(desc[21]), .Z(n_25028
		));
	notech_or4 i_136350678(.A(n_56081), .B(n_56114), .C(n_54089), .D(n_55342
		), .Z(n_1166));
	notech_reg desc_reg_22(.CP(n_62313), .D(n_25034), .CD(n_61125), .Q(desc[
		22]));
	notech_mux2 i_12358(.S(n_58532), .A(read_data[22]), .B(desc[22]), .Z(n_25034
		));
	notech_reg desc_reg_23(.CP(n_62313), .D(n_25040), .CD(n_61125), .Q(desc[
		23]));
	notech_mux2 i_12366(.S(n_58532), .A(read_data[23]), .B(desc[23]), .Z(n_25040
		));
	notech_nor2 i_136050681(.A(n_2666), .B(n_58960), .Z(n_1164));
	notech_reg desc_reg_24(.CP(n_62313), .D(n_25046), .CD(n_61125), .Q(desc[
		24]));
	notech_mux2 i_12374(.S(n_355776393), .A(read_data[24]), .B(desc[24]), .Z
		(n_25046));
	notech_or4 i_1820989(.A(n_1257), .B(n_1254), .C(n_1163), .D(n_1156), .Z(n_16801
		));
	notech_reg desc_reg_25(.CP(n_62313), .D(n_25052), .CD(n_61125), .Q(desc[
		25]));
	notech_mux2 i_12382(.S(n_355776393), .A(read_data[25]), .B(desc[25]), .Z
		(n_25052));
	notech_ao3 i_106650959(.A(opc_10[17]), .B(opcode_289113), .C(n_308418861
		), .Z(n_1163));
	notech_reg desc_reg_26(.CP(n_62371), .D(n_25058), .CD(n_61123), .Q(desc[
		26]));
	notech_mux2 i_12390(.S(n_355776393), .A(read_data[26]), .B(desc[26]), .Z
		(n_25058));
	notech_or4 i_106450961(.A(n_56196), .B(n_58660), .C(n_56369), .D(n_27583
		), .Z(n_1162));
	notech_reg desc_reg_27(.CP(n_62311), .D(n_25064), .CD(n_61120), .Q(desc[
		27]));
	notech_mux2 i_12398(.S(n_355776393), .A(read_data[27]), .B(desc[27]), .Z
		(n_25064));
	notech_reg desc_reg_28(.CP(n_62371), .D(n_25070), .CD(n_61120), .Q(desc[
		28]));
	notech_mux2 i_12406(.S(n_355776393), .A(read_data[28]), .B(desc[28]), .Z
		(n_25070));
	notech_reg desc_reg_29(.CP(n_62371), .D(n_25076), .CD(n_61120), .Q(desc[
		29]));
	notech_mux2 i_12414(.S(n_355776393), .A(read_data[29]), .B(desc[29]), .Z
		(n_25076));
	notech_reg desc_reg_30(.CP(n_62371), .D(n_25082), .CD(n_61120), .Q(desc[
		30]));
	notech_mux2 i_12422(.S(n_355776393), .A(read_data[30]), .B(desc[30]), .Z
		(n_25082));
	notech_reg desc_reg_31(.CP(n_62371), .D(n_25088), .CD(n_61120), .Q(desc[
		31]));
	notech_mux2 i_12430(.S(n_355776393), .A(read_data[31]), .B(desc[31]), .Z
		(n_25088));
	notech_or2 i_105950966(.A(n_55424), .B(n_58978), .Z(n_1157));
	notech_reg Daddrs_reg_0(.CP(n_62371), .D(n_25094), .CD(n_61120), .Q(Daddr
		[0]));
	notech_mux2 i_12438(.S(\nbus_11354[0] ), .A(Daddr[0]), .B(n_20843), .Z(n_25094
		));
	notech_nor2 i_106550960(.A(n_2648), .B(n_309618873), .Z(n_1156));
	notech_reg Daddrs_reg_1(.CP(n_62371), .D(n_25100), .CD(n_61120), .Q(Daddr
		[1]));
	notech_mux2 i_12447(.S(\nbus_11354[0] ), .A(Daddr[1]), .B(n_20849), .Z(n_25100
		));
	notech_or4 i_120716(.A(n_1154), .B(n_1250), .C(n_1155), .D(n_1148), .Z(n_19437
		));
	notech_reg Daddrs_reg_2(.CP(n_62371), .D(n_25106), .CD(n_61120), .Q(Daddr
		[2]));
	notech_mux2 i_12455(.S(\nbus_11354[0] ), .A(Daddr[2]), .B(n_20855), .Z(n_25106
		));
	notech_nor2 i_99551030(.A(n_2669), .B(n_55356), .Z(n_1155));
	notech_reg Daddrs_reg_3(.CP(n_62371), .D(n_25112), .CD(n_61120), .Q(Daddr
		[3]));
	notech_mux2 i_12463(.S(\nbus_11354[0] ), .A(Daddr[3]), .B(n_20861), .Z(n_25112
		));
	notech_nor2 i_99951026(.A(n_54468), .B(n_28986), .Z(n_1154));
	notech_reg Daddrs_reg_4(.CP(n_62371), .D(n_25118), .CD(n_61119), .Q(Daddr
		[4]));
	notech_mux2 i_12471(.S(\nbus_11354[0] ), .A(Daddr[4]), .B(n_20867), .Z(n_25118
		));
	notech_or2 i_99851027(.A(n_2699), .B(n_54428), .Z(n_1153));
	notech_reg Daddrs_reg_5(.CP(n_62371), .D(n_25124), .CD(n_61119), .Q(Daddr
		[5]));
	notech_mux2 i_12479(.S(\nbus_11354[0] ), .A(Daddr[5]), .B(n_20873), .Z(n_25124
		));
	notech_or4 i_100251023(.A(n_56177), .B(n_56163), .C(n_2688), .D(n_55827)
		, .Z(n_1152));
	notech_reg Daddrs_reg_6(.CP(n_62371), .D(n_25130), .CD(n_61119), .Q(Daddr
		[6]));
	notech_mux2 i_12487(.S(\nbus_11354[0] ), .A(Daddr[6]), .B(n_20879), .Z(n_25130
		));
	notech_nao3 i_100051025(.A(n_62427), .B(n_59113), .C(n_2684), .Z(n_1151)
		);
	notech_reg Daddrs_reg_7(.CP(n_62371), .D(n_25136), .CD(n_61119), .Q(Daddr
		[7]));
	notech_mux2 i_12495(.S(\nbus_11354[0] ), .A(Daddr[7]), .B(n_20885), .Z(n_25136
		));
	notech_reg Daddrs_reg_8(.CP(n_62371), .D(n_25142), .CD(n_61119), .Q(Daddr
		[8]));
	notech_mux2 i_12503(.S(\nbus_11354[0] ), .A(Daddr[8]), .B(n_20891), .Z(n_25142
		));
	notech_reg Daddrs_reg_9(.CP(n_62371), .D(n_25148), .CD(n_61119), .Q(Daddr
		[9]));
	notech_mux2 i_12511(.S(\nbus_11354[0] ), .A(Daddr[9]), .B(n_20897), .Z(n_25148
		));
	notech_and2 i_99651029(.A(n_2670), .B(opa[0]), .Z(n_1148));
	notech_reg Daddrs_reg_10(.CP(n_62371), .D(n_25154), .CD(n_61119), .Q(Daddr
		[10]));
	notech_mux2 i_12519(.S(\nbus_11354[0] ), .A(Daddr[10]), .B(n_20903), .Z(n_25154
		));
	notech_or4 i_1820733(.A(n_1146), .B(n_1243), .C(n_1147), .D(n_1140), .Z(n_19539
		));
	notech_reg Daddrs_reg_11(.CP(n_62371), .D(n_25160), .CD(n_61119), .Q(Daddr
		[11]));
	notech_mux2 i_12527(.S(\nbus_11354[0] ), .A(Daddr[11]), .B(n_20909), .Z(n_25160
		));
	notech_nor2 i_88351135(.A(n_2700), .B(n_2655), .Z(n_1147));
	notech_reg Daddrs_reg_12(.CP(n_62371), .D(n_25166), .CD(n_61119), .Q(Daddr
		[12]));
	notech_mux2 i_12535(.S(\nbus_11354[0] ), .A(Daddr[12]), .B(n_20915), .Z(n_25166
		));
	notech_nor2 i_88651132(.A(n_55068), .B(n_56784), .Z(n_1146));
	notech_reg Daddrs_reg_13(.CP(n_62371), .D(n_25172), .CD(n_61120), .Q(Daddr
		[13]));
	notech_mux2 i_12543(.S(\nbus_11354[0] ), .A(Daddr[13]), .B(n_20921), .Z(n_25172
		));
	notech_nor2 i_88751131(.A(n_55069), .B(n_55600), .Z(n_1145));
	notech_reg Daddrs_reg_14(.CP(n_62311), .D(n_25178), .CD(n_61121), .Q(Daddr
		[14]));
	notech_mux2 i_12551(.S(\nbus_11354[0] ), .A(Daddr[14]), .B(n_20927), .Z(n_25178
		));
	notech_ao3 i_88951129(.A(opc_10[17]), .B(opcode_289113), .C(n_2694), .Z(n_1144
		));
	notech_reg Daddrs_reg_15(.CP(n_62311), .D(n_25188), .CD(n_61121), .Q(Daddr
		[15]));
	notech_mux2 i_12559(.S(\nbus_11354[0] ), .A(Daddr[15]), .B(n_20933), .Z(n_25188
		));
	notech_nor2 i_88551133(.A(n_2648), .B(n_2674), .Z(n_1143));
	notech_reg Daddrs_reg_16(.CP(n_62311), .D(n_25194), .CD(n_61121), .Q(Daddr
		[16]));
	notech_mux2 i_12567(.S(n_54785), .A(Daddr[16]), .B(n_20939), .Z(n_25194)
		);
	notech_or2 i_88451134(.A(n_2672), .B(n_58978), .Z(n_1142));
	notech_reg Daddrs_reg_17(.CP(n_62311), .D(n_25203), .CD(n_61121), .Q(Daddr
		[17]));
	notech_mux2 i_12575(.S(n_54785), .A(Daddr[17]), .B(n_20945), .Z(n_25203)
		);
	notech_or4 i_88851130(.A(n_56177), .B(n_56163), .C(n_56369), .D(n_27583)
		, .Z(n_1141));
	notech_reg Daddrs_reg_18(.CP(n_62311), .D(n_25211), .CD(n_61121), .Q(Daddr
		[18]));
	notech_mux2 i_12583(.S(n_54785), .A(Daddr[18]), .B(n_20951), .Z(n_25211)
		);
	notech_and2 i_88251136(.A(\regs_13_14[17] ), .B(n_2652), .Z(n_1140));
	notech_reg Daddrs_reg_19(.CP(n_62311), .D(n_25225), .CD(n_61123), .Q(Daddr
		[19]));
	notech_mux2 i_12591(.S(n_54785), .A(Daddr[19]), .B(n_20957), .Z(n_25225)
		);
	notech_reg Daddrs_reg_20(.CP(n_62311), .D(n_25231), .CD(n_61123), .Q(Daddr
		[20]));
	notech_mux2 i_12599(.S(n_54785), .A(Daddr[20]), .B(n_20963), .Z(n_25231)
		);
	notech_reg Daddrs_reg_21(.CP(n_62311), .D(n_25240), .CD(n_61123), .Q(Daddr
		[21]));
	notech_mux2 i_12607(.S(n_54785), .A(Daddr[21]), .B(n_20969), .Z(n_25240)
		);
	notech_or4 i_86151155(.A(n_60752), .B(n_60739), .C(n_60768), .D(n_2693),
		 .Z(n_1137));
	notech_reg Daddrs_reg_22(.CP(n_62311), .D(n_25246), .CD(n_61123), .Q(Daddr
		[22]));
	notech_mux2 i_12615(.S(n_54785), .A(Daddr[22]), .B(n_20975), .Z(n_25246)
		);
	notech_reg Daddrs_reg_23(.CP(n_62227), .D(n_25252), .CD(n_61121), .Q(Daddr
		[23]));
	notech_mux2 i_12623(.S(n_54785), .A(Daddr[23]), .B(n_20981), .Z(n_25252)
		);
	notech_nand3 i_177057859(.A(calc_sz[0]), .B(n_205888855), .C(n_2041), .Z
		(n_1135));
	notech_reg Daddrs_reg_24(.CP(n_62227), .D(n_25258), .CD(n_61121), .Q(Daddr
		[24]));
	notech_mux2 i_12631(.S(n_54785), .A(Daddr[24]), .B(n_20987), .Z(n_25258)
		);
	notech_reg Daddrs_reg_25(.CP(n_62315), .D(n_25264), .CD(n_61120), .Q(Daddr
		[25]));
	notech_mux2 i_12639(.S(n_54785), .A(Daddr[25]), .B(n_20993), .Z(n_25264)
		);
	notech_reg Daddrs_reg_26(.CP(n_62229), .D(n_25270), .CD(n_61120), .Q(Daddr
		[26]));
	notech_mux2 i_12647(.S(n_54785), .A(Daddr[26]), .B(n_20999), .Z(n_25270)
		);
	notech_reg Daddrs_reg_27(.CP(n_62229), .D(n_25276), .CD(n_61121), .Q(Daddr
		[27]));
	notech_mux2 i_12655(.S(n_54785), .A(Daddr[27]), .B(n_21005), .Z(n_25276)
		);
	notech_reg Daddrs_reg_28(.CP(n_62229), .D(n_25282), .CD(n_61121), .Q(Daddr
		[28]));
	notech_mux2 i_12663(.S(n_54785), .A(Daddr[28]), .B(n_21011), .Z(n_25282)
		);
	notech_reg Daddrs_reg_29(.CP(n_62229), .D(n_25288), .CD(n_61121), .Q(Daddr
		[29]));
	notech_mux2 i_12671(.S(n_54785), .A(Daddr[29]), .B(n_21017), .Z(n_25288)
		);
	notech_reg Daddrs_reg_30(.CP(n_62229), .D(n_25294), .CD(n_61121), .Q(Daddr
		[30]));
	notech_mux2 i_12679(.S(n_54785), .A(Daddr[30]), .B(n_21023), .Z(n_25294)
		);
	notech_reg Daddrs_reg_31(.CP(n_62229), .D(n_25300), .CD(n_61121), .Q(Daddr
		[31]));
	notech_mux2 i_12687(.S(n_54785), .A(Daddr[31]), .B(n_21029), .Z(n_25300)
		);
	notech_reg read_req_reg(.CP(n_62229), .D(n_25307), .CD(n_61126), .Q(read_reqs
		));
	notech_mux2 i_12695(.S(n_18922), .A(read_reqs), .B(n_27296), .Z(n_25307)
		);
	notech_reg_set temp_ss_reg_0(.CP(n_62229), .D(n_25313), .SD(1'b1), .Q(temp_ss
		[0]));
	notech_mux2 i_12703(.S(\nbus_11327[0] ), .A(temp_ss[0]), .B(n_248085800)
		, .Z(n_25313));
	notech_reg_set temp_ss_reg_1(.CP(n_62229), .D(n_25319), .SD(1'b1), .Q(temp_ss
		[1]));
	notech_mux2 i_12711(.S(\nbus_11327[0] ), .A(temp_ss[1]), .B(n_248185801)
		, .Z(n_25319));
	notech_reg_set temp_ss_reg_2(.CP(n_62315), .D(n_25326), .SD(1'b1), .Q(temp_ss
		[2]));
	notech_mux2 i_12721(.S(\nbus_11327[0] ), .A(temp_ss[2]), .B(n_248285802)
		, .Z(n_25326));
	notech_reg_set temp_ss_reg_3(.CP(n_62315), .D(n_25334), .SD(1'b1), .Q(temp_ss
		[3]));
	notech_mux2 i_12729(.S(\nbus_11327[0] ), .A(temp_ss[3]), .B(n_248385803)
		, .Z(n_25334));
	notech_reg_set temp_ss_reg_4(.CP(n_62315), .D(n_25340), .SD(1'b1), .Q(temp_ss
		[4]));
	notech_mux2 i_12737(.S(\nbus_11327[0] ), .A(temp_ss[4]), .B(n_248485804)
		, .Z(n_25340));
	notech_reg_set temp_ss_reg_5(.CP(n_62315), .D(n_25346), .SD(1'b1), .Q(temp_ss
		[5]));
	notech_mux2 i_12745(.S(\nbus_11327[0] ), .A(temp_ss[5]), .B(n_248585805)
		, .Z(n_25346));
	notech_reg_set temp_ss_reg_6(.CP(n_62315), .D(n_25352), .SD(1'b1), .Q(temp_ss
		[6]));
	notech_mux2 i_12753(.S(\nbus_11327[0] ), .A(temp_ss[6]), .B(n_248685806)
		, .Z(n_25352));
	notech_reg_set temp_ss_reg_7(.CP(n_62315), .D(n_25358), .SD(1'b1), .Q(temp_ss
		[7]));
	notech_mux2 i_12761(.S(\nbus_11327[0] ), .A(temp_ss[7]), .B(n_248785807)
		, .Z(n_25358));
	notech_reg_set temp_ss_reg_8(.CP(n_62315), .D(n_25366), .SD(1'b1), .Q(temp_ss
		[8]));
	notech_mux2 i_12769(.S(\nbus_11327[0] ), .A(temp_ss[8]), .B(n_248885808)
		, .Z(n_25366));
	notech_nand3 i_820627(.A(n_1213), .B(n_1210), .C(n_1221), .Z(n_20153));
	notech_reg_set temp_ss_reg_9(.CP(n_62315), .D(n_25373), .SD(1'b1), .Q(temp_ss
		[9]));
	notech_mux2 i_12777(.S(\nbus_11327[0] ), .A(temp_ss[9]), .B(n_248985809)
		, .Z(n_25373));
	notech_reg_set temp_ss_reg_10(.CP(n_62315), .D(n_25379), .SD(1'b1), .Q(temp_ss
		[10]));
	notech_mux2 i_12785(.S(\nbus_11327[0] ), .A(temp_ss[10]), .B(n_249085810
		), .Z(n_25379));
	notech_reg_set temp_ss_reg_11(.CP(n_62315), .D(n_25385), .SD(1'b1), .Q(temp_ss
		[11]));
	notech_mux2 i_12793(.S(\nbus_11327[0] ), .A(temp_ss[11]), .B(n_249185811
		), .Z(n_25385));
	notech_nand2 i_62151380(.A(opa[7]), .B(n_2692), .Z(n_1115));
	notech_reg_set temp_ss_reg_12(.CP(n_62315), .D(n_25391), .SD(1'b1), .Q(temp_ss
		[12]));
	notech_mux2 i_12801(.S(\nbus_11327[0] ), .A(temp_ss[12]), .B(n_249285812
		), .Z(n_25391));
	notech_reg_set temp_ss_reg_13(.CP(n_62315), .D(n_25397), .SD(1'b1), .Q(temp_ss
		[13]));
	notech_mux2 i_12809(.S(\nbus_11327[0] ), .A(temp_ss[13]), .B(n_249385813
		), .Z(n_25397));
	notech_reg_set temp_ss_reg_14(.CP(n_62315), .D(n_25403), .SD(1'b1), .Q(temp_ss
		[14]));
	notech_mux2 i_12817(.S(\nbus_11327[0] ), .A(temp_ss[14]), .B(n_249485814
		), .Z(n_25403));
	notech_nao3 i_62351378(.A(opc_10[7]), .B(opcode_289113), .C(n_54526258),
		 .Z(n_1112));
	notech_reg_set temp_ss_reg_15(.CP(n_62315), .D(n_25409), .SD(1'b1), .Q(temp_ss
		[15]));
	notech_mux2 i_12825(.S(\nbus_11327[0] ), .A(temp_ss[15]), .B(n_249585815
		), .Z(n_25409));
	notech_nand2 i_61851383(.A(n_2676), .B(n_55819), .Z(n_1111));
	notech_reg_set temp_ss_reg_16(.CP(n_62315), .D(n_25415), .SD(1'b1), .Q(temp_ss
		[16]));
	notech_mux2 i_12833(.S(n_52529), .A(temp_ss[16]), .B(n_249685816), .Z(n_25415
		));
	notech_nand2 i_61651385(.A(sav_epc[7]), .B(n_60584), .Z(n_1110));
	notech_reg_set temp_ss_reg_17(.CP(n_62315), .D(n_25421), .SD(1'b1), .Q(temp_ss
		[17]));
	notech_mux2 i_12841(.S(n_52529), .A(temp_ss[17]), .B(n_249785817), .Z(n_25421
		));
	notech_reg_set temp_ss_reg_18(.CP(n_62315), .D(n_25427), .SD(1'b1), .Q(temp_ss
		[18]));
	notech_mux2 i_12849(.S(n_52529), .A(temp_ss[18]), .B(n_249885818), .Z(n_25427
		));
	notech_reg_set temp_ss_reg_19(.CP(n_62315), .D(n_25433), .SD(1'b1), .Q(temp_ss
		[19]));
	notech_mux2 i_12857(.S(n_52529), .A(temp_ss[19]), .B(n_249985819), .Z(n_25433
		));
	notech_reg_set temp_ss_reg_20(.CP(n_62229), .D(n_25439), .SD(1'b1), .Q(temp_ss
		[20]));
	notech_mux2 i_12865(.S(n_52529), .A(temp_ss[20]), .B(n_250085820), .Z(n_25439
		));
	notech_reg_set temp_ss_reg_21(.CP(n_62229), .D(n_25445), .SD(1'b1), .Q(temp_ss
		[21]));
	notech_mux2 i_12873(.S(n_52529), .A(temp_ss[21]), .B(n_250185821), .Z(n_25445
		));
	notech_and4 i_60751391(.A(n_55846), .B(n_1963), .C(n_55834), .D(n_55833)
		, .Z(n_1105));
	notech_reg_set temp_ss_reg_22(.CP(n_62231), .D(n_25451), .SD(1'b1), .Q(temp_ss
		[22]));
	notech_mux2 i_12881(.S(n_52529), .A(temp_ss[22]), .B(n_250285822), .Z(n_25451
		));
	notech_and3 i_55251442(.A(n_55667), .B(n_1079), .C(n_54668), .Z(n_1104)
		);
	notech_reg_set temp_ss_reg_23(.CP(n_62231), .D(n_25457), .SD(1'b1), .Q(temp_ss
		[23]));
	notech_mux2 i_12889(.S(n_52529), .A(temp_ss[23]), .B(n_250385823), .Z(n_25457
		));
	notech_reg_set temp_ss_reg_24(.CP(n_62231), .D(n_25463), .SD(1'b1), .Q(temp_ss
		[24]));
	notech_mux2 i_12897(.S(n_52529), .A(temp_ss[24]), .B(n_250485824), .Z(n_25463
		));
	notech_reg_set temp_ss_reg_25(.CP(n_62231), .D(n_25469), .SD(1'b1), .Q(temp_ss
		[25]));
	notech_mux2 i_12905(.S(n_52529), .A(temp_ss[25]), .B(n_250585825), .Z(n_25469
		));
	notech_reg_set temp_ss_reg_26(.CP(n_62231), .D(n_25475), .SD(1'b1), .Q(temp_ss
		[26]));
	notech_mux2 i_12913(.S(n_52529), .A(temp_ss[26]), .B(n_250685826), .Z(n_25475
		));
	notech_reg_set temp_ss_reg_27(.CP(n_62231), .D(n_25481), .SD(1'b1), .Q(temp_ss
		[27]));
	notech_mux2 i_12921(.S(n_52529), .A(temp_ss[27]), .B(n_250785827), .Z(n_25481
		));
	notech_reg_set temp_ss_reg_28(.CP(n_62231), .D(n_25487), .SD(1'b1), .Q(temp_ss
		[28]));
	notech_mux2 i_12929(.S(n_52529), .A(temp_ss[28]), .B(n_250885828), .Z(n_25487
		));
	notech_reg_set temp_ss_reg_29(.CP(n_62231), .D(n_25493), .SD(1'b1), .Q(temp_ss
		[29]));
	notech_mux2 i_12937(.S(n_52529), .A(temp_ss[29]), .B(n_250985829), .Z(n_25493
		));
	notech_reg_set temp_ss_reg_30(.CP(n_62231), .D(n_25499), .SD(1'b1), .Q(temp_ss
		[30]));
	notech_mux2 i_12945(.S(n_52529), .A(temp_ss[30]), .B(n_251085830), .Z(n_25499
		));
	notech_reg_set temp_ss_reg_31(.CP(n_62231), .D(n_25505), .SD(1'b1), .Q(temp_ss
		[31]));
	notech_mux2 i_12953(.S(n_52529), .A(temp_ss[31]), .B(n_251185831), .Z(n_25505
		));
	notech_reg errco_reg_0(.CP(n_62231), .D(n_25511), .CD(n_61133), .Q(errco
		[0]));
	notech_mux2 i_12961(.S(n_53864), .A(errco[0]), .B(n_67587010), .Z(n_25511
		));
	notech_reg errco_reg_1(.CP(n_62231), .D(n_25517), .CD(n_61133), .Q(errco
		[1]));
	notech_mux2 i_12969(.S(n_53864), .A(errco[1]), .B(wr_fault), .Z(n_25517)
		);
	notech_reg errco_reg_2(.CP(n_62231), .D(n_25523), .CD(n_61133), .Q(errco
		[2]));
	notech_mux2 i_12977(.S(n_53864), .A(errco[2]), .B(cs[1]), .Z(n_25523));
	notech_reg errco_reg_3(.CP(n_62231), .D(n_25532), .CD(n_61133), .Q(errco
		[3]));
	notech_ao3 i_12987(.A(n_59183), .B(errco[3]), .C(n_60415), .Z(n_25532)
		);
	notech_reg errco_reg_4(.CP(n_62231), .D(n_25535), .CD(n_61133), .Q(errco
		[4]));
	notech_mux2 i_12993(.S(n_53864), .A(errco[4]), .B(n_60415), .Z(n_25535)
		);
	notech_reg errco_reg_5(.CP(n_62231), .D(n_25544), .CD(n_61135), .Q(errco
		[5]));
	notech_ao3 i_13005(.A(n_59183), .B(errco[5]), .C(n_60415), .Z(n_25544)
		);
	notech_reg errco_reg_6(.CP(n_62231), .D(n_25550), .CD(n_61135), .Q(errco
		[6]));
	notech_ao3 i_13013(.A(n_59181), .B(errco[6]), .C(n_60423), .Z(n_25550)
		);
	notech_reg errco_reg_7(.CP(n_62231), .D(n_25557), .CD(n_61133), .Q(errco
		[7]));
	notech_ao3 i_13021(.A(n_59179), .B(errco[7]), .C(n_60415), .Z(n_25557)
		);
	notech_reg errco_reg_8(.CP(n_62231), .D(n_25566), .CD(n_61133), .Q(errco
		[8]));
	notech_ao3 i_13029(.A(n_59179), .B(errco[8]), .C(n_60415), .Z(n_25566)
		);
	notech_reg errco_reg_9(.CP(n_62165), .D(n_25574), .CD(n_61132), .Q(errco
		[9]));
	notech_ao3 i_13037(.A(n_59179), .B(errco[9]), .C(n_60415), .Z(n_25574)
		);
	notech_and3 i_27551702(.A(n_55667), .B(n_2651), .C(n_1073), .Z(n_1085)
		);
	notech_reg errco_reg_10(.CP(n_62165), .D(n_25584), .CD(n_61133), .Q(errco
		[10]));
	notech_ao3 i_13045(.A(n_59179), .B(errco[10]), .C(n_60415), .Z(n_25584)
		);
	notech_or2 i_27351704(.A(n_55580), .B(n_56144), .Z(n_1084));
	notech_reg errco_reg_11(.CP(n_62165), .D(n_25590), .CD(n_61132), .Q(errco
		[11]));
	notech_ao3 i_13053(.A(n_59179), .B(errco[11]), .C(n_60415), .Z(n_25590)
		);
	notech_or2 i_23951735(.A(n_56027), .B(n_2658), .Z(n_1083));
	notech_reg errco_reg_12(.CP(n_62165), .D(n_25596), .CD(n_61132), .Q(errco
		[12]));
	notech_ao3 i_13061(.A(n_59179), .B(errco[12]), .C(n_60415), .Z(n_25596)
		);
	notech_and3 i_180952006(.A(n_55658), .B(n_1081), .C(n_56029), .Z(n_54668
		));
	notech_reg errco_reg_13(.CP(n_62165), .D(n_25602), .CD(n_61133), .Q(errco
		[13]));
	notech_ao3 i_13069(.A(n_59179), .B(errco[13]), .C(n_60415), .Z(n_25602)
		);
	notech_or4 i_23651738(.A(n_2740), .B(n_1076), .C(n_54668), .D(n_60527), 
		.Z(n_1082));
	notech_reg errco_reg_14(.CP(n_62165), .D(n_25609), .CD(n_61133), .Q(errco
		[14]));
	notech_ao3 i_13077(.A(n_59179), .B(errco[14]), .C(n_60415), .Z(n_25609)
		);
	notech_or2 i_23351741(.A(n_56063), .B(n_26227), .Z(n_1081));
	notech_reg errco_reg_15(.CP(n_62165), .D(n_25615), .CD(n_61133), .Q(errco
		[15]));
	notech_ao3 i_13085(.A(n_59179), .B(errco[15]), .C(n_60415), .Z(n_25615)
		);
	notech_reg errco_reg_16(.CP(n_62165), .D(n_25621), .CD(n_61133), .Q(errco
		[16]));
	notech_ao3 i_13093(.A(n_59179), .B(errco[16]), .C(n_60415), .Z(n_25621)
		);
	notech_or2 i_21651757(.A(n_55858), .B(n_26227), .Z(n_1079));
	notech_reg errco_reg_17(.CP(n_62165), .D(n_25627), .CD(n_61133), .Q(errco
		[17]));
	notech_ao3 i_13101(.A(n_59179), .B(errco[17]), .C(n_60423), .Z(n_25627)
		);
	notech_reg errco_reg_18(.CP(n_62077), .D(n_25633), .CD(n_61135), .Q(errco
		[18]));
	notech_ao3 i_13109(.A(n_59179), .B(errco[18]), .C(n_60419), .Z(n_25633)
		);
	notech_nand3 i_20151772(.A(n_62409), .B(n_59375), .C(n_2689), .Z(n_1077)
		);
	notech_reg errco_reg_19(.CP(n_62165), .D(n_25639), .CD(n_61136), .Q(errco
		[19]));
	notech_ao3 i_13117(.A(n_59179), .B(errco[19]), .C(n_60419), .Z(n_25639)
		);
	notech_ao4 i_84051981(.A(n_59375), .B(opcode_289113), .C(n_2264), .D(n_26807
		), .Z(n_1076));
	notech_reg errco_reg_20(.CP(n_62263), .D(n_25645), .CD(n_61136), .Q(errco
		[20]));
	notech_ao3 i_13125(.A(n_59181), .B(errco[20]), .C(n_60419), .Z(n_25645)
		);
	notech_or2 i_20251771(.A(n_1076), .B(n_26315), .Z(n_1075));
	notech_reg errco_reg_21(.CP(n_62119), .D(n_25651), .CD(n_61135), .Q(errco
		[21]));
	notech_ao3 i_13133(.A(n_59181), .B(errco[21]), .C(n_60419), .Z(n_25651)
		);
	notech_reg errco_reg_22(.CP(n_62119), .D(n_25657), .CD(n_61136), .Q(errco
		[22]));
	notech_ao3 i_13141(.A(n_59181), .B(errco[22]), .C(n_60419), .Z(n_25657)
		);
	notech_or4 i_200352024(.A(n_1909), .B(n_1069), .C(n_59230), .D(n_60516),
		 .Z(n_54508));
	notech_reg errco_reg_23(.CP(n_62119), .D(n_25663), .CD(n_61136), .Q(errco
		[23]));
	notech_ao3 i_13149(.A(n_59181), .B(errco[23]), .C(n_60419), .Z(n_25663)
		);
	notech_and2 i_36352022(.A(n_55667), .B(n_1073), .Z(n_55986));
	notech_reg errco_reg_24(.CP(n_62191), .D(n_25670), .CD(n_61136), .Q(errco
		[24]));
	notech_ao3 i_13157(.A(n_59181), .B(errco[24]), .C(n_60419), .Z(n_25670)
		);
	notech_or2 i_18251791(.A(n_55858), .B(n_26574), .Z(n_1073));
	notech_reg errco_reg_25(.CP(n_62191), .D(n_25677), .CD(n_61136), .Q(errco
		[25]));
	notech_ao3 i_13165(.A(n_59181), .B(errco[25]), .C(n_60419), .Z(n_25677)
		);
	notech_reg errco_reg_26(.CP(n_62191), .D(n_25683), .CD(n_61136), .Q(errco
		[26]));
	notech_ao3 i_13173(.A(n_59181), .B(errco[26]), .C(n_60423), .Z(n_25683)
		);
	notech_or2 i_17951794(.A(n_55827), .B(n_26574), .Z(n_1071));
	notech_reg errco_reg_27(.CP(n_62191), .D(n_25689), .CD(n_61136), .Q(errco
		[27]));
	notech_ao3 i_13181(.A(n_59181), .B(errco[27]), .C(n_60423), .Z(n_25689)
		);
	notech_nand3 i_17551798(.A(n_62409), .B(n_59375), .C(n_56101), .Z(n_1070
		));
	notech_reg errco_reg_28(.CP(n_62191), .D(n_25695), .CD(n_61135), .Q(errco
		[28]));
	notech_ao3 i_13190(.A(n_59181), .B(errco[28]), .C(n_60423), .Z(n_25695)
		);
	notech_ao4 i_180551966(.A(n_59375), .B(opcode_289113), .C(n_2264), .D(n_26550
		), .Z(n_1069));
	notech_reg errco_reg_29(.CP(n_62191), .D(n_25701), .CD(n_61135), .Q(errco
		[29]));
	notech_ao3 i_13198(.A(n_59181), .B(errco[29]), .C(n_60423), .Z(n_25701)
		);
	notech_nand2 i_17651797(.A(n_56305), .B(n_28932), .Z(n_1068));
	notech_reg errco_reg_30(.CP(n_62191), .D(n_25707), .CD(n_61135), .Q(errco
		[30]));
	notech_ao3 i_13206(.A(n_59181), .B(errco[30]), .C(n_60419), .Z(n_25707)
		);
	notech_reg errco_reg_31(.CP(n_62191), .D(n_25713), .CD(n_61135), .Q(errco
		[31]));
	notech_ao3 i_13214(.A(n_59181), .B(errco[31]), .C(n_60419), .Z(n_25713)
		);
	notech_reg_set write_data_reg_0(.CP(n_62191), .D(n_25716), .SD(1'b1), .Q
		(write_data[0]));
	notech_mux2 i_13221(.S(n_27366), .A(write_data[0]), .B(n_18256), .Z(n_25716
		));
	notech_reg_set write_data_reg_1(.CP(n_62191), .D(n_25722), .SD(1'b1), .Q
		(write_data[1]));
	notech_mux2 i_13229(.S(n_27366), .A(write_data[1]), .B(n_18261), .Z(n_25722
		));
	notech_reg_set write_data_reg_2(.CP(n_62191), .D(n_25728), .SD(1'b1), .Q
		(write_data[2]));
	notech_mux2 i_13238(.S(n_27366), .A(write_data[2]), .B(n_18266), .Z(n_25728
		));
	notech_reg_set write_data_reg_3(.CP(n_62191), .D(n_25736), .SD(1'b1), .Q
		(write_data[3]));
	notech_mux2 i_13246(.S(n_27366), .A(write_data[3]), .B(n_18271), .Z(n_25736
		));
	notech_reg_set write_data_reg_4(.CP(n_62191), .D(n_25742), .SD(1'b1), .Q
		(write_data[4]));
	notech_mux2 i_13254(.S(n_27366), .A(write_data[4]), .B(n_18276), .Z(n_25742
		));
	notech_reg_set write_data_reg_5(.CP(n_62191), .D(n_25748), .SD(1'b1), .Q
		(write_data[5]));
	notech_mux2 i_13263(.S(n_27366), .A(write_data[5]), .B(n_18281), .Z(n_25748
		));
	notech_reg_set write_data_reg_6(.CP(n_62191), .D(n_25754), .SD(1'b1), .Q
		(write_data[6]));
	notech_mux2 i_13271(.S(n_27366), .A(write_data[6]), .B(n_18286), .Z(n_25754
		));
	notech_reg_set write_data_reg_7(.CP(n_62191), .D(n_25760), .SD(1'b1), .Q
		(write_data[7]));
	notech_mux2 i_13279(.S(n_27366), .A(write_data[7]), .B(n_18291), .Z(n_25760
		));
	notech_reg_set write_data_reg_8(.CP(n_62191), .D(n_25766), .SD(1'b1), .Q
		(write_data[8]));
	notech_mux2 i_13287(.S(n_27366), .A(write_data[8]), .B(n_18296), .Z(n_25766
		));
	notech_reg_set write_data_reg_9(.CP(n_62191), .D(n_25772), .SD(1'b1), .Q
		(write_data[9]));
	notech_mux2 i_13295(.S(n_27366), .A(write_data[9]), .B(n_18301), .Z(n_25772
		));
	notech_reg_set write_data_reg_10(.CP(n_62191), .D(n_25778), .SD(1'b1), .Q
		(write_data[10]));
	notech_mux2 i_13303(.S(n_27366), .A(write_data[10]), .B(n_18306), .Z(n_25778
		));
	notech_reg_set write_data_reg_11(.CP(n_62263), .D(n_25784), .SD(1'b1), .Q
		(write_data[11]));
	notech_mux2 i_13311(.S(n_27366), .A(write_data[11]), .B(n_18311), .Z(n_25784
		));
	notech_reg_set write_data_reg_12(.CP(n_62189), .D(n_25790), .SD(1'b1), .Q
		(write_data[12]));
	notech_mux2 i_13319(.S(n_27366), .A(write_data[12]), .B(n_18316), .Z(n_25790
		));
	notech_reg_set write_data_reg_13(.CP(n_62263), .D(n_25796), .SD(1'b1), .Q
		(write_data[13]));
	notech_mux2 i_13327(.S(n_27366), .A(write_data[13]), .B(n_18321), .Z(n_25796
		));
	notech_reg_set write_data_reg_14(.CP(n_62263), .D(n_25802), .SD(1'b1), .Q
		(write_data[14]));
	notech_mux2 i_13335(.S(n_27366), .A(write_data[14]), .B(n_18326), .Z(n_25802
		));
	notech_reg_set write_data_reg_15(.CP(n_62263), .D(n_25808), .SD(1'b1), .Q
		(write_data[15]));
	notech_mux2 i_13343(.S(n_27366), .A(write_data[15]), .B(n_18331), .Z(n_25808
		));
	notech_reg_set write_data_reg_16(.CP(n_62263), .D(n_25814), .SD(1'b1), .Q
		(write_data[16]));
	notech_mux2 i_13351(.S(n_53351), .A(write_data[16]), .B(n_18336), .Z(n_25814
		));
	notech_reg_set write_data_reg_17(.CP(n_62263), .D(n_25820), .SD(1'b1), .Q
		(write_data[17]));
	notech_mux2 i_13359(.S(n_53351), .A(write_data[17]), .B(n_18341), .Z(n_25820
		));
	notech_ao4 i_171556243(.A(n_2263), .B(n_26821), .C(n_1023), .D(n_26319),
		 .Z(n_1048));
	notech_reg_set write_data_reg_18(.CP(n_62263), .D(n_25826), .SD(1'b1), .Q
		(write_data[18]));
	notech_mux2 i_13367(.S(n_53351), .A(write_data[18]), .B(n_18346), .Z(n_25826
		));
	notech_reg_set write_data_reg_19(.CP(n_62263), .D(n_25832), .SD(1'b1), .Q
		(write_data[19]));
	notech_mux2 i_13375(.S(n_53351), .A(write_data[19]), .B(n_18351), .Z(n_25832
		));
	notech_ao4 i_171956239(.A(n_26591), .B(n_27019), .C(n_26230), .D(n_26189
		), .Z(n_1046));
	notech_reg_set write_data_reg_20(.CP(n_62263), .D(n_25838), .SD(1'b1), .Q
		(write_data[20]));
	notech_mux2 i_13383(.S(n_53351), .A(write_data[20]), .B(n_18356), .Z(n_25838
		));
	notech_reg_set write_data_reg_21(.CP(n_62263), .D(n_25846), .SD(1'b1), .Q
		(write_data[21]));
	notech_mux2 i_13391(.S(n_53351), .A(write_data[21]), .B(n_18361), .Z(n_25846
		));
	notech_ao4 i_172256236(.A(n_55959), .B(n_54505), .C(n_254834174), .D(eval_flag
		), .Z(n_1044));
	notech_reg_set write_data_reg_22(.CP(n_62263), .D(n_25854), .SD(1'b1), .Q
		(write_data[22]));
	notech_mux2 i_13399(.S(n_53351), .A(write_data[22]), .B(n_18366), .Z(n_25854
		));
	notech_reg_set write_data_reg_23(.CP(n_62263), .D(n_25860), .SD(1'b1), .Q
		(write_data[23]));
	notech_mux2 i_13407(.S(n_53351), .A(write_data[23]), .B(n_18371), .Z(n_25860
		));
	notech_reg_set write_data_reg_24(.CP(n_62263), .D(n_25879), .SD(1'b1), .Q
		(write_data[24]));
	notech_mux2 i_13415(.S(n_53351), .A(write_data[24]), .B(n_18376), .Z(n_25879
		));
	notech_or4 i_28522(.A(n_60752), .B(n_60739), .C(n_60768), .D(n_59369), .Z
		(n_1041));
	notech_reg_set write_data_reg_25(.CP(n_62263), .D(n_25892), .SD(1'b1), .Q
		(write_data[25]));
	notech_mux2 i_13423(.S(n_53351), .A(write_data[25]), .B(n_18381), .Z(n_25892
		));
	notech_or2 i_92456993(.A(n_55807), .B(n_55952), .Z(n_1040));
	notech_reg_set write_data_reg_26(.CP(n_62263), .D(n_25898), .SD(1'b1), .Q
		(write_data[26]));
	notech_mux2 i_13431(.S(n_53351), .A(write_data[26]), .B(n_18386), .Z(n_25898
		));
	notech_or4 i_92056997(.A(n_58931), .B(n_59369), .C(n_59899), .D(n_56551)
		, .Z(n_1039));
	notech_reg_set write_data_reg_27(.CP(n_62263), .D(n_25904), .SD(1'b1), .Q
		(write_data[27]));
	notech_mux2 i_13439(.S(n_53351), .A(write_data[27]), .B(n_18391), .Z(n_25904
		));
	notech_reg_set write_data_reg_28(.CP(n_62263), .D(n_25910), .SD(1'b1), .Q
		(write_data[28]));
	notech_mux2 i_13447(.S(n_53351), .A(write_data[28]), .B(n_18396), .Z(n_25910
		));
	notech_reg_set write_data_reg_29(.CP(n_62263), .D(n_25916), .SD(1'b1), .Q
		(write_data[29]));
	notech_mux2 i_13455(.S(n_53351), .A(write_data[29]), .B(n_18401), .Z(n_25916
		));
	notech_reg_set write_data_reg_30(.CP(n_62119), .D(n_25922), .SD(1'b1), .Q
		(write_data[30]));
	notech_mux2 i_13463(.S(n_53351), .A(write_data[30]), .B(n_18406), .Z(n_25922
		));
	notech_and2 i_91357004(.A(n_54953), .B(n_35829), .Z(n_1035));
	notech_reg_set write_data_reg_31(.CP(n_62189), .D(n_25928), .SD(1'b1), .Q
		(write_data[31]));
	notech_mux2 i_13471(.S(n_53351), .A(write_data[31]), .B(n_18411), .Z(n_25928
		));
	notech_reg writeio_req_reg(.CP(n_62189), .D(n_25934), .CD(n_61135), .Q(writeio_req
		));
	notech_mux2 i_13479(.S(n_17679), .A(writeio_req), .B(n_59819), .Z(n_25934
		));
	notech_reg write_sz_reg_0(.CP(n_62189), .D(n_25940), .CD(n_61135), .Q(write_sz
		[0]));
	notech_mux2 i_13487(.S(\nbus_11341[0] ), .A(write_sz[0]), .B(n_238885708
		), .Z(n_25940));
	notech_reg_set write_sz_reg_1(.CP(n_62119), .D(n_25946), .SD(n_61135), .Q
		(write_sz[1]));
	notech_mux2 i_13495(.S(\nbus_11341[0] ), .A(write_sz[1]), .B(n_27367), .Z
		(n_25946));
	notech_or4 i_31431(.A(n_58940), .B(n_60602), .C(n_57433), .D(n_273288723
		), .Z(n_1031));
	notech_reg flush_tlb_reg(.CP(n_62189), .D(n_25953), .CD(n_61135), .Q(flush_tlb
		));
	notech_mux2 i_13503(.S(n_17010), .A(flush_tlb), .B(n_59819), .Z(n_25953)
		);
	notech_reg flush_Dtlb_reg(.CP(n_62193), .D(n_25959), .CD(n_61135), .Q(flush_Dtlb
		));
	notech_mux2 i_13511(.S(n_14963), .A(flush_Dtlb), .B(n_238785707), .Z(n_25959
		));
	notech_reg_set terms_reg(.CP(n_62147), .D(n_25965), .SD(n_61132), .Q(terminate
		));
	notech_mux2 i_13519(.S(n_11472), .A(terminate), .B(n_11475), .Z(n_25965)
		);
	notech_reg writeio_data_reg_0(.CP(n_62147), .D(n_25971), .CD(n_61130), .Q
		(writeio_data[0]));
	notech_mux2 i_13527(.S(n_300186321), .A(opa[0]), .B(writeio_data[0]), .Z
		(n_25971));
	notech_ao3 i_93056987(.A(n_26887), .B(n_59819), .C(n_57374), .Z(n_1027)
		);
	notech_reg writeio_data_reg_1(.CP(n_62147), .D(n_25977), .CD(n_61130), .Q
		(writeio_data[1]));
	notech_mux2 i_13535(.S(n_300186321), .A(n_59708), .B(writeio_data[1]), .Z
		(n_25977));
	notech_reg writeio_data_reg_2(.CP(n_62193), .D(n_25983), .CD(n_61130), .Q
		(writeio_data[2]));
	notech_mux2 i_13543(.S(n_300186321), .A(n_59717), .B(writeio_data[2]), .Z
		(n_25983));
	notech_or4 i_23457904(.A(n_56487), .B(n_56478), .C(n_56440), .D(n_28966)
		, .Z(n_1025));
	notech_reg writeio_data_reg_3(.CP(n_62193), .D(n_25989), .CD(n_61130), .Q
		(writeio_data[3]));
	notech_mux2 i_13551(.S(n_300186321), .A(opa[3]), .B(writeio_data[3]), .Z
		(n_25989));
	notech_reg writeio_data_reg_4(.CP(n_62193), .D(n_25995), .CD(n_61130), .Q
		(writeio_data[4]));
	notech_mux2 i_13559(.S(n_300186321), .A(opa[4]), .B(writeio_data[4]), .Z
		(n_25995));
	notech_ao4 i_180157858(.A(n_59375), .B(opcode_289113), .C(n_2264), .D(n_26821
		), .Z(n_1023));
	notech_reg writeio_data_reg_5(.CP(n_62193), .D(n_26001), .CD(n_61130), .Q
		(writeio_data[5]));
	notech_mux2 i_13567(.S(n_300186321), .A(opa[5]), .B(writeio_data[5]), .Z
		(n_26001));
	notech_or2 i_90457012(.A(n_55858), .B(n_26805), .Z(n_1022));
	notech_reg writeio_data_reg_6(.CP(n_62193), .D(n_26007), .CD(n_61131), .Q
		(writeio_data[6]));
	notech_mux2 i_13575(.S(n_300186321), .A(opa[6]), .B(writeio_data[6]), .Z
		(n_26007));
	notech_or2 i_90357013(.A(n_55807), .B(n_26805), .Z(n_1021));
	notech_reg writeio_data_reg_7(.CP(n_62193), .D(n_26013), .CD(n_61130), .Q
		(writeio_data[7]));
	notech_mux2 i_13583(.S(n_300186321), .A(n_59744), .B(writeio_data[7]), .Z
		(n_26013));
	notech_or4 i_89357022(.A(n_26190), .B(n_55524), .C(n_60768), .D(n_60724)
		, .Z(n_1020));
	notech_reg writeio_data_reg_8(.CP(n_62193), .D(n_26019), .CD(n_61130), .Q
		(writeio_data[8]));
	notech_mux2 i_13591(.S(n_300186321), .A(opa[8]), .B(writeio_data[8]), .Z
		(n_26019));
	notech_and3 i_84957066(.A(n_55960), .B(n_55959), .C(n_55961), .Z(n_1019)
		);
	notech_reg writeio_data_reg_9(.CP(n_62193), .D(n_26025), .CD(n_61126), .Q
		(writeio_data[9]));
	notech_mux2 i_13599(.S(n_300186321), .A(opa[9]), .B(writeio_data[9]), .Z
		(n_26025));
	notech_reg writeio_data_reg_10(.CP(n_62193), .D(n_26031), .CD(n_61126), 
		.Q(writeio_data[10]));
	notech_mux2 i_13607(.S(n_300186321), .A(opa[10]), .B(writeio_data[10]), 
		.Z(n_26031));
	notech_or2 i_170257898(.A(n_55524), .B(n_26190), .Z(n_1017));
	notech_reg writeio_data_reg_11(.CP(n_62193), .D(n_26037), .CD(n_61126), 
		.Q(writeio_data[11]));
	notech_mux2 i_13615(.S(n_300186321), .A(opa[11]), .B(writeio_data[11]), 
		.Z(n_26037));
	notech_ao4 i_49157965(.A(n_26782), .B(n_26502), .C(n_26326), .D(n_35829)
		, .Z(n_1016));
	notech_reg writeio_data_reg_12(.CP(n_62193), .D(n_26043), .CD(n_61126), 
		.Q(writeio_data[12]));
	notech_mux2 i_13623(.S(n_300186321), .A(opa[12]), .B(writeio_data[12]), 
		.Z(n_26043));
	notech_reg writeio_data_reg_13(.CP(n_62193), .D(n_26049), .CD(n_61126), 
		.Q(writeio_data[13]));
	notech_mux2 i_13631(.S(n_300186321), .A(opa[13]), .B(writeio_data[13]), 
		.Z(n_26049));
	notech_ao4 i_167959002(.A(n_101413408), .B(n_28977), .C(n_57329), .D(n_101213406
		), .Z(n_1014));
	notech_reg writeio_data_reg_14(.CP(n_62193), .D(n_26055), .CD(n_61130), 
		.Q(writeio_data[14]));
	notech_mux2 i_13639(.S(n_300186321), .A(opa[14]), .B(writeio_data[14]), 
		.Z(n_26055));
	notech_reg writeio_data_reg_15(.CP(n_62193), .D(n_26061), .CD(n_61130), 
		.Q(writeio_data[15]));
	notech_mux2 i_13647(.S(n_59949), .A(opa[15]), .B(writeio_data[15]), .Z(n_26061
		));
	notech_ao4 i_168059001(.A(n_56216), .B(n_55249), .C(n_27552), .D(n_59819
		), .Z(n_1012));
	notech_reg writeio_data_reg_16(.CP(n_62147), .D(n_26067), .CD(n_61130), 
		.Q(writeio_data[16]));
	notech_mux2 i_13655(.S(n_59949), .A(opa[16]), .B(writeio_data[16]), .Z(n_26067
		));
	notech_ao4 i_169658986(.A(n_2263), .B(n_26304), .C(n_997), .D(n_26320), 
		.Z(n_1011));
	notech_reg writeio_data_reg_17(.CP(n_62193), .D(n_26073), .CD(n_61130), 
		.Q(writeio_data[17]));
	notech_mux2 i_13663(.S(n_59949), .A(opa[17]), .B(writeio_data[17]), .Z(n_26073
		));
	notech_reg writeio_data_reg_18(.CP(n_62193), .D(n_26079), .CD(n_61131), 
		.Q(writeio_data[18]));
	notech_mux2 i_13671(.S(n_59949), .A(opa[18]), .B(writeio_data[18]), .Z(n_26079
		));
	notech_reg writeio_data_reg_19(.CP(n_62193), .D(n_26085), .CD(n_61132), 
		.Q(writeio_data[19]));
	notech_mux2 i_13679(.S(n_59949), .A(opa[19]), .B(writeio_data[19]), .Z(n_26085
		));
	notech_reg writeio_data_reg_20(.CP(n_62147), .D(n_26091), .CD(n_61132), 
		.Q(writeio_data[20]));
	notech_mux2 i_13687(.S(n_59949), .A(opa[20]), .B(writeio_data[20]), .Z(n_26091
		));
	notech_reg writeio_data_reg_21(.CP(n_62193), .D(n_26097), .CD(n_61132), 
		.Q(writeio_data[21]));
	notech_mux2 i_13695(.S(n_59949), .A(opa[21]), .B(writeio_data[21]), .Z(n_26097
		));
	notech_or4 i_83459776(.A(n_56538), .B(n_205788856), .C(n_59898), .D(n_56892
		), .Z(n_1006));
	notech_reg writeio_data_reg_22(.CP(n_62147), .D(n_26103), .CD(n_61132), 
		.Q(writeio_data[22]));
	notech_mux2 i_13703(.S(n_59949), .A(opa[22]), .B(writeio_data[22]), .Z(n_26103
		));
	notech_reg writeio_data_reg_23(.CP(n_62147), .D(n_26109), .CD(n_61132), 
		.Q(writeio_data[23]));
	notech_mux2 i_13711(.S(n_59949), .A(opa[23]), .B(writeio_data[23]), .Z(n_26109
		));
	notech_reg writeio_data_reg_24(.CP(n_62147), .D(n_26115), .CD(n_61132), 
		.Q(writeio_data[24]));
	notech_mux2 i_13719(.S(n_59949), .A(opa[24]), .B(writeio_data[24]), .Z(n_26115
		));
	notech_reg writeio_data_reg_25(.CP(n_62147), .D(n_26121), .CD(n_61132), 
		.Q(writeio_data[25]));
	notech_mux2 i_13727(.S(n_59949), .A(opa[25]), .B(writeio_data[25]), .Z(n_26121
		));
	notech_reg writeio_data_reg_26(.CP(n_62147), .D(n_26127), .CD(n_61132), 
		.Q(writeio_data[26]));
	notech_mux2 i_13735(.S(n_300186321), .A(opa[26]), .B(writeio_data[26]), 
		.Z(n_26127));
	notech_reg writeio_data_reg_27(.CP(n_62147), .D(n_26133), .CD(n_61132), 
		.Q(writeio_data[27]));
	notech_mux2 i_13743(.S(n_59949), .A(opa[27]), .B(writeio_data[27]), .Z(n_26133
		));
	notech_reg writeio_data_reg_28(.CP(n_62147), .D(n_26139), .CD(n_61131), 
		.Q(writeio_data[28]));
	notech_mux2 i_13751(.S(n_59949), .A(opa[28]), .B(writeio_data[28]), .Z(n_26139
		));
	notech_reg writeio_data_reg_29(.CP(n_62147), .D(n_26145), .CD(n_61131), 
		.Q(writeio_data[29]));
	notech_mux2 i_13759(.S(n_59949), .A(opa[29]), .B(writeio_data[29]), .Z(n_26145
		));
	notech_reg writeio_data_reg_30(.CP(n_62147), .D(n_26151), .CD(n_61131), 
		.Q(writeio_data[30]));
	notech_mux2 i_13767(.S(n_59949), .A(opa[30]), .B(writeio_data[30]), .Z(n_26151
		));
	notech_ao4 i_180060553(.A(n_59375), .B(opcode_289113), .C(n_2264), .D(n_26304
		), .Z(n_997));
	notech_reg writeio_data_reg_31(.CP(n_62147), .D(n_26157), .CD(n_61131), 
		.Q(writeio_data[31]));
	notech_mux2 i_13775(.S(n_59949), .A(opa[31]), .B(writeio_data[31]), .Z(n_26157
		));
	notech_or2 i_84159769(.A(n_55807), .B(n_26582), .Z(n_996));
	notech_reg write_req_reg(.CP(n_62147), .D(n_26165), .CD(n_61131), .Q(write_reqs
		));
	notech_mux2 i_13783(.S(n_10124), .A(write_reqs), .B(n_27368), .Z(n_26165
		));
	notech_and3 i_82659784(.A(n_316988520), .B(n_320588484), .C(n_317688513)
		, .Z(n_995));
	notech_reg pc_req_reg(.CP(n_62147), .D(n_26171), .CD(n_61131), .Q(pc_req
		));
	notech_mux2 i_13791(.S(n_7558), .A(pc_req), .B(n_59819), .Z(n_26171));
	notech_or4 i_27591(.A(n_60768), .B(n_60724), .C(n_59141), .D(n_60584), .Z
		(n_994));
	notech_reg had_lgjmp_reg(.CP(n_62147), .D(n_26177), .CD(n_61131), .Q(had_lgjmp
		));
	notech_mux2 i_13799(.S(n_300686326), .A(\nbus_14523[31] ), .B(had_lgjmp)
		, .Z(n_26177));
	notech_reg readio_req_reg(.CP(n_62147), .D(n_26183), .CD(n_61131), .Q(readio_req
		));
	notech_mux2 i_13807(.S(n_7511), .A(readio_req), .B(n_59819), .Z(n_26183)
		);
	notech_inv i_29475(.A(n_55959), .Z(n_26189));
	notech_inv i_29476(.A(n_250134127), .Z(n_26190));
	notech_inv i_29477(.A(n_54711), .Z(n_26191));
	notech_inv i_29478(.A(n_193667756), .Z(n_26192));
	notech_inv i_29479(.A(n_193567755), .Z(n_26193));
	notech_inv i_29480(.A(n_238568190), .Z(n_26194));
	notech_inv i_29481(.A(n_192567745), .Z(n_26195));
	notech_inv i_29482(.A(n_239668201), .Z(n_26196));
	notech_inv i_29483(.A(n_192467744), .Z(n_26197));
	notech_inv i_29484(.A(n_241068215), .Z(n_26198));
	notech_inv i_29485(.A(n_242368222), .Z(n_26199));
	notech_inv i_29486(.A(n_243068229), .Z(n_26200));
	notech_inv i_29487(.A(n_250668305), .Z(n_26201));
	notech_inv i_29488(.A(n_186367683), .Z(n_26202));
	notech_inv i_29489(.A(n_2692), .Z(n_26203));
	notech_inv i_29490(.A(n_54949), .Z(n_26204));
	notech_inv i_29491(.A(n_277768576), .Z(n_26205));
	notech_inv i_29492(.A(n_296868767), .Z(n_26206));
	notech_inv i_29493(.A(n_102723014), .Z(n_26207));
	notech_inv i_29494(.A(n_297968778), .Z(n_26208));
	notech_inv i_29495(.A(n_298668785), .Z(n_26209));
	notech_inv i_29496(.A(n_299368792), .Z(n_26210));
	notech_inv i_29497(.A(n_300768806), .Z(n_26211));
	notech_inv i_29498(.A(n_302868827), .Z(n_26212));
	notech_inv i_29499(.A(n_304268841), .Z(n_26213));
	notech_inv i_29500(.A(n_306068859), .Z(n_26214));
	notech_inv i_29501(.A(n_313668935), .Z(n_26215));
	notech_inv i_29502(.A(n_314368942), .Z(n_26216));
	notech_inv i_29503(.A(n_315068949), .Z(n_26217));
	notech_inv i_29504(.A(n_315768956), .Z(n_26218));
	notech_inv i_29505(.A(n_316468963), .Z(n_26219));
	notech_inv i_29506(.A(n_322269021), .Z(n_26220));
	notech_inv i_29507(.A(n_322969028), .Z(n_26221));
	notech_inv i_29508(.A(n_323669035), .Z(n_26222));
	notech_inv i_29509(.A(n_324369042), .Z(n_26223));
	notech_inv i_29510(.A(n_326969068), .Z(n_26224));
	notech_inv i_29511(.A(n_55970), .Z(n_26225));
	notech_inv i_29513(.A(n_58487), .Z(n_26226));
	notech_inv i_29514(.A(n_55879), .Z(n_26227));
	notech_inv i_29515(.A(n_55934), .Z(n_26228));
	notech_inv i_29517(.A(n_2255), .Z(n_26229));
	notech_inv i_29519(.A(n_55961), .Z(n_26230));
	notech_inv i_29520(.A(n_55958), .Z(n_26231));
	notech_inv i_29522(.A(n_349465783), .Z(n_26232));
	notech_inv i_29523(.A(n_342969202), .Z(n_26233));
	notech_inv i_29525(.A(n_343969212), .Z(n_26234));
	notech_inv i_29526(.A(n_54936), .Z(n_26235));
	notech_inv i_29527(.A(n_243964756), .Z(n_26236));
	notech_inv i_29528(.A(n_352765816), .Z(n_26237));
	notech_inv i_29529(.A(n_212964463), .Z(n_26238));
	notech_inv i_29530(.A(n_351065799), .Z(n_26239));
	notech_inv i_29531(.A(n_185167671), .Z(n_26240));
	notech_inv i_29532(.A(n_324669045), .Z(n_26241));
	notech_inv i_29533(.A(n_55952), .Z(n_26242));
	notech_inv i_29534(.A(n_2192), .Z(n_26243));
	notech_inv i_29535(.A(n_337765679), .Z(n_26244));
	notech_inv i_29536(.A(n_337865680), .Z(n_26245));
	notech_inv i_29537(.A(n_250334129), .Z(n_26246));
	notech_inv i_29538(.A(n_239168196), .Z(n_26247));
	notech_inv i_29539(.A(n_56032), .Z(n_26248));
	notech_inv i_29540(.A(n_313168930), .Z(n_26249));
	notech_inv i_29541(.A(n_56009), .Z(n_26250));
	notech_inv i_29542(.A(n_56100), .Z(n_26251));
	notech_inv i_29543(.A(n_134170660), .Z(n_26252));
	notech_inv i_29544(.A(n_134570664), .Z(n_26253));
	notech_inv i_29545(.A(n_135470673), .Z(n_26254));
	notech_inv i_29546(.A(n_137670695), .Z(n_26255));
	notech_inv i_29547(.A(n_155270871), .Z(n_26256));
	notech_inv i_29548(.A(n_155970878), .Z(n_26257));
	notech_inv i_29549(.A(n_156670885), .Z(n_26258));
	notech_inv i_29550(.A(n_157770896), .Z(n_26259));
	notech_inv i_29551(.A(n_157970898), .Z(n_26260));
	notech_inv i_29552(.A(n_158170900), .Z(n_26261));
	notech_inv i_29553(.A(n_158570904), .Z(n_26262));
	notech_inv i_29554(.A(n_158770906), .Z(n_26263));
	notech_inv i_29555(.A(n_158970908), .Z(n_26264));
	notech_inv i_29556(.A(n_159370912), .Z(n_26265));
	notech_inv i_29557(.A(n_159570914), .Z(n_26266));
	notech_inv i_29558(.A(n_159770916), .Z(n_26268));
	notech_inv i_29559(.A(n_162070939), .Z(n_26269));
	notech_inv i_29560(.A(n_162770946), .Z(n_26270));
	notech_inv i_29561(.A(n_163470953), .Z(n_26271));
	notech_inv i_29562(.A(n_174471063), .Z(n_26272));
	notech_inv i_29563(.A(n_175171070), .Z(n_26273));
	notech_inv i_29564(.A(n_175871077), .Z(n_26274));
	notech_inv i_29565(.A(n_176571084), .Z(n_26275));
	notech_inv i_29566(.A(n_177271091), .Z(n_26276));
	notech_inv i_29567(.A(n_55988), .Z(n_26277));
	notech_inv i_29568(.A(n_183571146), .Z(n_26278));
	notech_inv i_29569(.A(n_186771178), .Z(n_26279));
	notech_inv i_29570(.A(n_187471185), .Z(n_26280));
	notech_inv i_29571(.A(n_326546823), .Z(n_26281));
	notech_inv i_29572(.A(n_326246826), .Z(n_26282));
	notech_inv i_29573(.A(n_326046828), .Z(n_26283));
	notech_inv i_29574(.A(n_3290), .Z(n_26284));
	notech_inv i_29575(.A(n_327646812), .Z(n_26285));
	notech_inv i_29576(.A(n_327446814), .Z(n_26286));
	notech_inv i_29577(.A(n_57177), .Z(n_26287));
	notech_inv i_29578(.A(n_2783), .Z(n_26288));
	notech_inv i_29579(.A(n_194271253), .Z(n_26289));
	notech_inv i_29580(.A(n_56067), .Z(n_26290));
	notech_inv i_29581(.A(n_55154), .Z(n_26291));
	notech_inv i_29582(.A(n_280472115), .Z(n_26292));
	notech_inv i_29583(.A(n_57399), .Z(n_26293));
	notech_inv i_29584(.A(n_57412), .Z(n_26294));
	notech_inv i_29585(.A(n_57410), .Z(n_26295));
	notech_inv i_29586(.A(n_274788710), .Z(n_26296));
	notech_inv i_29587(.A(n_275965076), .Z(n_26297));
	notech_inv i_29588(.A(n_275265069), .Z(n_26298));
	notech_inv i_29589(.A(n_273665053), .Z(n_26299));
	notech_inv i_29590(.A(n_239864717), .Z(n_26300));
	notech_inv i_29591(.A(n_234864667), .Z(n_26301));
	notech_inv i_29592(.A(n_233764656), .Z(n_26302));
	notech_inv i_29593(.A(n_229464617), .Z(n_26303));
	notech_inv i_29594(.A(n_263436789), .Z(n_26304));
	notech_inv i_29595(.A(n_56000), .Z(n_26305));
	notech_inv i_29596(.A(n_323588455), .Z(n_26306));
	notech_inv i_29597(.A(n_54665), .Z(n_26307));
	notech_inv i_29598(.A(n_173971058), .Z(n_26308));
	notech_inv i_29599(.A(n_55114), .Z(n_26309));
	notech_inv i_29601(.A(n_203164366), .Z(n_26310));
	notech_inv i_29602(.A(n_202264357), .Z(n_26311));
	notech_inv i_29603(.A(n_55972), .Z(n_26312));
	notech_inv i_29604(.A(n_56246), .Z(n_26313));
	notech_inv i_29605(.A(n_56235), .Z(n_26314));
	notech_inv i_29606(.A(n_57358), .Z(n_26315));
	notech_inv i_29607(.A(n_56226), .Z(n_26316));
	notech_inv i_29610(.A(n_57338), .Z(n_26317));
	notech_inv i_29611(.A(n_56296), .Z(n_26318));
	notech_inv i_29612(.A(n_56395), .Z(n_26319));
	notech_inv i_29613(.A(n_56285), .Z(n_26320));
	notech_inv i_29614(.A(n_59219), .Z(n_26321));
	notech_inv i_29617(.A(n_56255), .Z(n_26322));
	notech_inv i_29620(.A(n_145574323), .Z(n_26323));
	notech_inv i_29621(.A(n_142374291), .Z(n_26324));
	notech_inv i_29622(.A(n_147374341), .Z(n_26325));
	notech_inv i_29623(.A(n_56538), .Z(n_26326));
	notech_inv i_29624(.A(n_55302), .Z(n_26327));
	notech_inv i_29625(.A(n_186874736), .Z(n_26328));
	notech_inv i_29626(.A(n_188374751), .Z(n_26329));
	notech_inv i_29628(.A(n_177464112), .Z(n_26330));
	notech_inv i_29629(.A(n_177564113), .Z(n_26331));
	notech_inv i_29630(.A(n_189574763), .Z(n_26332));
	notech_inv i_29631(.A(n_190674774), .Z(n_26333));
	notech_inv i_29633(.A(n_191374781), .Z(n_26334));
	notech_inv i_29634(.A(n_192774795), .Z(n_26335));
	notech_inv i_29635(.A(n_193474802), .Z(n_26336));
	notech_inv i_29636(.A(n_194174809), .Z(n_26337));
	notech_inv i_29637(.A(n_196274830), .Z(n_26338));
	notech_inv i_29638(.A(n_168864026), .Z(n_26339));
	notech_inv i_29639(.A(n_201874886), .Z(n_26340));
	notech_inv i_29640(.A(n_208474952), .Z(n_26341));
	notech_inv i_29641(.A(n_321888472), .Z(n_26342));
	notech_inv i_29642(.A(n_221675077), .Z(n_26343));
	notech_inv i_29643(.A(n_237475227), .Z(n_26344));
	notech_inv i_29644(.A(n_238775240), .Z(n_26345));
	notech_inv i_29645(.A(n_240075253), .Z(n_26346));
	notech_inv i_29646(.A(n_267275511), .Z(n_26347));
	notech_inv i_29647(.A(n_268375522), .Z(n_26348));
	notech_inv i_29648(.A(n_269075529), .Z(n_26349));
	notech_inv i_29649(.A(n_269775536), .Z(n_26350));
	notech_inv i_29650(.A(n_270475543), .Z(n_26351));
	notech_inv i_29651(.A(n_271175550), .Z(n_26352));
	notech_inv i_29652(.A(n_271875557), .Z(n_26353));
	notech_inv i_29653(.A(n_272575564), .Z(n_26354));
	notech_inv i_29654(.A(n_273275571), .Z(n_26355));
	notech_inv i_29655(.A(n_273975578), .Z(n_26356));
	notech_inv i_29656(.A(n_274675585), .Z(n_26357));
	notech_inv i_29657(.A(n_304375882), .Z(n_26358));
	notech_inv i_29658(.A(n_305475893), .Z(n_26359));
	notech_inv i_29659(.A(n_306175900), .Z(n_26360));
	notech_inv i_29660(.A(n_134963687), .Z(n_26361));
	notech_inv i_29661(.A(n_307275911), .Z(n_26363));
	notech_inv i_29662(.A(n_308675925), .Z(n_26364));
	notech_inv i_29663(.A(n_309375932), .Z(n_26365));
	notech_inv i_29664(.A(n_310075939), .Z(n_26366));
	notech_inv i_29665(.A(n_133463672), .Z(n_26367));
	notech_inv i_29666(.A(n_310775946), .Z(n_26368));
	notech_inv i_29667(.A(n_132763665), .Z(n_26369));
	notech_inv i_29668(.A(n_312875967), .Z(n_26370));
	notech_inv i_29669(.A(n_313575974), .Z(n_26371));
	notech_inv i_29670(.A(n_314275981), .Z(n_26372));
	notech_inv i_29671(.A(n_314975988), .Z(n_26373));
	notech_inv i_29672(.A(n_57431), .Z(n_26374));
	notech_inv i_29673(.A(n_252861556), .Z(n_26375));
	notech_inv i_29674(.A(n_57441), .Z(n_26377));
	notech_inv i_29675(.A(n_323062234), .Z(n_26379));
	notech_inv i_29676(.A(n_57434), .Z(n_26380));
	notech_inv i_29677(.A(n_294261946), .Z(n_26381));
	notech_inv i_29678(.A(n_56420), .Z(n_26382));
	notech_inv i_29679(.A(n_151860600), .Z(n_26384));
	notech_inv i_29680(.A(n_56336), .Z(n_26385));
	notech_inv i_29681(.A(n_56511), .Z(n_26386));
	notech_inv i_29682(.A(n_56529), .Z(n_26387));
	notech_inv i_29684(.A(n_56327), .Z(n_26388));
	notech_inv i_29685(.A(n_341476251), .Z(n_26389));
	notech_inv i_29686(.A(n_59250), .Z(n_26390));
	notech_inv i_29687(.A(n_342176258), .Z(n_26391));
	notech_inv i_29688(.A(n_342976265), .Z(n_26393));
	notech_inv i_29689(.A(n_343676272), .Z(n_26394));
	notech_inv i_29690(.A(n_351288296), .Z(n_26395));
	notech_inv i_29691(.A(n_345776293), .Z(n_26396));
	notech_inv i_29692(.A(n_347176307), .Z(n_26397));
	notech_inv i_29693(.A(n_348676322), .Z(n_26398));
	notech_inv i_29694(.A(n_346488344), .Z(n_26399));
	notech_inv i_29695(.A(n_351976355), .Z(n_26400));
	notech_inv i_29696(.A(n_355276388), .Z(n_26401));
	notech_inv i_29697(.A(n_22579221), .Z(n_26403));
	notech_inv i_29698(.A(n_145974327), .Z(n_26404));
	notech_inv i_29699(.A(n_55729), .Z(n_26405));
	notech_inv i_29700(.A(n_57376), .Z(n_26406));
	notech_inv i_29701(.A(n_3314), .Z(n_26407));
	notech_inv i_29702(.A(n_188774755), .Z(n_26408));
	notech_inv i_29704(.A(n_189974767), .Z(n_26409));
	notech_inv i_29705(.A(n_322188469), .Z(n_26410));
	notech_inv i_29706(.A(n_323388457), .Z(n_26411));
	notech_inv i_29707(.A(n_264975488), .Z(n_26412));
	notech_inv i_29708(.A(n_265975498), .Z(n_26413));
	notech_inv i_29709(.A(n_267675515), .Z(n_26414));
	notech_inv i_29712(.A(n_323662240), .Z(n_26415));
	notech_inv i_29713(.A(n_304775886), .Z(n_26416));
	notech_inv i_29714(.A(n_306575904), .Z(n_26417));
	notech_inv i_29715(.A(n_57456), .Z(n_26418));
	notech_inv i_29716(.A(n_352376359), .Z(n_26419));
	notech_inv i_29717(.A(n_2224), .Z(n_26420));
	notech_inv i_29718(.A(n_149823485), .Z(n_26421));
	notech_inv i_29719(.A(n_54545), .Z(n_26422));
	notech_inv i_29720(.A(n_137177771), .Z(n_26423));
	notech_inv i_29721(.A(n_137677776), .Z(n_26424));
	notech_inv i_29722(.A(n_141477814), .Z(n_26425));
	notech_inv i_29723(.A(n_142177821), .Z(n_26426));
	notech_inv i_29724(.A(n_306062064), .Z(n_26427));
	notech_inv i_29725(.A(n_213278527), .Z(n_26428));
	notech_inv i_29726(.A(n_213578530), .Z(n_26429));
	notech_inv i_29727(.A(n_213778532), .Z(n_26430));
	notech_inv i_29728(.A(n_214578539), .Z(n_26431));
	notech_inv i_29729(.A(n_214878542), .Z(n_26432));
	notech_inv i_29730(.A(n_215078544), .Z(n_26433));
	notech_inv i_29731(.A(n_354069311), .Z(n_26434));
	notech_inv i_29732(.A(n_55819), .Z(n_26435));
	notech_inv i_29733(.A(n_237378763), .Z(n_26436));
	notech_inv i_29734(.A(n_271061738), .Z(n_26437));
	notech_inv i_29735(.A(n_239778787), .Z(n_26438));
	notech_inv i_29737(.A(n_241178801), .Z(n_26439));
	notech_inv i_29738(.A(n_241878808), .Z(n_26440));
	notech_inv i_29740(.A(n_247578865), .Z(n_26441));
	notech_inv i_29741(.A(n_260661634), .Z(n_26442));
	notech_inv i_29742(.A(n_301321900), .Z(n_26443));
	notech_inv i_29743(.A(n_2652), .Z(n_26444));
	notech_inv i_29744(.A(n_270588748), .Z(n_26445));
	notech_inv i_29745(.A(n_258678976), .Z(n_26446));
	notech_inv i_29746(.A(n_259278982), .Z(n_26447));
	notech_inv i_29747(.A(n_281779207), .Z(n_26448));
	notech_inv i_29748(.A(n_287979269), .Z(n_26449));
	notech_inv i_29749(.A(n_2701), .Z(n_26450));
	notech_inv i_29750(.A(n_322479614), .Z(n_26451));
	notech_inv i_29751(.A(n_323179621), .Z(n_26452));
	notech_inv i_29752(.A(n_323879628), .Z(n_26453));
	notech_inv i_29753(.A(n_324579635), .Z(n_26454));
	notech_inv i_29754(.A(n_331679706), .Z(n_26455));
	notech_inv i_29755(.A(n_332379713), .Z(n_26456));
	notech_inv i_29756(.A(n_333079720), .Z(n_26457));
	notech_inv i_29757(.A(n_333779727), .Z(n_26458));
	notech_inv i_29758(.A(n_188660960), .Z(n_26459));
	notech_inv i_29759(.A(n_190260976), .Z(n_26460));
	notech_inv i_29760(.A(n_189660970), .Z(n_26461));
	notech_inv i_29761(.A(n_344979797), .Z(n_26462));
	notech_inv i_29762(.A(n_152960611), .Z(n_26463));
	notech_inv i_29763(.A(n_220661279), .Z(n_26464));
	notech_inv i_29764(.A(n_155260634), .Z(n_26465));
	notech_inv i_29765(.A(n_219361266), .Z(n_26466));
	notech_inv i_29766(.A(n_154660628), .Z(n_26467));
	notech_inv i_29767(.A(n_55792), .Z(n_26468));
	notech_inv i_29768(.A(n_213361207), .Z(n_26469));
	notech_inv i_29769(.A(n_364079985), .Z(n_26470));
	notech_inv i_29770(.A(n_364379988), .Z(n_26471));
	notech_inv i_29771(.A(n_364579990), .Z(n_26472));
	notech_inv i_29772(.A(n_273388722), .Z(n_26473));
	notech_inv i_29773(.A(n_158660668), .Z(n_26474));
	notech_inv i_29774(.A(n_160060682), .Z(n_26475));
	notech_inv i_29775(.A(n_208061154), .Z(n_26476));
	notech_inv i_29776(.A(n_207661150), .Z(n_26477));
	notech_inv i_29777(.A(n_207361147), .Z(n_26478));
	notech_inv i_29778(.A(n_207061144), .Z(n_26480));
	notech_inv i_29779(.A(n_161460696), .Z(n_26481));
	notech_inv i_29780(.A(n_205261126), .Z(n_26483));
	notech_inv i_29781(.A(n_204561119), .Z(n_26484));
	notech_inv i_29782(.A(n_202061094), .Z(n_26485));
	notech_inv i_29783(.A(n_164860730), .Z(n_26486));
	notech_inv i_29784(.A(n_163760719), .Z(n_26487));
	notech_inv i_29785(.A(n_200561079), .Z(n_26488));
	notech_inv i_29786(.A(n_199761071), .Z(n_26489));
	notech_inv i_29787(.A(n_199461068), .Z(n_26490));
	notech_inv i_29788(.A(n_320179591), .Z(n_26491));
	notech_inv i_29789(.A(n_320579595), .Z(n_26492));
	notech_inv i_29790(.A(n_357479919), .Z(n_26493));
	notech_inv i_29791(.A(n_206841699), .Z(n_26494));
	notech_inv i_29792(.A(n_196861042), .Z(n_26495));
	notech_inv i_29793(.A(n_57442), .Z(n_26496));
	notech_inv i_29794(.A(n_275588702), .Z(n_26497));
	notech_inv i_29795(.A(n_2779), .Z(n_26498));
	notech_inv i_29796(.A(n_57432), .Z(n_26499));
	notech_inv i_29797(.A(n_55924), .Z(n_26500));
	notech_inv i_29798(.A(n_56033), .Z(n_26501));
	notech_inv i_29799(.A(n_57374), .Z(n_26502));
	notech_inv i_29800(.A(n_57378), .Z(n_26503));
	notech_inv i_29801(.A(n_54818), .Z(n_26504));
	notech_inv i_29802(.A(n_123981227), .Z(n_26505));
	notech_inv i_29803(.A(n_54874), .Z(n_26506));
	notech_inv i_29804(.A(n_166781655), .Z(n_26507));
	notech_inv i_29805(.A(n_54880), .Z(n_26508));
	notech_inv i_29806(.A(n_166981657), .Z(n_26509));
	notech_inv i_29807(.A(n_54770), .Z(n_26510));
	notech_inv i_29808(.A(n_55634), .Z(n_26511));
	notech_inv i_29809(.A(n_55893), .Z(n_26512));
	notech_inv i_29810(.A(n_55906), .Z(n_26513));
	notech_inv i_29811(.A(n_192861002), .Z(n_26514));
	notech_inv i_29812(.A(n_192560999), .Z(n_26515));
	notech_inv i_29813(.A(n_54507), .Z(n_26516));
	notech_inv i_29815(.A(n_172660808), .Z(n_26517));
	notech_inv i_29816(.A(n_189360967), .Z(n_26518));
	notech_inv i_29817(.A(n_164081628), .Z(n_26519));
	notech_inv i_29818(.A(n_172681714), .Z(n_26520));
	notech_inv i_29819(.A(n_187260946), .Z(n_26521));
	notech_inv i_29820(.A(n_174360825), .Z(n_26522));
	notech_inv i_29821(.A(n_185860932), .Z(n_26523));
	notech_inv i_29822(.A(n_185460928), .Z(n_26524));
	notech_inv i_29823(.A(n_184360917), .Z(n_26525));
	notech_inv i_29824(.A(n_183960913), .Z(n_26526));
	notech_inv i_29825(.A(n_175460836), .Z(n_26527));
	notech_inv i_29826(.A(n_180560886), .Z(n_26528));
	notech_inv i_29827(.A(n_180460885), .Z(n_26529));
	notech_inv i_29828(.A(n_179860879), .Z(n_26530));
	notech_inv i_29829(.A(n_178860870), .Z(n_26531));
	notech_inv i_29830(.A(n_178760869), .Z(n_26532));
	notech_inv i_29831(.A(n_178460866), .Z(n_26533));
	notech_inv i_29832(.A(n_178060862), .Z(n_26534));
	notech_inv i_29833(.A(n_177860860), .Z(n_26535));
	notech_inv i_29834(.A(n_2824), .Z(n_26536));
	notech_inv i_29838(.A(n_177060852), .Z(n_26538));
	notech_inv i_29839(.A(n_55752), .Z(n_26539));
	notech_inv i_29840(.A(n_135460436), .Z(n_26540));
	notech_inv i_29841(.A(n_141660498), .Z(n_26542));
	notech_inv i_29843(.A(n_54892), .Z(n_26543));
	notech_inv i_29845(.A(n_138860470), .Z(n_26544));
	notech_inv i_29846(.A(n_136660448), .Z(n_26545));
	notech_inv i_29848(.A(n_212282104), .Z(n_26546));
	notech_inv i_29849(.A(n_212382105), .Z(n_26547));
	notech_inv i_29852(.A(n_55268), .Z(n_26548));
	notech_inv i_29853(.A(n_323788453), .Z(n_26549));
	notech_inv i_29854(.A(n_56101), .Z(n_26550));
	notech_inv i_29856(.A(n_134860430), .Z(n_26551));
	notech_inv i_29857(.A(n_133760419), .Z(n_26552));
	notech_inv i_29858(.A(n_270488749), .Z(n_26553));
	notech_inv i_29859(.A(n_59163), .Z(n_26554));
	notech_inv i_29860(.A(n_56052), .Z(n_26555));
	notech_inv i_29863(.A(n_2190), .Z(n_26556));
	notech_inv i_29864(.A(n_216658447), .Z(n_26557));
	notech_inv i_29865(.A(n_323188459), .Z(n_26558));
	notech_inv i_29866(.A(n_322288468), .Z(n_26559));
	notech_inv i_29867(.A(n_208358369), .Z(n_26560));
	notech_inv i_29868(.A(n_320988480), .Z(n_26561));
	notech_inv i_29869(.A(n_183258118), .Z(n_26562));
	notech_inv i_29870(.A(n_182758113), .Z(n_26563));
	notech_inv i_29871(.A(n_318588504), .Z(n_26564));
	notech_inv i_29873(.A(n_352065809), .Z(n_26565));
	notech_inv i_29874(.A(n_270582680), .Z(n_26566));
	notech_inv i_29875(.A(n_271282687), .Z(n_26567));
	notech_inv i_29876(.A(n_271982694), .Z(n_26568));
	notech_inv i_29877(.A(n_272682701), .Z(n_26569));
	notech_inv i_29878(.A(n_55841), .Z(n_26570));
	notech_inv i_29879(.A(n_354869317), .Z(n_26571));
	notech_inv i_29880(.A(n_353065819), .Z(n_26572));
	notech_inv i_29881(.A(n_258958833), .Z(n_26573));
	notech_inv i_29882(.A(n_56144), .Z(n_26574));
	notech_inv i_29884(.A(n_311083085), .Z(n_26575));
	notech_inv i_29885(.A(n_56049), .Z(n_26576));
	notech_inv i_29886(.A(n_316783142), .Z(n_26577));
	notech_inv i_29887(.A(n_55102), .Z(n_26578));
	notech_inv i_29888(.A(n_55091), .Z(n_26579));
	notech_inv i_29889(.A(n_54822), .Z(n_26580));
	notech_inv i_29890(.A(n_56092), .Z(n_26581));
	notech_inv i_29891(.A(n_56126), .Z(n_26582));
	notech_inv i_29892(.A(n_55992), .Z(n_26583));
	notech_inv i_29893(.A(n_330483279), .Z(n_26584));
	notech_inv i_29894(.A(n_331183286), .Z(n_26585));
	notech_inv i_29895(.A(n_2269), .Z(n_26586));
	notech_inv i_29896(.A(n_56079), .Z(n_26587));
	notech_inv i_29897(.A(n_327546813), .Z(n_26588));
	notech_inv i_29898(.A(n_54968), .Z(n_26589));
	notech_inv i_29899(.A(n_494), .Z(n_26590));
	notech_inv i_29900(.A(n_56260), .Z(n_26591));
	notech_inv i_29901(.A(n_56551), .Z(n_26592));
	notech_inv i_29902(.A(n_54913), .Z(n_26593));
	notech_inv i_29903(.A(n_57438), .Z(n_26594));
	notech_inv i_29904(.A(n_27641995), .Z(n_26595));
	notech_inv i_29905(.A(n_54940), .Z(n_26596));
	notech_inv i_29906(.A(n_56409), .Z(n_26597));
	notech_inv i_29907(.A(n_54896), .Z(n_26598));
	notech_inv i_29908(.A(n_35829), .Z(n_26599));
	notech_inv i_29909(.A(n_56076), .Z(n_26600));
	notech_inv i_29910(.A(n_55657), .Z(n_26601));
	notech_inv i_29911(.A(n_210758392), .Z(n_26602));
	notech_inv i_29912(.A(n_204858334), .Z(n_26603));
	notech_inv i_29913(.A(n_275788700), .Z(n_26604));
	notech_inv i_29914(.A(n_56560), .Z(n_26605));
	notech_inv i_29915(.A(n_275888699), .Z(n_26606));
	notech_inv i_29916(.A(n_55324), .Z(n_26607));
	notech_inv i_29917(.A(n_55758), .Z(n_26608));
	notech_inv i_29918(.A(n_54967), .Z(n_26609));
	notech_inv i_29919(.A(n_264885968), .Z(n_26610));
	notech_inv i_29920(.A(n_57445), .Z(n_26611));
	notech_inv i_29921(.A(n_57444), .Z(n_26612));
	notech_inv i_29922(.A(n_55641), .Z(n_26613));
	notech_inv i_29923(.A(n_2823), .Z(n_26614));
	notech_inv i_29924(.A(n_275188706), .Z(n_26615));
	notech_inv i_29925(.A(n_273488721), .Z(n_26616));
	notech_inv i_29926(.A(n_280186121), .Z(n_26617));
	notech_inv i_29927(.A(n_310918886), .Z(n_26618));
	notech_inv i_29928(.A(n_58532), .Z(n_26619));
	notech_inv i_29929(.A(n_57372), .Z(n_26620));
	notech_inv i_29930(.A(n_60468), .Z(n_26621));
	notech_inv i_29931(.A(n_55625), .Z(n_26622));
	notech_inv i_29932(.A(n_93742656), .Z(n_26623));
	notech_inv i_29933(.A(n_55089), .Z(n_26624));
	notech_inv i_29934(.A(n_57446), .Z(n_26625));
	notech_inv i_29935(.A(n_189388132), .Z(n_26626));
	notech_inv i_29937(.A(\nbus_11334[0] ), .Z(n_26628));
	notech_inv i_29938(.A(n_59780), .Z(n_26629));
	notech_inv i_29939(.A(fecx), .Z(n_26630));
	notech_inv i_29940(.A(n_7487), .Z(n_26631));
	notech_inv i_29941(.A(sav_ecx[0]), .Z(n_26632));
	notech_inv i_29942(.A(sav_ecx[1]), .Z(n_26633));
	notech_inv i_29943(.A(sav_ecx[2]), .Z(n_26634));
	notech_inv i_29944(.A(sav_ecx[3]), .Z(n_26635));
	notech_inv i_29945(.A(sav_ecx[4]), .Z(n_26636));
	notech_inv i_29946(.A(sav_ecx[5]), .Z(n_26637));
	notech_inv i_29947(.A(sav_ecx[6]), .Z(n_26638));
	notech_inv i_29948(.A(sav_ecx[7]), .Z(n_26640));
	notech_inv i_29949(.A(sav_ecx[8]), .Z(n_26641));
	notech_inv i_29950(.A(sav_ecx[9]), .Z(n_26643));
	notech_inv i_29951(.A(sav_ecx[10]), .Z(n_26644));
	notech_inv i_29952(.A(sav_ecx[11]), .Z(n_26645));
	notech_inv i_29953(.A(sav_ecx[12]), .Z(n_26647));
	notech_inv i_29954(.A(sav_ecx[13]), .Z(n_26648));
	notech_inv i_29955(.A(sav_ecx[15]), .Z(n_26649));
	notech_inv i_29956(.A(n_2838), .Z(n_26650));
	notech_inv i_29957(.A(sav_ecx[18]), .Z(n_26651));
	notech_inv i_29958(.A(n_2837), .Z(n_26652));
	notech_inv i_29959(.A(sav_ecx[19]), .Z(n_26653));
	notech_inv i_29960(.A(sav_ecx[20]), .Z(n_26654));
	notech_inv i_29961(.A(sav_ecx[21]), .Z(n_26655));
	notech_inv i_29962(.A(sav_ecx[22]), .Z(n_26657));
	notech_inv i_29963(.A(sav_ecx[23]), .Z(n_26658));
	notech_inv i_29964(.A(sav_ecx[25]), .Z(n_26661));
	notech_inv i_29965(.A(n_231756227), .Z(n_26663));
	notech_inv i_29966(.A(sav_ecx[26]), .Z(n_26664));
	notech_inv i_29967(.A(n_2830), .Z(n_26666));
	notech_inv i_29968(.A(sav_ecx[27]), .Z(n_26673));
	notech_inv i_29969(.A(sav_ecx[28]), .Z(n_26674));
	notech_inv i_29970(.A(sav_ecx[29]), .Z(n_26676));
	notech_inv i_29971(.A(n_2826), .Z(n_26680));
	notech_inv i_29972(.A(sav_ecx[31]), .Z(n_26683));
	notech_inv i_29973(.A(fesp), .Z(n_26684));
	notech_inv i_29974(.A(sav_esp[0]), .Z(n_26685));
	notech_inv i_29975(.A(sav_esp[1]), .Z(n_26686));
	notech_inv i_29976(.A(sav_esp[2]), .Z(n_26687));
	notech_inv i_29979(.A(sav_esp[3]), .Z(n_26688));
	notech_inv i_29981(.A(sav_esp[4]), .Z(n_26689));
	notech_inv i_29982(.A(sav_esp[5]), .Z(n_26690));
	notech_inv i_29983(.A(sav_esp[6]), .Z(n_26691));
	notech_inv i_29985(.A(sav_esp[7]), .Z(n_26692));
	notech_inv i_29986(.A(sav_esp[8]), .Z(n_26693));
	notech_inv i_29987(.A(sav_esp[9]), .Z(n_26694));
	notech_inv i_29988(.A(sav_esp[10]), .Z(n_26695));
	notech_inv i_29989(.A(sav_esp[11]), .Z(n_26696));
	notech_inv i_29990(.A(sav_esp[12]), .Z(n_26697));
	notech_inv i_29991(.A(n_56972), .Z(n_26698));
	notech_inv i_29992(.A(sav_esp[13]), .Z(n_26699));
	notech_inv i_29993(.A(sav_esp[15]), .Z(n_26700));
	notech_inv i_29994(.A(sav_esp[16]), .Z(n_26701));
	notech_inv i_29995(.A(sav_esp[17]), .Z(n_26702));
	notech_inv i_29996(.A(sav_esp[18]), .Z(n_26703));
	notech_inv i_29997(.A(sav_esp[19]), .Z(n_26704));
	notech_inv i_29998(.A(sav_esp[20]), .Z(n_26705));
	notech_inv i_29999(.A(sav_esp[21]), .Z(n_26706));
	notech_inv i_30000(.A(sav_esp[22]), .Z(n_26707));
	notech_inv i_30001(.A(sav_esp[23]), .Z(n_26708));
	notech_inv i_30002(.A(sav_esp[24]), .Z(n_26709));
	notech_inv i_30003(.A(sav_esp[25]), .Z(n_26710));
	notech_inv i_30004(.A(sav_esp[26]), .Z(n_26711));
	notech_inv i_30005(.A(n_2792), .Z(n_26712));
	notech_inv i_30006(.A(sav_esp[27]), .Z(n_26713));
	notech_inv i_30007(.A(sav_esp[28]), .Z(n_26715));
	notech_inv i_30008(.A(sav_esi[0]), .Z(n_26716));
	notech_inv i_30009(.A(sav_esi[1]), .Z(n_26717));
	notech_inv i_30010(.A(sav_esi[2]), .Z(n_26718));
	notech_inv i_30011(.A(sav_esi[3]), .Z(n_26719));
	notech_inv i_30012(.A(sav_esi[4]), .Z(n_26720));
	notech_inv i_30013(.A(sav_esi[5]), .Z(n_26721));
	notech_inv i_30014(.A(sav_esi[6]), .Z(n_26722));
	notech_inv i_30015(.A(sav_esi[7]), .Z(n_26723));
	notech_inv i_30016(.A(sav_esi[9]), .Z(n_26724));
	notech_inv i_30017(.A(sav_esi[14]), .Z(n_26725));
	notech_inv i_30018(.A(sav_esi[17]), .Z(n_26726));
	notech_inv i_30019(.A(sav_esi[18]), .Z(n_26728));
	notech_inv i_30020(.A(sav_esi[19]), .Z(n_26729));
	notech_inv i_30021(.A(sav_esi[20]), .Z(n_26730));
	notech_inv i_30022(.A(sav_esi[21]), .Z(n_26731));
	notech_inv i_30024(.A(sav_esi[22]), .Z(n_26732));
	notech_inv i_30025(.A(sav_esi[23]), .Z(n_26733));
	notech_inv i_30026(.A(sav_esi[25]), .Z(n_26734));
	notech_inv i_30027(.A(sav_esi[26]), .Z(n_26735));
	notech_inv i_30028(.A(n_205888855), .Z(n_26736));
	notech_inv i_30029(.A(sav_esi[27]), .Z(n_26737));
	notech_inv i_30030(.A(sav_esi[28]), .Z(n_26738));
	notech_inv i_30031(.A(sav_esi[29]), .Z(n_26739));
	notech_inv i_30032(.A(sav_edi[1]), .Z(n_26740));
	notech_inv i_30033(.A(sav_edi[2]), .Z(n_26741));
	notech_inv i_30034(.A(sav_edi[3]), .Z(n_26742));
	notech_inv i_30035(.A(sav_edi[4]), .Z(n_26743));
	notech_inv i_30038(.A(sav_edi[5]), .Z(n_26744));
	notech_inv i_30039(.A(n_1915), .Z(n_26745));
	notech_inv i_30040(.A(sav_edi[6]), .Z(n_26746));
	notech_inv i_30041(.A(sav_edi[7]), .Z(n_26747));
	notech_inv i_30042(.A(sav_edi[8]), .Z(n_26748));
	notech_inv i_30043(.A(sav_edi[9]), .Z(n_26749));
	notech_inv i_30044(.A(sav_edi[10]), .Z(n_26750));
	notech_inv i_30045(.A(n_1919), .Z(n_26751));
	notech_inv i_30046(.A(sav_edi[11]), .Z(n_26752));
	notech_inv i_30048(.A(sav_edi[12]), .Z(n_26753));
	notech_inv i_30049(.A(sav_edi[13]), .Z(n_26754));
	notech_inv i_30050(.A(sav_edi[14]), .Z(n_26756));
	notech_inv i_30051(.A(sav_edi[15]), .Z(n_26757));
	notech_inv i_30052(.A(sav_edi[17]), .Z(n_26758));
	notech_inv i_30053(.A(sav_edi[18]), .Z(n_26759));
	notech_inv i_30054(.A(n_274688711), .Z(n_26760));
	notech_inv i_30055(.A(sav_edi[19]), .Z(n_26761));
	notech_inv i_30056(.A(sav_edi[20]), .Z(n_26762));
	notech_inv i_30058(.A(n_1911), .Z(n_26763));
	notech_inv i_30059(.A(sav_edi[21]), .Z(n_26764));
	notech_inv i_30060(.A(sav_edi[22]), .Z(n_26765));
	notech_inv i_30061(.A(sav_edi[23]), .Z(n_26766));
	notech_inv i_30062(.A(sav_edi[25]), .Z(n_26767));
	notech_inv i_30064(.A(sav_edi[26]), .Z(n_26769));
	notech_inv i_30065(.A(sav_edi[27]), .Z(n_26770));
	notech_inv i_30066(.A(sav_edi[28]), .Z(n_26771));
	notech_inv i_30067(.A(n_2739), .Z(n_26772));
	notech_inv i_30068(.A(n_206688847), .Z(n_26773));
	notech_inv i_30069(.A(sav_epc[8]), .Z(n_26774));
	notech_inv i_30070(.A(sav_epc[10]), .Z(n_26775));
	notech_inv i_30071(.A(n_190388902), .Z(n_26776));
	notech_inv i_30072(.A(sav_epc[11]), .Z(n_26777));
	notech_inv i_30073(.A(sav_epc[12]), .Z(n_26778));
	notech_inv i_30074(.A(sav_epc[13]), .Z(n_26779));
	notech_inv i_30075(.A(sav_epc[15]), .Z(n_26780));
	notech_inv i_30076(.A(sav_epc[16]), .Z(n_26781));
	notech_inv i_30077(.A(n_1900), .Z(n_26782));
	notech_inv i_30078(.A(sav_epc[18]), .Z(n_26783));
	notech_inv i_30079(.A(sav_epc[19]), .Z(n_26784));
	notech_inv i_30080(.A(n_2399), .Z(n_26785));
	notech_inv i_30082(.A(sav_epc[20]), .Z(n_26786));
	notech_inv i_30083(.A(sav_epc[21]), .Z(n_26787));
	notech_inv i_30084(.A(sav_epc[22]), .Z(n_26788));
	notech_inv i_30085(.A(sav_epc[23]), .Z(n_26789));
	notech_inv i_30086(.A(sav_epc[24]), .Z(n_26790));
	notech_inv i_30087(.A(sav_epc[25]), .Z(n_26791));
	notech_inv i_30088(.A(n_59958), .Z(n_26792));
	notech_inv i_30089(.A(sav_epc[26]), .Z(n_26793));
	notech_inv i_30090(.A(sav_epc[27]), .Z(n_26794));
	notech_inv i_30091(.A(n_106813462), .Z(n_26795));
	notech_inv i_30092(.A(sav_epc[30]), .Z(n_26796));
	notech_inv i_30093(.A(sav_epc[31]), .Z(n_26797));
	notech_inv i_30094(.A(\nbus_11284[0] ), .Z(n_26800));
	notech_inv i_30095(.A(n_7831), .Z(n_26801));
	notech_inv i_30096(.A(\nbus_11275[0] ), .Z(n_26803));
	notech_inv i_30097(.A(n_56386), .Z(n_26805));
	notech_inv i_30098(.A(n_271388742), .Z(n_26806));
	notech_inv i_30099(.A(n_2689), .Z(n_26807));
	notech_inv i_30100(.A(\nbus_11352[0] ), .Z(n_26808));
	notech_inv i_30102(.A(n_19785), .Z(n_26809));
	notech_inv i_30103(.A(n_19791), .Z(n_26810));
	notech_inv i_30104(.A(n_19797), .Z(n_26811));
	notech_inv i_30105(.A(n_19809), .Z(n_26812));
	notech_inv i_30106(.A(n_19821), .Z(n_26813));
	notech_inv i_30107(.A(n_19827), .Z(n_26814));
	notech_inv i_30109(.A(n_19845), .Z(n_26815));
	notech_inv i_30110(.A(n_19875), .Z(n_26816));
	notech_inv i_30111(.A(n_19917), .Z(n_26817));
	notech_inv i_30112(.A(n_19959), .Z(n_26818));
	notech_inv i_30113(.A(n_19965), .Z(n_26819));
	notech_inv i_30114(.A(n_19443), .Z(n_26820));
	notech_inv i_30115(.A(n_1025), .Z(n_26821));
	notech_inv i_30116(.A(n_19449), .Z(n_26822));
	notech_inv i_30117(.A(n_19461), .Z(n_26823));
	notech_inv i_30118(.A(n_19473), .Z(n_26824));
	notech_inv i_30119(.A(n_19479), .Z(n_26825));
	notech_inv i_30120(.A(n_1041), .Z(n_26826));
	notech_inv i_30121(.A(n_19485), .Z(n_26827));
	notech_inv i_30122(.A(n_19527), .Z(n_26828));
	notech_inv i_30123(.A(n_19569), .Z(n_26829));
	notech_inv i_30124(.A(n_19611), .Z(n_26830));
	notech_inv i_30125(.A(n_19617), .Z(n_26831));
	notech_inv i_30126(.A(n_19089), .Z(n_26832));
	notech_inv i_30127(.A(n_19095), .Z(n_26833));
	notech_inv i_30128(.A(n_19101), .Z(n_26834));
	notech_inv i_30129(.A(n_19113), .Z(n_26835));
	notech_inv i_30130(.A(n_19125), .Z(n_26836));
	notech_inv i_30131(.A(n_19131), .Z(n_26837));
	notech_inv i_30132(.A(n_19137), .Z(n_26838));
	notech_inv i_30133(.A(n_19149), .Z(n_26839));
	notech_inv i_30134(.A(n_19179), .Z(n_26840));
	notech_inv i_30135(.A(n_19221), .Z(n_26841));
	notech_inv i_30136(.A(n_19263), .Z(n_26842));
	notech_inv i_30137(.A(n_19269), .Z(n_26843));
	notech_inv i_30138(.A(\nbus_11349[0] ), .Z(n_26844));
	notech_inv i_30139(.A(n_8979), .Z(n_26845));
	notech_inv i_30140(.A(n_8985), .Z(n_26846));
	notech_inv i_30141(.A(n_8991), .Z(n_26847));
	notech_inv i_30142(.A(n_9003), .Z(n_26848));
	notech_inv i_30143(.A(n_9015), .Z(n_26849));
	notech_inv i_30144(.A(n_9021), .Z(n_26850));
	notech_inv i_30145(.A(n_9069), .Z(n_26851));
	notech_inv i_30146(.A(\nbus_11282[0] ), .Z(n_26852));
	notech_inv i_30147(.A(n_16699), .Z(n_26853));
	notech_inv i_30148(.A(n_16705), .Z(n_26854));
	notech_inv i_30149(.A(n_16711), .Z(n_26855));
	notech_inv i_30150(.A(n_2596), .Z(n_26856));
	notech_inv i_30151(.A(n_16717), .Z(n_26857));
	notech_inv i_30152(.A(n_16723), .Z(n_26858));
	notech_inv i_30153(.A(n_16735), .Z(n_26859));
	notech_inv i_30154(.A(n_16741), .Z(n_26860));
	notech_inv i_30155(.A(n_16747), .Z(n_26861));
	notech_inv i_30156(.A(n_2225), .Z(n_26862));
	notech_inv i_30157(.A(n_16753), .Z(n_26863));
	notech_inv i_30158(.A(n_16759), .Z(n_26864));
	notech_inv i_30159(.A(n_2573), .Z(n_26865));
	notech_inv i_30160(.A(n_16789), .Z(n_26866));
	notech_inv i_30161(.A(n_2586), .Z(n_26867));
	notech_inv i_30162(.A(n_16831), .Z(n_26868));
	notech_inv i_30163(.A(n_2385), .Z(n_26869));
	notech_inv i_30164(.A(n_16879), .Z(n_26870));
	notech_inv i_30165(.A(n_13815), .Z(n_26871));
	notech_inv i_30166(.A(n_13821), .Z(n_26872));
	notech_inv i_30167(.A(n_13827), .Z(n_26873));
	notech_inv i_30168(.A(n_13839), .Z(n_26874));
	notech_inv i_30169(.A(n_13851), .Z(n_26875));
	notech_inv i_30170(.A(n_13857), .Z(n_26876));
	notech_inv i_30171(.A(n_246156279), .Z(n_26877));
	notech_inv i_30172(.A(n_13905), .Z(n_26878));
	notech_inv i_30173(.A(n_13947), .Z(n_26879));
	notech_inv i_30174(.A(n_13989), .Z(n_26880));
	notech_inv i_30175(.A(\nbus_11311[0] ), .Z(n_26881));
	notech_inv i_30176(.A(n_13503), .Z(n_26882));
	notech_inv i_30177(.A(n_13509), .Z(n_26883));
	notech_inv i_30178(.A(n_13521), .Z(n_26884));
	notech_inv i_30179(.A(n_13527), .Z(n_26885));
	notech_inv i_30180(.A(pipe_mul[0]), .Z(n_26886));
	notech_inv i_30181(.A(eval_flag), .Z(n_26887));
	notech_inv i_30182(.A(rep_en1), .Z(n_26889));
	notech_inv i_30183(.A(rep_en4), .Z(n_26890));
	notech_inv i_30184(.A(nCF), .Z(n_26891));
	notech_inv i_30185(.A(nPF), .Z(n_26892));
	notech_inv i_30186(.A(n_8785), .Z(n_26893));
	notech_inv i_30187(.A(nSF), .Z(n_26894));
	notech_inv i_30188(.A(n_14933), .Z(n_26895));
	notech_inv i_30189(.A(n_20625), .Z(n_26896));
	notech_inv i_30190(.A(n_20649), .Z(n_26897));
	notech_inv i_30191(.A(\nbus_11353[10] ), .Z(n_26898));
	notech_inv i_30192(.A(n_20685), .Z(n_26899));
	notech_inv i_30193(.A(n_20751), .Z(n_26900));
	notech_inv i_30194(.A(n_20757), .Z(n_26901));
	notech_inv i_30195(.A(n_20763), .Z(n_26902));
	notech_inv i_30196(.A(n_20769), .Z(n_26903));
	notech_inv i_30197(.A(n_16368), .Z(n_26904));
	notech_inv i_30198(.A(n_16380), .Z(n_26905));
	notech_inv i_30199(.A(n_16386), .Z(n_26906));
	notech_inv i_30200(.A(n_16392), .Z(n_26907));
	notech_inv i_30201(.A(n_16404), .Z(n_26908));
	notech_inv i_30202(.A(n_16410), .Z(n_26909));
	notech_inv i_30203(.A(n_16434), .Z(n_26910));
	notech_inv i_30204(.A(n_16530), .Z(n_26911));
	notech_inv i_30205(.A(n_13115), .Z(n_26912));
	notech_inv i_30206(.A(n_13121), .Z(n_26913));
	notech_inv i_30208(.A(n_13127), .Z(n_26914));
	notech_inv i_30210(.A(n_13139), .Z(n_26915));
	notech_inv i_30211(.A(n_13151), .Z(n_26916));
	notech_inv i_30212(.A(n_13157), .Z(n_26917));
	notech_inv i_30213(.A(n_13205), .Z(n_26918));
	notech_inv i_30214(.A(n_13247), .Z(n_26919));
	notech_inv i_30215(.A(n_13295), .Z(n_26920));
	notech_inv i_30216(.A(n_14738), .Z(n_26921));
	notech_inv i_30217(.A(n_15018), .Z(n_26922));
	notech_inv i_30218(.A(temp_sp[0]), .Z(n_26923));
	notech_inv i_30219(.A(n_15023), .Z(n_26924));
	notech_inv i_30220(.A(temp_sp[1]), .Z(n_26925));
	notech_inv i_30221(.A(n_15028), .Z(n_26926));
	notech_inv i_30222(.A(temp_sp[2]), .Z(n_26927));
	notech_inv i_30223(.A(n_15033), .Z(n_26928));
	notech_inv i_30224(.A(temp_sp[3]), .Z(n_26929));
	notech_inv i_30225(.A(n_15038), .Z(n_26930));
	notech_inv i_30226(.A(temp_sp[4]), .Z(n_26931));
	notech_inv i_30227(.A(n_15043), .Z(n_26932));
	notech_inv i_30228(.A(temp_sp[5]), .Z(n_26933));
	notech_inv i_30229(.A(n_15048), .Z(n_26934));
	notech_inv i_30230(.A(temp_sp[6]), .Z(n_26935));
	notech_inv i_30231(.A(n_15053), .Z(n_26936));
	notech_inv i_30232(.A(temp_sp[7]), .Z(n_26937));
	notech_inv i_30233(.A(n_15058), .Z(n_26938));
	notech_inv i_30234(.A(temp_sp[8]), .Z(n_26939));
	notech_inv i_30235(.A(n_15063), .Z(n_26940));
	notech_inv i_30236(.A(temp_sp[9]), .Z(n_26941));
	notech_inv i_30237(.A(n_15068), .Z(n_26942));
	notech_inv i_30238(.A(temp_sp[10]), .Z(n_26943));
	notech_inv i_30239(.A(n_15073), .Z(n_26944));
	notech_inv i_30240(.A(temp_sp[11]), .Z(n_26945));
	notech_inv i_30241(.A(n_15078), .Z(n_26946));
	notech_inv i_30242(.A(temp_sp[12]), .Z(n_26947));
	notech_inv i_30243(.A(n_15083), .Z(n_26948));
	notech_inv i_30244(.A(temp_sp[13]), .Z(n_26949));
	notech_inv i_30245(.A(n_15088), .Z(n_26950));
	notech_inv i_30246(.A(temp_sp[14]), .Z(n_26951));
	notech_inv i_30247(.A(n_15093), .Z(n_26952));
	notech_inv i_30248(.A(temp_sp[15]), .Z(n_26953));
	notech_inv i_30249(.A(n_15098), .Z(n_26954));
	notech_inv i_30250(.A(temp_sp[16]), .Z(n_26955));
	notech_inv i_30251(.A(n_15103), .Z(n_26956));
	notech_inv i_30252(.A(temp_sp[17]), .Z(n_26957));
	notech_inv i_30253(.A(n_15108), .Z(n_26958));
	notech_inv i_30254(.A(temp_sp[18]), .Z(n_26959));
	notech_inv i_30255(.A(n_15113), .Z(n_26960));
	notech_inv i_30256(.A(temp_sp[19]), .Z(n_26961));
	notech_inv i_30257(.A(n_15118), .Z(n_26962));
	notech_inv i_30258(.A(temp_sp[20]), .Z(n_26963));
	notech_inv i_30259(.A(n_15123), .Z(n_26964));
	notech_inv i_30260(.A(temp_sp[21]), .Z(n_26965));
	notech_inv i_30261(.A(n_15128), .Z(n_26966));
	notech_inv i_30262(.A(temp_sp[22]), .Z(n_26967));
	notech_inv i_30263(.A(n_15133), .Z(n_26968));
	notech_inv i_30264(.A(temp_sp[23]), .Z(n_26969));
	notech_inv i_30265(.A(n_15138), .Z(n_26970));
	notech_inv i_30266(.A(temp_sp[24]), .Z(n_26971));
	notech_inv i_30267(.A(n_15143), .Z(n_26972));
	notech_inv i_30268(.A(temp_sp[25]), .Z(n_26973));
	notech_inv i_30269(.A(n_15148), .Z(n_26974));
	notech_inv i_30270(.A(temp_sp[26]), .Z(n_26975));
	notech_inv i_30271(.A(n_15153), .Z(n_26976));
	notech_inv i_30272(.A(temp_sp[27]), .Z(n_26977));
	notech_inv i_30273(.A(n_15158), .Z(n_26978));
	notech_inv i_30274(.A(temp_sp[28]), .Z(n_26979));
	notech_inv i_30275(.A(n_15163), .Z(n_26980));
	notech_inv i_30276(.A(temp_sp[29]), .Z(n_26983));
	notech_inv i_30277(.A(n_15168), .Z(n_26984));
	notech_inv i_30278(.A(temp_sp[30]), .Z(n_26985));
	notech_inv i_30279(.A(n_15173), .Z(n_26986));
	notech_inv i_30280(.A(temp_sp[31]), .Z(n_26987));
	notech_inv i_30281(.A(n_12773), .Z(n_26988));
	notech_inv i_30282(.A(n_12779), .Z(n_26989));
	notech_inv i_30284(.A(n_12785), .Z(n_26992));
	notech_inv i_30285(.A(n_12791), .Z(n_26993));
	notech_inv i_30286(.A(n_12797), .Z(n_26996));
	notech_inv i_30287(.A(n_12803), .Z(n_26997));
	notech_inv i_30288(.A(n_12809), .Z(n_26998));
	notech_inv i_30290(.A(\nbus_11308[0] ), .Z(n_27000));
	notech_inv i_30291(.A(n_12401), .Z(n_27002));
	notech_inv i_30292(.A(n_12407), .Z(n_27004));
	notech_inv i_30294(.A(n_12413), .Z(n_27005));
	notech_inv i_30295(.A(n_12425), .Z(n_27006));
	notech_inv i_30296(.A(n_12437), .Z(n_27007));
	notech_inv i_30297(.A(n_12443), .Z(n_27008));
	notech_inv i_30298(.A(n_12449), .Z(n_27009));
	notech_inv i_30299(.A(n_12461), .Z(n_27010));
	notech_inv i_30300(.A(n_12479), .Z(n_27011));
	notech_inv i_30301(.A(n_12491), .Z(n_27012));
	notech_inv i_30303(.A(n_12509), .Z(n_27013));
	notech_inv i_30304(.A(n_12515), .Z(n_27014));
	notech_inv i_30305(.A(n_12527), .Z(n_27015));
	notech_inv i_30306(.A(n_12533), .Z(n_27016));
	notech_inv i_30307(.A(n_12545), .Z(n_27017));
	notech_inv i_30308(.A(n_12557), .Z(n_27018));
	notech_inv i_30309(.A(n_2199), .Z(n_27019));
	notech_inv i_30310(.A(n_12569), .Z(n_27020));
	notech_inv i_30311(.A(n_12581), .Z(n_27021));
	notech_inv i_30312(.A(\nbus_11307[0] ), .Z(n_27022));
	notech_inv i_30313(.A(n_12055), .Z(n_27023));
	notech_inv i_30314(.A(n_12061), .Z(n_27024));
	notech_inv i_30315(.A(n_12073), .Z(n_27025));
	notech_inv i_30316(.A(n_12091), .Z(n_27026));
	notech_inv i_30317(.A(n_12097), .Z(n_27027));
	notech_inv i_30318(.A(n_12103), .Z(n_27028));
	notech_inv i_30319(.A(n_12109), .Z(n_27029));
	notech_inv i_30320(.A(n_12121), .Z(n_27030));
	notech_inv i_30321(.A(n_12163), .Z(n_27031));
	notech_inv i_30322(.A(n_12169), .Z(n_27032));
	notech_inv i_30323(.A(n_12187), .Z(n_27033));
	notech_inv i_30324(.A(n_12211), .Z(n_27034));
	notech_inv i_30325(.A(\nbus_11306[0] ), .Z(n_27035));
	notech_inv i_30326(.A(\nbus_14523[1] ), .Z(n_27036));
	notech_inv i_30327(.A(\nbus_14523[3] ), .Z(n_27037));
	notech_inv i_30328(.A(\nbus_14523[4] ), .Z(n_27038));
	notech_inv i_30329(.A(\nbus_14523[5] ), .Z(n_27039));
	notech_inv i_30330(.A(\nbus_14523[8] ), .Z(n_27040));
	notech_inv i_30331(.A(\nbus_14523[9] ), .Z(n_27041));
	notech_inv i_30332(.A(\nbus_14523[10] ), .Z(n_27042));
	notech_inv i_30333(.A(\nbus_14523[11] ), .Z(n_27043));
	notech_inv i_30334(.A(\nbus_14523[12] ), .Z(n_27044));
	notech_inv i_30335(.A(\nbus_14523[13] ), .Z(n_27045));
	notech_inv i_30336(.A(\nbus_14523[14] ), .Z(n_27046));
	notech_inv i_30337(.A(\nbus_14523[15] ), .Z(n_27047));
	notech_inv i_30338(.A(\nbus_14523[17] ), .Z(n_27048));
	notech_inv i_30339(.A(\nbus_14523[18] ), .Z(n_27049));
	notech_inv i_30340(.A(\nbus_14523[19] ), .Z(n_27050));
	notech_inv i_30341(.A(\nbus_14523[20] ), .Z(n_27051));
	notech_inv i_30342(.A(\nbus_14523[21] ), .Z(n_27052));
	notech_inv i_30343(.A(\nbus_14523[22] ), .Z(n_27053));
	notech_inv i_30344(.A(\nbus_14523[23] ), .Z(n_27054));
	notech_inv i_30345(.A(\nbus_14523[24] ), .Z(n_27055));
	notech_inv i_30346(.A(\nbus_14523[25] ), .Z(n_27056));
	notech_inv i_30347(.A(\nbus_14523[26] ), .Z(n_27057));
	notech_inv i_30348(.A(\nbus_14523[27] ), .Z(n_27058));
	notech_inv i_30349(.A(\nbus_14523[28] ), .Z(n_27059));
	notech_inv i_30350(.A(\nbus_14523[29] ), .Z(n_27060));
	notech_inv i_30351(.A(\nbus_14523[30] ), .Z(n_27061));
	notech_inv i_30352(.A(n_11415), .Z(n_27062));
	notech_inv i_30353(.A(n_11421), .Z(n_27063));
	notech_inv i_30354(.A(mask8b[1]), .Z(n_27064));
	notech_inv i_30355(.A(n_14092), .Z(n_27065));
	notech_inv i_30356(.A(n_14104), .Z(n_27066));
	notech_inv i_30357(.A(n_14110), .Z(n_27067));
	notech_inv i_30358(.A(n_14146), .Z(n_27068));
	notech_inv i_30359(.A(\nbus_11314[0] ), .Z(n_27069));
	notech_inv i_30360(.A(n_14188), .Z(n_27070));
	notech_inv i_30361(.A(n_14194), .Z(n_27071));
	notech_inv i_30362(.A(n_14272), .Z(n_27072));
	notech_inv i_30363(.A(n_14278), .Z(n_27073));
	notech_inv i_30364(.A(n_8477), .Z(n_27075));
	notech_inv i_30365(.A(n_8482), .Z(n_27077));
	notech_inv i_30366(.A(n_8487), .Z(n_27078));
	notech_inv i_30367(.A(n_8492), .Z(n_27079));
	notech_inv i_30368(.A(n_8497), .Z(n_27080));
	notech_inv i_30369(.A(n_206188852), .Z(n_27081));
	notech_inv i_30370(.A(n_8502), .Z(n_27082));
	notech_inv i_30371(.A(n_8507), .Z(n_27083));
	notech_inv i_30372(.A(n_8512), .Z(n_27084));
	notech_inv i_30373(.A(n_8517), .Z(n_27086));
	notech_inv i_30374(.A(n_8522), .Z(n_27087));
	notech_inv i_30375(.A(n_8527), .Z(n_27088));
	notech_inv i_30376(.A(n_8532), .Z(n_27089));
	notech_inv i_30377(.A(n_8537), .Z(n_27090));
	notech_inv i_30378(.A(n_8542), .Z(n_27091));
	notech_inv i_30379(.A(n_8547), .Z(n_27092));
	notech_inv i_30380(.A(n_8552), .Z(n_27094));
	notech_inv i_30381(.A(n_8557), .Z(n_27097));
	notech_inv i_30382(.A(n_8562), .Z(n_27098));
	notech_inv i_30383(.A(n_8567), .Z(n_27099));
	notech_inv i_30384(.A(n_8572), .Z(n_27100));
	notech_inv i_30385(.A(n_8577), .Z(n_27101));
	notech_inv i_30386(.A(n_8582), .Z(n_27102));
	notech_inv i_30387(.A(n_8587), .Z(n_27103));
	notech_inv i_30388(.A(n_8592), .Z(n_27104));
	notech_inv i_30389(.A(n_8597), .Z(n_27105));
	notech_inv i_30390(.A(n_8602), .Z(n_27106));
	notech_inv i_30391(.A(n_8607), .Z(n_27107));
	notech_inv i_30392(.A(n_8612), .Z(n_27108));
	notech_inv i_30393(.A(n_8617), .Z(n_27109));
	notech_inv i_30394(.A(n_8622), .Z(n_27110));
	notech_inv i_30397(.A(n_1944), .Z(n_27112));
	notech_inv i_30399(.A(n_21127), .Z(n_27114));
	notech_inv i_30400(.A(n_21152), .Z(n_27115));
	notech_inv i_30401(.A(n_21157), .Z(n_27116));
	notech_inv i_30402(.A(n_21162), .Z(n_27117));
	notech_inv i_30403(.A(n_21167), .Z(n_27118));
	notech_inv i_30404(.A(n_21172), .Z(n_27119));
	notech_inv i_30405(.A(n_21177), .Z(n_27120));
	notech_inv i_30406(.A(n_21182), .Z(n_27121));
	notech_inv i_30407(.A(n_21187), .Z(n_27122));
	notech_inv i_30408(.A(n_21192), .Z(n_27123));
	notech_inv i_30409(.A(n_21197), .Z(n_27124));
	notech_inv i_30410(.A(n_21277), .Z(n_27125));
	notech_inv i_30411(.A(n_11698), .Z(n_27126));
	notech_inv i_30412(.A(n_11704), .Z(n_27127));
	notech_inv i_30413(.A(n_11710), .Z(n_27128));
	notech_inv i_30414(.A(n_11716), .Z(n_27129));
	notech_inv i_30415(.A(n_11722), .Z(n_27130));
	notech_inv i_30416(.A(n_11728), .Z(n_27131));
	notech_inv i_30417(.A(n_11734), .Z(n_27132));
	notech_inv i_30418(.A(n_11746), .Z(n_27133));
	notech_inv i_30419(.A(n_11752), .Z(n_27134));
	notech_inv i_30420(.A(n_11806), .Z(n_27135));
	notech_inv i_30421(.A(n_11812), .Z(n_27136));
	notech_inv i_30422(.A(n_11830), .Z(n_27137));
	notech_inv i_30423(.A(n_11836), .Z(n_27138));
	notech_inv i_30424(.A(n_11842), .Z(n_27139));
	notech_inv i_30425(.A(n_11860), .Z(n_27140));
	notech_inv i_30426(.A(n_11872), .Z(n_27141));
	notech_inv i_30427(.A(\nbus_11286[0] ), .Z(n_27142));
	notech_inv i_30428(.A(\nbus_11286[5] ), .Z(n_27143));
	notech_inv i_30429(.A(\nbus_11286[8] ), .Z(n_27144));
	notech_inv i_30430(.A(\nbus_11286[16] ), .Z(n_27145));
	notech_inv i_30431(.A(nZF), .Z(n_27146));
	notech_inv i_30432(.A(n_15774), .Z(n_27147));
	notech_inv i_30433(.A(n_15798), .Z(n_27148));
	notech_inv i_30434(.A(n_15804), .Z(n_27149));
	notech_inv i_30435(.A(n_15810), .Z(n_27150));
	notech_inv i_30436(.A(n_15882), .Z(n_27151));
	notech_inv i_30437(.A(n_15888), .Z(n_27152));
	notech_inv i_30438(.A(n_15894), .Z(n_27153));
	notech_inv i_30439(.A(n_15900), .Z(n_27154));
	notech_inv i_30440(.A(n_15906), .Z(n_27155));
	notech_inv i_30441(.A(n_15912), .Z(n_27156));
	notech_inv i_30442(.A(n_15918), .Z(n_27157));
	notech_inv i_30443(.A(n_15924), .Z(n_27158));
	notech_inv i_30444(.A(n_15930), .Z(n_27159));
	notech_inv i_30445(.A(n_15936), .Z(n_27160));
	notech_inv i_30446(.A(n_15942), .Z(n_27161));
	notech_inv i_30447(.A(n_15948), .Z(n_27162));
	notech_inv i_30448(.A(\nbus_11330[0] ), .Z(n_27163));
	notech_inv i_30449(.A(nbus_14522[0]), .Z(n_27165));
	notech_inv i_30450(.A(nbus_14522[1]), .Z(n_27166));
	notech_inv i_30451(.A(nbus_14522[2]), .Z(n_27167));
	notech_inv i_30452(.A(nbus_14522[3]), .Z(n_27168));
	notech_inv i_30453(.A(nbus_14522[4]), .Z(n_27169));
	notech_inv i_30454(.A(nbus_14522[5]), .Z(n_27170));
	notech_inv i_30455(.A(nbus_14522[6]), .Z(n_27171));
	notech_inv i_30456(.A(nbus_14522[7]), .Z(n_27172));
	notech_inv i_30457(.A(nbus_14522[8]), .Z(n_27173));
	notech_inv i_30458(.A(nbus_14522[9]), .Z(n_27174));
	notech_inv i_30459(.A(nbus_14522[10]), .Z(n_27176));
	notech_inv i_30460(.A(nbus_14522[11]), .Z(n_27177));
	notech_inv i_30461(.A(nbus_14522[12]), .Z(n_27178));
	notech_inv i_30462(.A(nbus_14522[13]), .Z(n_27179));
	notech_inv i_30463(.A(nbus_14522[14]), .Z(n_27180));
	notech_inv i_30464(.A(nbus_14522[15]), .Z(n_27181));
	notech_inv i_30465(.A(nbus_14522[16]), .Z(n_27183));
	notech_inv i_30466(.A(nbus_14522[17]), .Z(n_27184));
	notech_inv i_30467(.A(nbus_14522[18]), .Z(n_27185));
	notech_inv i_30468(.A(nbus_14522[19]), .Z(n_27186));
	notech_inv i_30469(.A(nbus_14522[20]), .Z(n_27187));
	notech_inv i_30470(.A(nbus_14522[21]), .Z(n_27188));
	notech_inv i_30471(.A(nbus_14522[22]), .Z(n_27189));
	notech_inv i_30472(.A(nbus_14522[23]), .Z(n_27190));
	notech_inv i_30473(.A(nbus_14522[24]), .Z(n_27191));
	notech_inv i_30474(.A(nbus_14522[25]), .Z(n_27192));
	notech_inv i_30475(.A(nbus_14522[26]), .Z(n_27193));
	notech_inv i_30476(.A(nbus_14522[27]), .Z(n_27194));
	notech_inv i_30477(.A(nbus_14522[28]), .Z(n_27195));
	notech_inv i_30478(.A(nbus_14522[29]), .Z(n_27196));
	notech_inv i_30480(.A(nbus_14522[30]), .Z(n_27197));
	notech_inv i_30481(.A(nbus_14522[31]), .Z(n_27198));
	notech_inv i_30482(.A(cr2_reg[0]), .Z(n_27199));
	notech_inv i_30483(.A(cr2_reg[1]), .Z(n_27200));
	notech_inv i_30486(.A(cr2_reg[2]), .Z(n_27201));
	notech_inv i_30487(.A(cr2_reg[3]), .Z(n_27202));
	notech_inv i_30488(.A(cr2_reg[4]), .Z(n_27203));
	notech_inv i_30489(.A(cr2_reg[5]), .Z(n_27204));
	notech_inv i_30490(.A(cr2_reg[6]), .Z(n_27205));
	notech_inv i_30491(.A(cr2_reg[7]), .Z(n_27206));
	notech_inv i_30492(.A(cr2_reg[8]), .Z(n_27207));
	notech_inv i_30493(.A(cr2_reg[9]), .Z(n_27208));
	notech_inv i_30494(.A(cr2_reg[10]), .Z(n_27209));
	notech_inv i_30495(.A(cr2_reg[11]), .Z(n_27210));
	notech_inv i_30496(.A(cr2_reg[12]), .Z(n_27211));
	notech_inv i_30497(.A(cr2_reg[13]), .Z(n_27212));
	notech_inv i_30498(.A(cr2_reg[14]), .Z(n_27213));
	notech_inv i_30499(.A(cr2_reg[16]), .Z(n_27214));
	notech_inv i_30500(.A(cr2_reg[18]), .Z(n_27215));
	notech_inv i_30501(.A(cr2_reg[19]), .Z(n_27216));
	notech_inv i_30502(.A(cr2_reg[20]), .Z(n_27217));
	notech_inv i_30503(.A(cr2_reg[21]), .Z(n_27218));
	notech_inv i_30504(.A(cr2_reg[22]), .Z(n_27219));
	notech_inv i_30505(.A(cr2_reg[24]), .Z(n_27221));
	notech_inv i_30506(.A(cr2_reg[25]), .Z(n_27222));
	notech_inv i_30507(.A(cr2_reg[26]), .Z(n_27223));
	notech_inv i_30508(.A(cr2_reg[27]), .Z(n_27224));
	notech_inv i_30509(.A(cr2_reg[28]), .Z(n_27225));
	notech_inv i_30510(.A(cr2_reg[29]), .Z(n_27227));
	notech_inv i_30511(.A(cr2_reg[30]), .Z(n_27228));
	notech_inv i_30512(.A(cr2_reg[31]), .Z(n_27229));
	notech_inv i_30513(.A(\nbus_14521[0] ), .Z(n_27230));
	notech_inv i_30514(.A(\nbus_14521[1] ), .Z(n_27231));
	notech_inv i_30516(.A(\nbus_14521[2] ), .Z(n_27232));
	notech_inv i_30517(.A(\nbus_14521[3] ), .Z(n_27233));
	notech_inv i_30518(.A(\nbus_14521[4] ), .Z(n_27234));
	notech_inv i_30519(.A(\nbus_14521[5] ), .Z(n_27235));
	notech_inv i_30520(.A(\nbus_14521[6] ), .Z(n_27237));
	notech_inv i_30521(.A(\nbus_14521[7] ), .Z(n_27238));
	notech_inv i_30522(.A(n_17196), .Z(n_27239));
	notech_inv i_30523(.A(n_17202), .Z(n_27240));
	notech_inv i_30524(.A(n_17208), .Z(n_27241));
	notech_inv i_30525(.A(n_17214), .Z(n_27242));
	notech_inv i_30526(.A(n_17220), .Z(n_27243));
	notech_inv i_30527(.A(n_17226), .Z(n_27244));
	notech_inv i_30529(.A(n_17232), .Z(n_27245));
	notech_inv i_30530(.A(n_17238), .Z(n_27248));
	notech_inv i_30531(.A(\nbus_11339[0] ), .Z(n_27249));
	notech_inv i_30532(.A(n_17244), .Z(n_27250));
	notech_inv i_30533(.A(n_17250), .Z(n_27251));
	notech_inv i_30534(.A(n_17256), .Z(n_27252));
	notech_inv i_30535(.A(n_17262), .Z(n_27253));
	notech_inv i_30536(.A(n_17268), .Z(n_27254));
	notech_inv i_30537(.A(n_17280), .Z(n_27255));
	notech_inv i_30538(.A(n_17286), .Z(n_27256));
	notech_inv i_30539(.A(\nbus_11339[8] ), .Z(n_27257));
	notech_inv i_30540(.A(\nbus_11339[16] ), .Z(n_27258));
	notech_inv i_30541(.A(n_18841), .Z(n_27259));
	notech_inv i_30542(.A(n_18859), .Z(n_27261));
	notech_inv i_30543(.A(n_60739), .Z(n_27262));
	notech_inv i_30544(.A(n_14908), .Z(n_27263));
	notech_inv i_30545(.A(fsm[2]), .Z(n_27264));
	notech_inv i_30546(.A(n_60752), .Z(n_27265));
	notech_inv i_30547(.A(fsm[4]), .Z(n_27266));
	notech_inv i_30548(.A(vliw_pc[1]), .Z(n_27267));
	notech_inv i_30549(.A(vliw_pc[4]), .Z(n_27268));
	notech_inv i_30550(.A(Daddrgs[3]), .Z(n_27269));
	notech_inv i_30551(.A(Daddrgs[5]), .Z(n_27270));
	notech_inv i_30552(.A(Daddrgs[6]), .Z(n_27271));
	notech_inv i_30553(.A(Daddrgs[7]), .Z(n_27272));
	notech_inv i_30554(.A(Daddrgs[9]), .Z(n_27273));
	notech_inv i_30555(.A(Daddrgs[10]), .Z(n_27274));
	notech_inv i_30557(.A(Daddrgs[11]), .Z(n_27275));
	notech_inv i_30558(.A(Daddrgs[12]), .Z(n_27276));
	notech_inv i_30559(.A(Daddrgs[13]), .Z(n_27277));
	notech_inv i_30560(.A(Daddrgs[14]), .Z(n_27278));
	notech_inv i_30561(.A(Daddrgs[15]), .Z(n_27279));
	notech_inv i_30562(.A(Daddrgs[16]), .Z(n_27280));
	notech_inv i_30563(.A(Daddrgs[17]), .Z(n_27281));
	notech_inv i_30564(.A(Daddrgs[18]), .Z(n_27282));
	notech_inv i_30565(.A(Daddrgs[19]), .Z(n_27283));
	notech_inv i_30566(.A(Daddrgs[20]), .Z(n_27284));
	notech_inv i_30567(.A(Daddrgs[21]), .Z(n_27285));
	notech_inv i_30568(.A(Daddrgs[22]), .Z(n_27286));
	notech_inv i_30570(.A(Daddrgs[23]), .Z(n_27287));
	notech_inv i_30571(.A(Daddrgs[24]), .Z(n_27288));
	notech_inv i_30572(.A(Daddrgs[25]), .Z(n_27289));
	notech_inv i_30573(.A(Daddrgs[26]), .Z(n_27290));
	notech_inv i_30574(.A(Daddrgs[27]), .Z(n_27291));
	notech_inv i_30575(.A(Daddrgs[28]), .Z(n_27292));
	notech_inv i_30576(.A(Daddrgs[29]), .Z(n_27293));
	notech_inv i_30577(.A(Daddrgs[30]), .Z(n_27294));
	notech_inv i_30578(.A(Daddrgs[31]), .Z(n_27295));
	notech_inv i_30579(.A(n_18925), .Z(n_27296));
	notech_inv i_30580(.A(temp_ss[0]), .Z(n_27297));
	notech_inv i_30581(.A(temp_ss[1]), .Z(n_27298));
	notech_inv i_30582(.A(temp_ss[2]), .Z(n_27300));
	notech_inv i_30583(.A(temp_ss[3]), .Z(n_27301));
	notech_inv i_30584(.A(temp_ss[4]), .Z(n_27302));
	notech_inv i_30585(.A(temp_ss[5]), .Z(n_27304));
	notech_inv i_30586(.A(temp_ss[6]), .Z(n_27307));
	notech_inv i_30587(.A(temp_ss[7]), .Z(n_27308));
	notech_inv i_30588(.A(temp_ss[8]), .Z(n_27309));
	notech_inv i_30589(.A(temp_ss[9]), .Z(n_27310));
	notech_inv i_30590(.A(temp_ss[10]), .Z(n_27311));
	notech_inv i_30591(.A(temp_ss[11]), .Z(n_27312));
	notech_inv i_30592(.A(temp_ss[12]), .Z(n_27313));
	notech_inv i_30593(.A(temp_ss[13]), .Z(n_27314));
	notech_inv i_30594(.A(temp_ss[14]), .Z(n_27315));
	notech_inv i_30595(.A(temp_ss[15]), .Z(n_27316));
	notech_inv i_30596(.A(temp_ss[16]), .Z(n_27317));
	notech_inv i_30597(.A(temp_ss[17]), .Z(n_27318));
	notech_inv i_30598(.A(temp_ss[18]), .Z(n_27319));
	notech_inv i_30599(.A(temp_ss[19]), .Z(n_27320));
	notech_inv i_30600(.A(temp_ss[20]), .Z(n_27321));
	notech_inv i_30603(.A(temp_ss[21]), .Z(n_27322));
	notech_inv i_30607(.A(temp_ss[22]), .Z(n_27323));
	notech_inv i_30609(.A(temp_ss[23]), .Z(n_27324));
	notech_inv i_30610(.A(temp_ss[24]), .Z(n_27325));
	notech_inv i_30619(.A(temp_ss[25]), .Z(n_27326));
	notech_inv i_30620(.A(temp_ss[26]), .Z(n_27327));
	notech_inv i_30625(.A(temp_ss[27]), .Z(n_27328));
	notech_inv i_30626(.A(temp_ss[28]), .Z(n_27329));
	notech_inv i_30628(.A(temp_ss[29]), .Z(n_27330));
	notech_inv i_30629(.A(temp_ss[30]), .Z(n_27331));
	notech_inv i_30630(.A(temp_ss[31]), .Z(n_27332));
	notech_inv i_30631(.A(errco[0]), .Z(n_27333));
	notech_inv i_30632(.A(errco[1]), .Z(n_27334));
	notech_inv i_30633(.A(errco[2]), .Z(n_27335));
	notech_inv i_30634(.A(errco[3]), .Z(n_27336));
	notech_inv i_30635(.A(errco[4]), .Z(n_27337));
	notech_inv i_30636(.A(errco[5]), .Z(n_27338));
	notech_inv i_30638(.A(errco[6]), .Z(n_27339));
	notech_inv i_30639(.A(errco[7]), .Z(n_27340));
	notech_inv i_30640(.A(errco[8]), .Z(n_27341));
	notech_inv i_30642(.A(errco[9]), .Z(n_27342));
	notech_inv i_30643(.A(errco[10]), .Z(n_27343));
	notech_inv i_30645(.A(n_1266), .Z(n_27344));
	notech_inv i_30647(.A(errco[11]), .Z(n_27345));
	notech_inv i_30648(.A(errco[12]), .Z(n_27346));
	notech_inv i_30649(.A(errco[13]), .Z(n_27347));
	notech_inv i_30650(.A(errco[14]), .Z(n_27348));
	notech_inv i_30651(.A(errco[15]), .Z(n_27349));
	notech_inv i_30652(.A(errco[16]), .Z(n_27350));
	notech_inv i_30653(.A(errco[17]), .Z(n_27351));
	notech_inv i_30654(.A(errco[18]), .Z(n_27352));
	notech_inv i_30655(.A(errco[19]), .Z(n_27353));
	notech_inv i_30656(.A(errco[20]), .Z(n_27354));
	notech_inv i_30657(.A(errco[21]), .Z(n_27355));
	notech_inv i_30658(.A(errco[22]), .Z(n_27356));
	notech_inv i_30659(.A(errco[23]), .Z(n_27357));
	notech_inv i_30660(.A(errco[24]), .Z(n_27358));
	notech_inv i_30661(.A(errco[25]), .Z(n_27359));
	notech_inv i_30662(.A(errco[26]), .Z(n_27360));
	notech_inv i_30663(.A(errco[27]), .Z(n_27361));
	notech_inv i_30664(.A(errco[28]), .Z(n_27362));
	notech_inv i_30665(.A(errco[29]), .Z(n_27363));
	notech_inv i_30666(.A(errco[30]), .Z(n_27364));
	notech_inv i_30667(.A(errco[31]), .Z(n_27365));
	notech_inv i_30668(.A(\nbus_11345[0] ), .Z(n_27366));
	notech_inv i_30669(.A(n_17661), .Z(n_27367));
	notech_inv i_30670(.A(n_10127), .Z(n_27368));
	notech_inv i_30671(.A(\nbus_14523[31] ), .Z(n_27369));
	notech_inv i_30672(.A(ecx[0]), .Z(n_27370));
	notech_inv i_30673(.A(ecx[1]), .Z(n_27371));
	notech_inv i_30674(.A(ecx[2]), .Z(n_27372));
	notech_inv i_30675(.A(ecx[3]), .Z(n_27373));
	notech_inv i_30676(.A(ecx[4]), .Z(n_27374));
	notech_inv i_30677(.A(ecx[5]), .Z(n_27375));
	notech_inv i_30678(.A(ecx[6]), .Z(n_27376));
	notech_inv i_30679(.A(ecx[7]), .Z(n_27377));
	notech_inv i_30680(.A(ecx[8]), .Z(n_27378));
	notech_inv i_30681(.A(ecx[9]), .Z(n_27379));
	notech_inv i_30682(.A(ecx[10]), .Z(n_27380));
	notech_inv i_30683(.A(ecx[11]), .Z(n_27381));
	notech_inv i_30684(.A(ecx[12]), .Z(n_27382));
	notech_inv i_30685(.A(ecx[13]), .Z(n_27383));
	notech_inv i_30686(.A(ecx[14]), .Z(n_27384));
	notech_inv i_30687(.A(ecx[15]), .Z(n_27385));
	notech_inv i_30688(.A(ecx[16]), .Z(n_27386));
	notech_inv i_30689(.A(ecx[17]), .Z(n_27387));
	notech_inv i_30690(.A(ecx[18]), .Z(n_27388));
	notech_inv i_30691(.A(ecx[19]), .Z(n_27389));
	notech_inv i_30692(.A(ecx[20]), .Z(n_27390));
	notech_inv i_30693(.A(ecx[21]), .Z(n_27391));
	notech_inv i_30694(.A(ecx[22]), .Z(n_27392));
	notech_inv i_30695(.A(ecx[23]), .Z(n_27393));
	notech_inv i_30696(.A(ecx[24]), .Z(n_27394));
	notech_inv i_30697(.A(ecx[25]), .Z(n_27395));
	notech_inv i_30698(.A(ecx[26]), .Z(n_27396));
	notech_inv i_30699(.A(ecx[27]), .Z(n_27397));
	notech_inv i_30700(.A(ecx[28]), .Z(n_27398));
	notech_inv i_30701(.A(ecx[29]), .Z(n_27399));
	notech_inv i_30702(.A(ecx[30]), .Z(n_27400));
	notech_inv i_30703(.A(ecx[31]), .Z(n_27401));
	notech_inv i_30704(.A(calc_sz[0]), .Z(n_27402));
	notech_inv i_30705(.A(calc_sz[1]), .Z(n_27403));
	notech_inv i_30706(.A(calc_sz[3]), .Z(n_27404));
	notech_inv i_30707(.A(opa[0]), .Z(nbus_11273[0]));
	notech_inv i_30708(.A(n_59708), .Z(nbus_11273[1]));
	notech_inv i_30709(.A(n_59717), .Z(nbus_11273[2]));
	notech_inv i_30710(.A(opa[3]), .Z(nbus_11273[3]));
	notech_inv i_30711(.A(n_59726), .Z(nbus_11273[4]));
	notech_inv i_30712(.A(opa[5]), .Z(nbus_11273[5]));
	notech_inv i_30713(.A(n_59735), .Z(nbus_11273[6]));
	notech_inv i_30714(.A(n_59744), .Z(nbus_11273[7]));
	notech_inv i_30715(.A(opa[8]), .Z(nbus_11273[8]));
	notech_inv i_30716(.A(opa[9]), .Z(nbus_11273[9]));
	notech_inv i_30717(.A(opa[10]), .Z(nbus_11273[10]));
	notech_inv i_30718(.A(opa[11]), .Z(nbus_11273[11]));
	notech_inv i_30719(.A(opa[12]), .Z(nbus_11273[12]));
	notech_inv i_30720(.A(opa[13]), .Z(nbus_11273[13]));
	notech_inv i_30721(.A(opa[14]), .Z(nbus_11273[14]));
	notech_inv i_30722(.A(opa[15]), .Z(nbus_11273[15]));
	notech_inv i_30723(.A(opa[16]), .Z(nbus_11273[16]));
	notech_inv i_30724(.A(opa[17]), .Z(nbus_11273[17]));
	notech_inv i_30725(.A(opa[18]), .Z(nbus_11273[18]));
	notech_inv i_30726(.A(opa[19]), .Z(nbus_11273[19]));
	notech_inv i_30727(.A(opa[20]), .Z(nbus_11273[20]));
	notech_inv i_30728(.A(opa[21]), .Z(nbus_11273[21]));
	notech_inv i_30729(.A(opa[22]), .Z(nbus_11273[22]));
	notech_inv i_30730(.A(opa[23]), .Z(nbus_11273[23]));
	notech_inv i_30731(.A(opa[24]), .Z(nbus_11273[24]));
	notech_inv i_30732(.A(opa[25]), .Z(nbus_11273[25]));
	notech_inv i_30733(.A(opa[26]), .Z(nbus_11273[26]));
	notech_inv i_30734(.A(opa[27]), .Z(nbus_11273[27]));
	notech_inv i_30735(.A(opa[28]), .Z(nbus_11273[28]));
	notech_inv i_30736(.A(opa[29]), .Z(nbus_11273[29]));
	notech_inv i_30737(.A(opa[30]), .Z(nbus_11273[30]));
	notech_inv i_30738(.A(opa[31]), .Z(nbus_11273[31]));
	notech_inv i_30739(.A(opb[0]), .Z(\nbus_11276[0] ));
	notech_inv i_30740(.A(opb[1]), .Z(\nbus_11276[1] ));
	notech_inv i_30741(.A(opb[2]), .Z(\nbus_11276[2] ));
	notech_inv i_30742(.A(opb[3]), .Z(\nbus_11276[3] ));
	notech_inv i_30743(.A(opb[4]), .Z(\nbus_11276[4] ));
	notech_inv i_30744(.A(opb[5]), .Z(\nbus_11276[5] ));
	notech_inv i_30746(.A(opb[6]), .Z(\nbus_11276[6] ));
	notech_inv i_30747(.A(opb[7]), .Z(\nbus_11276[7] ));
	notech_inv i_30748(.A(opb[8]), .Z(\nbus_11276[8] ));
	notech_inv i_30749(.A(opb[9]), .Z(\nbus_11276[9] ));
	notech_inv i_30750(.A(opb[10]), .Z(\nbus_11276[10] ));
	notech_inv i_30751(.A(opb[11]), .Z(\nbus_11276[11] ));
	notech_inv i_30752(.A(opb[12]), .Z(\nbus_11276[12] ));
	notech_inv i_30753(.A(opb[13]), .Z(\nbus_11276[13] ));
	notech_inv i_30754(.A(opb[14]), .Z(\nbus_11276[14] ));
	notech_inv i_30755(.A(opb[15]), .Z(\nbus_11276[15] ));
	notech_inv i_30756(.A(opb[16]), .Z(\nbus_11276[16] ));
	notech_inv i_30757(.A(opb[17]), .Z(\nbus_11276[17] ));
	notech_inv i_30758(.A(opb[18]), .Z(\nbus_11276[18] ));
	notech_inv i_30759(.A(opb[19]), .Z(\nbus_11276[19] ));
	notech_inv i_30760(.A(opb[20]), .Z(\nbus_11276[20] ));
	notech_inv i_30761(.A(opb[21]), .Z(\nbus_11276[21] ));
	notech_inv i_30762(.A(opb[22]), .Z(\nbus_11276[22] ));
	notech_inv i_30763(.A(opb[23]), .Z(\nbus_11276[23] ));
	notech_inv i_30764(.A(opb[24]), .Z(\nbus_11276[24] ));
	notech_inv i_30765(.A(opb[25]), .Z(\nbus_11276[25] ));
	notech_inv i_30766(.A(opb[26]), .Z(\nbus_11276[26] ));
	notech_inv i_30767(.A(opb[27]), .Z(\nbus_11276[27] ));
	notech_inv i_30768(.A(opb[28]), .Z(\nbus_11276[28] ));
	notech_inv i_30769(.A(opb[29]), .Z(\nbus_11276[29] ));
	notech_inv i_30770(.A(opb[30]), .Z(\nbus_11276[30] ));
	notech_inv i_30771(.A(opb[31]), .Z(\nbus_11276[31] ));
	notech_inv i_30772(.A(n_59113), .Z(nbus_11326[0]));
	notech_inv i_30773(.A(opc[1]), .Z(nbus_11326[1]));
	notech_inv i_30774(.A(opc[2]), .Z(nbus_11326[2]));
	notech_inv i_30775(.A(opc[3]), .Z(nbus_11326[3]));
	notech_inv i_30776(.A(opc[4]), .Z(nbus_11326[4]));
	notech_inv i_30777(.A(opc[5]), .Z(nbus_11326[5]));
	notech_inv i_30778(.A(opc[6]), .Z(nbus_11326[6]));
	notech_inv i_30779(.A(opc[7]), .Z(nbus_11326[7]));
	notech_inv i_30780(.A(opc[8]), .Z(nbus_11326[8]));
	notech_inv i_30781(.A(opc[9]), .Z(nbus_11326[9]));
	notech_inv i_30782(.A(opc[10]), .Z(nbus_11326[10]));
	notech_inv i_30783(.A(opc[11]), .Z(nbus_11326[11]));
	notech_inv i_30784(.A(opc[12]), .Z(nbus_11326[12]));
	notech_inv i_30785(.A(opc[13]), .Z(nbus_11326[13]));
	notech_inv i_30786(.A(opc[14]), .Z(nbus_11326[14]));
	notech_inv i_30787(.A(opc[15]), .Z(nbus_11326[15]));
	notech_inv i_30788(.A(opc[16]), .Z(nbus_11326[16]));
	notech_inv i_30789(.A(opc[17]), .Z(nbus_11326[17]));
	notech_inv i_30790(.A(opc[18]), .Z(nbus_11326[18]));
	notech_inv i_30791(.A(opc[19]), .Z(nbus_11326[19]));
	notech_inv i_30792(.A(opc[20]), .Z(nbus_11326[20]));
	notech_inv i_30793(.A(opc[21]), .Z(nbus_11326[21]));
	notech_inv i_30794(.A(opc[22]), .Z(nbus_11326[22]));
	notech_inv i_30795(.A(opc[23]), .Z(nbus_11326[23]));
	notech_inv i_30796(.A(opc[24]), .Z(nbus_11326[24]));
	notech_inv i_30797(.A(opc[25]), .Z(nbus_11326[25]));
	notech_inv i_30798(.A(opc[26]), .Z(nbus_11326[26]));
	notech_inv i_30799(.A(opc[27]), .Z(nbus_11326[27]));
	notech_inv i_30800(.A(opc[28]), .Z(nbus_11326[28]));
	notech_inv i_30802(.A(opc[29]), .Z(nbus_11326[29]));
	notech_inv i_30803(.A(opc[30]), .Z(nbus_11326[30]));
	notech_inv i_30805(.A(opc[31]), .Z(nbus_11326[31]));
	notech_inv i_30806(.A(opz[0]), .Z(n_27517));
	notech_inv i_30807(.A(opz[1]), .Z(n_27518));
	notech_inv i_30808(.A(read_data[0]), .Z(n_27519));
	notech_inv i_30809(.A(read_data[1]), .Z(n_27520));
	notech_inv i_30810(.A(read_data[2]), .Z(n_27521));
	notech_inv i_30811(.A(read_data[3]), .Z(n_27522));
	notech_inv i_30812(.A(read_data[4]), .Z(n_27523));
	notech_inv i_30813(.A(read_data[5]), .Z(n_27524));
	notech_inv i_30814(.A(read_data[6]), .Z(n_27525));
	notech_inv i_30815(.A(read_data[7]), .Z(n_27526));
	notech_inv i_30816(.A(read_data[8]), .Z(n_27527));
	notech_inv i_30817(.A(read_data[9]), .Z(n_27528));
	notech_inv i_30818(.A(read_data[10]), .Z(n_27529));
	notech_inv i_30819(.A(read_data[11]), .Z(n_27530));
	notech_inv i_30820(.A(read_data[12]), .Z(n_27531));
	notech_inv i_30821(.A(read_data[13]), .Z(n_27532));
	notech_inv i_30822(.A(read_data[14]), .Z(n_27533));
	notech_inv i_30823(.A(read_data[15]), .Z(n_27534));
	notech_inv i_30824(.A(read_data[16]), .Z(n_27535));
	notech_inv i_30825(.A(read_data[17]), .Z(n_27537));
	notech_inv i_30826(.A(read_data[18]), .Z(n_27538));
	notech_inv i_30827(.A(read_data[19]), .Z(n_27539));
	notech_inv i_30828(.A(read_data[20]), .Z(n_27540));
	notech_inv i_30829(.A(read_data[21]), .Z(n_27541));
	notech_inv i_30830(.A(read_data[22]), .Z(n_27542));
	notech_inv i_30831(.A(read_data[23]), .Z(n_27545));
	notech_inv i_30832(.A(read_data[24]), .Z(n_27546));
	notech_inv i_30833(.A(read_data[25]), .Z(n_27548));
	notech_inv i_30834(.A(read_data[26]), .Z(n_27549));
	notech_inv i_30835(.A(read_data[27]), .Z(n_27550));
	notech_inv i_30836(.A(read_data[28]), .Z(n_27551));
	notech_inv i_30837(.A(read_data[29]), .Z(n_27552));
	notech_inv i_30838(.A(read_data[30]), .Z(n_27553));
	notech_inv i_30839(.A(read_data[31]), .Z(n_27554));
	notech_inv i_30840(.A(all_cnt[0]), .Z(n_27555));
	notech_inv i_30841(.A(all_cnt[1]), .Z(n_27556));
	notech_inv i_30842(.A(all_cnt[2]), .Z(n_27557));
	notech_inv i_30843(.A(all_cnt[3]), .Z(n_27558));
	notech_inv i_30844(.A(cs[0]), .Z(n_27559));
	notech_inv i_30845(.A(cs[1]), .Z(n_27560));
	notech_inv i_30846(.A(opd[0]), .Z(n_27561));
	notech_inv i_30847(.A(opd[1]), .Z(n_27562));
	notech_inv i_30848(.A(opd[2]), .Z(n_27563));
	notech_inv i_30849(.A(opd[3]), .Z(n_27564));
	notech_inv i_30850(.A(opd[4]), .Z(n_27565));
	notech_inv i_30851(.A(opd[5]), .Z(n_27566));
	notech_inv i_30852(.A(opd[6]), .Z(n_27568));
	notech_inv i_30853(.A(opd[7]), .Z(n_27570));
	notech_inv i_30854(.A(opd[8]), .Z(n_27571));
	notech_inv i_30855(.A(opd[9]), .Z(n_27574));
	notech_inv i_30856(.A(opd[10]), .Z(n_27575));
	notech_inv i_30857(.A(opd[11]), .Z(n_27576));
	notech_inv i_30858(.A(opd[12]), .Z(n_27577));
	notech_inv i_30859(.A(opd[13]), .Z(n_27578));
	notech_inv i_30860(.A(opd[14]), .Z(n_27579));
	notech_inv i_30861(.A(opd[15]), .Z(n_27581));
	notech_inv i_30862(.A(opd[16]), .Z(n_27582));
	notech_inv i_30863(.A(opd[17]), .Z(n_27583));
	notech_inv i_30864(.A(opd[18]), .Z(n_27584));
	notech_inv i_30865(.A(opd[19]), .Z(n_27585));
	notech_inv i_30866(.A(opd[20]), .Z(n_27586));
	notech_inv i_30867(.A(opd[21]), .Z(n_27588));
	notech_inv i_30868(.A(opd[22]), .Z(n_27589));
	notech_inv i_30869(.A(opd[23]), .Z(n_27590));
	notech_inv i_30870(.A(opd[24]), .Z(n_27592));
	notech_inv i_30871(.A(opd[25]), .Z(n_27593));
	notech_inv i_30872(.A(opd[26]), .Z(n_27594));
	notech_inv i_30873(.A(opd[27]), .Z(n_27595));
	notech_inv i_30874(.A(opd[28]), .Z(n_27596));
	notech_inv i_30875(.A(opd[29]), .Z(n_27597));
	notech_inv i_30876(.A(opd[30]), .Z(n_27599));
	notech_inv i_30877(.A(opd[31]), .Z(n_27601));
	notech_inv i_30878(.A(regs_12[0]), .Z(n_27602));
	notech_inv i_30879(.A(regs_12[1]), .Z(n_27605));
	notech_inv i_30880(.A(regs_12[2]), .Z(n_27608));
	notech_inv i_30882(.A(regs_12[3]), .Z(n_27609));
	notech_inv i_30883(.A(regs_12[4]), .Z(n_27610));
	notech_inv i_30884(.A(regs_12[5]), .Z(n_27611));
	notech_inv i_30885(.A(regs_12[6]), .Z(n_27612));
	notech_inv i_30886(.A(regs_12[7]), .Z(n_27613));
	notech_inv i_30887(.A(regs_12[8]), .Z(n_27614));
	notech_inv i_30888(.A(regs_12[9]), .Z(n_27615));
	notech_inv i_30889(.A(regs_12[10]), .Z(n_27616));
	notech_inv i_30890(.A(regs_12[11]), .Z(n_27617));
	notech_inv i_30891(.A(regs_12[12]), .Z(n_27618));
	notech_inv i_30892(.A(regs_12[13]), .Z(n_27619));
	notech_inv i_30893(.A(regs_12[14]), .Z(n_27620));
	notech_inv i_30895(.A(regs_12[15]), .Z(n_27621));
	notech_inv i_30896(.A(regs_12[16]), .Z(n_27622));
	notech_inv i_30897(.A(regs_12[17]), .Z(n_27623));
	notech_inv i_30898(.A(regs_12[18]), .Z(n_27624));
	notech_inv i_30899(.A(regs_12[19]), .Z(n_27625));
	notech_inv i_30901(.A(regs_12[20]), .Z(n_27626));
	notech_inv i_30902(.A(regs_12[21]), .Z(n_27627));
	notech_inv i_30903(.A(regs_12[22]), .Z(n_27628));
	notech_inv i_30904(.A(regs_12[23]), .Z(n_27629));
	notech_inv i_30905(.A(regs_12[24]), .Z(n_27630));
	notech_inv i_30906(.A(regs_12[25]), .Z(n_27631));
	notech_inv i_30908(.A(regs_12[26]), .Z(n_27632));
	notech_inv i_30909(.A(regs_12[27]), .Z(n_27633));
	notech_inv i_30910(.A(regs_12[28]), .Z(n_27634));
	notech_inv i_30911(.A(regs_12[29]), .Z(n_27635));
	notech_inv i_30912(.A(regs_12[30]), .Z(n_27636));
	notech_inv i_30913(.A(regs_12[31]), .Z(n_27638));
	notech_inv i_30914(.A(regs_8[0]), .Z(n_27639));
	notech_inv i_30915(.A(regs_8[1]), .Z(n_27640));
	notech_inv i_30916(.A(regs_8[2]), .Z(n_27641));
	notech_inv i_30917(.A(regs_8[3]), .Z(n_27642));
	notech_inv i_30918(.A(regs_8[4]), .Z(n_27643));
	notech_inv i_30919(.A(regs_8[5]), .Z(n_27644));
	notech_inv i_30922(.A(regs_8[6]), .Z(n_27646));
	notech_inv i_30923(.A(regs_8[7]), .Z(n_27647));
	notech_inv i_30924(.A(regs_8[8]), .Z(n_27649));
	notech_inv i_30925(.A(regs_8[9]), .Z(n_27650));
	notech_inv i_30926(.A(regs_8[10]), .Z(n_27652));
	notech_inv i_30927(.A(regs_8[11]), .Z(n_27653));
	notech_inv i_30928(.A(regs_8[12]), .Z(n_27654));
	notech_inv i_30929(.A(regs_8[13]), .Z(n_27655));
	notech_inv i_30930(.A(regs_8[14]), .Z(n_27657));
	notech_inv i_30931(.A(regs_8[15]), .Z(n_27658));
	notech_inv i_30932(.A(regs_8[16]), .Z(n_27659));
	notech_inv i_30933(.A(regs_8[17]), .Z(n_27660));
	notech_inv i_30934(.A(regs_8[18]), .Z(n_27661));
	notech_inv i_30935(.A(regs_8[19]), .Z(n_27662));
	notech_inv i_30936(.A(regs_8[20]), .Z(n_27666));
	notech_inv i_30937(.A(regs_8[21]), .Z(n_27667));
	notech_inv i_30938(.A(regs_8[22]), .Z(n_27669));
	notech_inv i_30939(.A(regs_8[23]), .Z(n_27670));
	notech_inv i_30940(.A(regs_8[24]), .Z(n_27671));
	notech_inv i_30941(.A(regs_8[25]), .Z(n_27672));
	notech_inv i_30942(.A(regs_8[26]), .Z(n_27673));
	notech_inv i_30943(.A(regs_8[27]), .Z(n_27674));
	notech_inv i_30944(.A(regs_8[28]), .Z(n_27676));
	notech_inv i_30945(.A(regs_8[29]), .Z(n_27677));
	notech_inv i_30946(.A(regs_8[30]), .Z(n_27679));
	notech_inv i_30947(.A(regs_8[31]), .Z(n_27680));
	notech_inv i_30948(.A(regs_6[0]), .Z(n_27681));
	notech_inv i_30949(.A(regs_6[1]), .Z(n_27682));
	notech_inv i_30950(.A(regs_6[2]), .Z(n_27685));
	notech_inv i_30951(.A(regs_6[3]), .Z(n_27686));
	notech_inv i_30952(.A(regs_6[4]), .Z(n_27687));
	notech_inv i_30953(.A(regs_6[5]), .Z(n_27688));
	notech_inv i_30954(.A(regs_6[6]), .Z(n_27689));
	notech_inv i_30955(.A(regs_6[7]), .Z(n_27690));
	notech_inv i_30956(.A(regs_6[8]), .Z(n_27691));
	notech_inv i_30957(.A(regs_6[9]), .Z(n_27692));
	notech_inv i_30958(.A(regs_6[10]), .Z(n_27693));
	notech_inv i_30959(.A(regs_6[11]), .Z(n_27694));
	notech_inv i_30960(.A(regs_6[12]), .Z(n_27695));
	notech_inv i_30961(.A(regs_6[13]), .Z(n_27696));
	notech_inv i_30962(.A(regs_6[14]), .Z(n_27697));
	notech_inv i_30963(.A(regs_6[15]), .Z(n_27698));
	notech_inv i_30964(.A(regs_6[16]), .Z(n_27699));
	notech_inv i_30965(.A(regs_6[17]), .Z(n_27700));
	notech_inv i_30966(.A(regs_6[18]), .Z(n_27701));
	notech_inv i_30967(.A(regs_6[19]), .Z(n_27702));
	notech_inv i_30968(.A(regs_6[20]), .Z(n_27703));
	notech_inv i_30969(.A(regs_6[21]), .Z(n_27704));
	notech_inv i_30970(.A(regs_6[22]), .Z(n_27705));
	notech_inv i_30971(.A(regs_6[23]), .Z(n_27706));
	notech_inv i_30972(.A(regs_6[24]), .Z(n_27707));
	notech_inv i_30973(.A(regs_6[25]), .Z(n_27708));
	notech_inv i_30974(.A(regs_6[26]), .Z(n_27709));
	notech_inv i_30975(.A(regs_6[27]), .Z(n_27710));
	notech_inv i_30976(.A(regs_6[28]), .Z(n_27711));
	notech_inv i_30977(.A(regs_6[29]), .Z(n_27712));
	notech_inv i_30978(.A(regs_6[30]), .Z(n_27713));
	notech_inv i_30979(.A(regs_6[31]), .Z(n_27714));
	notech_inv i_30980(.A(regs_5[0]), .Z(n_27715));
	notech_inv i_30981(.A(regs_5[1]), .Z(n_27716));
	notech_inv i_30982(.A(regs_5[2]), .Z(n_27717));
	notech_inv i_30983(.A(regs_5[3]), .Z(n_27718));
	notech_inv i_30984(.A(regs_5[4]), .Z(n_27719));
	notech_inv i_30985(.A(regs_5[5]), .Z(n_27720));
	notech_inv i_30986(.A(regs_5[6]), .Z(n_27721));
	notech_inv i_30987(.A(regs_5[7]), .Z(n_27722));
	notech_inv i_30988(.A(regs_5[8]), .Z(n_27723));
	notech_inv i_30989(.A(regs_5[9]), .Z(n_27724));
	notech_inv i_30990(.A(regs_5[10]), .Z(n_27725));
	notech_inv i_30991(.A(regs_5[11]), .Z(n_27726));
	notech_inv i_30992(.A(regs_5[12]), .Z(n_27727));
	notech_inv i_30993(.A(regs_5[13]), .Z(n_27728));
	notech_inv i_30994(.A(regs_5[14]), .Z(n_27729));
	notech_inv i_30995(.A(regs_5[15]), .Z(n_27730));
	notech_inv i_30996(.A(regs_5[16]), .Z(n_27731));
	notech_inv i_30997(.A(regs_5[17]), .Z(n_27732));
	notech_inv i_30998(.A(regs_5[18]), .Z(n_27733));
	notech_inv i_30999(.A(regs_5[19]), .Z(n_27734));
	notech_inv i_31000(.A(regs_5[20]), .Z(n_27735));
	notech_inv i_31001(.A(regs_5[21]), .Z(n_27736));
	notech_inv i_31002(.A(regs_5[22]), .Z(n_27737));
	notech_inv i_31003(.A(regs_5[23]), .Z(n_27738));
	notech_inv i_31004(.A(regs_5[24]), .Z(n_27739));
	notech_inv i_31005(.A(regs_5[25]), .Z(n_27740));
	notech_inv i_31006(.A(regs_5[26]), .Z(n_27741));
	notech_inv i_31007(.A(regs_5[27]), .Z(n_27742));
	notech_inv i_31008(.A(regs_5[28]), .Z(n_27743));
	notech_inv i_31009(.A(regs_5[29]), .Z(n_27744));
	notech_inv i_31010(.A(regs_5[30]), .Z(n_27745));
	notech_inv i_31011(.A(regs_5[31]), .Z(n_27746));
	notech_inv i_31012(.A(regs_3[0]), .Z(n_27747));
	notech_inv i_31013(.A(regs_3[1]), .Z(n_27748));
	notech_inv i_31014(.A(regs_3[2]), .Z(n_27749));
	notech_inv i_31015(.A(regs_3[3]), .Z(n_27750));
	notech_inv i_31017(.A(regs_3[4]), .Z(n_27751));
	notech_inv i_31018(.A(regs_3[5]), .Z(n_27752));
	notech_inv i_31019(.A(regs_3[6]), .Z(n_27753));
	notech_inv i_31020(.A(regs_3[7]), .Z(n_27754));
	notech_inv i_31021(.A(regs_3[8]), .Z(n_27755));
	notech_inv i_31022(.A(regs_3[9]), .Z(n_27756));
	notech_inv i_31023(.A(regs_3[10]), .Z(n_27757));
	notech_inv i_31024(.A(regs_3[11]), .Z(n_27758));
	notech_inv i_31025(.A(regs_3[12]), .Z(n_27760));
	notech_inv i_31026(.A(regs_3[13]), .Z(n_27761));
	notech_inv i_31027(.A(regs_3[14]), .Z(n_27763));
	notech_inv i_31028(.A(regs_3[15]), .Z(n_27764));
	notech_inv i_31029(.A(regs_3[16]), .Z(n_27766));
	notech_inv i_31030(.A(regs_3[17]), .Z(n_27768));
	notech_inv i_31031(.A(regs_3[18]), .Z(n_27769));
	notech_inv i_31032(.A(regs_3[19]), .Z(n_27770));
	notech_inv i_31033(.A(regs_3[20]), .Z(n_27772));
	notech_inv i_31034(.A(regs_3[21]), .Z(n_27773));
	notech_inv i_31035(.A(regs_3[22]), .Z(n_27774));
	notech_inv i_31036(.A(regs_3[23]), .Z(n_27777));
	notech_inv i_31037(.A(regs_3[24]), .Z(n_27778));
	notech_inv i_31038(.A(regs_3[25]), .Z(n_27779));
	notech_inv i_31039(.A(regs_3[26]), .Z(n_27780));
	notech_inv i_31040(.A(regs_3[27]), .Z(n_27781));
	notech_inv i_31041(.A(regs_3[28]), .Z(n_27782));
	notech_inv i_31042(.A(regs_3[29]), .Z(n_27783));
	notech_inv i_31043(.A(regs_3[30]), .Z(n_27784));
	notech_inv i_31044(.A(regs_3[31]), .Z(n_27785));
	notech_inv i_31045(.A(regs_14[0]), .Z(n_27786));
	notech_inv i_31046(.A(regs_14[1]), .Z(n_27787));
	notech_inv i_31047(.A(regs_14[2]), .Z(n_27788));
	notech_inv i_31048(.A(regs_14[3]), .Z(n_27789));
	notech_inv i_31049(.A(regs_14[4]), .Z(n_27790));
	notech_inv i_31050(.A(regs_14[5]), .Z(n_27791));
	notech_inv i_31051(.A(regs_14[6]), .Z(n_27792));
	notech_inv i_31052(.A(regs_14[7]), .Z(n_27793));
	notech_inv i_31053(.A(regs_14[8]), .Z(n_27794));
	notech_inv i_31054(.A(regs_14[9]), .Z(n_27795));
	notech_inv i_31055(.A(regs_14[10]), .Z(n_27796));
	notech_inv i_31056(.A(regs_14[11]), .Z(n_27797));
	notech_inv i_31057(.A(regs_14[12]), .Z(n_27798));
	notech_inv i_31058(.A(regs_14[13]), .Z(n_27799));
	notech_inv i_31059(.A(regs_14[14]), .Z(n_27800));
	notech_inv i_31060(.A(regs_14[15]), .Z(n_27801));
	notech_inv i_31061(.A(regs_14[16]), .Z(n_27802));
	notech_inv i_31062(.A(regs_14[17]), .Z(n_27803));
	notech_inv i_31063(.A(regs_14[18]), .Z(n_27804));
	notech_inv i_31064(.A(regs_14[19]), .Z(n_27805));
	notech_inv i_31065(.A(regs_14[20]), .Z(n_27806));
	notech_inv i_31066(.A(regs_14[21]), .Z(n_27807));
	notech_inv i_31067(.A(regs_14[22]), .Z(n_27808));
	notech_inv i_31068(.A(regs_14[23]), .Z(n_27809));
	notech_inv i_31069(.A(regs_14[24]), .Z(n_27810));
	notech_inv i_31070(.A(regs_14[25]), .Z(n_27811));
	notech_inv i_31071(.A(regs_14[26]), .Z(n_27812));
	notech_inv i_31072(.A(regs_14[27]), .Z(n_27813));
	notech_inv i_31073(.A(regs_14[28]), .Z(n_27814));
	notech_inv i_31074(.A(regs_14[29]), .Z(n_27815));
	notech_inv i_31075(.A(regs_14[30]), .Z(n_27816));
	notech_inv i_31076(.A(regs_14[31]), .Z(n_27817));
	notech_inv i_31077(.A(regs_2[0]), .Z(n_27818));
	notech_inv i_31078(.A(regs_2[1]), .Z(n_27819));
	notech_inv i_31079(.A(regs_2[2]), .Z(n_27820));
	notech_inv i_31080(.A(regs_2[3]), .Z(n_27821));
	notech_inv i_31081(.A(regs_2[4]), .Z(n_27822));
	notech_inv i_31082(.A(regs_2[5]), .Z(n_27823));
	notech_inv i_31083(.A(regs_2[6]), .Z(n_27824));
	notech_inv i_31084(.A(regs_2[7]), .Z(n_27825));
	notech_inv i_31085(.A(regs_2[8]), .Z(n_27826));
	notech_inv i_31086(.A(regs_2[9]), .Z(n_27827));
	notech_inv i_31087(.A(regs_2[10]), .Z(n_27828));
	notech_inv i_31088(.A(regs_2[11]), .Z(n_27829));
	notech_inv i_31089(.A(regs_2[12]), .Z(n_27830));
	notech_inv i_31090(.A(regs_2[13]), .Z(n_27831));
	notech_inv i_31091(.A(regs_2[14]), .Z(n_27832));
	notech_inv i_31092(.A(regs_2[15]), .Z(n_27833));
	notech_inv i_31093(.A(regs_2[16]), .Z(n_27834));
	notech_inv i_31094(.A(regs_2[17]), .Z(n_27835));
	notech_inv i_31095(.A(regs_2[18]), .Z(n_27836));
	notech_inv i_31096(.A(regs_2[19]), .Z(n_27837));
	notech_inv i_31097(.A(regs_2[20]), .Z(n_27838));
	notech_inv i_31098(.A(regs_2[21]), .Z(n_27839));
	notech_inv i_31099(.A(regs_2[22]), .Z(n_27840));
	notech_inv i_31100(.A(regs_2[23]), .Z(n_27841));
	notech_inv i_31101(.A(regs_2[24]), .Z(n_27842));
	notech_inv i_31102(.A(regs_2[25]), .Z(n_27843));
	notech_inv i_31103(.A(regs_2[26]), .Z(n_27844));
	notech_inv i_31104(.A(regs_2[27]), .Z(n_27845));
	notech_inv i_31105(.A(regs_2[28]), .Z(n_27846));
	notech_inv i_31106(.A(regs_2[29]), .Z(n_27847));
	notech_inv i_31107(.A(regs_2[30]), .Z(n_27848));
	notech_inv i_31108(.A(regs_2[31]), .Z(n_27849));
	notech_inv i_31109(.A(regs_10[0]), .Z(n_27850));
	notech_inv i_31110(.A(regs_10[1]), .Z(n_27851));
	notech_inv i_31111(.A(regs_10[2]), .Z(n_27852));
	notech_inv i_31112(.A(regs_10[3]), .Z(n_27853));
	notech_inv i_31113(.A(regs_10[4]), .Z(n_27854));
	notech_inv i_31114(.A(regs_10[5]), .Z(n_27855));
	notech_inv i_31115(.A(regs_10[6]), .Z(n_27856));
	notech_inv i_31116(.A(regs_10[7]), .Z(n_27857));
	notech_inv i_31117(.A(regs_10[8]), .Z(n_27858));
	notech_inv i_31118(.A(regs_10[9]), .Z(n_27859));
	notech_inv i_31119(.A(regs_10[10]), .Z(n_27860));
	notech_inv i_31120(.A(regs_10[11]), .Z(n_27861));
	notech_inv i_31122(.A(regs_10[12]), .Z(n_27862));
	notech_inv i_31123(.A(regs_10[13]), .Z(n_27863));
	notech_inv i_31124(.A(regs_10[14]), .Z(n_27864));
	notech_inv i_31125(.A(regs_10[15]), .Z(n_27866));
	notech_inv i_31126(.A(regs_10[16]), .Z(n_27867));
	notech_inv i_31127(.A(regs_10[17]), .Z(n_27868));
	notech_inv i_31128(.A(regs_10[18]), .Z(n_27870));
	notech_inv i_31129(.A(regs_10[19]), .Z(n_27871));
	notech_inv i_31130(.A(regs_10[20]), .Z(n_27872));
	notech_inv i_31131(.A(regs_10[21]), .Z(n_27873));
	notech_inv i_31132(.A(regs_10[22]), .Z(n_27874));
	notech_inv i_31133(.A(regs_10[23]), .Z(n_27875));
	notech_inv i_31134(.A(regs_10[24]), .Z(n_27877));
	notech_inv i_31136(.A(regs_10[25]), .Z(n_27878));
	notech_inv i_31137(.A(regs_10[26]), .Z(n_27879));
	notech_inv i_31138(.A(regs_10[27]), .Z(n_27880));
	notech_inv i_31139(.A(regs_10[28]), .Z(n_27881));
	notech_inv i_31140(.A(regs_10[29]), .Z(n_27882));
	notech_inv i_31141(.A(regs_10[30]), .Z(n_27883));
	notech_inv i_31142(.A(regs_10[31]), .Z(n_27884));
	notech_inv i_31143(.A(regs_0[0]), .Z(n_27885));
	notech_inv i_31144(.A(regs_0[1]), .Z(n_27886));
	notech_inv i_31145(.A(regs_0[2]), .Z(n_27887));
	notech_inv i_31146(.A(regs_0[3]), .Z(n_27888));
	notech_inv i_31147(.A(regs_0[4]), .Z(n_27889));
	notech_inv i_31148(.A(regs_0[5]), .Z(n_27891));
	notech_inv i_31149(.A(regs_0[6]), .Z(n_27893));
	notech_inv i_31150(.A(regs_0[7]), .Z(n_27894));
	notech_inv i_31151(.A(regs_0[8]), .Z(n_27895));
	notech_inv i_31152(.A(regs_0[9]), .Z(n_27896));
	notech_inv i_31153(.A(regs_0[10]), .Z(n_27897));
	notech_inv i_31154(.A(regs_0[11]), .Z(n_27898));
	notech_inv i_31155(.A(regs_0[12]), .Z(n_27899));
	notech_inv i_31156(.A(regs_0[13]), .Z(n_27900));
	notech_inv i_31157(.A(regs_0[14]), .Z(n_27901));
	notech_inv i_31158(.A(regs_0[15]), .Z(n_27902));
	notech_inv i_31159(.A(regs_0[16]), .Z(n_27903));
	notech_inv i_31160(.A(regs_0[17]), .Z(n_27904));
	notech_inv i_31161(.A(regs_0[18]), .Z(n_27905));
	notech_inv i_31162(.A(regs_0[19]), .Z(n_27906));
	notech_inv i_31163(.A(regs_0[20]), .Z(n_27907));
	notech_inv i_31164(.A(regs_0[21]), .Z(n_27908));
	notech_inv i_31165(.A(regs_0[22]), .Z(n_27909));
	notech_inv i_31166(.A(regs_0[23]), .Z(n_27910));
	notech_inv i_31167(.A(regs_0[24]), .Z(n_27911));
	notech_inv i_31168(.A(regs_0[25]), .Z(n_27912));
	notech_inv i_31169(.A(regs_0[26]), .Z(n_27913));
	notech_inv i_31170(.A(regs_0[27]), .Z(n_27914));
	notech_inv i_31171(.A(regs_0[28]), .Z(n_27915));
	notech_inv i_31172(.A(regs_0[29]), .Z(n_27916));
	notech_inv i_31173(.A(regs_0[30]), .Z(n_27917));
	notech_inv i_31174(.A(regs_0[31]), .Z(n_27918));
	notech_inv i_31175(.A(regs_11[0]), .Z(n_27919));
	notech_inv i_31176(.A(regs_11[1]), .Z(n_27920));
	notech_inv i_31177(.A(regs_11[2]), .Z(n_27921));
	notech_inv i_31178(.A(regs_11[3]), .Z(n_27922));
	notech_inv i_31179(.A(regs_11[4]), .Z(n_27923));
	notech_inv i_31180(.A(regs_11[5]), .Z(n_27924));
	notech_inv i_31181(.A(regs_11[6]), .Z(n_27925));
	notech_inv i_31182(.A(regs_11[7]), .Z(n_27926));
	notech_inv i_31183(.A(regs_11[8]), .Z(n_27927));
	notech_inv i_31184(.A(regs_11[9]), .Z(n_27928));
	notech_inv i_31185(.A(regs_11[10]), .Z(n_27929));
	notech_inv i_31186(.A(regs_11[11]), .Z(n_27930));
	notech_inv i_31187(.A(regs_11[12]), .Z(n_27931));
	notech_inv i_31188(.A(regs_11[13]), .Z(n_27932));
	notech_inv i_31189(.A(regs_11[14]), .Z(n_27933));
	notech_inv i_31190(.A(regs_11[15]), .Z(n_27934));
	notech_inv i_31191(.A(regs_11[16]), .Z(n_27935));
	notech_inv i_31192(.A(regs_11[17]), .Z(n_27937));
	notech_inv i_31193(.A(regs_11[18]), .Z(n_27938));
	notech_inv i_31194(.A(regs_11[19]), .Z(n_27939));
	notech_inv i_31195(.A(regs_11[20]), .Z(n_27940));
	notech_inv i_31196(.A(regs_11[21]), .Z(n_27942));
	notech_inv i_31197(.A(regs_11[22]), .Z(n_27943));
	notech_inv i_31198(.A(regs_11[23]), .Z(n_27944));
	notech_inv i_31199(.A(regs_11[24]), .Z(n_27945));
	notech_inv i_31200(.A(regs_11[25]), .Z(n_27946));
	notech_inv i_31201(.A(regs_11[26]), .Z(n_27947));
	notech_inv i_31202(.A(regs_11[27]), .Z(n_27948));
	notech_inv i_31203(.A(regs_11[28]), .Z(n_27949));
	notech_inv i_31204(.A(regs_11[29]), .Z(n_27950));
	notech_inv i_31205(.A(regs_11[30]), .Z(n_27951));
	notech_inv i_31206(.A(regs_11[31]), .Z(n_27952));
	notech_inv i_31207(.A(regs_4[0]), .Z(n_27953));
	notech_inv i_31208(.A(regs_4[1]), .Z(n_27954));
	notech_inv i_31209(.A(regs_4[2]), .Z(n_27955));
	notech_inv i_31210(.A(regs_4[3]), .Z(n_27956));
	notech_inv i_31211(.A(regs_4[4]), .Z(n_27957));
	notech_inv i_31212(.A(regs_4[5]), .Z(n_27958));
	notech_inv i_31213(.A(regs_4[6]), .Z(n_27959));
	notech_inv i_31214(.A(regs_4[7]), .Z(n_27960));
	notech_inv i_31215(.A(regs_4[8]), .Z(n_27961));
	notech_inv i_31216(.A(regs_4[9]), .Z(n_27962));
	notech_inv i_31217(.A(regs_4[10]), .Z(n_27963));
	notech_inv i_31218(.A(regs_4[11]), .Z(n_27964));
	notech_inv i_31219(.A(regs_4[12]), .Z(n_27965));
	notech_inv i_31220(.A(regs_4[13]), .Z(n_27966));
	notech_inv i_31221(.A(regs_4[14]), .Z(n_27967));
	notech_inv i_31222(.A(regs_4[15]), .Z(n_27968));
	notech_inv i_31223(.A(regs_4[16]), .Z(n_27969));
	notech_inv i_31224(.A(regs_4[17]), .Z(n_27970));
	notech_inv i_31225(.A(regs_4[18]), .Z(n_27971));
	notech_inv i_31226(.A(regs_4[19]), .Z(n_27972));
	notech_inv i_31227(.A(regs_4[20]), .Z(n_27973));
	notech_inv i_31228(.A(regs_4[21]), .Z(n_27974));
	notech_inv i_31229(.A(regs_4[22]), .Z(n_27975));
	notech_inv i_31230(.A(regs_4[23]), .Z(n_27976));
	notech_inv i_31231(.A(regs_4[24]), .Z(n_27977));
	notech_inv i_31232(.A(regs_4[25]), .Z(n_27978));
	notech_inv i_31233(.A(regs_4[26]), .Z(n_27979));
	notech_inv i_31234(.A(regs_4[27]), .Z(n_27980));
	notech_inv i_31235(.A(regs_4[28]), .Z(n_27981));
	notech_inv i_31236(.A(regs_4[29]), .Z(n_27982));
	notech_inv i_31237(.A(regs_4[30]), .Z(n_27983));
	notech_inv i_31238(.A(regs_4[31]), .Z(n_27984));
	notech_inv i_31239(.A(gs[0]), .Z(n_27985));
	notech_inv i_31240(.A(gs[1]), .Z(n_27986));
	notech_inv i_31241(.A(n_55322), .Z(n_27987));
	notech_inv i_31242(.A(gs[3]), .Z(n_27988));
	notech_inv i_31243(.A(gs[4]), .Z(n_27989));
	notech_inv i_31244(.A(gs[5]), .Z(n_27990));
	notech_inv i_31245(.A(gs[6]), .Z(n_27991));
	notech_inv i_31246(.A(gs[7]), .Z(n_27992));
	notech_inv i_31247(.A(gs[8]), .Z(n_27993));
	notech_inv i_31248(.A(gs[9]), .Z(n_27994));
	notech_inv i_31249(.A(gs[10]), .Z(n_27995));
	notech_inv i_31250(.A(gs[11]), .Z(n_27996));
	notech_inv i_31251(.A(gs[12]), .Z(n_27997));
	notech_inv i_31252(.A(gs[13]), .Z(n_27998));
	notech_inv i_31253(.A(gs[14]), .Z(n_27999));
	notech_inv i_31254(.A(gs[15]), .Z(n_28000));
	notech_inv i_31255(.A(gs[16]), .Z(n_28001));
	notech_inv i_31256(.A(gs[17]), .Z(n_28002));
	notech_inv i_31257(.A(gs[18]), .Z(n_28003));
	notech_inv i_31258(.A(gs[19]), .Z(n_28006));
	notech_inv i_31259(.A(gs[20]), .Z(n_28007));
	notech_inv i_31260(.A(gs[21]), .Z(n_28008));
	notech_inv i_31261(.A(gs[22]), .Z(n_28009));
	notech_inv i_31262(.A(gs[23]), .Z(n_28010));
	notech_inv i_31263(.A(gs[24]), .Z(n_28011));
	notech_inv i_31264(.A(gs[25]), .Z(n_28012));
	notech_inv i_31265(.A(gs[26]), .Z(n_28013));
	notech_inv i_31266(.A(gs[27]), .Z(n_28014));
	notech_inv i_31267(.A(gs[28]), .Z(n_28015));
	notech_inv i_31268(.A(gs[29]), .Z(n_28016));
	notech_inv i_31269(.A(gs[30]), .Z(n_28017));
	notech_inv i_31270(.A(gs[31]), .Z(n_28018));
	notech_inv i_31271(.A(regs_7[0]), .Z(n_28019));
	notech_inv i_31272(.A(regs_7[1]), .Z(n_28020));
	notech_inv i_31273(.A(regs_7[2]), .Z(n_28021));
	notech_inv i_31274(.A(regs_7[3]), .Z(n_28022));
	notech_inv i_31275(.A(regs_7[4]), .Z(n_28023));
	notech_inv i_31276(.A(regs_7[5]), .Z(n_28024));
	notech_inv i_31277(.A(regs_7[6]), .Z(n_28025));
	notech_inv i_31278(.A(regs_7[7]), .Z(n_28026));
	notech_inv i_31279(.A(regs_7[8]), .Z(n_28027));
	notech_inv i_31280(.A(regs_7[9]), .Z(n_28028));
	notech_inv i_31281(.A(regs_7[10]), .Z(n_28029));
	notech_inv i_31282(.A(regs_7[11]), .Z(n_28030));
	notech_inv i_31283(.A(regs_7[12]), .Z(n_28031));
	notech_inv i_31284(.A(regs_7[13]), .Z(n_28032));
	notech_inv i_31285(.A(regs_7[14]), .Z(n_28033));
	notech_inv i_31286(.A(regs_7[15]), .Z(n_28034));
	notech_inv i_31287(.A(regs_7[16]), .Z(n_28035));
	notech_inv i_31288(.A(regs_7[17]), .Z(n_28036));
	notech_inv i_31289(.A(regs_7[18]), .Z(n_28037));
	notech_inv i_31290(.A(regs_7[19]), .Z(n_28038));
	notech_inv i_31291(.A(regs_7[20]), .Z(n_28039));
	notech_inv i_31292(.A(regs_7[21]), .Z(n_28040));
	notech_inv i_31293(.A(regs_7[22]), .Z(n_28041));
	notech_inv i_31294(.A(regs_7[23]), .Z(n_28042));
	notech_inv i_31295(.A(regs_7[24]), .Z(n_28043));
	notech_inv i_31296(.A(regs_7[25]), .Z(n_28044));
	notech_inv i_31297(.A(regs_7[26]), .Z(n_28045));
	notech_inv i_31298(.A(regs_7[27]), .Z(n_28046));
	notech_inv i_31299(.A(regs_7[28]), .Z(n_28047));
	notech_inv i_31300(.A(regs_7[29]), .Z(n_28048));
	notech_inv i_31301(.A(regs_7[30]), .Z(n_28049));
	notech_inv i_31302(.A(regs_7[31]), .Z(n_28050));
	notech_inv i_31303(.A(opc_10[0]), .Z(n_28051));
	notech_inv i_31304(.A(opc_10[1]), .Z(n_28052));
	notech_inv i_31305(.A(opc_10[2]), .Z(n_28053));
	notech_inv i_31306(.A(opc_10[3]), .Z(n_28054));
	notech_inv i_31307(.A(opc_10[4]), .Z(n_28055));
	notech_inv i_31308(.A(opc_10[5]), .Z(n_28056));
	notech_inv i_31309(.A(opc_10[6]), .Z(n_28057));
	notech_inv i_31310(.A(opc_10[7]), .Z(n_28058));
	notech_inv i_31311(.A(opc_10[8]), .Z(n_28059));
	notech_inv i_31312(.A(opc_10[9]), .Z(n_28060));
	notech_inv i_31313(.A(opc_10[10]), .Z(n_28061));
	notech_inv i_31314(.A(opc_10[11]), .Z(n_28062));
	notech_inv i_31315(.A(opc_10[12]), .Z(n_28063));
	notech_inv i_31316(.A(opc_10[13]), .Z(n_28064));
	notech_inv i_31317(.A(opc_10[14]), .Z(n_28065));
	notech_inv i_31318(.A(opc_10[15]), .Z(n_28066));
	notech_inv i_31319(.A(opc_10[16]), .Z(n_28067));
	notech_inv i_31320(.A(opc_10[17]), .Z(n_28068));
	notech_inv i_31321(.A(opc_10[18]), .Z(n_28069));
	notech_inv i_31322(.A(opc_10[19]), .Z(n_28070));
	notech_inv i_31323(.A(opc_10[20]), .Z(n_28071));
	notech_inv i_31324(.A(opc_10[21]), .Z(n_28072));
	notech_inv i_31325(.A(opc_10[22]), .Z(n_28073));
	notech_inv i_31326(.A(opc_10[23]), .Z(n_28074));
	notech_inv i_31327(.A(opc_10[24]), .Z(n_28075));
	notech_inv i_31328(.A(opc_10[25]), .Z(n_28076));
	notech_inv i_31329(.A(opc_10[26]), .Z(n_28077));
	notech_inv i_31330(.A(opc_10[27]), .Z(n_28078));
	notech_inv i_31331(.A(opc_10[28]), .Z(n_28079));
	notech_inv i_31333(.A(opc_10[29]), .Z(n_28080));
	notech_inv i_31334(.A(opc_10[30]), .Z(n_28081));
	notech_inv i_31335(.A(opc_10[31]), .Z(n_28082));
	notech_inv i_31336(.A(nbus_11279[0]), .Z(n_28083));
	notech_inv i_31337(.A(nbus_11279[1]), .Z(n_28084));
	notech_inv i_31338(.A(nbus_11279[2]), .Z(n_28085));
	notech_inv i_31339(.A(nbus_11279[3]), .Z(n_28086));
	notech_inv i_31340(.A(nbus_11279[4]), .Z(n_28087));
	notech_inv i_31341(.A(nbus_11279[5]), .Z(n_28088));
	notech_inv i_31342(.A(nbus_11279[6]), .Z(n_28089));
	notech_inv i_31343(.A(nbus_11279[7]), .Z(n_28090));
	notech_inv i_31344(.A(nbus_11279[8]), .Z(n_28091));
	notech_inv i_31345(.A(nbus_11279[9]), .Z(n_28092));
	notech_inv i_31346(.A(nbus_11279[10]), .Z(n_28093));
	notech_inv i_31347(.A(nbus_11279[11]), .Z(n_28094));
	notech_inv i_31348(.A(nbus_11279[12]), .Z(n_28095));
	notech_inv i_31349(.A(nbus_11279[13]), .Z(n_28096));
	notech_inv i_31350(.A(nbus_11279[14]), .Z(n_28097));
	notech_inv i_31351(.A(nbus_11279[15]), .Z(n_28098));
	notech_inv i_31352(.A(nbus_11279[16]), .Z(n_28099));
	notech_inv i_31353(.A(nbus_11279[17]), .Z(n_28100));
	notech_inv i_31354(.A(nbus_11279[18]), .Z(n_28101));
	notech_inv i_31355(.A(nbus_11279[19]), .Z(n_28102));
	notech_inv i_31356(.A(nbus_11279[20]), .Z(n_28103));
	notech_inv i_31357(.A(nbus_11279[21]), .Z(n_28104));
	notech_inv i_31358(.A(nbus_11279[22]), .Z(n_28105));
	notech_inv i_31359(.A(nbus_11279[23]), .Z(n_28106));
	notech_inv i_31360(.A(nbus_11279[24]), .Z(n_28107));
	notech_inv i_31361(.A(nbus_11279[25]), .Z(n_28108));
	notech_inv i_31362(.A(nbus_11279[26]), .Z(n_28109));
	notech_inv i_31363(.A(nbus_11279[27]), .Z(n_28110));
	notech_inv i_31364(.A(nbus_11279[28]), .Z(n_28111));
	notech_inv i_31365(.A(nbus_11279[29]), .Z(n_28112));
	notech_inv i_31366(.A(nbus_11279[30]), .Z(n_28113));
	notech_inv i_31367(.A(nbus_11279[31]), .Z(n_28114));
	notech_inv i_31368(.A(nbus_136[0]), .Z(n_28115));
	notech_inv i_31369(.A(nbus_136[1]), .Z(n_28116));
	notech_inv i_31370(.A(nbus_136[2]), .Z(n_28117));
	notech_inv i_31371(.A(nbus_136[3]), .Z(n_28118));
	notech_inv i_31372(.A(nbus_136[4]), .Z(n_28119));
	notech_inv i_31373(.A(nbus_136[5]), .Z(n_28120));
	notech_inv i_31374(.A(nbus_136[6]), .Z(n_28121));
	notech_inv i_31375(.A(nbus_136[7]), .Z(n_28122));
	notech_inv i_31376(.A(nbus_136[8]), .Z(n_28123));
	notech_inv i_31377(.A(nbus_142[0]), .Z(n_28124));
	notech_inv i_31378(.A(nbus_142[1]), .Z(n_28125));
	notech_inv i_31379(.A(nbus_142[2]), .Z(n_28126));
	notech_inv i_31380(.A(nbus_142[3]), .Z(n_28127));
	notech_inv i_31381(.A(nbus_142[4]), .Z(n_28128));
	notech_inv i_31382(.A(nbus_142[5]), .Z(n_28129));
	notech_inv i_31383(.A(nbus_142[6]), .Z(n_28130));
	notech_inv i_31384(.A(nbus_142[7]), .Z(n_28131));
	notech_inv i_31385(.A(nbus_142[8]), .Z(n_28132));
	notech_inv i_31386(.A(nbus_142[9]), .Z(n_28133));
	notech_inv i_31387(.A(nbus_142[10]), .Z(n_28134));
	notech_inv i_31388(.A(nbus_142[11]), .Z(n_28135));
	notech_inv i_31389(.A(nbus_142[12]), .Z(n_28136));
	notech_inv i_31390(.A(nbus_142[14]), .Z(n_28137));
	notech_inv i_31391(.A(nbus_142[15]), .Z(n_28138));
	notech_inv i_31392(.A(nbus_142[16]), .Z(n_28139));
	notech_inv i_31393(.A(n_60130), .Z(n_28140));
	notech_inv i_31396(.A(cr0[2]), .Z(n_28141));
	notech_inv i_31398(.A(cr0[16]), .Z(n_28142));
	notech_inv i_31401(.A(readio_data[0]), .Z(n_28143));
	notech_inv i_31402(.A(readio_data[1]), .Z(n_28144));
	notech_inv i_31404(.A(readio_data[2]), .Z(n_28145));
	notech_inv i_31405(.A(readio_data[3]), .Z(n_28146));
	notech_inv i_31407(.A(readio_data[4]), .Z(n_28147));
	notech_inv i_31414(.A(readio_data[5]), .Z(n_28148));
	notech_inv i_31415(.A(readio_data[6]), .Z(n_28149));
	notech_inv i_31420(.A(readio_data[7]), .Z(n_28150));
	notech_inv i_31422(.A(readio_data[8]), .Z(n_28151));
	notech_inv i_31423(.A(readio_data[9]), .Z(n_28152));
	notech_inv i_31424(.A(readio_data[10]), .Z(n_28153));
	notech_inv i_31425(.A(readio_data[11]), .Z(n_28154));
	notech_inv i_31426(.A(readio_data[12]), .Z(n_28155));
	notech_inv i_31427(.A(readio_data[14]), .Z(n_28156));
	notech_inv i_31428(.A(readio_data[15]), .Z(n_28157));
	notech_inv i_31429(.A(readio_data[16]), .Z(n_28158));
	notech_inv i_31432(.A(readio_data[17]), .Z(n_28159));
	notech_inv i_31433(.A(readio_data[18]), .Z(n_28160));
	notech_inv i_31434(.A(readio_data[19]), .Z(n_28161));
	notech_inv i_31436(.A(readio_data[20]), .Z(n_28162));
	notech_inv i_31437(.A(readio_data[21]), .Z(n_28163));
	notech_inv i_31438(.A(readio_data[22]), .Z(n_28164));
	notech_inv i_31440(.A(readio_data[23]), .Z(n_28165));
	notech_inv i_31441(.A(readio_data[24]), .Z(n_28166));
	notech_inv i_31444(.A(readio_data[25]), .Z(n_28167));
	notech_inv i_31445(.A(readio_data[26]), .Z(n_28168));
	notech_inv i_31446(.A(readio_data[27]), .Z(n_28169));
	notech_inv i_31447(.A(readio_data[28]), .Z(n_28170));
	notech_inv i_31448(.A(readio_data[29]), .Z(n_28171));
	notech_inv i_31449(.A(readio_data[30]), .Z(n_28172));
	notech_inv i_31450(.A(readio_data[31]), .Z(n_28173));
	notech_inv i_31451(.A(resa_shiftbox[0]), .Z(n_28174));
	notech_inv i_31452(.A(resa_shiftbox[1]), .Z(n_28175));
	notech_inv i_31453(.A(resa_shiftbox[2]), .Z(n_28176));
	notech_inv i_31454(.A(resa_shiftbox[3]), .Z(n_28178));
	notech_inv i_31455(.A(resa_shiftbox[4]), .Z(n_28179));
	notech_inv i_31456(.A(resa_shiftbox[5]), .Z(n_28182));
	notech_inv i_31457(.A(resa_shiftbox[6]), .Z(n_28186));
	notech_inv i_31458(.A(resa_shiftbox[7]), .Z(n_28187));
	notech_inv i_31459(.A(resa_shiftbox[8]), .Z(n_28188));
	notech_inv i_31460(.A(resa_shiftbox[9]), .Z(n_28189));
	notech_inv i_31461(.A(resa_shiftbox[10]), .Z(n_28190));
	notech_inv i_31462(.A(resa_shiftbox[11]), .Z(n_28191));
	notech_inv i_31463(.A(resa_shiftbox[12]), .Z(n_28192));
	notech_inv i_31464(.A(resa_shiftbox[14]), .Z(n_28193));
	notech_inv i_31465(.A(resa_shiftbox[15]), .Z(n_28194));
	notech_inv i_31466(.A(resa_shiftbox[17]), .Z(n_28195));
	notech_inv i_31467(.A(resa_shiftbox[23]), .Z(n_28196));
	notech_inv i_31468(.A(cr3[13]), .Z(n_28198));
	notech_inv i_31469(.A(cr3[15]), .Z(n_28200));
	notech_inv i_31470(.A(cr3[17]), .Z(n_28202));
	notech_inv i_31471(.A(cr3[23]), .Z(n_28203));
	notech_inv i_31472(.A(resa_shift4box[0]), .Z(n_28204));
	notech_inv i_31473(.A(resa_shift4box[1]), .Z(n_28205));
	notech_inv i_31474(.A(resa_shift4box[2]), .Z(n_28206));
	notech_inv i_31475(.A(resa_shift4box[3]), .Z(n_28207));
	notech_inv i_31476(.A(resa_shift4box[4]), .Z(n_28208));
	notech_inv i_31477(.A(resa_shift4box[5]), .Z(n_28209));
	notech_inv i_31478(.A(resa_shift4box[6]), .Z(n_28210));
	notech_inv i_31479(.A(resa_shift4box[7]), .Z(n_28212));
	notech_inv i_31480(.A(resa_shift4box[8]), .Z(n_28213));
	notech_inv i_31481(.A(resa_shift4box[9]), .Z(n_28214));
	notech_inv i_31482(.A(resa_shift4box[10]), .Z(n_28215));
	notech_inv i_31483(.A(resa_shift4box[11]), .Z(n_28216));
	notech_inv i_31484(.A(resa_shift4box[12]), .Z(n_28217));
	notech_inv i_31485(.A(resa_shift4box[14]), .Z(n_28218));
	notech_inv i_31486(.A(resa_shift4box[15]), .Z(n_28219));
	notech_inv i_31487(.A(resa_shift4box[17]), .Z(n_28220));
	notech_inv i_31488(.A(resa_shift4box[23]), .Z(n_28221));
	notech_inv i_31489(.A(opa_0[0]), .Z(n_28222));
	notech_inv i_31490(.A(opa_0[1]), .Z(n_28223));
	notech_inv i_31491(.A(opa_0[2]), .Z(n_28224));
	notech_inv i_31492(.A(opa_0[3]), .Z(n_28225));
	notech_inv i_31493(.A(opa_0[4]), .Z(n_28226));
	notech_inv i_31494(.A(opa_0[5]), .Z(n_28227));
	notech_inv i_31495(.A(opa_0[6]), .Z(n_28228));
	notech_inv i_31496(.A(opa_0[7]), .Z(n_28229));
	notech_inv i_31497(.A(opa_0[8]), .Z(n_28230));
	notech_inv i_31498(.A(opa_0[9]), .Z(n_28231));
	notech_inv i_31499(.A(opa_0[10]), .Z(n_28232));
	notech_inv i_31500(.A(opa_0[11]), .Z(n_28233));
	notech_inv i_31501(.A(opa_0[12]), .Z(n_28234));
	notech_inv i_31502(.A(opa_0[14]), .Z(n_28235));
	notech_inv i_31503(.A(opa_0[15]), .Z(n_28236));
	notech_inv i_31504(.A(opa_0[16]), .Z(n_28237));
	notech_inv i_31505(.A(opa_0[17]), .Z(n_28238));
	notech_inv i_31506(.A(opa_0[18]), .Z(n_28239));
	notech_inv i_31507(.A(opa_0[19]), .Z(n_28240));
	notech_inv i_31508(.A(opa_0[20]), .Z(n_28241));
	notech_inv i_31509(.A(opa_0[21]), .Z(n_28242));
	notech_inv i_31510(.A(opa_0[22]), .Z(n_28243));
	notech_inv i_31511(.A(opa_0[23]), .Z(n_28244));
	notech_inv i_31512(.A(opa_0[24]), .Z(n_28245));
	notech_inv i_31513(.A(opa_0[25]), .Z(n_28246));
	notech_inv i_31514(.A(opa_0[26]), .Z(n_28247));
	notech_inv i_31515(.A(opa_0[27]), .Z(n_28248));
	notech_inv i_31516(.A(opa_0[28]), .Z(n_28249));
	notech_inv i_31517(.A(opa_0[29]), .Z(n_28250));
	notech_inv i_31518(.A(opa_0[30]), .Z(n_28251));
	notech_inv i_31519(.A(opa_0[31]), .Z(n_28252));
	notech_inv i_31520(.A(resa_arithbox[0]), .Z(n_28253));
	notech_inv i_31521(.A(resa_arithbox[1]), .Z(n_28254));
	notech_inv i_31522(.A(resa_arithbox[2]), .Z(n_28255));
	notech_inv i_31523(.A(resa_arithbox[3]), .Z(n_28256));
	notech_inv i_31524(.A(resa_arithbox[4]), .Z(n_28257));
	notech_inv i_31525(.A(resa_arithbox[5]), .Z(n_28258));
	notech_inv i_31526(.A(resa_arithbox[6]), .Z(n_28259));
	notech_inv i_31527(.A(resa_arithbox[7]), .Z(n_28260));
	notech_inv i_31528(.A(resa_arithbox[8]), .Z(n_28261));
	notech_inv i_31529(.A(resa_arithbox[9]), .Z(n_28262));
	notech_inv i_31530(.A(resa_arithbox[10]), .Z(n_28263));
	notech_inv i_31531(.A(resa_arithbox[11]), .Z(n_28264));
	notech_inv i_31532(.A(resa_arithbox[12]), .Z(n_28265));
	notech_inv i_31533(.A(resa_arithbox[14]), .Z(n_28266));
	notech_inv i_31534(.A(resa_arithbox[15]), .Z(n_28267));
	notech_inv i_31535(.A(nbus_139[0]), .Z(n_28268));
	notech_inv i_31536(.A(nbus_139[1]), .Z(n_28269));
	notech_inv i_31537(.A(nbus_139[2]), .Z(n_28270));
	notech_inv i_31538(.A(nbus_139[3]), .Z(n_28271));
	notech_inv i_31539(.A(nbus_139[4]), .Z(n_28272));
	notech_inv i_31540(.A(nbus_139[5]), .Z(n_28273));
	notech_inv i_31541(.A(nbus_139[6]), .Z(n_28274));
	notech_inv i_31542(.A(nbus_139[7]), .Z(n_28275));
	notech_inv i_31543(.A(nbus_139[8]), .Z(n_28276));
	notech_inv i_31544(.A(nbus_139[9]), .Z(n_28277));
	notech_inv i_31545(.A(nbus_139[10]), .Z(n_28278));
	notech_inv i_31546(.A(nbus_139[11]), .Z(n_28279));
	notech_inv i_31547(.A(nbus_139[12]), .Z(n_28280));
	notech_inv i_31548(.A(nbus_139[13]), .Z(n_28281));
	notech_inv i_31550(.A(nbus_139[14]), .Z(n_28282));
	notech_inv i_31551(.A(nbus_139[15]), .Z(n_28283));
	notech_inv i_31552(.A(nbus_139[16]), .Z(n_28284));
	notech_inv i_31554(.A(nbus_139[17]), .Z(n_28285));
	notech_inv i_31555(.A(nbus_139[18]), .Z(n_28286));
	notech_inv i_31556(.A(nbus_139[19]), .Z(n_28287));
	notech_inv i_31557(.A(nbus_139[20]), .Z(n_28288));
	notech_inv i_31558(.A(nbus_139[21]), .Z(n_28289));
	notech_inv i_31559(.A(nbus_139[22]), .Z(n_28292));
	notech_inv i_31560(.A(nbus_139[23]), .Z(n_28293));
	notech_inv i_31561(.A(nbus_139[24]), .Z(n_28294));
	notech_inv i_31562(.A(nbus_139[25]), .Z(n_28295));
	notech_inv i_31563(.A(nbus_139[26]), .Z(n_28296));
	notech_inv i_31564(.A(nbus_139[27]), .Z(n_28297));
	notech_inv i_31565(.A(nbus_139[28]), .Z(n_28298));
	notech_inv i_31566(.A(nbus_139[29]), .Z(n_28299));
	notech_inv i_31567(.A(nbus_139[30]), .Z(n_28300));
	notech_inv i_31568(.A(nbus_139[31]), .Z(n_28301));
	notech_inv i_31569(.A(nbus_139[32]), .Z(n_28302));
	notech_inv i_31570(.A(nbus_141[0]), .Z(n_28303));
	notech_inv i_31571(.A(nbus_141[1]), .Z(n_28304));
	notech_inv i_31572(.A(nbus_141[2]), .Z(n_28305));
	notech_inv i_31573(.A(nbus_141[3]), .Z(n_28306));
	notech_inv i_31574(.A(nbus_141[4]), .Z(n_28307));
	notech_inv i_31575(.A(nbus_141[5]), .Z(n_28308));
	notech_inv i_31576(.A(nbus_141[6]), .Z(n_28309));
	notech_inv i_31577(.A(nbus_141[7]), .Z(n_28310));
	notech_inv i_31578(.A(nbus_141[8]), .Z(n_28315));
	notech_inv i_31579(.A(nbus_141[9]), .Z(n_28316));
	notech_inv i_31580(.A(nbus_141[10]), .Z(n_28317));
	notech_inv i_31581(.A(nbus_141[11]), .Z(n_28318));
	notech_inv i_31582(.A(nbus_141[12]), .Z(n_28320));
	notech_inv i_31583(.A(nbus_141[13]), .Z(n_28321));
	notech_inv i_31584(.A(nbus_141[14]), .Z(n_28322));
	notech_inv i_31585(.A(nbus_141[15]), .Z(n_28323));
	notech_inv i_31586(.A(nbus_141[16]), .Z(n_28324));
	notech_inv i_31587(.A(nbus_141[17]), .Z(n_28325));
	notech_inv i_31588(.A(nbus_141[18]), .Z(n_28326));
	notech_inv i_31589(.A(nbus_141[19]), .Z(n_28327));
	notech_inv i_31590(.A(nbus_141[20]), .Z(n_28328));
	notech_inv i_31591(.A(nbus_141[21]), .Z(n_28329));
	notech_inv i_31592(.A(nbus_141[22]), .Z(n_28330));
	notech_inv i_31593(.A(nbus_141[23]), .Z(n_28331));
	notech_inv i_31594(.A(nbus_141[24]), .Z(n_28332));
	notech_inv i_31595(.A(nbus_141[25]), .Z(n_28333));
	notech_inv i_31596(.A(nbus_141[26]), .Z(n_28334));
	notech_inv i_31597(.A(nbus_141[27]), .Z(n_28335));
	notech_inv i_31598(.A(nbus_141[28]), .Z(n_28336));
	notech_inv i_31599(.A(nbus_141[29]), .Z(n_28337));
	notech_inv i_31600(.A(nbus_141[30]), .Z(n_28338));
	notech_inv i_31601(.A(nbus_141[31]), .Z(n_28339));
	notech_inv i_31602(.A(nbus_141[32]), .Z(n_28340));
	notech_inv i_31603(.A(nbus_134[0]), .Z(n_28341));
	notech_inv i_31604(.A(nbus_134[1]), .Z(n_28342));
	notech_inv i_31605(.A(nbus_134[2]), .Z(n_28343));
	notech_inv i_31606(.A(nbus_134[3]), .Z(n_28344));
	notech_inv i_31607(.A(nbus_134[4]), .Z(n_28345));
	notech_inv i_31608(.A(nbus_134[5]), .Z(n_28346));
	notech_inv i_31609(.A(nbus_134[6]), .Z(n_28347));
	notech_inv i_31610(.A(nbus_134[7]), .Z(n_28348));
	notech_inv i_31611(.A(nbus_134[8]), .Z(n_28349));
	notech_inv i_31613(.A(nbus_134[9]), .Z(n_28350));
	notech_inv i_31614(.A(nbus_134[10]), .Z(n_28351));
	notech_inv i_31616(.A(nbus_134[11]), .Z(n_28352));
	notech_inv i_31617(.A(nbus_134[12]), .Z(n_28353));
	notech_inv i_31618(.A(nbus_134[13]), .Z(n_28354));
	notech_inv i_31619(.A(nbus_134[14]), .Z(n_28355));
	notech_inv i_31620(.A(nbus_134[15]), .Z(n_28356));
	notech_inv i_31621(.A(nbus_134[16]), .Z(n_28357));
	notech_inv i_31622(.A(nbus_134[18]), .Z(n_28358));
	notech_inv i_31623(.A(nbus_134[19]), .Z(n_28359));
	notech_inv i_31624(.A(nbus_134[20]), .Z(n_28360));
	notech_inv i_31625(.A(nbus_134[21]), .Z(n_28361));
	notech_inv i_31626(.A(nbus_134[22]), .Z(n_28362));
	notech_inv i_31627(.A(nbus_134[24]), .Z(n_28363));
	notech_inv i_31628(.A(nbus_134[25]), .Z(n_28364));
	notech_inv i_31629(.A(nbus_134[26]), .Z(n_28365));
	notech_inv i_31630(.A(nbus_134[27]), .Z(n_28366));
	notech_inv i_31631(.A(nbus_134[28]), .Z(n_28367));
	notech_inv i_31632(.A(nbus_134[29]), .Z(n_28368));
	notech_inv i_31633(.A(nbus_134[30]), .Z(n_28369));
	notech_inv i_31634(.A(nbus_134[31]), .Z(n_28370));
	notech_inv i_31635(.A(nbus_134[32]), .Z(n_28371));
	notech_inv i_31636(.A(nbus_140[0]), .Z(n_28372));
	notech_inv i_31637(.A(nbus_140[1]), .Z(n_28373));
	notech_inv i_31638(.A(nbus_140[2]), .Z(n_28374));
	notech_inv i_31639(.A(nbus_140[3]), .Z(n_28375));
	notech_inv i_31640(.A(nbus_140[4]), .Z(n_28376));
	notech_inv i_31641(.A(nbus_140[5]), .Z(n_28377));
	notech_inv i_31642(.A(nbus_140[6]), .Z(n_28378));
	notech_inv i_31643(.A(nbus_140[7]), .Z(n_28379));
	notech_inv i_31644(.A(nbus_140[8]), .Z(n_28380));
	notech_inv i_31645(.A(nbus_140[9]), .Z(n_28381));
	notech_inv i_31646(.A(nbus_140[10]), .Z(n_28382));
	notech_inv i_31647(.A(nbus_140[11]), .Z(n_28383));
	notech_inv i_31648(.A(nbus_140[12]), .Z(n_28384));
	notech_inv i_31649(.A(nbus_140[14]), .Z(n_28385));
	notech_inv i_31650(.A(nbus_140[15]), .Z(n_28386));
	notech_inv i_31651(.A(nbus_135[0]), .Z(n_28387));
	notech_inv i_31652(.A(nbus_135[1]), .Z(n_28388));
	notech_inv i_31653(.A(nbus_135[2]), .Z(n_28389));
	notech_inv i_31654(.A(nbus_135[3]), .Z(n_28390));
	notech_inv i_31655(.A(nbus_135[4]), .Z(n_28391));
	notech_inv i_31656(.A(nbus_135[5]), .Z(n_28392));
	notech_inv i_31657(.A(nbus_135[6]), .Z(n_28393));
	notech_inv i_31658(.A(nbus_135[7]), .Z(n_28394));
	notech_inv i_31659(.A(nbus_135[8]), .Z(n_28395));
	notech_inv i_31660(.A(nbus_135[9]), .Z(n_28396));
	notech_inv i_31661(.A(nbus_135[10]), .Z(n_28397));
	notech_inv i_31662(.A(nbus_135[11]), .Z(n_28398));
	notech_inv i_31663(.A(nbus_135[12]), .Z(n_28399));
	notech_inv i_31664(.A(nbus_135[13]), .Z(n_28400));
	notech_inv i_31665(.A(nbus_135[14]), .Z(n_28401));
	notech_inv i_31666(.A(nbus_135[15]), .Z(n_28402));
	notech_inv i_31667(.A(nbus_138[0]), .Z(n_28403));
	notech_inv i_31668(.A(nbus_138[1]), .Z(n_28404));
	notech_inv i_31669(.A(nbus_138[3]), .Z(n_28405));
	notech_inv i_31670(.A(nbus_138[4]), .Z(n_28406));
	notech_inv i_31671(.A(nbus_138[5]), .Z(n_28407));
	notech_inv i_31672(.A(nbus_138[6]), .Z(n_28408));
	notech_inv i_31673(.A(nbus_138[7]), .Z(n_28409));
	notech_inv i_31674(.A(nbus_138[9]), .Z(n_28410));
	notech_inv i_31675(.A(nbus_138[15]), .Z(n_28411));
	notech_inv i_31676(.A(nbus_138[16]), .Z(n_28412));
	notech_inv i_31677(.A(over_seg[5]), .Z(n_28413));
	notech_inv i_31678(.A(regs_4_2[0]), .Z(n_28414));
	notech_inv i_31680(.A(regs_4_2[1]), .Z(n_28415));
	notech_inv i_31681(.A(regs_4_2[2]), .Z(n_28416));
	notech_inv i_31682(.A(regs_4_2[3]), .Z(n_28417));
	notech_inv i_31683(.A(regs_4_2[4]), .Z(n_28418));
	notech_inv i_31684(.A(regs_4_2[5]), .Z(n_28419));
	notech_inv i_31685(.A(regs_4_2[6]), .Z(n_28420));
	notech_inv i_31686(.A(regs_4_2[7]), .Z(n_28421));
	notech_inv i_31687(.A(regs_4_2[8]), .Z(n_28422));
	notech_inv i_31688(.A(regs_4_2[9]), .Z(n_28423));
	notech_inv i_31689(.A(regs_4_2[10]), .Z(n_28424));
	notech_inv i_31690(.A(regs_4_2[11]), .Z(n_28425));
	notech_inv i_31691(.A(regs_4_2[12]), .Z(n_28426));
	notech_inv i_31692(.A(regs_4_2[13]), .Z(n_28427));
	notech_inv i_31693(.A(regs_4_2[14]), .Z(n_28428));
	notech_inv i_31694(.A(regs_4_2[15]), .Z(n_28429));
	notech_inv i_31695(.A(regs_4_2[16]), .Z(n_28430));
	notech_inv i_31696(.A(regs_4_2[17]), .Z(n_28431));
	notech_inv i_31697(.A(regs_4_2[18]), .Z(n_28432));
	notech_inv i_31698(.A(regs_4_2[19]), .Z(n_28433));
	notech_inv i_31699(.A(regs_4_2[20]), .Z(n_28434));
	notech_inv i_31700(.A(regs_4_2[21]), .Z(n_28435));
	notech_inv i_31701(.A(regs_4_2[22]), .Z(n_28436));
	notech_inv i_31702(.A(regs_4_2[23]), .Z(n_28437));
	notech_inv i_31703(.A(regs_4_2[24]), .Z(n_28438));
	notech_inv i_31704(.A(regs_4_2[25]), .Z(n_28439));
	notech_inv i_31705(.A(regs_4_2[26]), .Z(n_28440));
	notech_inv i_31706(.A(regs_4_2[27]), .Z(n_28441));
	notech_inv i_31707(.A(regs_4_2[28]), .Z(n_28442));
	notech_inv i_31708(.A(regs_4_2[29]), .Z(n_28443));
	notech_inv i_31709(.A(regs_4_2[30]), .Z(n_28444));
	notech_inv i_31711(.A(regs_4_2[31]), .Z(n_28445));
	notech_inv i_31712(.A(Daddrs_1[1]), .Z(n_28446));
	notech_inv i_31713(.A(Daddrs_1[2]), .Z(n_28447));
	notech_inv i_31714(.A(Daddrs_1[3]), .Z(n_28448));
	notech_inv i_31715(.A(Daddrs_1[4]), .Z(n_28449));
	notech_inv i_31716(.A(Daddrs_1[5]), .Z(n_28450));
	notech_inv i_31717(.A(Daddrs_1[6]), .Z(n_28451));
	notech_inv i_31718(.A(Daddrs_1[7]), .Z(n_28452));
	notech_inv i_31721(.A(Daddrs_1[8]), .Z(n_28453));
	notech_inv i_31722(.A(Daddrs_1[31]), .Z(n_28454));
	notech_inv i_31724(.A(Daddrs_8[31]), .Z(n_28455));
	notech_inv i_31725(.A(Daddrs_3[0]), .Z(n_28456));
	notech_inv i_31726(.A(Daddrs_3[1]), .Z(n_28457));
	notech_inv i_31727(.A(Daddrs_3[2]), .Z(n_28459));
	notech_inv i_31728(.A(Daddrs_3[3]), .Z(n_28460));
	notech_inv i_31729(.A(Daddrs_3[4]), .Z(n_28461));
	notech_inv i_31730(.A(Daddrs_3[5]), .Z(n_28462));
	notech_inv i_31731(.A(Daddrs_3[6]), .Z(n_28463));
	notech_inv i_31732(.A(Daddrs_3[7]), .Z(n_28464));
	notech_inv i_31733(.A(Daddrs_3[8]), .Z(n_28466));
	notech_inv i_31734(.A(Daddrs_3[9]), .Z(n_28467));
	notech_inv i_31735(.A(Daddrs_3[10]), .Z(n_28468));
	notech_inv i_31736(.A(Daddrs_3[11]), .Z(n_28469));
	notech_inv i_31737(.A(Daddrs_3[12]), .Z(n_28470));
	notech_inv i_31738(.A(Daddrs_3[13]), .Z(n_28474));
	notech_inv i_31739(.A(Daddrs_3[14]), .Z(n_28475));
	notech_inv i_31740(.A(Daddrs_3[15]), .Z(n_28476));
	notech_inv i_31741(.A(Daddrs_3[16]), .Z(n_28478));
	notech_inv i_31742(.A(Daddrs_3[17]), .Z(n_28481));
	notech_inv i_31743(.A(Daddrs_3[18]), .Z(n_28486));
	notech_inv i_31744(.A(Daddrs_3[19]), .Z(n_28487));
	notech_inv i_31745(.A(Daddrs_3[20]), .Z(n_28488));
	notech_inv i_31746(.A(Daddrs_3[21]), .Z(n_28489));
	notech_inv i_31747(.A(Daddrs_3[22]), .Z(n_28490));
	notech_inv i_31748(.A(Daddrs_3[23]), .Z(n_28491));
	notech_inv i_31749(.A(Daddrs_3[24]), .Z(n_28492));
	notech_inv i_31750(.A(Daddrs_3[25]), .Z(n_28493));
	notech_inv i_31751(.A(Daddrs_3[26]), .Z(n_28494));
	notech_inv i_31752(.A(Daddrs_3[27]), .Z(n_28495));
	notech_inv i_31753(.A(Daddrs_3[28]), .Z(n_28496));
	notech_inv i_31754(.A(Daddrs_3[29]), .Z(n_28497));
	notech_inv i_31755(.A(Daddrs_3[30]), .Z(n_28498));
	notech_inv i_31756(.A(instrc[0]), .Z(n_28499));
	notech_inv i_31757(.A(instrc[1]), .Z(n_28500));
	notech_inv i_31758(.A(instrc[2]), .Z(n_28501));
	notech_inv i_31759(.A(instrc[3]), .Z(n_28502));
	notech_inv i_31760(.A(instrc[4]), .Z(n_28503));
	notech_inv i_31761(.A(instrc[5]), .Z(n_28504));
	notech_inv i_31762(.A(instrc[6]), .Z(n_28505));
	notech_inv i_31763(.A(instrc[7]), .Z(n_28506));
	notech_inv i_31764(.A(instrc[8]), .Z(n_28507));
	notech_inv i_31765(.A(instrc[9]), .Z(n_28508));
	notech_inv i_31766(.A(instrc[10]), .Z(n_28509));
	notech_inv i_31767(.A(instrc[11]), .Z(n_28510));
	notech_inv i_31768(.A(instrc[12]), .Z(n_28511));
	notech_inv i_31769(.A(instrc[13]), .Z(n_28512));
	notech_inv i_31770(.A(instrc[14]), .Z(n_28513));
	notech_inv i_31771(.A(instrc[15]), .Z(n_28514));
	notech_inv i_31772(.A(instrc[16]), .Z(n_28515));
	notech_inv i_31773(.A(instrc[17]), .Z(n_28516));
	notech_inv i_31774(.A(instrc[18]), .Z(n_28517));
	notech_inv i_31775(.A(instrc[19]), .Z(n_28518));
	notech_inv i_31776(.A(instrc[20]), .Z(n_28519));
	notech_inv i_31777(.A(instrc[21]), .Z(n_28520));
	notech_inv i_31778(.A(instrc[22]), .Z(n_28521));
	notech_inv i_31779(.A(instrc[23]), .Z(n_28522));
	notech_inv i_31780(.A(instrc[24]), .Z(n_28523));
	notech_inv i_31781(.A(instrc[25]), .Z(n_28524));
	notech_inv i_31782(.A(instrc[26]), .Z(n_28525));
	notech_inv i_31783(.A(instrc[27]), .Z(n_28526));
	notech_inv i_31784(.A(instrc[28]), .Z(n_28527));
	notech_inv i_31785(.A(instrc[29]), .Z(n_28528));
	notech_inv i_31786(.A(instrc[30]), .Z(n_28529));
	notech_inv i_31787(.A(instrc[31]), .Z(n_28530));
	notech_inv i_31788(.A(instrc[32]), .Z(n_28531));
	notech_inv i_31789(.A(instrc[33]), .Z(n_28532));
	notech_inv i_31790(.A(instrc[34]), .Z(n_28533));
	notech_inv i_31791(.A(instrc[35]), .Z(n_28534));
	notech_inv i_31792(.A(instrc[36]), .Z(n_28535));
	notech_inv i_31793(.A(instrc[37]), .Z(n_28536));
	notech_inv i_31794(.A(instrc[38]), .Z(n_28537));
	notech_inv i_31795(.A(instrc[39]), .Z(n_28538));
	notech_inv i_31796(.A(instrc[40]), .Z(n_28539));
	notech_inv i_31797(.A(instrc[41]), .Z(n_28540));
	notech_inv i_31798(.A(instrc[42]), .Z(n_28541));
	notech_inv i_31799(.A(instrc[43]), .Z(n_28542));
	notech_inv i_31800(.A(instrc[44]), .Z(n_28543));
	notech_inv i_31801(.A(instrc[45]), .Z(n_28544));
	notech_inv i_31802(.A(instrc[46]), .Z(n_28545));
	notech_inv i_31803(.A(instrc[47]), .Z(n_28546));
	notech_inv i_31804(.A(instrc[48]), .Z(n_28547));
	notech_inv i_31805(.A(instrc[49]), .Z(n_28548));
	notech_inv i_31806(.A(instrc[50]), .Z(n_28549));
	notech_inv i_31807(.A(instrc[51]), .Z(n_28550));
	notech_inv i_31808(.A(instrc[52]), .Z(n_28551));
	notech_inv i_31809(.A(instrc[53]), .Z(n_28552));
	notech_inv i_31810(.A(instrc[55]), .Z(n_28553));
	notech_inv i_31811(.A(instrc[72]), .Z(n_28554));
	notech_inv i_31812(.A(instrc[73]), .Z(n_28555));
	notech_inv i_31813(.A(instrc[74]), .Z(n_28556));
	notech_inv i_31814(.A(instrc[75]), .Z(n_28557));
	notech_inv i_31815(.A(instrc[76]), .Z(n_28558));
	notech_inv i_31816(.A(instrc[77]), .Z(n_28559));
	notech_inv i_31817(.A(instrc[78]), .Z(n_28560));
	notech_inv i_31818(.A(instrc[79]), .Z(n_28561));
	notech_inv i_31819(.A(instrc[108]), .Z(n_28562));
	notech_inv i_31820(.A(instrc[109]), .Z(n_28563));
	notech_inv i_31821(.A(n_59290), .Z(n_28564));
	notech_inv i_31822(.A(n_59263), .Z(n_28565));
	notech_inv i_31823(.A(instrc[120]), .Z(n_28566));
	notech_inv i_31824(.A(n_60516), .Z(n_28567));
	notech_inv i_31826(.A(mul64[7]), .Z(n_28569));
	notech_inv i_31827(.A(imm[14]), .Z(n_28570));
	notech_inv i_31828(.A(imm[7]), .Z(n_28571));
	notech_inv i_31829(.A(imm[30]), .Z(n_28572));
	notech_inv i_31830(.A(imm[13]), .Z(n_28573));
	notech_inv i_31831(.A(imm[12]), .Z(n_28576));
	notech_inv i_31832(.A(imm[11]), .Z(n_28577));
	notech_inv i_31833(.A(imm[10]), .Z(n_28578));
	notech_inv i_31834(.A(imm[8]), .Z(n_28579));
	notech_inv i_31835(.A(imm[38]), .Z(n_28580));
	notech_inv i_31836(.A(imm[5]), .Z(n_28581));
	notech_inv i_31837(.A(imm[37]), .Z(n_28582));
	notech_inv i_31838(.A(imm[4]), .Z(n_28583));
	notech_inv i_31839(.A(imm[36]), .Z(n_28584));
	notech_inv i_31840(.A(imm[3]), .Z(n_28585));
	notech_inv i_31841(.A(imm[35]), .Z(n_28586));
	notech_inv i_31842(.A(imm[2]), .Z(n_28587));
	notech_inv i_31843(.A(imm[0]), .Z(n_28588));
	notech_inv i_31844(.A(imm[32]), .Z(n_28589));
	notech_inv i_31845(.A(imm[1]), .Z(n_28590));
	notech_inv i_31846(.A(imm[9]), .Z(n_28591));
	notech_inv i_31847(.A(imm[16]), .Z(n_28592));
	notech_inv i_31848(.A(imm[15]), .Z(n_28593));
	notech_inv i_31849(.A(imm[47]), .Z(n_28594));
	notech_inv i_31850(.A(imm[31]), .Z(n_28595));
	notech_inv i_31851(.A(imm[17]), .Z(n_28596));
	notech_inv i_31852(.A(imm[29]), .Z(n_28598));
	notech_inv i_31853(.A(imm[28]), .Z(n_28599));
	notech_inv i_31854(.A(imm[27]), .Z(n_28600));
	notech_inv i_31855(.A(imm[26]), .Z(n_28602));
	notech_inv i_31856(.A(imm[25]), .Z(n_28603));
	notech_inv i_31857(.A(imm[24]), .Z(n_28604));
	notech_inv i_31858(.A(imm[23]), .Z(n_28605));
	notech_inv i_31859(.A(imm[22]), .Z(n_28606));
	notech_inv i_31860(.A(imm[21]), .Z(n_28607));
	notech_inv i_31861(.A(imm[20]), .Z(n_28608));
	notech_inv i_31862(.A(imm[19]), .Z(n_28609));
	notech_inv i_31863(.A(imm[18]), .Z(n_28610));
	notech_inv i_31864(.A(add_src[0]), .Z(n_28611));
	notech_inv i_31865(.A(add_src[1]), .Z(n_28612));
	notech_inv i_31866(.A(add_src[2]), .Z(n_28613));
	notech_inv i_31867(.A(add_src[3]), .Z(n_28614));
	notech_inv i_31868(.A(add_src[4]), .Z(n_28615));
	notech_inv i_31869(.A(add_src[5]), .Z(n_28616));
	notech_inv i_31870(.A(add_src[6]), .Z(n_28617));
	notech_inv i_31871(.A(add_src[7]), .Z(n_28618));
	notech_inv i_31872(.A(add_src[8]), .Z(n_28619));
	notech_inv i_31873(.A(add_src[9]), .Z(n_28620));
	notech_inv i_31875(.A(add_src[10]), .Z(n_28621));
	notech_inv i_31876(.A(add_src[11]), .Z(n_28622));
	notech_inv i_31877(.A(add_src[12]), .Z(n_28623));
	notech_inv i_31878(.A(add_src[13]), .Z(n_28624));
	notech_inv i_31879(.A(add_src[14]), .Z(n_28625));
	notech_inv i_31880(.A(add_src[15]), .Z(n_28626));
	notech_inv i_31881(.A(add_src[16]), .Z(n_28627));
	notech_inv i_31882(.A(add_src[17]), .Z(n_28628));
	notech_inv i_31883(.A(add_src[18]), .Z(n_28629));
	notech_inv i_31884(.A(add_src[19]), .Z(n_28630));
	notech_inv i_31885(.A(add_src[20]), .Z(n_28631));
	notech_inv i_31886(.A(add_src[21]), .Z(n_28632));
	notech_inv i_31887(.A(add_src[22]), .Z(n_28633));
	notech_inv i_31888(.A(add_src[23]), .Z(n_28634));
	notech_inv i_31889(.A(add_src[24]), .Z(n_28635));
	notech_inv i_31890(.A(add_src[25]), .Z(n_28636));
	notech_inv i_31891(.A(add_src[26]), .Z(n_28637));
	notech_inv i_31892(.A(add_src[27]), .Z(n_28638));
	notech_inv i_31893(.A(add_src[28]), .Z(n_28639));
	notech_inv i_31894(.A(add_src[29]), .Z(n_28640));
	notech_inv i_31895(.A(add_src[30]), .Z(n_28641));
	notech_inv i_31896(.A(add_src[31]), .Z(n_28642));
	notech_inv i_31897(.A(divq[0]), .Z(n_28643));
	notech_inv i_31898(.A(divq[1]), .Z(n_28644));
	notech_inv i_31899(.A(divq[2]), .Z(n_28645));
	notech_inv i_31900(.A(divq[3]), .Z(n_28647));
	notech_inv i_31901(.A(divq[4]), .Z(n_28648));
	notech_inv i_31902(.A(divq[5]), .Z(n_28649));
	notech_inv i_31903(.A(divq[6]), .Z(n_28650));
	notech_inv i_31904(.A(divq[7]), .Z(n_28651));
	notech_inv i_31905(.A(divq[8]), .Z(n_28652));
	notech_inv i_31906(.A(divq[9]), .Z(n_28653));
	notech_inv i_31907(.A(divq[10]), .Z(n_28654));
	notech_inv i_31908(.A(divq[11]), .Z(n_28655));
	notech_inv i_31909(.A(divq[12]), .Z(n_28656));
	notech_inv i_31910(.A(divq[13]), .Z(n_28657));
	notech_inv i_31911(.A(divq[14]), .Z(n_28658));
	notech_inv i_31912(.A(divq[15]), .Z(n_28659));
	notech_inv i_31913(.A(divq[16]), .Z(n_28660));
	notech_inv i_31914(.A(divq[17]), .Z(n_28661));
	notech_inv i_31915(.A(divq[18]), .Z(n_28662));
	notech_inv i_31916(.A(divq[19]), .Z(n_28663));
	notech_inv i_31917(.A(divq[20]), .Z(n_28664));
	notech_inv i_31918(.A(divq[21]), .Z(n_28665));
	notech_inv i_31919(.A(divq[22]), .Z(n_28666));
	notech_inv i_31920(.A(divq[23]), .Z(n_28667));
	notech_inv i_31921(.A(divq[24]), .Z(n_28668));
	notech_inv i_31922(.A(divq[25]), .Z(n_28669));
	notech_inv i_31923(.A(divq[26]), .Z(n_28670));
	notech_inv i_31924(.A(divq[27]), .Z(n_28671));
	notech_inv i_31925(.A(divq[28]), .Z(n_28672));
	notech_inv i_31926(.A(divq[29]), .Z(n_28673));
	notech_inv i_31927(.A(divq[30]), .Z(n_28674));
	notech_inv i_31928(.A(divq[31]), .Z(n_28675));
	notech_inv i_31929(.A(divq[32]), .Z(n_28676));
	notech_inv i_31930(.A(divq[33]), .Z(n_28677));
	notech_inv i_31931(.A(divq[34]), .Z(n_28678));
	notech_inv i_31932(.A(divq[35]), .Z(n_28679));
	notech_inv i_31933(.A(divq[36]), .Z(n_28680));
	notech_inv i_31934(.A(divq[37]), .Z(n_28681));
	notech_inv i_31935(.A(divq[38]), .Z(n_28682));
	notech_inv i_31936(.A(divq[39]), .Z(n_28683));
	notech_inv i_31937(.A(divq[40]), .Z(n_28684));
	notech_inv i_31938(.A(divq[41]), .Z(n_28685));
	notech_inv i_31939(.A(divq[42]), .Z(n_28686));
	notech_inv i_31940(.A(divq[43]), .Z(n_28687));
	notech_inv i_31941(.A(divq[44]), .Z(n_28688));
	notech_inv i_31942(.A(divq[45]), .Z(n_28689));
	notech_inv i_31943(.A(divq[46]), .Z(n_28690));
	notech_inv i_31944(.A(divq[47]), .Z(n_28691));
	notech_inv i_31945(.A(divq[48]), .Z(n_28692));
	notech_inv i_31946(.A(divq[49]), .Z(n_28693));
	notech_inv i_31947(.A(divq[50]), .Z(n_28694));
	notech_inv i_31948(.A(divq[51]), .Z(n_28695));
	notech_inv i_31949(.A(divq[52]), .Z(n_28696));
	notech_inv i_31950(.A(divq[53]), .Z(n_28697));
	notech_inv i_31951(.A(divq[54]), .Z(n_28698));
	notech_inv i_31953(.A(divq[55]), .Z(n_28699));
	notech_inv i_31954(.A(divq[56]), .Z(n_28700));
	notech_inv i_31955(.A(divq[57]), .Z(n_28701));
	notech_inv i_31956(.A(divq[58]), .Z(n_28702));
	notech_inv i_31957(.A(divq[59]), .Z(n_28703));
	notech_inv i_31958(.A(divq[60]), .Z(n_28704));
	notech_inv i_31959(.A(divq[61]), .Z(n_28705));
	notech_inv i_31961(.A(divq[62]), .Z(n_28706));
	notech_inv i_31962(.A(divq[63]), .Z(n_28707));
	notech_inv i_31963(.A(tsc[0]), .Z(n_28708));
	notech_inv i_31964(.A(tsc[14]), .Z(n_28709));
	notech_inv i_31965(.A(tsc[16]), .Z(n_28710));
	notech_inv i_31966(.A(tsc[17]), .Z(n_28711));
	notech_inv i_31967(.A(tsc[30]), .Z(n_28712));
	notech_inv i_31968(.A(tsc[31]), .Z(n_28713));
	notech_inv i_31969(.A(tsc[32]), .Z(n_28714));
	notech_inv i_31970(.A(tsc[34]), .Z(n_28715));
	notech_inv i_31971(.A(tsc[35]), .Z(n_28716));
	notech_inv i_31972(.A(tsc[37]), .Z(n_28717));
	notech_inv i_31973(.A(tsc[49]), .Z(n_28718));
	notech_inv i_31974(.A(tsc[51]), .Z(n_28719));
	notech_inv i_31975(.A(tsc[52]), .Z(n_28720));
	notech_inv i_31976(.A(tsc[55]), .Z(n_28721));
	notech_inv i_31977(.A(tsc[59]), .Z(n_28722));
	notech_inv i_31978(.A(nbus_144[0]), .Z(n_28723));
	notech_inv i_31979(.A(nbus_144[1]), .Z(n_28724));
	notech_inv i_31980(.A(nbus_144[2]), .Z(n_28725));
	notech_inv i_31982(.A(nbus_144[3]), .Z(n_28726));
	notech_inv i_31983(.A(nbus_144[4]), .Z(n_28727));
	notech_inv i_31984(.A(nbus_144[5]), .Z(n_28728));
	notech_inv i_31985(.A(nbus_144[7]), .Z(n_28729));
	notech_inv i_31986(.A(nbus_144[8]), .Z(n_28730));
	notech_inv i_31987(.A(nbus_143[0]), .Z(n_28731));
	notech_inv i_31988(.A(nbus_143[1]), .Z(n_28732));
	notech_inv i_31989(.A(nbus_143[2]), .Z(n_28733));
	notech_inv i_31990(.A(nbus_143[3]), .Z(n_28734));
	notech_inv i_31991(.A(nbus_143[4]), .Z(n_28735));
	notech_inv i_31992(.A(nbus_143[5]), .Z(n_28736));
	notech_inv i_31993(.A(nbus_143[6]), .Z(n_28737));
	notech_inv i_31994(.A(nbus_143[7]), .Z(n_28738));
	notech_inv i_31995(.A(nbus_143[8]), .Z(n_28739));
	notech_inv i_31996(.A(nbus_143[9]), .Z(n_28740));
	notech_inv i_31997(.A(nbus_143[10]), .Z(n_28741));
	notech_inv i_31998(.A(nbus_143[11]), .Z(n_28742));
	notech_inv i_31999(.A(nbus_143[12]), .Z(n_28743));
	notech_inv i_32000(.A(nbus_143[13]), .Z(n_28744));
	notech_inv i_32001(.A(nbus_143[14]), .Z(n_28745));
	notech_inv i_32002(.A(nbus_143[15]), .Z(n_28746));
	notech_inv i_32003(.A(nbus_143[16]), .Z(n_28747));
	notech_inv i_32004(.A(nbus_143[17]), .Z(n_28748));
	notech_inv i_32005(.A(nbus_143[18]), .Z(n_28749));
	notech_inv i_32006(.A(nbus_143[19]), .Z(n_28750));
	notech_inv i_32007(.A(nbus_143[20]), .Z(n_28751));
	notech_inv i_32008(.A(nbus_143[21]), .Z(n_28752));
	notech_inv i_32009(.A(nbus_143[22]), .Z(n_28753));
	notech_inv i_32010(.A(nbus_143[23]), .Z(n_28754));
	notech_inv i_32011(.A(nbus_143[24]), .Z(n_28755));
	notech_inv i_32012(.A(nbus_143[25]), .Z(n_28756));
	notech_inv i_32013(.A(nbus_143[26]), .Z(n_28757));
	notech_inv i_32014(.A(nbus_143[27]), .Z(n_28758));
	notech_inv i_32015(.A(nbus_143[28]), .Z(n_28763));
	notech_inv i_32016(.A(nbus_143[29]), .Z(n_28764));
	notech_inv i_32017(.A(nbus_143[30]), .Z(n_28766));
	notech_inv i_32018(.A(nbus_143[31]), .Z(n_28767));
	notech_inv i_32019(.A(nbus_143[32]), .Z(n_28768));
	notech_inv i_32020(.A(resb_shiftbox[0]), .Z(n_28769));
	notech_inv i_32021(.A(resb_shiftbox[2]), .Z(n_28770));
	notech_inv i_32022(.A(resb_shiftbox[3]), .Z(n_28775));
	notech_inv i_32023(.A(resb_shiftbox[4]), .Z(n_28778));
	notech_inv i_32024(.A(resb_shiftbox[5]), .Z(n_28779));
	notech_inv i_32025(.A(resb_shiftbox[6]), .Z(n_28780));
	notech_inv i_32026(.A(resb_shiftbox[7]), .Z(n_28781));
	notech_inv i_32027(.A(resb_shiftbox[8]), .Z(n_28782));
	notech_inv i_32028(.A(resb_shiftbox[9]), .Z(n_28783));
	notech_inv i_32029(.A(resb_shiftbox[10]), .Z(n_28784));
	notech_inv i_32030(.A(resb_shiftbox[11]), .Z(n_28785));
	notech_inv i_32031(.A(resb_shiftbox[12]), .Z(n_28786));
	notech_inv i_32032(.A(resb_shiftbox[13]), .Z(n_28787));
	notech_inv i_32033(.A(resb_shiftbox[14]), .Z(n_28788));
	notech_inv i_32034(.A(resb_shiftbox[15]), .Z(n_28789));
	notech_inv i_32035(.A(resb_shiftbox[16]), .Z(n_28790));
	notech_inv i_32036(.A(resb_shiftbox[17]), .Z(n_28791));
	notech_inv i_32037(.A(resb_shiftbox[19]), .Z(n_28792));
	notech_inv i_32038(.A(resb_shiftbox[21]), .Z(n_28793));
	notech_inv i_32039(.A(resb_shiftbox[23]), .Z(n_28794));
	notech_inv i_32040(.A(resb_shiftbox[24]), .Z(n_28795));
	notech_inv i_32041(.A(resb_shiftbox[26]), .Z(n_28796));
	notech_inv i_32042(.A(resb_shiftbox[27]), .Z(n_28797));
	notech_inv i_32043(.A(resb_shiftbox[29]), .Z(n_28798));
	notech_inv i_32044(.A(resb_shiftbox[30]), .Z(n_28799));
	notech_inv i_32046(.A(resb_shiftbox[31]), .Z(n_28800));
	notech_inv i_32047(.A(resb_shift4box[0]), .Z(n_28801));
	notech_inv i_32048(.A(resb_shift4box[1]), .Z(n_28802));
	notech_inv i_32049(.A(resb_shift4box[2]), .Z(n_28803));
	notech_inv i_32050(.A(resb_shift4box[3]), .Z(n_28804));
	notech_inv i_32051(.A(resb_shift4box[4]), .Z(n_28805));
	notech_inv i_32052(.A(resb_shift4box[5]), .Z(n_28806));
	notech_inv i_32053(.A(resb_shift4box[6]), .Z(n_28807));
	notech_inv i_32054(.A(resb_shift4box[7]), .Z(n_28808));
	notech_inv i_32055(.A(resb_shift4box[8]), .Z(n_28809));
	notech_inv i_32056(.A(resb_shift4box[9]), .Z(n_28810));
	notech_inv i_32057(.A(resb_shift4box[10]), .Z(n_28811));
	notech_inv i_32058(.A(resb_shift4box[11]), .Z(n_28812));
	notech_inv i_32059(.A(resb_shift4box[12]), .Z(n_28813));
	notech_inv i_32062(.A(resb_shift4box[13]), .Z(n_28814));
	notech_inv i_32064(.A(resb_shift4box[14]), .Z(n_28815));
	notech_inv i_32066(.A(resb_shift4box[15]), .Z(n_28816));
	notech_inv i_32067(.A(resb_shift4box[18]), .Z(n_28817));
	notech_inv i_32070(.A(resb_shift4box[19]), .Z(n_28818));
	notech_inv i_32072(.A(resb_shift4box[20]), .Z(n_28819));
	notech_inv i_32073(.A(resb_shift4box[21]), .Z(n_28821));
	notech_inv i_32074(.A(resb_shift4box[22]), .Z(n_28822));
	notech_inv i_32076(.A(resb_shift4box[23]), .Z(n_28823));
	notech_inv i_32078(.A(resb_shift4box[24]), .Z(n_28824));
	notech_inv i_32079(.A(resb_shift4box[25]), .Z(n_28825));
	notech_inv i_32080(.A(resb_shift4box[26]), .Z(n_28826));
	notech_inv i_32082(.A(resb_shift4box[27]), .Z(n_28827));
	notech_inv i_32083(.A(resb_shift4box[28]), .Z(n_28828));
	notech_inv i_32084(.A(resb_shift4box[29]), .Z(n_28829));
	notech_inv i_32085(.A(nbus_137[0]), .Z(n_28830));
	notech_inv i_32088(.A(nbus_137[1]), .Z(n_28831));
	notech_inv i_32089(.A(nbus_137[2]), .Z(n_28832));
	notech_inv i_32090(.A(nbus_137[3]), .Z(n_28833));
	notech_inv i_32091(.A(nbus_137[4]), .Z(n_28834));
	notech_inv i_32092(.A(nbus_137[5]), .Z(n_28835));
	notech_inv i_32093(.A(nbus_137[6]), .Z(n_28836));
	notech_inv i_32094(.A(nbus_137[7]), .Z(n_28837));
	notech_inv i_32095(.A(nbus_137[8]), .Z(n_28838));
	notech_inv i_32097(.A(nbus_137[9]), .Z(n_28839));
	notech_inv i_32098(.A(nbus_137[10]), .Z(n_28840));
	notech_inv i_32100(.A(nbus_137[11]), .Z(n_28841));
	notech_inv i_32103(.A(nbus_137[12]), .Z(n_28842));
	notech_inv i_32105(.A(nbus_137[13]), .Z(n_28843));
	notech_inv i_32106(.A(nbus_137[14]), .Z(n_28844));
	notech_inv i_32107(.A(nbus_137[15]), .Z(n_28845));
	notech_inv i_32108(.A(nbus_137[16]), .Z(n_28846));
	notech_inv i_32109(.A(nbus_137[17]), .Z(n_28847));
	notech_inv i_32110(.A(nbus_137[19]), .Z(n_28848));
	notech_inv i_32111(.A(nbus_137[21]), .Z(n_28849));
	notech_inv i_32112(.A(nbus_137[23]), .Z(n_28850));
	notech_inv i_32113(.A(nbus_137[26]), .Z(n_28851));
	notech_inv i_32114(.A(nbus_137[27]), .Z(n_28852));
	notech_inv i_32115(.A(nbus_137[29]), .Z(n_28853));
	notech_inv i_32116(.A(nbus_137[30]), .Z(n_28854));
	notech_inv i_32117(.A(nbus_137[31]), .Z(n_28855));
	notech_inv i_32118(.A(nbus_137[32]), .Z(n_28856));
	notech_inv i_32119(.A(nbus_11313[6]), .Z(n_28857));
	notech_inv i_32120(.A(nbus_11313[8]), .Z(n_28858));
	notech_inv i_32121(.A(nbus_11313[9]), .Z(n_28859));
	notech_inv i_32122(.A(nbus_11313[10]), .Z(n_28860));
	notech_inv i_32123(.A(nbus_11313[11]), .Z(n_28861));
	notech_inv i_32124(.A(nbus_11313[12]), .Z(n_28862));
	notech_inv i_32125(.A(nbus_11313[13]), .Z(n_28863));
	notech_inv i_32126(.A(nbus_11313[14]), .Z(n_28864));
	notech_inv i_32127(.A(nbus_11313[15]), .Z(n_28865));
	notech_inv i_32128(.A(nbus_11313[31]), .Z(n_28866));
	notech_inv i_32129(.A(from_acu[0]), .Z(n_28867));
	notech_inv i_32130(.A(from_acu[1]), .Z(n_28868));
	notech_inv i_32131(.A(from_acu[2]), .Z(n_28869));
	notech_inv i_32132(.A(from_acu[3]), .Z(n_28870));
	notech_inv i_32133(.A(from_acu[4]), .Z(n_28871));
	notech_inv i_32134(.A(from_acu[5]), .Z(n_28872));
	notech_inv i_32135(.A(from_acu[6]), .Z(n_28873));
	notech_inv i_32136(.A(write_data_33[1]), .Z(n_28875));
	notech_inv i_32137(.A(write_data_33[2]), .Z(n_28876));
	notech_inv i_32138(.A(write_data_33[3]), .Z(n_28878));
	notech_inv i_32139(.A(write_data_33[4]), .Z(n_28879));
	notech_inv i_32140(.A(write_data_33[5]), .Z(n_28880));
	notech_inv i_32141(.A(write_data_33[6]), .Z(n_28881));
	notech_inv i_32142(.A(write_data_33[7]), .Z(n_28882));
	notech_inv i_32143(.A(write_data_33[8]), .Z(n_28883));
	notech_inv i_32144(.A(write_data_33[9]), .Z(n_28884));
	notech_inv i_32145(.A(write_data_33[10]), .Z(n_28885));
	notech_inv i_32146(.A(write_data_33[11]), .Z(n_28886));
	notech_inv i_32147(.A(write_data_33[12]), .Z(n_28887));
	notech_inv i_32148(.A(write_data_33[13]), .Z(n_28888));
	notech_inv i_32149(.A(write_data_33[14]), .Z(n_28889));
	notech_inv i_32150(.A(write_data_33[15]), .Z(n_28890));
	notech_inv i_32151(.A(write_data_33[16]), .Z(n_28891));
	notech_inv i_32152(.A(write_data_33[17]), .Z(n_28892));
	notech_inv i_32153(.A(write_data_33[18]), .Z(n_28893));
	notech_inv i_32154(.A(write_data_33[19]), .Z(n_28894));
	notech_inv i_32155(.A(write_data_33[20]), .Z(n_28897));
	notech_inv i_32156(.A(write_data_33[21]), .Z(n_28898));
	notech_inv i_32157(.A(opc_14[0]), .Z(n_28901));
	notech_inv i_32158(.A(opc_14[1]), .Z(n_28902));
	notech_inv i_32159(.A(opc_14[2]), .Z(n_28903));
	notech_inv i_32160(.A(opc_14[3]), .Z(n_28904));
	notech_inv i_32161(.A(opc_14[4]), .Z(n_28905));
	notech_inv i_32162(.A(opc_14[6]), .Z(n_28906));
	notech_inv i_32163(.A(opc_14[7]), .Z(n_28907));
	notech_inv i_32164(.A(opc_14[8]), .Z(n_28908));
	notech_inv i_32165(.A(opc_14[9]), .Z(n_28909));
	notech_inv i_32166(.A(opc_14[10]), .Z(n_28910));
	notech_inv i_32167(.A(opc_14[11]), .Z(n_28911));
	notech_inv i_32168(.A(opc_14[12]), .Z(n_28912));
	notech_inv i_32169(.A(opc_14[13]), .Z(n_28913));
	notech_inv i_32170(.A(opc_14[14]), .Z(n_28914));
	notech_inv i_32171(.A(opc_14[15]), .Z(n_28915));
	notech_inv i_32172(.A(opc_14[16]), .Z(n_28916));
	notech_inv i_32173(.A(opc_14[17]), .Z(n_28917));
	notech_inv i_32174(.A(opc_14[18]), .Z(n_28918));
	notech_inv i_32175(.A(opc_14[19]), .Z(n_28919));
	notech_inv i_32176(.A(opc_14[20]), .Z(n_28920));
	notech_inv i_32177(.A(opc_14[21]), .Z(n_28921));
	notech_inv i_32178(.A(opc_14[22]), .Z(n_28922));
	notech_inv i_32179(.A(opc_14[23]), .Z(n_28923));
	notech_inv i_32180(.A(opc_14[24]), .Z(n_28924));
	notech_inv i_32181(.A(opc_14[25]), .Z(n_28925));
	notech_inv i_32182(.A(opc_14[26]), .Z(n_28926));
	notech_inv i_32183(.A(opc_14[27]), .Z(n_28927));
	notech_inv i_32184(.A(opc_14[28]), .Z(n_28928));
	notech_inv i_32185(.A(opc_14[29]), .Z(n_28929));
	notech_inv i_32186(.A(opc_14[30]), .Z(n_28930));
	notech_inv i_32187(.A(opc_14[31]), .Z(n_28931));
	notech_inv i_32188(.A(n_1069), .Z(n_28932));
	notech_inv i_32189(.A(divr[0]), .Z(nbus_11348[0]));
	notech_inv i_32190(.A(divr[1]), .Z(nbus_11348[1]));
	notech_inv i_32191(.A(divr[2]), .Z(nbus_11348[2]));
	notech_inv i_32192(.A(divr[3]), .Z(nbus_11348[3]));
	notech_inv i_32193(.A(divr[4]), .Z(nbus_11348[4]));
	notech_inv i_32194(.A(divr[5]), .Z(nbus_11348[5]));
	notech_inv i_32195(.A(divr[6]), .Z(nbus_11348[6]));
	notech_inv i_32196(.A(divr[7]), .Z(nbus_11348[7]));
	notech_inv i_32197(.A(divr[8]), .Z(nbus_11348[8]));
	notech_inv i_32198(.A(divr[9]), .Z(nbus_11348[9]));
	notech_inv i_32199(.A(divr[10]), .Z(nbus_11348[10]));
	notech_inv i_32200(.A(divr[11]), .Z(nbus_11348[11]));
	notech_inv i_32201(.A(divr[12]), .Z(nbus_11348[12]));
	notech_inv i_32202(.A(divr[13]), .Z(nbus_11348[13]));
	notech_inv i_32203(.A(divr[14]), .Z(nbus_11348[14]));
	notech_inv i_32204(.A(divr[15]), .Z(nbus_11348[15]));
	notech_inv i_32205(.A(divr[16]), .Z(nbus_11348[16]));
	notech_inv i_3220695047(.A(divr[17]), .Z(nbus_11348[17]));
	notech_inv i_32207(.A(divr[18]), .Z(nbus_11348[18]));
	notech_inv i_32208(.A(divr[19]), .Z(nbus_11348[19]));
	notech_inv i_32209(.A(divr[20]), .Z(nbus_11348[20]));
	notech_inv i_32210(.A(divr[21]), .Z(nbus_11348[21]));
	notech_inv i_3221195046(.A(divr[22]), .Z(nbus_11348[22]));
	notech_inv i_32212(.A(divr[23]), .Z(nbus_11348[23]));
	notech_inv i_32213(.A(divr[24]), .Z(nbus_11348[24]));
	notech_inv i_32214(.A(divr[25]), .Z(nbus_11348[25]));
	notech_inv i_32215(.A(divr[26]), .Z(nbus_11348[26]));
	notech_inv i_3221695045(.A(divr[27]), .Z(nbus_11348[27]));
	notech_inv i_32217(.A(divr[28]), .Z(nbus_11348[28]));
	notech_inv i_32218(.A(divr[29]), .Z(nbus_11348[29]));
	notech_inv i_32219(.A(divr[30]), .Z(nbus_11348[30]));
	notech_inv i_32220(.A(divr[31]), .Z(nbus_11348[31]));
	notech_inv i_3222195044(.A(n_56460), .Z(n_28966));
	notech_inv i_32222(.A(n_56478), .Z(n_28967));
	notech_inv i_32223(.A(readio_ack), .Z(n_28968));
	notech_inv i_32224(.A(n_62437), .Z(n_28969));
	notech_inv i_32225(.A(instrc[126]), .Z(n_28970));
	notech_inv i_3222695043(.A(instrc[102]), .Z(n_28971));
	notech_inv i_32227(.A(instrc[94]), .Z(n_28972));
	notech_inv i_32228(.A(instrc[86]), .Z(n_28973));
	notech_inv i_32229(.A(n_62395), .Z(n_28974));
	notech_inv i_32230(.A(\opcode[3] ), .Z(n_28975));
	notech_inv i_3223195042(.A(n_62433), .Z(n_28976));
	notech_inv i_32232(.A(\regs_13_14[29] ), .Z(n_28977));
	notech_inv i_32233(.A(\nbus_14524[17] ), .Z(n_28978));
	notech_inv i_32234(.A(\eflags[17] ), .Z(n_28979));
	notech_inv i_32235(.A(\nbus_14524[7] ), .Z(n_28980));
	notech_inv i_32236(.A(\eflags[7] ), .Z(n_28981));
	notech_inv i_32237(.A(n_6801), .Z(n_28982));
	notech_inv i_32238(.A(\opa_12[7] ), .Z(n_28983));
	notech_inv i_32239(.A(n_60584), .Z(n_28984));
	notech_inv i_32240(.A(\eflags[0] ), .Z(n_28985));
	notech_inv i_32241(.A(\opa_12[0] ), .Z(n_28986));
	notech_inv i_32242(.A(\regs_13_14[17] ), .Z(n_28987));
	notech_inv i_32243(.A(\eflags[30] ), .Z(n_28988));
	notech_inv i_32244(.A(\nbus_14524[30] ), .Z(n_28989));
	notech_inv i_32245(.A(\eflags[31] ), .Z(n_28990));
	notech_inv i_32246(.A(\nbus_14524[31] ), .Z(n_28991));
	notech_inv i_32247(.A(\nbus_14524[29] ), .Z(n_28992));
	notech_inv i_32248(.A(\eflags[29] ), .Z(n_28993));
	notech_inv i_32249(.A(n_3409), .Z(n_28994));
	notech_inv i_32250(.A(n_3408), .Z(n_28995));
	notech_inv i_32251(.A(\regs_13_14[31] ), .Z(n_28996));
	notech_inv i_32252(.A(\regs_13_14[30] ), .Z(n_28997));
	notech_inv i_32253(.A(n_3407), .Z(n_28998));
	notech_inv i_32254(.A(n_3406), .Z(n_28999));
	notech_inv i_32255(.A(\eflags[14] ), .Z(n_29000));
	notech_inv i_32256(.A(\nbus_14524[14] ), .Z(n_29001));
	notech_inv i_32257(.A(\eflags[16] ), .Z(n_29002));
	notech_inv i_32258(.A(\nbus_14524[16] ), .Z(n_29003));
	notech_inv i_32259(.A(\regs_13_14[16] ), .Z(n_29004));
	notech_inv i_32260(.A(n_6810), .Z(n_29005));
	notech_inv i_32261(.A(\opa_12[14] ), .Z(n_29006));
	notech_inv i_32263(.A(n_4689), .Z(n_29007));
	notech_inv i_32264(.A(n_57162), .Z(n_29008));
	notech_inv i_32265(.A(start_up), .Z(n_29009));
	notech_inv i_32266(.A(n_56469), .Z(n_29010));
	notech_inv i_32267(.A(n_1046), .Z(n_29011));
	notech_inv i_32268(.A(n_1011), .Z(n_29012));
	notech_inv i_32270(.A(instrc[98]), .Z(n_29013));
	notech_inv i_32271(.A(instrc[90]), .Z(n_29014));
	notech_inv i_32272(.A(instrc[82]), .Z(n_29015));
	notech_inv i_32274(.A(instrc[99]), .Z(n_29016));
	notech_inv i_32275(.A(instrc[91]), .Z(n_29017));
	notech_inv i_32276(.A(instrc[83]), .Z(n_29018));
	notech_inv i_32277(.A(instrc[96]), .Z(n_29019));
	notech_inv i_32279(.A(instrc[88]), .Z(n_29020));
	notech_inv i_32280(.A(instrc[80]), .Z(n_29021));
	notech_inv i_32281(.A(instrc[97]), .Z(n_29022));
	notech_inv i_32283(.A(instrc[89]), .Z(n_29023));
	notech_inv i_32284(.A(instrc[81]), .Z(n_29024));
	notech_inv i_32285(.A(instrc[101]), .Z(n_29025));
	notech_inv i_32286(.A(instrc[93]), .Z(n_29026));
	notech_inv i_32287(.A(instrc[85]), .Z(n_29027));
	notech_inv i_32289(.A(instrc[127]), .Z(n_29028));
	notech_inv i_32290(.A(instrc[103]), .Z(n_29029));
	notech_inv i_32291(.A(instrc[95]), .Z(n_29030));
	notech_inv i_32292(.A(instrc[87]), .Z(n_29031));
	notech_inv i_32293(.A(instrc[124]), .Z(n_29032));
	notech_inv i_32294(.A(instrc[100]), .Z(n_29033));
	notech_inv i_32295(.A(instrc[92]), .Z(n_29034));
	notech_inv i_32296(.A(instrc[84]), .Z(n_29035));
	notech_inv i_32297(.A(n_6296), .Z(n_29036));
	notech_inv i_32298(.A(\opa_12[13] ), .Z(n_29037));
	notech_inv i_32299(.A(\opa_1[13] ), .Z(n_29038));
	notech_inv i_32300(.A(mul64[13]), .Z(n_29039));
	notech_inv i_32301(.A(instrc[107]), .Z(n_29040));
	notech_inv i_32302(.A(n_4678), .Z(n_29041));
	notech_inv i_32303(.A(\opa_12[3] ), .Z(n_29043));
	notech_inv i_32304(.A(n_4683), .Z(n_29044));
	notech_inv i_32305(.A(\opa_12[8] ), .Z(n_29045));
	notech_inv i_32306(.A(n_4684), .Z(n_29046));
	notech_inv i_32307(.A(\regs_1[9] ), .Z(n_29047));
	notech_inv i_32309(.A(\opa_12[9] ), .Z(n_29048));
	notech_inv i_32310(.A(\opa_12[1] ), .Z(n_29049));
	notech_inv i_32311(.A(\opa_12[2] ), .Z(n_29050));
	notech_inv i_32312(.A(n_5169), .Z(n_29051));
	notech_inv i_32313(.A(n_4676), .Z(n_29053));
	notech_inv i_32314(.A(n_4677), .Z(n_29056));
	notech_inv i_32315(.A(n_4679), .Z(n_29058));
	notech_inv i_32316(.A(\regs_1[4] ), .Z(n_29059));
	notech_inv i_32317(.A(\opa_12[4] ), .Z(n_29063));
	notech_inv i_32318(.A(n_4680), .Z(n_29064));
	notech_inv i_32319(.A(\opa_12[5] ), .Z(n_29065));
	notech_inv i_32320(.A(n_4681), .Z(n_29066));
	notech_inv i_32322(.A(\opa_12[6] ), .Z(n_29068));
	notech_inv i_32323(.A(\regs_1[7] ), .Z(n_29076));
	notech_inv i_32324(.A(\opa_12[10] ), .Z(n_29077));
	notech_inv i_32325(.A(n_4685), .Z(n_29078));
	notech_inv i_32326(.A(\regs_1[10] ), .Z(n_29079));
	notech_inv i_32327(.A(\opa_12[11] ), .Z(n_29080));
	notech_inv i_32328(.A(n_4686), .Z(n_29081));
	notech_inv i_32329(.A(n_4687), .Z(n_29082));
	notech_inv i_32330(.A(\regs_1[12] ), .Z(n_29083));
	notech_inv i_32331(.A(\opa_12[12] ), .Z(n_29084));
	notech_inv i_32332(.A(n_4688), .Z(n_29085));
	notech_inv i_32333(.A(\regs_1[13] ), .Z(n_29086));
	notech_inv i_32334(.A(\opa_12[15] ), .Z(n_29087));
	notech_inv i_32335(.A(n_4690), .Z(n_29088));
	notech_inv i_32336(.A(\add_len_pc[10] ), .Z(n_29089));
	notech_inv i_32337(.A(\nbus_14524[10] ), .Z(n_29090));
	notech_inv i_32338(.A(n_55460), .Z(n_29091));
	notech_inv i_32339(.A(\add_len_pc[11] ), .Z(n_29092));
	notech_inv i_32340(.A(\nbus_14524[11] ), .Z(n_29093));
	notech_inv i_32341(.A(\eflags[11] ), .Z(n_29094));
	notech_inv i_32342(.A(\add_len_pc[12] ), .Z(n_29095));
	notech_inv i_32343(.A(\nbus_14524[12] ), .Z(n_29096));
	notech_inv i_32344(.A(\eflags[12] ), .Z(n_29097));
	notech_inv i_32345(.A(\add_len_pc[13] ), .Z(n_29098));
	notech_inv i_32346(.A(\nbus_14524[13] ), .Z(n_29099));
	notech_inv i_32347(.A(\eflags[13] ), .Z(n_29100));
	notech_inv i_32348(.A(\nbus_14524[8] ), .Z(n_29101));
	notech_inv i_32349(.A(\eflags[8] ), .Z(n_29102));
	notech_inv i_32350(.A(\nbus_14524[4] ), .Z(n_29103));
	notech_inv i_32351(.A(\eflags[4] ), .Z(n_29104));
	notech_inv i_32352(.A(\nbus_14524[6] ), .Z(n_29105));
	notech_inv i_32353(.A(\eflags[6] ), .Z(n_29106));
	notech_inv i_32354(.A(n_6800), .Z(n_29107));
	notech_inv i_32355(.A(n_6798), .Z(n_29108));
	notech_inv i_32356(.A(n_2414), .Z(n_29109));
	notech_inv i_32357(.A(n_2415), .Z(n_29110));
	notech_inv i_32358(.A(n_3346), .Z(n_29111));
	notech_inv i_32359(.A(\regs_1_0[17] ), .Z(n_29112));
	notech_inv i_32360(.A(mul64[17]), .Z(n_29113));
	notech_inv i_32361(.A(n_4693), .Z(n_29114));
	notech_inv i_32362(.A(\nbus_14524[2] ), .Z(n_29115));
	notech_inv i_32363(.A(\eflags[3] ), .Z(n_29116));
	notech_inv i_32364(.A(\nbus_14524[3] ), .Z(n_29117));
	notech_inv i_32365(.A(\eflags[5] ), .Z(n_29118));
	notech_inv i_32366(.A(\nbus_14524[5] ), .Z(n_29119));
	notech_inv i_32367(.A(instrc[104]), .Z(n_29120));
	notech_inv i_32368(.A(\eflags[2] ), .Z(n_29121));
	notech_inv i_32369(.A(instrc[105]), .Z(n_29122));
	notech_inv i_32370(.A(n_61131), .Z(n_29123));
	notech_inv i_32371(.A(n_613), .Z(n_29124));
	notech_inv i_32372(.A(n_6697), .Z(n_29125));
	notech_inv i_32373(.A(n_6646), .Z(n_29126));
	notech_inv i_32374(.A(n_6621), .Z(n_29127));
	notech_inv i_32375(.A(n_6588), .Z(n_29128));
	notech_inv i_32376(.A(n_6541), .Z(n_29129));
	notech_inv i_32377(.A(read_ack), .Z(n_29130));
	notech_inv i_32378(.A(n_2449), .Z(n_29131));
	notech_inv i_32379(.A(n_2448), .Z(n_29132));
	notech_inv i_32380(.A(n_2427), .Z(n_29133));
	notech_inv i_32381(.A(n_2429), .Z(n_29134));
	notech_inv i_32382(.A(n_2432), .Z(n_29135));
	notech_inv i_32383(.A(n_2433), .Z(n_29136));
	notech_inv i_32384(.A(\regs_13_14[24] ), .Z(n_29137));
	notech_inv i_32385(.A(n_2435), .Z(n_29138));
	notech_inv i_32386(.A(n_2437), .Z(n_29139));
	notech_inv i_32387(.A(n_2441), .Z(n_29140));
	notech_inv i_32388(.A(n_2463), .Z(n_29141));
	notech_inv i_32389(.A(\nbus_14524[24] ), .Z(n_29142));
	notech_inv i_32390(.A(\eflags[24] ), .Z(n_29143));
	notech_inv i_32391(.A(n_2476), .Z(n_29144));
	notech_inv i_32392(.A(n_2477), .Z(n_29145));
	notech_inv i_32393(.A(n_2474), .Z(n_29146));
	notech_inv i_32394(.A(n_2475), .Z(n_29147));
	notech_inv i_32395(.A(n_2472), .Z(n_29148));
	notech_inv i_32396(.A(n_2473), .Z(n_29149));
	notech_inv i_32397(.A(n_3445), .Z(n_29150));
	notech_inv i_32398(.A(n_2461), .Z(n_29151));
	notech_inv i_32399(.A(\regs_13_14[23] ), .Z(n_29152));
	notech_inv i_32400(.A(n_2469), .Z(n_29153));
	notech_inv i_32401(.A(\regs_13_14[27] ), .Z(n_29154));
	notech_inv i_32402(.A(n_6820), .Z(n_29155));
	notech_inv i_32403(.A(\regs_13_14[26] ), .Z(n_29156));
	notech_inv i_32404(.A(\add_len_pc[26] ), .Z(n_29157));
	notech_inv i_32405(.A(\nbus_14524[26] ), .Z(n_29158));
	notech_inv i_32406(.A(\eflags[26] ), .Z(n_29159));
	notech_inv i_32407(.A(n_6821), .Z(n_29160));
	notech_inv i_32408(.A(\add_len_pc[27] ), .Z(n_29161));
	notech_inv i_32409(.A(\eflags[27] ), .Z(n_29162));
	notech_inv i_32410(.A(\nbus_14524[27] ), .Z(n_29163));
	notech_inv i_32411(.A(n_2451), .Z(n_29164));
	notech_inv i_32412(.A(\regs_13_14[18] ), .Z(n_29165));
	notech_inv i_32413(.A(n_2453), .Z(n_29166));
	notech_inv i_32414(.A(\regs_13_14[19] ), .Z(n_29167));
	notech_inv i_32415(.A(n_2455), .Z(n_29168));
	notech_inv i_32416(.A(\regs_13_14[20] ), .Z(n_29169));
	notech_inv i_32417(.A(n_2457), .Z(n_29170));
	notech_inv i_32418(.A(\regs_13_14[21] ), .Z(n_29172));
	notech_inv i_32419(.A(n_2459), .Z(n_29173));
	notech_inv i_32420(.A(\regs_13_14[22] ), .Z(n_29174));
	notech_inv i_32421(.A(n_6814), .Z(n_29175));
	notech_inv i_32422(.A(\add_len_pc[20] ), .Z(n_29176));
	notech_inv i_32423(.A(\nbus_14524[20] ), .Z(n_29177));
	notech_inv i_32424(.A(\eflags[20] ), .Z(n_29178));
	notech_inv i_32425(.A(n_6815), .Z(n_29179));
	notech_inv i_32426(.A(\add_len_pc[21] ), .Z(n_29180));
	notech_inv i_32427(.A(\nbus_14524[21] ), .Z(n_29181));
	notech_inv i_32428(.A(\eflags[21] ), .Z(n_29182));
	notech_inv i_32429(.A(n_2446), .Z(n_29183));
	notech_inv i_32430(.A(n_2447), .Z(n_29184));
	notech_inv i_32431(.A(n_2442), .Z(n_29185));
	notech_inv i_32432(.A(n_2443), .Z(n_29186));
	notech_inv i_32433(.A(n_614), .Z(n_29187));
	notech_inv i_32434(.A(n_3416), .Z(n_29188));
	notech_inv i_32435(.A(n_3419), .Z(n_29189));
	notech_inv i_32436(.A(\regs_1_0[29] ), .Z(n_29190));
	notech_inv i_32437(.A(n_3415), .Z(n_29191));
	notech_inv i_32438(.A(n_3417), .Z(n_29194));
	notech_inv i_32439(.A(n_3418), .Z(n_29195));
	notech_inv i_32440(.A(n_3420), .Z(n_29198));
	notech_inv i_32441(.A(n_3421), .Z(n_29199));
	notech_inv i_32442(.A(n_3356), .Z(n_29200));
	notech_inv i_32443(.A(n_3357), .Z(n_29201));
	notech_inv i_32444(.A(n_2425), .Z(n_29202));
	notech_inv i_32445(.A(n_3426), .Z(n_29203));
	notech_inv i_32446(.A(n_3429), .Z(n_29204));
	notech_inv i_32447(.A(\nbus_14524[15] ), .Z(n_29205));
	notech_inv i_32448(.A(\eflags[15] ), .Z(n_29206));
	notech_inv i_32449(.A(n_6799), .Z(n_29207));
	notech_inv i_32450(.A(n_3414), .Z(n_29208));
	notech_inv i_32451(.A(n_6825), .Z(n_29209));
	notech_inv i_32452(.A(n_6824), .Z(n_29210));
	notech_inv i_32453(.A(n_6823), .Z(n_29211));
	notech_inv i_32454(.A(n_3444), .Z(n_29212));
	notech_inv i_32455(.A(\regs_1_0[31] ), .Z(n_29213));
	notech_inv i_32456(.A(\regs_1_0[25] ), .Z(n_29214));
	notech_inv i_32457(.A(\regs_13_14[25] ), .Z(n_29215));
	notech_inv i_32458(.A(\regs_1_0[26] ), .Z(n_29216));
	notech_inv i_32459(.A(\regs_1_0[27] ), .Z(n_29217));
	notech_inv i_32460(.A(\regs_1_0[28] ), .Z(n_29218));
	notech_inv i_32461(.A(\regs_13_14[28] ), .Z(n_29219));
	notech_inv i_32462(.A(n_6817), .Z(n_29220));
	notech_inv i_32463(.A(\add_len_pc[23] ), .Z(n_29221));
	notech_inv i_32464(.A(\nbus_14524[23] ), .Z(n_29222));
	notech_inv i_32465(.A(\eflags[23] ), .Z(n_29223));
	notech_inv i_32466(.A(n_6819), .Z(n_29224));
	notech_inv i_32467(.A(\add_len_pc[25] ), .Z(n_29225));
	notech_inv i_32468(.A(\nbus_14524[25] ), .Z(n_29226));
	notech_inv i_32469(.A(\eflags[25] ), .Z(n_29227));
	notech_inv i_32470(.A(\eflags[28] ), .Z(n_29228));
	notech_inv i_32471(.A(\nbus_14524[28] ), .Z(n_29229));
	notech_inv i_32472(.A(\regs_1_0[18] ), .Z(n_29230));
	notech_inv i_32473(.A(n_6812), .Z(n_29231));
	notech_inv i_32474(.A(\add_len_pc[18] ), .Z(n_29232));
	notech_inv i_32475(.A(\nbus_14524[18] ), .Z(n_29233));
	notech_inv i_32476(.A(\eflags[18] ), .Z(n_29234));
	notech_inv i_32477(.A(n_6813), .Z(n_29235));
	notech_inv i_32478(.A(\add_len_pc[19] ), .Z(n_29236));
	notech_inv i_32479(.A(\nbus_14524[19] ), .Z(n_29237));
	notech_inv i_32480(.A(\eflags[19] ), .Z(n_29238));
	notech_inv i_32481(.A(n_6816), .Z(n_29239));
	notech_inv i_32482(.A(\add_len_pc[22] ), .Z(n_29240));
	notech_inv i_32483(.A(\eflags[22] ), .Z(n_29241));
	notech_inv i_32484(.A(\nbus_14524[22] ), .Z(n_29242));
	notech_inv i_32486(.A(n_3430), .Z(n_29243));
	notech_inv i_32487(.A(n_3428), .Z(n_29244));
	notech_inv i_32488(.A(\regs_1_0[16] ), .Z(n_29245));
	notech_inv i_32489(.A(\add_len_pc[28] ), .Z(n_29246));
	notech_inv i_32490(.A(n_2421), .Z(n_29247));
	notech_inv i_32491(.A(n_3348), .Z(n_29248));
	notech_inv i_32492(.A(n_3349), .Z(n_29249));
	notech_inv i_32493(.A(n_3350), .Z(n_29250));
	notech_inv i_32494(.A(n_3351), .Z(n_29251));
	notech_inv i_32495(.A(n_3353), .Z(n_29252));
	notech_inv i_32496(.A(n_3352), .Z(n_29253));
	notech_inv i_32497(.A(n_3364), .Z(n_29254));
	notech_inv i_32498(.A(n_3365), .Z(n_29255));
	notech_inv i_32499(.A(n_2417), .Z(n_29256));
	notech_inv i_32500(.A(n_2419), .Z(n_29257));
	notech_inv i_32501(.A(n_3362), .Z(n_29258));
	notech_inv i_32502(.A(n_3366), .Z(n_29259));
	notech_inv i_32503(.A(n_3368), .Z(n_29260));
	notech_inv i_32504(.A(n_3370), .Z(n_29261));
	notech_inv i_32505(.A(n_3372), .Z(n_29262));
	notech_inv i_32506(.A(n_3376), .Z(n_29263));
	notech_inv i_32507(.A(\nbus_14524[9] ), .Z(n_29264));
	notech_inv i_32508(.A(ie), .Z(n_29265));
	notech_inv i_32509(.A(\eflags[1] ), .Z(n_29266));
	notech_inv i_32510(.A(n_6811), .Z(n_29267));
	notech_inv i_32511(.A(n_6803), .Z(n_29268));
	notech_inv i_32512(.A(n_353169303), .Z(n_29269));
	notech_inv i_32513(.A(n_6797), .Z(n_29270));
	notech_inv i_32514(.A(n_6796), .Z(n_29271));
	notech_inv i_32515(.A(n_6795), .Z(n_29272));
	notech_inv i_32516(.A(n_6794), .Z(n_29273));
	notech_inv i_32517(.A(n_3443), .Z(n_29274));
	notech_inv i_32518(.A(mul64[29]), .Z(n_29275));
	notech_inv i_32519(.A(n_4705), .Z(n_29276));
	notech_inv i_32520(.A(mul64[45]), .Z(n_29277));
	notech_inv i_32521(.A(\opc_5[13] ), .Z(n_29278));
	notech_inv i_32522(.A(n_3381), .Z(n_29279));
	notech_inv i_32523(.A(n_3380), .Z(n_29280));
	notech_inv i_32524(.A(n_3379), .Z(n_29281));
	notech_inv i_32525(.A(n_3378), .Z(n_29282));
	notech_inv i_32526(.A(n_3375), .Z(n_29283));
	notech_inv i_32527(.A(n_3374), .Z(n_29284));
	notech_inv i_32528(.A(n_5880), .Z(n_29285));
	notech_inv i_32529(.A(n_5881), .Z(n_29286));
	notech_inv i_32530(.A(n_5882), .Z(n_29287));
	notech_inv i_32531(.A(nCF_shiftbox), .Z(n_29288));
	notech_inv i_32532(.A(n_6283), .Z(n_29289));
	notech_inv i_32533(.A(n_6284), .Z(n_29290));
	notech_inv i_32534(.A(n_6285), .Z(n_29291));
	notech_inv i_32535(.A(n_6286), .Z(n_29292));
	notech_inv i_32536(.A(n_6287), .Z(n_29293));
	notech_inv i_32537(.A(n_6288), .Z(n_29294));
	notech_inv i_32538(.A(n_6289), .Z(n_29295));
	notech_inv i_32539(.A(\opa_1[7] ), .Z(n_29296));
	notech_inv i_32540(.A(n_6290), .Z(n_29297));
	notech_inv i_32541(.A(\opa_1[8] ), .Z(n_29298));
	notech_inv i_32542(.A(mul64[8]), .Z(n_29299));
	notech_inv i_32543(.A(n_6291), .Z(n_29300));
	notech_inv i_32544(.A(\opa_1[9] ), .Z(n_29301));
	notech_inv i_32545(.A(mul64[9]), .Z(n_29302));
	notech_inv i_32546(.A(n_6292), .Z(n_29303));
	notech_inv i_32547(.A(\opa_1[10] ), .Z(n_29304));
	notech_inv i_32548(.A(mul64[10]), .Z(n_29305));
	notech_inv i_32549(.A(n_6293), .Z(n_29306));
	notech_inv i_32550(.A(\opa_1[11] ), .Z(n_29307));
	notech_inv i_32551(.A(mul64[11]), .Z(n_29308));
	notech_inv i_32552(.A(n_6294), .Z(n_29309));
	notech_inv i_32553(.A(\opa_1[12] ), .Z(n_29310));
	notech_inv i_32554(.A(mul64[12]), .Z(n_29311));
	notech_inv i_32555(.A(n_6295), .Z(n_29312));
	notech_inv i_32556(.A(\opa_1[14] ), .Z(n_29313));
	notech_inv i_32557(.A(mul64[14]), .Z(n_29314));
	notech_inv i_32558(.A(n_6297), .Z(n_29315));
	notech_inv i_32559(.A(\opa_1[15] ), .Z(n_29316));
	notech_inv i_32560(.A(mul64[15]), .Z(n_29317));
	notech_inv i_32561(.A(n_6298), .Z(n_29318));
	notech_inv i_32562(.A(n_6299), .Z(n_29319));
	notech_inv i_32563(.A(mul64[16]), .Z(n_29320));
	notech_inv i_32564(.A(n_6300), .Z(n_29321));
	notech_inv i_32565(.A(n_6301), .Z(n_29322));
	notech_inv i_32566(.A(mul64[18]), .Z(n_29323));
	notech_inv i_32567(.A(n_6302), .Z(n_29324));
	notech_inv i_32568(.A(mul64[19]), .Z(n_29325));
	notech_inv i_32569(.A(n_6303), .Z(n_29326));
	notech_inv i_32570(.A(mul64[20]), .Z(n_29327));
	notech_inv i_32571(.A(n_6304), .Z(n_29328));
	notech_inv i_32572(.A(mul64[21]), .Z(n_29329));
	notech_inv i_32573(.A(n_6305), .Z(n_29330));
	notech_inv i_32574(.A(mul64[22]), .Z(n_29331));
	notech_inv i_32575(.A(n_6306), .Z(n_29332));
	notech_inv i_32576(.A(mul64[23]), .Z(n_29333));
	notech_inv i_32577(.A(n_6307), .Z(n_29334));
	notech_inv i_32578(.A(mul64[24]), .Z(n_29335));
	notech_inv i_32579(.A(n_6308), .Z(n_29336));
	notech_inv i_32580(.A(mul64[25]), .Z(n_29337));
	notech_inv i_32581(.A(n_6309), .Z(n_29338));
	notech_inv i_32582(.A(mul64[26]), .Z(n_29339));
	notech_inv i_32583(.A(n_6310), .Z(n_29340));
	notech_inv i_32584(.A(mul64[27]), .Z(n_29341));
	notech_inv i_32585(.A(n_6311), .Z(n_29342));
	notech_inv i_32586(.A(mul64[28]), .Z(n_29343));
	notech_inv i_32587(.A(n_6312), .Z(n_29344));
	notech_inv i_32588(.A(n_6313), .Z(n_29345));
	notech_inv i_32589(.A(mul64[30]), .Z(n_29346));
	notech_inv i_32590(.A(n_6314), .Z(n_29347));
	notech_inv i_32591(.A(mul64[31]), .Z(n_29348));
	notech_inv i_32592(.A(n_3360), .Z(n_29349));
	notech_inv i_32593(.A(n_3361), .Z(n_29350));
	notech_inv i_32594(.A(n_2423), .Z(n_29351));
	notech_inv i_32595(.A(n_3424), .Z(n_29352));
	notech_inv i_32596(.A(n_2431), .Z(n_29354));
	notech_inv i_32597(.A(n_2439), .Z(n_29355));
	notech_inv i_32598(.A(n_2445), .Z(n_29356));
	notech_inv i_32599(.A(n_4718), .Z(n_29357));
	notech_inv i_32600(.A(mul64[58]), .Z(n_29358));
	notech_inv i_32601(.A(\opc_5[26] ), .Z(n_29359));
	notech_inv i_32602(.A(n_4716), .Z(n_29360));
	notech_inv i_32603(.A(mul64[56]), .Z(n_29361));
	notech_inv i_32604(.A(\opc_5[24] ), .Z(n_29362));
	notech_inv i_32605(.A(n_4702), .Z(n_29363));
	notech_inv i_32606(.A(mul64[42]), .Z(n_29364));
	notech_inv i_32607(.A(n_4700), .Z(n_29367));
	notech_inv i_32608(.A(mul64[40]), .Z(n_29368));
	notech_inv i_32609(.A(n_4695), .Z(n_29369));
	notech_inv i_32610(.A(n_4694), .Z(n_29370));
	notech_inv i_32611(.A(n_4692), .Z(n_29371));
	notech_inv i_32612(.A(n_2465), .Z(n_29372));
	notech_inv i_32613(.A(n_2467), .Z(n_29373));
	notech_inv i_32614(.A(n_2471), .Z(n_29374));
	notech_inv i_32615(.A(n_6808), .Z(n_29375));
	notech_inv i_32616(.A(write_ack), .Z(n_29376));
	notech_inv i_32617(.A(n_3423), .Z(n_29377));
	notech_inv i_32618(.A(n_3431), .Z(n_29378));
	notech_inv i_32619(.A(n_3358), .Z(n_29379));
	notech_inv i_32620(.A(n_3359), .Z(n_29380));
	notech_inv i_32621(.A(n_3405), .Z(n_29381));
	notech_inv i_32622(.A(n_6351), .Z(n_29382));
	notech_inv i_32623(.A(n_6352), .Z(n_29383));
	notech_inv i_32625(.A(n_6353), .Z(n_29384));
	notech_inv i_32626(.A(n_6354), .Z(n_29385));
	notech_inv i_32627(.A(n_5156), .Z(n_29386));
	notech_inv i_32628(.A(n_6357), .Z(n_29387));
	notech_inv i_32629(.A(n_6358), .Z(n_29388));
	notech_inv i_32630(.A(n_5158), .Z(n_29389));
	notech_inv i_32631(.A(n_5159), .Z(n_29390));
	notech_inv i_32632(.A(n_5160), .Z(n_29391));
	notech_inv i_32633(.A(n_6365), .Z(n_29392));
	notech_inv i_32634(.A(n_6366), .Z(n_29393));
	notech_inv i_32635(.A(n_5162), .Z(n_29394));
	notech_inv i_32636(.A(n_6368), .Z(n_29395));
	notech_inv i_32637(.A(n_5163), .Z(n_29396));
	notech_inv i_32638(.A(n_5164), .Z(n_29397));
	notech_inv i_32639(.A(n_5165), .Z(n_29398));
	notech_inv i_32640(.A(n_5166), .Z(n_29399));
	notech_inv i_32641(.A(n_5167), .Z(n_29400));
	notech_inv i_32642(.A(n_5168), .Z(n_29401));
	notech_inv i_32643(.A(n_5170), .Z(n_29402));
	notech_inv i_32644(.A(n_5171), .Z(n_29403));
	notech_inv i_32645(.A(n_5172), .Z(n_29404));
	notech_inv i_32646(.A(n_5173), .Z(n_29405));
	notech_inv i_32647(.A(n_5174), .Z(n_29406));
	notech_inv i_32648(.A(n_5175), .Z(n_29407));
	notech_inv i_32649(.A(n_5176), .Z(n_29408));
	notech_inv i_32650(.A(n_5177), .Z(n_29409));
	notech_inv i_32651(.A(n_5178), .Z(n_29410));
	notech_inv i_32652(.A(n_5179), .Z(n_29411));
	notech_inv i_32653(.A(n_5180), .Z(n_29412));
	notech_inv i_32654(.A(n_5181), .Z(n_29413));
	notech_inv i_32655(.A(n_5182), .Z(n_29414));
	notech_inv i_32656(.A(n_5183), .Z(n_29415));
	notech_inv i_32657(.A(\regs_1_0[24] ), .Z(n_29416));
	notech_inv i_32658(.A(n_3422), .Z(n_29417));
	notech_inv i_32659(.A(n_3425), .Z(n_29418));
	notech_inv i_32660(.A(n_3427), .Z(n_29419));
	notech_inv i_32661(.A(n_3438), .Z(n_29420));
	notech_inv i_32662(.A(n_3394), .Z(n_29421));
	notech_inv i_32663(.A(\opc_1[4] ), .Z(n_29422));
	notech_inv i_32664(.A(n_4729), .Z(n_29423));
	notech_inv i_32665(.A(n_4696), .Z(n_29424));
	notech_inv i_32666(.A(mul64[36]), .Z(n_29425));
	notech_inv i_32667(.A(\regs_1_0[23] ), .Z(n_29426));
	notech_inv i_32668(.A(n_3437), .Z(n_29427));
	notech_inv i_32669(.A(n_3439), .Z(n_29428));
	notech_inv i_32670(.A(n_3440), .Z(n_29429));
	notech_inv i_32671(.A(n_3441), .Z(n_29430));
	notech_inv i_32672(.A(n_3442), .Z(n_29431));
	notech_inv i_32673(.A(n_3392), .Z(n_29432));
	notech_inv i_32674(.A(n_3396), .Z(n_29433));
	notech_inv i_32675(.A(n_3398), .Z(n_29434));
	notech_inv i_32676(.A(n_3400), .Z(n_29435));
	notech_inv i_32677(.A(n_3402), .Z(n_29436));
	notech_inv i_32678(.A(\regs_1_0[19] ), .Z(n_29437));
	notech_inv i_32679(.A(\regs_1_0[20] ), .Z(n_29438));
	notech_inv i_32680(.A(\regs_1_0[21] ), .Z(n_29439));
	notech_inv i_32681(.A(\regs_1_0[22] ), .Z(n_29440));
	notech_inv i_32682(.A(n_3432), .Z(n_29441));
	notech_inv i_32683(.A(n_3433), .Z(n_29442));
	notech_inv i_32684(.A(n_3434), .Z(n_29443));
	notech_inv i_32685(.A(n_3435), .Z(n_29444));
	notech_inv i_32686(.A(n_3436), .Z(n_29447));
	notech_inv i_32687(.A(n_3382), .Z(n_29448));
	notech_inv i_32688(.A(n_3384), .Z(n_29449));
	notech_inv i_32689(.A(n_3386), .Z(n_29450));
	notech_inv i_32690(.A(n_3388), .Z(n_29451));
	notech_inv i_32691(.A(n_3390), .Z(n_29452));
	notech_inv i_32694(.A(n_6350), .Z(n_29453));
	notech_inv i_32695(.A(n_6349), .Z(n_29454));
	notech_inv i_32696(.A(n_6412), .Z(n_29455));
	notech_inv i_32697(.A(n_5184), .Z(n_29456));
	notech_inv i_32698(.A(n_6411), .Z(n_29457));
	notech_inv i_32699(.A(mul64[62]), .Z(n_29458));
	notech_inv i_32700(.A(mul64[60]), .Z(n_29459));
	notech_inv i_32701(.A(mul64[63]), .Z(n_29460));
	notech_inv i_32702(.A(mul64[59]), .Z(n_29461));
	notech_inv i_32703(.A(mul64[61]), .Z(n_29462));
	notech_inv i_32704(.A(mul64[48]), .Z(n_29463));
	notech_inv i_32705(.A(mul64[57]), .Z(n_29464));
	notech_inv i_32706(.A(mul64[55]), .Z(n_29465));
	notech_inv i_32707(.A(mul64[54]), .Z(n_29470));
	notech_inv i_32708(.A(mul64[53]), .Z(n_29471));
	notech_inv i_32709(.A(mul64[52]), .Z(n_29472));
	notech_inv i_32710(.A(mul64[51]), .Z(n_29473));
	notech_inv i_32711(.A(mul64[50]), .Z(n_29475));
	notech_inv i_32712(.A(mul64[49]), .Z(n_29476));
	notech_inv i_32713(.A(mul64[47]), .Z(n_29477));
	notech_inv i_32714(.A(mul64[46]), .Z(n_29478));
	notech_inv i_32715(.A(mul64[44]), .Z(n_29479));
	notech_inv i_32716(.A(mul64[43]), .Z(n_29480));
	notech_inv i_32717(.A(mul64[41]), .Z(n_29481));
	notech_inv i_32718(.A(mul64[39]), .Z(n_29482));
	notech_inv i_32719(.A(mul64[38]), .Z(n_29483));
	notech_inv i_32720(.A(mul64[37]), .Z(n_29484));
	notech_inv i_32721(.A(n_572), .Z(n_29485));
	notech_inv i_32722(.A(n_573), .Z(n_29486));
	notech_inv i_32723(.A(n_578), .Z(n_29487));
	notech_inv i_32724(.A(n_5802), .Z(n_29488));
	notech_inv i_32725(.A(n_5800), .Z(n_29489));
	notech_inv i_32726(.A(n_5810), .Z(n_29490));
	notech_inv i_32727(.A(n_5811), .Z(n_29491));
	notech_inv i_32728(.A(n_5815), .Z(n_29492));
	notech_inv i_32729(.A(n_5816), .Z(n_29493));
	notech_inv i_32730(.A(n_5817), .Z(n_29494));
	notech_inv i_32731(.A(n_5821), .Z(n_29495));
	notech_inv i_32732(.A(n_5822), .Z(n_29496));
	notech_inv i_32733(.A(n_5830), .Z(n_29497));
	notech_inv i_32734(.A(n_5831), .Z(n_29498));
	notech_inv i_32735(.A(n_5832), .Z(n_29499));
	notech_inv i_32736(.A(n_5845), .Z(n_29500));
	notech_inv i_32737(.A(n_5846), .Z(n_29501));
	notech_inv i_32738(.A(n_5847), .Z(n_29502));
	notech_inv i_32739(.A(n_5850), .Z(n_29503));
	notech_inv i_32740(.A(n_5851), .Z(n_29504));
	notech_inv i_32741(.A(n_5852), .Z(n_29505));
	notech_inv i_32742(.A(n_5855), .Z(n_29506));
	notech_inv i_32743(.A(n_5856), .Z(n_29507));
	notech_inv i_32744(.A(n_5857), .Z(n_29508));
	notech_inv i_32745(.A(n_5860), .Z(n_29509));
	notech_inv i_32746(.A(n_5861), .Z(n_29510));
	notech_inv i_32747(.A(n_5862), .Z(n_29511));
	notech_inv i_32748(.A(n_5865), .Z(n_29512));
	notech_inv i_32749(.A(n_5866), .Z(n_29513));
	notech_inv i_32750(.A(n_5867), .Z(n_29514));
	notech_inv i_32751(.A(n_5870), .Z(n_29515));
	notech_inv i_32752(.A(n_5871), .Z(n_29516));
	notech_inv i_32753(.A(n_5872), .Z(n_29517));
	notech_inv i_32754(.A(n_5875), .Z(n_29518));
	notech_inv i_32755(.A(n_5876), .Z(n_29519));
	notech_inv i_32756(.A(n_5877), .Z(n_29520));
	notech_inv i_32757(.A(n_5885), .Z(n_29521));
	notech_inv i_32758(.A(n_5886), .Z(n_29522));
	notech_inv i_32759(.A(n_5887), .Z(n_29523));
	notech_inv i_32760(.A(n_5890), .Z(n_29524));
	notech_inv i_32761(.A(n_5891), .Z(n_29525));
	notech_inv i_32762(.A(n_5892), .Z(n_29526));
	notech_inv i_32763(.A(n_5895), .Z(n_29527));
	notech_inv i_32764(.A(n_5896), .Z(n_29528));
	notech_inv i_32765(.A(n_5897), .Z(n_29529));
	notech_inv i_32766(.A(n_5900), .Z(n_29530));
	notech_inv i_32768(.A(n_5901), .Z(n_29531));
	notech_inv i_32770(.A(n_5902), .Z(n_29532));
	notech_inv i_32771(.A(n_5905), .Z(n_29533));
	notech_inv i_32772(.A(n_5906), .Z(n_29534));
	notech_inv i_32775(.A(n_5907), .Z(n_29535));
	notech_inv i_32777(.A(n_5910), .Z(n_29536));
	notech_inv i_32778(.A(n_5911), .Z(n_29537));
	notech_inv i_32779(.A(n_5912), .Z(n_29538));
	notech_inv i_32780(.A(n_5915), .Z(n_29539));
	notech_inv i_32782(.A(n_5916), .Z(n_29540));
	notech_inv i_32783(.A(n_5917), .Z(n_29541));
	notech_inv i_32785(.A(n_5920), .Z(n_29542));
	notech_inv i_32787(.A(n_5921), .Z(n_29543));
	notech_inv i_32788(.A(n_5922), .Z(n_29544));
	notech_inv i_32789(.A(n_5925), .Z(n_29545));
	notech_inv i_32790(.A(n_5926), .Z(n_29546));
	notech_inv i_32791(.A(n_5927), .Z(n_29547));
	notech_inv i_32792(.A(n_5930), .Z(n_29548));
	notech_inv i_32793(.A(n_5931), .Z(n_29549));
	notech_inv i_32794(.A(n_5932), .Z(n_29550));
	notech_inv i_32795(.A(n_5935), .Z(n_29551));
	notech_inv i_32796(.A(n_5936), .Z(n_29552));
	notech_inv i_32797(.A(n_5937), .Z(n_29553));
	notech_inv i_32798(.A(n_5940), .Z(n_29554));
	notech_inv i_32799(.A(n_5941), .Z(n_29555));
	notech_inv i_32800(.A(n_5942), .Z(n_29556));
	notech_inv i_32801(.A(n_5945), .Z(n_29557));
	notech_inv i_32802(.A(n_5946), .Z(n_29558));
	notech_inv i_32803(.A(n_5947), .Z(n_29559));
	notech_inv i_32804(.A(n_5950), .Z(n_29560));
	notech_inv i_32805(.A(n_5951), .Z(n_29561));
	notech_inv i_32806(.A(n_5952), .Z(n_29562));
	notech_inv i_32807(.A(n_5955), .Z(n_29563));
	notech_inv i_32808(.A(n_5957), .Z(n_29564));
	notech_inv i_32809(.A(n_4242), .Z(n_29565));
	notech_inv i_32810(.A(n_4243), .Z(n_29566));
	notech_inv i_32811(.A(n_4244), .Z(n_29567));
	notech_inv i_32812(.A(n_4245), .Z(n_29568));
	notech_inv i_32813(.A(n_4246), .Z(n_29569));
	notech_inv i_32814(.A(n_4247), .Z(n_29570));
	notech_inv i_32815(.A(n_4248), .Z(n_29571));
	notech_inv i_32816(.A(n_4249), .Z(n_29572));
	notech_inv i_32817(.A(n_4250), .Z(n_29573));
	notech_inv i_32818(.A(n_4251), .Z(n_29574));
	notech_inv i_32819(.A(n_4252), .Z(n_29575));
	notech_inv i_32820(.A(n_4253), .Z(n_29576));
	notech_inv i_32821(.A(n_4254), .Z(n_29577));
	notech_inv i_32822(.A(n_4255), .Z(n_29578));
	notech_inv i_32823(.A(n_4256), .Z(n_29579));
	notech_inv i_32824(.A(n_4257), .Z(n_29580));
	notech_inv i_32825(.A(n_4258), .Z(n_29581));
	notech_inv i_32826(.A(n_4259), .Z(n_29582));
	notech_inv i_32827(.A(n_4260), .Z(n_29583));
	notech_inv i_32828(.A(n_4261), .Z(n_29584));
	notech_inv i_32829(.A(n_4262), .Z(n_29585));
	notech_inv i_32830(.A(n_4263), .Z(n_29586));
	notech_inv i_32831(.A(n_4264), .Z(n_29587));
	notech_inv i_32832(.A(n_4265), .Z(n_29588));
	notech_inv i_32833(.A(n_4266), .Z(n_29589));
	notech_inv i_32834(.A(n_4267), .Z(n_29590));
	notech_inv i_32835(.A(n_4268), .Z(n_29591));
	notech_inv i_32836(.A(n_4269), .Z(n_29592));
	notech_inv i_32837(.A(n_4270), .Z(n_29593));
	notech_inv i_32838(.A(n_4271), .Z(n_29594));
	notech_inv i_32839(.A(n_4272), .Z(n_29595));
	notech_inv i_32840(.A(n_4273), .Z(n_29596));
	notech_inv i_32841(.A(n_4274), .Z(n_29597));
	notech_inv i_32842(.A(n_5841), .Z(n_29598));
	notech_inv i_32843(.A(n_5842), .Z(n_29599));
	notech_inv i_32844(.A(n_3354), .Z(n_29600));
	notech_inv i_32845(.A(n_3355), .Z(n_29601));
	notech_inv i_32846(.A(n_4717), .Z(n_29602));
	notech_inv i_32847(.A(\opc_5[25] ), .Z(n_29603));
	notech_inv i_32848(.A(n_4715), .Z(n_29604));
	notech_inv i_32849(.A(\opc_5[23] ), .Z(n_29605));
	notech_inv i_32850(.A(n_4714), .Z(n_29606));
	notech_inv i_32851(.A(\opc_5[22] ), .Z(n_29607));
	notech_inv i_32852(.A(n_4713), .Z(n_29608));
	notech_inv i_32853(.A(\opc_5[21] ), .Z(n_29609));
	notech_inv i_32854(.A(n_4712), .Z(n_29610));
	notech_inv i_32855(.A(\opc_5[20] ), .Z(n_29611));
	notech_inv i_32856(.A(n_4711), .Z(n_29612));
	notech_inv i_32857(.A(\opc_5[19] ), .Z(n_29614));
	notech_inv i_32858(.A(n_4710), .Z(n_29615));
	notech_inv i_32859(.A(\opc_5[18] ), .Z(n_29616));
	notech_inv i_32860(.A(n_4709), .Z(n_29617));
	notech_inv i_32861(.A(\opc_5[17] ), .Z(n_29618));
	notech_inv i_32862(.A(n_4707), .Z(n_29619));
	notech_inv i_32863(.A(\opc_5[15] ), .Z(n_29621));
	notech_inv i_32864(.A(n_4706), .Z(n_29622));
	notech_inv i_32865(.A(\opc_5[14] ), .Z(n_29623));
	notech_inv i_32866(.A(n_4704), .Z(n_29624));
	notech_inv i_32867(.A(n_4703), .Z(n_29625));
	notech_inv i_32868(.A(n_4701), .Z(n_29628));
	notech_inv i_32869(.A(\opc_1[6] ), .Z(n_29630));
	notech_inv i_32870(.A(\opc_5[6] ), .Z(n_29632));
	notech_inv i_32871(.A(n_4698), .Z(n_29633));
	notech_inv i_32872(.A(\opc_1[7] ), .Z(n_29634));
	notech_inv i_32873(.A(\opc_5[7] ), .Z(n_29638));
	notech_inv i_32874(.A(n_5836), .Z(n_29641));
	notech_inv i_32875(.A(\opc_5[5] ), .Z(n_29642));
	notech_inv i_32876(.A(\opc_1[5] ), .Z(n_29643));
	notech_inv i_32877(.A(n_4697), .Z(n_29644));
	notech_inv i_32878(.A(n_5805), .Z(n_29645));
	notech_inv i_32879(.A(n_5806), .Z(n_29646));
	notech_inv i_32880(.A(n_5825), .Z(n_29647));
	notech_inv i_32881(.A(n_5826), .Z(n_29648));
	notech_inv i_32882(.A(n_6635), .Z(n_29649));
	notech_inv i_32883(.A(n_6634), .Z(n_29650));
	notech_inv i_32884(.A(n_6633), .Z(n_29651));
	notech_inv i_32885(.A(n_6632), .Z(n_29652));
	notech_inv i_32886(.A(n_6631), .Z(n_29653));
	notech_inv i_32887(.A(n_6630), .Z(n_29654));
	notech_inv i_32888(.A(n_6629), .Z(n_29655));
	notech_inv i_32889(.A(n_6628), .Z(n_29656));
	notech_inv i_32890(.A(n_6627), .Z(n_29657));
	notech_inv i_32891(.A(n_6626), .Z(n_29658));
	notech_inv i_32892(.A(n_6625), .Z(n_29659));
	notech_inv i_32893(.A(n_6624), .Z(n_29660));
	notech_inv i_32894(.A(n_6623), .Z(n_29661));
	notech_inv i_32895(.A(n_6622), .Z(n_29662));
	notech_inv i_32896(.A(n_6620), .Z(n_29663));
	notech_inv i_32897(.A(n_6619), .Z(n_29664));
	notech_inv i_32898(.A(n_6618), .Z(n_29665));
	notech_inv i_32899(.A(n_6617), .Z(n_29666));
	notech_inv i_32900(.A(n_6616), .Z(n_29667));
	notech_inv i_32901(.A(n_6615), .Z(n_29668));
	notech_inv i_32902(.A(n_6614), .Z(n_29669));
	notech_inv i_32904(.A(n_6613), .Z(n_29670));
	notech_inv i_32905(.A(n_6612), .Z(n_29671));
	notech_inv i_32906(.A(n_6611), .Z(n_29672));
	notech_inv i_32907(.A(n_6610), .Z(n_29673));
	notech_inv i_32908(.A(n_6609), .Z(n_29674));
	notech_inv i_32909(.A(n_6608), .Z(n_29675));
	notech_inv i_32910(.A(n_6607), .Z(n_29676));
	notech_inv i_32911(.A(n_6606), .Z(n_29677));
	notech_inv i_32912(.A(n_6605), .Z(n_29678));
	notech_inv i_32913(.A(n_6572), .Z(n_29679));
	notech_inv i_32915(.A(n_6571), .Z(n_29680));
	notech_inv i_32917(.A(n_6570), .Z(n_29681));
	notech_inv i_32918(.A(n_6569), .Z(n_29682));
	notech_inv i_32920(.A(n_6568), .Z(n_29683));
	notech_inv i_32921(.A(n_6567), .Z(n_29684));
	notech_inv i_32922(.A(n_6566), .Z(n_29685));
	notech_inv i_32923(.A(n_6565), .Z(n_29686));
	notech_inv i_32924(.A(n_6564), .Z(n_29687));
	notech_inv i_32925(.A(n_6563), .Z(n_29688));
	notech_inv i_32926(.A(n_6562), .Z(n_29689));
	notech_inv i_32927(.A(n_6561), .Z(n_29690));
	notech_inv i_32928(.A(n_6560), .Z(n_29691));
	notech_inv i_32929(.A(n_6559), .Z(n_29693));
	notech_inv i_32930(.A(n_6558), .Z(n_29694));
	notech_inv i_32931(.A(n_6557), .Z(n_29695));
	notech_inv i_32932(.A(n_6556), .Z(n_29696));
	notech_inv i_32933(.A(n_6555), .Z(n_29697));
	notech_inv i_32934(.A(n_6554), .Z(n_29698));
	notech_inv i_32935(.A(n_6553), .Z(n_29699));
	notech_inv i_32936(.A(n_6552), .Z(n_29700));
	notech_inv i_32937(.A(n_6551), .Z(n_29701));
	notech_inv i_32938(.A(n_6550), .Z(n_29702));
	notech_inv i_32939(.A(n_6549), .Z(n_29703));
	notech_inv i_32940(.A(n_6548), .Z(n_29704));
	notech_inv i_32941(.A(n_6547), .Z(n_29705));
	notech_inv i_32942(.A(n_6546), .Z(n_29706));
	notech_inv i_32943(.A(n_6545), .Z(n_29707));
	notech_inv i_32944(.A(n_6544), .Z(n_29708));
	notech_inv i_32945(.A(n_6543), .Z(n_29709));
	notech_inv i_32946(.A(n_4178), .Z(n_29710));
	notech_inv i_32947(.A(n_4179), .Z(n_29711));
	notech_inv i_32948(.A(n_4180), .Z(n_29712));
	notech_inv i_32949(.A(n_4181), .Z(n_29713));
	notech_inv i_32950(.A(n_4182), .Z(n_29714));
	notech_inv i_32951(.A(n_4183), .Z(n_29715));
	notech_inv i_32952(.A(n_4184), .Z(n_29716));
	notech_inv i_32953(.A(n_4185), .Z(n_29717));
	notech_inv i_32954(.A(n_4186), .Z(n_29718));
	notech_inv i_32955(.A(n_4187), .Z(n_29719));
	notech_inv i_32956(.A(n_4188), .Z(n_29720));
	notech_inv i_32957(.A(n_4189), .Z(n_29721));
	notech_inv i_32958(.A(n_4190), .Z(n_29722));
	notech_inv i_32959(.A(n_4191), .Z(n_29723));
	notech_inv i_32960(.A(n_4192), .Z(n_29724));
	notech_inv i_32961(.A(n_4193), .Z(n_29725));
	notech_inv i_32962(.A(n_4194), .Z(n_29726));
	notech_inv i_32963(.A(n_4195), .Z(n_29727));
	notech_inv i_32964(.A(n_4196), .Z(n_29728));
	notech_inv i_32965(.A(n_4197), .Z(n_29729));
	notech_inv i_32966(.A(n_4198), .Z(n_29730));
	notech_inv i_32967(.A(n_4199), .Z(n_29731));
	notech_inv i_32968(.A(n_4200), .Z(n_29732));
	notech_inv i_32969(.A(n_4201), .Z(n_29733));
	notech_inv i_32970(.A(n_4202), .Z(n_29734));
	notech_inv i_32971(.A(n_4203), .Z(n_29735));
	notech_inv i_32972(.A(n_4204), .Z(n_29736));
	notech_inv i_32973(.A(n_4205), .Z(n_29737));
	notech_inv i_32974(.A(n_4206), .Z(n_29738));
	notech_inv i_32975(.A(n_4207), .Z(n_29739));
	notech_inv i_32976(.A(n_4208), .Z(n_29740));
	notech_inv i_32977(.A(n_4209), .Z(n_29741));
	notech_inv i_32978(.A(n_4210), .Z(n_29742));
	notech_inv i_32979(.A(n_4211), .Z(n_29743));
	notech_inv i_32980(.A(n_4212), .Z(n_29744));
	notech_inv i_32981(.A(n_4213), .Z(n_29745));
	notech_inv i_32982(.A(n_4214), .Z(n_29746));
	notech_inv i_32983(.A(n_4215), .Z(n_29747));
	notech_inv i_32984(.A(n_4216), .Z(n_29748));
	notech_inv i_32985(.A(n_4217), .Z(n_29749));
	notech_inv i_32986(.A(n_4218), .Z(n_29750));
	notech_inv i_32987(.A(n_4219), .Z(n_29751));
	notech_inv i_32988(.A(n_4220), .Z(n_29752));
	notech_inv i_32989(.A(n_4221), .Z(n_29753));
	notech_inv i_32991(.A(n_4222), .Z(n_29754));
	notech_inv i_32992(.A(n_4223), .Z(n_29755));
	notech_inv i_32993(.A(n_4224), .Z(n_29756));
	notech_inv i_32994(.A(n_4225), .Z(n_29757));
	notech_inv i_32996(.A(n_4226), .Z(n_29758));
	notech_inv i_32997(.A(n_4227), .Z(n_29759));
	notech_inv i_32998(.A(n_4228), .Z(n_29762));
	notech_inv i_32999(.A(n_4229), .Z(n_29763));
	notech_inv i_33000(.A(n_4230), .Z(n_29764));
	notech_inv i_33001(.A(n_4231), .Z(n_29765));
	notech_inv i_33002(.A(n_4232), .Z(n_29766));
	notech_inv i_33003(.A(n_4233), .Z(n_29767));
	notech_inv i_33004(.A(n_4234), .Z(n_29768));
	notech_inv i_33005(.A(n_4235), .Z(n_29769));
	notech_inv i_33006(.A(n_4236), .Z(n_29770));
	notech_inv i_33007(.A(n_4237), .Z(n_29771));
	notech_inv i_33009(.A(n_4238), .Z(n_29773));
	notech_inv i_33010(.A(n_4239), .Z(n_29774));
	notech_inv i_33011(.A(n_4240), .Z(n_29775));
	notech_inv i_33012(.A(n_4241), .Z(n_29777));
	notech_inv i_33013(.A(n_6636), .Z(n_29778));
	notech_inv i_33014(.A(n_6542), .Z(n_29779));
	notech_inv i_33015(.A(n_4723), .Z(n_29780));
	notech_inv i_33016(.A(\opc_5[31] ), .Z(n_29781));
	notech_inv i_33017(.A(n_4722), .Z(n_29782));
	notech_inv i_33018(.A(\opc_5[30] ), .Z(n_29783));
	notech_inv i_33019(.A(n_4721), .Z(n_29784));
	notech_inv i_33020(.A(\opc_5[29] ), .Z(n_29785));
	notech_inv i_33021(.A(n_4720), .Z(n_29786));
	notech_inv i_33022(.A(\opc_5[28] ), .Z(n_29787));
	notech_inv i_33023(.A(n_4719), .Z(n_29788));
	notech_inv i_33024(.A(\opc_5[27] ), .Z(n_29789));
	notech_inv i_33025(.A(n_4708), .Z(n_29790));
	notech_inv i_33026(.A(\opc_5[16] ), .Z(n_29791));
	notech_inv i_33027(.A(n_60419), .Z(n_29792));
	notech_inv i_33028(.A(n_6700), .Z(n_29793));
	notech_inv i_33029(.A(n_6699), .Z(n_29794));
	notech_inv i_33030(.A(n_6698), .Z(n_29795));
	notech_inv i_33031(.A(n_6696), .Z(n_29796));
	notech_inv i_33032(.A(n_6695), .Z(n_29797));
	notech_inv i_33033(.A(n_6694), .Z(n_29799));
	notech_inv i_33034(.A(n_6693), .Z(n_29800));
	notech_inv i_33035(.A(n_6692), .Z(n_29801));
	notech_inv i_33036(.A(n_6691), .Z(n_29803));
	notech_inv i_33037(.A(n_6690), .Z(n_29804));
	notech_inv i_33038(.A(n_6689), .Z(n_29805));
	notech_inv i_33039(.A(n_6688), .Z(n_29806));
	notech_inv i_33040(.A(n_6687), .Z(n_29807));
	notech_inv i_33041(.A(n_6686), .Z(n_29808));
	notech_inv i_33042(.A(n_6685), .Z(n_29809));
	notech_inv i_33043(.A(n_6684), .Z(n_29811));
	notech_inv i_33044(.A(n_6683), .Z(n_29812));
	notech_inv i_33045(.A(n_6682), .Z(n_29815));
	notech_inv i_33046(.A(n_6681), .Z(n_29817));
	notech_inv i_33047(.A(n_6680), .Z(n_29819));
	notech_inv i_33048(.A(n_6679), .Z(n_29820));
	notech_inv i_33049(.A(n_6678), .Z(n_29821));
	notech_inv i_33050(.A(n_6677), .Z(n_29822));
	notech_inv i_33051(.A(n_6676), .Z(n_29824));
	notech_inv i_33052(.A(n_6675), .Z(n_29825));
	notech_inv i_33053(.A(n_6674), .Z(n_29827));
	notech_inv i_33054(.A(n_6673), .Z(n_29828));
	notech_inv i_33055(.A(n_6672), .Z(n_29829));
	notech_inv i_33056(.A(n_6671), .Z(n_29830));
	notech_inv i_33057(.A(n_6670), .Z(n_29831));
	notech_inv i_33058(.A(n_6668), .Z(n_29832));
	notech_inv i_33059(.A(n_6666), .Z(n_29833));
	notech_inv i_33060(.A(n_6665), .Z(n_29835));
	notech_inv i_33061(.A(n_6664), .Z(n_29836));
	notech_inv i_33062(.A(n_6663), .Z(n_29837));
	notech_inv i_33063(.A(n_6662), .Z(n_29838));
	notech_inv i_33064(.A(n_6661), .Z(n_29839));
	notech_inv i_33065(.A(n_6660), .Z(n_29840));
	notech_inv i_33066(.A(n_6659), .Z(n_29841));
	notech_inv i_33067(.A(n_6658), .Z(n_29842));
	notech_inv i_33068(.A(n_6657), .Z(n_29843));
	notech_inv i_33069(.A(n_6656), .Z(n_29844));
	notech_inv i_33070(.A(n_6655), .Z(n_29845));
	notech_inv i_33071(.A(n_6654), .Z(n_29846));
	notech_inv i_33072(.A(n_6653), .Z(n_29847));
	notech_inv i_33073(.A(n_6652), .Z(n_29848));
	notech_inv i_33074(.A(n_6651), .Z(n_29849));
	notech_inv i_33075(.A(n_6650), .Z(n_29850));
	notech_inv i_33076(.A(n_6649), .Z(n_29851));
	notech_inv i_33077(.A(n_6648), .Z(n_29852));
	notech_inv i_33078(.A(n_6647), .Z(n_29853));
	notech_inv i_33079(.A(n_6645), .Z(n_29854));
	notech_inv i_33080(.A(n_6644), .Z(n_29855));
	notech_inv i_33081(.A(n_6643), .Z(n_29856));
	notech_inv i_33082(.A(n_6642), .Z(n_29858));
	notech_inv i_33083(.A(n_6641), .Z(n_29859));
	notech_inv i_33084(.A(n_6640), .Z(n_29860));
	notech_inv i_33085(.A(n_6639), .Z(n_29863));
	notech_inv i_33086(.A(n_6638), .Z(n_29864));
	notech_inv i_33087(.A(n_6637), .Z(n_29867));
	notech_inv i_33088(.A(n_6603), .Z(n_29868));
	notech_inv i_33089(.A(n_6602), .Z(n_29870));
	notech_inv i_33090(.A(n_6601), .Z(n_29871));
	notech_inv i_33091(.A(n_6600), .Z(n_29872));
	notech_inv i_33092(.A(n_6599), .Z(n_29873));
	notech_inv i_33093(.A(n_6598), .Z(n_29874));
	notech_inv i_33094(.A(n_6597), .Z(n_29875));
	notech_inv i_33095(.A(n_6596), .Z(n_29876));
	notech_inv i_33096(.A(n_6595), .Z(n_29877));
	notech_inv i_33097(.A(n_6594), .Z(n_29878));
	notech_inv i_33098(.A(n_6593), .Z(n_29879));
	notech_inv i_33099(.A(n_6592), .Z(n_29880));
	notech_inv i_33100(.A(n_6591), .Z(n_29881));
	notech_inv i_33101(.A(n_6590), .Z(n_29882));
	notech_inv i_33102(.A(n_6589), .Z(n_29883));
	notech_inv i_33103(.A(n_6587), .Z(n_29884));
	notech_inv i_33104(.A(n_6586), .Z(n_29885));
	notech_inv i_33105(.A(n_6585), .Z(n_29886));
	notech_inv i_33106(.A(n_6584), .Z(n_29887));
	notech_inv i_33107(.A(n_6583), .Z(n_29888));
	notech_inv i_33108(.A(n_6582), .Z(n_29889));
	notech_inv i_33109(.A(n_6581), .Z(n_29890));
	notech_inv i_33110(.A(n_6580), .Z(n_29891));
	notech_inv i_33111(.A(n_6579), .Z(n_29892));
	notech_inv i_33112(.A(n_6578), .Z(n_29893));
	notech_inv i_33113(.A(n_6577), .Z(n_29894));
	notech_inv i_33114(.A(n_6576), .Z(n_29895));
	notech_inv i_33115(.A(n_6575), .Z(n_29896));
	notech_inv i_33116(.A(n_6574), .Z(n_29897));
	notech_inv i_33117(.A(n_6573), .Z(n_29898));
	notech_inv i_33118(.A(n_6669), .Z(n_29899));
	notech_inv i_33119(.A(n_6667), .Z(n_29900));
	notech_inv i_33120(.A(n_6604), .Z(n_29901));
	AWMUX_16_32_7 i_32206(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14524[31] , \nbus_14524[30] , \nbus_14524[29] , \nbus_14524[28] 
		, \nbus_14524[27] , \nbus_14524[26] , \nbus_14524[25] , \nbus_14524[24] 
		, \nbus_14524[23] , \nbus_14524[22] , \nbus_14524[21] , \nbus_14524[20] 
		, \nbus_14524[19] , \nbus_14524[18] , \nbus_14524[17] , \nbus_14524[16] 
		, \nbus_14524[15] , \nbus_14524[14] , \nbus_14524[13] , \nbus_14524[12] 
		, \nbus_14524[11] , \nbus_14524[10] , \nbus_14524[9] , \nbus_14524[8] 
		, \nbus_14524[7] , \nbus_14524[6] , \nbus_14524[5] , \nbus_14524[4] 
		, \nbus_14524[3] , \nbus_14524[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_55315, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, n_55460, ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[107], n_57157, instrc[105], instrc[104]}), .O0({n_6572
		, n_6571, n_6570, n_6569, n_6568, n_6567, n_6566, n_6565, n_6564
		, n_6563, n_6562, n_6561, n_6560, n_6559, n_6558, n_6557, n_6556
		, n_6555, n_6554, n_6553, n_6552, n_6551, n_6550, n_6549, n_6548
		, n_6547, n_6546, n_6545, n_6544, n_6543, n_6542, n_6541}));
	AWMUX_16_32_6 i_32211(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14524[31] , \nbus_14524[30] , \nbus_14524[29] , \nbus_14524[28] 
		, \nbus_14524[27] , \nbus_14524[26] , \nbus_14524[25] , \nbus_14524[24] 
		, \nbus_14524[23] , \nbus_14524[22] , \nbus_14524[21] , \nbus_14524[20] 
		, \nbus_14524[19] , \nbus_14524[18] , \nbus_14524[17] , \nbus_14524[16] 
		, \nbus_14524[15] , \nbus_14524[14] , \nbus_14524[13] , \nbus_14524[12] 
		, \nbus_14524[11] , \nbus_14524[10] , \nbus_14524[9] , \nbus_14524[8] 
		, \nbus_14524[7] , \nbus_14524[6] , \nbus_14524[5] , \nbus_14524[4] 
		, \nbus_14524[3] , \nbus_14524[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_55315, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, n_55460, ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[103], instrc[102], instrc[101], instrc[100]}), .O0
		({n_6604, n_6603, n_6602, n_6601, n_6600, n_6599, n_6598, n_6597
		, n_6596, n_6595, n_6594, n_6593, n_6592, n_6591, n_6590, n_6589
		, n_6588, n_6587, n_6586, n_6585, n_6584, n_6583, n_6582, n_6581
		, n_6580, n_6579, n_6578, n_6577, n_6576, n_6575, n_6574, n_6573
		}));
	AWMUX_16_32_5 i_32216(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14524[31] , \nbus_14524[30] , \nbus_14524[29] , \nbus_14524[28] 
		, \nbus_14524[27] , \nbus_14524[26] , \nbus_14524[25] , \nbus_14524[24] 
		, \nbus_14524[23] , \nbus_14524[22] , \nbus_14524[21] , \nbus_14524[20] 
		, \nbus_14524[19] , \nbus_14524[18] , \nbus_14524[17] , \nbus_14524[16] 
		, \nbus_14524[15] , \nbus_14524[14] , \nbus_14524[13] , \nbus_14524[12] 
		, \nbus_14524[11] , \nbus_14524[10] , \nbus_14524[9] , \nbus_14524[8] 
		, \nbus_14524[7] , \nbus_14524[6] , \nbus_14524[5] , \nbus_14524[4] 
		, \nbus_14524[3] , \nbus_14524[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_55315, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, n_55460, ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[99], instrc[98], instrc[97], instrc[96]}), .O0({n_6636
		, n_6635, n_6634, n_6633, n_6632, n_6631, n_6630, n_6629, n_6628
		, n_6627, n_6626, n_6625, n_6624, n_6623, n_6622, n_6621, n_6620
		, n_6619, n_6618, n_6617, n_6616, n_6615, n_6614, n_6613, n_6612
		, n_6611, n_6610, n_6609, n_6608, n_6607, n_6606, n_6605}));
	AWMUX_16_32_4 i_32221(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14524[31] , \nbus_14524[30] , \nbus_14524[29] , \nbus_14524[28] 
		, \nbus_14524[27] , \nbus_14524[26] , \nbus_14524[25] , \nbus_14524[24] 
		, \nbus_14524[23] , \nbus_14524[22] , \nbus_14524[21] , \nbus_14524[20] 
		, \nbus_14524[19] , \nbus_14524[18] , \nbus_14524[17] , \nbus_14524[16] 
		, \nbus_14524[15] , \nbus_14524[14] , \nbus_14524[13] , \nbus_14524[12] 
		, \nbus_14524[11] , \nbus_14524[10] , \nbus_14524[9] , \nbus_14524[8] 
		, \nbus_14524[7] , \nbus_14524[6] , \nbus_14524[5] , \nbus_14524[4] 
		, \nbus_14524[3] , \nbus_14524[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_55315, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, n_55460, ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[95], instrc[94], instrc[93], instrc[92]}), .O0({n_6668
		, n_6667, n_6666, n_6665, n_6664, n_6663, n_6662, n_6661, n_6660
		, n_6659, n_6658, n_6657, n_6656, n_6655, n_6654, n_6653, n_6652
		, n_6651, n_6650, n_6649, n_6648, n_6647, n_6646, n_6645, n_6644
		, n_6643, n_6642, n_6641, n_6640, n_6639, n_6638, n_6637}));
	AWMUX_16_32_3 i_32226(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14524[31] , \nbus_14524[30] , \nbus_14524[29] , \nbus_14524[28] 
		, \nbus_14524[27] , \nbus_14524[26] , \nbus_14524[25] , \nbus_14524[24] 
		, \nbus_14524[23] , \nbus_14524[22] , \nbus_14524[21] , \nbus_14524[20] 
		, \nbus_14524[19] , \nbus_14524[18] , \nbus_14524[17] , \nbus_14524[16] 
		, \nbus_14524[15] , \nbus_14524[14] , \nbus_14524[13] , \nbus_14524[12] 
		, \nbus_14524[11] , \nbus_14524[10] , \nbus_14524[9] , \nbus_14524[8] 
		, \nbus_14524[7] , \nbus_14524[6] , \nbus_14524[5] , \nbus_14524[4] 
		, \nbus_14524[3] , \nbus_14524[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_55315, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, n_55460, ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[91], instrc[90], instrc[89], instrc[88]}), .O0({n_6700
		, n_6699, n_6698, n_6697, n_6696, n_6695, n_6694, n_6693, n_6692
		, n_6691, n_6690, n_6689, n_6688, n_6687, n_6686, n_6685, n_6684
		, n_6683, n_6682, n_6681, n_6680, n_6679, n_6678, n_6677, n_6676
		, n_6675, n_6674, n_6673, n_6672, n_6671, n_6670, n_6669}));
	AWMUX_16_32_2 i_32231(.I0(write_data_25), .I1(write_data_26), .I2(write_data_27
		), .I3(write_data_28), .I4(write_data_29), .I5(write_data_30), .I6
		(write_data_31), .I7(write_data_32), .S(all_cnt), .O0(write_data_33
		));
	AWMUX_16_32_1 i_55548(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14524[31] , \nbus_14524[30] , \nbus_14524[29] , \nbus_14524[28] 
		, \nbus_14524[27] , \nbus_14524[26] , \nbus_14524[25] , \nbus_14524[24] 
		, \nbus_14524[23] , \nbus_14524[22] , \nbus_14524[21] , \nbus_14524[20] 
		, \nbus_14524[19] , \nbus_14524[18] , \nbus_14524[17] , \nbus_14524[16] 
		, \nbus_14524[15] , \nbus_14524[14] , \nbus_14524[13] , \nbus_14524[12] 
		, \nbus_14524[11] , \nbus_14524[10] , \nbus_14524[9] , \nbus_14524[8] 
		, \nbus_14524[7] , \nbus_14524[6] , \nbus_14524[5] , \nbus_14524[4] 
		, \nbus_14524[3] , \nbus_14524[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_55315, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, n_55460, ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({instrc[127], instrc[126], instrc[125], instrc[124]}), .O0
		({\regs_13_14[31] , \regs_13_14[30] , \regs_13_14[29] , \regs_13_14[28] 
		, \regs_13_14[27] , \regs_13_14[26] , \regs_13_14[25] , \regs_13_14[24] 
		, \regs_13_14[23] , \regs_13_14[22] , \regs_13_14[21] , \regs_13_14[20] 
		, \regs_13_14[19] , \regs_13_14[18] , \regs_13_14[17] , \regs_13_14[16] 
		, \opa_12[15] , \opa_12[14] , \opa_12[13] , \opa_12[12] , \opa_12[11] 
		, \opa_12[10] , \opa_12[9] , \opa_12[8] , \opa_12[7] , \opa_12[6] 
		, \opa_12[5] , \opa_12[4] , \opa_12[3] , \opa_12[2] , \opa_12[1] 
		, \opa_12[0] }));
	AWMUX_16_32_0 i_55999(.I0(regs_0), .I1(ecx), .I2(regs_2), .I3(regs_3), .I4
		(regs_4), .I5(regs_5), .I6(regs_6), .I7(regs_7), .I8(regs_8), .I9
		({\nbus_14524[31] , \nbus_14524[30] , \nbus_14524[29] , \nbus_14524[28] 
		, \nbus_14524[27] , \nbus_14524[26] , \nbus_14524[25] , \nbus_14524[24] 
		, \nbus_14524[23] , \nbus_14524[22] , \nbus_14524[21] , \nbus_14524[20] 
		, \nbus_14524[19] , \nbus_14524[18] , \nbus_14524[17] , \nbus_14524[16] 
		, \nbus_14524[15] , \nbus_14524[14] , \nbus_14524[13] , \nbus_14524[12] 
		, \nbus_14524[11] , \nbus_14524[10] , \nbus_14524[9] , \nbus_14524[8] 
		, \nbus_14524[7] , \nbus_14524[6] , \nbus_14524[5] , \nbus_14524[4] 
		, \nbus_14524[3] , \nbus_14524[2] , cs[1], cs[0]}), .I10(regs_10
		), .I11(regs_11), .I12(regs_12), .I13({gs[31], gs[30], gs[29], gs
		[28], gs[27], gs[26], gs[25], gs[24], gs[23], gs[22], gs[21], gs
		[20], gs[19], gs[18], gs[17], gs[16], gs[15], gs[14], gs[13], gs
		[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs[6], gs[5], gs[4], gs
		[3], n_55315, gs[1], gs[0]}), .I14(regs_14), .I15({\eflags[31] ,
		 \eflags[30] , \eflags[29] , \eflags[28] , \eflags[27] , \eflags[26] 
		, \eflags[25] , \eflags[24] , \eflags[23] , \eflags[22] , \eflags[21] 
		, \eflags[20] , \eflags[19] , \eflags[18] , \eflags[17] , \eflags[16] 
		, \eflags[15] , \eflags[14] , \eflags[13] , \eflags[12] , \eflags[11] 
		, n_55460, ie, \eflags[8] , \eflags[7] , \eflags[6] , \eflags[5] 
		, \eflags[4] , \eflags[3] , \eflags[2] , \eflags[1] , \eflags[0] 
		}), .S({n_56469, n_56478, n_56487, n_56458}), .O0(opc_10));
	AWDP_INC_201 i_1049(.O0({n_489, n_487, n_485, n_483, n_481, n_479, n_477
		, n_475, n_473, n_471, n_469, n_467, n_465, n_463, n_461, n_459,
		 n_457, n_455, n_453, n_451, n_449, n_447, n_445, n_443, n_441, n_439
		, n_437, n_435, n_433, n_431, n_429, n_427, n_425, n_423, n_421,
		 n_419, n_417, n_415, n_413, n_411, n_409, n_407, n_405, n_403, n_401
		, n_399, n_397, n_395, n_393, n_391, n_389, n_387, n_385, n_383,
		 n_381, n_379, n_377, n_375, n_373, n_371, n_369, n_367, n_365, n_363
		}), .tsc(tsc));
	AWDP_SUB_233 i_999(.O0(regs_4_2), .regs_4(regs_4), .calc_sz({calc_sz[2],
		 calc_sz[1], calc_sz[0]}));
	AWDP_ADD_14 i_998(.O0({n_3445, n_3444, n_3443, n_3442, n_3441, n_3440, n_3439
		, n_3438, n_3437, n_3436, n_3435, n_3434, n_3433, n_3432, n_3431
		, n_3430, n_3429, n_3428, n_3427, n_3426, n_3425, n_3424, n_3423
		, n_3422, n_3421, n_3420, n_3419, n_3418, n_3417, n_3416, n_3415
		, n_3414}), .regs_4(regs_4), .calc_sz({calc_sz[2], calc_sz[1], calc_sz
		[0]}));
	AWDP_ADD_13 i_995(.O0({n_2476, n_2474, n_2472, n_2470, n_2468, n_2466, n_2464
		, n_2462, n_2460, n_2458, n_2456, n_2454, n_2452, n_2450, n_2448
		, n_2446, n_2444, n_2442, n_2440, n_2438, n_2436, n_2434, n_2432
		, n_2430, n_2428, n_2426, n_2424, n_2422, n_2420, n_2418, n_2416
		, n_2414}), .regs_7(regs_7), .opd({opd[31], opd[30], opd[29], opd
		[28], opd[27], opd[26], opd[25], opd[24], opd[23], opd[22], opd[
		21], opd[20], opd[19], opd[18], opd[17], opd[16], opd[15], opd[
		14], opd[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7],
		 opd[6], opd[5], opd[4], opd[3], opd[2], opd[1], n_55341}));
	AWDP_SUB_29 i_994(.O0({n_2477, n_2475, n_2473, n_2471, n_2469, n_2467, n_2465
		, n_2463, n_2461, n_2459, n_2457, n_2455, n_2453, n_2451, n_2449
		, n_2447, n_2445, n_2443, n_2441, n_2439, n_2437, n_2435, n_2433
		, n_2431, n_2429, n_2427, n_2425, n_2423, n_2421, n_2419, n_2417
		, n_2415}), .regs_7(regs_7), .opd(opd));
	shiftbox shiftbox(.shiftop({\opcode[3] , opcode_289113, \opcode[1] , \opcode[0] 
		}), .calc_sz(calc_sz), .ci(\eflags[0] ), .co(nCF_shiftbox), .co4
		(nCF_shift4box), .opa({opa[31], opa[30], opa[29], opa[28], opa[
		27], opa[26], opa[25], opa[24], opa[23], opa[22], opa[21], opa[
		20], opa[19], opa[18], opa[17], opa[16], opa[15], opa[14], opa[
		13], opa[12], opa[11], opa[10], opa[9], opa[8], n_59744, n_59735
		, opa[5], n_59726, opa[3], n_59717, n_59708, n_59699}), .opb(opb
		), .resa(resa_shiftbox), .resb(resb_shiftbox), .resa4(resa_shift4box
		), .resb4(resb_shift4box));
	AWMUX_16_1 i_978(.I0(\eflags[11] ), .I2(\eflags[0] ), .I4(\eflags[6] ), 
		.I6(\cond[6] ), .I8(\eflags[7] ), .I10(\eflags[2] ), .I12(\cond[12] 
		), .I14(\cond[14] ), .S({\opcode[3] , n_62409, n_62437, n_62395}
		), .O0(cond_1));
	AWDP_ADD_97 i_976(.add_len_pc32(add_len_pc32), .regs_14(regs_14), .lenpc
		(lenpc));
	AWDP_ADD_25 i_975(.add_len_pc16({n_571, n_570, n_569, n_568, n_567, n_566
		, n_565, n_564, n_563, n_562, n_561, n_560, n_559, n_558, n_557,
		 n_556}), .regs_14({regs_14[15], regs_14[14], regs_14[13], regs_14
		[12], regs_14[11], regs_14[10], regs_14[9], regs_14[8], regs_14[
		7], regs_14[6], regs_14[5], regs_14[4], regs_14[3], regs_14[2], regs_14
		[1], regs_14[0]}), .lenpc({lenpc[15], lenpc[14], lenpc[13], lenpc
		[12], lenpc[11], lenpc[10], lenpc[9], lenpc[8], lenpc[7], lenpc[
		6], lenpc[5], lenpc[4], lenpc[3], lenpc[2], lenpc[1], lenpc[0]})
		);
	AWDP_ADD_198 i_974(.O0({n_6825, n_6824, n_6823, n_6822, n_6821, n_6820, n_6819
		, n_6818, n_6817, n_6816, n_6815, n_6814, n_6813, n_6812, n_6811
		, n_6810, n_6809, n_6808, n_6807, n_6806, n_6805, n_6804, n_6803
		, n_6802, n_6801, n_6800, n_6799, n_6798, n_6797, n_6796, n_6795
		, n_6794}), .I0(nbus_11313), .add_len_pc({\add_len_pc[31] , n_352565814
		, n_352465813, \add_len_pc[28] , \add_len_pc[27] , \add_len_pc[26] 
		, \add_len_pc[25] , \add_len_pc[24] , \add_len_pc[23] , \add_len_pc[22] 
		, \add_len_pc[21] , \add_len_pc[20] , \add_len_pc[19] , \add_len_pc[18] 
		, \add_len_pc[17] , n_271788738, \add_len_pc[15] , \add_len_pc[14] 
		, \add_len_pc[13] , \add_len_pc[12] , \add_len_pc[11] , \add_len_pc[10] 
		, n_353169303, \add_len_pc[8] , n_2676, n_319788492, \add_len_pc[5] 
		, n_319688493, \add_len_pc[3] , \add_len_pc[2] , \add_len_pc[1] 
		, \add_len_pc[0] }));
	AWDP_EQ_86 i_950(.O0({n_572}), .mul64({mul64[63], mul64[62], mul64[61], mul64
		[60], mul64[59], mul64[58], mul64[57], mul64[56], mul64[55], mul64
		[54], mul64[53], mul64[52], mul64[51], mul64[50], mul64[49], mul64
		[48], mul64[47], mul64[46], mul64[45], mul64[44], mul64[43], mul64
		[42], mul64[41], mul64[40], mul64[39], mul64[38], mul64[37], mul64
		[36], mul64[35], mul64[34], mul64[33], mul64[32], mul64[31], mul64
		[30], mul64[29], mul64[28], mul64[27], mul64[26], mul64[25], mul64
		[24], mul64[23], mul64[22], mul64[21], mul64[20], mul64[19], mul64
		[18], mul64[17], mul64[16], mul64[15], mul64[14], mul64[13], mul64
		[12], mul64[11], mul64[10], mul64[9], mul64[8]}));
	AWDP_EQ_130 i_949(.O0({n_573}), .mul64({mul64[63], mul64[62], mul64[61],
		 mul64[60], mul64[59], mul64[58], mul64[57], mul64[56], mul64[55
		], mul64[54], mul64[53], mul64[52], mul64[51], mul64[50], mul64[
		49], mul64[48], mul64[47], mul64[46], mul64[45], mul64[44], mul64
		[43], mul64[42], mul64[41], mul64[40], mul64[39], mul64[38], mul64
		[37], mul64[36], mul64[35], mul64[34], mul64[33], mul64[32], mul64
		[31], mul64[30], mul64[29], mul64[28], mul64[27], mul64[26], mul64
		[25], mul64[24], mul64[23], mul64[22], mul64[21], mul64[20], mul64
		[19], mul64[18], mul64[17], mul64[16]}));
	AWDP_EQ_58112339 i_946(.O0({n_576}), .mul64({mul64[63], mul64[62], mul64
		[61], mul64[60], mul64[59], mul64[58], mul64[57], mul64[56], mul64
		[55], mul64[54], mul64[53], mul64[52], mul64[51], mul64[50], mul64
		[49], mul64[48], mul64[47], mul64[46], mul64[45], mul64[44], mul64
		[43], mul64[42], mul64[41], mul64[40], mul64[39], mul64[38], mul64
		[37], mul64[36], mul64[35], mul64[34], mul64[33], mul64[32], mul64
		[31], mul64[30], mul64[29], mul64[28], mul64[27], mul64[26], mul64
		[25], mul64[24], mul64[23], mul64[22], mul64[21], mul64[20], mul64
		[19], mul64[18], mul64[17], mul64[16], mul64[15], mul64[14], mul64
		[13], mul64[12], mul64[11], mul64[10], mul64[9], mul64[8]}));
	AWDP_EQ_153 i_944(.O0({n_578}), .mul64({mul64[63], mul64[62], mul64[61],
		 mul64[60], mul64[59], mul64[58], mul64[57], mul64[56], mul64[55
		], mul64[54], mul64[53], mul64[52], mul64[51], mul64[50], mul64[
		49], mul64[48], mul64[47], mul64[46], mul64[45], mul64[44], mul64
		[43], mul64[42], mul64[41], mul64[40], mul64[39], mul64[38], mul64
		[37], mul64[36], mul64[35], mul64[34], mul64[33], mul64[32], mul64
		[31], mul64[30], mul64[29], mul64[28], mul64[27], mul64[26], mul64
		[25], mul64[24], mul64[23], mul64[22], mul64[21], mul64[20], mul64
		[19], mul64[18], mul64[17], mul64[16]}));
	AWDP_EQ_125 i_942(.O0({n_580}), .mul64({mul64[63], mul64[62], mul64[61],
		 mul64[60], mul64[59], mul64[58], mul64[57], mul64[56], mul64[55
		], mul64[54], mul64[53], mul64[52], mul64[51], mul64[50], mul64[
		49], mul64[48], mul64[47], mul64[46], mul64[45], mul64[44], mul64
		[43], mul64[42], mul64[41], mul64[40], mul64[39], mul64[38], mul64
		[37], mul64[36], mul64[35], mul64[34], mul64[33], mul64[32]}));
	AWDP_ADD_122 i_936(.O0(nbus_134), .opa({opa[31], opa[30], opa[29], opa[
		28], opa[27], opa[26], opa[25], opa[24], opa[23], opa[22], opa[
		21], opa[20], opa[19], opa[18], opa[17], opa[16], opa[15], opa[
		14], opa[13], opa[12], opa[11], opa[10], opa[9], opa[8], n_59744
		, n_59735, opa[5], n_59726, opa[3], n_59717, n_59708, n_59699}),
		 .opd({opd[31], opd[30], opd[29], opd[28], opd[27], opd[26], opd
		[25], opd[24], opd[23], opd[22], opd[21], opd[20], opd[19], opd[
		18], opd[17], opd[16], opd[15], opd[14], opd[13], opd[12], opd[
		11], opd[10], opd[9], opd[8], opd[7], opd[6], opd[5], n_58547, n_58566
		, n_55298, n_55330, n_55341}));
	AWDP_ADD_139 i_934(.O0(nbus_135), .opa({opa[15], opa[14], opa[13], opa[
		12], opa[11], opa[10], opa[9], opa[8], n_59744, n_59735, opa[5],
		 n_59726, opa[3], n_59717, n_59708, n_59699}), .opd({opd[15], opd
		[14], opd[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7]
		, opd[6], opd[5], n_58547, n_58566, n_55298, n_55330, n_55341})
		);
	AWDP_ADD_194 i_933(.O0(nbus_136), .opa({n_59744, n_59735, opa[5], n_59726
		, opa[3], n_59717, n_59708, n_59699}), .opd({opd[7], opd[6], opd
		[5], opd[4], opd[3], opd[2], opd[1], opd[0]}));
	AWDP_ADD_100 i_932(.O0(nbus_137), .opb(opb), .I0({UNCONNECTED_000, 
		UNCONNECTED_001, UNCONNECTED_002, UNCONNECTED_003, 
		UNCONNECTED_004, UNCONNECTED_005, UNCONNECTED_006, 
		UNCONNECTED_007, UNCONNECTED_008, UNCONNECTED_009, 
		UNCONNECTED_010, UNCONNECTED_011, UNCONNECTED_012, n_57157, 
		UNCONNECTED_013, UNCONNECTED_014, UNCONNECTED_015, 
		UNCONNECTED_016, UNCONNECTED_017, UNCONNECTED_018, 
		UNCONNECTED_019, UNCONNECTED_020, UNCONNECTED_021, 
		UNCONNECTED_022, UNCONNECTED_023, UNCONNECTED_024, 
		UNCONNECTED_025, UNCONNECTED_026, UNCONNECTED_027, 
		UNCONNECTED_028, instrc[105], instrc[104]}));
	AWDP_ADD_60 i_931(.O0(nbus_138), .opb({opb[15], opb[14], opb[13], opb[12
		], opb[11], opb[10], opb[9], opb[8], opb[7], opb[6], opb[5], opb
		[4], opb[3], opb[2], opb[1], opb[0]}), .I0({n_57161, 
		UNCONNECTED_029, UNCONNECTED_030, UNCONNECTED_031, 
		UNCONNECTED_032, UNCONNECTED_033, UNCONNECTED_034, 
		UNCONNECTED_035, UNCONNECTED_036, UNCONNECTED_037, 
		UNCONNECTED_038, UNCONNECTED_039, UNCONNECTED_040, 
		UNCONNECTED_041, instrc[105], instrc[104]}));
	AWDP_ADD_47 i_930(.O0(nbus_139), .opa({opa[31], opa[30], opa[29], opa[28
		], opa[27], opa[26], opa[25], opa[24], opa[23], opa[22], opa[21]
		, opa[20], opa[19], opa[18], opa[17], opa[16], opa[15], opa[14],
		 opa[13], opa[12], opa[11], opa[10], opa[9], opa[8], n_59744, n_59735
		, opa[5], n_59726, opa[3], n_59717, n_59708, n_59699}), .I0({
		UNCONNECTED_042, UNCONNECTED_043, UNCONNECTED_044, 
		UNCONNECTED_045, UNCONNECTED_046, UNCONNECTED_047, 
		UNCONNECTED_048, UNCONNECTED_049, UNCONNECTED_050, 
		UNCONNECTED_051, UNCONNECTED_052, UNCONNECTED_053, n_57162, 
		UNCONNECTED_054, UNCONNECTED_055, UNCONNECTED_056, 
		UNCONNECTED_057, UNCONNECTED_058, UNCONNECTED_059, 
		UNCONNECTED_060, UNCONNECTED_061, UNCONNECTED_062, 
		UNCONNECTED_063, UNCONNECTED_064, UNCONNECTED_065, 
		UNCONNECTED_066, UNCONNECTED_067, UNCONNECTED_068, 
		UNCONNECTED_069, UNCONNECTED_070, instrc[105], instrc[104]}));
	AWDP_ADD_136 i_929(.O0(nbus_140), .opa({opa[15], opa[14], opa[13], opa[
		12], opa[11], opa[10], opa[9], opa[8], n_59744, n_59735, opa[5],
		 n_59726, opa[3], n_59717, n_59708, n_59699}), .I0({
		UNCONNECTED_071, UNCONNECTED_072, n_57156, UNCONNECTED_073, 
		UNCONNECTED_074, UNCONNECTED_075, UNCONNECTED_076, 
		UNCONNECTED_077, UNCONNECTED_078, UNCONNECTED_079, 
		UNCONNECTED_080, UNCONNECTED_081, UNCONNECTED_082, 
		UNCONNECTED_083, instrc[105], instrc[104]}));
	AWDP_SUB_41 i_928(.O0(nbus_141), .opa({opa[31], opa[30], opa[29], opa[28
		], opa[27], opa[26], opa[25], opa[24], opa[23], opa[22], opa[21]
		, opa[20], opa[19], opa[18], opa[17], opa[16], opa[15], opa[14],
		 opa[13], opa[12], opa[11], opa[10], opa[9], opa[8], n_59744, n_59735
		, opa[5], n_59726, opa[3], n_59717, n_59708, n_59699}), .I0({
		UNCONNECTED_084, UNCONNECTED_085, UNCONNECTED_086, 
		UNCONNECTED_087, UNCONNECTED_088, UNCONNECTED_089, 
		UNCONNECTED_090, UNCONNECTED_091, UNCONNECTED_092, 
		UNCONNECTED_093, UNCONNECTED_094, UNCONNECTED_095, n_57157, 
		UNCONNECTED_096, UNCONNECTED_097, UNCONNECTED_098, 
		UNCONNECTED_099, UNCONNECTED_100, UNCONNECTED_101, 
		UNCONNECTED_102, UNCONNECTED_103, UNCONNECTED_104, 
		UNCONNECTED_105, UNCONNECTED_106, UNCONNECTED_107, 
		UNCONNECTED_108, UNCONNECTED_109, UNCONNECTED_110, 
		UNCONNECTED_111, UNCONNECTED_112, instrc[105], instrc[104]}));
	AWDP_SUB_205 i_927(.O0(nbus_142), .opa({opa[15], opa[14], opa[13], opa[
		12], opa[11], opa[10], opa[9], opa[8], n_59744, n_59735, opa[5],
		 n_59726, opa[3], n_59717, n_59708, n_59699}), .I0({
		UNCONNECTED_113, UNCONNECTED_114, n_57157, UNCONNECTED_115, 
		UNCONNECTED_116, UNCONNECTED_117, UNCONNECTED_118, 
		UNCONNECTED_119, UNCONNECTED_120, UNCONNECTED_121, 
		UNCONNECTED_122, UNCONNECTED_123, UNCONNECTED_124, 
		UNCONNECTED_125, instrc[105], instrc[104]}));
	AWDP_ADD_81 i_926(.O0(nbus_143), .opd({opd[31], opd[30], opd[29], opd[28
		], opd[27], opd[26], opd[25], opd[24], opd[23], opd[22], opd[21]
		, opd[20], opd[19], opd[18], opd[17], opd[16], opd[15], opd[14],
		 opd[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7], opd
		[6], opd[5], n_58547, n_58566, n_55298, n_55330, n_55341}), .I0(
		{UNCONNECTED_126, UNCONNECTED_127, UNCONNECTED_128, 
		UNCONNECTED_129, UNCONNECTED_130, UNCONNECTED_131, 
		UNCONNECTED_132, UNCONNECTED_133, UNCONNECTED_134, 
		UNCONNECTED_135, UNCONNECTED_136, UNCONNECTED_137, 
		UNCONNECTED_138, UNCONNECTED_139, UNCONNECTED_140, 
		UNCONNECTED_141, UNCONNECTED_142, UNCONNECTED_143, 
		UNCONNECTED_144, UNCONNECTED_145, UNCONNECTED_146, 
		UNCONNECTED_147, UNCONNECTED_148, UNCONNECTED_149, 
		UNCONNECTED_150, UNCONNECTED_151, UNCONNECTED_152, n_57155, 
		UNCONNECTED_153, UNCONNECTED_154, instrc[105], instrc[104]}));
	AWDP_ADD_6 i_925(.O0(nbus_144), .opd({opd[15], opd[14], opd[13], opd[12]
		, opd[11], opd[10], opd[9], opd[8], opd[7], opd[6], opd[5], n_58547
		, n_58566, n_55298, n_55330, n_55341}), .I0({UNCONNECTED_155, 
		UNCONNECTED_156, UNCONNECTED_157, UNCONNECTED_158, 
		UNCONNECTED_159, UNCONNECTED_160, UNCONNECTED_161, 
		UNCONNECTED_162, UNCONNECTED_163, UNCONNECTED_164, 
		UNCONNECTED_165, n_57155, UNCONNECTED_166, UNCONNECTED_167, instrc
		[105], instrc[104]}));
	AWDP_LSH_43 i_924(.O0(nbus_11279), .opb({opb[4], opb[3], opb[2], opb[1],
		 opb[0]}));
	AWDP_ADD_207 i_809(.O0({n_3408, n_3406, n_3404, n_3402, n_3400, n_3398, n_3396
		, n_3394, n_3392, n_3390, n_3388, n_3386, n_3384, n_3382, n_3380
		, n_3378, n_3376, n_3374, n_3372, n_3370, n_3368, n_3366, n_3364
		, n_3362, n_3360, n_3358, n_3356, n_3354, n_3352, n_3350, n_3348
		, n_3346}), .regs_6(regs_6), .opd(opd));
	AWDP_SUB_17 i_808(.O0({n_3409, n_3407, n_3405, n_3403, n_3401, n_3399, n_3397
		, n_3395, n_3393, n_3391, n_3389, n_3387, n_3385, n_3383, n_3381
		, n_3379, n_3377, n_3375, n_3373, n_3371, n_3369, n_3367, n_3365
		, n_3363, n_3361, n_3359, n_3357, n_3355, n_3353, n_3351, n_3349
		, n_3347}), .regs_6(regs_6), .opd({opd[31], opd[30], opd[29], opd
		[28], opd[27], opd[26], opd[25], opd[24], opd[23], opd[22], opd[
		21], opd[20], opd[19], opd[18], opd[17], opd[16], opd[15], opd[
		14], opd[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7],
		 opd[6], opd[5], n_58547, opd[3], opd[2], n_55330, n_55341}));
	AWDP_ADD_185 i_778(.O0({n_5955, n_5950, n_5945, n_5940, n_5935, n_5930, n_5925
		, n_5920, n_5915, n_5910, n_5905, n_5900, n_5895, n_5890, n_5885
		, n_5880, n_5875, n_5870, n_5865, n_5860, n_5855, n_5850, n_5845
		, n_5840, n_5835, n_5830, n_5825, n_5820, n_5815, n_5810, n_5805
		, n_5800}), .opb(opb), .I0({UNCONNECTED_168, UNCONNECTED_169, 
		UNCONNECTED_170, UNCONNECTED_171, UNCONNECTED_172, 
		UNCONNECTED_173, UNCONNECTED_174, UNCONNECTED_175, 
		UNCONNECTED_176, UNCONNECTED_177, UNCONNECTED_178, 
		UNCONNECTED_179, UNCONNECTED_180, UNCONNECTED_181, 
		UNCONNECTED_182, UNCONNECTED_183, UNCONNECTED_184, 
		UNCONNECTED_185, UNCONNECTED_186, UNCONNECTED_187, 
		UNCONNECTED_188, UNCONNECTED_189, UNCONNECTED_190, 
		UNCONNECTED_191, n_59744, n_59735, opa[5], n_59726, opa[3], n_59717
		, n_59708, n_59699}));
	AWDP_ADD_0 i_776(.O0({n_5957, n_5951, n_5946, n_5941, n_5936, n_5931, n_5926
		, n_5921, n_5916, n_5911, n_5906, n_5901, n_5896, n_5891, n_5886
		, n_5881, n_5876, n_5871, n_5866, n_5861, n_5856, n_5851, n_5846
		, n_5841, n_5836, n_5831, n_5826, n_5821, n_5816, n_5811, n_5806
		, n_5801}), .opd({opd[31], opd[30], opd[29], opd[28], opd[27], opd
		[26], opd[25], opd[24], opd[23], opd[22], opd[21], opd[20], opd[
		19], opd[18], opd[17], opd[16], opd[15], opd[14], opd[13], opd[
		12], opd[11], opd[10], opd[9], opd[8], opd[7], opd[6], opd[5], n_58547
		, n_58566, opd[2], n_55330, n_55341}), .I0({UNCONNECTED_192, 
		UNCONNECTED_193, UNCONNECTED_194, opc[31], opc[30], opc[29], opc
		[28], opc[27], opc[26], opc[25], opc[24], opc[23], opc[22], opc[
		21], opc[20], opc[19], opc[18], opc[17], opc[16], opc[15], opc[
		14], opc[13], opc[12], opc[11], opc[10], opc[9], opc[8], opc[7],
		 opc[6], opc[5], UNCONNECTED_195, UNCONNECTED_196}));
	AWDP_ADD_36 i_775(.O0({n_5958, n_5952, n_5947, n_5942, n_5937, n_5932, n_5927
		, n_5922, n_5917, n_5912, n_5907, n_5902, n_5897, n_5892, n_5887
		, n_5882, n_5877, n_5872, n_5867, n_5862, n_5857, n_5852, n_5847
		, n_5842, n_5837, n_5832, n_5827, n_5822, n_5817, n_5812, n_5807
		, n_5802}), .opd({opd[31], opd[30], opd[29], opd[28], opd[27], opd
		[26], opd[25], opd[24], opd[23], opd[22], opd[21], opd[20], opd[
		19], opd[18], opd[17], opd[16], opd[15], opd[14], opd[13], opd[
		12], opd[11], opd[10], opd[9], opd[8], opd[7], opd[6], opd[5], n_58547
		, n_58566, n_55298, n_55330, n_55341}));
	AWDP_INC_148 i_772(.O0({n_4241, n_4240, n_4239, n_4238, n_4237, n_4236, n_4235
		, n_4234, n_4233, n_4232, n_4231, n_4230, n_4229, n_4228, n_4227
		, n_4226, n_4225, n_4224, n_4223, n_4222, n_4221, n_4220, n_4219
		, n_4218, n_4217, n_4216, n_4215, n_4214, n_4213, n_4212, n_4211
		, n_4210, n_4209, n_4208, n_4207, n_4206, n_4205, n_4204, n_4203
		, n_4202, n_4201, n_4200, n_4199, n_4198, n_4197, n_4196, n_4195
		, n_4194, n_4193, n_4192, n_4191, n_4190, n_4189, n_4188, n_4187
		, n_4186, n_4185, n_4184, n_4183, n_4182, n_4181, n_4180, n_4179
		, n_4178}), .I0({n_59095, n_59050, n_59104, n_59077, n_59059, n_59068
		, n_59023, n_59086, n_59041, n_59032, n_58996, n_59005, n_59014,
		 n_58969, n_58978, n_58987, nbus_11326[15], nbus_11326[14], nbus_11326
		[13], nbus_11326[12], nbus_11326[11], nbus_11326[10], nbus_11326
		[9], nbus_11326[8], nbus_11326[7], nbus_11326[6], nbus_11326[5],
		 nbus_11326[4], nbus_11326[3], nbus_11326[2], nbus_11326[1], nbus_11326
		[0], n_58951, n_56901, n_56892, n_56883, n_56874, n_56865, n_56856
		, n_56847, n_56838, n_56829, n_56820, n_56811, n_56802, n_56793,
		 n_56784, n_56775, n_56766, n_56757, n_56748, n_56739, n_56730, n_56721
		, n_56712, n_56703, n_57326, n_56694, n_56685, n_56676, n_56667,
		 n_56658, n_56649, n_58960}));
	AWDP_INC_99 i_769(.O0({UNCONNECTED_197, UNCONNECTED_198, UNCONNECTED_199
		, UNCONNECTED_200, UNCONNECTED_201, UNCONNECTED_202, 
		UNCONNECTED_203, UNCONNECTED_204, UNCONNECTED_205, 
		UNCONNECTED_206, UNCONNECTED_207, UNCONNECTED_208, 
		UNCONNECTED_209, UNCONNECTED_210, UNCONNECTED_211, 
		UNCONNECTED_212, UNCONNECTED_213, UNCONNECTED_214, 
		UNCONNECTED_215, UNCONNECTED_216, UNCONNECTED_217, 
		UNCONNECTED_218, UNCONNECTED_219, UNCONNECTED_220, 
		UNCONNECTED_221, UNCONNECTED_222, UNCONNECTED_223, 
		UNCONNECTED_224, UNCONNECTED_225, UNCONNECTED_226, 
		UNCONNECTED_227, n_4274, n_4273, n_4272, n_4271, n_4270, n_4269,
		 n_4268, n_4267, n_4266, n_4265, n_4264, n_4263, n_4262, n_4261,
		 n_4260, n_4259, n_4258, n_4257, n_4256, n_4255, n_4254, n_4253,
		 n_4252, n_4251, n_4250, n_4249, n_4248, n_4247, n_4246, n_4245,
		 n_4244, n_4243, n_4242}), .I0({UNCONNECTED_228, UNCONNECTED_229
		, UNCONNECTED_230, UNCONNECTED_231, UNCONNECTED_232, 
		UNCONNECTED_233, UNCONNECTED_234, UNCONNECTED_235, 
		UNCONNECTED_236, UNCONNECTED_237, UNCONNECTED_238, 
		UNCONNECTED_239, UNCONNECTED_240, UNCONNECTED_241, 
		UNCONNECTED_242, UNCONNECTED_243, UNCONNECTED_244, 
		UNCONNECTED_245, UNCONNECTED_246, UNCONNECTED_247, 
		UNCONNECTED_248, UNCONNECTED_249, UNCONNECTED_250, 
		UNCONNECTED_251, UNCONNECTED_252, UNCONNECTED_253, 
		UNCONNECTED_254, UNCONNECTED_255, UNCONNECTED_256, 
		UNCONNECTED_257, UNCONNECTED_258, UNCONNECTED_259, n_56943, n_55234
		, n_55249, n_55261, n_59328, n_59337, n_59346, n_56207, n_59319,
		 n_55647, n_59310, n_55631, n_55620, n_55609, n_55600, n_55590, n_55578
		, n_55566, n_55552, n_55542, n_55469, n_55438, n_55425, n_55413,
		 n_55400, n_55387, n_55375, n_55365, n_55277, n_55289, n_59753, n_55356
		}));
	AWDP_GE_12 i_766(.O0({n_613}), .divr(divr), .divq(divq));
	AWDP_SUB_174 i_765(.O0(divr_0), .divr(divr), .divq(divq));
	AWDP_LE_209 i_763(.O0({n_614}), .divq(divq), .I0({UNCONNECTED_260, divr[
		63], divr[62], divr[61], divr[60], divr[59], divr[58], divr[57],
		 divr[56], divr[55], divr[54], divr[53], divr[52], divr[51], divr
		[50], divr[49], divr[48], divr[47], divr[46], divr[45], divr[44]
		, divr[43], divr[42], divr[41], divr[40], divr[39], divr[38], divr
		[37], divr[36], divr[35], divr[34], divr[33], divr[32], divr[31]
		, divr[30], divr[29], divr[28], divr[27], divr[26], divr[25], divr
		[24], divr[23], divr[22], divr[21], divr[20], divr[19], divr[18]
		, divr[17], divr[16], divr[15], divr[14], divr[13], divr[12], divr
		[11], divr[10], divr[9], divr[8], divr[7], divr[6], divr[5], divr
		[4], divr[3], divr[2], divr[1]}));
	AWDP_DEC_166 i_759(.O0({\regs_1_0[31] , \regs_1_0[30] , \regs_1_0[29] , \regs_1_0[28] 
		, \regs_1_0[27] , \regs_1_0[26] , \regs_1_0[25] , \regs_1_0[24] 
		, \regs_1_0[23] , \regs_1_0[22] , \regs_1_0[21] , \regs_1_0[20] 
		, \regs_1_0[19] , \regs_1_0[18] , \regs_1_0[17] , \regs_1_0[16] 
		, n_4690, n_4689, n_4688, n_4687, n_4686, n_4685, n_4684, n_4683
		, n_4682, n_4681, n_4680, n_4679, n_4678, n_4677, n_4676, n_4675
		}), .ecx(ecx));
	AWDP_DEC_162 i_758(.O0({\regs_1[15] , \regs_1[14] , \regs_1[13] , \regs_1[12] 
		, \regs_1[11] , \regs_1[10] , \regs_1[9] , \regs_1[8] , \regs_1[7] 
		, \regs_1[6] , \regs_1[5] , \regs_1[4] , \regs_1[3] , \regs_1[2] 
		, \regs_1[1] , \regs_1[0] }), .cx({ecx[15], ecx[14], ecx[13], ecx
		[12], ecx[11], ecx[10], ecx[9], ecx[8], ecx[7], ecx[6], ecx[5], ecx
		[4], ecx[3], ecx[2], ecx[1], ecx[0]}));
	AWDP_LSH_196 i_756(.O0(nbus_11304), .opd({opd[5], n_58547, n_58566, n_55298
		, n_55330, n_55341}));
	AWDP_ADD_195 i_755(.O0(opc_14), .opc({opc[31], opc[30], opc[29], opc[28]
		, opc[27], opc[26], opc[25], opc[24], opc[23], opc[22], opc[21],
		 opc[20], opc[19], opc[18], opc[17], opc[16], opc[15], opc[14], opc
		[13], opc[12], opc[11], opc[10], opc[9], opc[8], opc[7], opc[6],
		 opc[5], opc[4], opc[3], opc[2], opc[1], n_59113}), .I0(nbus_11304
		));
	AWDP_INC_26 i_749(.O0({n_4723, n_4722, n_4721, n_4720, n_4719, n_4718, n_4717
		, n_4716, n_4715, n_4714, n_4713, n_4712, n_4711, n_4710, n_4709
		, n_4708, n_4707, n_4706, n_4705, n_4704, n_4703, n_4702, n_4701
		, n_4700, n_4699, n_4698, n_4697, n_4696, n_4695, n_4694, n_4693
		, n_4692}), .I0(nbus_11348));
	AWDP_DEC_7 i_746(.O0({\opc_1[7] , \opc_1[6] , \opc_1[5] , \opc_1[4] , \opc_1[3] 
		, \opc_1[2] , \opc_1[1] , \opc_1[0] }), .opc({opc[7], opc[6], opc
		[5], opc[4], opc[3], opc[2], opc[1], n_59113}));
	AWDP_DEC_2 i_743(.O0({\opc_5[31] , \opc_5[30] , \opc_5[29] , \opc_5[28] 
		, \opc_5[27] , \opc_5[26] , \opc_5[25] , \opc_5[24] , \opc_5[23] 
		, \opc_5[22] , \opc_5[21] , \opc_5[20] , \opc_5[19] , \opc_5[18] 
		, \opc_5[17] , \opc_5[16] , \opc_5[15] , \opc_5[14] , \opc_5[13] 
		, \opc_5[12] , \opc_5[11] , \opc_5[10] , \opc_5[9] , \opc_5[8] ,
		 \opc_5[7] , \opc_5[6] , \opc_5[5] , n_4729, n_4728, n_4727, n_4726
		, n_4725}), .opc({opc[31], opc[30], opc[29], opc[28], opc[27], opc
		[26], opc[25], opc[24], opc[23], opc[22], opc[21], opc[20], opc[
		19], opc[18], opc[17], opc[16], opc[15], opc[14], opc[13], opc[
		12], opc[11], opc[10], opc[9], opc[8], opc[7], opc[6], opc[5], opc
		[4], opc[3], opc[2], opc[1], n_59113}));
	AWDP_EQ_218 i_738(.O0({n_620}), .I0({opb[31], opb[30], opb[29], opb[28],
		 opb[27], opb[26], opb[25], opb[24], opb[23], opb[22], opb[21], opb
		[20], opb[19], opb[18], opb[17], opb[16], opb[15], opb[14], opb[
		13], opb[12], opb[11], opb[10], opb[9], opb[8], opb[7], opb[6], opb
		[5], opb[4], opb[3], opb[2], opb[1], opb[0], opc[31], opc[30], opc
		[29], opc[28], opc[27], opc[26], opc[25], opc[24], opc[23], opc[
		22], opc[21], opc[20], opc[19], opc[18], opc[17], opc[16], opc[
		15], opc[14], opc[13], opc[12], opc[11], opc[10], opc[9], opc[8]
		, opc[7], opc[6], opc[5], opc[4], opc[3], opc[2], opc[1], n_59113
		}), .I1({regs_2[31], regs_2[30], regs_2[29], regs_2[28], regs_2[
		27], regs_2[26], regs_2[25], regs_2[24], regs_2[23], regs_2[22],
		 regs_2[21], regs_2[20], regs_2[19], regs_2[18], regs_2[17], regs_2
		[16], regs_2[15], regs_2[14], regs_2[13], regs_2[12], regs_2[11]
		, regs_2[10], regs_2[9], regs_2[8], regs_2[7], regs_2[6], regs_2
		[5], regs_2[4], regs_2[3], regs_2[2], regs_2[1], regs_2[0], regs_0
		[31], regs_0[30], regs_0[29], regs_0[28], regs_0[27], regs_0[26]
		, regs_0[25], regs_0[24], regs_0[23], regs_0[22], regs_0[21], regs_0
		[20], regs_0[19], regs_0[18], regs_0[17], regs_0[16], regs_0[15]
		, regs_0[14], regs_0[13], regs_0[12], regs_0[11], regs_0[10], regs_0
		[9], regs_0[8], regs_0[7], regs_0[6], regs_0[5], regs_0[4], regs_0
		[3], regs_0[2], regs_0[1], regs_0[0]}));
	AWDP_INC_235 i_730(.O0(opa_0), .I0({n_58951, n_56901, n_56892, n_56883, n_56874
		, n_56865, n_56856, n_56847, n_56838, n_56829, n_56820, n_56811,
		 n_56802, n_56793, n_56784, n_56775, n_56766, n_56757, n_56748, n_56739
		, n_56730, n_56721, n_56712, n_56703, n_57326, n_56694, n_56685,
		 n_56676, n_56667, n_56658, n_56649, n_58960}));
	AWDP_INC_77 i_728(.O0({\opa_1[15] , \opa_1[14] , \opa_1[13] , \opa_1[12] 
		, \opa_1[11] , \opa_1[10] , \opa_1[9] , \opa_1[8] , \opa_1[7] , \opa_1[6] 
		, \opa_1[5] , \opa_1[4] , \opa_1[3] , \opa_1[2] , \opa_1[1] , \opa_1[0] 
		}), .I0({n_56766, n_56757, n_56748, n_56739, n_56730, n_56721, n_56712
		, n_56703, n_57326, n_56694, n_56685, n_56676, n_56667, n_56658,
		 n_56649, n_58960}));
	AWDP_INC_78 i_717(.O0({n_6314, n_6313, n_6312, n_6311, n_6310, n_6309, n_6308
		, n_6307, n_6306, n_6305, n_6304, n_6303, n_6302, n_6301, n_6300
		, n_6299, n_6298, n_6297, n_6296, n_6295, n_6294, n_6293, n_6292
		, n_6291, n_6290, n_6289, n_6288, n_6287, n_6286, n_6285, n_6284
		, n_6283}), .I0({n_59095, n_59050, n_59104, n_59077, n_59059, n_59068
		, n_59023, n_59086, n_59041, n_59032, n_58996, n_59005, n_59014,
		 n_58969, n_58978, n_58987, nbus_11326[15], nbus_11326[14], nbus_11326
		[13], nbus_11326[12], nbus_11326[11], nbus_11326[10], nbus_11326
		[9], nbus_11326[8], nbus_11326[7], nbus_11326[6], nbus_11326[5],
		 nbus_11326[4], nbus_11326[3], nbus_11326[2], nbus_11326[1], nbus_11326
		[0]}));
	arithbox arithbox(.arithop({\opcode[3] , opcode_289113, \opcode[1] , \opcode[0] 
		}), .calc_sz(calc_sz), .ci(\eflags[0] ), .co(nCF_arithbox), .af(nAF_arithbox
		), .ai(\eflags[4] ), .sa(opas_arithbox), .sb(opbs_arithbox), .opa
		({opa[31], opa[30], opa[29], opa[28], opa[27], opa[26], opa[25],
		 opa[24], opa[23], opa[22], opa[21], opa[20], opa[19], opa[18], opa
		[17], opa[16], opa[15], opa[14], opa[13], opa[12], opa[11], opa[
		10], opa[9], opa[8], n_59744, n_59735, opa[5], n_59726, opa[3], n_59717
		, n_59708, opa[0]}), .opb(opb), .resa(resa_arithbox), .cmp(tcmp_arithbox
		));
	synthetic_op synthetic_op(.clk(clk), .sel({opcode_289113, \opcode[1] , \opcode[0] 
		}), .opa32({opa[31], opa[30], opa[29], opa[28], opa[27], opa[26]
		, opa[25], opa[24], opa[23], opa[22], opa[21], opa[20], opa[19],
		 opa[18], opa[17], opa[16], opa[15], opa[14], opa[13], opa[12], opa
		[11], opa[10], opa[9], opa[8], n_59744, n_59735, opa[5], n_59726
		, opa[3], n_59717, n_59708, opa[0]}), .opb32(opb), .res64(mul64)
		);
	AWDP_ADD_69 i_679(.O0({n_851, n_849, n_847, n_845, n_843, n_841, n_839, n_837
		, n_835, n_833, n_831, n_829, n_827, n_825, n_823, n_821, n_819,
		 n_817, n_815, n_813, n_811, n_809, n_807, n_805, n_803, n_801, n_799
		, n_797, n_795, n_793, n_791, n_789}), .ldtr(ldtr), .I0({gs[31],
		 gs[30], gs[29], gs[28], gs[27], gs[26], gs[25], gs[24], gs[23],
		 gs[22], gs[21], gs[20], gs[19], gs[18], gs[17], gs[16], gs[15],
		 gs[14], gs[13], gs[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs
		[6], gs[5], gs[4], gs[3], UNCONNECTED_261, UNCONNECTED_262, 
		UNCONNECTED_263}));
	AWDP_ADD_22 i_677(.O0({n_852, n_850, n_848, n_846, n_844, n_842, n_840, n_838
		, n_836, n_834, n_832, n_830, n_828, n_826, n_824, n_822, n_820,
		 n_818, n_816, n_814, n_812, n_810, n_808, n_806, n_804, n_802, n_800
		, n_798, n_796, n_794, n_792, n_790}), .gdtr(gdtr), .I0({gs[31],
		 gs[30], gs[29], gs[28], gs[27], gs[26], gs[25], gs[24], gs[23],
		 gs[22], gs[21], gs[20], gs[19], gs[18], gs[17], gs[16], gs[15],
		 gs[14], gs[13], gs[12], gs[11], gs[10], gs[9], gs[8], gs[7], gs
		[6], gs[5], gs[4], gs[3], UNCONNECTED_264, UNCONNECTED_265, 
		UNCONNECTED_266}));
	AWDP_ADD_181 i_674(.O0({n_6411, n_6409, n_6407, n_6405, n_6403, n_6401, n_6399
		, n_6397, n_6395, n_6393, n_6391, n_6389, n_6387, n_6385, n_6383
		, n_6381, n_6379, n_6377, n_6375, n_6373, n_6371, n_6369, n_6367
		, n_6365, n_6363, n_6361, n_6359, n_6357, n_6355, n_6353, n_6351
		, n_6349}), .idtr(idtr), .I0({instrc[95], instrc[94], instrc[93]
		, instrc[92], instrc[91], instrc[90], instrc[89], instrc[88], instrc
		[87], instrc[86], instrc[85], instrc[84], instrc[83], instrc[82]
		, instrc[81], instrc[80], UNCONNECTED_267, UNCONNECTED_268, 
		UNCONNECTED_269}));
	AWDP_ADD_238 i_672(.O0({n_6412, n_6410, n_6408, n_6406, n_6404, n_6402, n_6400
		, n_6398, n_6396, n_6394, n_6392, n_6390, n_6388, n_6386, n_6384
		, n_6382, n_6380, n_6378, n_6376, n_6374, n_6372, n_6370, n_6368
		, n_6366, n_6364, n_6362, n_6360, n_6358, n_6356, n_6354, n_6352
		, n_6350}), .gdtr(gdtr), .I0({\tr[15] , \tr[14] , \tr[13] , \tr[12] 
		, \tr[11] , \tr[10] , \tr[9] , \tr[8] , \tr[7] , \tr[6] , \tr[5] 
		, \tr[4] , \tr[3] , UNCONNECTED_270, UNCONNECTED_271, 
		UNCONNECTED_272}));
	AWDP_SUB_200 i_671(.O0(Daddrs_8), .opd({opd[31], opd[30], opd[29], opd[
		28], opd[27], opd[26], opd[25], opd[24], opd[23], opd[22], opd[
		21], opd[20], opd[19], opd[18], opd[17], opd[16], opd[15], opd[
		14], opd[13], opd[12], opd[11], opd[10], opd[9], opd[8], opd[7],
		 opd[6], opd[5], n_58547, n_58566, n_55298, n_55330, n_55341})
		);
	AWDP_ADD_239 i_670(.O0(Daddrs_1), .Daddrs(Daddr));
	AWDP_ADD_8 i_669(.O0(Daddrs_3), .Daddrs(Daddr));
	AWDP_ADD_241 i_667(.O0({n_5184, n_5183, n_5182, n_5181, n_5180, n_5179, n_5178
		, n_5177, n_5176, n_5175, n_5174, n_5173, n_5172, n_5171, n_5170
		, n_5169, n_5168, n_5167, n_5166, n_5165, n_5164, n_5163, n_5162
		, n_5161, n_5160, n_5159, n_5158, n_5157, n_5156, n_5155, n_5154
		, n_5153}), .opd({opd[31], opd[30], opd[29], opd[28], opd[27], opd
		[26], opd[25], opd[24], opd[23], opd[22], opd[21], opd[20], opd[
		19], opd[18], opd[17], opd[16], opd[15], opd[14], opd[13], opd[
		12], opd[11], opd[10], opd[9], opd[8], opd[7], opd[6], opd[5], n_58547
		, n_58566, n_55298, n_55330, n_55341}), .desc(desc));
	AWDP_ADD_40 i_606(.O0({n_1476, n_1475, n_1474, n_1473, n_1472, n_1471, n_1470
		, n_1469, n_1468, n_1467, n_1466, n_1465, n_1464, n_1463, n_1462
		, n_1461, n_1460, n_1459, n_1458, n_1457, n_1456, n_1455, n_1454
		, n_1453, n_1452, n_1451, n_1450, n_1449, n_1448, n_1447, n_1446
		, n_1445}), .I0({UNCONNECTED_273, UNCONNECTED_274, 
		UNCONNECTED_275, UNCONNECTED_276, UNCONNECTED_277, 
		UNCONNECTED_278, UNCONNECTED_279, UNCONNECTED_280, 
		UNCONNECTED_281, UNCONNECTED_282, UNCONNECTED_283, 
		UNCONNECTED_284, UNCONNECTED_285, UNCONNECTED_286, 
		UNCONNECTED_287, UNCONNECTED_288, regs_14[15], regs_14[14], regs_14
		[13], regs_14[12], regs_14[11], regs_14[10], regs_14[9], regs_14
		[8], regs_14[7], regs_14[6], regs_14[5], regs_14[4], regs_14[3],
		 regs_14[2], regs_14[1], regs_14[0]}), .I1({\nbus_14524[27] , \nbus_14524[26] 
		, \nbus_14524[25] , \nbus_14524[24] , \nbus_14524[23] , \nbus_14524[22] 
		, \nbus_14524[21] , \nbus_14524[20] , \nbus_14524[19] , \nbus_14524[18] 
		, \nbus_14524[17] , \nbus_14524[16] , \nbus_14524[15] , \nbus_14524[14] 
		, \nbus_14524[13] , \nbus_14524[12] , \nbus_14524[11] , \nbus_14524[10] 
		, \nbus_14524[9] , \nbus_14524[8] , \nbus_14524[7] , \nbus_14524[6] 
		, \nbus_14524[5] , \nbus_14524[4] , \nbus_14524[3] , \nbus_14524[2] 
		, cs[1], cs[0], UNCONNECTED_289, UNCONNECTED_290, 
		UNCONNECTED_291, UNCONNECTED_292}));
endmodule
module cpu(clk, rstn, iack, int_cpu, ivect, cr0, cr2, icr2, cr3, cs, pg_fault, ipg_fault
		, useq_ptr, valid_len, queue, pg_en, pc_out, pc_req, read_req, write_req
		, read_ack, write_ack, flush_Itlb, flush_Dtlb, readio_req, writeio_req
		, readio_ack, writeio_ack, write_data, writeio_data, read_data, readio_data
		, write_sz, read_sz, io_add, Daddr, pt_fault, wr_fault);

	input clk;
	input rstn;
	output iack;
	input int_cpu;
	input [7:0] ivect;
	output [31:0] cr0;
	input [31:0] cr2;
	input [31:0] icr2;
	output [31:0] cr3;
	output [31:0] cs;
	input pg_fault;
	input ipg_fault;
	output [3:0] useq_ptr;
	input [5:0] valid_len;
	input [127:0] queue;
	output pg_en;
	output [31:0] pc_out;
	output pc_req;
	output read_req;
	output write_req;
	input read_ack;
	input write_ack;
	output flush_Itlb;
	output flush_Dtlb;
	output readio_req;
	output writeio_req;
	input readio_ack;
	input writeio_ack;
	output [31:0] write_data;
	output [31:0] writeio_data;
	input [31:0] read_data;
	input [31:0] readio_data;
	output [1:0] write_sz;
	output [1:0] read_sz;
	output [31:0] io_add;
	output [31:0] Daddr;
	input pt_fault;
	input wr_fault;

	wire [2:0] reps;
	wire [2:0] opz;
	wire [127:0] dec2vliw;
	wire [31:0] lenpc;
	wire [31:0] add_src;
	wire [7:0] from_acu;
	wire [63:0] to_acu;
	wire [210:0] deco2acu;



	vliw i_vliw(.clk(clk), .rstn(rstn), .instrc(dec2vliw), .ie(ie), .readio_data
		(readio_data), .io_add({UNCONNECTED_000, UNCONNECTED_001, 
		UNCONNECTED_002, UNCONNECTED_003, UNCONNECTED_004, 
		UNCONNECTED_005, UNCONNECTED_006, UNCONNECTED_007, 
		UNCONNECTED_008, UNCONNECTED_009, UNCONNECTED_010, 
		UNCONNECTED_011, UNCONNECTED_012, UNCONNECTED_013, 
		UNCONNECTED_014, UNCONNECTED_015, io_add[15], io_add[14], io_add
		[13], io_add[12], io_add[11], io_add[10], io_add[9], io_add[8], io_add
		[7], io_add[6], io_add[5], io_add[4], io_add[3], io_add[2], io_add
		[1], io_add[0]}), .writeio_data(writeio_data), .writeio_req(writeio_req
		), .readio_req(readio_req), .writeio_ack(writeio_ack), .readio_ack
		(readio_ack), .read_reqs(read_req), .read_ack(read_ack), .read_data
		(read_data), .over_seg({\over_seg[5] , UNCONNECTED_016, 
		UNCONNECTED_017, UNCONNECTED_018, UNCONNECTED_019, 
		UNCONNECTED_020}), .cr3({cr3[31], cr3[30], cr3[29], cr3[28], cr3
		[27], cr3[26], cr3[25], cr3[24], cr3[23], cr3[22], cr3[21], cr3[
		20], cr3[19], cr3[18], cr3[17], cr3[16], cr3[15], cr3[14], cr3[
		13], cr3[12], UNCONNECTED_021, UNCONNECTED_022, UNCONNECTED_023,
		 UNCONNECTED_024, UNCONNECTED_025, UNCONNECTED_026, 
		UNCONNECTED_027, UNCONNECTED_028, UNCONNECTED_029, 
		UNCONNECTED_030, UNCONNECTED_031, UNCONNECTED_032}), .cr2(cr2), 
		.icr2(icr2), .cr0({UNCONNECTED_033, UNCONNECTED_034, 
		UNCONNECTED_035, UNCONNECTED_036, UNCONNECTED_037, 
		UNCONNECTED_038, UNCONNECTED_039, UNCONNECTED_040, 
		UNCONNECTED_041, UNCONNECTED_042, UNCONNECTED_043, 
		UNCONNECTED_044, UNCONNECTED_045, UNCONNECTED_046, 
		UNCONNECTED_047, cr0[16], UNCONNECTED_048, UNCONNECTED_049, 
		UNCONNECTED_050, UNCONNECTED_051, UNCONNECTED_052, 
		UNCONNECTED_053, UNCONNECTED_054, UNCONNECTED_055, 
		UNCONNECTED_056, UNCONNECTED_057, UNCONNECTED_058, 
		UNCONNECTED_059, UNCONNECTED_060, \cr0[2] , UNCONNECTED_061, \cr0[0] 
		}), .write_reqs(write_req), .write_ack(write_ack), .write_data(write_data
		), .Daddr(Daddr), .write_sz(write_sz), .cs({UNCONNECTED_062, 
		UNCONNECTED_063, UNCONNECTED_064, UNCONNECTED_065, 
		UNCONNECTED_066, UNCONNECTED_067, UNCONNECTED_068, 
		UNCONNECTED_069, UNCONNECTED_070, UNCONNECTED_071, 
		UNCONNECTED_072, UNCONNECTED_073, UNCONNECTED_074, 
		UNCONNECTED_075, UNCONNECTED_076, UNCONNECTED_077, 
		UNCONNECTED_078, UNCONNECTED_079, UNCONNECTED_080, 
		UNCONNECTED_081, UNCONNECTED_082, UNCONNECTED_083, 
		UNCONNECTED_084, UNCONNECTED_085, UNCONNECTED_086, 
		UNCONNECTED_087, UNCONNECTED_088, UNCONNECTED_089, 
		UNCONNECTED_090, UNCONNECTED_091, cs[1], cs[0]}), .add_src(add_src
		), .from_acu(from_acu), .to_acu(to_acu), .pg_en(pg_en), .imm({
		UNCONNECTED_092, UNCONNECTED_093, UNCONNECTED_094, 
		UNCONNECTED_095, UNCONNECTED_096, UNCONNECTED_097, 
		UNCONNECTED_098, UNCONNECTED_099, UNCONNECTED_100, 
		UNCONNECTED_101, UNCONNECTED_102, UNCONNECTED_103, 
		UNCONNECTED_104, UNCONNECTED_105, UNCONNECTED_106, 
		UNCONNECTED_107, \imm[47] , \imm[46] , \imm[45] , \imm[44] , \imm[43] 
		, \imm[42] , \imm[41] , \imm[40] , \imm[39] , \imm[38] , \imm[37] 
		, \imm[36] , \imm[35] , \imm[34] , \imm[33] , \imm[32] , \imm[31] 
		, \imm[30] , \imm[29] , \imm[28] , \imm[27] , \imm[26] , \imm[25] 
		, \imm[24] , \imm[23] , \imm[22] , \imm[21] , \imm[20] , \imm[19] 
		, \imm[18] , \imm[17] , \imm[16] , \imm[15] , \imm[14] , \imm[13] 
		, \imm[12] , \imm[11] , \imm[10] , \imm[9] , \imm[8] , \imm[7] ,
		 \imm[6] , \imm[5] , \imm[4] , \imm[3] , \imm[2] , \imm[1] , \imm[0] 
		}), .lenpc(lenpc), .pc_out(pc_out), .pc_req(pc_req), .opz(opz), 
		.reps(reps), .flush_tlb(flush_Itlb), .flush_Dtlb(flush_Dtlb), .terminate
		(term), .start_up(st), .pg_fault(pg_fault), .ipg_fault(ipg_fault
		), .wr_fault(wr_fault), .pt_fault(pt_fault));
	acu i_acu(.clk(clk), .rstn(rstn), .from_regf(to_acu), .add_src(add_src),
		 .to_regf(from_acu), .from_dec(deco2acu), .db67(\cr0[0] ));
	deco i_deco(.clk(clk), .rstn(rstn), .useq_ptr(useq_ptr), .in128(queue), 
		.adz(\cr0[0] ), .pc_req(pc_req), .ivect(ivect), .int_main(int_cpu
		), .iack(iack), .ie(ie), .pg_fault(pg_fault), .ipg_fault(ipg_fault
		), .cpl({cs[1], cs[0]}), .cr0({UNCONNECTED_108, UNCONNECTED_109,
		 UNCONNECTED_110, UNCONNECTED_111, UNCONNECTED_112, 
		UNCONNECTED_113, UNCONNECTED_114, UNCONNECTED_115, 
		UNCONNECTED_116, UNCONNECTED_117, UNCONNECTED_118, 
		UNCONNECTED_119, UNCONNECTED_120, UNCONNECTED_121, 
		UNCONNECTED_122, UNCONNECTED_123, UNCONNECTED_124, 
		UNCONNECTED_125, UNCONNECTED_126, UNCONNECTED_127, 
		UNCONNECTED_128, UNCONNECTED_129, UNCONNECTED_130, 
		UNCONNECTED_131, UNCONNECTED_132, UNCONNECTED_133, 
		UNCONNECTED_134, UNCONNECTED_135, UNCONNECTED_136, \cr0[2] , 
		UNCONNECTED_137, UNCONNECTED_138}), .valid_len(valid_len), .to_vliw
		(dec2vliw), .lenpc_out(lenpc), .immediate({UNCONNECTED_139, 
		UNCONNECTED_140, UNCONNECTED_141, UNCONNECTED_142, 
		UNCONNECTED_143, UNCONNECTED_144, UNCONNECTED_145, 
		UNCONNECTED_146, UNCONNECTED_147, UNCONNECTED_148, 
		UNCONNECTED_149, UNCONNECTED_150, UNCONNECTED_151, 
		UNCONNECTED_152, UNCONNECTED_153, UNCONNECTED_154, \imm[47] , \imm[46] 
		, \imm[45] , \imm[44] , \imm[43] , \imm[42] , \imm[41] , \imm[40] 
		, \imm[39] , \imm[38] , \imm[37] , \imm[36] , \imm[35] , \imm[34] 
		, \imm[33] , \imm[32] , \imm[31] , \imm[30] , \imm[29] , \imm[28] 
		, \imm[27] , \imm[26] , \imm[25] , \imm[24] , \imm[23] , \imm[22] 
		, \imm[21] , \imm[20] , \imm[19] , \imm[18] , \imm[17] , \imm[16] 
		, \imm[15] , \imm[14] , \imm[13] , \imm[12] , \imm[11] , \imm[10] 
		, \imm[9] , \imm[8] , \imm[7] , \imm[6] , \imm[5] , \imm[4] , \imm[3] 
		, \imm[2] , \imm[1] , \imm[0] }), .to_acu(deco2acu), .operand_size
		(opz), .reps(reps), .over_seg({\over_seg[5] , UNCONNECTED_155, 
		UNCONNECTED_156, UNCONNECTED_157, UNCONNECTED_158, 
		UNCONNECTED_159}), .term(term), .start(st));
endmodule
module AWDP_ADD_12(O0, addrshft, useq_ptr);
    output [6:0] O0;
    input [5:0] addrshft;
    input [3:0] useq_ptr;
    // Line 58
    wire [6:0] O0;
    // Line 81
    wire [6:0] N874;

    // Line 58
    assign O0 = N874;
    // Line 81
    assign N874 = useq_ptr + addrshft;
endmodule

module AWDP_ADD_2(O0, addr);

	output [31:0] O0;
	input [31:0] addr;

	wire \addr[4] ;
	wire \addr[5] ;
	wire \addr[6] ;
	wire \addr[7] ;
	wire \addr[8] ;
	wire \addr[9] ;
	wire \addr[10] ;
	wire \addr[11] ;
	wire \addr[12] ;
	wire \addr[13] ;
	wire \addr[14] ;
	wire \addr[15] ;
	wire \addr[16] ;
	wire \addr[17] ;
	wire \addr[18] ;
	wire \addr[19] ;
	wire \addr[20] ;
	wire \addr[21] ;
	wire \addr[22] ;
	wire \addr[23] ;
	wire \addr[24] ;
	wire \addr[25] ;
	wire \addr[26] ;
	wire \addr[27] ;
	wire \addr[28] ;
	wire \addr[29] ;
	wire \addr[30] ;
	wire \addr[31] ;


	assign O0[0] = addr[0];
	assign O0[1] = addr[1];
	assign O0[2] = addr[2];
	assign O0[3] = addr[3];
	assign \addr[4]  = addr[4];
	assign \addr[5]  = addr[5];
	assign \addr[6]  = addr[6];
	assign \addr[7]  = addr[7];
	assign \addr[8]  = addr[8];
	assign \addr[9]  = addr[9];
	assign \addr[10]  = addr[10];
	assign \addr[11]  = addr[11];
	assign \addr[12]  = addr[12];
	assign \addr[13]  = addr[13];
	assign \addr[14]  = addr[14];
	assign \addr[15]  = addr[15];
	assign \addr[16]  = addr[16];
	assign \addr[17]  = addr[17];
	assign \addr[18]  = addr[18];
	assign \addr[19]  = addr[19];
	assign \addr[20]  = addr[20];
	assign \addr[21]  = addr[21];
	assign \addr[22]  = addr[22];
	assign \addr[23]  = addr[23];
	assign \addr[24]  = addr[24];
	assign \addr[25]  = addr[25];
	assign \addr[26]  = addr[26];
	assign \addr[27]  = addr[27];
	assign \addr[28]  = addr[28];
	assign \addr[29]  = addr[29];
	assign \addr[30]  = addr[30];
	assign \addr[31]  = addr[31];

	notech_ha2 i_27(.A(\addr[31] ), .B(n_300), .Z(O0[31]));
	notech_ha2 i_26(.A(\addr[30] ), .B(n_298), .Z(O0[30]), .CO(n_300));
	notech_ha2 i_25(.A(\addr[29] ), .B(n_296), .Z(O0[29]), .CO(n_298));
	notech_ha2 i_24(.A(\addr[28] ), .B(n_294), .Z(O0[28]), .CO(n_296));
	notech_ha2 i_23(.A(\addr[27] ), .B(n_292), .Z(O0[27]), .CO(n_294));
	notech_ha2 i_22(.A(\addr[26] ), .B(n_290), .Z(O0[26]), .CO(n_292));
	notech_ha2 i_21(.A(\addr[25] ), .B(n_288), .Z(O0[25]), .CO(n_290));
	notech_ha2 i_20(.A(\addr[24] ), .B(n_286), .Z(O0[24]), .CO(n_288));
	notech_ha2 i_19(.A(\addr[23] ), .B(n_284), .Z(O0[23]), .CO(n_286));
	notech_ha2 i_18(.A(\addr[22] ), .B(n_282), .Z(O0[22]), .CO(n_284));
	notech_ha2 i_17(.A(\addr[21] ), .B(n_280), .Z(O0[21]), .CO(n_282));
	notech_ha2 i_16(.A(\addr[20] ), .B(n_278), .Z(O0[20]), .CO(n_280));
	notech_ha2 i_15(.A(\addr[19] ), .B(n_276), .Z(O0[19]), .CO(n_278));
	notech_ha2 i_14(.A(\addr[18] ), .B(n_274), .Z(O0[18]), .CO(n_276));
	notech_ha2 i_13(.A(\addr[17] ), .B(n_272), .Z(O0[17]), .CO(n_274));
	notech_ha2 i_12(.A(\addr[16] ), .B(n_270), .Z(O0[16]), .CO(n_272));
	notech_ha2 i_11(.A(\addr[15] ), .B(n_268), .Z(O0[15]), .CO(n_270));
	notech_ha2 i_10(.A(\addr[14] ), .B(n_266), .Z(O0[14]), .CO(n_268));
	notech_ha2 i_9(.A(\addr[13] ), .B(n_264), .Z(O0[13]), .CO(n_266));
	notech_ha2 i_8(.A(\addr[12] ), .B(n_262), .Z(O0[12]), .CO(n_264));
	notech_ha2 i_7(.A(\addr[11] ), .B(n_260), .Z(O0[11]), .CO(n_262));
	notech_ha2 i_6(.A(\addr[10] ), .B(n_258), .Z(O0[10]), .CO(n_260));
	notech_ha2 i_5(.A(\addr[9] ), .B(n_256), .Z(O0[9]), .CO(n_258));
	notech_ha2 i_4(.A(\addr[8] ), .B(n_254), .Z(O0[8]), .CO(n_256));
	notech_ha2 i_3(.A(\addr[7] ), .B(n_252), .Z(O0[7]), .CO(n_254));
	notech_ha2 i_2(.A(\addr[6] ), .B(n_250), .Z(O0[6]), .CO(n_252));
	notech_ha2 i_1(.A(\addr[5] ), .B(\addr[4] ), .Z(O0[5]), .CO(n_250));
	notech_inv i_0(.A(\addr[4] ), .Z(O0[4]));
endmodule
module AWDP_EQ_46(O0, addr, addrf);
    output [0:0] O0;
    input [31:0] addr;
    input [31:0] addrf;
    // Line 85
    wire [0:0] N900;
    // Line 58
    wire [0:0] O0;

    // Line 85
    assign N900 = addr == addrf;
    // Line 58
    assign O0 = N900;
endmodule

module AWDP_EQ_715217(O0, tagA, addr);
    output [0:0] O0;
    input [17:0] tagA;
    input [31:14] addr;
    // Line 128
    wire [0:0] N907;
    // Line 128
    wire [0:0] O0;

    // Line 128
    assign N907 = tagA == addr;
    // Line 128
    assign O0 = N907;
endmodule

module AWDP_INC_1(O0, purge_cnt);

	output [10:0] O0;
	input [10:0] purge_cnt;




	notech_ha2 i_10(.A(purge_cnt[10]), .B(n_106), .Z(O0[10]));
	notech_ha2 i_9(.A(purge_cnt[9]), .B(n_104), .Z(O0[9]), .CO(n_106));
	notech_ha2 i_8(.A(purge_cnt[8]), .B(n_102), .Z(O0[8]), .CO(n_104));
	notech_ha2 i_7(.A(purge_cnt[7]), .B(n_100), .Z(O0[7]), .CO(n_102));
	notech_ha2 i_6(.A(purge_cnt[6]), .B(n_98), .Z(O0[6]), .CO(n_100));
	notech_ha2 i_5(.A(purge_cnt[5]), .B(n_96), .Z(O0[5]), .CO(n_98));
	notech_ha2 i_4(.A(purge_cnt[4]), .B(n_94), .Z(O0[4]), .CO(n_96));
	notech_ha2 i_3(.A(purge_cnt[3]), .B(n_92), .Z(O0[3]), .CO(n_94));
	notech_ha2 i_2(.A(purge_cnt[2]), .B(n_90), .Z(O0[2]), .CO(n_92));
	notech_ha2 i_1(.A(purge_cnt[1]), .B(purge_cnt[0]), .Z(O0[1]), .CO(n_90)
		);
	notech_inv i_0(.A(purge_cnt[0]), .Z(O0[0]));
endmodule
module useq(iaddr, idata, code_req, code_ack, clk, rstn, useq_ptr, squeue, pc_in
		, pc_req, cs, pg_en, pg_fault, pc_pg_fault, valid_len, busy_ram
		);

	output [31:0] iaddr;
	input [127:0] idata;
	output code_req;
	input code_ack;
	input clk;
	input rstn;
	input [3:0] useq_ptr;
	output [127:0] squeue;
	input [31:0] pc_in;
	input pc_req;
	input [31:0] cs;
	input pg_en;
	input pg_fault;
	output pc_pg_fault;
	output [5:0] valid_len;
	input busy_ram;

	wire [1:0] wptr;
	wire [255:0] queue;
	wire [1:0] fault_wptr;
	wire [3:0] tagV;
	wire [17:0] tagA;
	wire [31:0] addr_0;
	wire [9:0] cacheA;
	wire [149:0] cacheD;
	wire [6:0] nbus_12105;
	wire [5:0] addrshft;
	wire [10:0] purge_cnt;
	wire [31:0] addrf;

	supply0 AMBIT_GND;
	supply1 AMBIT_VDD;


	notech_inv i_16042(.A(n_62374), .Z(n_62375));
	notech_inv i_16041(.A(n_62325), .Z(n_62374));
	notech_inv i_16000(.A(n_62332), .Z(n_62333));
	notech_inv i_15999(.A(n_62257), .Z(n_62332));
	notech_inv i_15998(.A(n_62330), .Z(n_62331));
	notech_inv i_15997(.A(n_62251), .Z(n_62330));
	notech_inv i_15996(.A(n_62328), .Z(n_62329));
	notech_inv i_15995(.A(n_62247), .Z(n_62328));
	notech_inv i_15994(.A(n_62326), .Z(n_62327));
	notech_inv i_15993(.A(n_62245), .Z(n_62326));
	notech_inv i_15992(.A(n_62324), .Z(n_62325));
	notech_inv i_15991(.A(n_62327), .Z(n_62324));
	notech_inv i_15928(.A(n_62260), .Z(n_62261));
	notech_inv i_15927(.A(n_62185), .Z(n_62260));
	notech_inv i_15926(.A(n_62258), .Z(n_62259));
	notech_inv i_15925(.A(n_62183), .Z(n_62258));
	notech_inv i_15924(.A(n_62256), .Z(n_62257));
	notech_inv i_15923(.A(n_62259), .Z(n_62256));
	notech_inv i_15922(.A(n_62254), .Z(n_62255));
	notech_inv i_15921(.A(n_62179), .Z(n_62254));
	notech_inv i_15920(.A(n_62252), .Z(n_62253));
	notech_inv i_15919(.A(n_62177), .Z(n_62252));
	notech_inv i_15918(.A(n_62250), .Z(n_62251));
	notech_inv i_15917(.A(n_62253), .Z(n_62250));
	notech_inv i_15916(.A(n_62248), .Z(n_62249));
	notech_inv i_15915(.A(n_62175), .Z(n_62248));
	notech_inv i_15914(.A(n_62246), .Z(n_62247));
	notech_inv i_15913(.A(n_62249), .Z(n_62246));
	notech_inv i_15912(.A(n_62244), .Z(n_62245));
	notech_inv i_15911(.A(n_62329), .Z(n_62244));
	notech_inv i_15854(.A(n_62186), .Z(n_62187));
	notech_inv i_15853(.A(clk), .Z(n_62186));
	notech_inv i_15852(.A(n_62184), .Z(n_62185));
	notech_inv i_15851(.A(n_62187), .Z(n_62184));
	notech_inv i_15850(.A(n_62182), .Z(n_62183));
	notech_inv i_15849(.A(n_62261), .Z(n_62182));
	notech_inv i_15848(.A(n_62180), .Z(n_62181));
	notech_inv i_15847(.A(n_62087), .Z(n_62180));
	notech_inv i_15846(.A(n_62178), .Z(n_62179));
	notech_inv i_15845(.A(n_62181), .Z(n_62178));
	notech_inv i_15844(.A(n_62176), .Z(n_62177));
	notech_inv i_15843(.A(n_62255), .Z(n_62176));
	notech_inv i_15842(.A(n_62174), .Z(n_62175));
	notech_inv i_15841(.A(n_62331), .Z(n_62174));
	notech_inv i_15753(.A(n_62086), .Z(n_62087));
	notech_inv i_15752(.A(n_62333), .Z(n_62086));
	notech_inv i_15221(.A(n_61542), .Z(n_61558));
	notech_inv i_15219(.A(n_61542), .Z(n_61556));
	notech_inv i_15218(.A(n_61542), .Z(n_61555));
	notech_inv i_15214(.A(n_61542), .Z(n_61551));
	notech_inv i_15212(.A(n_61542), .Z(n_61549));
	notech_inv i_15209(.A(n_61542), .Z(n_61546));
	notech_inv i_15207(.A(n_61542), .Z(n_61544));
	notech_inv i_15206(.A(n_61542), .Z(code_req));
	notech_inv i_15205(.A(n_61560), .Z(n_61542));
	notech_inv i_14353(.A(n_60972), .Z(n_60995));
	notech_inv i_14352(.A(n_60972), .Z(n_60994));
	notech_inv i_14351(.A(n_60972), .Z(n_60993));
	notech_inv i_14350(.A(n_60972), .Z(n_60992));
	notech_inv i_14349(.A(n_60972), .Z(n_60991));
	notech_inv i_14347(.A(n_60972), .Z(n_60989));
	notech_inv i_14346(.A(n_60972), .Z(n_60988));
	notech_inv i_14345(.A(n_60972), .Z(n_60987));
	notech_inv i_14344(.A(n_60972), .Z(n_60986));
	notech_inv i_14343(.A(n_60972), .Z(n_60985));
	notech_inv i_14341(.A(n_60972), .Z(n_60983));
	notech_inv i_14340(.A(n_60972), .Z(n_60982));
	notech_inv i_14339(.A(n_60972), .Z(n_60981));
	notech_inv i_14338(.A(n_60972), .Z(n_60980));
	notech_inv i_14337(.A(n_60972), .Z(n_60979));
	notech_inv i_14335(.A(n_60972), .Z(n_60977));
	notech_inv i_14334(.A(n_60972), .Z(n_60976));
	notech_inv i_14333(.A(n_60972), .Z(n_60975));
	notech_inv i_14332(.A(n_60972), .Z(n_60974));
	notech_inv i_14331(.A(n_60972), .Z(n_60973));
	notech_inv i_14330(.A(rstn), .Z(n_60972));
	notech_inv i_14329(.A(n_60966), .Z(n_60971));
	notech_inv i_14328(.A(n_60966), .Z(n_60970));
	notech_inv i_14327(.A(n_60966), .Z(n_60969));
	notech_inv i_14326(.A(n_60966), .Z(n_60968));
	notech_inv i_14325(.A(n_60966), .Z(n_60967));
	notech_inv i_14324(.A(rstn), .Z(n_60966));
	notech_inv i_13797(.A(n_60395), .Z(n_60400));
	notech_inv i_13793(.A(n_60395), .Z(n_60396));
	notech_inv i_13792(.A(pc_req), .Z(n_60395));
	notech_inv i_13778(.A(n_60270), .Z(n_60286));
	notech_inv i_13776(.A(n_60270), .Z(n_60284));
	notech_inv i_13775(.A(n_60270), .Z(n_60283));
	notech_inv i_13771(.A(n_60270), .Z(n_60279));
	notech_inv i_13769(.A(n_60270), .Z(n_60277));
	notech_inv i_13766(.A(n_60270), .Z(n_60274));
	notech_inv i_13764(.A(n_60270), .Z(n_60272));
	notech_inv i_13763(.A(n_60270), .Z(n_60271));
	notech_inv i_13762(.A(wptr[1]), .Z(n_60270));
	notech_inv i_13755(.A(n_60257), .Z(n_60262));
	notech_inv i_13751(.A(n_60257), .Z(n_60258));
	notech_inv i_13750(.A(n_3078), .Z(n_60257));
	notech_inv i_13748(.A(n_60238), .Z(n_60254));
	notech_inv i_13746(.A(n_60238), .Z(n_60252));
	notech_inv i_13745(.A(n_60238), .Z(n_60251));
	notech_inv i_13741(.A(n_60238), .Z(n_60247));
	notech_inv i_13739(.A(n_60238), .Z(n_60245));
	notech_inv i_13737(.A(n_60238), .Z(n_60243));
	notech_inv i_13735(.A(n_60238), .Z(n_60241));
	notech_inv i_13733(.A(n_60238), .Z(n_60239));
	notech_inv i_13732(.A(n_142753060), .Z(n_60238));
	notech_inv i_13725(.A(n_60229), .Z(n_60230));
	notech_inv i_13724(.A(n_141853051), .Z(n_60229));
	notech_inv i_13720(.A(n_60229), .Z(n_60225));
	notech_inv i_13716(.A(n_60229), .Z(n_60221));
	notech_inv i_13711(.A(n_60229), .Z(n_60216));
	notech_inv i_13707(.A(n_60229), .Z(n_60212));
	notech_inv i_13697(.A(n_60201), .Z(n_60202));
	notech_inv i_13696(.A(n_60182), .Z(n_60201));
	notech_inv i_13692(.A(n_60201), .Z(n_60197));
	notech_inv i_13688(.A(n_60201), .Z(n_60193));
	notech_inv i_13683(.A(n_60201), .Z(n_60188));
	notech_inv i_13679(.A(n_60201), .Z(n_60184));
	notech_inv i_13677(.A(n_60229), .Z(n_60182));
	notech_inv i_13669(.A(n_60173), .Z(n_60174));
	notech_inv i_13668(.A(n_60154), .Z(n_60173));
	notech_inv i_13664(.A(n_60173), .Z(n_60169));
	notech_inv i_13660(.A(n_60173), .Z(n_60165));
	notech_inv i_13655(.A(n_60173), .Z(n_60160));
	notech_inv i_13651(.A(n_60173), .Z(n_60156));
	notech_inv i_13649(.A(n_60229), .Z(n_60154));
	notech_inv i_13639(.A(n_60142), .Z(n_60143));
	notech_inv i_13638(.A(\nbus_12117[0] ), .Z(n_60142));
	notech_inv i_13516(.A(n_60243), .Z(n_60010));
	notech_inv i_13514(.A(n_60243), .Z(n_60008));
	notech_inv i_13513(.A(n_60243), .Z(n_60007));
	notech_inv i_13509(.A(n_60243), .Z(n_60003));
	notech_inv i_13507(.A(n_60243), .Z(n_60001));
	notech_inv i_13504(.A(n_60243), .Z(n_59998));
	notech_inv i_13502(.A(n_60243), .Z(n_59996));
	notech_inv i_13501(.A(n_60243), .Z(n_59995));
	notech_inv i_11877(.A(n_58374), .Z(n_58379));
	notech_inv i_11873(.A(n_58374), .Z(n_58375));
	notech_inv i_11872(.A(n_3074), .Z(n_58374));
	notech_inv i_11870(.A(n_58358), .Z(n_58371));
	notech_inv i_11868(.A(n_58358), .Z(n_58369));
	notech_inv i_11864(.A(n_58358), .Z(n_58365));
	notech_inv i_11858(.A(n_58358), .Z(n_58359));
	notech_inv i_11857(.A(n_1304), .Z(n_58358));
	notech_inv i_11855(.A(n_58342), .Z(n_58355));
	notech_inv i_11853(.A(n_58342), .Z(n_58353));
	notech_inv i_11849(.A(n_58342), .Z(n_58349));
	notech_inv i_11843(.A(n_58342), .Z(n_58343));
	notech_inv i_11842(.A(n_1305), .Z(n_58342));
	notech_inv i_11840(.A(n_58326), .Z(n_58339));
	notech_inv i_11838(.A(n_58326), .Z(n_58337));
	notech_inv i_11834(.A(n_58326), .Z(n_58333));
	notech_inv i_11828(.A(n_58326), .Z(n_58327));
	notech_inv i_11827(.A(n_1296), .Z(n_58326));
	notech_inv i_11825(.A(n_58310), .Z(n_58323));
	notech_inv i_11823(.A(n_58310), .Z(n_58321));
	notech_inv i_11819(.A(n_58310), .Z(n_58317));
	notech_inv i_11813(.A(n_58310), .Z(n_58311));
	notech_inv i_11812(.A(n_1297), .Z(n_58310));
	notech_inv i_11810(.A(n_58294), .Z(n_58307));
	notech_inv i_11808(.A(n_58294), .Z(n_58305));
	notech_inv i_11804(.A(n_58294), .Z(n_58301));
	notech_inv i_11798(.A(n_58294), .Z(n_58295));
	notech_inv i_11797(.A(n_1300), .Z(n_58294));
	notech_inv i_11795(.A(n_58278), .Z(n_58291));
	notech_inv i_11793(.A(n_58278), .Z(n_58289));
	notech_inv i_11789(.A(n_58278), .Z(n_58285));
	notech_inv i_11783(.A(n_58278), .Z(n_58279));
	notech_inv i_11782(.A(n_1301), .Z(n_58278));
	notech_inv i_11779(.A(n_58259), .Z(n_58274));
	notech_inv i_11777(.A(n_58259), .Z(n_58272));
	notech_inv i_11772(.A(n_58259), .Z(n_58267));
	notech_inv i_11771(.A(n_58259), .Z(n_58266));
	notech_inv i_11765(.A(n_58259), .Z(n_58260));
	notech_inv i_11764(.A(n_1290), .Z(n_58259));
	notech_inv i_11762(.A(n_58240), .Z(n_58256));
	notech_inv i_11760(.A(n_58240), .Z(n_58254));
	notech_inv i_11759(.A(n_58240), .Z(n_58253));
	notech_inv i_11755(.A(n_58240), .Z(n_58249));
	notech_inv i_11753(.A(n_58240), .Z(n_58247));
	notech_inv i_11750(.A(n_58240), .Z(n_58244));
	notech_inv i_11748(.A(n_58240), .Z(n_58242));
	notech_inv i_11747(.A(n_58240), .Z(n_58241));
	notech_inv i_11746(.A(n_1291), .Z(n_58240));
	notech_inv i_11744(.A(n_58221), .Z(n_58237));
	notech_inv i_11742(.A(n_58221), .Z(n_58235));
	notech_inv i_11741(.A(n_58221), .Z(n_58234));
	notech_inv i_11737(.A(n_58221), .Z(n_58230));
	notech_inv i_11735(.A(n_58221), .Z(n_58228));
	notech_inv i_11732(.A(n_58221), .Z(n_58225));
	notech_inv i_11730(.A(n_58221), .Z(n_58223));
	notech_inv i_11729(.A(n_58221), .Z(n_58222));
	notech_inv i_11728(.A(n_1292), .Z(n_58221));
	notech_inv i_11726(.A(n_58202), .Z(n_58218));
	notech_inv i_11724(.A(n_58202), .Z(n_58216));
	notech_inv i_11723(.A(n_58202), .Z(n_58215));
	notech_inv i_11719(.A(n_58202), .Z(n_58211));
	notech_inv i_11717(.A(n_58202), .Z(n_58209));
	notech_inv i_11714(.A(n_58202), .Z(n_58206));
	notech_inv i_11712(.A(n_58202), .Z(n_58204));
	notech_inv i_11711(.A(n_58202), .Z(n_58203));
	notech_inv i_11710(.A(n_1982), .Z(n_58202));
	notech_inv i_11703(.A(n_58189), .Z(n_58194));
	notech_inv i_11699(.A(n_58189), .Z(n_58190));
	notech_inv i_11698(.A(n_1999), .Z(n_58189));
	notech_inv i_11691(.A(n_58176), .Z(n_58181));
	notech_inv i_11687(.A(n_58176), .Z(n_58177));
	notech_inv i_11686(.A(n_1998), .Z(n_58176));
	notech_inv i_11679(.A(n_58163), .Z(n_58168));
	notech_inv i_11675(.A(n_58163), .Z(n_58164));
	notech_inv i_11674(.A(n_1996), .Z(n_58163));
	notech_inv i_11667(.A(n_58150), .Z(n_58155));
	notech_inv i_11663(.A(n_58150), .Z(n_58151));
	notech_inv i_11662(.A(n_1995), .Z(n_58150));
	notech_inv i_11655(.A(n_58137), .Z(n_58142));
	notech_inv i_11651(.A(n_58137), .Z(n_58138));
	notech_inv i_11650(.A(n_1979), .Z(n_58137));
	notech_inv i_11643(.A(n_58124), .Z(n_58129));
	notech_inv i_11639(.A(n_58124), .Z(n_58125));
	notech_inv i_11638(.A(n_1978), .Z(n_58124));
	notech_inv i_11631(.A(n_58111), .Z(n_58116));
	notech_inv i_11627(.A(n_58111), .Z(n_58112));
	notech_inv i_11626(.A(n_1984), .Z(n_58111));
	notech_inv i_11619(.A(n_58098), .Z(n_58103));
	notech_inv i_11615(.A(n_58098), .Z(n_58099));
	notech_inv i_11614(.A(n_1983), .Z(n_58098));
	notech_inv i_11607(.A(n_58085), .Z(n_58090));
	notech_inv i_11603(.A(n_58085), .Z(n_58086));
	notech_inv i_11602(.A(n_1991), .Z(n_58085));
	notech_inv i_11595(.A(n_58072), .Z(n_58077));
	notech_inv i_11591(.A(n_58072), .Z(n_58073));
	notech_inv i_11590(.A(n_1990), .Z(n_58072));
	notech_inv i_11583(.A(n_58059), .Z(n_58064));
	notech_inv i_11579(.A(n_58059), .Z(n_58060));
	notech_inv i_11578(.A(n_1988), .Z(n_58059));
	notech_inv i_11571(.A(n_58046), .Z(n_58051));
	notech_inv i_11567(.A(n_58046), .Z(n_58047));
	notech_inv i_11566(.A(n_1987), .Z(n_58046));
	notech_inv i_11564(.A(n_58030), .Z(n_58043));
	notech_inv i_11562(.A(n_58030), .Z(n_58041));
	notech_inv i_11558(.A(n_58030), .Z(n_58037));
	notech_inv i_11552(.A(n_58030), .Z(n_58031));
	notech_inv i_11551(.A(n_1318), .Z(n_58030));
	notech_inv i_11549(.A(n_58014), .Z(n_58027));
	notech_inv i_11547(.A(n_58014), .Z(n_58025));
	notech_inv i_11543(.A(n_58014), .Z(n_58021));
	notech_inv i_11537(.A(n_58014), .Z(n_58015));
	notech_inv i_11536(.A(n_1321), .Z(n_58014));
	notech_inv i_11534(.A(n_57998), .Z(n_58011));
	notech_inv i_11532(.A(n_57998), .Z(n_58009));
	notech_inv i_11528(.A(n_57998), .Z(n_58005));
	notech_inv i_11522(.A(n_57998), .Z(n_57999));
	notech_inv i_11521(.A(n_1310), .Z(n_57998));
	notech_inv i_11519(.A(n_57982), .Z(n_57995));
	notech_inv i_11517(.A(n_57982), .Z(n_57993));
	notech_inv i_11513(.A(n_57982), .Z(n_57989));
	notech_inv i_11507(.A(n_57982), .Z(n_57983));
	notech_inv i_11506(.A(n_1311), .Z(n_57982));
	notech_inv i_11504(.A(n_57966), .Z(n_57979));
	notech_inv i_11502(.A(n_57966), .Z(n_57977));
	notech_inv i_11498(.A(n_57966), .Z(n_57973));
	notech_inv i_11492(.A(n_57966), .Z(n_57967));
	notech_inv i_11491(.A(n_1314), .Z(n_57966));
	notech_inv i_11489(.A(n_57950), .Z(n_57963));
	notech_inv i_11487(.A(n_57950), .Z(n_57961));
	notech_inv i_11483(.A(n_57950), .Z(n_57957));
	notech_inv i_11477(.A(n_57950), .Z(n_57951));
	notech_inv i_11476(.A(n_1315), .Z(n_57950));
	notech_inv i_11474(.A(n_57929), .Z(n_57947));
	notech_inv i_11472(.A(n_57929), .Z(n_57945));
	notech_inv i_11469(.A(n_57929), .Z(n_57942));
	notech_inv i_11467(.A(n_57929), .Z(n_57940));
	notech_inv i_11464(.A(n_57929), .Z(n_57937));
	notech_inv i_11462(.A(n_57929), .Z(n_57935));
	notech_inv i_11459(.A(n_57929), .Z(n_57932));
	notech_inv i_11457(.A(n_57929), .Z(n_57930));
	notech_inv i_11456(.A(n_3073), .Z(n_57929));
	notech_inv i_8422(.A(\nbus_12116[0] ), .Z(n_54331));
	notech_inv i_8420(.A(\nbus_12116[0] ), .Z(n_54329));
	notech_inv i_8417(.A(\nbus_12116[0] ), .Z(n_54326));
	notech_inv i_8415(.A(\nbus_12116[0] ), .Z(n_54324));
	notech_inv i_8412(.A(\nbus_12116[0] ), .Z(n_54321));
	notech_inv i_8410(.A(\nbus_12116[0] ), .Z(n_54319));
	notech_inv i_8407(.A(\nbus_12116[0] ), .Z(n_54316));
	notech_inv i_8405(.A(\nbus_12116[0] ), .Z(n_54314));
	notech_inv i_8402(.A(\nbus_12116[128] ), .Z(n_54310));
	notech_inv i_8400(.A(\nbus_12116[128] ), .Z(n_54308));
	notech_inv i_8397(.A(\nbus_12116[128] ), .Z(n_54305));
	notech_inv i_8395(.A(\nbus_12116[128] ), .Z(n_54303));
	notech_inv i_8392(.A(\nbus_12116[128] ), .Z(n_54300));
	notech_inv i_8390(.A(\nbus_12116[128] ), .Z(n_54298));
	notech_inv i_8387(.A(\nbus_12116[128] ), .Z(n_54295));
	notech_inv i_8385(.A(\nbus_12116[128] ), .Z(n_54293));
	notech_inv i_8382(.A(n_54271), .Z(n_54289));
	notech_inv i_8380(.A(n_54271), .Z(n_54287));
	notech_inv i_8377(.A(n_54271), .Z(n_54284));
	notech_inv i_8375(.A(n_54271), .Z(n_54282));
	notech_inv i_8372(.A(n_54271), .Z(n_54279));
	notech_inv i_8370(.A(n_54271), .Z(n_54277));
	notech_inv i_8367(.A(n_54271), .Z(n_54274));
	notech_inv i_8365(.A(n_54271), .Z(n_54272));
	notech_inv i_8364(.A(n_49596963), .Z(n_54271));
	notech_and4 i_129277399(.A(n_2535), .B(n_2537), .C(n_2539), .D(n_1778), 
		.Z(n_2540));
	notech_ao4 i_128377408(.A(n_1988), .B(n_42252), .C(n_1987), .D(n_42268),
		 .Z(n_2541));
	notech_ao4 i_128477407(.A(n_1991), .B(n_42276), .C(n_1990), .D(n_42260),
		 .Z(n_2542));
	notech_and3 i_129077401(.A(n_2542), .B(n_2541), .C(n_1791), .Z(n_2544)
		);
	notech_ao4 i_128777404(.A(n_1996), .B(n_42297), .C(n_1995), .D(n_42361),
		 .Z(n_2545));
	notech_ao4 i_128877403(.A(n_1999), .B(n_42329), .C(n_1998), .D(n_42313),
		 .Z(n_2546));
	notech_ao4 i_131177380(.A(n_58253), .B(n_42221), .C(n_58234), .D(n_42229
		), .Z(n_2549));
	notech_ao4 i_131377378(.A(n_1979), .B(n_42237), .C(n_1978), .D(n_42245),
		 .Z(n_2551));
	notech_ao4 i_132077371(.A(n_1984), .B(n_42285), .C(n_1983), .D(n_42347),
		 .Z(n_2553));
	notech_and4 i_132377368(.A(n_2549), .B(n_2551), .C(n_2553), .D(n_1794), 
		.Z(n_2554));
	notech_ao4 i_131477377(.A(n_1988), .B(n_42253), .C(n_1987), .D(n_42269),
		 .Z(n_2555));
	notech_ao4 i_131577376(.A(n_1991), .B(n_42277), .C(n_1990), .D(n_42261),
		 .Z(n_2556));
	notech_and3 i_132177370(.A(n_2556), .B(n_2555), .C(n_1807), .Z(n_2558)
		);
	notech_ao4 i_131877373(.A(n_1996), .B(n_42299), .C(n_1995), .D(n_42363),
		 .Z(n_2559));
	notech_ao4 i_131977372(.A(n_1999), .B(n_42331), .C(n_1998), .D(n_42315),
		 .Z(n_2560));
	notech_ao4 i_134277349(.A(n_58253), .B(n_42222), .C(n_58234), .D(n_42230
		), .Z(n_2563));
	notech_ao4 i_134477347(.A(n_1979), .B(n_42238), .C(n_1978), .D(n_42246),
		 .Z(n_2565));
	notech_ao4 i_135177340(.A(n_1984), .B(n_42286), .C(n_1983), .D(n_42349),
		 .Z(n_2567));
	notech_and4 i_135477337(.A(n_2563), .B(n_2565), .C(n_2567), .D(n_1810), 
		.Z(n_2568));
	notech_ao4 i_134577346(.A(n_58064), .B(n_42254), .C(n_58051), .D(n_42270
		), .Z(n_2569));
	notech_ao4 i_134677345(.A(n_58090), .B(n_42278), .C(n_58077), .D(n_42262
		), .Z(n_2570));
	notech_and3 i_135277339(.A(n_2570), .B(n_2569), .C(n_1823), .Z(n_2572)
		);
	notech_ao4 i_134977342(.A(n_58168), .B(n_42301), .C(n_58155), .D(n_42365
		), .Z(n_2573));
	notech_ao4 i_135077341(.A(n_58194), .B(n_42333), .C(n_58181), .D(n_42317
		), .Z(n_2574));
	notech_ao4 i_137377318(.A(n_58253), .B(n_42223), .C(n_58234), .D(n_42231
		), .Z(n_2577));
	notech_ao4 i_137577316(.A(n_58142), .B(n_42239), .C(n_58129), .D(n_42247
		), .Z(n_2579));
	notech_ao4 i_138277309(.A(n_58116), .B(n_42287), .C(n_58103), .D(n_42351
		), .Z(n_2581));
	notech_and4 i_138577306(.A(n_2577), .B(n_2579), .C(n_2581), .D(n_1826), 
		.Z(n_2582));
	notech_ao4 i_137677315(.A(n_1988), .B(n_42255), .C(n_1987), .D(n_42271),
		 .Z(n_2583));
	notech_ao4 i_137777314(.A(n_1991), .B(n_42279), .C(n_1990), .D(n_42263),
		 .Z(n_2584));
	notech_and3 i_138377308(.A(n_2584), .B(n_2583), .C(n_1839), .Z(n_2586)
		);
	notech_ao4 i_138077311(.A(n_1996), .B(n_42303), .C(n_1995), .D(n_42367),
		 .Z(n_2587));
	notech_ao4 i_138177310(.A(n_1999), .B(n_42335), .C(n_1998), .D(n_42319),
		 .Z(n_2588));
	notech_ao4 i_140477287(.A(n_58253), .B(n_42224), .C(n_58234), .D(n_42232
		), .Z(n_2591));
	notech_ao4 i_140677285(.A(n_1979), .B(n_42240), .C(n_1978), .D(n_42248),
		 .Z(n_2593));
	notech_ao4 i_141377278(.A(n_1984), .B(n_42288), .C(n_1983), .D(n_42353),
		 .Z(n_2595));
	notech_and4 i_141677275(.A(n_2591), .B(n_2593), .C(n_2595), .D(n_1842), 
		.Z(n_2596));
	notech_ao4 i_140777284(.A(n_1988), .B(n_42256), .C(n_1987), .D(n_42272),
		 .Z(n_2597));
	notech_ao4 i_140877283(.A(n_1991), .B(n_42280), .C(n_1990), .D(n_42264),
		 .Z(n_2598));
	notech_and3 i_141477277(.A(n_2598), .B(n_2597), .C(n_1855), .Z(n_2600)
		);
	notech_ao4 i_141177280(.A(n_1996), .B(n_42305), .C(n_1995), .D(n_42369),
		 .Z(n_2601));
	notech_ao4 i_141277279(.A(n_1999), .B(n_42337), .C(n_1998), .D(n_42321),
		 .Z(n_2602));
	notech_ao4 i_143577256(.A(n_58234), .B(n_42233), .C(n_58272), .D(n_42217
		), .Z(n_2605));
	notech_ao4 i_143777254(.A(n_1979), .B(n_42241), .C(n_1978), .D(n_42249),
		 .Z(n_2607));
	notech_ao4 i_144477247(.A(n_1984), .B(n_42291), .C(n_1983), .D(n_42355),
		 .Z(n_2609));
	notech_and4 i_144777244(.A(n_2605), .B(n_2607), .C(n_2609), .D(n_1858), 
		.Z(n_2610));
	notech_ao4 i_143877253(.A(n_1988), .B(n_42257), .C(n_1987), .D(n_42273),
		 .Z(n_2611));
	notech_ao4 i_143977252(.A(n_1991), .B(n_42281), .C(n_1990), .D(n_42265),
		 .Z(n_2612));
	notech_and3 i_144577246(.A(n_2612), .B(n_2611), .C(n_1871), .Z(n_2614)
		);
	notech_ao4 i_144277249(.A(n_1996), .B(n_42307), .C(n_1995), .D(n_42371),
		 .Z(n_2615));
	notech_ao4 i_144377248(.A(n_1999), .B(n_42339), .C(n_1998), .D(n_42323),
		 .Z(n_2616));
	notech_ao4 i_146677225(.A(n_58253), .B(n_42226), .C(n_58234), .D(n_42234
		), .Z(n_2619));
	notech_ao4 i_146877223(.A(n_1979), .B(n_42242), .C(n_1978), .D(n_42250),
		 .Z(n_2621));
	notech_ao4 i_147577216(.A(n_1984), .B(n_42293), .C(n_1983), .D(n_42357),
		 .Z(n_2623));
	notech_and4 i_147877213(.A(n_2619), .B(n_2621), .C(n_2623), .D(n_1874), 
		.Z(n_2624));
	notech_ao4 i_146977222(.A(n_58064), .B(n_42258), .C(n_58051), .D(n_42274
		), .Z(n_2625));
	notech_ao4 i_147077221(.A(n_58090), .B(n_42282), .C(n_58077), .D(n_42266
		), .Z(n_2626));
	notech_and3 i_147677215(.A(n_2626), .B(n_2625), .C(n_1887), .Z(n_2628)
		);
	notech_ao4 i_147377218(.A(n_58168), .B(n_42309), .C(n_58155), .D(n_42373
		), .Z(n_2629));
	notech_ao4 i_147477217(.A(n_58194), .B(n_42341), .C(n_58181), .D(n_42325
		), .Z(n_2630));
	notech_ao4 i_149777194(.A(n_58253), .B(n_42227), .C(n_58234), .D(n_42235
		), .Z(n_2633));
	notech_ao4 i_149977192(.A(n_58142), .B(n_42243), .C(n_58129), .D(n_42251
		), .Z(n_2635));
	notech_ao4 i_150677185(.A(n_58116), .B(n_42295), .C(n_58103), .D(n_42359
		), .Z(n_2637));
	notech_and4 i_150977182(.A(n_2633), .B(n_2635), .C(n_2637), .D(n_1890), 
		.Z(n_2638));
	notech_ao4 i_150077191(.A(n_58064), .B(n_42259), .C(n_58051), .D(n_42275
		), .Z(n_2639));
	notech_ao4 i_150177190(.A(n_58090), .B(n_42283), .C(n_58077), .D(n_42267
		), .Z(n_2640));
	notech_and3 i_150777184(.A(n_2640), .B(n_2639), .C(n_1903), .Z(n_2642)
		);
	notech_ao4 i_150477187(.A(n_58168), .B(n_42311), .C(n_58155), .D(n_42375
		), .Z(n_2643));
	notech_ao4 i_150577186(.A(n_58194), .B(n_42343), .C(n_58181), .D(n_42327
		), .Z(n_2644));
	notech_ao4 i_152877163(.A(n_58253), .B(n_42228), .C(n_58234), .D(n_42236
		), .Z(n_2647));
	notech_ao4 i_153077161(.A(n_58142), .B(n_42244), .C(n_58129), .D(n_42252
		), .Z(n_2649));
	notech_ao4 i_153777154(.A(n_58116), .B(n_42297), .C(n_58103), .D(n_42361
		), .Z(n_2651));
	notech_and4 i_154077151(.A(n_2647), .B(n_2649), .C(n_2651), .D(n_1906), 
		.Z(n_2652));
	notech_ao4 i_153177160(.A(n_58064), .B(n_42260), .C(n_58051), .D(n_42276
		), .Z(n_2653));
	notech_ao4 i_153277159(.A(n_58090), .B(n_42284), .C(n_58077), .D(n_42268
		), .Z(n_2654));
	notech_and3 i_153877153(.A(n_2654), .B(n_2653), .C(n_1919), .Z(n_2656)
		);
	notech_ao4 i_153577156(.A(n_58168), .B(n_42313), .C(n_58155), .D(n_42377
		), .Z(n_2657));
	notech_ao4 i_153677155(.A(n_58194), .B(n_42345), .C(n_58181), .D(n_42329
		), .Z(n_2658));
	notech_ao4 i_155977132(.A(n_58253), .B(n_42229), .C(n_58235), .D(n_42237
		), .Z(n_2661));
	notech_ao4 i_156177130(.A(n_58142), .B(n_42245), .C(n_58129), .D(n_42253
		), .Z(n_2663));
	notech_ao4 i_156877123(.A(n_58116), .B(n_42299), .C(n_58103), .D(n_42363
		), .Z(n_2665));
	notech_and4 i_157177120(.A(n_2661), .B(n_2663), .C(n_2665), .D(n_1922), 
		.Z(n_2666));
	notech_ao4 i_156277129(.A(n_58064), .B(n_42261), .C(n_58051), .D(n_42277
		), .Z(n_2667));
	notech_ao4 i_156377128(.A(n_58090), .B(n_42285), .C(n_58077), .D(n_42269
		), .Z(n_2668));
	notech_and3 i_156977122(.A(n_2668), .B(n_2667), .C(n_1935), .Z(n_2670)
		);
	notech_ao4 i_156677125(.A(n_58168), .B(n_42315), .C(n_58155), .D(n_42379
		), .Z(n_2671));
	notech_ao4 i_156777124(.A(n_58194), .B(n_42347), .C(n_58181), .D(n_42331
		), .Z(n_2672));
	notech_ao4 i_159077101(.A(n_58254), .B(n_42230), .C(n_58235), .D(n_42238
		), .Z(n_2675));
	notech_ao4 i_159277099(.A(n_58142), .B(n_42246), .C(n_58129), .D(n_42254
		), .Z(n_2677));
	notech_ao4 i_159977092(.A(n_58116), .B(n_42301), .C(n_58103), .D(n_42365
		), .Z(n_2679));
	notech_and4 i_160277089(.A(n_2675), .B(n_2677), .C(n_2679), .D(n_1938), 
		.Z(n_2680));
	notech_ao4 i_159377098(.A(n_58064), .B(n_42262), .C(n_58051), .D(n_42278
		), .Z(n_2681));
	notech_ao4 i_159477097(.A(n_58090), .B(n_42286), .C(n_58077), .D(n_42270
		), .Z(n_2682));
	notech_and3 i_160077091(.A(n_2682), .B(n_2681), .C(n_1951), .Z(n_2684)
		);
	notech_ao4 i_159777094(.A(n_58168), .B(n_42317), .C(n_58155), .D(n_42381
		), .Z(n_2685));
	notech_ao4 i_159877093(.A(n_58194), .B(n_42349), .C(n_58181), .D(n_42333
		), .Z(n_2686));
	notech_ao4 i_162177070(.A(n_58254), .B(n_42242), .C(n_58235), .D(n_42250
		), .Z(n_2689));
	notech_ao4 i_162377068(.A(n_58142), .B(n_42258), .C(n_58129), .D(n_42266
		), .Z(n_2691));
	notech_ao4 i_163077061(.A(n_58116), .B(n_42325), .C(n_58103), .D(n_42389
		), .Z(n_2693));
	notech_and4 i_163377058(.A(n_2689), .B(n_2691), .C(n_2693), .D(n_1954), 
		.Z(n_2694));
	notech_ao4 i_162477067(.A(n_58064), .B(n_42274), .C(n_58051), .D(n_42293
		), .Z(n_2695));
	notech_ao4 i_162577066(.A(n_58090), .B(n_42309), .C(n_58077), .D(n_42282
		), .Z(n_2696));
	notech_and3 i_163177060(.A(n_2696), .B(n_2695), .C(n_1967), .Z(n_2698)
		);
	notech_ao4 i_162877063(.A(n_58168), .B(n_42341), .C(n_58155), .D(n_42405
		), .Z(n_2699));
	notech_ao4 i_162977062(.A(n_58194), .B(n_42373), .C(n_58181), .D(n_42357
		), .Z(n_2700));
	notech_ao4 i_214876543(.A(n_60212), .B(n_42629), .C(n_60003), .D(n_42343
		), .Z(n_2703));
	notech_ao4 i_218176510(.A(n_60212), .B(n_42621), .C(n_60003), .D(n_42327
		), .Z(n_2704));
	notech_ao4 i_221376478(.A(n_60212), .B(n_42613), .C(n_60003), .D(n_42311
		), .Z(n_2705));
	notech_ao4 i_224576446(.A(n_60212), .B(n_42605), .C(n_60003), .D(n_42295
		), .Z(n_2706));
	notech_ao4 i_128977402(.A(n_58116), .B(n_42284), .C(n_58103), .D(n_42345
		), .Z(n_2539));
	notech_nand3 i_68(.A(n_57942), .B(n_58215), .C(queue[14]), .Z(n_2707));
	notech_or2 i_69(.A(n_58235), .B(n_42199), .Z(n_2722));
	notech_nand3 i_1524994(.A(n_3096), .B(n_3089), .C(n_2707), .Z(squeue[14]
		));
	notech_nand3 i_99(.A(n_57942), .B(n_58215), .C(queue[29]), .Z(n_2723));
	notech_or2 i_100(.A(n_58234), .B(n_42214), .Z(n_2738));
	notech_nand3 i_3025009(.A(n_3110), .B(n_3103), .C(n_2723), .Z(squeue[29]
		));
	notech_nand3 i_130(.A(n_57942), .B(n_58215), .C(queue[37]), .Z(n_2739)
		);
	notech_or2 i_131(.A(n_58234), .B(n_42222), .Z(n_2754));
	notech_nand3 i_3825017(.A(n_3124), .B(n_3117), .C(n_2739), .Z(squeue[37]
		));
	notech_nand3 i_161(.A(n_57942), .B(n_58215), .C(queue[54]), .Z(n_2755)
		);
	notech_or2 i_162(.A(n_58234), .B(n_42239), .Z(n_2770));
	notech_nand3 i_5525034(.A(n_3138), .B(n_3131), .C(n_2755), .Z(squeue[54]
		));
	notech_nand3 i_378(.A(n_57942), .B(n_58215), .C(queue[61]), .Z(n_2771)
		);
	notech_or2 i_379(.A(n_58234), .B(n_42246), .Z(n_2786));
	notech_nand3 i_6225041(.A(n_3152), .B(n_3145), .C(n_2771), .Z(squeue[61]
		));
	notech_nand3 i_409(.A(n_57942), .B(n_58215), .C(queue[62]), .Z(n_2787)
		);
	notech_or2 i_410(.A(n_58230), .B(n_42247), .Z(n_2802));
	notech_nand3 i_6325042(.A(n_3166), .B(n_3159), .C(n_2787), .Z(squeue[62]
		));
	notech_nand3 i_471(.A(n_57942), .B(n_58215), .C(queue[64]), .Z(n_2803)
		);
	notech_or2 i_472(.A(n_58230), .B(n_42249), .Z(n_2818));
	notech_nand3 i_6525044(.A(n_3180), .B(n_3173), .C(n_2803), .Z(squeue[64]
		));
	notech_nand3 i_595(.A(n_57942), .B(n_58215), .C(queue[69]), .Z(n_2819)
		);
	notech_or2 i_596(.A(n_58230), .B(n_42254), .Z(n_2834));
	notech_nand3 i_7025049(.A(n_3194), .B(n_3187), .C(n_2819), .Z(squeue[69]
		));
	notech_nand3 i_626(.A(n_57942), .B(n_58215), .C(queue[70]), .Z(n_2835)
		);
	notech_or2 i_627(.A(n_58230), .B(n_42255), .Z(n_2850));
	notech_nand3 i_7125050(.A(n_3208), .B(n_3201), .C(n_2835), .Z(squeue[70]
		));
	notech_nand3 i_843(.A(n_57942), .B(n_58215), .C(queue[77]), .Z(n_2851)
		);
	notech_or2 i_844(.A(n_58230), .B(n_42262), .Z(n_2866));
	notech_nand3 i_7825057(.A(n_3222), .B(n_3215), .C(n_2851), .Z(squeue[77]
		));
	notech_nand3 i_874(.A(n_57942), .B(n_58216), .C(queue[78]), .Z(n_2867)
		);
	notech_or2 i_875(.A(n_58230), .B(n_42263), .Z(n_2882));
	notech_nand3 i_7925058(.A(n_3236), .B(n_3229), .C(n_2867), .Z(squeue[78]
		));
	notech_nand3 i_1091(.A(n_57942), .B(n_58216), .C(queue[85]), .Z(n_2883)
		);
	notech_or2 i_1092(.A(n_58230), .B(n_42270), .Z(n_2898));
	notech_nand3 i_8625065(.A(n_3250), .B(n_3243), .C(n_2883), .Z(squeue[85]
		));
	notech_nand3 i_1122(.A(n_57942), .B(n_58215), .C(queue[86]), .Z(n_2899)
		);
	notech_or2 i_1123(.A(n_58230), .B(n_42271), .Z(n_2914));
	notech_nand3 i_8725066(.A(n_3264), .B(n_3257), .C(n_2899), .Z(squeue[86]
		));
	notech_nand3 i_1339(.A(n_57942), .B(n_58215), .C(queue[93]), .Z(n_2915)
		);
	notech_or2 i_1340(.A(n_58234), .B(n_42278), .Z(n_2930));
	notech_nand3 i_9425073(.A(n_3278), .B(n_3271), .C(n_2915), .Z(squeue[93]
		));
	notech_nand3 i_1370(.A(n_57942), .B(n_58215), .C(queue[94]), .Z(n_2931)
		);
	notech_or2 i_1371(.A(n_58234), .B(n_42279), .Z(n_2948));
	notech_nand3 i_9525074(.A(n_3292), .B(n_3285), .C(n_2931), .Z(squeue[94]
		));
	notech_nand3 i_1587(.A(n_57942), .B(n_58215), .C(queue[101]), .Z(n_2949)
		);
	notech_or2 i_1588(.A(n_58234), .B(n_42286), .Z(n_296493405));
	notech_nand3 i_10225081(.A(n_3306), .B(n_3299), .C(n_2949), .Z(squeue[
		101]));
	notech_nand3 i_1618(.A(n_57940), .B(n_58215), .C(queue[102]), .Z(n_2965)
		);
	notech_or2 i_1619(.A(n_58234), .B(n_42287), .Z(n_298096992));
	notech_nand3 i_10325082(.A(n_3320), .B(n_3313), .C(n_2965), .Z(squeue[
		102]));
	notech_nand3 i_1835(.A(n_57940), .B(n_58211), .C(queue[109]), .Z(n_2981)
		);
	notech_or2 i_1836(.A(n_58230), .B(n_42301), .Z(n_2996));
	notech_nand3 i_11025089(.A(n_3334), .B(n_3327), .C(n_2981), .Z(squeue[
		109]));
	notech_nand3 i_1866(.A(n_57940), .B(n_58211), .C(queue[110]), .Z(n_2997)
		);
	notech_or2 i_1867(.A(n_58230), .B(n_42303), .Z(n_3012));
	notech_nand3 i_11125090(.A(n_3348), .B(n_3341), .C(n_2997), .Z(squeue[
		110]));
	notech_nand3 i_2083(.A(n_57940), .B(n_58211), .C(queue[117]), .Z(n_3013)
		);
	notech_or2 i_2084(.A(n_58234), .B(n_42317), .Z(n_3028));
	notech_nand3 i_11825097(.A(n_3362), .B(n_3355), .C(n_3013), .Z(squeue[
		117]));
	notech_nand3 i_2114(.A(n_57940), .B(n_58211), .C(queue[118]), .Z(n_3029)
		);
	notech_or2 i_2115(.A(n_58234), .B(n_42319), .Z(n_3044));
	notech_nand3 i_11925098(.A(n_3376), .B(n_3369), .C(n_3029), .Z(squeue[
		118]));
	notech_nand3 i_2362(.A(n_57940), .B(n_58211), .C(queue[126]), .Z(n_3045)
		);
	notech_or2 i_2363(.A(n_58237), .B(n_42335), .Z(n_3060));
	notech_nand3 i_12725106(.A(n_3390), .B(n_3383), .C(n_3045), .Z(squeue[
		126]));
	notech_and2 i_1(.A(addrshft[1]), .B(n_42549), .Z(n_3061));
	notech_nor2 i_60(.A(addrshft[5]), .B(addrshft[4]), .Z(n_3062));
	notech_and3 i_6(.A(addrshft[0]), .B(n_3062), .C(addrshft[3]), .Z(n_3064)
		);
	notech_nao3 i_1331172(.A(addrshft[1]), .B(n_3064), .C(addrshft[2]), .Z(n_1321
		));
	notech_ao3 i_9(.A(addrshft[3]), .B(n_3062), .C(addrshft[0]), .Z(n_3066)
		);
	notech_nao3 i_1331167(.A(addrshft[1]), .B(n_3066), .C(addrshft[2]), .Z(n_1318
		));
	notech_and2 i_5(.A(addrshft[1]), .B(addrshft[2]), .Z(n_3068));
	notech_nand3 i_1331192(.A(addrshft[1]), .B(addrshft[2]), .C(n_3064), .Z(n_1315
		));
	notech_nand3 i_1331187(.A(addrshft[1]), .B(addrshft[2]), .C(n_3066), .Z(n_1314
		));
	notech_and2 i_7(.A(addrshft[2]), .B(n_42548), .Z(n_3070));
	notech_nao3 i_1331182(.A(addrshft[2]), .B(n_3064), .C(addrshft[1]), .Z(n_1311
		));
	notech_nao3 i_1331177(.A(addrshft[2]), .B(n_3066), .C(addrshft[1]), .Z(n_1310
		));
	notech_and4 i_18(.A(n_58009), .B(n_57993), .C(n_57977), .D(n_57961), .Z(n_3072
		));
	notech_and3 i_5295(.A(n_58041), .B(n_58025), .C(n_3072), .Z(n_3073));
	notech_ao3 i_2(.A(addrshft[0]), .B(n_3062), .C(addrshft[3]), .Z(n_3074)
		);
	notech_nand3 i_1331152(.A(n_3074), .B(addrshft[1]), .C(addrshft[2]), .Z(n_1305
		));
	notech_nand3 i_1331142(.A(n_58379), .B(addrshft[2]), .C(n_42548), .Z(n_1304
		));
	notech_or4 i_10(.A(addrshft[5]), .B(addrshft[4]), .C(addrshft[0]), .D(addrshft
		[3]), .Z(n_3076));
	notech_nao3 i_1331147(.A(addrshft[1]), .B(addrshft[2]), .C(n_3076), .Z(n_1301
		));
	notech_nao3 i_1331137(.A(addrshft[2]), .B(n_42548), .C(n_3076), .Z(n_1300
		));
	notech_and2 i_8(.A(n_42548), .B(n_42549), .Z(n_3078));
	notech_nand2 i_1331162(.A(n_3078), .B(n_3064), .Z(n_1297));
	notech_nand2 i_1331157(.A(n_60262), .B(n_3066), .Z(n_1296));
	notech_and4 i_14(.A(n_58337), .B(n_58321), .C(n_58305), .D(n_58289), .Z(n_3080
		));
	notech_nand3 i_3(.A(n_3074), .B(addrshft[1]), .C(n_42549), .Z(n_1292));
	notech_nao3 i_1331127(.A(addrshft[1]), .B(n_42549), .C(n_3076), .Z(n_1291
		));
	notech_nand3 i_1331122(.A(n_3074), .B(n_42548), .C(n_42549), .Z(n_1290)
		);
	notech_and3 i_5314(.A(n_58272), .B(n_58254), .C(n_58237), .Z(n_3083));
	notech_ao4 i_70(.A(n_58305), .B(n_42207), .C(n_58289), .D(n_42223), .Z(n_3084
		));
	notech_ao4 i_71(.A(n_58254), .B(n_42191), .C(n_57961), .D(n_42303), .Z(n_3086
		));
	notech_ao4 i_72(.A(n_57993), .B(n_42279), .C(n_57977), .D(n_42287), .Z(n_3087
		));
	notech_and4 i_81(.A(n_3087), .B(n_3086), .C(n_3084), .D(n_2722), .Z(n_3089
		));
	notech_ao4 i_73(.A(n_58025), .B(n_42263), .C(n_58009), .D(n_42271), .Z(n_3090
		));
	notech_ao4 i_74(.A(n_58321), .B(n_42247), .C(n_58041), .D(n_42255), .Z(n_3091
		));
	notech_ao4 i_75(.A(n_58353), .B(n_42231), .C(n_58337), .D(n_42239), .Z(n_3093
		));
	notech_ao4 i_76(.A(n_58272), .B(n_42183), .C(n_58369), .D(n_42215), .Z(n_3094
		));
	notech_and4 i_82(.A(n_3094), .B(n_3093), .C(n_3091), .D(n_3090), .Z(n_3096
		));
	notech_ao4 i_101(.A(n_58301), .B(n_42222), .C(n_58285), .D(n_42238), .Z(n_3098
		));
	notech_ao4 i_102(.A(n_58253), .B(n_42206), .C(n_57957), .D(n_42333), .Z(n_3100
		));
	notech_ao4 i_103(.A(n_57989), .B(n_42301), .C(n_57973), .D(n_42317), .Z(n_3101
		));
	notech_and4 i_112(.A(n_3101), .B(n_3100), .C(n_3098), .D(n_2738), .Z(n_3103
		));
	notech_ao4 i_104(.A(n_58021), .B(n_42278), .C(n_58005), .D(n_42286), .Z(n_3104
		));
	notech_ao4 i_105(.A(n_58317), .B(n_42262), .C(n_58037), .D(n_42270), .Z(n_3105
		));
	notech_ao4 i_106(.A(n_58353), .B(n_42246), .C(n_58333), .D(n_42254), .Z(n_3107
		));
	notech_ao4 i_107(.A(n_58272), .B(n_42198), .C(n_58369), .D(n_42230), .Z(n_3108
		));
	notech_and4 i_113(.A(n_3108), .B(n_3107), .C(n_3105), .D(n_3104), .Z(n_3110
		));
	notech_ao4 i_132(.A(n_58305), .B(n_42230), .C(n_58289), .D(n_42246), .Z(n_3112
		));
	notech_ao4 i_133(.A(n_58253), .B(n_42214), .C(n_57961), .D(n_42349), .Z(n_3114
		));
	notech_ao4 i_134(.A(n_57993), .B(n_42317), .C(n_57977), .D(n_42333), .Z(n_3115
		));
	notech_and4 i_143(.A(n_3115), .B(n_3114), .C(n_3112), .D(n_2754), .Z(n_3117
		));
	notech_ao4 i_135(.A(n_58025), .B(n_42286), .C(n_58009), .D(n_42301), .Z(n_3118
		));
	notech_ao4 i_136(.A(n_58321), .B(n_42270), .C(n_58041), .D(n_42278), .Z(n_3119
		));
	notech_ao4 i_137(.A(n_58349), .B(n_42254), .C(n_58337), .D(n_42262), .Z(n_3121
		));
	notech_ao4 i_138(.A(n_58272), .B(n_42206), .C(n_58365), .D(n_42238), .Z(n_3122
		));
	notech_and4 i_144(.A(n_3122), .B(n_3121), .C(n_3119), .D(n_3118), .Z(n_3124
		));
	notech_ao4 i_163(.A(n_58305), .B(n_42247), .C(n_58289), .D(n_42263), .Z(n_3126
		));
	notech_ao4 i_164(.A(n_58253), .B(n_42231), .C(n_57961), .D(n_42383), .Z(n_3128
		));
	notech_ao4 i_165(.A(n_57993), .B(n_42351), .C(n_57977), .D(n_42367), .Z(n_3129
		));
	notech_and4 i_174(.A(n_3129), .B(n_3128), .C(n_3126), .D(n_2770), .Z(n_3131
		));
	notech_ao4 i_166(.A(n_58025), .B(n_42319), .C(n_58009), .D(n_42335), .Z(n_3132
		));
	notech_ao4 i_167(.A(n_58321), .B(n_42287), .C(n_58041), .D(n_42303), .Z(n_3133
		));
	notech_ao4 i_168(.A(n_58353), .B(n_42271), .C(n_58337), .D(n_42279), .Z(n_3135
		));
	notech_ao4 i_169(.A(n_58272), .B(n_42223), .C(n_58369), .D(n_42255), .Z(n_3136
		));
	notech_and4 i_175(.A(n_3136), .B(n_3135), .C(n_3133), .D(n_3132), .Z(n_3138
		));
	notech_ao4 i_380(.A(n_58305), .B(n_42254), .C(n_58289), .D(n_42270), .Z(n_3140
		));
	notech_ao4 i_381(.A(n_58253), .B(n_42238), .C(n_57961), .D(n_42397), .Z(n_3142
		));
	notech_ao4 i_382(.A(n_57993), .B(n_42365), .C(n_57977), .D(n_42381), .Z(n_3143
		));
	notech_and4 i_391(.A(n_3143), .B(n_3142), .C(n_3140), .D(n_2786), .Z(n_3145
		));
	notech_ao4 i_383(.A(n_58025), .B(n_42333), .C(n_58009), .D(n_42349), .Z(n_3146
		));
	notech_ao4 i_384(.A(n_58321), .B(n_42301), .C(n_58041), .D(n_42317), .Z(n_3147
		));
	notech_ao4 i_385(.A(n_58353), .B(n_42278), .C(n_58337), .D(n_42286), .Z(n_3149
		));
	notech_ao4 i_386(.A(n_58272), .B(n_42230), .C(n_58369), .D(n_42262), .Z(n_3150
		));
	notech_and4 i_392(.A(n_3150), .B(n_3149), .C(n_3147), .D(n_3146), .Z(n_3152
		));
	notech_ao4 i_411(.A(n_58305), .B(n_42255), .C(n_58289), .D(n_42271), .Z(n_3154
		));
	notech_ao4 i_412(.A(n_58249), .B(n_42239), .C(n_57961), .D(n_42399), .Z(n_3156
		));
	notech_ao4 i_413(.A(n_57993), .B(n_42367), .C(n_57977), .D(n_42383), .Z(n_3157
		));
	notech_and4 i_422(.A(n_3157), .B(n_3156), .C(n_3154), .D(n_2802), .Z(n_3159
		));
	notech_ao4 i_414(.A(n_58025), .B(n_42335), .C(n_58009), .D(n_42351), .Z(n_3160
		));
	notech_ao4 i_415(.A(n_58321), .B(n_42303), .C(n_58041), .D(n_42319), .Z(n_3161
		));
	notech_ao4 i_416(.A(n_58353), .B(n_42279), .C(n_58337), .D(n_42287), .Z(n_3163
		));
	notech_ao4 i_417(.A(n_58272), .B(n_42231), .C(n_58369), .D(n_42263), .Z(n_3164
		));
	notech_and4 i_423(.A(n_3164), .B(n_3163), .C(n_3161), .D(n_3160), .Z(n_3166
		));
	notech_ao4 i_473(.A(n_58305), .B(n_42257), .C(n_58289), .D(n_42273), .Z(n_3168
		));
	notech_ao4 i_474(.A(n_58249), .B(n_42241), .C(n_57961), .D(n_42403), .Z(n_3170
		));
	notech_ao4 i_475(.A(n_57993), .B(n_42371), .C(n_57977), .D(n_42387), .Z(n_3171
		));
	notech_and4 i_484(.A(n_3171), .B(n_3170), .C(n_3168), .D(n_2818), .Z(n_3173
		));
	notech_ao4 i_476(.A(n_58025), .B(n_42339), .C(n_58009), .D(n_42355), .Z(n_3174
		));
	notech_ao4 i_477(.A(n_58321), .B(n_42307), .C(n_58041), .D(n_42323), .Z(n_3175
		));
	notech_ao4 i_478(.A(n_58353), .B(n_42281), .C(n_58337), .D(n_42291), .Z(n_3177
		));
	notech_ao4 i_479(.A(n_58272), .B(n_42233), .C(n_58369), .D(n_42265), .Z(n_3178
		));
	notech_and4 i_485(.A(n_3178), .B(n_3177), .C(n_3175), .D(n_3174), .Z(n_3180
		));
	notech_ao4 i_597(.A(n_58305), .B(n_42262), .C(n_58289), .D(n_42278), .Z(n_3182
		));
	notech_ao4 i_598(.A(n_58249), .B(n_42246), .C(n_57961), .D(n_42413), .Z(n_3184
		));
	notech_ao4 i_599(.A(n_57993), .B(n_42381), .C(n_57977), .D(n_42397), .Z(n_3185
		));
	notech_and4 i_608(.A(n_3185), .B(n_3184), .C(n_3182), .D(n_2834), .Z(n_3187
		));
	notech_ao4 i_600(.A(n_58025), .B(n_42349), .C(n_58009), .D(n_42365), .Z(n_3188
		));
	notech_ao4 i_601(.A(n_58321), .B(n_42317), .C(n_58041), .D(n_42333), .Z(n_3189
		));
	notech_ao4 i_602(.A(n_58353), .B(n_42286), .C(n_58337), .D(n_42301), .Z(n_3191
		));
	notech_ao4 i_603(.A(n_58272), .B(n_42238), .C(n_58369), .D(n_42270), .Z(n_3192
		));
	notech_and4 i_609(.A(n_3192), .B(n_3191), .C(n_3189), .D(n_3188), .Z(n_3194
		));
	notech_ao4 i_628(.A(n_58301), .B(n_42263), .C(n_58285), .D(n_42279), .Z(n_3196
		));
	notech_ao4 i_629(.A(n_58249), .B(n_42247), .C(n_57957), .D(n_42415), .Z(n_3198
		));
	notech_ao4 i_630(.A(n_57989), .B(n_42383), .C(n_57973), .D(n_42399), .Z(n_3199
		));
	notech_and4 i_639(.A(n_3199), .B(n_3198), .C(n_3196), .D(n_2850), .Z(n_3201
		));
	notech_ao4 i_631(.A(n_58021), .B(n_42351), .C(n_58005), .D(n_42367), .Z(n_3202
		));
	notech_ao4 i_632(.A(n_58317), .B(n_42319), .C(n_58037), .D(n_42335), .Z(n_3203
		));
	notech_ao4 i_633(.A(n_58353), .B(n_42287), .C(n_58333), .D(n_42303), .Z(n_3205
		));
	notech_ao4 i_634(.A(n_58272), .B(n_42239), .C(n_58369), .D(n_42271), .Z(n_3206
		));
	notech_and4 i_640(.A(n_3206), .B(n_3205), .C(n_3203), .D(n_3202), .Z(n_3208
		));
	notech_ao4 i_845(.A(n_58301), .B(n_42270), .C(n_58285), .D(n_42286), .Z(n_3210
		));
	notech_ao4 i_846(.A(n_58249), .B(n_42254), .C(n_57957), .D(n_42429), .Z(n_3212
		));
	notech_ao4 i_847(.A(n_57989), .B(n_42397), .C(n_57973), .D(n_42413), .Z(n_3213
		));
	notech_and4 i_856(.A(n_3213), .B(n_3212), .C(n_3210), .D(n_2866), .Z(n_3215
		));
	notech_ao4 i_848(.A(n_58021), .B(n_42365), .C(n_58005), .D(n_42381), .Z(n_3216
		));
	notech_ao4 i_849(.A(n_58317), .B(n_42333), .C(n_58037), .D(n_42349), .Z(n_3217
		));
	notech_ao4 i_850(.A(n_58349), .B(n_42301), .C(n_58333), .D(n_42317), .Z(n_3219
		));
	notech_ao4 i_851(.A(n_58267), .B(n_42246), .C(n_58365), .D(n_42278), .Z(n_3220
		));
	notech_and4 i_857(.A(n_3220), .B(n_3219), .C(n_3217), .D(n_3216), .Z(n_3222
		));
	notech_ao4 i_876(.A(n_58301), .B(n_42271), .C(n_58285), .D(n_42287), .Z(n_3224
		));
	notech_ao4 i_877(.A(n_58249), .B(n_42255), .C(n_57957), .D(n_42431), .Z(n_3226
		));
	notech_ao4 i_878(.A(n_57989), .B(n_42399), .C(n_57973), .D(n_42415), .Z(n_3227
		));
	notech_and4 i_887(.A(n_3227), .B(n_3226), .C(n_3224), .D(n_2882), .Z(n_3229
		));
	notech_ao4 i_879(.A(n_58021), .B(n_42367), .C(n_58005), .D(n_42383), .Z(n_3230
		));
	notech_ao4 i_880(.A(n_58317), .B(n_42335), .C(n_58037), .D(n_42351), .Z(n_3231
		));
	notech_ao4 i_881(.A(n_58349), .B(n_42303), .C(n_58333), .D(n_42319), .Z(n_3233
		));
	notech_ao4 i_882(.A(n_58267), .B(n_42247), .C(n_58365), .D(n_42279), .Z(n_3234
		));
	notech_and4 i_888(.A(n_3234), .B(n_3233), .C(n_3231), .D(n_3230), .Z(n_3236
		));
	notech_ao4 i_1093(.A(n_58301), .B(n_42278), .C(n_58285), .D(n_42301), .Z
		(n_3238));
	notech_ao4 i_1094(.A(n_58249), .B(n_42262), .C(n_57957), .D(n_42445), .Z
		(n_3240));
	notech_ao4 i_1095(.A(n_57989), .B(n_42413), .C(n_57973), .D(n_42429), .Z
		(n_3241));
	notech_and4 i_1104(.A(n_3241), .B(n_3240), .C(n_3238), .D(n_2898), .Z(n_3243
		));
	notech_ao4 i_1096(.A(n_58021), .B(n_42381), .C(n_58005), .D(n_42397), .Z
		(n_3244));
	notech_ao4 i_1097(.A(n_58317), .B(n_42349), .C(n_58037), .D(n_42365), .Z
		(n_3245));
	notech_ao4 i_1098(.A(n_58349), .B(n_42317), .C(n_58333), .D(n_42333), .Z
		(n_3247));
	notech_ao4 i_1099(.A(n_58267), .B(n_42254), .C(n_58365), .D(n_42286), .Z
		(n_3248));
	notech_and4 i_1105(.A(n_3248), .B(n_3247), .C(n_3245), .D(n_3244), .Z(n_3250
		));
	notech_ao4 i_1124(.A(n_58301), .B(n_42279), .C(n_58285), .D(n_42303), .Z
		(n_3252));
	notech_ao4 i_1125(.A(n_58249), .B(n_42263), .C(n_57957), .D(n_42447), .Z
		(n_3254));
	notech_ao4 i_1126(.A(n_57989), .B(n_42415), .C(n_57973), .D(n_42431), .Z
		(n_3255));
	notech_and4 i_1135(.A(n_3255), .B(n_3254), .C(n_3252), .D(n_2914), .Z(n_3257
		));
	notech_ao4 i_1127(.A(n_58021), .B(n_42383), .C(n_58005), .D(n_42399), .Z
		(n_3258));
	notech_ao4 i_1128(.A(n_58317), .B(n_42351), .C(n_58037), .D(n_42367), .Z
		(n_3259));
	notech_ao4 i_1129(.A(n_58349), .B(n_42319), .C(n_58333), .D(n_42335), .Z
		(n_3261));
	notech_ao4 i_1130(.A(n_58267), .B(n_42255), .C(n_58365), .D(n_42287), .Z
		(n_3262));
	notech_and4 i_1136(.A(n_3262), .B(n_3261), .C(n_3259), .D(n_3258), .Z(n_3264
		));
	notech_ao4 i_1341(.A(n_58301), .B(n_42286), .C(n_58285), .D(n_42317), .Z
		(n_3266));
	notech_ao4 i_1342(.A(n_58253), .B(n_42270), .C(n_57957), .D(n_42461), .Z
		(n_3268));
	notech_ao4 i_1343(.A(n_57989), .B(n_42429), .C(n_57973), .D(n_42445), .Z
		(n_3269));
	notech_and4 i_1352(.A(n_3269), .B(n_3268), .C(n_3266), .D(n_2930), .Z(n_3271
		));
	notech_ao4 i_1344(.A(n_58021), .B(n_42397), .C(n_58005), .D(n_42413), .Z
		(n_3272));
	notech_ao4 i_1345(.A(n_58317), .B(n_42365), .C(n_58037), .D(n_42381), .Z
		(n_3273));
	notech_ao4 i_1346(.A(n_58349), .B(n_42333), .C(n_58333), .D(n_42349), .Z
		(n_3275));
	notech_ao4 i_1347(.A(n_58267), .B(n_42262), .C(n_58365), .D(n_42301), .Z
		(n_3276));
	notech_and4 i_1353(.A(n_3276), .B(n_3275), .C(n_3273), .D(n_3272), .Z(n_3278
		));
	notech_ao4 i_1372(.A(n_58301), .B(n_42287), .C(n_58285), .D(n_42319), .Z
		(n_3280));
	notech_ao4 i_1373(.A(n_58253), .B(n_42271), .C(n_57957), .D(n_42463), .Z
		(n_3282));
	notech_ao4 i_1374(.A(n_57989), .B(n_42431), .C(n_57973), .D(n_42447), .Z
		(n_3283));
	notech_and4 i_1383(.A(n_3283), .B(n_3282), .C(n_3280), .D(n_2948), .Z(n_3285
		));
	notech_ao4 i_1375(.A(n_58021), .B(n_42399), .C(n_58005), .D(n_42415), .Z
		(n_3286));
	notech_ao4 i_1376(.A(n_58317), .B(n_42367), .C(n_58037), .D(n_42383), .Z
		(n_3287));
	notech_ao4 i_1377(.A(n_58349), .B(n_42335), .C(n_58333), .D(n_42351), .Z
		(n_3289));
	notech_ao4 i_1378(.A(n_58267), .B(n_42263), .C(n_58365), .D(n_42303), .Z
		(n_3290));
	notech_and4 i_1384(.A(n_3290), .B(n_3289), .C(n_3287), .D(n_3286), .Z(n_3292
		));
	notech_ao4 i_1589(.A(n_58301), .B(n_42301), .C(n_58285), .D(n_42333), .Z
		(n_3294));
	notech_ao4 i_1590(.A(n_58253), .B(n_42278), .C(n_57957), .D(n_42477), .Z
		(n_3296));
	notech_ao4 i_1591(.A(n_57989), .B(n_42445), .C(n_57973), .D(n_42461), .Z
		(n_3297));
	notech_and4 i_1600(.A(n_3297), .B(n_3296), .C(n_3294), .D(n_296493405), 
		.Z(n_3299));
	notech_ao4 i_1592(.A(n_58021), .B(n_42413), .C(n_58005), .D(n_42429), .Z
		(n_3300));
	notech_ao4 i_1593(.A(n_58317), .B(n_42381), .C(n_58037), .D(n_42397), .Z
		(n_3301));
	notech_ao4 i_1594(.A(n_58349), .B(n_42349), .C(n_58333), .D(n_42365), .Z
		(n_3303));
	notech_ao4 i_1595(.A(n_58272), .B(n_42270), .C(n_58365), .D(n_42317), .Z
		(n_3304));
	notech_and4 i_1601(.A(n_3304), .B(n_3303), .C(n_3301), .D(n_3300), .Z(n_3306
		));
	notech_ao4 i_1620(.A(n_58301), .B(n_42303), .C(n_58285), .D(n_42335), .Z
		(n_3308));
	notech_ao4 i_1621(.A(n_58253), .B(n_42279), .C(n_57957), .D(n_42479), .Z
		(n_3310));
	notech_ao4 i_1622(.A(n_57989), .B(n_42447), .C(n_57973), .D(n_42463), .Z
		(n_3311));
	notech_and4 i_1631(.A(n_3311), .B(n_3310), .C(n_3308), .D(n_298096992), 
		.Z(n_3313));
	notech_ao4 i_1623(.A(n_58021), .B(n_42415), .C(n_58005), .D(n_42431), .Z
		(n_3314));
	notech_ao4 i_1624(.A(n_58317), .B(n_42383), .C(n_58037), .D(n_42399), .Z
		(n_3315));
	notech_ao4 i_1625(.A(n_58349), .B(n_42351), .C(n_58333), .D(n_42367), .Z
		(n_3317));
	notech_ao4 i_1626(.A(n_58272), .B(n_42271), .C(n_58365), .D(n_42319), .Z
		(n_3318));
	notech_and4 i_1632(.A(n_3318), .B(n_3317), .C(n_3315), .D(n_3314), .Z(n_3320
		));
	notech_ao4 i_1837(.A(n_58301), .B(n_42317), .C(n_58285), .D(n_42349), .Z
		(n_3322));
	notech_ao4 i_1838(.A(n_58249), .B(n_42286), .C(n_57957), .D(n_42493), .Z
		(n_3324));
	notech_ao4 i_1839(.A(n_57989), .B(n_42461), .C(n_57973), .D(n_42477), .Z
		(n_3325));
	notech_and4 i_1848(.A(n_3325), .B(n_3324), .C(n_3322), .D(n_2996), .Z(n_3327
		));
	notech_ao4 i_1840(.A(n_58021), .B(n_42429), .C(n_58005), .D(n_42445), .Z
		(n_3328));
	notech_ao4 i_1841(.A(n_58317), .B(n_42397), .C(n_58037), .D(n_42413), .Z
		(n_3329));
	notech_ao4 i_1842(.A(n_58349), .B(n_42365), .C(n_58333), .D(n_42381), .Z
		(n_3331));
	notech_ao4 i_1843(.A(n_58267), .B(n_42278), .C(n_58365), .D(n_42333), .Z
		(n_3332));
	notech_and4 i_1849(.A(n_3332), .B(n_3331), .C(n_3329), .D(n_3328), .Z(n_3334
		));
	notech_ao4 i_1868(.A(n_58305), .B(n_42319), .C(n_58289), .D(n_42351), .Z
		(n_3336));
	notech_ao4 i_1869(.A(n_58249), .B(n_42287), .C(n_57961), .D(n_42495), .Z
		(n_3338));
	notech_ao4 i_1870(.A(n_57993), .B(n_42463), .C(n_57977), .D(n_42479), .Z
		(n_3339));
	notech_and4 i_1879(.A(n_3339), .B(n_3338), .C(n_3336), .D(n_3012), .Z(n_3341
		));
	notech_ao4 i_1871(.A(n_58025), .B(n_42431), .C(n_58009), .D(n_42447), .Z
		(n_3342));
	notech_ao4 i_1872(.A(n_58321), .B(n_42399), .C(n_58041), .D(n_42415), .Z
		(n_3343));
	notech_ao4 i_1873(.A(n_58349), .B(n_42367), .C(n_58337), .D(n_42383), .Z
		(n_3345));
	notech_ao4 i_1874(.A(n_58267), .B(n_42279), .C(n_58365), .D(n_42335), .Z
		(n_3346));
	notech_and4 i_1880(.A(n_3346), .B(n_3345), .C(n_3343), .D(n_3342), .Z(n_3348
		));
	notech_ao4 i_2085(.A(n_58307), .B(n_42333), .C(n_58291), .D(n_42365), .Z
		(n_3350));
	notech_ao4 i_2086(.A(n_58253), .B(n_42301), .C(n_57963), .D(n_42509), .Z
		(n_3352));
	notech_ao4 i_2087(.A(n_57995), .B(n_42477), .C(n_57979), .D(n_42493), .Z
		(n_3353));
	notech_and4 i_2096(.A(n_3353), .B(n_3352), .C(n_3350), .D(n_3028), .Z(n_3355
		));
	notech_ao4 i_2088(.A(n_58027), .B(n_42445), .C(n_58011), .D(n_42461), .Z
		(n_3356));
	notech_ao4 i_2089(.A(n_58323), .B(n_42413), .C(n_58043), .D(n_42429), .Z
		(n_3357));
	notech_ao4 i_2090(.A(n_58353), .B(n_42381), .C(n_58339), .D(n_42397), .Z
		(n_3359));
	notech_ao4 i_2091(.A(n_58267), .B(n_42286), .C(n_58369), .D(n_42349), .Z
		(n_3360));
	notech_and4 i_2097(.A(n_3360), .B(n_3359), .C(n_3357), .D(n_3356), .Z(n_3362
		));
	notech_ao4 i_2116(.A(n_58307), .B(n_42335), .C(n_58291), .D(n_42367), .Z
		(n_3364));
	notech_ao4 i_2117(.A(n_58253), .B(n_42303), .C(n_57963), .D(n_42511), .Z
		(n_3366));
	notech_ao4 i_2118(.A(n_57995), .B(n_42479), .C(n_57979), .D(n_42495), .Z
		(n_3367));
	notech_and4 i_2127(.A(n_3367), .B(n_3366), .C(n_3364), .D(n_3044), .Z(n_3369
		));
	notech_ao4 i_2119(.A(n_58027), .B(n_42447), .C(n_58011), .D(n_42463), .Z
		(n_3370));
	notech_ao4 i_2120(.A(n_58323), .B(n_42415), .C(n_58043), .D(n_42431), .Z
		(n_3371));
	notech_ao4 i_2121(.A(n_58355), .B(n_42383), .C(n_58339), .D(n_42399), .Z
		(n_3373));
	notech_ao4 i_2122(.A(n_58272), .B(n_42287), .C(n_58371), .D(n_42351), .Z
		(n_3374));
	notech_and4 i_2128(.A(n_3374), .B(n_3373), .C(n_3371), .D(n_3370), .Z(n_3376
		));
	notech_ao4 i_2364(.A(n_58307), .B(n_42351), .C(n_58291), .D(n_42383), .Z
		(n_3378));
	notech_ao4 i_2365(.A(n_58256), .B(n_42319), .C(n_57963), .D(n_42527), .Z
		(n_3380));
	notech_ao4 i_2366(.A(n_57995), .B(n_42495), .C(n_57979), .D(n_42511), .Z
		(n_3381));
	notech_and4 i_2375(.A(n_3381), .B(n_3380), .C(n_3378), .D(n_3060), .Z(n_3383
		));
	notech_ao4 i_2367(.A(n_58027), .B(n_42463), .C(n_58011), .D(n_42479), .Z
		(n_3384));
	notech_ao4 i_2368(.A(n_58323), .B(n_42431), .C(n_58043), .D(n_42447), .Z
		(n_3385));
	notech_ao4 i_2369(.A(n_58355), .B(n_42399), .C(n_58339), .D(n_42415), .Z
		(n_3387));
	notech_ao4 i_2370(.A(n_58274), .B(n_42303), .C(n_58371), .D(n_42367), .Z
		(n_3388));
	notech_and4 i_2376(.A(n_3388), .B(n_3387), .C(n_3385), .D(n_3384), .Z(n_3390
		));
	notech_ao4 i_227172(.A(n_1119), .B(addrshft[1]), .C(n_112493391), .D(n_112593392
		), .Z(valid_len_197052));
	notech_ao4 i_327173(.A(n_3392), .B(addrshft[2]), .C(n_112493391), .D(n_1112
		), .Z(valid_len_297051));
	notech_ao4 i_427174(.A(n_1119), .B(addrshft[3]), .C(n_112493391), .D(n_1107
		), .Z(valid_len_397050));
	notech_ao3 i_627176(.A(n_60283), .B(addrshft[5]), .C(wptr[0]), .Z(valid_len
		[5]));
	notech_or2 i_331094(.A(wptr[0]), .B(n_42170), .Z(n_3392));
	notech_ao4 i_128277409(.A(n_58142), .B(n_42236), .C(n_58129), .D(n_42244
		), .Z(n_2537));
	notech_ao4 i_128077411(.A(n_58256), .B(n_42220), .C(n_58237), .D(n_42228
		), .Z(n_2535));
	notech_ao4 i_125777434(.A(n_1999), .B(n_42327), .C(n_1998), .D(n_42311),
		 .Z(n_2532));
	notech_ao4 i_125677435(.A(n_1996), .B(n_42295), .C(n_1995), .D(n_42359),
		 .Z(n_2531));
	notech_and3 i_125977432(.A(n_2528), .B(n_2527), .C(n_1775), .Z(n_2530)
		);
	notech_ao4 i_125377438(.A(n_1991), .B(n_42275), .C(n_1990), .D(n_42259),
		 .Z(n_2528));
	notech_ao4 i_125277439(.A(n_1988), .B(n_42251), .C(n_1987), .D(n_42267),
		 .Z(n_2527));
	notech_and4 i_126177430(.A(n_2521), .B(n_2523), .C(n_2525), .D(n_1762), 
		.Z(n_2526));
	notech_ao4 i_125877433(.A(n_1984), .B(n_42283), .C(n_1983), .D(n_42343),
		 .Z(n_2525));
	notech_ao4 i_125177440(.A(n_1979), .B(n_42235), .C(n_1978), .D(n_42243),
		 .Z(n_2523));
	notech_ao4 i_124977442(.A(n_58256), .B(n_42219), .C(n_58237), .D(n_42227
		), .Z(n_2521));
	notech_ao4 i_122677465(.A(n_1999), .B(n_42325), .C(n_1998), .D(n_42309),
		 .Z(n_2518));
	notech_ao4 i_122577466(.A(n_1996), .B(n_42293), .C(n_1995), .D(n_42357),
		 .Z(n_2517));
	notech_and3 i_122877463(.A(n_2514), .B(n_2513), .C(n_1759), .Z(n_2516)
		);
	notech_ao4 i_122277469(.A(n_1991), .B(n_42274), .C(n_1990), .D(n_42258),
		 .Z(n_2514));
	notech_ao4 i_122177470(.A(n_1988), .B(n_42250), .C(n_1987), .D(n_42266),
		 .Z(n_2513));
	notech_and4 i_123077461(.A(n_2507), .B(n_2509), .C(n_2511), .D(n_1746), 
		.Z(n_2512));
	notech_ao4 i_122777464(.A(n_1984), .B(n_42282), .C(n_1983), .D(n_42341),
		 .Z(n_2511));
	notech_ao4 i_122077471(.A(n_1979), .B(n_42234), .C(n_1978), .D(n_42242),
		 .Z(n_2509));
	notech_ao4 i_121877473(.A(n_58256), .B(n_42218), .C(n_58237), .D(n_42226
		), .Z(n_2507));
	notech_ao4 i_119577496(.A(n_1999), .B(n_42323), .C(n_1998), .D(n_42307),
		 .Z(n_2504));
	notech_ao4 i_119477497(.A(n_1996), .B(n_42291), .C(n_1995), .D(n_42355),
		 .Z(n_2503));
	notech_and3 i_119777494(.A(n_2500), .B(n_2499), .C(n_1743), .Z(n_2502)
		);
	notech_ao4 i_119177500(.A(n_1991), .B(n_42273), .C(n_1990), .D(n_42257),
		 .Z(n_2500));
	notech_ao4 i_119077501(.A(n_1988), .B(n_42249), .C(n_1987), .D(n_42265),
		 .Z(n_2499));
	notech_and4 i_119977492(.A(n_2493), .B(n_2495), .C(n_2497), .D(n_1730), 
		.Z(n_2498));
	notech_ao4 i_119677495(.A(n_1984), .B(n_42281), .C(n_1983), .D(n_42339),
		 .Z(n_2497));
	notech_ao4 i_118977502(.A(n_1979), .B(n_42233), .C(n_1978), .D(n_42241),
		 .Z(n_2495));
	notech_ao4 i_118777504(.A(n_58256), .B(n_42217), .C(n_58274), .D(n_42209
		), .Z(n_2493));
	notech_ao4 i_116477527(.A(n_1999), .B(n_42321), .C(n_1998), .D(n_42305),
		 .Z(n_2490));
	notech_ao4 i_116377528(.A(n_1996), .B(n_42288), .C(n_1995), .D(n_42353),
		 .Z(n_2489));
	notech_and3 i_116677525(.A(n_2486), .B(n_2485), .C(n_1727), .Z(n_2488)
		);
	notech_ao4 i_116077531(.A(n_1991), .B(n_42272), .C(n_1990), .D(n_42256),
		 .Z(n_2486));
	notech_ao4 i_115977532(.A(n_1988), .B(n_42248), .C(n_1987), .D(n_42264),
		 .Z(n_2485));
	notech_and4 i_116877523(.A(n_2479), .B(n_2481), .C(n_2483), .D(n_1714), 
		.Z(n_2484));
	notech_ao4 i_116577526(.A(n_1984), .B(n_42280), .C(n_1983), .D(n_42337),
		 .Z(n_2483));
	notech_ao4 i_115877533(.A(n_1979), .B(n_42232), .C(n_1978), .D(n_42240),
		 .Z(n_2481));
	notech_ao4 i_115677535(.A(n_58256), .B(n_42216), .C(n_58237), .D(n_42224
		), .Z(n_2479));
	notech_ao4 i_113377558(.A(n_1999), .B(n_42319), .C(n_1998), .D(n_42303),
		 .Z(n_2476));
	notech_ao4 i_113277559(.A(n_1996), .B(n_42287), .C(n_1995), .D(n_42351),
		 .Z(n_2475));
	notech_and3 i_113577556(.A(n_2472), .B(n_2471), .C(n_1711), .Z(n_2474)
		);
	notech_ao4 i_112977562(.A(n_1991), .B(n_42271), .C(n_1990), .D(n_42255),
		 .Z(n_2472));
	notech_ao4 i_112877563(.A(n_1988), .B(n_42247), .C(n_1987), .D(n_42263),
		 .Z(n_2471));
	notech_and4 i_113777554(.A(n_2465), .B(n_2467), .C(n_2469), .D(n_1698), 
		.Z(n_2470));
	notech_ao4 i_113477557(.A(n_1984), .B(n_42279), .C(n_1983), .D(n_42335),
		 .Z(n_2469));
	notech_ao4 i_112777564(.A(n_1979), .B(n_42231), .C(n_1978), .D(n_42239),
		 .Z(n_2467));
	notech_ao4 i_112577566(.A(n_58256), .B(n_42215), .C(n_58237), .D(n_42223
		), .Z(n_2465));
	notech_ao4 i_110277589(.A(n_1999), .B(n_42315), .C(n_1998), .D(n_42299),
		 .Z(n_2462));
	notech_ao4 i_110177590(.A(n_1996), .B(n_42285), .C(n_1995), .D(n_42347),
		 .Z(n_2461));
	notech_and3 i_110477587(.A(n_2458), .B(n_2457), .C(n_1695), .Z(n_2460)
		);
	notech_ao4 i_109877593(.A(n_1991), .B(n_42269), .C(n_1990), .D(n_42253),
		 .Z(n_2458));
	notech_ao4 i_109777594(.A(n_1988), .B(n_42245), .C(n_1987), .D(n_42261),
		 .Z(n_2457));
	notech_and4 i_110677585(.A(n_2451), .B(n_2453), .C(n_2455), .D(n_1682), 
		.Z(n_2456));
	notech_ao4 i_110377588(.A(n_1984), .B(n_42277), .C(n_1983), .D(n_42331),
		 .Z(n_2455));
	notech_ao4 i_109677595(.A(n_1979), .B(n_42229), .C(n_1978), .D(n_42237),
		 .Z(n_2453));
	notech_ao4 i_109477597(.A(n_58256), .B(n_42213), .C(n_58237), .D(n_42221
		), .Z(n_2451));
	notech_ao4 i_107177620(.A(n_1999), .B(n_42313), .C(n_1998), .D(n_42297),
		 .Z(n_2448));
	notech_ao4 i_107077621(.A(n_1996), .B(n_42284), .C(n_1995), .D(n_42345),
		 .Z(n_2447));
	notech_and3 i_107377618(.A(n_2444), .B(n_2443), .C(n_1679), .Z(n_2446)
		);
	notech_ao4 i_106777624(.A(n_1991), .B(n_42268), .C(n_1990), .D(n_42252),
		 .Z(n_2444));
	notech_ao4 i_106677625(.A(n_1988), .B(n_42244), .C(n_1987), .D(n_42260),
		 .Z(n_2443));
	notech_and4 i_107577616(.A(n_2437), .B(n_2439), .C(n_2441), .D(n_1666), 
		.Z(n_2442));
	notech_ao4 i_107277619(.A(n_1984), .B(n_42276), .C(n_1983), .D(n_42329),
		 .Z(n_2441));
	notech_ao4 i_106577626(.A(n_1979), .B(n_42228), .C(n_1978), .D(n_42236),
		 .Z(n_2439));
	notech_ao4 i_106377628(.A(n_58256), .B(n_42212), .C(n_58237), .D(n_42220
		), .Z(n_2437));
	notech_ao4 i_104077651(.A(n_1999), .B(n_42311), .C(n_1998), .D(n_42295),
		 .Z(n_2434));
	notech_ao4 i_103977652(.A(n_1996), .B(n_42283), .C(n_1995), .D(n_42343),
		 .Z(n_2433));
	notech_and3 i_104277649(.A(n_2430), .B(n_2429), .C(n_1663), .Z(n_2432)
		);
	notech_ao4 i_103677655(.A(n_1991), .B(n_42267), .C(n_1990), .D(n_42251),
		 .Z(n_2430));
	notech_ao4 i_103577656(.A(n_1988), .B(n_42243), .C(n_1987), .D(n_42259),
		 .Z(n_2429));
	notech_and4 i_104477647(.A(n_2423), .B(n_2425), .C(n_2427), .D(n_1650), 
		.Z(n_2428));
	notech_ao4 i_104177650(.A(n_1984), .B(n_42275), .C(n_1983), .D(n_42327),
		 .Z(n_2427));
	notech_ao4 i_103477657(.A(n_1979), .B(n_42227), .C(n_1978), .D(n_42235),
		 .Z(n_2425));
	notech_ao4 i_103277659(.A(n_58256), .B(n_42211), .C(n_58237), .D(n_42219
		), .Z(n_2423));
	notech_ao4 i_100977682(.A(n_1999), .B(n_42309), .C(n_1998), .D(n_42293),
		 .Z(n_2420));
	notech_ao4 i_100877683(.A(n_1996), .B(n_42282), .C(n_1995), .D(n_42341),
		 .Z(n_2419));
	notech_and3 i_101177680(.A(n_2416), .B(n_2415), .C(n_1647), .Z(n_2418)
		);
	notech_ao4 i_100577686(.A(n_1991), .B(n_42266), .C(n_1990), .D(n_42250),
		 .Z(n_2416));
	notech_ao4 i_100477687(.A(n_1988), .B(n_42242), .C(n_1987), .D(n_42258),
		 .Z(n_2415));
	notech_and4 i_101377678(.A(n_2409), .B(n_2411), .C(n_2413), .D(n_1634), 
		.Z(n_2414));
	notech_ao4 i_101077681(.A(n_1984), .B(n_42274), .C(n_1983), .D(n_42325),
		 .Z(n_2413));
	notech_ao4 i_100377688(.A(n_1979), .B(n_42226), .C(n_1978), .D(n_42234),
		 .Z(n_2411));
	notech_ao4 i_100177690(.A(n_58256), .B(n_42210), .C(n_58237), .D(n_42218
		), .Z(n_2409));
	notech_ao4 i_97877713(.A(n_1999), .B(n_42307), .C(n_1998), .D(n_42291), 
		.Z(n_2406));
	notech_ao4 i_97777714(.A(n_1996), .B(n_42281), .C(n_1995), .D(n_42339), 
		.Z(n_2405));
	notech_and3 i_98077711(.A(n_2402), .B(n_2401), .C(n_1631), .Z(n_2404));
	notech_ao4 i_97477717(.A(n_1991), .B(n_42265), .C(n_1990), .D(n_42249), 
		.Z(n_2402));
	notech_ao4 i_97377718(.A(n_1988), .B(n_42241), .C(n_1987), .D(n_42257), 
		.Z(n_2401));
	notech_and4 i_98277709(.A(n_2395), .B(n_2397), .C(n_2399), .D(n_1618), .Z
		(n_2400));
	notech_ao4 i_97977712(.A(n_1984), .B(n_42273), .C(n_1983), .D(n_42323), 
		.Z(n_2399));
	notech_ao4 i_97277719(.A(n_1979), .B(n_42225), .C(n_1978), .D(n_42233), 
		.Z(n_2397));
	notech_ao4 i_97077721(.A(n_58237), .B(n_42217), .C(n_58256), .D(n_42209)
		, .Z(n_2395));
	notech_ao4 i_94777744(.A(n_1999), .B(n_42305), .C(n_1998), .D(n_42288), 
		.Z(n_2392));
	notech_ao4 i_94677745(.A(n_1996), .B(n_42280), .C(n_1995), .D(n_42337), 
		.Z(n_2391));
	notech_and3 i_94977742(.A(n_2388), .B(n_2387), .C(n_1615), .Z(n_2390));
	notech_ao4 i_94377748(.A(n_1991), .B(n_42264), .C(n_1990), .D(n_42248), 
		.Z(n_2388));
	notech_ao4 i_94277749(.A(n_1988), .B(n_42240), .C(n_1987), .D(n_42256), 
		.Z(n_2387));
	notech_and4 i_95177740(.A(n_2381), .B(n_2383), .C(n_2385), .D(n_1602), .Z
		(n_2386));
	notech_ao4 i_94877743(.A(n_1984), .B(n_42272), .C(n_1983), .D(n_42321), 
		.Z(n_2385));
	notech_ao4 i_94177750(.A(n_1979), .B(n_42224), .C(n_1978), .D(n_42232), 
		.Z(n_2383));
	notech_ao4 i_93977752(.A(n_58256), .B(n_42208), .C(n_58237), .D(n_42216)
		, .Z(n_2381));
	notech_ao4 i_91677775(.A(n_1999), .B(n_42303), .C(n_1998), .D(n_42287), 
		.Z(n_2378));
	notech_ao4 i_91577776(.A(n_1996), .B(n_42279), .C(n_1995), .D(n_42335), 
		.Z(n_2377));
	notech_and3 i_91877773(.A(n_2374), .B(n_2373), .C(n_1599), .Z(n_2376));
	notech_ao4 i_91277779(.A(n_1991), .B(n_42263), .C(n_1990), .D(n_42247), 
		.Z(n_2374));
	notech_ao4 i_91177780(.A(n_1988), .B(n_42239), .C(n_1987), .D(n_42255), 
		.Z(n_2373));
	notech_and4 i_92077771(.A(n_2367), .B(n_2369), .C(n_2371), .D(n_1586), .Z
		(n_2372));
	notech_ao4 i_91777774(.A(n_1984), .B(n_42271), .C(n_1983), .D(n_42319), 
		.Z(n_2371));
	notech_ao4 i_91077781(.A(n_1979), .B(n_42223), .C(n_1978), .D(n_42231), 
		.Z(n_2369));
	notech_ao4 i_90877783(.A(n_58256), .B(n_42207), .C(n_58237), .D(n_42215)
		, .Z(n_2367));
	notech_ao4 i_88577806(.A(n_1999), .B(n_42299), .C(n_1998), .D(n_42285), 
		.Z(n_2364));
	notech_ao4 i_88477807(.A(n_1996), .B(n_42277), .C(n_1995), .D(n_42331), 
		.Z(n_2363));
	notech_and3 i_88777804(.A(n_2360), .B(n_2359), .C(n_1583), .Z(n_2362));
	notech_ao4 i_88177810(.A(n_1991), .B(n_42261), .C(n_1990), .D(n_42245), 
		.Z(n_2360));
	notech_ao4 i_88077811(.A(n_1988), .B(n_42237), .C(n_1987), .D(n_42253), 
		.Z(n_2359));
	notech_and4 i_88977802(.A(n_2353), .B(n_2355), .C(n_2357), .D(n_1570), .Z
		(n_2358));
	notech_ao4 i_88677805(.A(n_1984), .B(n_42269), .C(n_1983), .D(n_42315), 
		.Z(n_2357));
	notech_ao4 i_87977812(.A(n_1979), .B(n_42221), .C(n_1978), .D(n_42229), 
		.Z(n_2355));
	notech_ao4 i_87777814(.A(n_58256), .B(n_42205), .C(n_58237), .D(n_42213)
		, .Z(n_2353));
	notech_ao4 i_85477837(.A(n_58194), .B(n_42297), .C(n_58181), .D(n_42284)
		, .Z(n_2350));
	notech_ao4 i_85377838(.A(n_58168), .B(n_42276), .C(n_58155), .D(n_42329)
		, .Z(n_2349));
	notech_and3 i_85677835(.A(n_2346), .B(n_2345), .C(n_1567), .Z(n_2348));
	notech_ao4 i_85077841(.A(n_58090), .B(n_42260), .C(n_58077), .D(n_42244)
		, .Z(n_2346));
	notech_ao4 i_84977842(.A(n_58064), .B(n_42236), .C(n_58051), .D(n_42252)
		, .Z(n_2345));
	notech_and4 i_85877833(.A(n_2339), .B(n_2341), .C(n_2343), .D(n_1554), .Z
		(n_2344));
	notech_ao4 i_85577836(.A(n_58116), .B(n_42268), .C(n_58103), .D(n_42313)
		, .Z(n_2343));
	notech_ao4 i_84877843(.A(n_58142), .B(n_42220), .C(n_58129), .D(n_42228)
		, .Z(n_2341));
	notech_ao4 i_84677845(.A(n_58256), .B(n_42204), .C(n_58237), .D(n_42212)
		, .Z(n_2339));
	notech_ao4 i_82377868(.A(n_58190), .B(n_42295), .C(n_58177), .D(n_42283)
		, .Z(n_2336));
	notech_ao4 i_82277869(.A(n_58164), .B(n_42275), .C(n_58151), .D(n_42327)
		, .Z(n_2335));
	notech_and3 i_82577866(.A(n_2332), .B(n_2331), .C(n_1551), .Z(n_2334));
	notech_ao4 i_81977872(.A(n_58086), .B(n_42259), .C(n_58073), .D(n_42243)
		, .Z(n_2332));
	notech_ao4 i_81877873(.A(n_58060), .B(n_42235), .C(n_58047), .D(n_42251)
		, .Z(n_2331));
	notech_and4 i_82777864(.A(n_2325), .B(n_2327), .C(n_2329), .D(n_1538), .Z
		(n_2330));
	notech_ao4 i_82477867(.A(n_58112), .B(n_42267), .C(n_58099), .D(n_42311)
		, .Z(n_2329));
	notech_ao4 i_81777874(.A(n_58138), .B(n_42219), .C(n_58125), .D(n_42227)
		, .Z(n_2327));
	notech_ao4 i_81577876(.A(n_58254), .B(n_42203), .C(n_58235), .D(n_42211)
		, .Z(n_2325));
	notech_ao4 i_79277899(.A(n_58190), .B(n_42293), .C(n_58177), .D(n_42282)
		, .Z(n_2322));
	notech_ao4 i_79177900(.A(n_58164), .B(n_42274), .C(n_58151), .D(n_42325)
		, .Z(n_2321));
	notech_and3 i_79477897(.A(n_2318), .B(n_2317), .C(n_1535), .Z(n_2320));
	notech_ao4 i_78877903(.A(n_58086), .B(n_42258), .C(n_58073), .D(n_42242)
		, .Z(n_2318));
	notech_ao4 i_78777904(.A(n_58060), .B(n_42234), .C(n_58047), .D(n_42250)
		, .Z(n_2317));
	notech_and4 i_79677895(.A(n_2311), .B(n_2313), .C(n_2315), .D(n_1522), .Z
		(n_2316));
	notech_ao4 i_79377898(.A(n_58112), .B(n_42266), .C(n_58099), .D(n_42309)
		, .Z(n_2315));
	notech_ao4 i_78677905(.A(n_58138), .B(n_42218), .C(n_58125), .D(n_42226)
		, .Z(n_2313));
	notech_ao4 i_78477907(.A(n_58254), .B(n_42202), .C(n_58235), .D(n_42210)
		, .Z(n_2311));
	notech_ao4 i_76177930(.A(n_58190), .B(n_42291), .C(n_58177), .D(n_42281)
		, .Z(n_2308));
	notech_ao4 i_76077931(.A(n_58164), .B(n_42273), .C(n_58151), .D(n_42323)
		, .Z(n_2307));
	notech_and3 i_76377928(.A(n_2304), .B(n_2303), .C(n_1519), .Z(n_2306));
	notech_ao4 i_75777934(.A(n_58086), .B(n_42257), .C(n_58073), .D(n_42241)
		, .Z(n_2304));
	notech_ao4 i_75677935(.A(n_58060), .B(n_42233), .C(n_58047), .D(n_42249)
		, .Z(n_2303));
	notech_and4 i_76577926(.A(n_2297), .B(n_2299), .C(n_2301), .D(n_1506), .Z
		(n_2302));
	notech_ao4 i_76277929(.A(n_58112), .B(n_42265), .C(n_58099), .D(n_42307)
		, .Z(n_2301));
	notech_ao4 i_75577936(.A(n_58138), .B(n_42217), .C(n_58125), .D(n_42225)
		, .Z(n_2299));
	notech_ao4 i_75377938(.A(n_58254), .B(n_42201), .C(n_58235), .D(n_42209)
		, .Z(n_2297));
	notech_ao4 i_73077961(.A(n_58190), .B(n_42288), .C(n_58177), .D(n_42280)
		, .Z(n_2294));
	notech_ao4 i_72977962(.A(n_58164), .B(n_42272), .C(n_58151), .D(n_42321)
		, .Z(n_2293));
	notech_and3 i_73277959(.A(n_2290), .B(n_2289), .C(n_1503), .Z(n_2292));
	notech_ao4 i_72677965(.A(n_58086), .B(n_42256), .C(n_58073), .D(n_42240)
		, .Z(n_2290));
	notech_ao4 i_72577966(.A(n_58060), .B(n_42232), .C(n_58047), .D(n_42248)
		, .Z(n_2289));
	notech_and4 i_73477957(.A(n_2283), .B(n_2285), .C(n_2287), .D(n_1490), .Z
		(n_2288));
	notech_ao4 i_73177960(.A(n_58112), .B(n_42264), .C(n_58099), .D(n_42305)
		, .Z(n_2287));
	notech_ao4 i_72477967(.A(n_58138), .B(n_42216), .C(n_58125), .D(n_42224)
		, .Z(n_2285));
	notech_ao4 i_72277969(.A(n_58254), .B(n_42200), .C(n_58235), .D(n_42208)
		, .Z(n_2283));
	notech_ao4 i_69977992(.A(n_58190), .B(n_42287), .C(n_58177), .D(n_42279)
		, .Z(n_2280));
	notech_ao4 i_69877993(.A(n_58164), .B(n_42271), .C(n_58151), .D(n_42319)
		, .Z(n_2279));
	notech_and3 i_70177990(.A(n_2276), .B(n_2275), .C(n_1487), .Z(n_2278));
	notech_ao4 i_69577996(.A(n_58086), .B(n_42255), .C(n_58073), .D(n_42239)
		, .Z(n_2276));
	notech_ao4 i_69477997(.A(n_58060), .B(n_42231), .C(n_58047), .D(n_42247)
		, .Z(n_2275));
	notech_and4 i_70377988(.A(n_2269), .B(n_2271), .C(n_2273), .D(n_1474), .Z
		(n_2274));
	notech_ao4 i_70077991(.A(n_58112), .B(n_42263), .C(n_58099), .D(n_42303)
		, .Z(n_2273));
	notech_ao4 i_69377998(.A(n_58138), .B(n_42215), .C(n_58125), .D(n_42223)
		, .Z(n_2271));
	notech_ao4 i_69178000(.A(n_58254), .B(n_42199), .C(n_58235), .D(n_42207)
		, .Z(n_2269));
	notech_ao4 i_66878023(.A(n_58190), .B(n_42286), .C(n_58177), .D(n_42278)
		, .Z(n_2266));
	notech_ao4 i_66778024(.A(n_58164), .B(n_42270), .C(n_58151), .D(n_42317)
		, .Z(n_2265));
	notech_and3 i_67078021(.A(n_2262), .B(n_2261), .C(n_1471), .Z(n_2264));
	notech_ao4 i_66478027(.A(n_58086), .B(n_42254), .C(n_58073), .D(n_42238)
		, .Z(n_2262));
	notech_ao4 i_66378028(.A(n_58060), .B(n_42230), .C(n_58047), .D(n_42246)
		, .Z(n_2261));
	notech_and4 i_67278019(.A(n_2255), .B(n_2257), .C(n_2259), .D(n_1458), .Z
		(n_2260));
	notech_ao4 i_66978022(.A(n_58112), .B(n_42262), .C(n_58099), .D(n_42301)
		, .Z(n_2259));
	notech_ao4 i_66278029(.A(n_58138), .B(n_42214), .C(n_58125), .D(n_42222)
		, .Z(n_2257));
	notech_ao4 i_66078031(.A(n_58254), .B(n_42198), .C(n_58235), .D(n_42206)
		, .Z(n_2255));
	notech_ao4 i_63778054(.A(n_58190), .B(n_42285), .C(n_58177), .D(n_42277)
		, .Z(n_2252));
	notech_ao4 i_63678055(.A(n_58164), .B(n_42269), .C(n_58151), .D(n_42315)
		, .Z(n_2251));
	notech_and3 i_63978052(.A(n_2248), .B(n_2247), .C(n_1455), .Z(n_2250));
	notech_ao4 i_63378058(.A(n_58086), .B(n_42253), .C(n_58073), .D(n_42237)
		, .Z(n_2248));
	notech_ao4 i_63278059(.A(n_58060), .B(n_42229), .C(n_58047), .D(n_42245)
		, .Z(n_2247));
	notech_and4 i_64178050(.A(n_2241), .B(n_2243), .C(n_2245), .D(n_1442), .Z
		(n_2246));
	notech_ao4 i_63878053(.A(n_58112), .B(n_42261), .C(n_58099), .D(n_42299)
		, .Z(n_2245));
	notech_ao4 i_63178060(.A(n_58138), .B(n_42213), .C(n_58125), .D(n_42221)
		, .Z(n_2243));
	notech_ao4 i_62978062(.A(n_58254), .B(n_42197), .C(n_58235), .D(n_42205)
		, .Z(n_2241));
	notech_ao4 i_60678085(.A(n_58190), .B(n_42284), .C(n_58177), .D(n_42276)
		, .Z(n_2238));
	notech_ao4 i_60578086(.A(n_58164), .B(n_42268), .C(n_58151), .D(n_42313)
		, .Z(n_2237));
	notech_and3 i_60878083(.A(n_2234), .B(n_2233), .C(n_1439), .Z(n_2236));
	notech_ao4 i_60278089(.A(n_58086), .B(n_42252), .C(n_58073), .D(n_42236)
		, .Z(n_2234));
	notech_ao4 i_60178090(.A(n_58060), .B(n_42228), .C(n_58047), .D(n_42244)
		, .Z(n_2233));
	notech_and4 i_61078081(.A(n_2227), .B(n_2229), .C(n_2231), .D(n_1426), .Z
		(n_2232));
	notech_ao4 i_60778084(.A(n_58112), .B(n_42260), .C(n_58099), .D(n_42297)
		, .Z(n_2231));
	notech_ao4 i_60078091(.A(n_58138), .B(n_42212), .C(n_58125), .D(n_42220)
		, .Z(n_2229));
	notech_ao4 i_59878093(.A(n_58254), .B(n_42196), .C(n_58235), .D(n_42204)
		, .Z(n_2227));
	notech_ao4 i_57578116(.A(n_58190), .B(n_42283), .C(n_58177), .D(n_42275)
		, .Z(n_2224));
	notech_ao4 i_57478117(.A(n_58164), .B(n_42267), .C(n_58151), .D(n_42311)
		, .Z(n_2223));
	notech_and3 i_57778114(.A(n_2220), .B(n_2219), .C(n_1423), .Z(n_2222));
	notech_ao4 i_57178120(.A(n_58086), .B(n_42251), .C(n_58073), .D(n_42235)
		, .Z(n_2220));
	notech_ao4 i_57078121(.A(n_58060), .B(n_42227), .C(n_58047), .D(n_42243)
		, .Z(n_2219));
	notech_and4 i_57978112(.A(n_2213), .B(n_2215), .C(n_2217), .D(n_1410), .Z
		(n_2218));
	notech_ao4 i_57678115(.A(n_58112), .B(n_42259), .C(n_58099), .D(n_42295)
		, .Z(n_2217));
	notech_ao4 i_56978122(.A(n_58138), .B(n_42211), .C(n_58125), .D(n_42219)
		, .Z(n_2215));
	notech_ao4 i_56778124(.A(n_58254), .B(n_42195), .C(n_58235), .D(n_42203)
		, .Z(n_2213));
	notech_ao4 i_54478147(.A(n_58190), .B(n_42282), .C(n_58177), .D(n_42274)
		, .Z(n_2210));
	notech_ao4 i_54378148(.A(n_58164), .B(n_42266), .C(n_58151), .D(n_42309)
		, .Z(n_2209));
	notech_and3 i_54678145(.A(n_2206), .B(n_2205), .C(n_1407), .Z(n_2208));
	notech_ao4 i_54078151(.A(n_58086), .B(n_42250), .C(n_58073), .D(n_42234)
		, .Z(n_2206));
	notech_ao4 i_53978152(.A(n_58060), .B(n_42226), .C(n_58047), .D(n_42242)
		, .Z(n_2205));
	notech_and4 i_54878143(.A(n_2199), .B(n_2201), .C(n_2203), .D(n_1394), .Z
		(n_2204));
	notech_ao4 i_54578146(.A(n_58112), .B(n_42258), .C(n_58099), .D(n_42293)
		, .Z(n_2203));
	notech_ao4 i_53878153(.A(n_58138), .B(n_42210), .C(n_58125), .D(n_42218)
		, .Z(n_2201));
	notech_ao4 i_53678155(.A(n_58254), .B(n_42194), .C(n_58235), .D(n_42202)
		, .Z(n_2199));
	notech_ao4 i_51378178(.A(n_58190), .B(n_42281), .C(n_58177), .D(n_42273)
		, .Z(n_2196));
	notech_ao4 i_51278179(.A(n_58164), .B(n_42265), .C(n_58151), .D(n_42307)
		, .Z(n_2195));
	notech_and3 i_51578176(.A(n_2192), .B(n_2191), .C(n_1391), .Z(n_2194));
	notech_ao4 i_50978182(.A(n_58086), .B(n_42249), .C(n_58073), .D(n_42233)
		, .Z(n_2192));
	notech_ao4 i_50878183(.A(n_58060), .B(n_42225), .C(n_58047), .D(n_42241)
		, .Z(n_2191));
	notech_and4 i_51778174(.A(n_2185), .B(n_2187), .C(n_2189), .D(n_1378), .Z
		(n_2190));
	notech_ao4 i_51478177(.A(n_58112), .B(n_42257), .C(n_58099), .D(n_42291)
		, .Z(n_2189));
	notech_ao4 i_50778184(.A(n_58138), .B(n_42209), .C(n_58125), .D(n_42217)
		, .Z(n_2187));
	notech_ao4 i_50578186(.A(n_58237), .B(n_42201), .C(n_58274), .D(n_42185)
		, .Z(n_2185));
	notech_ao4 i_48278209(.A(n_42280), .B(n_58190), .C(n_42272), .D(n_58177)
		, .Z(n_2182));
	notech_ao4 i_48178210(.A(n_42264), .B(n_58164), .C(n_42305), .D(n_58151)
		, .Z(n_2181));
	notech_and3 i_48478207(.A(n_2178), .B(n_2177), .C(n_1375), .Z(n_2180));
	notech_ao4 i_47878213(.A(n_42248), .B(n_58086), .C(n_42232), .D(n_58073)
		, .Z(n_2178));
	notech_ao4 i_47778214(.A(n_42224), .B(n_58060), .C(n_42240), .D(n_58047)
		, .Z(n_2177));
	notech_and4 i_48678205(.A(n_2171), .B(n_2173), .C(n_2175), .D(n_1362), .Z
		(n_2176));
	notech_ao4 i_48378208(.A(n_42256), .B(n_58112), .C(n_42288), .D(n_58099)
		, .Z(n_2175));
	notech_ao4 i_47678215(.A(n_42208), .B(n_58138), .C(n_42216), .D(n_58125)
		, .Z(n_2173));
	notech_ao4 i_47478217(.A(n_58256), .B(n_42192), .C(n_58237), .D(n_42200)
		, .Z(n_2171));
	notech_ao4 i_45178240(.A(n_58190), .B(n_42278), .C(n_58177), .D(n_42270)
		, .Z(n_2168));
	notech_ao4 i_45078241(.A(n_58164), .B(n_42262), .C(n_58151), .D(n_42301)
		, .Z(n_2167));
	notech_and3 i_45378238(.A(n_2164), .B(n_2163), .C(n_1359), .Z(n_2166));
	notech_ao4 i_44778244(.A(n_58086), .B(n_42246), .C(n_58073), .D(n_42230)
		, .Z(n_2164));
	notech_ao4 i_44678245(.A(n_58060), .B(n_42222), .C(n_58047), .D(n_42238)
		, .Z(n_2163));
	notech_and4 i_45578236(.A(n_2157), .B(n_2159), .C(n_2161), .D(n_1346), .Z
		(n_2162));
	notech_ao4 i_45278239(.A(n_58112), .B(n_42254), .C(n_58099), .D(n_42286)
		, .Z(n_2161));
	notech_ao4 i_44578246(.A(n_58138), .B(n_42206), .C(n_58125), .D(n_42214)
		, .Z(n_2159));
	notech_ao4 i_44378248(.A(n_58256), .B(n_42190), .C(n_58235), .D(n_42198)
		, .Z(n_2157));
	notech_ao4 i_42078271(.A(n_58194), .B(n_42277), .C(n_58181), .D(n_42269)
		, .Z(n_2154));
	notech_ao4 i_41978272(.A(n_58168), .B(n_42261), .C(n_58155), .D(n_42299)
		, .Z(n_2153));
	notech_and3 i_42278269(.A(n_2150), .B(n_2149), .C(n_1343), .Z(n_2152));
	notech_ao4 i_41678275(.A(n_58090), .B(n_42245), .C(n_58077), .D(n_42229)
		, .Z(n_2150));
	notech_ao4 i_41578276(.A(n_58064), .B(n_42221), .C(n_58051), .D(n_42237)
		, .Z(n_2149));
	notech_and4 i_42478267(.A(n_2143), .B(n_2145), .C(n_2147), .D(n_1330), .Z
		(n_2148));
	notech_ao4 i_42178270(.A(n_58116), .B(n_42253), .C(n_58103), .D(n_42285)
		, .Z(n_2147));
	notech_ao4 i_41478277(.A(n_58142), .B(n_42205), .C(n_58129), .D(n_42213)
		, .Z(n_2145));
	notech_ao4 i_41278279(.A(n_58254), .B(n_42189), .C(n_58235), .D(n_42197)
		, .Z(n_2143));
	notech_ao4 i_38978302(.A(n_58194), .B(n_42276), .C(n_58181), .D(n_42268)
		, .Z(n_2140));
	notech_ao4 i_38878303(.A(n_58168), .B(n_42260), .C(n_58155), .D(n_42297)
		, .Z(n_2139));
	notech_and3 i_39178300(.A(n_2136), .B(n_2135), .C(n_1327), .Z(n_2138));
	notech_ao4 i_38578306(.A(n_58090), .B(n_42244), .C(n_58077), .D(n_42228)
		, .Z(n_2136));
	notech_ao4 i_38478307(.A(n_58064), .B(n_42220), .C(n_58051), .D(n_42236)
		, .Z(n_2135));
	notech_and4 i_39378298(.A(n_2129), .B(n_2131), .C(n_2133), .D(n_1308), .Z
		(n_2134));
	notech_ao4 i_39078301(.A(n_58116), .B(n_42252), .C(n_58103), .D(n_42284)
		, .Z(n_2133));
	notech_ao4 i_38378308(.A(n_58142), .B(n_42204), .C(n_58129), .D(n_42212)
		, .Z(n_2131));
	notech_ao4 i_38178310(.A(n_58254), .B(n_42188), .C(n_58235), .D(n_42196)
		, .Z(n_2129));
	notech_ao4 i_35878333(.A(n_58194), .B(n_42275), .C(n_58181), .D(n_42267)
		, .Z(n_2126));
	notech_ao4 i_35778334(.A(n_58168), .B(n_42259), .C(n_58155), .D(n_42295)
		, .Z(n_2125));
	notech_and3 i_36078331(.A(n_2122), .B(n_2121), .C(n_1303), .Z(n_2124));
	notech_ao4 i_35478337(.A(n_58090), .B(n_42243), .C(n_58077), .D(n_42227)
		, .Z(n_2122));
	notech_ao4 i_35378338(.A(n_58064), .B(n_42219), .C(n_58051), .D(n_42235)
		, .Z(n_2121));
	notech_and4 i_36278329(.A(n_2115), .B(n_2117), .C(n_2119), .D(n_1282), .Z
		(n_2120));
	notech_ao4 i_35978332(.A(n_58116), .B(n_42251), .C(n_58103), .D(n_42283)
		, .Z(n_2119));
	notech_ao4 i_35278339(.A(n_58142), .B(n_42203), .C(n_58129), .D(n_42211)
		, .Z(n_2117));
	notech_ao4 i_35078341(.A(n_58254), .B(n_42187), .C(n_58235), .D(n_42195)
		, .Z(n_2115));
	notech_ao4 i_32778364(.A(n_58194), .B(n_42274), .C(n_58181), .D(n_42266)
		, .Z(n_2112));
	notech_ao4 i_32678365(.A(n_58168), .B(n_42258), .C(n_58155), .D(n_42293)
		, .Z(n_2111));
	notech_and3 i_32978362(.A(n_2108), .B(n_2107), .C(n_1279), .Z(n_2110));
	notech_ao4 i_32378368(.A(n_58090), .B(n_42242), .C(n_58077), .D(n_42226)
		, .Z(n_2108));
	notech_ao4 i_32278369(.A(n_58064), .B(n_42218), .C(n_58051), .D(n_42234)
		, .Z(n_2107));
	notech_and4 i_33178360(.A(n_2101), .B(n_2103), .C(n_2105), .D(n_1266), .Z
		(n_2106));
	notech_ao4 i_32878363(.A(n_58116), .B(n_42250), .C(n_58103), .D(n_42282)
		, .Z(n_2105));
	notech_ao4 i_32178370(.A(n_58142), .B(n_42202), .C(n_58129), .D(n_42210)
		, .Z(n_2103));
	notech_ao4 i_31978372(.A(n_58254), .B(n_42186), .C(n_58230), .D(n_42194)
		, .Z(n_2101));
	notech_ao4 i_29678395(.A(n_58194), .B(n_42273), .C(n_58181), .D(n_42265)
		, .Z(n_2098));
	notech_ao4 i_29578396(.A(n_58168), .B(n_42257), .C(n_58155), .D(n_42291)
		, .Z(n_2097));
	notech_and3 i_29878393(.A(n_2094), .B(n_2093), .C(n_1263), .Z(n_2096));
	notech_ao4 i_29278399(.A(n_58090), .B(n_42241), .C(n_58077), .D(n_42225)
		, .Z(n_2094));
	notech_ao4 i_29178400(.A(n_58064), .B(n_42217), .C(n_58051), .D(n_42233)
		, .Z(n_2093));
	notech_and4 i_30078391(.A(n_2087), .B(n_2089), .C(n_2091), .D(n_1250), .Z
		(n_2092));
	notech_ao4 i_29778394(.A(n_58116), .B(n_42249), .C(n_58103), .D(n_42281)
		, .Z(n_2091));
	notech_ao4 i_29078401(.A(n_58142), .B(n_42201), .C(n_58129), .D(n_42209)
		, .Z(n_2089));
	notech_ao4 i_28878403(.A(n_58274), .B(n_42177), .C(n_58249), .D(n_42185)
		, .Z(n_2087));
	notech_ao4 i_26578426(.A(n_58194), .B(n_42271), .C(n_58181), .D(n_42263)
		, .Z(n_2084));
	notech_ao4 i_26478427(.A(n_58168), .B(n_42255), .C(n_58155), .D(n_42287)
		, .Z(n_2083));
	notech_and3 i_26778424(.A(n_2080), .B(n_2079), .C(n_1247), .Z(n_2082));
	notech_ao4 i_26178430(.A(n_58090), .B(n_42239), .C(n_58077), .D(n_42223)
		, .Z(n_2080));
	notech_ao4 i_26078431(.A(n_58064), .B(n_42215), .C(n_58051), .D(n_42231)
		, .Z(n_2079));
	notech_and4 i_26978422(.A(n_2073), .B(n_2075), .C(n_2077), .D(n_1234), .Z
		(n_2078));
	notech_ao4 i_26678425(.A(n_58116), .B(n_42247), .C(n_58103), .D(n_42279)
		, .Z(n_2077));
	notech_ao4 i_25978432(.A(n_58142), .B(n_42199), .C(n_58129), .D(n_42207)
		, .Z(n_2075));
	notech_ao4 i_25778434(.A(n_58242), .B(n_42183), .C(n_58223), .D(n_42191)
		, .Z(n_2073));
	notech_ao4 i_23478457(.A(n_58194), .B(n_42270), .C(n_58181), .D(n_42262)
		, .Z(n_2070));
	notech_ao4 i_23378458(.A(n_58168), .B(n_42254), .C(n_58155), .D(n_42286)
		, .Z(n_2069));
	notech_and3 i_23678455(.A(n_2066), .B(n_2065), .C(n_1231), .Z(n_2068));
	notech_ao4 i_23078461(.A(n_58090), .B(n_42238), .C(n_58077), .D(n_42222)
		, .Z(n_2066));
	notech_ao4 i_22978462(.A(n_58064), .B(n_42214), .C(n_58051), .D(n_42230)
		, .Z(n_2065));
	notech_and4 i_23878453(.A(n_2059), .B(n_2061), .C(n_2063), .D(n_1218), .Z
		(n_2064));
	notech_ao4 i_23578456(.A(n_58116), .B(n_42246), .C(n_58103), .D(n_42278)
		, .Z(n_2063));
	notech_ao4 i_22878463(.A(n_58142), .B(n_42198), .C(n_58129), .D(n_42206)
		, .Z(n_2061));
	notech_ao4 i_22678465(.A(n_58242), .B(n_42182), .C(n_58223), .D(n_42190)
		, .Z(n_2059));
	notech_ao4 i_20378488(.A(n_58190), .B(n_42269), .C(n_58177), .D(n_42261)
		, .Z(n_2056));
	notech_ao4 i_20278489(.A(n_58164), .B(n_42253), .C(n_58151), .D(n_42285)
		, .Z(n_2055));
	notech_and3 i_20578486(.A(n_2052), .B(n_2051), .C(n_1215), .Z(n_2054));
	notech_ao4 i_19978492(.A(n_58086), .B(n_42237), .C(n_58073), .D(n_42221)
		, .Z(n_2052));
	notech_ao4 i_19878493(.A(n_58060), .B(n_42213), .C(n_58047), .D(n_42229)
		, .Z(n_2051));
	notech_and4 i_20778484(.A(n_2045), .B(n_2047), .C(n_2049), .D(n_1201), .Z
		(n_2050));
	notech_ao4 i_20478487(.A(n_58112), .B(n_42245), .C(n_58099), .D(n_42277)
		, .Z(n_2049));
	notech_ao4 i_19778494(.A(n_58138), .B(n_42197), .C(n_58125), .D(n_42205)
		, .Z(n_2047));
	notech_ao4 i_19578496(.A(n_58242), .B(n_42181), .C(n_58223), .D(n_42189)
		, .Z(n_2045));
	notech_ao4 i_17278519(.A(n_58190), .B(n_42268), .C(n_58177), .D(n_42260)
		, .Z(n_2042));
	notech_ao4 i_17178520(.A(n_58164), .B(n_42252), .C(n_58151), .D(n_42284)
		, .Z(n_2041));
	notech_and3 i_17478517(.A(n_2038), .B(n_2037), .C(n_1198), .Z(n_2040));
	notech_ao4 i_16878523(.A(n_58086), .B(n_42236), .C(n_58073), .D(n_42220)
		, .Z(n_2038));
	notech_ao4 i_16778524(.A(n_58060), .B(n_42212), .C(n_58047), .D(n_42228)
		, .Z(n_2037));
	notech_and4 i_17678515(.A(n_2031), .B(n_2033), .C(n_2035), .D(n_1185), .Z
		(n_2036));
	notech_ao4 i_17378518(.A(n_58112), .B(n_42244), .C(n_58099), .D(n_42276)
		, .Z(n_2035));
	notech_ao4 i_16678525(.A(n_58138), .B(n_42196), .C(n_58125), .D(n_42204)
		, .Z(n_2033));
	notech_ao4 i_16478527(.A(n_58242), .B(n_42180), .C(n_58223), .D(n_42188)
		, .Z(n_2031));
	notech_ao4 i_14178550(.A(n_58194), .B(n_42267), .C(n_58181), .D(n_42259)
		, .Z(n_2028));
	notech_ao4 i_14078551(.A(n_58168), .B(n_42251), .C(n_58155), .D(n_42283)
		, .Z(n_2027));
	notech_and3 i_14378548(.A(n_2024), .B(n_2023), .C(n_1182), .Z(n_2026));
	notech_ao4 i_13778554(.A(n_58090), .B(n_42235), .C(n_58077), .D(n_42219)
		, .Z(n_2024));
	notech_ao4 i_13678555(.A(n_58064), .B(n_42211), .C(n_58051), .D(n_42227)
		, .Z(n_2023));
	notech_and4 i_14578546(.A(n_2017), .B(n_2019), .C(n_2021), .D(n_1169), .Z
		(n_2022));
	notech_ao4 i_14278549(.A(n_58116), .B(n_42243), .C(n_58103), .D(n_42275)
		, .Z(n_2021));
	notech_ao4 i_13578556(.A(n_58142), .B(n_42195), .C(n_58129), .D(n_42203)
		, .Z(n_2019));
	notech_ao4 i_13378558(.A(n_58242), .B(n_42179), .C(n_58223), .D(n_42187)
		, .Z(n_2017));
	notech_ao4 i_11078581(.A(n_58194), .B(n_42266), .C(n_58181), .D(n_42258)
		, .Z(n_2014));
	notech_ao4 i_10978582(.A(n_58168), .B(n_42250), .C(n_58155), .D(n_42282)
		, .Z(n_2013));
	notech_and3 i_11278579(.A(n_2010), .B(n_2009), .C(n_1166), .Z(n_2012));
	notech_ao4 i_10678585(.A(n_58090), .B(n_42234), .C(n_58077), .D(n_42218)
		, .Z(n_2010));
	notech_ao4 i_10578586(.A(n_58064), .B(n_42210), .C(n_58051), .D(n_42226)
		, .Z(n_2009));
	notech_and4 i_11478577(.A(n_2003), .B(n_2005), .C(n_2007), .D(n_1153), .Z
		(n_2008));
	notech_ao4 i_11178580(.A(n_58116), .B(n_42242), .C(n_58103), .D(n_42274)
		, .Z(n_2007));
	notech_ao4 i_10478587(.A(n_58142), .B(n_42194), .C(n_58129), .D(n_42202)
		, .Z(n_2005));
	notech_ao4 i_10278589(.A(n_58242), .B(n_42178), .C(n_58223), .D(n_42186)
		, .Z(n_2003));
	notech_ao4 i_7878612(.A(n_58194), .B(n_42265), .C(n_58181), .D(n_42257),
		 .Z(n_2000));
	notech_nand3 i_1078673(.A(n_58211), .B(n_3070), .C(n_3064), .Z(n_1999)
		);
	notech_nand3 i_978674(.A(n_3070), .B(n_3066), .C(n_58211), .Z(n_1998));
	notech_ao4 i_7778613(.A(n_58168), .B(n_42249), .C(n_58155), .D(n_42281),
		 .Z(n_1997));
	notech_nand3 i_878675(.A(n_3064), .B(n_3061), .C(n_58211), .Z(n_1996));
	notech_nand3 i_478679(.A(n_3068), .B(n_3064), .C(n_58215), .Z(n_1995));
	notech_and3 i_8178610(.A(n_1992), .B(n_1989), .C(n_1150), .Z(n_1994));
	notech_ao4 i_7478616(.A(n_58090), .B(n_42233), .C(n_58077), .D(n_42217),
		 .Z(n_1992));
	notech_nand3 i_778676(.A(n_3078), .B(n_3064), .C(n_3083), .Z(n_1991));
	notech_nand3 i_678677(.A(n_3074), .B(n_3068), .C(n_3083), .Z(n_1990));
	notech_ao4 i_7378617(.A(n_58064), .B(n_42209), .C(n_58051), .D(n_42225),
		 .Z(n_1989));
	notech_nao3 i_578678(.A(n_3068), .B(n_3083), .C(n_3076), .Z(n_1988));
	notech_nand3 i_378680(.A(n_3078), .B(n_3066), .C(n_3083), .Z(n_1987));
	notech_and4 i_8378608(.A(n_1976), .B(n_1980), .C(n_1985), .D(n_113293395
		), .Z(n_1986));
	notech_ao4 i_7978611(.A(n_58116), .B(n_42241), .C(n_58103), .D(n_42273),
		 .Z(n_1985));
	notech_nand3 i_1278671(.A(n_3066), .B(n_58211), .C(n_3061), .Z(n_1984)
		);
	notech_nand3 i_1178672(.A(n_58215), .B(n_3068), .C(n_3066), .Z(n_1983)
		);
	notech_and4 i_1778666(.A(n_58371), .B(n_58355), .C(n_3080), .D(n_3083), 
		.Z(n_1982));
	notech_ao4 i_7278618(.A(n_58142), .B(n_42193), .C(n_58129), .D(n_42201),
		 .Z(n_1980));
	notech_nao3 i_178681(.A(n_3070), .B(n_3083), .C(n_3076), .Z(n_1979));
	notech_nand3 i_078682(.A(n_58379), .B(n_3070), .C(n_3083), .Z(n_1978));
	notech_ao4 i_6778620(.A(n_58242), .B(n_42177), .C(n_58223), .D(n_42185),
		 .Z(n_1976));
	notech_nand2 i_328403(.A(n_2706), .B(n_1974), .Z(n_35087));
	notech_or4 i_224376448(.A(n_61555), .B(n_60283), .C(n_60251), .D(n_42739
		), .Z(n_1974));
	notech_nand2 i_1128411(.A(n_2705), .B(n_1972), .Z(n_35135));
	notech_or4 i_221176480(.A(n_61555), .B(n_60283), .C(n_60251), .D(n_42738
		), .Z(n_1972));
	notech_nand2 i_1928419(.A(n_2704), .B(n_1970), .Z(n_35183));
	notech_or4 i_217976512(.A(n_61555), .B(n_60283), .C(n_60251), .D(n_42737
		), .Z(n_1970));
	notech_nand2 i_2728427(.A(n_2703), .B(n_1968), .Z(n_35231));
	notech_or4 i_214676545(.A(n_61555), .B(n_60283), .C(n_60251), .D(n_42736
		), .Z(n_1968));
	notech_and4 i_6625045(.A(n_2700), .B(n_2699), .C(n_2694), .D(n_2698), .Z
		(squeue_6597053));
	notech_nand3 i_162077071(.A(n_57940), .B(n_58215), .C(queue[65]), .Z(n_1967
		));
	notech_nand3 i_160777084(.A(n_3078), .B(n_58379), .C(queue[73]), .Z(n_1954
		));
	notech_and4 i_5425033(.A(n_2686), .B(n_2685), .C(n_2680), .D(n_2684), .Z
		(squeue_5397054));
	notech_nand3 i_158977102(.A(n_57940), .B(n_58211), .C(queue[53]), .Z(n_1951
		));
	notech_nand3 i_157677115(.A(n_60262), .B(n_58379), .C(queue[61]), .Z(n_1938
		));
	notech_and4 i_5325032(.A(n_2672), .B(n_2671), .C(n_2666), .D(n_2670), .Z
		(squeue_5297055));
	notech_nand3 i_155877133(.A(n_57940), .B(n_58211), .C(queue[52]), .Z(n_1935
		));
	notech_nand3 i_154577146(.A(n_60262), .B(n_58379), .C(queue[60]), .Z(n_1922
		));
	notech_and4 i_5225031(.A(n_2658), .B(n_2657), .C(n_2652), .D(n_2656), .Z
		(squeue_5197056));
	notech_nand3 i_152777164(.A(n_57940), .B(n_58211), .C(queue[51]), .Z(n_1919
		));
	notech_nand3 i_151477177(.A(n_60262), .B(n_58379), .C(queue[59]), .Z(n_1906
		));
	notech_and4 i_5125030(.A(n_2644), .B(n_2643), .C(n_2638), .D(n_2642), .Z
		(squeue_5097057));
	notech_nand3 i_149677195(.A(n_57940), .B(n_58211), .C(queue[50]), .Z(n_1903
		));
	notech_nand3 i_148377208(.A(n_60262), .B(n_58379), .C(queue[58]), .Z(n_1890
		));
	notech_and4 i_5025029(.A(n_2630), .B(n_2629), .C(n_2624), .D(n_2628), .Z
		(squeue_4997058));
	notech_nand3 i_146577226(.A(n_57940), .B(n_58216), .C(queue[49]), .Z(n_1887
		));
	notech_nand3 i_145277239(.A(n_60262), .B(n_3074), .C(queue[57]), .Z(n_1874
		));
	notech_and4 i_4925028(.A(n_2616), .B(n_2615), .C(n_2610), .D(n_2614), .Z
		(squeue_4897059));
	notech_nand3 i_143477257(.A(n_57940), .B(n_58218), .C(queue[48]), .Z(n_1871
		));
	notech_or2 i_142177270(.A(n_58242), .B(n_42225), .Z(n_1858));
	notech_and4 i_4825027(.A(n_2602), .B(n_2601), .C(n_2596), .D(n_2600), .Z
		(squeue_4797060));
	notech_nand3 i_140377288(.A(n_57940), .B(n_58218), .C(queue[47]), .Z(n_1855
		));
	notech_or2 i_139077301(.A(n_58274), .B(n_42216), .Z(n_1842));
	notech_and4 i_4725026(.A(n_2588), .B(n_2587), .C(n_2582), .D(n_2586), .Z
		(squeue_4697061));
	notech_nand3 i_137277319(.A(n_57940), .B(n_58218), .C(queue[46]), .Z(n_1839
		));
	notech_or2 i_135977332(.A(n_58274), .B(n_42215), .Z(n_1826));
	notech_and4 i_4625025(.A(n_2574), .B(n_2573), .C(n_2568), .D(n_2572), .Z
		(squeue_4597062));
	notech_nand3 i_134177350(.A(n_57940), .B(n_58218), .C(queue[45]), .Z(n_1823
		));
	notech_nand3 i_132877363(.A(n_60262), .B(n_3074), .C(queue[53]), .Z(n_1810
		));
	notech_and4 i_4525024(.A(n_2560), .B(n_2559), .C(n_2554), .D(n_2558), .Z
		(squeue_4497063));
	notech_nand3 i_131077381(.A(n_57947), .B(n_58218), .C(queue[44]), .Z(n_1807
		));
	notech_nand3 i_129777394(.A(n_3078), .B(n_3074), .C(queue[52]), .Z(n_1794
		));
	notech_and4 i_4425023(.A(n_2546), .B(n_2545), .C(n_2540), .D(n_2544), .Z
		(squeue_4397064));
	notech_nand3 i_127977412(.A(n_57947), .B(n_58218), .C(queue[43]), .Z(n_1791
		));
	notech_nand3 i_126677425(.A(n_3078), .B(n_3074), .C(queue[51]), .Z(n_1778
		));
	notech_and4 i_4325022(.A(n_2532), .B(n_2531), .C(n_2526), .D(n_2530), .Z
		(squeue_4297065));
	notech_nand3 i_124877443(.A(n_57947), .B(n_58218), .C(queue[42]), .Z(n_1775
		));
	notech_nand3 i_123577456(.A(n_3078), .B(n_3074), .C(queue[50]), .Z(n_1762
		));
	notech_and4 i_4225021(.A(n_2518), .B(n_2517), .C(n_2512), .D(n_2516), .Z
		(squeue_4197066));
	notech_nand3 i_121777474(.A(n_57947), .B(n_58218), .C(queue[41]), .Z(n_1759
		));
	notech_nand3 i_120477487(.A(n_3078), .B(n_3074), .C(queue[49]), .Z(n_1746
		));
	notech_and4 i_4125020(.A(n_2504), .B(n_2503), .C(n_2498), .D(n_2502), .Z
		(squeue_4097067));
	notech_nand3 i_118677505(.A(n_57947), .B(n_58218), .C(queue[40]), .Z(n_1743
		));
	notech_or2 i_117377518(.A(n_58223), .B(n_42225), .Z(n_1730));
	notech_and4 i_4025019(.A(n_2490), .B(n_2489), .C(n_2484), .D(n_2488), .Z
		(squeue_3997068));
	notech_nand3 i_115577536(.A(n_57947), .B(n_58218), .C(queue[39]), .Z(n_1727
		));
	notech_or2 i_114277549(.A(n_58274), .B(n_42208), .Z(n_1714));
	notech_and4 i_3925018(.A(n_2476), .B(n_2475), .C(n_2470), .D(n_2474), .Z
		(squeue_3897069));
	notech_nand3 i_112477567(.A(n_57947), .B(n_58218), .C(queue[38]), .Z(n_1711
		));
	notech_or2 i_111177580(.A(n_58274), .B(n_42207), .Z(n_1698));
	notech_and4 i_3725016(.A(n_2462), .B(n_2461), .C(n_2456), .D(n_2460), .Z
		(squeue_3697070));
	notech_nand3 i_109377598(.A(n_57947), .B(n_58218), .C(queue[36]), .Z(n_1695
		));
	notech_nand3 i_108077611(.A(n_3078), .B(n_3074), .C(queue[44]), .Z(n_1682
		));
	notech_and4 i_3625015(.A(n_2448), .B(n_2447), .C(n_2442), .D(n_2446), .Z
		(squeue_3597071));
	notech_nand3 i_106277629(.A(n_57947), .B(n_58218), .C(queue[35]), .Z(n_1679
		));
	notech_nand3 i_104977642(.A(n_3078), .B(n_3074), .C(queue[43]), .Z(n_1666
		));
	notech_and4 i_3525014(.A(n_2434), .B(n_2433), .C(n_2428), .D(n_2432), .Z
		(squeue_3497072));
	notech_nand3 i_103177660(.A(n_57947), .B(n_58218), .C(queue[34]), .Z(n_1663
		));
	notech_nand3 i_101877673(.A(n_3078), .B(n_3074), .C(queue[42]), .Z(n_1650
		));
	notech_and4 i_3425013(.A(n_2420), .B(n_2419), .C(n_2414), .D(n_2418), .Z
		(squeue_3397073));
	notech_nand3 i_100077691(.A(n_57947), .B(n_58218), .C(queue[33]), .Z(n_1647
		));
	notech_nand3 i_98777704(.A(n_3078), .B(n_3074), .C(queue[41]), .Z(n_1634
		));
	notech_and4 i_3325012(.A(n_2406), .B(n_2405), .C(n_2400), .D(n_2404), .Z
		(squeue_3297074));
	notech_nand3 i_96977722(.A(n_57947), .B(n_58218), .C(queue[32]), .Z(n_1631
		));
	notech_nand3 i_95677735(.A(n_3078), .B(n_3074), .C(queue[40]), .Z(n_1618
		));
	notech_and4 i_3225011(.A(n_2392), .B(n_2391), .C(n_2386), .D(n_2390), .Z
		(squeue_3197075));
	notech_nand3 i_93877753(.A(n_57947), .B(n_58218), .C(queue[31]), .Z(n_1615
		));
	notech_or2 i_28078943(.A(n_99694400), .B(n_307096441), .Z(n_99594399));
	notech_ao4 i_3579183(.A(n_60212), .B(n_309696467), .C(n_100494408), .D(n_100594409
		), .Z(n_99694400));
	notech_or4 i_27778946(.A(n_60003), .B(n_307096441), .C(n_42165), .D(n_42163
		), .Z(n_99894402));
	notech_nao3 i_27878945(.A(n_140853041), .B(pg_fault), .C(n_307096441), .Z
		(n_99994403));
	notech_ao3 i_28278941(.A(n_42165), .B(n_60251), .C(n_307096441), .Z(n_100094404
		));
	notech_nao3 i_46178762(.A(n_8288), .B(n_140853041), .C(pg_fault), .Z(n_100494408
		));
	notech_nand2 i_45978764(.A(n_34674), .B(n_42740), .Z(n_100594409));
	notech_nand2 i_7263(.A(n_34674), .B(n_42164), .Z(n_3855342));
	notech_nand2 i_2078663(.A(n_309596466), .B(n_8293), .Z(n_101094414));
	notech_nor2 i_6878687(.A(fault_wptr[1]), .B(fault_wptr[0]), .Z(n_7792)
		);
	notech_nao3 i_211485(.A(tagV[2]), .B(n_35018), .C(n_127594669), .Z(n_8288
		));
	notech_ao4 i_4578641(.A(n_127694670), .B(n_3855342), .C(n_309696467), .D
		(n_60212), .Z(n_101194415));
	notech_or2 i_7078685(.A(wptr[0]), .B(n_60283), .Z(n_7790));
	notech_or4 i_173676955(.A(n_61555), .B(n_60283), .C(n_60251), .D(n_42744
		), .Z(n_101494418));
	notech_nand2 i_12728527(.A(n_127794671), .B(n_101494418), .Z(n_35831));
	notech_or4 i_174476947(.A(n_61555), .B(n_60283), .C(n_60251), .D(n_42745
		), .Z(n_101694420));
	notech_nand2 i_12528525(.A(n_127894672), .B(n_101694420), .Z(n_35819));
	notech_or4 i_174876943(.A(n_61555), .B(n_60283), .C(n_60251), .D(n_42746
		), .Z(n_101894422));
	notech_nand2 i_12428524(.A(n_127994673), .B(n_101894422), .Z(n_35813));
	notech_or4 i_175276939(.A(n_61555), .B(n_60283), .C(n_60251), .D(n_42747
		), .Z(n_102094424));
	notech_nand2 i_12328523(.A(n_128094674), .B(n_102094424), .Z(n_35807));
	notech_or4 i_175676935(.A(n_61556), .B(n_60284), .C(n_60251), .D(n_42748
		), .Z(n_102294426));
	notech_nand2 i_12228522(.A(n_128194675), .B(n_102294426), .Z(n_35801));
	notech_or4 i_176076931(.A(n_61556), .B(n_60284), .C(n_60252), .D(n_42749
		), .Z(n_102494428));
	notech_nand2 i_12128521(.A(n_128294676), .B(n_102494428), .Z(n_35795));
	notech_or4 i_176476927(.A(n_61556), .B(n_60283), .C(n_60252), .D(n_42750
		), .Z(n_102694430));
	notech_nand2 i_12028520(.A(n_128394677), .B(n_102694430), .Z(n_35789));
	notech_or4 i_176876923(.A(n_61556), .B(n_60283), .C(n_60251), .D(n_42751
		), .Z(n_102894432));
	notech_nand2 i_11928519(.A(n_128494678), .B(n_102894432), .Z(n_35783));
	notech_or4 i_177276919(.A(n_61555), .B(n_60283), .C(n_60251), .D(n_42752
		), .Z(n_103094434));
	notech_nand2 i_11828518(.A(n_128594679), .B(n_103094434), .Z(n_35777));
	notech_or4 i_177676915(.A(n_61555), .B(n_60283), .C(n_60251), .D(n_42753
		), .Z(n_103294436));
	notech_nand2 i_11728517(.A(n_128794680), .B(n_103294436), .Z(n_35771));
	notech_or4 i_178076911(.A(n_61555), .B(n_60283), .C(n_60251), .D(n_42754
		), .Z(n_103494438));
	notech_nand2 i_11628516(.A(n_128894681), .B(n_103494438), .Z(n_35765));
	notech_or4 i_178476907(.A(n_61555), .B(n_60279), .C(n_60251), .D(n_42755
		), .Z(n_103694440));
	notech_nand2 i_11528515(.A(n_128994682), .B(n_103694440), .Z(n_35759));
	notech_or4 i_178876903(.A(n_61555), .B(n_60279), .C(n_60247), .D(n_42756
		), .Z(n_103894442));
	notech_nand2 i_11428514(.A(n_129394683), .B(n_103894442), .Z(n_35753));
	notech_or4 i_179276899(.A(n_61551), .B(n_60279), .C(n_60247), .D(n_42757
		), .Z(n_104094444));
	notech_nand2 i_11328513(.A(n_129494684), .B(n_104094444), .Z(n_35747));
	notech_or4 i_179676895(.A(n_61551), .B(n_60279), .C(n_60247), .D(n_42758
		), .Z(n_104294446));
	notech_nand2 i_11228512(.A(n_129594685), .B(n_104294446), .Z(n_35741));
	notech_or4 i_180076891(.A(n_61551), .B(n_60279), .C(n_60247), .D(n_42759
		), .Z(n_104494448));
	notech_nand2 i_11128511(.A(n_129894686), .B(n_104494448), .Z(n_35735));
	notech_or4 i_180476887(.A(n_61551), .B(n_60279), .C(n_60247), .D(n_42760
		), .Z(n_104694450));
	notech_nand2 i_11028510(.A(n_129994687), .B(n_104694450), .Z(n_35729));
	notech_or4 i_180876883(.A(n_61551), .B(n_60279), .C(n_60247), .D(n_42761
		), .Z(n_104894452));
	notech_nand2 i_10928509(.A(n_130294688), .B(n_104894452), .Z(n_35723));
	notech_or4 i_181276879(.A(n_61551), .B(n_60279), .C(n_60247), .D(n_42762
		), .Z(n_105094454));
	notech_nand2 i_10828508(.A(n_130394689), .B(n_105094454), .Z(n_35717));
	notech_or4 i_181676875(.A(n_61551), .B(n_60283), .C(n_60247), .D(n_42763
		), .Z(n_105294456));
	notech_nand2 i_10728507(.A(n_130694690), .B(n_105294456), .Z(n_35711));
	notech_or4 i_182076871(.A(n_61551), .B(n_60279), .C(n_60251), .D(n_42764
		), .Z(n_105494458));
	notech_nand2 i_10628506(.A(n_130794691), .B(n_105494458), .Z(n_35705));
	notech_or4 i_182476867(.A(n_61555), .B(n_60283), .C(n_60247), .D(n_42765
		), .Z(n_105694460));
	notech_nand2 i_10528505(.A(n_130894692), .B(n_105694460), .Z(n_35699));
	notech_or4 i_182876863(.A(n_61555), .B(n_60283), .C(n_60251), .D(n_42766
		), .Z(n_105894462));
	notech_nand2 i_10428504(.A(n_130994693), .B(n_105894462), .Z(n_35693));
	notech_or4 i_183276859(.A(n_61555), .B(n_60279), .C(n_60251), .D(n_42767
		), .Z(n_106094464));
	notech_nand2 i_10328503(.A(n_131294694), .B(n_106094464), .Z(n_35687));
	notech_or4 i_183676855(.A(n_61555), .B(n_60279), .C(n_60247), .D(n_42768
		), .Z(n_106294466));
	notech_nand2 i_10228502(.A(n_131394695), .B(n_106294466), .Z(n_35681));
	notech_or4 i_184076851(.A(n_61551), .B(n_60279), .C(n_60247), .D(n_42769
		), .Z(n_106494468));
	notech_nand2 i_10128501(.A(n_131694696), .B(n_106494468), .Z(n_35675));
	notech_or4 i_184576846(.A(n_61551), .B(n_60279), .C(n_60247), .D(n_42770
		), .Z(n_106794471));
	notech_nand2 i_10028500(.A(n_131794697), .B(n_106794471), .Z(n_35669));
	notech_or4 i_184976842(.A(n_61555), .B(n_60284), .C(n_60247), .D(n_42771
		), .Z(n_106994473));
	notech_nand2 i_9928499(.A(n_131994698), .B(n_106994473), .Z(n_35663));
	notech_or4 i_185376838(.A(n_61551), .B(n_60286), .C(n_60252), .D(n_42772
		), .Z(n_107194475));
	notech_nand2 i_9828498(.A(n_132094699), .B(n_107194475), .Z(n_35657));
	notech_or4 i_185876833(.A(n_61556), .B(n_60286), .C(n_60254), .D(n_42773
		), .Z(n_107494478));
	notech_nand2 i_9728497(.A(n_132294700), .B(n_107494478), .Z(n_35651));
	notech_or4 i_186276829(.A(n_61558), .B(n_60286), .C(n_60254), .D(n_42774
		), .Z(n_107694480));
	notech_nand2 i_9628496(.A(n_132394701), .B(n_107694480), .Z(n_35645));
	notech_or4 i_186776824(.A(n_61558), .B(n_60286), .C(n_60254), .D(n_42775
		), .Z(n_107994483));
	notech_nand2 i_9528495(.A(n_132494702), .B(n_107994483), .Z(n_35639));
	notech_or4 i_187276819(.A(n_61558), .B(n_60286), .C(n_60254), .D(n_42776
		), .Z(n_108294486));
	notech_nand2 i_9428494(.A(n_132594703), .B(n_108294486), .Z(n_35633));
	notech_or4 i_187676815(.A(n_61558), .B(n_60286), .C(n_60254), .D(n_42777
		), .Z(n_108494488));
	notech_nand2 i_9328493(.A(n_132694704), .B(n_108494488), .Z(n_35627));
	notech_or4 i_188176810(.A(n_61558), .B(n_60286), .C(n_60254), .D(n_42778
		), .Z(n_108794491));
	notech_nand2 i_9228492(.A(n_132794705), .B(n_108794491), .Z(n_35621));
	notech_or4 i_188676805(.A(n_61558), .B(n_60286), .C(n_60254), .D(n_42779
		), .Z(n_109094494));
	notech_nand2 i_9128491(.A(n_132894706), .B(n_109094494), .Z(n_35615));
	notech_or4 i_189176800(.A(n_61558), .B(n_60286), .C(n_60254), .D(n_42780
		), .Z(n_109394497));
	notech_nand2 i_9028490(.A(n_132994707), .B(n_109394497), .Z(n_35609));
	notech_or4 i_190176790(.A(n_61558), .B(n_60286), .C(n_60254), .D(n_42781
		), .Z(n_109694500));
	notech_nand2 i_8828488(.A(n_133094708), .B(n_109694500), .Z(n_35597));
	notech_or4 i_190676785(.A(n_61558), .B(n_60286), .C(n_60254), .D(n_42782
		), .Z(n_109994503));
	notech_nand2 i_8728487(.A(n_133194709), .B(n_109994503), .Z(n_35591));
	notech_or4 i_191076781(.A(n_61558), .B(n_60286), .C(n_60254), .D(n_42783
		), .Z(n_110194505));
	notech_nand2 i_8628486(.A(n_133294710), .B(n_110194505), .Z(n_35585));
	notech_or4 i_191476777(.A(n_61558), .B(n_60286), .C(n_60254), .D(n_42784
		), .Z(n_110394507));
	notech_nand2 i_8528485(.A(n_133394711), .B(n_110394507), .Z(n_35579));
	notech_or4 i_191876773(.A(n_61558), .B(n_60286), .C(n_60254), .D(n_42785
		), .Z(n_110594509));
	notech_nand2 i_8428484(.A(n_133494712), .B(n_110594509), .Z(n_35573));
	notech_or4 i_192276769(.A(n_61558), .B(n_60286), .C(n_60254), .D(n_42786
		), .Z(n_110794511));
	notech_nand2 i_8328483(.A(n_133594713), .B(n_110794511), .Z(n_35567));
	notech_or4 i_192676765(.A(n_61558), .B(n_60286), .C(n_60254), .D(n_42787
		), .Z(n_110994513));
	notech_nand2 i_8228482(.A(n_133694714), .B(n_110994513), .Z(n_35561));
	notech_or4 i_193076761(.A(n_61558), .B(n_60286), .C(n_60254), .D(n_42788
		), .Z(n_111194515));
	notech_nand2 i_8128481(.A(n_133794715), .B(n_111194515), .Z(n_35555));
	notech_or4 i_193476757(.A(n_61558), .B(n_60284), .C(n_60254), .D(n_42789
		), .Z(n_111394517));
	notech_nand2 i_8028480(.A(n_133894716), .B(n_111394517), .Z(n_35549));
	notech_or4 i_193876753(.A(n_61558), .B(n_60284), .C(n_60252), .D(n_42790
		), .Z(n_111594519));
	notech_nand2 i_7928479(.A(n_133994717), .B(n_111594519), .Z(n_35543));
	notech_or4 i_194276749(.A(n_61556), .B(n_60284), .C(n_60252), .D(n_42791
		), .Z(n_111894521));
	notech_nand2 i_7828478(.A(n_134094718), .B(n_111894521), .Z(n_35537));
	notech_or4 i_194676745(.A(n_61556), .B(n_60284), .C(n_60252), .D(n_42792
		), .Z(n_112294523));
	notech_nand2 i_7728477(.A(n_134194719), .B(n_112294523), .Z(n_35531));
	notech_or4 i_195076741(.A(n_61556), .B(n_60284), .C(n_60252), .D(n_42793
		), .Z(n_112494525));
	notech_nand2 i_7628476(.A(n_134294720), .B(n_112494525), .Z(n_35525));
	notech_or4 i_195476737(.A(n_61556), .B(n_60284), .C(n_60252), .D(n_42794
		), .Z(n_112694526));
	notech_nand2 i_7528475(.A(n_134394721), .B(n_112694526), .Z(n_35519));
	notech_or4 i_195876733(.A(n_61556), .B(n_60284), .C(n_60252), .D(n_42795
		), .Z(n_112894528));
	notech_nand2 i_7428474(.A(n_134494722), .B(n_112894528), .Z(n_35513));
	notech_or4 i_196276729(.A(n_61556), .B(n_60284), .C(n_60252), .D(n_42796
		), .Z(n_113094530));
	notech_nand2 i_7328473(.A(n_134594723), .B(n_113094530), .Z(n_35507));
	notech_or4 i_196676725(.A(n_61556), .B(n_60284), .C(n_60252), .D(n_42797
		), .Z(n_113294532));
	notech_nand2 i_7228472(.A(n_134694724), .B(n_113294532), .Z(n_35501));
	notech_or4 i_197476717(.A(n_61556), .B(n_60284), .C(n_60252), .D(n_42798
		), .Z(n_113494534));
	notech_nand2 i_7028470(.A(n_134794725), .B(n_113494534), .Z(n_35489));
	notech_or4 i_197876713(.A(n_61558), .B(n_60286), .C(n_60252), .D(n_42799
		), .Z(n_113794536));
	notech_nand2 i_6928469(.A(n_134894726), .B(n_113794536), .Z(n_35483));
	notech_or4 i_198276709(.A(n_61556), .B(n_60284), .C(n_60254), .D(n_42800
		), .Z(n_114294538));
	notech_nand2 i_6828468(.A(n_134994727), .B(n_114294538), .Z(n_35477));
	notech_or4 i_198676705(.A(n_61558), .B(n_60284), .C(n_60252), .D(n_42801
		), .Z(n_114494540));
	notech_nand2 i_6728467(.A(n_135094728), .B(n_114494540), .Z(n_35471));
	notech_or4 i_199076701(.A(n_61558), .B(n_60284), .C(n_60252), .D(n_42802
		), .Z(n_114694542));
	notech_nand2 i_6628466(.A(n_135194729), .B(n_114694542), .Z(n_35465));
	notech_or4 i_199476697(.A(n_61556), .B(n_60284), .C(n_60252), .D(n_42803
		), .Z(n_114894544));
	notech_nand2 i_6528465(.A(n_135294730), .B(n_114894544), .Z(n_35459));
	notech_or4 i_199876693(.A(n_61556), .B(n_60284), .C(n_60252), .D(n_42804
		), .Z(n_115094546));
	notech_nand2 i_6428464(.A(n_135394731), .B(n_115094546), .Z(n_35453));
	notech_or4 i_200276689(.A(n_61556), .B(n_60272), .C(n_60252), .D(n_42805
		), .Z(n_115294548));
	notech_nand2 i_6328463(.A(n_135494732), .B(n_115294548), .Z(n_35447));
	notech_or4 i_200676685(.A(n_61556), .B(n_60272), .C(n_60247), .D(n_42806
		), .Z(n_115494550));
	notech_nand2 i_6228462(.A(n_135594733), .B(n_115494550), .Z(n_35441));
	notech_or4 i_201076681(.A(n_61544), .B(n_60272), .C(n_60241), .D(n_42807
		), .Z(n_115694552));
	notech_nand2 i_6128461(.A(n_135694734), .B(n_115694552), .Z(n_35435));
	notech_or4 i_201476677(.A(n_61544), .B(n_60272), .C(n_60241), .D(n_42808
		), .Z(n_115894554));
	notech_nand2 i_6028460(.A(n_135794735), .B(n_115894554), .Z(n_35429));
	notech_or4 i_202276669(.A(n_61546), .B(n_60272), .C(n_60241), .D(n_42809
		), .Z(n_116094556));
	notech_nand2 i_5828458(.A(n_135894736), .B(n_116094556), .Z(n_35417));
	notech_or4 i_202676665(.A(n_61546), .B(n_60272), .C(n_60241), .D(n_42810
		), .Z(n_116294558));
	notech_nand2 i_5728457(.A(n_135994737), .B(n_116294558), .Z(n_35411));
	notech_or4 i_203076661(.A(n_61544), .B(n_60272), .C(n_60241), .D(n_42811
		), .Z(n_116494560));
	notech_nand2 i_5628456(.A(n_136094738), .B(n_116494560), .Z(n_35405));
	notech_or4 i_203476657(.A(n_61544), .B(n_60272), .C(n_60239), .D(n_42812
		), .Z(n_116694562));
	notech_nand2 i_5528455(.A(n_136194739), .B(n_116694562), .Z(n_35399));
	notech_or4 i_203876653(.A(n_61544), .B(n_60274), .C(n_60241), .D(n_42813
		), .Z(n_116894564));
	notech_nand2 i_5428454(.A(n_136294740), .B(n_116894564), .Z(n_35393));
	notech_or4 i_204276649(.A(n_61544), .B(n_60274), .C(n_60241), .D(n_42814
		), .Z(n_117094566));
	notech_nand2 i_5328453(.A(n_136394741), .B(n_117094566), .Z(n_35387));
	notech_or4 i_204676645(.A(n_61546), .B(n_60274), .C(n_60241), .D(n_42815
		), .Z(n_117294568));
	notech_nand2 i_5228452(.A(n_136494742), .B(n_117294568), .Z(n_35381));
	notech_or4 i_205076641(.A(n_61546), .B(n_60274), .C(n_60241), .D(n_42816
		), .Z(n_117494570));
	notech_nand2 i_5128451(.A(n_136594743), .B(n_117494570), .Z(n_35375));
	notech_or4 i_205476637(.A(n_61546), .B(n_60274), .C(n_60241), .D(n_42817
		), .Z(n_117694572));
	notech_nand2 i_5028450(.A(n_136694744), .B(n_117694572), .Z(n_35369));
	notech_or4 i_205876633(.A(n_61546), .B(n_60272), .C(n_60241), .D(n_42818
		), .Z(n_117894574));
	notech_nand2 i_4928449(.A(n_136794745), .B(n_117894574), .Z(n_35363));
	notech_or4 i_206276629(.A(n_61546), .B(n_60274), .C(n_60241), .D(n_42819
		), .Z(n_118094576));
	notech_nand2 i_4828448(.A(n_136894746), .B(n_118094576), .Z(n_35357));
	notech_or4 i_206676625(.A(n_61546), .B(n_60274), .C(n_60241), .D(n_42820
		), .Z(n_118294578));
	notech_nand2 i_4728447(.A(n_136994747), .B(n_118294578), .Z(n_35351));
	notech_or4 i_207076621(.A(n_61546), .B(n_60272), .C(n_60241), .D(n_42821
		), .Z(n_118494580));
	notech_nand2 i_4628446(.A(n_137094748), .B(n_118494580), .Z(n_35345));
	notech_or4 i_207476617(.A(n_61546), .B(n_60271), .C(n_60241), .D(n_42822
		), .Z(n_118694582));
	notech_nand2 i_4528445(.A(n_137194749), .B(n_118694582), .Z(n_35339));
	notech_or4 i_207876613(.A(n_61544), .B(n_60271), .C(n_60239), .D(n_42823
		), .Z(n_118894584));
	notech_nand2 i_4428444(.A(n_137294750), .B(n_118894584), .Z(n_35333));
	notech_or4 i_208276609(.A(n_61544), .B(n_60271), .C(n_60239), .D(n_42824
		), .Z(n_119094586));
	notech_nand2 i_4328443(.A(n_137394751), .B(n_119094586), .Z(n_35327));
	notech_or4 i_208676605(.A(code_req), .B(n_60271), .C(n_60239), .D(n_42825
		), .Z(n_119294588));
	notech_nand2 i_4228442(.A(n_137494752), .B(n_119294588), .Z(n_35321));
	notech_or4 i_209076601(.A(n_61544), .B(n_60271), .C(n_60239), .D(n_42826
		), .Z(n_119494590));
	notech_nand2 i_4128441(.A(n_137594753), .B(n_119494590), .Z(n_35315));
	notech_or4 i_209476597(.A(n_61544), .B(n_60271), .C(n_60239), .D(n_42827
		), .Z(n_119694592));
	notech_nand2 i_4028440(.A(n_137694754), .B(n_119694592), .Z(n_35309));
	notech_or4 i_209876593(.A(code_req), .B(n_60271), .C(n_60239), .D(n_42828
		), .Z(n_119894594));
	notech_nand2 i_3928439(.A(n_137794755), .B(n_119894594), .Z(n_35303));
	notech_or4 i_210276589(.A(code_req), .B(n_60271), .C(n_60239), .D(n_42829
		), .Z(n_120094596));
	notech_nand2 i_3828438(.A(n_137894756), .B(n_120094596), .Z(n_35297));
	notech_or4 i_210676585(.A(code_req), .B(n_60272), .C(n_60239), .D(n_42830
		), .Z(n_120294598));
	notech_nand2 i_3728437(.A(n_137994757), .B(n_120294598), .Z(n_35291));
	notech_or4 i_211076581(.A(code_req), .B(n_60272), .C(n_60239), .D(n_42831
		), .Z(n_120494600));
	notech_nand2 i_3628436(.A(n_138094758), .B(n_120494600), .Z(n_35285));
	notech_or4 i_211476577(.A(n_61544), .B(n_60272), .C(n_60239), .D(n_42832
		), .Z(n_120694602));
	notech_nand2 i_3528435(.A(n_138194759), .B(n_120694602), .Z(n_35279));
	notech_or4 i_211876573(.A(n_61544), .B(n_60272), .C(n_60239), .D(n_42833
		), .Z(n_120894604));
	notech_nand2 i_3428434(.A(n_138294760), .B(n_120894604), .Z(n_35273));
	notech_or4 i_212276569(.A(n_61544), .B(n_60272), .C(n_60239), .D(n_42834
		), .Z(n_121094606));
	notech_nand2 i_3328433(.A(n_138394761), .B(n_121094606), .Z(n_35267));
	notech_or4 i_212676565(.A(n_61544), .B(n_60272), .C(n_60239), .D(n_42835
		), .Z(n_121394608));
	notech_nand2 i_3228432(.A(n_138494762), .B(n_121394608), .Z(n_35261));
	notech_or4 i_213076561(.A(n_61544), .B(n_60272), .C(n_60239), .D(n_42836
		), .Z(n_121594610));
	notech_nand2 i_3128431(.A(n_138594763), .B(n_121594610), .Z(n_35255));
	notech_or4 i_213476557(.A(n_61544), .B(n_60272), .C(n_60239), .D(n_42837
		), .Z(n_121794611));
	notech_nand2 i_3028430(.A(n_138694764), .B(n_121794611), .Z(n_35249));
	notech_or4 i_213876553(.A(n_61544), .B(n_60274), .C(n_60239), .D(n_42838
		), .Z(n_121994613));
	notech_nand2 i_2928429(.A(n_138794765), .B(n_121994613), .Z(n_35243));
	notech_or4 i_214276549(.A(n_61544), .B(n_60277), .C(n_60239), .D(n_42839
		), .Z(n_122194615));
	notech_nand2 i_2828428(.A(n_138894766), .B(n_122194615), .Z(n_35237));
	notech_or4 i_215076541(.A(n_61549), .B(n_60277), .C(n_60241), .D(n_42840
		), .Z(n_122394617));
	notech_nand2 i_2628426(.A(n_138994767), .B(n_122394617), .Z(n_35225));
	notech_or4 i_215476537(.A(n_61549), .B(n_60277), .C(n_60245), .D(n_42841
		), .Z(n_122594619));
	notech_nand2 i_2528425(.A(n_139094768), .B(n_122594619), .Z(n_35219));
	notech_or4 i_215876533(.A(n_61549), .B(n_60277), .C(n_60245), .D(n_42842
		), .Z(n_122794621));
	notech_nand2 i_2428424(.A(n_139194769), .B(n_122794621), .Z(n_35213));
	notech_or4 i_216276529(.A(n_61549), .B(n_60277), .C(n_60245), .D(n_42843
		), .Z(n_122994623));
	notech_nand2 i_2328423(.A(n_139294770), .B(n_122994623), .Z(n_35207));
	notech_or4 i_216676525(.A(n_61549), .B(n_60277), .C(n_60245), .D(n_42844
		), .Z(n_123194625));
	notech_nand2 i_2228422(.A(n_139394771), .B(n_123194625), .Z(n_35201));
	notech_or4 i_217076521(.A(n_61549), .B(n_60277), .C(n_60245), .D(n_42845
		), .Z(n_123394627));
	notech_nand2 i_2128421(.A(n_139494772), .B(n_123394627), .Z(n_35195));
	notech_or4 i_217576516(.A(n_61549), .B(n_60277), .C(n_60245), .D(n_42846
		), .Z(n_123694630));
	notech_nand2 i_2028420(.A(n_139594773), .B(n_123694630), .Z(n_35189));
	notech_or4 i_218376508(.A(n_61549), .B(n_60279), .C(n_60245), .D(n_42847
		), .Z(n_123894632));
	notech_nand2 i_1828418(.A(n_139694774), .B(n_123894632), .Z(n_35177));
	notech_or4 i_218776504(.A(n_61551), .B(n_60279), .C(n_60245), .D(n_42848
		), .Z(n_124094634));
	notech_nand2 i_1728417(.A(n_139794775), .B(n_124094634), .Z(n_35171));
	notech_or4 i_219176500(.A(n_61551), .B(n_60279), .C(n_60247), .D(n_42849
		), .Z(n_124294636));
	notech_nand2 i_1628416(.A(n_139894776), .B(n_124294636), .Z(n_35165));
	notech_or4 i_219576496(.A(n_61551), .B(n_60279), .C(n_60247), .D(n_42850
		), .Z(n_124494638));
	notech_nand2 i_1528415(.A(n_139994777), .B(n_124494638), .Z(n_35159));
	notech_or4 i_219976492(.A(n_61551), .B(n_60277), .C(n_60247), .D(n_42851
		), .Z(n_124694640));
	notech_nand2 i_1428414(.A(n_140094778), .B(n_124694640), .Z(n_35153));
	notech_or4 i_220376488(.A(n_61551), .B(n_60277), .C(n_60247), .D(n_42852
		), .Z(n_124894642));
	notech_nand2 i_1328413(.A(n_140194779), .B(n_124894642), .Z(n_35147));
	notech_or4 i_220776484(.A(n_61549), .B(n_60279), .C(n_60245), .D(n_42853
		), .Z(n_125094644));
	notech_nand2 i_1228412(.A(n_140294780), .B(n_125094644), .Z(n_35141));
	notech_or4 i_221576476(.A(n_61551), .B(n_60277), .C(n_60245), .D(n_42854
		), .Z(n_125294646));
	notech_nand2 i_1028410(.A(n_140394781), .B(n_125294646), .Z(n_35129));
	notech_or4 i_221976472(.A(n_61551), .B(n_60277), .C(n_60245), .D(n_42855
		), .Z(n_125494648));
	notech_nand2 i_928409(.A(n_140494782), .B(n_125494648), .Z(n_35123));
	notech_or4 i_222376468(.A(n_61549), .B(n_60274), .C(n_60245), .D(n_42856
		), .Z(n_125694650));
	notech_nand2 i_828408(.A(n_140594783), .B(n_125694650), .Z(n_35117));
	notech_or4 i_222776464(.A(n_61546), .B(n_60274), .C(n_60245), .D(n_42857
		), .Z(n_125894652));
	notech_nand2 i_728407(.A(n_140694784), .B(n_125894652), .Z(n_35111));
	notech_or4 i_223176460(.A(n_61546), .B(n_60274), .C(n_60243), .D(n_42858
		), .Z(n_126094654));
	notech_nand2 i_628406(.A(n_140794785), .B(n_126094654), .Z(n_35105));
	notech_or4 i_223576456(.A(n_61546), .B(n_60274), .C(n_60243), .D(n_42859
		), .Z(n_126294656));
	notech_nand2 i_528405(.A(n_140894786), .B(n_126294656), .Z(n_35099));
	notech_or4 i_223976452(.A(n_61546), .B(n_60274), .C(n_60243), .D(n_42860
		), .Z(n_126494658));
	notech_nand2 i_428404(.A(n_140994787), .B(n_126494658), .Z(n_35093));
	notech_or4 i_224776444(.A(n_61546), .B(n_60274), .C(n_60243), .D(n_42861
		), .Z(n_126694660));
	notech_nand2 i_228402(.A(n_141094788), .B(n_126694660), .Z(n_35081));
	notech_or4 i_225176440(.A(n_61546), .B(n_60274), .C(n_60241), .D(n_42862
		), .Z(n_126894662));
	notech_nand2 i_128401(.A(n_141194789), .B(n_126894662), .Z(n_35075));
	notech_and2 i_1678667(.A(n_42743), .B(n_42170), .Z(n_141953052));
	notech_or4 i_4378643(.A(tagV[1]), .B(tagV[0]), .C(tagV[3]), .D(purge), .Z
		(n_127594669));
	notech_or4 i_1878665(.A(n_61546), .B(pg_fault), .C(n_60274), .D(n_60241)
		, .Z(n_127694670));
	notech_ao4 i_173876953(.A(n_60212), .B(n_42729), .C(n_60003), .D(n_42543
		), .Z(n_127794671));
	notech_ao4 i_174676945(.A(n_60212), .B(n_42727), .C(n_60003), .D(n_42539
		), .Z(n_127894672));
	notech_ao4 i_175076941(.A(n_60182), .B(n_42726), .C(n_60003), .D(n_42537
		), .Z(n_127994673));
	notech_ao4 i_175476937(.A(n_60182), .B(n_42725), .C(n_60003), .D(n_42535
		), .Z(n_128094674));
	notech_ao4 i_175876933(.A(n_60182), .B(n_42724), .C(n_60007), .D(n_42533
		), .Z(n_128194675));
	notech_ao4 i_176276929(.A(n_60182), .B(n_42723), .C(n_60007), .D(n_42531
		), .Z(n_128294676));
	notech_ao4 i_176676925(.A(n_60182), .B(n_42722), .C(n_60007), .D(n_42529
		), .Z(n_128394677));
	notech_ao4 i_177076921(.A(n_60212), .B(n_42721), .C(n_60007), .D(n_42527
		), .Z(n_128494678));
	notech_ao4 i_177476917(.A(n_60182), .B(n_42720), .C(n_60007), .D(n_42525
		), .Z(n_128594679));
	notech_ao4 i_177876913(.A(n_60182), .B(n_42719), .C(n_60007), .D(n_42523
		), .Z(n_128794680));
	notech_ao4 i_178276909(.A(n_60216), .B(n_42718), .C(n_60007), .D(n_42521
		), .Z(n_128894681));
	notech_ao4 i_178676905(.A(n_60216), .B(n_42717), .C(n_60007), .D(n_42519
		), .Z(n_128994682));
	notech_ao4 i_179076901(.A(n_60216), .B(n_42716), .C(n_60001), .D(n_42517
		), .Z(n_129394683));
	notech_ao4 i_179476897(.A(n_60216), .B(n_42715), .C(n_60001), .D(n_42515
		), .Z(n_129494684));
	notech_ao4 i_179876893(.A(n_60216), .B(n_42714), .C(n_60001), .D(n_42513
		), .Z(n_129594685));
	notech_ao4 i_180276889(.A(n_60216), .B(n_42713), .C(n_60001), .D(n_42511
		), .Z(n_129894686));
	notech_ao4 i_180676885(.A(n_60216), .B(n_42712), .C(n_60001), .D(n_42509
		), .Z(n_129994687));
	notech_ao4 i_181076881(.A(n_60216), .B(n_42711), .C(n_60001), .D(n_42507
		), .Z(n_130294688));
	notech_ao4 i_181476877(.A(n_60212), .B(n_42710), .C(n_60001), .D(n_42505
		), .Z(n_130394689));
	notech_ao4 i_181876873(.A(n_60212), .B(n_42709), .C(n_60001), .D(n_42503
		), .Z(n_130694690));
	notech_ao4 i_182276869(.A(n_60212), .B(n_42708), .C(n_60001), .D(n_42501
		), .Z(n_130794691));
	notech_ao4 i_182676865(.A(n_60212), .B(n_42707), .C(n_60003), .D(n_42499
		), .Z(n_130894692));
	notech_ao4 i_183076861(.A(n_60216), .B(n_42706), .C(n_60003), .D(n_42497
		), .Z(n_130994693));
	notech_ao4 i_183476857(.A(n_60216), .B(n_42705), .C(n_60003), .D(n_42495
		), .Z(n_131294694));
	notech_ao4 i_183876853(.A(n_60212), .B(n_42704), .C(n_60003), .D(n_42493
		), .Z(n_131394695));
	notech_ao4 i_184376848(.A(n_60001), .B(n_42491), .C(n_60212), .D(n_42703
		), .Z(n_131694696));
	notech_ao4 i_184776844(.A(n_60202), .B(n_42702), .C(n_60001), .D(n_42489
		), .Z(n_131794697));
	notech_ao4 i_185176840(.A(n_60202), .B(n_42701), .C(n_60003), .D(n_42487
		), .Z(n_131994698));
	notech_ao4 i_185676835(.A(n_60001), .B(n_42485), .C(n_60197), .D(n_42700
		), .Z(n_132094699));
	notech_ao4 i_186076831(.A(n_60202), .B(n_42699), .C(n_60010), .D(n_42483
		), .Z(n_132294700));
	notech_ao4 i_186576826(.A(n_60010), .B(n_42481), .C(n_60202), .D(n_42698
		), .Z(n_132394701));
	notech_ao4 i_187076821(.A(n_60010), .B(n_42479), .C(n_60202), .D(n_42697
		), .Z(n_132494702));
	notech_ao4 i_187476817(.A(n_60202), .B(n_42696), .C(n_60010), .D(n_42477
		), .Z(n_132594703));
	notech_ao4 i_187976812(.A(n_60008), .B(n_42475), .C(n_60202), .D(n_42695
		), .Z(n_132694704));
	notech_ao4 i_188476807(.A(n_60008), .B(n_42473), .C(n_60197), .D(n_42694
		), .Z(n_132794705));
	notech_ao4 i_188976802(.A(n_60010), .B(n_42471), .C(n_60197), .D(n_42693
		), .Z(n_132894706));
	notech_ao4 i_189476797(.A(n_60008), .B(n_42469), .C(n_60197), .D(n_42692
		), .Z(n_132994707));
	notech_ao4 i_190476787(.A(n_60010), .B(n_42465), .C(n_60197), .D(n_42690
		), .Z(n_133094708));
	notech_ao4 i_190876783(.A(n_60197), .B(n_42689), .C(n_60010), .D(n_42463
		), .Z(n_133194709));
	notech_ao4 i_191276779(.A(n_60197), .B(n_42688), .C(n_60010), .D(n_42461
		), .Z(n_133294710));
	notech_ao4 i_191676775(.A(n_60197), .B(n_42687), .C(n_60010), .D(n_42459
		), .Z(n_133394711));
	notech_ao4 i_192076771(.A(n_60197), .B(n_42686), .C(n_60010), .D(n_42457
		), .Z(n_133494712));
	notech_ao4 i_192476767(.A(n_60182), .B(n_42685), .C(n_60010), .D(n_42455
		), .Z(n_133594713));
	notech_ao4 i_192876763(.A(n_60182), .B(n_42684), .C(n_60010), .D(n_42453
		), .Z(n_133694714));
	notech_ao4 i_193276759(.A(n_60182), .B(n_42683), .C(n_60010), .D(n_42451
		), .Z(n_133794715));
	notech_ao4 i_193676755(.A(n_60182), .B(n_42682), .C(n_60010), .D(n_42449
		), .Z(n_133894716));
	notech_ao4 i_194076751(.A(n_60182), .B(n_42681), .C(n_60007), .D(n_42447
		), .Z(n_133994717));
	notech_ao4 i_194476747(.A(n_60182), .B(n_42680), .C(n_60007), .D(n_42445
		), .Z(n_134094718));
	notech_ao4 i_194876743(.A(n_60182), .B(n_42679), .C(n_60008), .D(n_42443
		), .Z(n_134194719));
	notech_ao4 i_195276739(.A(n_60182), .B(n_42678), .C(n_60008), .D(n_42441
		), .Z(n_134294720));
	notech_ao4 i_195676735(.A(n_60202), .B(n_42677), .C(n_60007), .D(n_42439
		), .Z(n_134394721));
	notech_ao4 i_196076731(.A(n_60202), .B(n_42676), .C(n_60007), .D(n_42437
		), .Z(n_134494722));
	notech_ao4 i_196476727(.A(n_60202), .B(n_42675), .C(n_60007), .D(n_42435
		), .Z(n_134594723));
	notech_ao4 i_196876723(.A(n_60202), .B(n_42674), .C(n_60007), .D(n_42433
		), .Z(n_134694724));
	notech_ao4 i_197676715(.A(n_60202), .B(n_42672), .C(n_60008), .D(n_42429
		), .Z(n_134794725));
	notech_ao4 i_198076711(.A(n_60202), .B(n_42671), .C(n_60008), .D(n_42427
		), .Z(n_134894726));
	notech_ao4 i_198476707(.A(n_60202), .B(n_42670), .C(n_60008), .D(n_42425
		), .Z(n_134994727));
	notech_ao4 i_198876703(.A(n_60202), .B(n_42669), .C(n_60008), .D(n_42423
		), .Z(n_135094728));
	notech_ao4 i_199276699(.A(n_60216), .B(n_42668), .C(n_60008), .D(n_42421
		), .Z(n_135194729));
	notech_ao4 i_199676695(.A(n_60230), .B(n_42667), .C(n_60008), .D(n_42419
		), .Z(n_135294730));
	notech_ao4 i_200076691(.A(n_60230), .B(n_42666), .C(n_60008), .D(n_42417
		), .Z(n_135394731));
	notech_ao4 i_200476687(.A(n_60230), .B(n_42665), .C(n_60008), .D(n_42415
		), .Z(n_135494732));
	notech_ao4 i_200876683(.A(n_60230), .B(n_42664), .C(n_60008), .D(n_42413
		), .Z(n_135594733));
	notech_ao4 i_201276679(.A(n_60230), .B(n_42663), .C(n_60001), .D(n_42411
		), .Z(n_135694734));
	notech_ao4 i_201676675(.A(n_60230), .B(n_42662), .C(n_60001), .D(n_42409
		), .Z(n_135794735));
	notech_ao4 i_202476667(.A(n_60230), .B(n_42660), .C(n_59995), .D(n_42405
		), .Z(n_135894736));
	notech_ao4 i_202876663(.A(n_60230), .B(n_42659), .C(n_60001), .D(n_42403
		), .Z(n_135994737));
	notech_ao4 i_203276659(.A(n_60230), .B(n_42658), .C(n_60001), .D(n_42401
		), .Z(n_136094738));
	notech_ao4 i_203676655(.A(n_60230), .B(n_42657), .C(n_60003), .D(n_42399
		), .Z(n_136194739));
	notech_ao4 i_204076651(.A(n_60225), .B(n_42656), .C(n_60001), .D(n_42397
		), .Z(n_136294740));
	notech_ao4 i_204476647(.A(n_60225), .B(n_42655), .C(n_60001), .D(n_42395
		), .Z(n_136394741));
	notech_ao4 i_204876643(.A(n_60230), .B(n_42654), .C(n_59995), .D(n_42393
		), .Z(n_136494742));
	notech_ao4 i_205276639(.A(n_60230), .B(n_42653), .C(n_59995), .D(n_42391
		), .Z(n_136594743));
	notech_ao4 i_205676635(.A(n_60230), .B(n_42652), .C(n_59995), .D(n_42389
		), .Z(n_136694744));
	notech_ao4 i_206076631(.A(n_60230), .B(n_42651), .C(n_59995), .D(n_42387
		), .Z(n_136794745));
	notech_ao4 i_206476627(.A(n_141853051), .B(n_42650), .C(n_59995), .D(n_42385
		), .Z(n_136894746));
	notech_ao4 i_206876623(.A(n_141853051), .B(n_42649), .C(n_59995), .D(n_42383
		), .Z(n_136994747));
	notech_ao4 i_207276619(.A(n_141853051), .B(n_42648), .C(n_59995), .D(n_42381
		), .Z(n_137094748));
	notech_ao4 i_207676615(.A(n_141853051), .B(n_42647), .C(n_59995), .D(n_42379
		), .Z(n_137194749));
	notech_ao4 i_208076611(.A(n_141853051), .B(n_42646), .C(n_59995), .D(n_42377
		), .Z(n_137294750));
	notech_ao4 i_208476607(.A(n_141853051), .B(n_42645), .C(n_60008), .D(n_42375
		), .Z(n_137394751));
	notech_ao4 i_208876603(.A(n_141853051), .B(n_42644), .C(n_60008), .D(n_42373
		), .Z(n_137494752));
	notech_ao4 i_209276599(.A(n_141853051), .B(n_42643), .C(n_60010), .D(n_42371
		), .Z(n_137594753));
	notech_ao4 i_209676595(.A(n_141853051), .B(n_42642), .C(n_60010), .D(n_42369
		), .Z(n_137694754));
	notech_ao4 i_210076591(.A(n_141853051), .B(n_42641), .C(n_60008), .D(n_42367
		), .Z(n_137794755));
	notech_ao4 i_210476587(.A(n_60230), .B(n_42640), .C(n_60008), .D(n_42365
		), .Z(n_137894756));
	notech_ao4 i_210876583(.A(n_141853051), .B(n_42639), .C(n_60008), .D(n_42363
		), .Z(n_137994757));
	notech_ao4 i_211276579(.A(n_141853051), .B(n_42638), .C(n_60008), .D(n_42361
		), .Z(n_138094758));
	notech_ao4 i_211676575(.A(n_141853051), .B(n_42637), .C(n_60010), .D(n_42359
		), .Z(n_138194759));
	notech_ao4 i_212076571(.A(n_141853051), .B(n_42636), .C(n_60003), .D(n_42357
		), .Z(n_138294760));
	notech_ao4 i_212476567(.A(n_141853051), .B(n_42635), .C(n_60003), .D(n_42355
		), .Z(n_138394761));
	notech_ao4 i_212876563(.A(n_60221), .B(n_42634), .C(n_60003), .D(n_42353
		), .Z(n_138494762));
	notech_ao4 i_213276559(.A(n_60221), .B(n_42633), .C(n_60003), .D(n_42351
		), .Z(n_138594763));
	notech_ao4 i_213676555(.A(n_60221), .B(n_42632), .C(n_60010), .D(n_42349
		), .Z(n_138694764));
	notech_ao4 i_214076551(.A(n_60221), .B(n_42631), .C(n_60010), .D(n_42347
		), .Z(n_138794765));
	notech_ao4 i_214476547(.A(n_60221), .B(n_42630), .C(n_60003), .D(n_42345
		), .Z(n_138894766));
	notech_ao4 i_215276539(.A(n_60221), .B(n_42628), .C(n_60010), .D(n_42341
		), .Z(n_138994767));
	notech_ao4 i_215676535(.A(n_60221), .B(n_42627), .C(n_59998), .D(n_42339
		), .Z(n_139094768));
	notech_ao4 i_216076531(.A(n_60221), .B(n_42626), .C(n_59998), .D(n_42337
		), .Z(n_139194769));
	notech_ao4 i_216476527(.A(n_60216), .B(n_42625), .C(n_59998), .D(n_42335
		), .Z(n_139294770));
	notech_ao4 i_216876523(.A(n_60216), .B(n_42624), .C(n_59998), .D(n_42333
		), .Z(n_139394771));
	notech_ao4 i_217376518(.A(n_59998), .B(n_42331), .C(n_60216), .D(n_42623
		), .Z(n_139494772));
	notech_ao4 i_217776514(.A(n_60216), .B(n_42622), .C(n_59996), .D(n_42329
		), .Z(n_139594773));
	notech_ao4 i_218576506(.A(n_60221), .B(n_42620), .C(n_59998), .D(n_42325
		), .Z(n_139694774));
	notech_ao4 i_218976502(.A(n_60221), .B(n_42619), .C(n_59998), .D(n_42323
		), .Z(n_139794775));
	notech_ao4 i_219376498(.A(n_60221), .B(n_42618), .C(n_59998), .D(n_42321
		), .Z(n_139894776));
	notech_ao4 i_219776494(.A(n_60221), .B(n_42617), .C(n_59998), .D(n_42319
		), .Z(n_139994777));
	notech_ao4 i_220176490(.A(n_60225), .B(n_42616), .C(n_59998), .D(n_42317
		), .Z(n_140094778));
	notech_ao4 i_220576486(.A(n_60225), .B(n_42615), .C(n_60001), .D(n_42315
		), .Z(n_140194779));
	notech_ao4 i_220976482(.A(n_60225), .B(n_42614), .C(n_60001), .D(n_42313
		), .Z(n_140294780));
	notech_ao4 i_221776474(.A(n_60225), .B(n_42612), .C(n_59998), .D(n_42309
		), .Z(n_140394781));
	notech_ao4 i_222176470(.A(n_60225), .B(n_42611), .C(n_59998), .D(n_42307
		), .Z(n_140494782));
	notech_ao4 i_222576466(.A(n_60225), .B(n_42610), .C(n_59998), .D(n_42305
		), .Z(n_140594783));
	notech_ao4 i_222976462(.A(n_60225), .B(n_42609), .C(n_59998), .D(n_42303
		), .Z(n_140694784));
	notech_ao4 i_223376458(.A(n_60225), .B(n_42608), .C(n_59996), .D(n_42301
		), .Z(n_140794785));
	notech_ao4 i_223776454(.A(n_60221), .B(n_42607), .C(n_59996), .D(n_42299
		), .Z(n_140894786));
	notech_ao4 i_224176450(.A(n_60225), .B(n_42606), .C(n_59996), .D(n_42297
		), .Z(n_140994787));
	notech_ao4 i_224976442(.A(n_60221), .B(n_42604), .C(n_59996), .D(n_42293
		), .Z(n_141094788));
	notech_ao4 i_225376438(.A(n_60221), .B(n_42603), .C(n_59995), .D(n_42291
		), .Z(n_141194789));
	notech_nand3 i_3593499(.A(n_58216), .B(queue[7]), .C(n_57947), .Z(n_141294790
		));
	notech_or2 i_3693514(.A(n_58225), .B(n_42192), .Z(n_142794805));
	notech_nand3 i_824987(.A(n_230495682), .B(n_229795675), .C(n_141294790),
		 .Z(squeue[7]));
	notech_nand3 i_19293515(.A(n_57947), .B(n_58216), .C(queue[55]), .Z(n_142894806
		));
	notech_or2 i_19393530(.A(n_58225), .B(n_42240), .Z(n_144394821));
	notech_nand3 i_5625035(.A(n_231895696), .B(n_231195689), .C(n_142894806)
		, .Z(squeue[55]));
	notech_nand3 i_22393531(.A(n_57947), .B(n_58216), .C(queue[56]), .Z(n_144494822
		));
	notech_or2 i_22493546(.A(n_58225), .B(n_42241), .Z(n_145994837));
	notech_nand3 i_5725036(.A(n_233295710), .B(n_232595703), .C(n_144494822)
		, .Z(squeue[56]));
	notech_nand3 i_25493547(.A(n_57945), .B(n_58216), .C(queue[57]), .Z(n_146094838
		));
	notech_or2 i_25593562(.A(n_58225), .B(n_42242), .Z(n_147594853));
	notech_nand3 i_5825037(.A(n_234695724), .B(n_233995717), .C(n_146094838)
		, .Z(squeue[57]));
	notech_nand3 i_28593563(.A(n_57945), .B(n_58216), .C(queue[58]), .Z(n_147694854
		));
	notech_or2 i_28693578(.A(n_58225), .B(n_42243), .Z(n_149194869));
	notech_nand3 i_5925038(.A(n_236095738), .B(n_235395731), .C(n_147694854)
		, .Z(squeue[58]));
	notech_nand3 i_31693579(.A(n_57945), .B(n_58216), .C(queue[59]), .Z(n_149294870
		));
	notech_or2 i_31793594(.A(n_58225), .B(n_42244), .Z(n_150794885));
	notech_nand3 i_6025039(.A(n_237495752), .B(n_236795745), .C(n_149294870)
		, .Z(squeue[59]));
	notech_nand3 i_34793595(.A(n_57945), .B(n_58216), .C(queue[60]), .Z(n_150894886
		));
	notech_or2 i_34893610(.A(n_58225), .B(n_42245), .Z(n_152394901));
	notech_nand3 i_6125040(.A(n_238895766), .B(n_238195759), .C(n_150894886)
		, .Z(squeue[60]));
	notech_nand3 i_44093611(.A(n_57945), .B(n_58216), .C(queue[63]), .Z(n_152494902
		));
	notech_or2 i_44193626(.A(n_58225), .B(n_42248), .Z(n_153994917));
	notech_nand3 i_6425043(.A(n_240295780), .B(n_239595773), .C(n_152494902)
		, .Z(squeue[63]));
	notech_nand3 i_50293627(.A(n_57945), .B(n_58216), .C(queue[66]), .Z(n_154094918
		));
	notech_or2 i_50393642(.A(n_58222), .B(n_42251), .Z(n_155594933));
	notech_nand3 i_6725046(.A(n_241695794), .B(n_240995787), .C(n_154094918)
		, .Z(squeue[66]));
	notech_nand3 i_53393643(.A(n_57945), .B(n_58216), .C(queue[67]), .Z(n_155694934
		));
	notech_or2 i_53493658(.A(n_58222), .B(n_42252), .Z(n_157194949));
	notech_nand3 i_6825047(.A(n_243095808), .B(n_242395801), .C(n_155694934)
		, .Z(squeue[67]));
	notech_nand3 i_56493659(.A(n_57945), .B(n_58218), .C(queue[68]), .Z(n_157294950
		));
	notech_or2 i_56593674(.A(n_58222), .B(n_42253), .Z(n_158794965));
	notech_nand3 i_6925048(.A(n_244495822), .B(n_243795815), .C(n_157294950)
		, .Z(squeue[68]));
	notech_nand3 i_65793675(.A(n_57945), .B(n_58216), .C(queue[71]), .Z(n_158894966
		));
	notech_or2 i_65893690(.A(n_58222), .B(n_42256), .Z(n_160394981));
	notech_nand3 i_7225051(.A(n_245895836), .B(n_245195829), .C(n_158894966)
		, .Z(squeue[71]));
	notech_nand3 i_68893691(.A(n_57945), .B(n_58216), .C(queue[72]), .Z(n_160494982
		));
	notech_or2 i_68993706(.A(n_58222), .B(n_42257), .Z(n_161994997));
	notech_nand3 i_7325052(.A(n_247295850), .B(n_246595843), .C(n_160494982)
		, .Z(squeue[72]));
	notech_nand3 i_71993707(.A(n_57945), .B(n_58216), .C(queue[73]), .Z(n_162094998
		));
	notech_or2 i_72093722(.A(n_58222), .B(n_42258), .Z(n_163595013));
	notech_nand3 i_7425053(.A(n_248695864), .B(n_247995857), .C(n_162094998)
		, .Z(squeue[73]));
	notech_nand3 i_75093723(.A(n_57945), .B(n_58216), .C(queue[74]), .Z(n_163695014
		));
	notech_or2 i_75193738(.A(n_58222), .B(n_42259), .Z(n_165195029));
	notech_nand3 i_7525054(.A(n_250095878), .B(n_249395871), .C(n_163695014)
		, .Z(squeue[74]));
	notech_nand3 i_78193739(.A(n_57945), .B(n_58216), .C(queue[75]), .Z(n_165295030
		));
	notech_or2 i_78293754(.A(n_58222), .B(n_42260), .Z(n_166795045));
	notech_nand3 i_7625055(.A(n_251495892), .B(n_250795885), .C(n_165295030)
		, .Z(squeue[75]));
	notech_nand3 i_81293755(.A(n_57945), .B(n_58204), .C(queue[76]), .Z(n_166895046
		));
	notech_or2 i_81393770(.A(n_58223), .B(n_42261), .Z(n_168395061));
	notech_nand3 i_7725056(.A(n_252895906), .B(n_252195899), .C(n_166895046)
		, .Z(squeue[76]));
	notech_nand3 i_90593771(.A(n_57945), .B(n_58204), .C(queue[79]), .Z(n_168495062
		));
	notech_or2 i_90693786(.A(n_58223), .B(n_42264), .Z(n_169995077));
	notech_nand3 i_8025059(.A(n_254295920), .B(n_253595913), .C(n_168495062)
		, .Z(squeue[79]));
	notech_nand3 i_93693787(.A(n_57945), .B(n_58204), .C(queue[80]), .Z(n_170095078
		));
	notech_or2 i_93793802(.A(n_58223), .B(n_42265), .Z(n_171595093));
	notech_nand3 i_8125060(.A(n_255695934), .B(n_254995927), .C(n_170095078)
		, .Z(squeue[80]));
	notech_nand3 i_96793803(.A(n_57932), .B(n_58204), .C(queue[81]), .Z(n_171695094
		));
	notech_or2 i_96893818(.A(n_58223), .B(n_42266), .Z(n_173195109));
	notech_nand3 i_8225061(.A(n_257095948), .B(n_256395941), .C(n_171695094)
		, .Z(squeue[81]));
	notech_nand3 i_99893819(.A(n_57932), .B(n_58204), .C(queue[82]), .Z(n_173295110
		));
	notech_or2 i_99993834(.A(n_58223), .B(n_42267), .Z(n_174795125));
	notech_nand3 i_8325062(.A(n_258495962), .B(n_257795955), .C(n_173295110)
		, .Z(squeue[82]));
	notech_nand3 i_102993835(.A(n_57932), .B(n_58204), .C(queue[83]), .Z(n_174895126
		));
	notech_or2 i_103093850(.A(n_58223), .B(n_42268), .Z(n_176395141));
	notech_nand3 i_8425063(.A(n_259895976), .B(n_259195969), .C(n_174895126)
		, .Z(squeue[83]));
	notech_nand3 i_106093851(.A(n_57932), .B(n_58204), .C(queue[84]), .Z(n_176495142
		));
	notech_or2 i_106193866(.A(n_58223), .B(n_42269), .Z(n_177995157));
	notech_nand3 i_8525064(.A(n_261295990), .B(n_260595983), .C(n_176495142)
		, .Z(squeue[84]));
	notech_nand3 i_115393867(.A(n_57932), .B(n_58204), .C(queue[87]), .Z(n_178095158
		));
	notech_or2 i_115493882(.A(n_58223), .B(n_42272), .Z(n_179595173));
	notech_nand3 i_8825067(.A(n_262696004), .B(n_261995997), .C(n_178095158)
		, .Z(squeue[87]));
	notech_nand3 i_118493883(.A(n_57932), .B(n_58206), .C(queue[88]), .Z(n_179695174
		));
	notech_or2 i_118593898(.A(n_58228), .B(n_42273), .Z(n_181195189));
	notech_nand3 i_8925068(.A(n_264096018), .B(n_263396011), .C(n_179695174)
		, .Z(squeue[88]));
	notech_nand3 i_121593899(.A(n_57932), .B(n_58206), .C(queue[89]), .Z(n_181295190
		));
	notech_or2 i_121693914(.A(n_58228), .B(n_42274), .Z(n_182795205));
	notech_nand3 i_9025069(.A(n_265496032), .B(n_264796025), .C(n_181295190)
		, .Z(squeue[89]));
	notech_nand3 i_124693915(.A(n_57932), .B(n_58206), .C(queue[90]), .Z(n_182895206
		));
	notech_or2 i_124793930(.A(n_58228), .B(n_42275), .Z(n_184395221));
	notech_nand3 i_9125070(.A(n_266896046), .B(n_266196039), .C(n_182895206)
		, .Z(squeue[90]));
	notech_nand3 i_127793931(.A(n_57932), .B(n_58206), .C(queue[91]), .Z(n_184495222
		));
	notech_or2 i_127893946(.A(n_58228), .B(n_42276), .Z(n_185995237));
	notech_nand3 i_9225071(.A(n_268296060), .B(n_267596053), .C(n_184495222)
		, .Z(squeue[91]));
	notech_nand3 i_130893947(.A(n_57932), .B(n_58206), .C(queue[92]), .Z(n_186095238
		));
	notech_or2 i_130993962(.A(n_58228), .B(n_42277), .Z(n_187595253));
	notech_nand3 i_9325072(.A(n_269696074), .B(n_268996067), .C(n_186095238)
		, .Z(squeue[92]));
	notech_nand3 i_140193963(.A(n_57932), .B(n_58204), .C(queue[95]), .Z(n_187695254
		));
	notech_or2 i_140293978(.A(n_58228), .B(n_42280), .Z(n_189195269));
	notech_nand3 i_9625075(.A(n_271096088), .B(n_270396081), .C(n_187695254)
		, .Z(squeue[95]));
	notech_nand3 i_143293979(.A(n_57932), .B(n_58206), .C(queue[96]), .Z(n_189295270
		));
	notech_or2 i_143393994(.A(n_58228), .B(n_42281), .Z(n_190795285));
	notech_nand3 i_9725076(.A(n_272496102), .B(n_271796095), .C(n_189295270)
		, .Z(squeue[96]));
	notech_nand3 i_146393995(.A(n_57932), .B(n_58206), .C(queue[97]), .Z(n_190895286
		));
	notech_or2 i_146494010(.A(n_58228), .B(n_42282), .Z(n_192395301));
	notech_nand3 i_9825077(.A(n_273896116), .B(n_273196109), .C(n_190895286)
		, .Z(squeue[97]));
	notech_nand3 i_149494011(.A(n_57932), .B(n_58204), .C(queue[98]), .Z(n_192495302
		));
	notech_or2 i_149594026(.A(n_58230), .B(n_42283), .Z(n_193995317));
	notech_nand3 i_9925078(.A(n_275296130), .B(n_274596123), .C(n_192495302)
		, .Z(squeue[98]));
	notech_nand3 i_152594027(.A(n_57932), .B(n_58203), .C(queue[99]), .Z(n_194095318
		));
	notech_or2 i_152694042(.A(n_58230), .B(n_42284), .Z(n_195595333));
	notech_nand3 i_10025079(.A(n_276696144), .B(n_275996137), .C(n_194095318
		), .Z(squeue[99]));
	notech_nand3 i_155694043(.A(n_57932), .B(n_58203), .C(queue[100]), .Z(n_195695334
		));
	notech_or2 i_155794058(.A(n_58230), .B(n_42285), .Z(n_197195349));
	notech_nand3 i_10125080(.A(n_278096158), .B(n_277396151), .C(n_195695334
		), .Z(squeue[100]));
	notech_nand3 i_1649(.A(n_57930), .B(n_58203), .C(queue[103]), .Z(n_197295350
		));
	notech_or2 i_1650(.A(n_58230), .B(n_42288), .Z(n_198795365));
	notech_nand3 i_10425083(.A(n_279496172), .B(n_278796165), .C(n_197295350
		), .Z(squeue[103]));
	notech_nand3 i_1680(.A(n_57930), .B(n_58203), .C(queue[104]), .Z(n_198895366
		));
	notech_or2 i_1681(.A(n_58230), .B(n_42291), .Z(n_200395381));
	notech_nand3 i_10525084(.A(n_280896186), .B(n_280196179), .C(n_198895366
		), .Z(squeue[104]));
	notech_nand3 i_1711(.A(n_57930), .B(n_58203), .C(queue[105]), .Z(n_200495382
		));
	notech_or2 i_1712(.A(n_58228), .B(n_42293), .Z(n_201995397));
	notech_nand3 i_10625085(.A(n_282296200), .B(n_281596193), .C(n_200495382
		), .Z(squeue[105]));
	notech_nand3 i_1742(.A(n_57930), .B(n_58203), .C(queue[106]), .Z(n_202095398
		));
	notech_or2 i_1743(.A(n_58230), .B(n_42295), .Z(n_203595413));
	notech_nand3 i_10725086(.A(n_283696214), .B(n_282996207), .C(n_202095398
		), .Z(squeue[106]));
	notech_nand3 i_1773(.A(n_57930), .B(n_58203), .C(queue[107]), .Z(n_203695414
		));
	notech_or2 i_1774(.A(n_58230), .B(n_42297), .Z(n_205195429));
	notech_nand3 i_10825087(.A(n_285096228), .B(n_284396221), .C(n_203695414
		), .Z(squeue[107]));
	notech_nand3 i_1804(.A(n_57930), .B(n_58203), .C(queue[108]), .Z(n_205295430
		));
	notech_or2 i_1805(.A(n_58225), .B(n_42299), .Z(n_206795445));
	notech_nand3 i_10925088(.A(n_286496242), .B(n_285796235), .C(n_205295430
		), .Z(squeue[108]));
	notech_nand3 i_1897(.A(n_57930), .B(n_58204), .C(queue[111]), .Z(n_206895446
		));
	notech_or2 i_1898(.A(n_58225), .B(n_42305), .Z(n_208395461));
	notech_nand3 i_11225091(.A(n_287896256), .B(n_287196249), .C(n_206895446
		), .Z(squeue[111]));
	notech_nand3 i_1928(.A(n_57930), .B(n_58204), .C(queue[112]), .Z(n_208495462
		));
	notech_or2 i_1929(.A(n_58225), .B(n_42307), .Z(n_209995477));
	notech_nand3 i_11325092(.A(n_289296270), .B(n_288596263), .C(n_208495462
		), .Z(squeue[112]));
	notech_nand3 i_1959(.A(n_57930), .B(n_58204), .C(queue[113]), .Z(n_210095478
		));
	notech_or2 i_1960(.A(n_58225), .B(n_42309), .Z(n_211595493));
	notech_nand3 i_11425093(.A(n_290696284), .B(n_289996277), .C(n_210095478
		), .Z(squeue[113]));
	notech_nand3 i_1990(.A(n_57930), .B(n_58204), .C(queue[114]), .Z(n_211695494
		));
	notech_or2 i_1991(.A(n_58225), .B(n_42311), .Z(n_213195509));
	notech_nand3 i_11525094(.A(n_292096298), .B(n_291396291), .C(n_211695494
		), .Z(squeue[114]));
	notech_nand3 i_2021(.A(n_57930), .B(n_58204), .C(queue[115]), .Z(n_213295510
		));
	notech_or2 i_2022(.A(n_58225), .B(n_42313), .Z(n_214795525));
	notech_nand3 i_11625095(.A(n_293596312), .B(n_292796305), .C(n_213295510
		), .Z(squeue[115]));
	notech_nand3 i_2052(.A(n_57930), .B(n_58204), .C(queue[116]), .Z(n_214895526
		));
	notech_or2 i_2053(.A(n_58225), .B(n_42315), .Z(n_216395541));
	notech_nand3 i_11725096(.A(n_295496326), .B(n_294496319), .C(n_214895526
		), .Z(squeue[116]));
	notech_nand3 i_2145(.A(n_57930), .B(n_58204), .C(queue[119]), .Z(n_216495542
		));
	notech_or2 i_2146(.A(n_58225), .B(n_42321), .Z(n_217995557));
	notech_nand3 i_12025099(.A(n_296996340), .B(n_296196333), .C(n_216495542
		), .Z(squeue[119]));
	notech_nand3 i_2176(.A(n_57930), .B(n_58204), .C(queue[120]), .Z(n_218095558
		));
	notech_or2 i_2177(.A(n_58228), .B(n_42323), .Z(n_219595573));
	notech_nand3 i_12125100(.A(n_298396354), .B(n_297696347), .C(n_218095558
		), .Z(squeue[120]));
	notech_nand3 i_2207(.A(n_57930), .B(n_58206), .C(queue[121]), .Z(n_219695574
		));
	notech_or2 i_2208(.A(n_58228), .B(n_42325), .Z(n_221195589));
	notech_nand3 i_12225101(.A(n_299796368), .B(n_299096361), .C(n_219695574
		), .Z(squeue[121]));
	notech_nand3 i_2238(.A(n_57930), .B(n_58209), .C(queue[122]), .Z(n_221295590
		));
	notech_or2 i_2239(.A(n_58228), .B(n_42327), .Z(n_222795605));
	notech_nand3 i_12325102(.A(n_301196382), .B(n_300496375), .C(n_221295590
		), .Z(squeue[122]));
	notech_nand3 i_2269(.A(n_57937), .B(n_58209), .C(queue[123]), .Z(n_222895606
		));
	notech_or2 i_2270(.A(n_58228), .B(n_42329), .Z(n_224395621));
	notech_nand3 i_12425103(.A(n_302596396), .B(n_301896389), .C(n_222895606
		), .Z(squeue[123]));
	notech_nand3 i_2300(.A(n_57937), .B(n_58209), .C(queue[124]), .Z(n_224495622
		));
	notech_or2 i_2301(.A(n_58228), .B(n_42331), .Z(n_225995637));
	notech_nand3 i_12525104(.A(n_303996410), .B(n_303296403), .C(n_224495622
		), .Z(squeue[124]));
	notech_nand3 i_2331(.A(n_57937), .B(n_58209), .C(queue[125]), .Z(n_226095638
		));
	notech_or2 i_2332(.A(n_58228), .B(n_42333), .Z(n_227595653));
	notech_nand3 i_12625105(.A(n_305396424), .B(n_304696417), .C(n_226095638
		), .Z(squeue[125]));
	notech_nand3 i_2393(.A(n_57937), .B(n_58209), .C(queue[127]), .Z(n_227695654
		));
	notech_or2 i_2394(.A(n_58228), .B(n_42337), .Z(n_229195669));
	notech_nand3 i_12825107(.A(n_306796438), .B(n_306096431), .C(n_227695654
		), .Z(squeue[127]));
	notech_ao4 i_3794059(.A(n_58307), .B(n_42200), .C(n_58291), .D(n_42216),
		 .Z(n_229295670));
	notech_ao4 i_3894061(.A(n_58244), .B(n_42184), .C(n_42288), .D(n_57963),
		 .Z(n_229495672));
	notech_ao4 i_3994062(.A(n_42272), .B(n_57995), .C(n_42280), .D(n_57979),
		 .Z(n_229595673));
	notech_and4 i_4894064(.A(n_229595673), .B(n_229495672), .C(n_229295670),
		 .D(n_142794805), .Z(n_229795675));
	notech_ao4 i_4094065(.A(n_42256), .B(n_58027), .C(n_42264), .D(n_58011),
		 .Z(n_229895676));
	notech_ao4 i_4194066(.A(n_42240), .B(n_58323), .C(n_42248), .D(n_58043),
		 .Z(n_229995677));
	notech_ao4 i_4294068(.A(n_42224), .B(n_58355), .C(n_58339), .D(n_42232),
		 .Z(n_230195679));
	notech_ao4 i_4394069(.A(n_58274), .B(n_42176), .C(n_58371), .D(n_42208),
		 .Z(n_230295680));
	notech_and4 i_4994071(.A(n_230295680), .B(n_230195679), .C(n_229995677),
		 .D(n_229895676), .Z(n_230495682));
	notech_ao4 i_19494073(.A(n_58307), .B(n_42248), .C(n_58291), .D(n_42264)
		, .Z(n_230695684));
	notech_ao4 i_19594075(.A(n_58244), .B(n_42232), .C(n_57963), .D(n_42385)
		, .Z(n_230895686));
	notech_ao4 i_19694076(.A(n_57995), .B(n_42353), .C(n_57979), .D(n_42369)
		, .Z(n_230995687));
	notech_and4 i_20594078(.A(n_230995687), .B(n_230895686), .C(n_230695684)
		, .D(n_144394821), .Z(n_231195689));
	notech_ao4 i_19794079(.A(n_58027), .B(n_42321), .C(n_58011), .D(n_42337)
		, .Z(n_231295690));
	notech_ao4 i_19894080(.A(n_58323), .B(n_42288), .C(n_58043), .D(n_42305)
		, .Z(n_231395691));
	notech_ao4 i_19994082(.A(n_58355), .B(n_42272), .C(n_58339), .D(n_42280)
		, .Z(n_231595693));
	notech_ao4 i_20094083(.A(n_58274), .B(n_42224), .C(n_58371), .D(n_42256)
		, .Z(n_231695694));
	notech_and4 i_20694085(.A(n_231695694), .B(n_231595693), .C(n_231395691)
		, .D(n_231295690), .Z(n_231895696));
	notech_ao4 i_22594087(.A(n_58307), .B(n_42249), .C(n_58291), .D(n_42265)
		, .Z(n_232095698));
	notech_ao4 i_22694089(.A(n_58244), .B(n_42233), .C(n_57963), .D(n_42387)
		, .Z(n_232295700));
	notech_ao4 i_22794090(.A(n_57995), .B(n_42355), .C(n_57979), .D(n_42371)
		, .Z(n_232395701));
	notech_and4 i_23694092(.A(n_232395701), .B(n_232295700), .C(n_232095698)
		, .D(n_145994837), .Z(n_232595703));
	notech_ao4 i_22894093(.A(n_58027), .B(n_42323), .C(n_58011), .D(n_42339)
		, .Z(n_232695704));
	notech_ao4 i_22994094(.A(n_58323), .B(n_42291), .C(n_58043), .D(n_42307)
		, .Z(n_232795705));
	notech_ao4 i_23094096(.A(n_58355), .B(n_42273), .C(n_58339), .D(n_42281)
		, .Z(n_232995707));
	notech_ao4 i_23194097(.A(n_58274), .B(n_42225), .C(n_58371), .D(n_42257)
		, .Z(n_233095708));
	notech_and4 i_23794099(.A(n_233095708), .B(n_232995707), .C(n_232795705)
		, .D(n_232695704), .Z(n_233295710));
	notech_ao4 i_25694101(.A(n_58307), .B(n_42250), .C(n_58291), .D(n_42266)
		, .Z(n_233495712));
	notech_ao4 i_25779461(.A(n_58244), .B(n_42234), .C(n_57963), .D(n_42389)
		, .Z(n_233695714));
	notech_ao4 i_25894103(.A(n_57995), .B(n_42357), .C(n_57979), .D(n_42373)
		, .Z(n_233795715));
	notech_and4 i_26794105(.A(n_233795715), .B(n_233695714), .C(n_233495712)
		, .D(n_147594853), .Z(n_233995717));
	notech_ao4 i_25994106(.A(n_58027), .B(n_42325), .C(n_58011), .D(n_42341)
		, .Z(n_234095718));
	notech_ao4 i_26094107(.A(n_58323), .B(n_42293), .C(n_58043), .D(n_42309)
		, .Z(n_234195719));
	notech_ao4 i_26194109(.A(n_58355), .B(n_42274), .C(n_58339), .D(n_42282)
		, .Z(n_234395721));
	notech_ao4 i_26294110(.A(n_58272), .B(n_42226), .C(n_58371), .D(n_42258)
		, .Z(n_234495722));
	notech_and4 i_26894112(.A(n_234495722), .B(n_234395721), .C(n_234195719)
		, .D(n_234095718), .Z(n_234695724));
	notech_ao4 i_28794114(.A(n_58307), .B(n_42251), .C(n_58291), .D(n_42267)
		, .Z(n_234895726));
	notech_ao4 i_28894116(.A(n_58244), .B(n_42235), .C(n_57963), .D(n_42391)
		, .Z(n_235095728));
	notech_ao4 i_28994117(.A(n_57995), .B(n_42359), .C(n_57979), .D(n_42375)
		, .Z(n_235195729));
	notech_and4 i_29894119(.A(n_235195729), .B(n_235095728), .C(n_234895726)
		, .D(n_149194869), .Z(n_235395731));
	notech_ao4 i_29094120(.A(n_58027), .B(n_42327), .C(n_58011), .D(n_42343)
		, .Z(n_235495732));
	notech_ao4 i_29194121(.A(n_58323), .B(n_42295), .C(n_58043), .D(n_42311)
		, .Z(n_235595733));
	notech_ao4 i_29294123(.A(n_58355), .B(n_42275), .C(n_58339), .D(n_42283)
		, .Z(n_235795735));
	notech_ao4 i_29394124(.A(n_58274), .B(n_42227), .C(n_58371), .D(n_42259)
		, .Z(n_235895736));
	notech_and4 i_29994126(.A(n_235895736), .B(n_235795735), .C(n_235595733)
		, .D(n_235495732), .Z(n_236095738));
	notech_ao4 i_31894128(.A(n_58307), .B(n_42252), .C(n_58291), .D(n_42268)
		, .Z(n_236295740));
	notech_ao4 i_31994130(.A(n_58244), .B(n_42236), .C(n_57963), .D(n_42393)
		, .Z(n_236495742));
	notech_ao4 i_32094131(.A(n_57995), .B(n_42361), .C(n_57979), .D(n_42377)
		, .Z(n_236595743));
	notech_and4 i_32994133(.A(n_236595743), .B(n_236495742), .C(n_236295740)
		, .D(n_150794885), .Z(n_236795745));
	notech_ao4 i_32194134(.A(n_58027), .B(n_42329), .C(n_58011), .D(n_42345)
		, .Z(n_236895746));
	notech_ao4 i_32294135(.A(n_58323), .B(n_42297), .C(n_58043), .D(n_42313)
		, .Z(n_236995747));
	notech_ao4 i_32394137(.A(n_58355), .B(n_42276), .C(n_58339), .D(n_42284)
		, .Z(n_237195749));
	notech_ao4 i_32494138(.A(n_58272), .B(n_42228), .C(n_58371), .D(n_42260)
		, .Z(n_237295750));
	notech_and4 i_33094140(.A(n_237295750), .B(n_237195749), .C(n_236995747)
		, .D(n_236895746), .Z(n_237495752));
	notech_ao4 i_34994142(.A(n_58307), .B(n_42253), .C(n_58291), .D(n_42269)
		, .Z(n_237695754));
	notech_ao4 i_35094144(.A(n_58244), .B(n_42237), .C(n_57963), .D(n_42395)
		, .Z(n_237895756));
	notech_ao4 i_35194145(.A(n_57995), .B(n_42363), .C(n_57979), .D(n_42379)
		, .Z(n_237995757));
	notech_and4 i_36094147(.A(n_237995757), .B(n_237895756), .C(n_237695754)
		, .D(n_152394901), .Z(n_238195759));
	notech_ao4 i_35294148(.A(n_58027), .B(n_42331), .C(n_58011), .D(n_42347)
		, .Z(n_238295760));
	notech_ao4 i_35394149(.A(n_58323), .B(n_42299), .C(n_58043), .D(n_42315)
		, .Z(n_238395761));
	notech_ao4 i_35494151(.A(n_58355), .B(n_42277), .C(n_58339), .D(n_42285)
		, .Z(n_238595763));
	notech_ao4 i_35594152(.A(n_58272), .B(n_42229), .C(n_58371), .D(n_42261)
		, .Z(n_238695764));
	notech_and4 i_36194154(.A(n_238695764), .B(n_238595763), .C(n_238395761)
		, .D(n_238295760), .Z(n_238895766));
	notech_ao4 i_44294156(.A(n_58305), .B(n_42256), .C(n_58289), .D(n_42272)
		, .Z(n_239095768));
	notech_ao4 i_44394158(.A(n_58244), .B(n_42240), .C(n_57961), .D(n_42401)
		, .Z(n_239295770));
	notech_ao4 i_44494159(.A(n_57993), .B(n_42369), .C(n_57977), .D(n_42385)
		, .Z(n_239395771));
	notech_and4 i_45394161(.A(n_239395771), .B(n_239295770), .C(n_239095768)
		, .D(n_153994917), .Z(n_239595773));
	notech_ao4 i_44594162(.A(n_58025), .B(n_42337), .C(n_58009), .D(n_42353)
		, .Z(n_239695774));
	notech_ao4 i_44694163(.A(n_58321), .B(n_42305), .C(n_58041), .D(n_42321)
		, .Z(n_239795775));
	notech_ao4 i_44794165(.A(n_58353), .B(n_42280), .C(n_58337), .D(n_42288)
		, .Z(n_239995777));
	notech_ao4 i_44894166(.A(n_58272), .B(n_42232), .C(n_58369), .D(n_42264)
		, .Z(n_240095778));
	notech_and4 i_45494168(.A(n_240095778), .B(n_239995777), .C(n_239795775)
		, .D(n_239695774), .Z(n_240295780));
	notech_ao4 i_50494170(.A(n_58305), .B(n_42259), .C(n_58289), .D(n_42275)
		, .Z(n_240495782));
	notech_ao4 i_50594172(.A(n_58241), .B(n_42243), .C(n_57961), .D(n_42407)
		, .Z(n_240695784));
	notech_ao4 i_50694173(.A(n_57993), .B(n_42375), .C(n_57977), .D(n_42391)
		, .Z(n_240795785));
	notech_and4 i_51594175(.A(n_240795785), .B(n_240695784), .C(n_240495782)
		, .D(n_155594933), .Z(n_240995787));
	notech_ao4 i_50794176(.A(n_58025), .B(n_42343), .C(n_58009), .D(n_42359)
		, .Z(n_241095788));
	notech_ao4 i_50894177(.A(n_58321), .B(n_42311), .C(n_58041), .D(n_42327)
		, .Z(n_241195789));
	notech_ao4 i_50994179(.A(n_58353), .B(n_42283), .C(n_58337), .D(n_42295)
		, .Z(n_241395791));
	notech_ao4 i_51094180(.A(n_58274), .B(n_42235), .C(n_58369), .D(n_42267)
		, .Z(n_241495792));
	notech_and4 i_51694182(.A(n_241495792), .B(n_241395791), .C(n_241195789)
		, .D(n_241095788), .Z(n_241695794));
	notech_ao4 i_53594184(.A(n_58305), .B(n_42260), .C(n_58289), .D(n_42276)
		, .Z(n_241895796));
	notech_ao4 i_53694186(.A(n_58241), .B(n_42244), .C(n_57961), .D(n_42409)
		, .Z(n_242095798));
	notech_ao4 i_53794187(.A(n_57993), .B(n_42377), .C(n_57977), .D(n_42393)
		, .Z(n_242195799));
	notech_and4 i_54694189(.A(n_242195799), .B(n_242095798), .C(n_241895796)
		, .D(n_157194949), .Z(n_242395801));
	notech_ao4 i_53894190(.A(n_58025), .B(n_42345), .C(n_58009), .D(n_42361)
		, .Z(n_242495802));
	notech_ao4 i_53994191(.A(n_58321), .B(n_42313), .C(n_58041), .D(n_42329)
		, .Z(n_242595803));
	notech_ao4 i_54094193(.A(n_58353), .B(n_42284), .C(n_58337), .D(n_42297)
		, .Z(n_242795805));
	notech_ao4 i_54194194(.A(n_58274), .B(n_42236), .C(n_58369), .D(n_42268)
		, .Z(n_242895806));
	notech_and4 i_54794196(.A(n_242895806), .B(n_242795805), .C(n_242595803)
		, .D(n_242495802), .Z(n_243095808));
	notech_ao4 i_56694198(.A(n_58305), .B(n_42261), .C(n_58289), .D(n_42277)
		, .Z(n_243295810));
	notech_ao4 i_56794200(.A(n_58241), .B(n_42245), .C(n_57961), .D(n_42411)
		, .Z(n_243495812));
	notech_ao4 i_56894201(.A(n_57993), .B(n_42379), .C(n_57977), .D(n_42395)
		, .Z(n_243595813));
	notech_and4 i_57794203(.A(n_243595813), .B(n_243495812), .C(n_243295810)
		, .D(n_158794965), .Z(n_243795815));
	notech_ao4 i_56994204(.A(n_58025), .B(n_42347), .C(n_58009), .D(n_42363)
		, .Z(n_243895816));
	notech_ao4 i_57094205(.A(n_58321), .B(n_42315), .C(n_58041), .D(n_42331)
		, .Z(n_243995817));
	notech_ao4 i_57194207(.A(n_58353), .B(n_42285), .C(n_58337), .D(n_42299)
		, .Z(n_244195819));
	notech_ao4 i_57294208(.A(n_58274), .B(n_42237), .C(n_58369), .D(n_42269)
		, .Z(n_244295820));
	notech_and4 i_57894210(.A(n_244295820), .B(n_244195819), .C(n_243995817)
		, .D(n_243895816), .Z(n_244495822));
	notech_ao4 i_65994212(.A(n_58305), .B(n_42264), .C(n_58289), .D(n_42280)
		, .Z(n_244695824));
	notech_ao4 i_66094214(.A(n_58241), .B(n_42248), .C(n_57961), .D(n_42417)
		, .Z(n_244895826));
	notech_ao4 i_66194215(.A(n_57993), .B(n_42385), .C(n_57977), .D(n_42401)
		, .Z(n_244995827));
	notech_and4 i_67094217(.A(n_244995827), .B(n_244895826), .C(n_244695824)
		, .D(n_160394981), .Z(n_245195829));
	notech_ao4 i_66294218(.A(n_58025), .B(n_42353), .C(n_58009), .D(n_42369)
		, .Z(n_245295830));
	notech_ao4 i_66394219(.A(n_58321), .B(n_42321), .C(n_58041), .D(n_42337)
		, .Z(n_245395831));
	notech_ao4 i_66494221(.A(n_58353), .B(n_42288), .C(n_58337), .D(n_42305)
		, .Z(n_245595833));
	notech_ao4 i_66594222(.A(n_58274), .B(n_42240), .C(n_58369), .D(n_42272)
		, .Z(n_245695834));
	notech_and4 i_67194224(.A(n_245695834), .B(n_245595833), .C(n_245395831)
		, .D(n_245295830), .Z(n_245895836));
	notech_ao4 i_69094226(.A(n_58307), .B(n_42265), .C(n_58291), .D(n_42281)
		, .Z(n_246095838));
	notech_ao4 i_69194228(.A(n_58241), .B(n_42249), .C(n_57963), .D(n_42419)
		, .Z(n_246295840));
	notech_ao4 i_69294229(.A(n_57995), .B(n_42387), .C(n_57979), .D(n_42403)
		, .Z(n_246395841));
	notech_and4 i_70194231(.A(n_246395841), .B(n_246295840), .C(n_246095838)
		, .D(n_161994997), .Z(n_246595843));
	notech_ao4 i_69394232(.A(n_58027), .B(n_42355), .C(n_58011), .D(n_42371)
		, .Z(n_246695844));
	notech_ao4 i_69494233(.A(n_58323), .B(n_42323), .C(n_58043), .D(n_42339)
		, .Z(n_246795845));
	notech_ao4 i_69594235(.A(n_58355), .B(n_42291), .C(n_58339), .D(n_42307)
		, .Z(n_246995847));
	notech_ao4 i_69694236(.A(n_58274), .B(n_42241), .C(n_58371), .D(n_42273)
		, .Z(n_247095848));
	notech_and4 i_70294238(.A(n_247095848), .B(n_246995847), .C(n_246795845)
		, .D(n_246695844), .Z(n_247295850));
	notech_ao4 i_72194240(.A(n_58307), .B(n_42266), .C(n_58291), .D(n_42282)
		, .Z(n_247495852));
	notech_ao4 i_72294242(.A(n_58241), .B(n_42250), .C(n_57963), .D(n_42421)
		, .Z(n_247695854));
	notech_ao4 i_72394243(.A(n_57995), .B(n_42389), .C(n_57979), .D(n_42405)
		, .Z(n_247795855));
	notech_and4 i_73294245(.A(n_247795855), .B(n_247695854), .C(n_247495852)
		, .D(n_163595013), .Z(n_247995857));
	notech_ao4 i_72494246(.A(n_58027), .B(n_42357), .C(n_58011), .D(n_42373)
		, .Z(n_248095858));
	notech_ao4 i_72594247(.A(n_58323), .B(n_42325), .C(n_58043), .D(n_42341)
		, .Z(n_248195859));
	notech_ao4 i_72694249(.A(n_58355), .B(n_42293), .C(n_58339), .D(n_42309)
		, .Z(n_248395861));
	notech_ao4 i_72794250(.A(n_58274), .B(n_42242), .C(n_58371), .D(n_42274)
		, .Z(n_248495862));
	notech_and4 i_73394252(.A(n_248495862), .B(n_248395861), .C(n_248195859)
		, .D(n_248095858), .Z(n_248695864));
	notech_ao4 i_75294254(.A(n_58307), .B(n_42267), .C(n_58291), .D(n_42283)
		, .Z(n_248895866));
	notech_ao4 i_75394256(.A(n_58241), .B(n_42251), .C(n_57963), .D(n_42423)
		, .Z(n_249095868));
	notech_ao4 i_75494257(.A(n_57995), .B(n_42391), .C(n_57979), .D(n_42407)
		, .Z(n_249195869));
	notech_and4 i_76394259(.A(n_249195869), .B(n_249095868), .C(n_248895866)
		, .D(n_165195029), .Z(n_249395871));
	notech_ao4 i_75594260(.A(n_58027), .B(n_42359), .C(n_58011), .D(n_42375)
		, .Z(n_249495872));
	notech_ao4 i_75694261(.A(n_58323), .B(n_42327), .C(n_58043), .D(n_42343)
		, .Z(n_249595873));
	notech_ao4 i_75794263(.A(n_58355), .B(n_42295), .C(n_58339), .D(n_42311)
		, .Z(n_249795875));
	notech_ao4 i_75894264(.A(n_58260), .B(n_42243), .C(n_58371), .D(n_42275)
		, .Z(n_249895876));
	notech_and4 i_76494266(.A(n_249895876), .B(n_249795875), .C(n_249595873)
		, .D(n_249495872), .Z(n_250095878));
	notech_ao4 i_78394268(.A(n_58307), .B(n_42268), .C(n_58291), .D(n_42284)
		, .Z(n_250295880));
	notech_ao4 i_78494270(.A(n_58241), .B(n_42252), .C(n_57963), .D(n_42425)
		, .Z(n_250495882));
	notech_ao4 i_78594271(.A(n_57995), .B(n_42393), .C(n_57979), .D(n_42409)
		, .Z(n_250595883));
	notech_and4 i_79494273(.A(n_250595883), .B(n_250495882), .C(n_250295880)
		, .D(n_166795045), .Z(n_250795885));
	notech_ao4 i_78694274(.A(n_58027), .B(n_42361), .C(n_58011), .D(n_42377)
		, .Z(n_250895886));
	notech_ao4 i_78794275(.A(n_58323), .B(n_42329), .C(n_58043), .D(n_42345)
		, .Z(n_250995887));
	notech_ao4 i_78894277(.A(n_58355), .B(n_42297), .C(n_58339), .D(n_42313)
		, .Z(n_251195889));
	notech_ao4 i_78994278(.A(n_58260), .B(n_42244), .C(n_58371), .D(n_42276)
		, .Z(n_251295890));
	notech_and4 i_79594280(.A(n_251295890), .B(n_251195889), .C(n_250995887)
		, .D(n_250895886), .Z(n_251495892));
	notech_ao4 i_81494282(.A(n_58295), .B(n_42269), .C(n_58279), .D(n_42285)
		, .Z(n_251695894));
	notech_ao4 i_81594284(.A(n_58242), .B(n_42253), .C(n_57951), .D(n_42427)
		, .Z(n_251895896));
	notech_ao4 i_81694285(.A(n_57983), .B(n_42395), .C(n_57967), .D(n_42411)
		, .Z(n_251995897));
	notech_and4 i_82594287(.A(n_251995897), .B(n_251895896), .C(n_251695894)
		, .D(n_168395061), .Z(n_252195899));
	notech_ao4 i_81794288(.A(n_58015), .B(n_42363), .C(n_57999), .D(n_42379)
		, .Z(n_252295900));
	notech_ao4 i_81894289(.A(n_58311), .B(n_42331), .C(n_58031), .D(n_42347)
		, .Z(n_252395901));
	notech_ao4 i_81994291(.A(n_58343), .B(n_42299), .C(n_58327), .D(n_42315)
		, .Z(n_252595903));
	notech_ao4 i_82094292(.A(n_58260), .B(n_42245), .C(n_58359), .D(n_42277)
		, .Z(n_252695904));
	notech_and4 i_82694294(.A(n_252695904), .B(n_252595903), .C(n_252395901)
		, .D(n_252295900), .Z(n_252895906));
	notech_ao4 i_90794296(.A(n_58295), .B(n_42272), .C(n_58279), .D(n_42288)
		, .Z(n_253095908));
	notech_ao4 i_90894298(.A(n_58242), .B(n_42256), .C(n_57951), .D(n_42433)
		, .Z(n_253295910));
	notech_ao4 i_90994299(.A(n_57983), .B(n_42401), .C(n_57967), .D(n_42417)
		, .Z(n_253395911));
	notech_and4 i_91894301(.A(n_253395911), .B(n_253295910), .C(n_253095908)
		, .D(n_169995077), .Z(n_253595913));
	notech_ao4 i_91094302(.A(n_58015), .B(n_42369), .C(n_57999), .D(n_42385)
		, .Z(n_253695914));
	notech_ao4 i_91194303(.A(n_58311), .B(n_42337), .C(n_58031), .D(n_42353)
		, .Z(n_253795915));
	notech_ao4 i_91294305(.A(n_58343), .B(n_42305), .C(n_58327), .D(n_42321)
		, .Z(n_253995917));
	notech_ao4 i_91394306(.A(n_58260), .B(n_42248), .C(n_58359), .D(n_42280)
		, .Z(n_254095918));
	notech_and4 i_91994308(.A(n_254095918), .B(n_253995917), .C(n_253795915)
		, .D(n_253695914), .Z(n_254295920));
	notech_ao4 i_93894310(.A(n_58295), .B(n_42273), .C(n_58279), .D(n_42291)
		, .Z(n_254495922));
	notech_ao4 i_93994312(.A(n_58242), .B(n_42257), .C(n_57951), .D(n_42435)
		, .Z(n_254695924));
	notech_ao4 i_94094313(.A(n_57983), .B(n_42403), .C(n_57967), .D(n_42419)
		, .Z(n_254795925));
	notech_and4 i_94994315(.A(n_254795925), .B(n_254695924), .C(n_254495922)
		, .D(n_171595093), .Z(n_254995927));
	notech_ao4 i_94194316(.A(n_58015), .B(n_42371), .C(n_57999), .D(n_42387)
		, .Z(n_255095928));
	notech_ao4 i_94294317(.A(n_58311), .B(n_42339), .C(n_58031), .D(n_42355)
		, .Z(n_255195929));
	notech_ao4 i_94394319(.A(n_58343), .B(n_42307), .C(n_58327), .D(n_42323)
		, .Z(n_255395931));
	notech_ao4 i_94494320(.A(n_58260), .B(n_42249), .C(n_58359), .D(n_42281)
		, .Z(n_255495932));
	notech_and4 i_95094322(.A(n_255495932), .B(n_255395931), .C(n_255195929)
		, .D(n_255095928), .Z(n_255695934));
	notech_ao4 i_96994324(.A(n_58295), .B(n_42274), .C(n_58279), .D(n_42293)
		, .Z(n_255895936));
	notech_ao4 i_97094326(.A(n_58242), .B(n_42258), .C(n_57951), .D(n_42437)
		, .Z(n_256095938));
	notech_ao4 i_97194327(.A(n_57983), .B(n_42405), .C(n_57967), .D(n_42421)
		, .Z(n_256195939));
	notech_and4 i_98094329(.A(n_256195939), .B(n_256095938), .C(n_255895936)
		, .D(n_173195109), .Z(n_256395941));
	notech_ao4 i_97294330(.A(n_58015), .B(n_42373), .C(n_57999), .D(n_42389)
		, .Z(n_256495942));
	notech_ao4 i_97394331(.A(n_58311), .B(n_42341), .C(n_58031), .D(n_42357)
		, .Z(n_256595943));
	notech_ao4 i_97494333(.A(n_58343), .B(n_42309), .C(n_58327), .D(n_42325)
		, .Z(n_256795945));
	notech_ao4 i_97594334(.A(n_58260), .B(n_42250), .C(n_58359), .D(n_42282)
		, .Z(n_256895946));
	notech_and4 i_98194336(.A(n_256895946), .B(n_256795945), .C(n_256595943)
		, .D(n_256495942), .Z(n_257095948));
	notech_ao4 i_100094338(.A(n_58295), .B(n_42275), .C(n_58279), .D(n_42295
		), .Z(n_257295950));
	notech_ao4 i_100194340(.A(n_58242), .B(n_42259), .C(n_57951), .D(n_42439
		), .Z(n_257495952));
	notech_ao4 i_100294341(.A(n_57983), .B(n_42407), .C(n_57967), .D(n_42423
		), .Z(n_257595953));
	notech_and4 i_101194343(.A(n_257595953), .B(n_257495952), .C(n_257295950
		), .D(n_174795125), .Z(n_257795955));
	notech_ao4 i_100394344(.A(n_58015), .B(n_42375), .C(n_57999), .D(n_42391
		), .Z(n_257895956));
	notech_ao4 i_100494345(.A(n_58311), .B(n_42343), .C(n_58031), .D(n_42359
		), .Z(n_257995957));
	notech_ao4 i_100594347(.A(n_58343), .B(n_42311), .C(n_58327), .D(n_42327
		), .Z(n_258195959));
	notech_ao4 i_100694348(.A(n_58266), .B(n_42251), .C(n_58359), .D(n_42283
		), .Z(n_258295960));
	notech_and4 i_101294350(.A(n_258295960), .B(n_258195959), .C(n_257995957
		), .D(n_257895956), .Z(n_258495962));
	notech_ao4 i_103194352(.A(n_58295), .B(n_42276), .C(n_58279), .D(n_42297
		), .Z(n_258695964));
	notech_ao4 i_103294354(.A(n_58242), .B(n_42260), .C(n_57951), .D(n_42441
		), .Z(n_258895966));
	notech_ao4 i_103394355(.A(n_57983), .B(n_42409), .C(n_57967), .D(n_42425
		), .Z(n_258995967));
	notech_and4 i_104294357(.A(n_258995967), .B(n_258895966), .C(n_258695964
		), .D(n_176395141), .Z(n_259195969));
	notech_ao4 i_103494358(.A(n_58015), .B(n_42377), .C(n_57999), .D(n_42393
		), .Z(n_259295970));
	notech_ao4 i_103594359(.A(n_58311), .B(n_42345), .C(n_58031), .D(n_42361
		), .Z(n_259395971));
	notech_ao4 i_103694361(.A(n_58343), .B(n_42313), .C(n_58327), .D(n_42329
		), .Z(n_259595973));
	notech_ao4 i_103794362(.A(n_58266), .B(n_42252), .C(n_58359), .D(n_42284
		), .Z(n_259695974));
	notech_and4 i_104394364(.A(n_259695974), .B(n_259595973), .C(n_259395971
		), .D(n_259295970), .Z(n_259895976));
	notech_ao4 i_106294366(.A(n_58305), .B(n_42277), .C(n_58289), .D(n_42299
		), .Z(n_260095978));
	notech_ao4 i_106394368(.A(n_58242), .B(n_42261), .C(n_57961), .D(n_42443
		), .Z(n_260295980));
	notech_ao4 i_106494369(.A(n_57993), .B(n_42411), .C(n_57977), .D(n_42427
		), .Z(n_260395981));
	notech_and4 i_107394371(.A(n_260395981), .B(n_260295980), .C(n_260095978
		), .D(n_177995157), .Z(n_260595983));
	notech_ao4 i_106594372(.A(n_58025), .B(n_42379), .C(n_58009), .D(n_42395
		), .Z(n_260695984));
	notech_ao4 i_106694373(.A(n_58321), .B(n_42347), .C(n_58041), .D(n_42363
		), .Z(n_260795985));
	notech_ao4 i_106794375(.A(n_58353), .B(n_42315), .C(n_58337), .D(n_42331
		), .Z(n_260995987));
	notech_ao4 i_106894376(.A(n_58266), .B(n_42253), .C(n_58369), .D(n_42285
		), .Z(n_261095988));
	notech_and4 i_107494378(.A(n_261095988), .B(n_260995987), .C(n_260795985
		), .D(n_260695984), .Z(n_261295990));
	notech_ao4 i_115594380(.A(n_58295), .B(n_42280), .C(n_58279), .D(n_42305
		), .Z(n_261495992));
	notech_ao4 i_115694382(.A(n_58242), .B(n_42264), .C(n_57951), .D(n_42449
		), .Z(n_261695994));
	notech_ao4 i_115794383(.A(n_57983), .B(n_42417), .C(n_57967), .D(n_42433
		), .Z(n_261795995));
	notech_and4 i_116694385(.A(n_261795995), .B(n_261695994), .C(n_261495992
		), .D(n_179595173), .Z(n_261995997));
	notech_ao4 i_115894386(.A(n_58015), .B(n_42385), .C(n_57999), .D(n_42401
		), .Z(n_262095998));
	notech_ao4 i_115994387(.A(n_58311), .B(n_42353), .C(n_58031), .D(n_42369
		), .Z(n_262195999));
	notech_ao4 i_116094389(.A(n_58343), .B(n_42321), .C(n_58327), .D(n_42337
		), .Z(n_262396001));
	notech_ao4 i_116194390(.A(n_58260), .B(n_42256), .C(n_58359), .D(n_42288
		), .Z(n_262496002));
	notech_and4 i_116794392(.A(n_262496002), .B(n_262396001), .C(n_262195999
		), .D(n_262095998), .Z(n_262696004));
	notech_ao4 i_118694394(.A(n_58295), .B(n_42281), .C(n_58279), .D(n_42307
		), .Z(n_262896006));
	notech_ao4 i_118794396(.A(n_58247), .B(n_42265), .C(n_57951), .D(n_42451
		), .Z(n_263096008));
	notech_ao4 i_118894397(.A(n_57983), .B(n_42419), .C(n_57967), .D(n_42435
		), .Z(n_263196009));
	notech_and4 i_119794399(.A(n_263196009), .B(n_263096008), .C(n_262896006
		), .D(n_181195189), .Z(n_263396011));
	notech_ao4 i_118994400(.A(n_58015), .B(n_42387), .C(n_57999), .D(n_42403
		), .Z(n_263496012));
	notech_ao4 i_119094401(.A(n_58311), .B(n_42355), .C(n_58031), .D(n_42371
		), .Z(n_263596013));
	notech_ao4 i_119194403(.A(n_58343), .B(n_42323), .C(n_58327), .D(n_42339
		), .Z(n_263796015));
	notech_ao4 i_119294404(.A(n_58266), .B(n_42257), .C(n_58359), .D(n_42291
		), .Z(n_263896016));
	notech_and4 i_119894406(.A(n_263896016), .B(n_263796015), .C(n_263596013
		), .D(n_263496012), .Z(n_264096018));
	notech_ao4 i_121794408(.A(n_58295), .B(n_42282), .C(n_58279), .D(n_42309
		), .Z(n_264296020));
	notech_ao4 i_121894410(.A(n_58247), .B(n_42266), .C(n_57951), .D(n_42453
		), .Z(n_264496022));
	notech_ao4 i_121994411(.A(n_57983), .B(n_42421), .C(n_57967), .D(n_42437
		), .Z(n_264596023));
	notech_and4 i_122894413(.A(n_264596023), .B(n_264496022), .C(n_264296020
		), .D(n_182795205), .Z(n_264796025));
	notech_ao4 i_122094414(.A(n_58015), .B(n_42389), .C(n_57999), .D(n_42405
		), .Z(n_264896026));
	notech_ao4 i_122194415(.A(n_58311), .B(n_42357), .C(n_58031), .D(n_42373
		), .Z(n_264996027));
	notech_ao4 i_122294417(.A(n_58343), .B(n_42325), .C(n_58327), .D(n_42341
		), .Z(n_265196029));
	notech_ao4 i_122394418(.A(n_58260), .B(n_42258), .C(n_58359), .D(n_42293
		), .Z(n_265296030));
	notech_and4 i_122994420(.A(n_265296030), .B(n_265196029), .C(n_264996027
		), .D(n_264896026), .Z(n_265496032));
	notech_ao4 i_124894422(.A(n_58295), .B(n_42283), .C(n_58279), .D(n_42311
		), .Z(n_265696034));
	notech_ao4 i_124994424(.A(n_58247), .B(n_42267), .C(n_57951), .D(n_42455
		), .Z(n_265896036));
	notech_ao4 i_125094425(.A(n_57983), .B(n_42423), .C(n_57967), .D(n_42439
		), .Z(n_265996037));
	notech_and4 i_125994427(.A(n_265996037), .B(n_265896036), .C(n_265696034
		), .D(n_184395221), .Z(n_266196039));
	notech_ao4 i_125194428(.A(n_58015), .B(n_42391), .C(n_57999), .D(n_42407
		), .Z(n_266296040));
	notech_ao4 i_125294429(.A(n_58311), .B(n_42359), .C(n_58031), .D(n_42375
		), .Z(n_266396041));
	notech_ao4 i_125394431(.A(n_58343), .B(n_42327), .C(n_58327), .D(n_42343
		), .Z(n_266596043));
	notech_ao4 i_125494432(.A(n_58260), .B(n_42259), .C(n_58359), .D(n_42295
		), .Z(n_266696044));
	notech_and4 i_126094434(.A(n_266696044), .B(n_266596043), .C(n_266396041
		), .D(n_266296040), .Z(n_266896046));
	notech_ao4 i_127994436(.A(n_58295), .B(n_42284), .C(n_58279), .D(n_42313
		), .Z(n_267096048));
	notech_ao4 i_128094438(.A(n_58247), .B(n_42268), .C(n_57951), .D(n_42457
		), .Z(n_267296050));
	notech_ao4 i_128194439(.A(n_57983), .B(n_42425), .C(n_57967), .D(n_42441
		), .Z(n_267396051));
	notech_and4 i_129094441(.A(n_267396051), .B(n_267296050), .C(n_267096048
		), .D(n_185995237), .Z(n_267596053));
	notech_ao4 i_128294442(.A(n_58015), .B(n_42393), .C(n_57999), .D(n_42409
		), .Z(n_267696054));
	notech_ao4 i_128394443(.A(n_58311), .B(n_42361), .C(n_58031), .D(n_42377
		), .Z(n_267796055));
	notech_ao4 i_128494445(.A(n_58343), .B(n_42329), .C(n_58327), .D(n_42345
		), .Z(n_267996057));
	notech_ao4 i_128594446(.A(n_58260), .B(n_42260), .C(n_58359), .D(n_42297
		), .Z(n_268096058));
	notech_and4 i_129194448(.A(n_268096058), .B(n_267996057), .C(n_267796055
		), .D(n_267696054), .Z(n_268296060));
	notech_ao4 i_131094450(.A(n_58295), .B(n_42285), .C(n_58279), .D(n_42315
		), .Z(n_268496062));
	notech_ao4 i_131194452(.A(n_58247), .B(n_42269), .C(n_57951), .D(n_42459
		), .Z(n_268696064));
	notech_ao4 i_131294453(.A(n_57983), .B(n_42427), .C(n_57967), .D(n_42443
		), .Z(n_268796065));
	notech_and4 i_132194455(.A(n_268796065), .B(n_268696064), .C(n_268496062
		), .D(n_187595253), .Z(n_268996067));
	notech_ao4 i_131394456(.A(n_58015), .B(n_42395), .C(n_57999), .D(n_42411
		), .Z(n_269096068));
	notech_ao4 i_131494457(.A(n_58311), .B(n_42363), .C(n_58031), .D(n_42379
		), .Z(n_269196069));
	notech_ao4 i_131594459(.A(n_58343), .B(n_42331), .C(n_58327), .D(n_42347
		), .Z(n_269396071));
	notech_ao4 i_131694460(.A(n_58260), .B(n_42261), .C(n_58359), .D(n_42299
		), .Z(n_269496072));
	notech_and4 i_132294462(.A(n_269496072), .B(n_269396071), .C(n_269196069
		), .D(n_269096068), .Z(n_269696074));
	notech_ao4 i_140394464(.A(n_58295), .B(n_42288), .C(n_58279), .D(n_42321
		), .Z(n_269896076));
	notech_ao4 i_140494466(.A(n_58247), .B(n_42272), .C(n_57951), .D(n_42465
		), .Z(n_270096078));
	notech_ao4 i_140594467(.A(n_57983), .B(n_42433), .C(n_57967), .D(n_42449
		), .Z(n_270196079));
	notech_and4 i_141494469(.A(n_270196079), .B(n_270096078), .C(n_269896076
		), .D(n_189195269), .Z(n_270396081));
	notech_ao4 i_140694470(.A(n_58015), .B(n_42401), .C(n_57999), .D(n_42417
		), .Z(n_270496082));
	notech_ao4 i_140794471(.A(n_58311), .B(n_42369), .C(n_58031), .D(n_42385
		), .Z(n_270596083));
	notech_ao4 i_140894473(.A(n_58343), .B(n_42337), .C(n_58327), .D(n_42353
		), .Z(n_270796085));
	notech_ao4 i_140994474(.A(n_58260), .B(n_42264), .C(n_58359), .D(n_42305
		), .Z(n_270896086));
	notech_and4 i_141594476(.A(n_270896086), .B(n_270796085), .C(n_270596083
		), .D(n_270496082), .Z(n_271096088));
	notech_ao4 i_143494478(.A(n_58295), .B(n_42291), .C(n_58279), .D(n_42323
		), .Z(n_271296090));
	notech_ao4 i_143594480(.A(n_58247), .B(n_42273), .C(n_57951), .D(n_42467
		), .Z(n_271496092));
	notech_ao4 i_143694481(.A(n_57983), .B(n_42435), .C(n_57967), .D(n_42451
		), .Z(n_271596093));
	notech_and4 i_144594483(.A(n_271596093), .B(n_271496092), .C(n_271296090
		), .D(n_190795285), .Z(n_271796095));
	notech_ao4 i_143794484(.A(n_58015), .B(n_42403), .C(n_57999), .D(n_42419
		), .Z(n_271896096));
	notech_ao4 i_143894485(.A(n_58311), .B(n_42371), .C(n_58031), .D(n_42387
		), .Z(n_271996097));
	notech_ao4 i_143994487(.A(n_58343), .B(n_42339), .C(n_58327), .D(n_42355
		), .Z(n_272196099));
	notech_ao4 i_144094488(.A(n_58260), .B(n_42265), .C(n_58359), .D(n_42307
		), .Z(n_272296100));
	notech_and4 i_144694490(.A(n_272296100), .B(n_272196099), .C(n_271996097
		), .D(n_271896096), .Z(n_272496102));
	notech_ao4 i_146594492(.A(n_58295), .B(n_42293), .C(n_58279), .D(n_42325
		), .Z(n_272696104));
	notech_ao4 i_146694494(.A(n_58247), .B(n_42274), .C(n_57951), .D(n_42469
		), .Z(n_272896106));
	notech_ao4 i_146794495(.A(n_57983), .B(n_42437), .C(n_57967), .D(n_42453
		), .Z(n_272996107));
	notech_and4 i_147694497(.A(n_272996107), .B(n_272896106), .C(n_272696104
		), .D(n_192395301), .Z(n_273196109));
	notech_ao4 i_146894498(.A(n_58015), .B(n_42405), .C(n_57999), .D(n_42421
		), .Z(n_273296110));
	notech_ao4 i_146994499(.A(n_58311), .B(n_42373), .C(n_58031), .D(n_42389
		), .Z(n_273396111));
	notech_ao4 i_147094501(.A(n_58343), .B(n_42341), .C(n_58327), .D(n_42357
		), .Z(n_273596113));
	notech_ao4 i_147194502(.A(n_58260), .B(n_42266), .C(n_58359), .D(n_42309
		), .Z(n_273696114));
	notech_and4 i_147794504(.A(n_273696114), .B(n_273596113), .C(n_273396111
		), .D(n_273296110), .Z(n_273896116));
	notech_ao4 i_149694506(.A(n_58295), .B(n_42295), .C(n_58279), .D(n_42327
		), .Z(n_274096118));
	notech_ao4 i_149794508(.A(n_58249), .B(n_42275), .C(n_57951), .D(n_42471
		), .Z(n_274296120));
	notech_ao4 i_149894509(.A(n_57983), .B(n_42439), .C(n_57967), .D(n_42455
		), .Z(n_274396121));
	notech_and4 i_150794511(.A(n_274396121), .B(n_274296120), .C(n_274096118
		), .D(n_193995317), .Z(n_274596123));
	notech_ao4 i_149994512(.A(n_58015), .B(n_42407), .C(n_57999), .D(n_42423
		), .Z(n_274696124));
	notech_ao4 i_150094513(.A(n_58311), .B(n_42375), .C(n_58031), .D(n_42391
		), .Z(n_274796125));
	notech_ao4 i_150194515(.A(n_58343), .B(n_42343), .C(n_58327), .D(n_42359
		), .Z(n_274996127));
	notech_ao4 i_150294516(.A(n_58260), .B(n_42267), .C(n_58359), .D(n_42311
		), .Z(n_275096128));
	notech_and4 i_150894518(.A(n_275096128), .B(n_274996127), .C(n_274796125
		), .D(n_274696124), .Z(n_275296130));
	notech_ao4 i_152794520(.A(n_58295), .B(n_42297), .C(n_58279), .D(n_42329
		), .Z(n_275496132));
	notech_ao4 i_152894522(.A(n_58249), .B(n_42276), .C(n_57951), .D(n_42473
		), .Z(n_275696134));
	notech_ao4 i_152994523(.A(n_57983), .B(n_42441), .C(n_57967), .D(n_42457
		), .Z(n_275796135));
	notech_and4 i_153894525(.A(n_275796135), .B(n_275696134), .C(n_275496132
		), .D(n_195595333), .Z(n_275996137));
	notech_ao4 i_153094526(.A(n_58015), .B(n_42409), .C(n_57999), .D(n_42425
		), .Z(n_276096138));
	notech_ao4 i_153194527(.A(n_58311), .B(n_42377), .C(n_58031), .D(n_42393
		), .Z(n_276196139));
	notech_ao4 i_153294529(.A(n_58343), .B(n_42345), .C(n_58327), .D(n_42361
		), .Z(n_276396141));
	notech_ao4 i_153394530(.A(n_58260), .B(n_42268), .C(n_58359), .D(n_42313
		), .Z(n_276496142));
	notech_and4 i_153994532(.A(n_276496142), .B(n_276396141), .C(n_276196139
		), .D(n_276096138), .Z(n_276696144));
	notech_ao4 i_155894534(.A(n_58295), .B(n_42299), .C(n_58279), .D(n_42331
		), .Z(n_276896146));
	notech_ao4 i_155994535(.A(n_58249), .B(n_42277), .C(n_57951), .D(n_42475
		), .Z(n_277096148));
	notech_ao4 i_156094536(.A(n_57983), .B(n_42443), .C(n_57967), .D(n_42459
		), .Z(n_277196149));
	notech_and4 i_1569(.A(n_277196149), .B(n_277096148), .C(n_276896146), .D
		(n_197195349), .Z(n_277396151));
	notech_ao4 i_156194537(.A(n_58015), .B(n_42411), .C(n_57999), .D(n_42427
		), .Z(n_277496152));
	notech_ao4 i_156294538(.A(n_58311), .B(n_42379), .C(n_58031), .D(n_42395
		), .Z(n_277596153));
	notech_ao4 i_1563(.A(n_58343), .B(n_42347), .C(n_58327), .D(n_42363), .Z
		(n_277796155));
	notech_ao4 i_1564(.A(n_58260), .B(n_42269), .C(n_58359), .D(n_42315), .Z
		(n_277896156));
	notech_and4 i_1570(.A(n_277896156), .B(n_277796155), .C(n_277596153), .D
		(n_277496152), .Z(n_278096158));
	notech_ao4 i_1651(.A(n_58305), .B(n_42305), .C(n_58289), .D(n_42337), .Z
		(n_278296160));
	notech_ao4 i_1652(.A(n_58249), .B(n_42280), .C(n_57961), .D(n_42481), .Z
		(n_278496162));
	notech_ao4 i_1653(.A(n_57993), .B(n_42449), .C(n_57977), .D(n_42465), .Z
		(n_278596163));
	notech_and4 i_1662(.A(n_278596163), .B(n_278496162), .C(n_278296160), .D
		(n_198795365), .Z(n_278796165));
	notech_ao4 i_1654(.A(n_58025), .B(n_42417), .C(n_58009), .D(n_42433), .Z
		(n_278896166));
	notech_ao4 i_1655(.A(n_58321), .B(n_42385), .C(n_58041), .D(n_42401), .Z
		(n_278996167));
	notech_ao4 i_1656(.A(n_58353), .B(n_42353), .C(n_58337), .D(n_42369), .Z
		(n_279196169));
	notech_ao4 i_1657(.A(n_58260), .B(n_42272), .C(n_58369), .D(n_42321), .Z
		(n_279296170));
	notech_and4 i_1663(.A(n_279296170), .B(n_279196169), .C(n_278996167), .D
		(n_278896166), .Z(n_279496172));
	notech_ao4 i_1682(.A(n_58301), .B(n_42307), .C(n_58285), .D(n_42339), .Z
		(n_279696174));
	notech_ao4 i_1683(.A(n_58249), .B(n_42281), .C(n_57957), .D(n_42483), .Z
		(n_279896176));
	notech_ao4 i_1684(.A(n_57989), .B(n_42451), .C(n_57973), .D(n_42467), .Z
		(n_279996177));
	notech_and4 i_1693(.A(n_279996177), .B(n_279896176), .C(n_279696174), .D
		(n_200395381), .Z(n_280196179));
	notech_ao4 i_1685(.A(n_58021), .B(n_42419), .C(n_58005), .D(n_42435), .Z
		(n_280296180));
	notech_ao4 i_1686(.A(n_58317), .B(n_42387), .C(n_58037), .D(n_42403), .Z
		(n_280396181));
	notech_ao4 i_1687(.A(n_58349), .B(n_42355), .C(n_58333), .D(n_42371), .Z
		(n_280596183));
	notech_ao4 i_1688(.A(n_58266), .B(n_42273), .C(n_58365), .D(n_42323), .Z
		(n_280696184));
	notech_and4 i_1694(.A(n_280696184), .B(n_280596183), .C(n_280396181), .D
		(n_280296180), .Z(n_280896186));
	notech_ao4 i_1713(.A(n_58301), .B(n_42309), .C(n_58285), .D(n_42341), .Z
		(n_281096188));
	notech_ao4 i_1714(.A(n_58247), .B(n_42282), .C(n_57957), .D(n_42485), .Z
		(n_281296190));
	notech_ao4 i_1715(.A(n_57989), .B(n_42453), .C(n_57973), .D(n_42469), .Z
		(n_281396191));
	notech_and4 i_1724(.A(n_281396191), .B(n_281296190), .C(n_281096188), .D
		(n_201995397), .Z(n_281596193));
	notech_ao4 i_1716(.A(n_58021), .B(n_42421), .C(n_58005), .D(n_42437), .Z
		(n_281696194));
	notech_ao4 i_1717(.A(n_58317), .B(n_42389), .C(n_58037), .D(n_42405), .Z
		(n_281796195));
	notech_ao4 i_1718(.A(n_58349), .B(n_42357), .C(n_58333), .D(n_42373), .Z
		(n_281996197));
	notech_ao4 i_1719(.A(n_58267), .B(n_42274), .C(n_58365), .D(n_42325), .Z
		(n_282096198));
	notech_and4 i_1725(.A(n_282096198), .B(n_281996197), .C(n_281796195), .D
		(n_281696194), .Z(n_282296200));
	notech_ao4 i_1744(.A(n_58301), .B(n_42311), .C(n_58285), .D(n_42343), .Z
		(n_282496202));
	notech_ao4 i_1745(.A(n_58249), .B(n_42283), .C(n_57957), .D(n_42487), .Z
		(n_282696204));
	notech_ao4 i_1746(.A(n_57989), .B(n_42455), .C(n_57973), .D(n_42471), .Z
		(n_282796205));
	notech_and4 i_1755(.A(n_282796205), .B(n_282696204), .C(n_282496202), .D
		(n_203595413), .Z(n_282996207));
	notech_ao4 i_1747(.A(n_58021), .B(n_42423), .C(n_58005), .D(n_42439), .Z
		(n_283096208));
	notech_ao4 i_1748(.A(n_58317), .B(n_42391), .C(n_58037), .D(n_42407), .Z
		(n_283196209));
	notech_ao4 i_1749(.A(n_58349), .B(n_42359), .C(n_58333), .D(n_42375), .Z
		(n_283396211));
	notech_ao4 i_1750(.A(n_58267), .B(n_42275), .C(n_58365), .D(n_42327), .Z
		(n_283496212));
	notech_and4 i_1756(.A(n_283496212), .B(n_283396211), .C(n_283196209), .D
		(n_283096208), .Z(n_283696214));
	notech_ao4 i_1775(.A(n_58301), .B(n_42313), .C(n_58285), .D(n_42345), .Z
		(n_283896216));
	notech_ao4 i_1776(.A(n_58249), .B(n_42284), .C(n_57957), .D(n_42489), .Z
		(n_284096218));
	notech_ao4 i_1777(.A(n_57989), .B(n_42457), .C(n_57973), .D(n_42473), .Z
		(n_284196219));
	notech_and4 i_1786(.A(n_284196219), .B(n_284096218), .C(n_283896216), .D
		(n_205195429), .Z(n_284396221));
	notech_ao4 i_1778(.A(n_58021), .B(n_42425), .C(n_58005), .D(n_42441), .Z
		(n_284496222));
	notech_ao4 i_1779(.A(n_58317), .B(n_42393), .C(n_58037), .D(n_42409), .Z
		(n_284596223));
	notech_ao4 i_1780(.A(n_58349), .B(n_42361), .C(n_58333), .D(n_42377), .Z
		(n_284796225));
	notech_ao4 i_1781(.A(n_58267), .B(n_42276), .C(n_58365), .D(n_42329), .Z
		(n_284896226));
	notech_and4 i_1787(.A(n_284896226), .B(n_284796225), .C(n_284596223), .D
		(n_284496222), .Z(n_285096228));
	notech_ao4 i_1806(.A(n_58301), .B(n_42315), .C(n_58285), .D(n_42347), .Z
		(n_285296230));
	notech_ao4 i_1807(.A(n_58244), .B(n_42285), .C(n_57957), .D(n_42491), .Z
		(n_285496232));
	notech_ao4 i_1808(.A(n_57989), .B(n_42459), .C(n_57973), .D(n_42475), .Z
		(n_285596233));
	notech_and4 i_1817(.A(n_285596233), .B(n_285496232), .C(n_285296230), .D
		(n_206795445), .Z(n_285796235));
	notech_ao4 i_1809(.A(n_58021), .B(n_42427), .C(n_58005), .D(n_42443), .Z
		(n_285896236));
	notech_ao4 i_1810(.A(n_58317), .B(n_42395), .C(n_58037), .D(n_42411), .Z
		(n_285996237));
	notech_ao4 i_1811(.A(n_58349), .B(n_42363), .C(n_58333), .D(n_42379), .Z
		(n_286196239));
	notech_ao4 i_1812(.A(n_58266), .B(n_42277), .C(n_58365), .D(n_42331), .Z
		(n_286296240));
	notech_and4 i_1818(.A(n_286296240), .B(n_286196239), .C(n_285996237), .D
		(n_285896236), .Z(n_286496242));
	notech_ao4 i_1899(.A(n_58301), .B(n_42321), .C(n_58285), .D(n_42353), .Z
		(n_286696244));
	notech_ao4 i_1900(.A(n_58244), .B(n_42288), .C(n_57957), .D(n_42497), .Z
		(n_286896246));
	notech_ao4 i_1901(.A(n_57989), .B(n_42465), .C(n_57973), .D(n_42481), .Z
		(n_286996247));
	notech_and4 i_1910(.A(n_286996247), .B(n_286896246), .C(n_286696244), .D
		(n_208395461), .Z(n_287196249));
	notech_ao4 i_1902(.A(n_58021), .B(n_42433), .C(n_58005), .D(n_42449), .Z
		(n_287296250));
	notech_ao4 i_1903(.A(n_58317), .B(n_42401), .C(n_58037), .D(n_42417), .Z
		(n_287396251));
	notech_ao4 i_1904(.A(n_58349), .B(n_42369), .C(n_58333), .D(n_42385), .Z
		(n_287596253));
	notech_ao4 i_1905(.A(n_58266), .B(n_42280), .C(n_58365), .D(n_42337), .Z
		(n_287696254));
	notech_and4 i_1911(.A(n_287696254), .B(n_287596253), .C(n_287396251), .D
		(n_287296250), .Z(n_287896256));
	notech_ao4 i_1930(.A(n_58301), .B(n_42323), .C(n_58285), .D(n_42355), .Z
		(n_288096258));
	notech_ao4 i_1931(.A(n_58244), .B(n_42291), .C(n_57957), .D(n_42499), .Z
		(n_288296260));
	notech_ao4 i_1932(.A(n_57989), .B(n_42467), .C(n_57973), .D(n_42483), .Z
		(n_288396261));
	notech_and4 i_1941(.A(n_288396261), .B(n_288296260), .C(n_288096258), .D
		(n_209995477), .Z(n_288596263));
	notech_ao4 i_1933(.A(n_58021), .B(n_42435), .C(n_58005), .D(n_42451), .Z
		(n_288696264));
	notech_ao4 i_1934(.A(n_58317), .B(n_42403), .C(n_58037), .D(n_42419), .Z
		(n_288796265));
	notech_ao4 i_1935(.A(n_58349), .B(n_42371), .C(n_58333), .D(n_42387), .Z
		(n_288996267));
	notech_ao4 i_1936(.A(n_58267), .B(n_42281), .C(n_58365), .D(n_42339), .Z
		(n_289096268));
	notech_and4 i_1942(.A(n_289096268), .B(n_288996267), .C(n_288796265), .D
		(n_288696264), .Z(n_289296270));
	notech_ao4 i_1961(.A(n_58301), .B(n_42325), .C(n_58285), .D(n_42357), .Z
		(n_289496272));
	notech_ao4 i_1962(.A(n_58244), .B(n_42293), .C(n_57957), .D(n_42501), .Z
		(n_289696274));
	notech_ao4 i_1963(.A(n_57989), .B(n_42469), .C(n_57973), .D(n_42485), .Z
		(n_289796275));
	notech_and4 i_1972(.A(n_289796275), .B(n_289696274), .C(n_289496272), .D
		(n_211595493), .Z(n_289996277));
	notech_ao4 i_1964(.A(n_58021), .B(n_42437), .C(n_58005), .D(n_42453), .Z
		(n_290096278));
	notech_ao4 i_1965(.A(n_58317), .B(n_42405), .C(n_58037), .D(n_42421), .Z
		(n_290196279));
	notech_ao4 i_1966(.A(n_58349), .B(n_42373), .C(n_58333), .D(n_42389), .Z
		(n_290396281));
	notech_ao4 i_1967(.A(n_58267), .B(n_42282), .C(n_58365), .D(n_42341), .Z
		(n_290496282));
	notech_and4 i_1973(.A(n_290496282), .B(n_290396281), .C(n_290196279), .D
		(n_290096278), .Z(n_290696284));
	notech_ao4 i_1992(.A(n_58301), .B(n_42327), .C(n_58285), .D(n_42359), .Z
		(n_290896286));
	notech_ao4 i_1993(.A(n_58244), .B(n_42295), .C(n_57957), .D(n_42503), .Z
		(n_291096288));
	notech_ao4 i_1994(.A(n_57989), .B(n_42471), .C(n_57973), .D(n_42487), .Z
		(n_291196289));
	notech_and4 i_2003(.A(n_291196289), .B(n_291096288), .C(n_290896286), .D
		(n_213195509), .Z(n_291396291));
	notech_ao4 i_1995(.A(n_58021), .B(n_42439), .C(n_58005), .D(n_42455), .Z
		(n_291496292));
	notech_ao4 i_1996(.A(n_58317), .B(n_42407), .C(n_58037), .D(n_42423), .Z
		(n_291596293));
	notech_ao4 i_1997(.A(n_58349), .B(n_42375), .C(n_58333), .D(n_42391), .Z
		(n_291796295));
	notech_ao4 i_1998(.A(n_58267), .B(n_42283), .C(n_58365), .D(n_42343), .Z
		(n_291896296));
	notech_and4 i_2004(.A(n_291896296), .B(n_291796295), .C(n_291596293), .D
		(n_291496292), .Z(n_292096298));
	notech_ao4 i_2023(.A(n_58307), .B(n_42329), .C(n_58291), .D(n_42361), .Z
		(n_292296300));
	notech_ao4 i_2024(.A(n_58244), .B(n_42297), .C(n_57963), .D(n_42505), .Z
		(n_292496302));
	notech_ao4 i_2025(.A(n_57995), .B(n_42473), .C(n_57979), .D(n_42489), .Z
		(n_292596303));
	notech_and4 i_2034(.A(n_292596303), .B(n_292496302), .C(n_292296300), .D
		(n_214795525), .Z(n_292796305));
	notech_ao4 i_2026(.A(n_58027), .B(n_42441), .C(n_58011), .D(n_42457), .Z
		(n_292896306));
	notech_ao4 i_2027(.A(n_58323), .B(n_42409), .C(n_58043), .D(n_42425), .Z
		(n_292996307));
	notech_ao4 i_2028(.A(n_58355), .B(n_42377), .C(n_58339), .D(n_42393), .Z
		(n_293196309));
	notech_ao4 i_2029(.A(n_58267), .B(n_42284), .C(n_58371), .D(n_42345), .Z
		(n_293296310));
	notech_and4 i_2035(.A(n_293296310), .B(n_293196309), .C(n_292996307), .D
		(n_292896306), .Z(n_293596312));
	notech_ao4 i_2054(.A(n_58305), .B(n_42331), .C(n_58289), .D(n_42363), .Z
		(n_293796314));
	notech_ao4 i_2055(.A(n_58244), .B(n_42299), .C(n_57961), .D(n_42507), .Z
		(n_293996316));
	notech_ao4 i_2056(.A(n_57993), .B(n_42475), .C(n_57977), .D(n_42491), .Z
		(n_294096317));
	notech_and4 i_2065(.A(n_294096317), .B(n_293996316), .C(n_293796314), .D
		(n_216395541), .Z(n_294496319));
	notech_ao4 i_2057(.A(n_58025), .B(n_42443), .C(n_58009), .D(n_42459), .Z
		(n_294796320));
	notech_ao4 i_2058(.A(n_58321), .B(n_42411), .C(n_58041), .D(n_42427), .Z
		(n_294896321));
	notech_ao4 i_2059(.A(n_58353), .B(n_42379), .C(n_58337), .D(n_42395), .Z
		(n_295096323));
	notech_ao4 i_2060(.A(n_58267), .B(n_42285), .C(n_58369), .D(n_42347), .Z
		(n_295196324));
	notech_and4 i_2066(.A(n_295196324), .B(n_295096323), .C(n_294896321), .D
		(n_294796320), .Z(n_295496326));
	notech_ao4 i_2147(.A(n_58305), .B(n_42337), .C(n_58289), .D(n_42369), .Z
		(n_295696328));
	notech_ao4 i_2148(.A(n_58244), .B(n_42305), .C(n_57961), .D(n_42513), .Z
		(n_295896330));
	notech_ao4 i_2149(.A(n_57993), .B(n_42481), .C(n_57977), .D(n_42497), .Z
		(n_295996331));
	notech_and4 i_2158(.A(n_295996331), .B(n_295896330), .C(n_295696328), .D
		(n_217995557), .Z(n_296196333));
	notech_ao4 i_2150(.A(n_58025), .B(n_42449), .C(n_58009), .D(n_42465), .Z
		(n_296296334));
	notech_ao4 i_2151(.A(n_58321), .B(n_42417), .C(n_58041), .D(n_42433), .Z
		(n_296396335));
	notech_ao4 i_2152(.A(n_58353), .B(n_42385), .C(n_58337), .D(n_42401), .Z
		(n_296696337));
	notech_ao4 i_2153(.A(n_58267), .B(n_42288), .C(n_58369), .D(n_42353), .Z
		(n_296796338));
	notech_and4 i_2159(.A(n_296796338), .B(n_296696337), .C(n_296396335), .D
		(n_296296334), .Z(n_296996340));
	notech_ao4 i_2178(.A(n_58305), .B(n_42339), .C(n_58289), .D(n_42371), .Z
		(n_297196342));
	notech_ao4 i_2179(.A(n_58247), .B(n_42307), .C(n_57961), .D(n_42515), .Z
		(n_297396344));
	notech_ao4 i_2180(.A(n_57993), .B(n_42483), .C(n_57977), .D(n_42499), .Z
		(n_297496345));
	notech_and4 i_2189(.A(n_297496345), .B(n_297396344), .C(n_297196342), .D
		(n_219595573), .Z(n_297696347));
	notech_ao4 i_2181(.A(n_58025), .B(n_42451), .C(n_58009), .D(n_42467), .Z
		(n_297796348));
	notech_ao4 i_2182(.A(n_58321), .B(n_42419), .C(n_58041), .D(n_42435), .Z
		(n_297896349));
	notech_ao4 i_2183(.A(n_58353), .B(n_42387), .C(n_58337), .D(n_42403), .Z
		(n_298096351));
	notech_ao4 i_2184(.A(n_58266), .B(n_42291), .C(n_58369), .D(n_42355), .Z
		(n_298196352));
	notech_and4 i_2190(.A(n_298196352), .B(n_298096351), .C(n_297896349), .D
		(n_297796348), .Z(n_298396354));
	notech_ao4 i_2209(.A(n_58305), .B(n_42341), .C(n_58289), .D(n_42373), .Z
		(n_298596356));
	notech_ao4 i_2210(.A(n_58247), .B(n_42309), .C(n_57961), .D(n_42517), .Z
		(n_298796358));
	notech_ao4 i_2211(.A(n_57993), .B(n_42485), .C(n_57977), .D(n_42501), .Z
		(n_298896359));
	notech_and4 i_2220(.A(n_298896359), .B(n_298796358), .C(n_298596356), .D
		(n_221195589), .Z(n_299096361));
	notech_ao4 i_2212(.A(n_58025), .B(n_42453), .C(n_58009), .D(n_42469), .Z
		(n_299196362));
	notech_ao4 i_2213(.A(n_58321), .B(n_42421), .C(n_58041), .D(n_42437), .Z
		(n_299296363));
	notech_ao4 i_2214(.A(n_58353), .B(n_42389), .C(n_58337), .D(n_42405), .Z
		(n_299496365));
	notech_ao4 i_2215(.A(n_58266), .B(n_42293), .C(n_58369), .D(n_42357), .Z
		(n_299596366));
	notech_and4 i_2221(.A(n_299596366), .B(n_299496365), .C(n_299296363), .D
		(n_299196362), .Z(n_299796368));
	notech_ao4 i_2240(.A(n_58307), .B(n_42343), .C(n_58291), .D(n_42375), .Z
		(n_299996370));
	notech_ao4 i_2241(.A(n_58247), .B(n_42311), .C(n_57963), .D(n_42519), .Z
		(n_300196372));
	notech_ao4 i_2242(.A(n_57995), .B(n_42487), .C(n_57979), .D(n_42503), .Z
		(n_300296373));
	notech_and4 i_2251(.A(n_300296373), .B(n_300196372), .C(n_299996370), .D
		(n_222795605), .Z(n_300496375));
	notech_ao4 i_2243(.A(n_58027), .B(n_42455), .C(n_58011), .D(n_42471), .Z
		(n_300596376));
	notech_ao4 i_2244(.A(n_58323), .B(n_42423), .C(n_58043), .D(n_42439), .Z
		(n_300696377));
	notech_ao4 i_2245(.A(n_58355), .B(n_42391), .C(n_58339), .D(n_42407), .Z
		(n_300896379));
	notech_ao4 i_2246(.A(n_58266), .B(n_42295), .C(n_58371), .D(n_42359), .Z
		(n_300996380));
	notech_and4 i_2252(.A(n_300996380), .B(n_300896379), .C(n_300696377), .D
		(n_300596376), .Z(n_301196382));
	notech_ao4 i_2271(.A(n_58307), .B(n_42345), .C(n_58291), .D(n_42377), .Z
		(n_301396384));
	notech_ao4 i_2272(.A(n_58247), .B(n_42313), .C(n_57963), .D(n_42521), .Z
		(n_301596386));
	notech_ao4 i_2273(.A(n_57995), .B(n_42489), .C(n_57979), .D(n_42505), .Z
		(n_301696387));
	notech_and4 i_2282(.A(n_301696387), .B(n_301596386), .C(n_301396384), .D
		(n_224395621), .Z(n_301896389));
	notech_ao4 i_2274(.A(n_58027), .B(n_42457), .C(n_58011), .D(n_42473), .Z
		(n_301996390));
	notech_ao4 i_2275(.A(n_58323), .B(n_42425), .C(n_58043), .D(n_42441), .Z
		(n_302096391));
	notech_ao4 i_2276(.A(n_58355), .B(n_42393), .C(n_58339), .D(n_42409), .Z
		(n_302296393));
	notech_ao4 i_2277(.A(n_58266), .B(n_42297), .C(n_58371), .D(n_42361), .Z
		(n_302396394));
	notech_and4 i_2283(.A(n_302396394), .B(n_302296393), .C(n_302096391), .D
		(n_301996390), .Z(n_302596396));
	notech_ao4 i_2302(.A(n_58307), .B(n_42347), .C(n_58291), .D(n_42379), .Z
		(n_302796398));
	notech_ao4 i_2303(.A(n_58247), .B(n_42315), .C(n_57963), .D(n_42523), .Z
		(n_302996400));
	notech_ao4 i_2304(.A(n_57995), .B(n_42491), .C(n_57979), .D(n_42507), .Z
		(n_303096401));
	notech_and4 i_2313(.A(n_303096401), .B(n_302996400), .C(n_302796398), .D
		(n_225995637), .Z(n_303296403));
	notech_ao4 i_2305(.A(n_58027), .B(n_42459), .C(n_58011), .D(n_42475), .Z
		(n_303396404));
	notech_ao4 i_2306(.A(n_58323), .B(n_42427), .C(n_58043), .D(n_42443), .Z
		(n_303496405));
	notech_ao4 i_2307(.A(n_58355), .B(n_42395), .C(n_58339), .D(n_42411), .Z
		(n_303696407));
	notech_ao4 i_2308(.A(n_58266), .B(n_42299), .C(n_58371), .D(n_42363), .Z
		(n_303796408));
	notech_and4 i_2314(.A(n_303796408), .B(n_303696407), .C(n_303496405), .D
		(n_303396404), .Z(n_303996410));
	notech_ao4 i_2333(.A(n_58307), .B(n_42349), .C(n_58291), .D(n_42381), .Z
		(n_304196412));
	notech_ao4 i_2334(.A(n_58247), .B(n_42317), .C(n_57963), .D(n_42525), .Z
		(n_304396414));
	notech_ao4 i_2335(.A(n_57995), .B(n_42493), .C(n_57979), .D(n_42509), .Z
		(n_304496415));
	notech_and4 i_2344(.A(n_304496415), .B(n_304396414), .C(n_304196412), .D
		(n_227595653), .Z(n_304696417));
	notech_ao4 i_2336(.A(n_58027), .B(n_42461), .C(n_58011), .D(n_42477), .Z
		(n_304796418));
	notech_ao4 i_2337(.A(n_58323), .B(n_42429), .C(n_58043), .D(n_42445), .Z
		(n_304896419));
	notech_ao4 i_2338(.A(n_58355), .B(n_42397), .C(n_58339), .D(n_42413), .Z
		(n_305096421));
	notech_ao4 i_2339(.A(n_58266), .B(n_42301), .C(n_58371), .D(n_42365), .Z
		(n_305196422));
	notech_and4 i_2345(.A(n_305196422), .B(n_305096421), .C(n_304896419), .D
		(n_304796418), .Z(n_305396424));
	notech_ao4 i_2395(.A(n_58307), .B(n_42353), .C(n_58291), .D(n_42385), .Z
		(n_305596426));
	notech_ao4 i_2396(.A(n_58247), .B(n_42321), .C(n_57963), .D(n_42529), .Z
		(n_305796428));
	notech_ao4 i_2397(.A(n_57995), .B(n_42497), .C(n_57979), .D(n_42513), .Z
		(n_305896429));
	notech_and4 i_2406(.A(n_305896429), .B(n_305796428), .C(n_305596426), .D
		(n_229195669), .Z(n_306096431));
	notech_ao4 i_2398(.A(n_58027), .B(n_42465), .C(n_58011), .D(n_42481), .Z
		(n_306196432));
	notech_ao4 i_2399(.A(n_58323), .B(n_42433), .C(n_58043), .D(n_42449), .Z
		(n_306296433));
	notech_ao4 i_2400(.A(n_58355), .B(n_42401), .C(n_58339), .D(n_42417), .Z
		(n_306496435));
	notech_ao4 i_2401(.A(n_58266), .B(n_42305), .C(n_58371), .D(n_42369), .Z
		(n_306596436));
	notech_and4 i_2407(.A(n_306596436), .B(n_306496435), .C(n_306296433), .D
		(n_306196432), .Z(n_306796438));
	notech_nao3 i_65346(.A(n_32555629), .B(n_7789), .C(n_100094404), .Z(\nbus_12117[0] 
		));
	notech_nand3 i_65453(.A(n_99594399), .B(n_8293), .C(n_32555629), .Z(n_36824
		));
	notech_and4 i_64510(.A(n_7789), .B(n_32555629), .C(n_99894402), .D(n_99994403
		), .Z(\nbus_12114[0] ));
	notech_nand3 i_6679210(.A(n_309596466), .B(n_8293), .C(n_60400), .Z(n_32555629
		));
	notech_or4 i_6578717(.A(n_60400), .B(n_42167), .C(n_42168), .D(n_59995),
		 .Z(n_306996440));
	notech_nand3 i_2278661(.A(n_8293), .B(n_42741), .C(n_309596466), .Z(n_307096441
		));
	notech_and3 i_4278684(.A(n_42743), .B(n_42170), .C(n_59995), .Z(n_140853041
		));
	notech_nao3 i_7258(.A(pg_fault), .B(n_42742), .C(fault_wptr_en), .Z(n_8293
		));
	notech_or2 i_7178686(.A(n_101194415), .B(n_307096441), .Z(n_7789));
	notech_or4 i_3878683(.A(nbus_12105[5]), .B(nbus_12105[4]), .C(nbus_12105
		[6]), .D(n_141953052), .Z(n_141853051));
	notech_nand2 i_7259(.A(fault_wptr_en), .B(n_7792), .Z(n_309596466));
	notech_nao3 i_7261(.A(n_42602), .B(n_42601), .C(nbus_12105[6]), .Z(n_142753060
		));
	notech_nand2 i_211483(.A(code_ack), .B(n_61546), .Z(n_309696467));
	notech_nand2 i_1478669(.A(n_8293), .B(n_42741), .Z(n_142353056));
	notech_or2 i_92577766(.A(n_58266), .B(n_42200), .Z(n_1602));
	notech_and4 i_3125010(.A(n_2378), .B(n_2377), .C(n_2372), .D(n_2376), .Z
		(squeue_3097076));
	notech_nand3 i_90777784(.A(n_57937), .B(n_58209), .C(queue[30]), .Z(n_1599
		));
	notech_or2 i_89477797(.A(n_58266), .B(n_42199), .Z(n_1586));
	notech_and4 i_2925008(.A(n_2364), .B(n_2363), .C(n_2358), .D(n_2362), .Z
		(squeue_2897077));
	notech_nand3 i_87677815(.A(n_57937), .B(n_58209), .C(queue[28]), .Z(n_1583
		));
	notech_nand3 i_4279176(.A(code_ack), .B(n_61549), .C(n_8288), .Z(n_7796545
		));
	notech_ao3 i_17579048(.A(n_60243), .B(n_42741), .C(nbus_12105[4]), .Z(n_20596673
		));
	notech_xor2 i_3979179(.A(addrshft[4]), .B(n_46296930), .Z(n_26296730));
	notech_and2 i_27478949(.A(purge_cnt[10]), .B(purge), .Z(n_28996757));
	notech_or4 i_27678947(.A(n_59995), .B(n_307096441), .C(n_42165), .D(n_7792
		), .Z(n_29196759));
	notech_or4 i_3679182(.A(useq_ptr[3]), .B(useq_ptr[2]), .C(useq_ptr[1]), 
		.D(useq_ptr[0]), .Z(n_29296760));
	notech_and2 i_5013(.A(n_34630), .B(n_46396931), .Z(n_29396761));
	notech_and2 i_5014(.A(n_34632), .B(n_46396931), .Z(n_29496762));
	notech_and2 i_5015(.A(n_34634), .B(n_46396931), .Z(n_29596763));
	notech_and2 i_5016(.A(n_34636), .B(n_46396931), .Z(n_29696764));
	notech_and2 i_5017(.A(n_34638), .B(n_46396931), .Z(n_29796765));
	notech_and2 i_5018(.A(n_34640), .B(n_46396931), .Z(n_29896766));
	notech_and2 i_5019(.A(n_34642), .B(n_46396931), .Z(n_29996767));
	notech_and2 i_5020(.A(n_34644), .B(n_46396931), .Z(n_30096768));
	notech_and2 i_5021(.A(n_34646), .B(n_46396931), .Z(n_30196769));
	notech_and2 i_5022(.A(n_34648), .B(n_46396931), .Z(n_30296770));
	notech_and2 i_5023(.A(n_34650), .B(n_46396931), .Z(n_30396771));
	notech_nor2 i_5024(.A(n_60400), .B(wptr[0]), .Z(n_30496772));
	notech_and2 i_5037(.A(addr_0[0]), .B(n_42741), .Z(n_30596773));
	notech_and2 i_5041(.A(addr_0[1]), .B(n_42741), .Z(n_30696774));
	notech_and2 i_5042(.A(addr_0[2]), .B(n_42741), .Z(n_30796775));
	notech_and2 i_5043(.A(addr_0[3]), .B(n_42741), .Z(n_30896776));
	notech_and2 i_5047(.A(cacheD[148]), .B(n_7796545), .Z(codeWEN));
	notech_and2 i_333279212(.A(idata[0]), .B(cacheD[148]), .Z(cacheD[0]));
	notech_and2 i_333179213(.A(idata[1]), .B(cacheD[148]), .Z(cacheD[1]));
	notech_and2 i_333079214(.A(idata[2]), .B(cacheD[148]), .Z(cacheD[2]));
	notech_and2 i_332979215(.A(idata[3]), .B(cacheD[148]), .Z(cacheD[3]));
	notech_and2 i_332879216(.A(idata[4]), .B(cacheD[148]), .Z(cacheD[4]));
	notech_and2 i_332779217(.A(idata[5]), .B(cacheD[148]), .Z(cacheD[5]));
	notech_and2 i_332679218(.A(idata[6]), .B(cacheD[148]), .Z(cacheD[6]));
	notech_and2 i_332579219(.A(idata[7]), .B(cacheD[148]), .Z(cacheD[7]));
	notech_and2 i_332479220(.A(idata[8]), .B(cacheD[148]), .Z(cacheD[8]));
	notech_and2 i_332379221(.A(idata[9]), .B(cacheD[148]), .Z(cacheD[9]));
	notech_and2 i_332279222(.A(idata[10]), .B(cacheD[148]), .Z(cacheD[10])
		);
	notech_and2 i_332179223(.A(idata[11]), .B(cacheD[148]), .Z(cacheD[11])
		);
	notech_and2 i_332079224(.A(idata[12]), .B(cacheD[148]), .Z(cacheD[12])
		);
	notech_and2 i_331979225(.A(idata[13]), .B(cacheD[148]), .Z(cacheD[13])
		);
	notech_and2 i_331879226(.A(idata[14]), .B(cacheD[148]), .Z(cacheD[14])
		);
	notech_and2 i_331779227(.A(idata[15]), .B(cacheD[148]), .Z(cacheD[15])
		);
	notech_and2 i_331679228(.A(idata[16]), .B(cacheD[148]), .Z(cacheD[16])
		);
	notech_and2 i_331579229(.A(idata[17]), .B(cacheD[148]), .Z(cacheD[17])
		);
	notech_and2 i_331479230(.A(idata[18]), .B(cacheD[148]), .Z(cacheD[18])
		);
	notech_and2 i_331379231(.A(idata[19]), .B(cacheD[148]), .Z(cacheD[19])
		);
	notech_and2 i_331279232(.A(idata[20]), .B(cacheD[148]), .Z(cacheD[20])
		);
	notech_and2 i_331179233(.A(idata[21]), .B(cacheD[148]), .Z(cacheD[21])
		);
	notech_and2 i_331079234(.A(idata[22]), .B(cacheD[148]), .Z(cacheD[22])
		);
	notech_and2 i_330979235(.A(idata[23]), .B(cacheD[148]), .Z(cacheD[23])
		);
	notech_and2 i_330879236(.A(idata[24]), .B(cacheD[148]), .Z(cacheD[24])
		);
	notech_and2 i_330779237(.A(idata[25]), .B(cacheD[148]), .Z(cacheD[25])
		);
	notech_and2 i_330679238(.A(idata[26]), .B(cacheD[148]), .Z(cacheD[26])
		);
	notech_and2 i_330579239(.A(idata[27]), .B(cacheD[148]), .Z(cacheD[27])
		);
	notech_and2 i_330479240(.A(idata[28]), .B(cacheD[148]), .Z(cacheD[28])
		);
	notech_and2 i_330379241(.A(idata[29]), .B(cacheD[148]), .Z(cacheD[29])
		);
	notech_and2 i_330279242(.A(idata[30]), .B(cacheD[148]), .Z(cacheD[30])
		);
	notech_and2 i_330179243(.A(idata[31]), .B(cacheD[148]), .Z(cacheD[31])
		);
	notech_and2 i_330079244(.A(idata[32]), .B(cacheD[148]), .Z(cacheD[32])
		);
	notech_and2 i_329979245(.A(idata[33]), .B(cacheD[148]), .Z(cacheD[33])
		);
	notech_and2 i_329879246(.A(idata[34]), .B(cacheD[148]), .Z(cacheD[34])
		);
	notech_and2 i_329779247(.A(idata[35]), .B(cacheD[148]), .Z(cacheD[35])
		);
	notech_and2 i_329679248(.A(idata[36]), .B(cacheD[148]), .Z(cacheD[36])
		);
	notech_and2 i_329579249(.A(idata[37]), .B(cacheD[148]), .Z(cacheD[37])
		);
	notech_and2 i_329479250(.A(idata[38]), .B(cacheD[148]), .Z(cacheD[38])
		);
	notech_and2 i_329379251(.A(idata[39]), .B(cacheD[148]), .Z(cacheD[39])
		);
	notech_and2 i_329279252(.A(idata[40]), .B(cacheD[148]), .Z(cacheD[40])
		);
	notech_and2 i_329179253(.A(idata[41]), .B(cacheD[148]), .Z(cacheD[41])
		);
	notech_and2 i_329079254(.A(idata[42]), .B(cacheD[148]), .Z(cacheD[42])
		);
	notech_and2 i_328979255(.A(idata[43]), .B(cacheD[148]), .Z(cacheD[43])
		);
	notech_and2 i_328879256(.A(idata[44]), .B(cacheD[148]), .Z(cacheD[44])
		);
	notech_and2 i_328779257(.A(idata[45]), .B(cacheD[148]), .Z(cacheD[45])
		);
	notech_and2 i_328679258(.A(idata[46]), .B(cacheD[148]), .Z(cacheD[46])
		);
	notech_and2 i_328579259(.A(idata[47]), .B(cacheD[148]), .Z(cacheD[47])
		);
	notech_and2 i_328479260(.A(idata[48]), .B(cacheD[148]), .Z(cacheD[48])
		);
	notech_and2 i_328379261(.A(idata[49]), .B(cacheD[148]), .Z(cacheD[49])
		);
	notech_and2 i_328279262(.A(idata[50]), .B(cacheD[148]), .Z(cacheD[50])
		);
	notech_and2 i_328179263(.A(idata[51]), .B(cacheD[148]), .Z(cacheD[51])
		);
	notech_and2 i_328079264(.A(idata[52]), .B(cacheD[148]), .Z(cacheD[52])
		);
	notech_and2 i_327979265(.A(idata[53]), .B(cacheD[148]), .Z(cacheD[53])
		);
	notech_and2 i_327879266(.A(idata[54]), .B(cacheD[148]), .Z(cacheD[54])
		);
	notech_and2 i_327779267(.A(idata[55]), .B(cacheD[148]), .Z(cacheD[55])
		);
	notech_and2 i_327679268(.A(idata[56]), .B(cacheD[148]), .Z(cacheD[56])
		);
	notech_and2 i_327579269(.A(idata[57]), .B(cacheD[148]), .Z(cacheD[57])
		);
	notech_and2 i_327479270(.A(idata[58]), .B(cacheD[148]), .Z(cacheD[58])
		);
	notech_and2 i_327379271(.A(idata[59]), .B(cacheD[148]), .Z(cacheD[59])
		);
	notech_and2 i_327279272(.A(idata[60]), .B(cacheD[148]), .Z(cacheD[60])
		);
	notech_and2 i_327179273(.A(idata[61]), .B(cacheD[148]), .Z(cacheD[61])
		);
	notech_and2 i_327079274(.A(idata[62]), .B(cacheD[148]), .Z(cacheD[62])
		);
	notech_and2 i_326979275(.A(idata[63]), .B(cacheD[148]), .Z(cacheD[63])
		);
	notech_and2 i_326879276(.A(idata[64]), .B(cacheD[148]), .Z(cacheD[64])
		);
	notech_and2 i_326779277(.A(idata[65]), .B(cacheD[148]), .Z(cacheD[65])
		);
	notech_and2 i_326679278(.A(idata[66]), .B(cacheD[148]), .Z(cacheD[66])
		);
	notech_and2 i_326579279(.A(idata[67]), .B(cacheD[148]), .Z(cacheD[67])
		);
	notech_and2 i_326479280(.A(idata[68]), .B(cacheD[148]), .Z(cacheD[68])
		);
	notech_and2 i_326379281(.A(idata[69]), .B(cacheD[148]), .Z(cacheD[69])
		);
	notech_and2 i_326279282(.A(idata[70]), .B(cacheD[148]), .Z(cacheD[70])
		);
	notech_and2 i_326179283(.A(idata[71]), .B(cacheD[148]), .Z(cacheD[71])
		);
	notech_and2 i_326079284(.A(idata[72]), .B(cacheD[148]), .Z(cacheD[72])
		);
	notech_and2 i_325979285(.A(idata[73]), .B(cacheD[148]), .Z(cacheD[73])
		);
	notech_and2 i_325879286(.A(idata[74]), .B(cacheD[148]), .Z(cacheD[74])
		);
	notech_and2 i_325779287(.A(idata[75]), .B(cacheD[148]), .Z(cacheD[75])
		);
	notech_and2 i_325679288(.A(idata[76]), .B(cacheD[148]), .Z(cacheD[76])
		);
	notech_and2 i_325579289(.A(idata[77]), .B(cacheD[148]), .Z(cacheD[77])
		);
	notech_and2 i_325479290(.A(idata[78]), .B(cacheD[148]), .Z(cacheD[78])
		);
	notech_and2 i_325379291(.A(idata[79]), .B(cacheD[148]), .Z(cacheD[79])
		);
	notech_and2 i_325279292(.A(idata[80]), .B(cacheD[148]), .Z(cacheD[80])
		);
	notech_and2 i_325179293(.A(idata[81]), .B(cacheD[148]), .Z(cacheD[81])
		);
	notech_and2 i_325079294(.A(idata[82]), .B(cacheD[148]), .Z(cacheD[82])
		);
	notech_and2 i_324979295(.A(idata[83]), .B(cacheD[148]), .Z(cacheD[83])
		);
	notech_and2 i_324879296(.A(idata[84]), .B(cacheD[148]), .Z(cacheD[84])
		);
	notech_and2 i_324779297(.A(idata[85]), .B(cacheD[148]), .Z(cacheD[85])
		);
	notech_and2 i_324679298(.A(idata[86]), .B(cacheD[148]), .Z(cacheD[86])
		);
	notech_and2 i_324579299(.A(idata[87]), .B(cacheD[148]), .Z(cacheD[87])
		);
	notech_and2 i_324479300(.A(idata[88]), .B(cacheD[148]), .Z(cacheD[88])
		);
	notech_and2 i_324379301(.A(idata[89]), .B(cacheD[148]), .Z(cacheD[89])
		);
	notech_and2 i_324279302(.A(idata[90]), .B(cacheD[148]), .Z(cacheD[90])
		);
	notech_and2 i_324179303(.A(idata[91]), .B(cacheD[148]), .Z(cacheD[91])
		);
	notech_and2 i_324079304(.A(idata[92]), .B(cacheD[148]), .Z(cacheD[92])
		);
	notech_and2 i_323979305(.A(idata[93]), .B(cacheD[148]), .Z(cacheD[93])
		);
	notech_and2 i_323879306(.A(idata[94]), .B(cacheD[148]), .Z(cacheD[94])
		);
	notech_and2 i_323779307(.A(idata[95]), .B(cacheD[148]), .Z(cacheD[95])
		);
	notech_and2 i_323679308(.A(idata[96]), .B(cacheD[148]), .Z(cacheD[96])
		);
	notech_and2 i_323579309(.A(idata[97]), .B(cacheD[148]), .Z(cacheD[97])
		);
	notech_and2 i_323479310(.A(idata[98]), .B(cacheD[148]), .Z(cacheD[98])
		);
	notech_and2 i_323379311(.A(idata[99]), .B(cacheD[148]), .Z(cacheD[99])
		);
	notech_and2 i_323279312(.A(idata[100]), .B(cacheD[148]), .Z(cacheD[100])
		);
	notech_and2 i_323179313(.A(idata[101]), .B(cacheD[148]), .Z(cacheD[101])
		);
	notech_and2 i_323079314(.A(idata[102]), .B(cacheD[148]), .Z(cacheD[102])
		);
	notech_and2 i_322979315(.A(idata[103]), .B(cacheD[148]), .Z(cacheD[103])
		);
	notech_and2 i_322879316(.A(idata[104]), .B(cacheD[148]), .Z(cacheD[104])
		);
	notech_and2 i_322779317(.A(idata[105]), .B(cacheD[148]), .Z(cacheD[105])
		);
	notech_and2 i_322679318(.A(idata[106]), .B(cacheD[148]), .Z(cacheD[106])
		);
	notech_and2 i_322579319(.A(idata[107]), .B(cacheD[148]), .Z(cacheD[107])
		);
	notech_and2 i_322479320(.A(idata[108]), .B(cacheD[148]), .Z(cacheD[108])
		);
	notech_and2 i_322379321(.A(idata[109]), .B(cacheD[148]), .Z(cacheD[109])
		);
	notech_and2 i_322279322(.A(idata[110]), .B(cacheD[148]), .Z(cacheD[110])
		);
	notech_and2 i_322179323(.A(idata[111]), .B(cacheD[148]), .Z(cacheD[111])
		);
	notech_and2 i_322079324(.A(idata[112]), .B(cacheD[148]), .Z(cacheD[112])
		);
	notech_and2 i_321979325(.A(idata[113]), .B(cacheD[148]), .Z(cacheD[113])
		);
	notech_and2 i_321879326(.A(idata[114]), .B(cacheD[148]), .Z(cacheD[114])
		);
	notech_and2 i_321779327(.A(idata[115]), .B(cacheD[148]), .Z(cacheD[115])
		);
	notech_and2 i_321679328(.A(idata[116]), .B(cacheD[148]), .Z(cacheD[116])
		);
	notech_and2 i_321579329(.A(idata[117]), .B(cacheD[148]), .Z(cacheD[117])
		);
	notech_and2 i_321479330(.A(idata[118]), .B(cacheD[148]), .Z(cacheD[118])
		);
	notech_and2 i_321379331(.A(idata[119]), .B(cacheD[148]), .Z(cacheD[119])
		);
	notech_and2 i_321279332(.A(idata[120]), .B(cacheD[148]), .Z(cacheD[120])
		);
	notech_and2 i_321179333(.A(idata[121]), .B(cacheD[148]), .Z(cacheD[121])
		);
	notech_and2 i_321079334(.A(idata[122]), .B(cacheD[148]), .Z(cacheD[122])
		);
	notech_and2 i_320979335(.A(idata[123]), .B(cacheD[148]), .Z(cacheD[123])
		);
	notech_and2 i_320879336(.A(idata[124]), .B(cacheD[148]), .Z(cacheD[124])
		);
	notech_and2 i_320779337(.A(idata[125]), .B(cacheD[148]), .Z(cacheD[125])
		);
	notech_and2 i_320679338(.A(idata[126]), .B(cacheD[148]), .Z(cacheD[126])
		);
	notech_and2 i_320579339(.A(idata[127]), .B(cacheD[148]), .Z(cacheD[127])
		);
	notech_and2 i_320479340(.A(iaddr[14]), .B(cacheD[148]), .Z(cacheD[128])
		);
	notech_and2 i_320379341(.A(iaddr[15]), .B(cacheD[148]), .Z(cacheD[129])
		);
	notech_and2 i_320279342(.A(iaddr[16]), .B(cacheD[148]), .Z(cacheD[130])
		);
	notech_and2 i_320179343(.A(iaddr[17]), .B(cacheD[148]), .Z(cacheD[131])
		);
	notech_and2 i_320079344(.A(iaddr[18]), .B(cacheD[148]), .Z(cacheD[132])
		);
	notech_and2 i_319979345(.A(iaddr[19]), .B(cacheD[148]), .Z(cacheD[133])
		);
	notech_and2 i_319879346(.A(iaddr[20]), .B(cacheD[148]), .Z(cacheD[134])
		);
	notech_and2 i_319779347(.A(iaddr[21]), .B(cacheD[148]), .Z(cacheD[135])
		);
	notech_and2 i_319679348(.A(iaddr[22]), .B(cacheD[148]), .Z(cacheD[136])
		);
	notech_and2 i_319579349(.A(iaddr[23]), .B(cacheD[148]), .Z(cacheD[137])
		);
	notech_and2 i_319479350(.A(iaddr[24]), .B(cacheD[148]), .Z(cacheD[138])
		);
	notech_and2 i_319379351(.A(iaddr[25]), .B(cacheD[148]), .Z(cacheD[139])
		);
	notech_and2 i_319279352(.A(iaddr[26]), .B(cacheD[148]), .Z(cacheD[140])
		);
	notech_and2 i_319179353(.A(iaddr[27]), .B(cacheD[148]), .Z(cacheD[141])
		);
	notech_and2 i_319079354(.A(iaddr[28]), .B(cacheD[148]), .Z(cacheD[142])
		);
	notech_and2 i_318979355(.A(iaddr[29]), .B(cacheD[148]), .Z(cacheD[143])
		);
	notech_and2 i_318879356(.A(iaddr[30]), .B(cacheD[148]), .Z(cacheD[144])
		);
	notech_and2 i_318779357(.A(iaddr[31]), .B(cacheD[148]), .Z(cacheD[145])
		);
	notech_nao3 i_27978944(.A(n_29296760), .B(n_59996), .C(n_307096441), .Z(n_45696924
		));
	notech_or4 i_4079178(.A(addrshft[0]), .B(addrshft[1]), .C(addrshft[3]), 
		.D(addrshft[2]), .Z(n_46296930));
	notech_nor2 i_6279186(.A(pc_pg_fault), .B(purge_cnt[10]), .Z(n_46396931)
		);
	notech_xor2 i_3178652(.A(nbus_12105[5]), .B(nbus_12105[4]), .Z(n_46496932
		));
	notech_ao4 i_64565(.A(n_7789), .B(n_7790), .C(n_59996), .D(n_307096441),
		 .Z(\nbus_12116[0] ));
	notech_mux2 i_822067(.S(n_60400), .A(addr_0[7]), .B(pc_in[7]), .Z(n_36666
		));
	notech_mux2 i_222688(.S(n_51396981), .A(n_51196979), .B(n_51296980), .Z(n_35007
		));
	notech_ao4 i_222684(.A(n_142353056), .B(n_51496982), .C(n_8293), .D(n_42170
		), .Z(n_35037));
	notech_ao4 i_22928629(.A(n_60225), .B(n_42703), .C(n_54284), .D(n_42769)
		, .Z(n_36443));
	notech_ao4 i_22628626(.A(n_60225), .B(n_42700), .C(n_54284), .D(n_42772)
		, .Z(n_36425));
	notech_ao4 i_22428624(.A(n_60225), .B(n_42698), .C(n_54284), .D(n_42774)
		, .Z(n_36413));
	notech_ao4 i_22328623(.A(n_60225), .B(n_42697), .C(n_54284), .D(n_42775)
		, .Z(n_36407));
	notech_ao4 i_22128621(.A(n_60169), .B(n_42695), .C(n_54284), .D(n_42777)
		, .Z(n_36395));
	notech_ao4 i_22028620(.A(n_60169), .B(n_42694), .C(n_54284), .D(n_42778)
		, .Z(n_36389));
	notech_ao4 i_21928619(.A(n_60169), .B(n_42693), .C(n_54284), .D(n_42779)
		, .Z(n_36383));
	notech_ao4 i_21828618(.A(n_60169), .B(n_42692), .C(n_54284), .D(n_42780)
		, .Z(n_36377));
	notech_ao4 i_21728617(.A(n_60169), .B(n_42691), .C(n_54284), .D(n_42867)
		, .Z(n_36371));
	notech_ao4 i_21628616(.A(n_60169), .B(n_42690), .C(n_54284), .D(n_42781)
		, .Z(n_36365));
	notech_nor2 i_3778715(.A(n_140853041), .B(n_60243), .Z(n_49596963));
	notech_ao4 i_14928549(.A(n_60169), .B(n_42623), .C(n_54284), .D(n_42845)
		, .Z(n_35963));
	notech_or4 i_173276959(.A(n_61549), .B(n_60277), .C(n_60245), .D(n_42866
		), .Z(n_49796965));
	notech_nand2 i_12828528(.A(n_51596983), .B(n_49796965), .Z(n_35837));
	notech_or4 i_174076951(.A(n_61549), .B(n_60277), .C(n_60245), .D(n_42865
		), .Z(n_50096968));
	notech_nand2 i_12628526(.A(n_51696984), .B(n_50096968), .Z(n_35825));
	notech_or4 i_189676795(.A(n_61549), .B(n_60277), .C(n_60245), .D(n_42867
		), .Z(n_50396971));
	notech_nand2 i_8928489(.A(n_51796985), .B(n_50396971), .Z(n_35603));
	notech_or4 i_197076721(.A(n_61549), .B(n_60277), .C(n_60245), .D(n_42864
		), .Z(n_50596973));
	notech_nand2 i_7128471(.A(n_51896986), .B(n_50596973), .Z(n_35495));
	notech_or4 i_201876673(.A(n_61549), .B(n_60274), .C(n_60243), .D(n_42863
		), .Z(n_50796975));
	notech_nand2 i_5928459(.A(n_51996987), .B(n_50796975), .Z(n_35423));
	notech_and2 i_2378660(.A(n_60243), .B(n_42741), .Z(n_51196979));
	notech_and2 i_2678657(.A(n_59996), .B(n_42741), .Z(n_51296980));
	notech_xor2 i_2178662(.A(wptr[0]), .B(n_60274), .Z(n_51396981));
	notech_nand2 i_169177000(.A(fault_wptr[1]), .B(fault_wptr[0]), .Z(n_51496982
		));
	notech_ao4 i_173476957(.A(n_59996), .B(n_42545), .C(n_60169), .D(n_42730
		), .Z(n_51596983));
	notech_ao4 i_174276949(.A(n_59996), .B(n_42541), .C(n_60165), .D(n_42728
		), .Z(n_51696984));
	notech_ao4 i_189976792(.A(n_59996), .B(n_42467), .C(n_60165), .D(n_42691
		), .Z(n_51796985));
	notech_ao4 i_197276719(.A(n_60165), .B(n_42673), .C(n_59996), .D(n_42431
		), .Z(n_51896986));
	notech_ao4 i_202076671(.A(n_60165), .B(n_42661), .C(n_59996), .D(n_42407
		), .Z(n_51996987));
	notech_nao3 i_64520(.A(n_32555629), .B(n_8293), .C(n_42167), .Z(n_35014)
		);
	notech_nand3 i_65536(.A(n_32555629), .B(n_45696924), .C(n_306996440), .Z
		(\nbus_12119[0] ));
	notech_nand3 i_64530(.A(n_8293), .B(n_32555629), .C(n_29196759), .Z(\nbus_12115[0] 
		));
	notech_ao4 i_64539(.A(n_101094414), .B(n_42741), .C(n_42168), .D(n_309596466
		), .Z(n_35044));
	notech_or2 i_65491(.A(pc_pg_fault), .B(purge), .Z(\nbus_12118[0] ));
	notech_or2 i_65557(.A(pc_pg_fault), .B(n_28996757), .Z(n_36952));
	notech_ao4 i_64566(.A(n_7789), .B(n_52196989), .C(n_59996), .D(n_307096441
		), .Z(\nbus_12116[128] ));
	notech_mux2 i_179460(.S(purge), .A(iaddr[4]), .B(purge_cnt[0]), .Z(cacheA
		[0]));
	notech_mux2 i_211494(.S(purge), .A(iaddr[5]), .B(purge_cnt[1]), .Z(cacheA
		[1]));
	notech_mux2 i_379459(.S(purge), .A(iaddr[6]), .B(purge_cnt[2]), .Z(cacheA
		[2]));
	notech_mux2 i_479458(.S(purge), .A(iaddr[7]), .B(purge_cnt[3]), .Z(cacheA
		[3]));
	notech_mux2 i_511495(.S(purge), .A(iaddr[8]), .B(purge_cnt[4]), .Z(cacheA
		[4]));
	notech_mux2 i_679457(.S(purge), .A(iaddr[9]), .B(purge_cnt[5]), .Z(cacheA
		[5]));
	notech_mux2 i_779456(.S(purge), .A(iaddr[10]), .B(purge_cnt[6]), .Z(cacheA
		[6]));
	notech_mux2 i_879455(.S(purge), .A(iaddr[11]), .B(purge_cnt[7]), .Z(cacheA
		[7]));
	notech_mux2 i_979454(.S(purge), .A(iaddr[12]), .B(purge_cnt[8]), .Z(cacheA
		[8]));
	notech_mux2 i_1079453(.S(purge), .A(iaddr[13]), .B(purge_cnt[9]), .Z(cacheA
		[9]));
	notech_mux2 i_127171(.S(addrshft[0]), .A(n_3392), .B(n_112493391), .Z(valid_len_097049
		));
	notech_ao4 i_527175(.A(addrshft[4]), .B(n_3392), .C(n_26296730), .D(n_112493391
		), .Z(valid_len_497048));
	notech_mux2 i_3279209(.S(n_60400), .A(addr_0[31]), .B(pc_in[31]), .Z(n_36810
		));
	notech_mux2 i_3179208(.S(n_60400), .A(addr_0[30]), .B(pc_in[30]), .Z(n_36804
		));
	notech_mux2 i_3079207(.S(n_60400), .A(addr_0[29]), .B(pc_in[29]), .Z(n_36798
		));
	notech_mux2 i_2979206(.S(n_60400), .A(addr_0[28]), .B(pc_in[28]), .Z(n_36792
		));
	notech_mux2 i_2879205(.S(n_60400), .A(addr_0[27]), .B(pc_in[27]), .Z(n_36786
		));
	notech_mux2 i_2779204(.S(n_60400), .A(addr_0[26]), .B(pc_in[26]), .Z(n_36780
		));
	notech_mux2 i_2679203(.S(n_60400), .A(addr_0[25]), .B(pc_in[25]), .Z(n_36774
		));
	notech_mux2 i_2579202(.S(n_60400), .A(addr_0[24]), .B(pc_in[24]), .Z(n_36768
		));
	notech_mux2 i_2479201(.S(n_60400), .A(addr_0[23]), .B(pc_in[23]), .Z(n_36762
		));
	notech_mux2 i_2379200(.S(n_60400), .A(addr_0[22]), .B(pc_in[22]), .Z(n_36756
		));
	notech_mux2 i_2279199(.S(n_60400), .A(addr_0[21]), .B(pc_in[21]), .Z(n_36750
		));
	notech_mux2 i_2179198(.S(n_60400), .A(addr_0[20]), .B(pc_in[20]), .Z(n_36744
		));
	notech_mux2 i_2079197(.S(n_60400), .A(addr_0[19]), .B(pc_in[19]), .Z(n_36738
		));
	notech_mux2 i_1979196(.S(n_60400), .A(addr_0[18]), .B(pc_in[18]), .Z(n_36732
		));
	notech_mux2 i_1879195(.S(n_60396), .A(addr_0[17]), .B(pc_in[17]), .Z(n_36726
		));
	notech_mux2 i_1779194(.S(n_60396), .A(addr_0[16]), .B(pc_in[16]), .Z(n_36720
		));
	notech_mux2 i_1679193(.S(n_60396), .A(addr_0[15]), .B(pc_in[15]), .Z(n_36714
		));
	notech_mux2 i_1579192(.S(n_60396), .A(addr_0[14]), .B(pc_in[14]), .Z(n_36708
		));
	notech_mux2 i_1479191(.S(n_60396), .A(addr_0[13]), .B(pc_in[13]), .Z(n_36702
		));
	notech_mux2 i_1379190(.S(n_60396), .A(addr_0[12]), .B(pc_in[12]), .Z(n_36696
		));
	notech_mux2 i_1279189(.S(n_60396), .A(addr_0[11]), .B(pc_in[11]), .Z(n_36690
		));
	notech_mux2 i_1179188(.S(n_60396), .A(addr_0[10]), .B(pc_in[10]), .Z(n_36684
		));
	notech_mux2 i_1022069(.S(n_60396), .A(addr_0[9]), .B(pc_in[9]), .Z(n_36678
		));
	notech_mux2 i_922068(.S(n_60396), .A(addr_0[8]), .B(pc_in[8]), .Z(n_36672
		));
	notech_mux2 i_722066(.S(n_60396), .A(addr_0[6]), .B(pc_in[6]), .Z(n_36660
		));
	notech_mux2 i_622065(.S(n_60396), .A(addr_0[5]), .B(pc_in[5]), .Z(n_36654
		));
	notech_mux2 i_522064(.S(n_60396), .A(addr_0[4]), .B(pc_in[4]), .Z(n_36648
		));
	notech_mux2 i_427186(.S(n_60396), .A(nbus_12105[3]), .B(pc_in[3]), .Z(n_36931
		));
	notech_mux2 i_327185(.S(n_60396), .A(nbus_12105[2]), .B(pc_in[2]), .Z(n_36925
		));
	notech_mux2 i_227184(.S(n_60396), .A(nbus_12105[1]), .B(pc_in[1]), .Z(n_36919
		));
	notech_mux2 i_127183(.S(n_60396), .A(nbus_12105[0]), .B(pc_in[0]), .Z(n_36913
		));
	notech_ao4 i_122683(.A(n_142353056), .B(fault_wptr[0]), .C(n_8293), .D(n_42169
		), .Z(n_35031));
	notech_ao4 i_25628656(.A(n_60169), .B(n_42730), .C(n_54284), .D(n_42866)
		, .Z(n_36605));
	notech_ao4 i_25528655(.A(n_54284), .B(n_42744), .C(n_60169), .D(n_42729)
		, .Z(n_36599));
	notech_ao4 i_25428654(.A(n_60165), .B(n_42728), .C(n_54284), .D(n_42865)
		, .Z(n_36593));
	notech_ao4 i_25328653(.A(n_54284), .B(n_42745), .C(n_60169), .D(n_42727)
		, .Z(n_36587));
	notech_ao4 i_25228652(.A(n_54284), .B(n_42746), .C(n_60174), .D(n_42726)
		, .Z(n_36581));
	notech_ao4 i_25128651(.A(n_54282), .B(n_42747), .C(n_60174), .D(n_42725)
		, .Z(n_36575));
	notech_ao4 i_25028650(.A(n_54282), .B(n_42748), .C(n_60174), .D(n_42724)
		, .Z(n_36569));
	notech_ao4 i_24928649(.A(n_54282), .B(n_42749), .C(n_60174), .D(n_42723)
		, .Z(n_36563));
	notech_ao4 i_24828648(.A(n_54282), .B(n_42750), .C(n_60174), .D(n_42722)
		, .Z(n_36557));
	notech_ao4 i_24728647(.A(n_54282), .B(n_42751), .C(n_60174), .D(n_42721)
		, .Z(n_36551));
	notech_ao4 i_24628646(.A(n_54282), .B(n_42752), .C(n_60174), .D(n_42720)
		, .Z(n_36545));
	notech_ao4 i_24528645(.A(n_60174), .B(n_42719), .C(n_54282), .D(n_42753)
		, .Z(n_36539));
	notech_ao4 i_24428644(.A(n_54282), .B(n_42754), .C(n_60174), .D(n_42718)
		, .Z(n_36533));
	notech_ao4 i_24328643(.A(n_54282), .B(n_42755), .C(n_60174), .D(n_42717)
		, .Z(n_36527));
	notech_ao4 i_24228642(.A(n_54282), .B(n_42756), .C(n_60169), .D(n_42716)
		, .Z(n_36521));
	notech_ao4 i_24128641(.A(n_54282), .B(n_42757), .C(n_60169), .D(n_42715)
		, .Z(n_36515));
	notech_ao4 i_24028640(.A(n_54282), .B(n_42758), .C(n_60174), .D(n_42714)
		, .Z(n_36509));
	notech_ao4 i_23928639(.A(n_54282), .B(n_42759), .C(n_60174), .D(n_42713)
		, .Z(n_36503));
	notech_ao4 i_23828638(.A(n_54282), .B(n_42760), .C(n_60174), .D(n_42712)
		, .Z(n_36497));
	notech_ao4 i_23728637(.A(n_54282), .B(n_42761), .C(n_60174), .D(n_42711)
		, .Z(n_36491));
	notech_ao4 i_23628636(.A(n_54282), .B(n_42762), .C(n_60156), .D(n_42710)
		, .Z(n_36485));
	notech_ao4 i_23528635(.A(n_54289), .B(n_42763), .C(n_60156), .D(n_42709)
		, .Z(n_36479));
	notech_ao4 i_23428634(.A(n_54289), .B(n_42764), .C(n_60156), .D(n_42708)
		, .Z(n_36473));
	notech_ao4 i_23328633(.A(n_54289), .B(n_42765), .C(n_60156), .D(n_42707)
		, .Z(n_36467));
	notech_ao4 i_23228632(.A(n_54289), .B(n_42766), .C(n_60160), .D(n_42706)
		, .Z(n_36461));
	notech_ao4 i_23128631(.A(n_60160), .B(n_42705), .C(n_54289), .D(n_42767)
		, .Z(n_36455));
	notech_ao4 i_23028630(.A(n_60156), .B(n_42704), .C(n_54289), .D(n_42768)
		, .Z(n_36449));
	notech_ao4 i_22828628(.A(n_60160), .B(n_42702), .C(n_54289), .D(n_42770)
		, .Z(n_36437));
	notech_ao4 i_22728627(.A(n_60156), .B(n_42701), .C(n_54289), .D(n_42771)
		, .Z(n_36431));
	notech_ao4 i_22528625(.A(n_60156), .B(n_42699), .C(n_54289), .D(n_42773)
		, .Z(n_36419));
	notech_ao4 i_22228622(.A(n_60156), .B(n_42696), .C(n_54289), .D(n_42776)
		, .Z(n_36401));
	notech_ao4 i_21528615(.A(n_60156), .B(n_42689), .C(n_54289), .D(n_42782)
		, .Z(n_36359));
	notech_ao4 i_21428614(.A(n_60156), .B(n_42688), .C(n_54289), .D(n_42783)
		, .Z(n_36353));
	notech_ao4 i_21328613(.A(n_60156), .B(n_42687), .C(n_54289), .D(n_42784)
		, .Z(n_36347));
	notech_ao4 i_21228612(.A(n_60156), .B(n_42686), .C(n_54289), .D(n_42785)
		, .Z(n_36341));
	notech_ao4 i_21128611(.A(n_60156), .B(n_42685), .C(n_54289), .D(n_42786)
		, .Z(n_36335));
	notech_ao4 i_21028610(.A(n_60165), .B(n_42684), .C(n_54289), .D(n_42787)
		, .Z(n_36329));
	notech_ao4 i_20928609(.A(n_60165), .B(n_42683), .C(n_54287), .D(n_42788)
		, .Z(n_36323));
	notech_ao4 i_20828608(.A(n_60160), .B(n_42682), .C(n_54287), .D(n_42789)
		, .Z(n_36317));
	notech_ao4 i_20728607(.A(n_60165), .B(n_42681), .C(n_54287), .D(n_42790)
		, .Z(n_36311));
	notech_ao4 i_20628606(.A(n_60165), .B(n_42680), .C(n_54287), .D(n_42791)
		, .Z(n_36305));
	notech_ao4 i_20528605(.A(n_60165), .B(n_42679), .C(n_54287), .D(n_42792)
		, .Z(n_36299));
	notech_ao4 i_20428604(.A(n_60165), .B(n_42678), .C(n_54287), .D(n_42793)
		, .Z(n_36293));
	notech_ao4 i_20328603(.A(n_60165), .B(n_42677), .C(n_54287), .D(n_42794)
		, .Z(n_36287));
	notech_ao4 i_20228602(.A(n_60160), .B(n_42676), .C(n_54287), .D(n_42795)
		, .Z(n_36281));
	notech_ao4 i_20128601(.A(n_60160), .B(n_42675), .C(n_54287), .D(n_42796)
		, .Z(n_36275));
	notech_ao4 i_20028600(.A(n_60160), .B(n_42674), .C(n_54287), .D(n_42797)
		, .Z(n_36269));
	notech_ao4 i_19928599(.A(n_60160), .B(n_42673), .C(n_54287), .D(n_42864)
		, .Z(n_36263));
	notech_ao4 i_19828598(.A(n_60160), .B(n_42672), .C(n_54287), .D(n_42798)
		, .Z(n_36257));
	notech_ao4 i_19728597(.A(n_60160), .B(n_42671), .C(n_54287), .D(n_42799)
		, .Z(n_36251));
	notech_ao4 i_19628596(.A(n_60160), .B(n_42670), .C(n_54287), .D(n_42800)
		, .Z(n_36245));
	notech_ao4 i_19528595(.A(n_60160), .B(n_42669), .C(n_54287), .D(n_42801)
		, .Z(n_36239));
	notech_ao4 i_19428594(.A(n_60174), .B(n_42668), .C(n_54287), .D(n_42802)
		, .Z(n_36233));
	notech_ao4 i_19328593(.A(n_60188), .B(n_42667), .C(n_54274), .D(n_42803)
		, .Z(n_36227));
	notech_ao4 i_19228592(.A(n_60193), .B(n_42666), .C(n_54274), .D(n_42804)
		, .Z(n_36221));
	notech_ao4 i_19128591(.A(n_60188), .B(n_42665), .C(n_54274), .D(n_42805)
		, .Z(n_36215));
	notech_ao4 i_19028590(.A(n_60188), .B(n_42664), .C(n_54274), .D(n_42806)
		, .Z(n_36209));
	notech_ao4 i_18928589(.A(n_60193), .B(n_42663), .C(n_54274), .D(n_42807)
		, .Z(n_36203));
	notech_ao4 i_18828588(.A(n_60193), .B(n_42662), .C(n_54274), .D(n_42808)
		, .Z(n_36197));
	notech_ao4 i_18728587(.A(n_60193), .B(n_42661), .C(n_54274), .D(n_42863)
		, .Z(n_36191));
	notech_ao4 i_18628586(.A(n_60193), .B(n_42660), .C(n_54274), .D(n_42809)
		, .Z(n_36185));
	notech_ao4 i_18528585(.A(n_60188), .B(n_42659), .C(n_54274), .D(n_42810)
		, .Z(n_36179));
	notech_ao4 i_18428584(.A(n_60188), .B(n_42658), .C(n_54274), .D(n_42811)
		, .Z(n_36173));
	notech_ao4 i_18328583(.A(n_54274), .B(n_42812), .C(n_60188), .D(n_42657)
		, .Z(n_36167));
	notech_ao4 i_18228582(.A(n_60188), .B(n_42656), .C(n_54274), .D(n_42813)
		, .Z(n_36161));
	notech_ao4 i_18128581(.A(n_60188), .B(n_42655), .C(n_54274), .D(n_42814)
		, .Z(n_36155));
	notech_ao4 i_18028580(.A(n_60188), .B(n_42654), .C(n_54274), .D(n_42815)
		, .Z(n_36149));
	notech_ao4 i_17928579(.A(n_60188), .B(n_42653), .C(n_54274), .D(n_42816)
		, .Z(n_36143));
	notech_ao4 i_17828578(.A(n_60188), .B(n_42652), .C(n_54274), .D(n_42817)
		, .Z(n_36137));
	notech_ao4 i_17728577(.A(n_60197), .B(n_42651), .C(n_54272), .D(n_42818)
		, .Z(n_36131));
	notech_ao4 i_17628576(.A(n_60197), .B(n_42650), .C(n_54272), .D(n_42819)
		, .Z(n_36125));
	notech_ao4 i_17528575(.A(n_60193), .B(n_42649), .C(n_54272), .D(n_42820)
		, .Z(n_36119));
	notech_ao4 i_17428574(.A(n_60193), .B(n_42648), .C(n_54272), .D(n_42821)
		, .Z(n_36113));
	notech_ao4 i_17328573(.A(n_60197), .B(n_42647), .C(n_54272), .D(n_42822)
		, .Z(n_36107));
	notech_ao4 i_17228572(.A(n_60197), .B(n_42646), .C(n_54272), .D(n_42823)
		, .Z(n_36101));
	notech_ao4 i_17128571(.A(n_60197), .B(n_42645), .C(n_54272), .D(n_42824)
		, .Z(n_36095));
	notech_ao4 i_17028570(.A(n_60197), .B(n_42644), .C(n_54272), .D(n_42825)
		, .Z(n_36089));
	notech_ao4 i_16928569(.A(n_60193), .B(n_42643), .C(n_54272), .D(n_42826)
		, .Z(n_36083));
	notech_ao4 i_16828568(.A(n_60193), .B(n_42642), .C(n_54272), .D(n_42827)
		, .Z(n_36077));
	notech_ao4 i_16728567(.A(n_60193), .B(n_42641), .C(n_54272), .D(n_42828)
		, .Z(n_36071));
	notech_ao4 i_16628566(.A(n_60193), .B(n_42640), .C(n_54272), .D(n_42829)
		, .Z(n_36065));
	notech_ao4 i_16528565(.A(n_60193), .B(n_42639), .C(n_54272), .D(n_42830)
		, .Z(n_36059));
	notech_ao4 i_16428564(.A(n_60193), .B(n_42638), .C(n_54272), .D(n_42831)
		, .Z(n_36053));
	notech_ao4 i_16328563(.A(n_60193), .B(n_42637), .C(n_54272), .D(n_42832)
		, .Z(n_36047));
	notech_ao4 i_16228562(.A(n_60193), .B(n_42636), .C(n_54272), .D(n_42833)
		, .Z(n_36041));
	notech_ao4 i_16128561(.A(n_60154), .B(n_42635), .C(n_54279), .D(n_42834)
		, .Z(n_36035));
	notech_ao4 i_16028560(.A(n_60154), .B(n_42634), .C(n_54279), .D(n_42835)
		, .Z(n_36029));
	notech_ao4 i_15928559(.A(n_60154), .B(n_42633), .C(n_54279), .D(n_42836)
		, .Z(n_36023));
	notech_ao4 i_15828558(.A(n_60154), .B(n_42632), .C(n_54279), .D(n_42837)
		, .Z(n_36017));
	notech_ao4 i_15728557(.A(n_60184), .B(n_42631), .C(n_54279), .D(n_42838)
		, .Z(n_36011));
	notech_ao4 i_15628556(.A(n_60184), .B(n_42630), .C(n_54279), .D(n_42839)
		, .Z(n_36005));
	notech_ao4 i_15528555(.A(n_60154), .B(n_42629), .C(n_54279), .D(n_42736)
		, .Z(n_35999));
	notech_ao4 i_15428554(.A(n_60184), .B(n_42628), .C(n_54279), .D(n_42840)
		, .Z(n_35993));
	notech_ao4 i_15328553(.A(n_60154), .B(n_42627), .C(n_54279), .D(n_42841)
		, .Z(n_35987));
	notech_ao4 i_15228552(.A(n_60154), .B(n_42626), .C(n_54279), .D(n_42842)
		, .Z(n_35981));
	notech_ao4 i_15128551(.A(n_60154), .B(n_42625), .C(n_54279), .D(n_42843)
		, .Z(n_35975));
	notech_ao4 i_15028550(.A(n_60154), .B(n_42624), .C(n_54279), .D(n_42844)
		, .Z(n_35969));
	notech_ao4 i_14828548(.A(n_60154), .B(n_42622), .C(n_54279), .D(n_42846)
		, .Z(n_35957));
	notech_ao4 i_14728547(.A(n_60154), .B(n_42621), .C(n_54279), .D(n_42737)
		, .Z(n_35951));
	notech_ao4 i_14628546(.A(n_60154), .B(n_42620), .C(n_54279), .D(n_42847)
		, .Z(n_35945));
	notech_ao4 i_14528545(.A(n_60154), .B(n_42619), .C(n_54279), .D(n_42848)
		, .Z(n_35939));
	notech_ao4 i_14428544(.A(n_60184), .B(n_42618), .C(n_54277), .D(n_42849)
		, .Z(n_35933));
	notech_ao4 i_14328543(.A(n_60184), .B(n_42617), .C(n_54277), .D(n_42850)
		, .Z(n_35927));
	notech_ao4 i_14228542(.A(n_60184), .B(n_42616), .C(n_54277), .D(n_42851)
		, .Z(n_35921));
	notech_ao4 i_14128541(.A(n_60184), .B(n_42615), .C(n_54277), .D(n_42852)
		, .Z(n_35915));
	notech_ao4 i_14028540(.A(n_60188), .B(n_42614), .C(n_54277), .D(n_42853)
		, .Z(n_35909));
	notech_ao4 i_13928539(.A(n_60188), .B(n_42613), .C(n_54277), .D(n_42738)
		, .Z(n_35903));
	notech_ao4 i_13828538(.A(n_54277), .B(n_42854), .C(n_60188), .D(n_42612)
		, .Z(n_35897));
	notech_ao4 i_13728537(.A(n_60188), .B(n_42611), .C(n_54277), .D(n_42855)
		, .Z(n_35891));
	notech_ao4 i_13628536(.A(n_60184), .B(n_42610), .C(n_54277), .D(n_42856)
		, .Z(n_35885));
	notech_ao4 i_13528535(.A(n_60184), .B(n_42609), .C(n_54277), .D(n_42857)
		, .Z(n_35879));
	notech_ao4 i_13428534(.A(n_60184), .B(n_42608), .C(n_54277), .D(n_42858)
		, .Z(n_35873));
	notech_ao4 i_13328533(.A(n_60184), .B(n_42607), .C(n_54277), .D(n_42859)
		, .Z(n_35867));
	notech_ao4 i_13228532(.A(n_60184), .B(n_42606), .C(n_54277), .D(n_42860)
		, .Z(n_35861));
	notech_ao4 i_13128531(.A(n_60184), .B(n_42605), .C(n_54277), .D(n_42739)
		, .Z(n_35855));
	notech_ao4 i_13028530(.A(n_60184), .B(n_42604), .C(n_54277), .D(n_42861)
		, .Z(n_35849));
	notech_ao4 i_12928529(.A(n_60184), .B(n_42603), .C(n_54277), .D(n_42862)
		, .Z(n_35843));
	notech_nand3 i_86377828(.A(n_3078), .B(n_58379), .C(queue[36]), .Z(n_1570
		));
	notech_and4 i_2825007(.A(n_2350), .B(n_2349), .C(n_2344), .D(n_2348), .Z
		(squeue_2797078));
	notech_nand3 i_84577846(.A(n_57937), .B(n_58209), .C(queue[27]), .Z(n_1567
		));
	notech_nand3 i_83277859(.A(n_3078), .B(n_58375), .C(queue[35]), .Z(n_1554
		));
	notech_and4 i_2725006(.A(n_2336), .B(n_2335), .C(n_2330), .D(n_2334), .Z
		(squeue_2697079));
	notech_nand3 i_81477877(.A(n_57937), .B(n_58211), .C(queue[26]), .Z(n_1551
		));
	notech_nand3 i_80177890(.A(n_60258), .B(n_58375), .C(queue[34]), .Z(n_1538
		));
	notech_and4 i_2625005(.A(n_2322), .B(n_2321), .C(n_2316), .D(n_2320), .Z
		(squeue_2597080));
	notech_nand3 i_78377908(.A(n_57937), .B(n_58211), .C(queue[25]), .Z(n_1535
		));
	notech_nand3 i_77077921(.A(n_60258), .B(n_58375), .C(queue[33]), .Z(n_1522
		));
	notech_and4 i_2525004(.A(n_2308), .B(n_2307), .C(n_2302), .D(n_2306), .Z
		(squeue_2497081));
	notech_nand3 i_75277939(.A(n_57937), .B(n_58211), .C(queue[24]), .Z(n_1519
		));
	notech_nand3 i_73977952(.A(n_60258), .B(n_58379), .C(queue[32]), .Z(n_1506
		));
	notech_and4 i_2425003(.A(n_2294), .B(n_2293), .C(n_2288), .D(n_2292), .Z
		(squeue_2397082));
	notech_nand3 i_72177970(.A(n_57937), .B(n_58211), .C(queue[23]), .Z(n_1503
		));
	notech_or2 i_70877983(.A(n_58266), .B(n_42192), .Z(n_1490));
	notech_and4 i_2325002(.A(n_2280), .B(n_2279), .C(n_2274), .D(n_2278), .Z
		(squeue_2297083));
	notech_nand3 i_69078001(.A(n_57937), .B(n_58209), .C(queue[22]), .Z(n_1487
		));
	notech_nand3 i_67778014(.A(n_60262), .B(n_58375), .C(queue[30]), .Z(n_1474
		));
	notech_and4 i_2225001(.A(n_2266), .B(n_2265), .C(n_2260), .D(n_2264), .Z
		(squeue_2197084));
	notech_nand3 i_65978032(.A(n_57937), .B(n_58209), .C(queue[21]), .Z(n_1471
		));
	notech_nand3 i_64678045(.A(n_60262), .B(n_58375), .C(queue[29]), .Z(n_1458
		));
	notech_and4 i_2125000(.A(n_2252), .B(n_2251), .C(n_2246), .D(n_2250), .Z
		(squeue_2097085));
	notech_nand3 i_62878063(.A(n_57937), .B(n_58211), .C(queue[20]), .Z(n_1455
		));
	notech_nand3 i_61578076(.A(n_60258), .B(n_58375), .C(queue[28]), .Z(n_1442
		));
	notech_and4 i_2024999(.A(n_2238), .B(n_2237), .C(n_2232), .D(n_2236), .Z
		(squeue_1997086));
	notech_nand3 i_59778094(.A(n_57937), .B(n_58209), .C(queue[19]), .Z(n_1439
		));
	notech_nand3 i_58478107(.A(n_60258), .B(n_58375), .C(queue[27]), .Z(n_1426
		));
	notech_and4 i_1924998(.A(n_2224), .B(n_2223), .C(n_2218), .D(n_2222), .Z
		(squeue_1897087));
	notech_nand3 i_56678125(.A(n_57937), .B(n_58209), .C(queue[18]), .Z(n_1423
		));
	notech_nand2 i_8078716(.A(wptr[0]), .B(n_42170), .Z(n_52196989));
	notech_ao3 i_627188(.A(n_60245), .B(n_42741), .C(n_46496932), .Z(n_52296990
		));
	notech_ao3 i_5033(.A(n_42170), .B(n_42743), .C(n_142353056), .Z(n_52396991
		));
	notech_reg fault_wptr_en_reg(.CP(n_62087), .D(n_40221), .CD(n_60986), .Q
		(fault_wptr_en));
	notech_mux2 i_53164(.S(n_35014), .A(fault_wptr_en), .B(n_42168), .Z(n_40221
		));
	notech_reg addr_reg_0(.CP(n_62087), .D(n_40227), .CD(n_60986), .Q(iaddr[
		0]));
	notech_mux2 i_53172(.S(\nbus_12117[0] ), .A(iaddr[0]), .B(n_30596773), .Z
		(n_40227));
	notech_reg addr_reg_1(.CP(n_62087), .D(n_40233), .CD(n_60986), .Q(iaddr[
		1]));
	notech_mux2 i_53180(.S(\nbus_12117[0] ), .A(iaddr[1]), .B(n_30696774), .Z
		(n_40233));
	notech_reg addr_reg_2(.CP(n_62087), .D(n_40239), .CD(n_60986), .Q(iaddr[
		2]));
	notech_mux2 i_53188(.S(\nbus_12117[0] ), .A(iaddr[2]), .B(n_30796775), .Z
		(n_40239));
	notech_reg addr_reg_3(.CP(n_62087), .D(n_40245), .CD(n_60986), .Q(iaddr[
		3]));
	notech_mux2 i_53196(.S(\nbus_12117[0] ), .A(iaddr[3]), .B(n_30896776), .Z
		(n_40245));
	notech_reg addr_reg_4(.CP(n_62087), .D(n_40251), .CD(n_60987), .Q(iaddr[
		4]));
	notech_mux2 i_53204(.S(\nbus_12117[0] ), .A(iaddr[4]), .B(n_36648), .Z(n_40251
		));
	notech_reg addr_reg_5(.CP(n_62087), .D(n_40257), .CD(n_60987), .Q(iaddr[
		5]));
	notech_mux2 i_53212(.S(\nbus_12117[0] ), .A(iaddr[5]), .B(n_36654), .Z(n_40257
		));
	notech_reg addr_reg_6(.CP(n_62087), .D(n_40263), .CD(n_60987), .Q(iaddr[
		6]));
	notech_mux2 i_53220(.S(\nbus_12117[0] ), .A(iaddr[6]), .B(n_36660), .Z(n_40263
		));
	notech_reg addr_reg_7(.CP(n_62087), .D(n_40269), .CD(n_60986), .Q(iaddr[
		7]));
	notech_mux2 i_53228(.S(\nbus_12117[0] ), .A(iaddr[7]), .B(n_36666), .Z(n_40269
		));
	notech_reg addr_reg_8(.CP(n_62087), .D(n_40275), .CD(n_60987), .Q(iaddr[
		8]));
	notech_mux2 i_53236(.S(\nbus_12117[0] ), .A(iaddr[8]), .B(n_36672), .Z(n_40275
		));
	notech_nand3 i_55378138(.A(n_60258), .B(n_58375), .C(queue[26]), .Z(n_1410
		));
	notech_reg addr_reg_9(.CP(n_62087), .D(n_40281), .CD(n_60986), .Q(iaddr[
		9]));
	notech_mux2 i_53244(.S(\nbus_12117[0] ), .A(iaddr[9]), .B(n_36678), .Z(n_40281
		));
	notech_reg_set addr_reg_10(.CP(n_62181), .D(n_40287), .SD(n_60986), .Q(iaddr
		[10]));
	notech_mux2 i_53252(.S(\nbus_12117[0] ), .A(iaddr[10]), .B(n_36684), .Z(n_40287
		));
	notech_reg_set addr_reg_11(.CP(n_62181), .D(n_40293), .SD(n_60986), .Q(iaddr
		[11]));
	notech_mux2 i_53260(.S(\nbus_12117[0] ), .A(iaddr[11]), .B(n_36690), .Z(n_40293
		));
	notech_and4 i_1824997(.A(n_2210), .B(n_2209), .C(n_2204), .D(n_2208), .Z
		(squeue_1797088));
	notech_reg_set addr_reg_12(.CP(n_62181), .D(n_40299), .SD(n_60985), .Q(iaddr
		[12]));
	notech_mux2 i_53268(.S(\nbus_12117[0] ), .A(iaddr[12]), .B(n_36696), .Z(n_40299
		));
	notech_nand3 i_53578156(.A(n_57935), .B(n_58206), .C(queue[17]), .Z(n_1407
		));
	notech_reg_set addr_reg_13(.CP(n_62181), .D(n_40305), .SD(n_60985), .Q(iaddr
		[13]));
	notech_mux2 i_53276(.S(\nbus_12117[0] ), .A(iaddr[13]), .B(n_36702), .Z(n_40305
		));
	notech_reg_set addr_reg_14(.CP(n_62181), .D(n_40311), .SD(n_60985), .Q(iaddr
		[14]));
	notech_mux2 i_53284(.S(\nbus_12117[0] ), .A(iaddr[14]), .B(n_36708), .Z(n_40311
		));
	notech_reg_set addr_reg_15(.CP(n_62181), .D(n_40317), .SD(n_60986), .Q(iaddr
		[15]));
	notech_mux2 i_53292(.S(\nbus_12117[0] ), .A(iaddr[15]), .B(n_36714), .Z(n_40317
		));
	notech_reg_set addr_reg_16(.CP(n_62181), .D(n_40323), .SD(n_60986), .Q(iaddr
		[16]));
	notech_mux2 i_53300(.S(n_60143), .A(iaddr[16]), .B(n_36720), .Z(n_40323)
		);
	notech_reg_set addr_reg_17(.CP(n_62181), .D(n_40329), .SD(n_60986), .Q(iaddr
		[17]));
	notech_mux2 i_53308(.S(n_60143), .A(iaddr[17]), .B(n_36726), .Z(n_40329)
		);
	notech_reg_set addr_reg_18(.CP(n_62181), .D(n_40335), .SD(n_60986), .Q(iaddr
		[18]));
	notech_mux2 i_53316(.S(n_60143), .A(iaddr[18]), .B(n_36732), .Z(n_40335)
		);
	notech_reg_set addr_reg_19(.CP(n_62181), .D(n_40341), .SD(n_60986), .Q(iaddr
		[19]));
	notech_mux2 i_53324(.S(n_60143), .A(iaddr[19]), .B(n_36738), .Z(n_40341)
		);
	notech_reg addr_reg_20(.CP(n_62181), .D(n_40347), .CD(n_60987), .Q(iaddr
		[20]));
	notech_mux2 i_53332(.S(n_60143), .A(iaddr[20]), .B(n_36744), .Z(n_40347)
		);
	notech_reg addr_reg_21(.CP(n_62181), .D(n_40353), .CD(n_60988), .Q(iaddr
		[21]));
	notech_mux2 i_53340(.S(n_60143), .A(iaddr[21]), .B(n_36750), .Z(n_40353)
		);
	notech_reg addr_reg_22(.CP(n_62181), .D(n_40359), .CD(n_60988), .Q(iaddr
		[22]));
	notech_mux2 i_53348(.S(n_60143), .A(iaddr[22]), .B(n_36756), .Z(n_40359)
		);
	notech_reg addr_reg_23(.CP(n_62181), .D(n_40365), .CD(n_60988), .Q(iaddr
		[23]));
	notech_mux2 i_53356(.S(n_60143), .A(iaddr[23]), .B(n_36762), .Z(n_40365)
		);
	notech_reg addr_reg_24(.CP(n_62181), .D(n_40371), .CD(n_60988), .Q(iaddr
		[24]));
	notech_mux2 i_53364(.S(n_60143), .A(iaddr[24]), .B(n_36768), .Z(n_40371)
		);
	notech_reg addr_reg_25(.CP(n_62181), .D(n_40377), .CD(n_60988), .Q(iaddr
		[25]));
	notech_mux2 i_53372(.S(n_60143), .A(iaddr[25]), .B(n_36774), .Z(n_40377)
		);
	notech_nand3 i_52278169(.A(n_60258), .B(n_58375), .C(queue[25]), .Z(n_1394
		));
	notech_reg addr_reg_26(.CP(n_62181), .D(n_40383), .CD(n_60988), .Q(iaddr
		[26]));
	notech_mux2 i_53380(.S(n_60143), .A(iaddr[26]), .B(n_36780), .Z(n_40383)
		);
	notech_reg addr_reg_27(.CP(n_62181), .D(n_40389), .CD(n_60988), .Q(iaddr
		[27]));
	notech_mux2 i_53388(.S(n_60143), .A(iaddr[27]), .B(n_36786), .Z(n_40389)
		);
	notech_reg addr_reg_28(.CP(n_62181), .D(n_40395), .CD(n_60988), .Q(iaddr
		[28]));
	notech_mux2 i_53396(.S(n_60143), .A(iaddr[28]), .B(n_36792), .Z(n_40395)
		);
	notech_and4 i_1724996(.A(n_2196), .B(n_2195), .C(n_2190), .D(n_2194), .Z
		(squeue_1697089));
	notech_reg addr_reg_29(.CP(n_62179), .D(n_40401), .CD(n_60988), .Q(iaddr
		[29]));
	notech_mux2 i_53404(.S(n_60143), .A(iaddr[29]), .B(n_36798), .Z(n_40401)
		);
	notech_nand3 i_50478187(.A(n_57935), .B(n_58206), .C(queue[16]), .Z(n_1391
		));
	notech_reg addr_reg_30(.CP(n_62179), .D(n_40407), .CD(n_60988), .Q(iaddr
		[30]));
	notech_mux2 i_53412(.S(n_60143), .A(iaddr[30]), .B(n_36804), .Z(n_40407)
		);
	notech_reg addr_reg_31(.CP(n_62255), .D(n_40413), .CD(n_60988), .Q(iaddr
		[31]));
	notech_mux2 i_53420(.S(n_60143), .A(iaddr[31]), .B(n_36810), .Z(n_40413)
		);
	notech_reg code_req_reg(.CP(n_62255), .D(n_40419), .CD(n_60987), .Q(n_61560
		));
	notech_mux2 i_53428(.S(n_36824), .A(n_61549), .B(n_52396991), .Z(n_40419
		));
	notech_reg addrshft_reg_0(.CP(n_62255), .D(n_40425), .CD(n_60987), .Q(addrshft
		[0]));
	notech_mux2 i_53436(.S(\nbus_12119[0] ), .A(addrshft[0]), .B(n_36913), .Z
		(n_40425));
	notech_reg addrshft_reg_1(.CP(n_62255), .D(n_40431), .CD(n_60987), .Q(addrshft
		[1]));
	notech_mux2 i_53444(.S(\nbus_12119[0] ), .A(addrshft[1]), .B(n_36919), .Z
		(n_40431));
	notech_reg addrshft_reg_2(.CP(n_62255), .D(n_40437), .CD(n_60987), .Q(addrshft
		[2]));
	notech_mux2 i_53452(.S(\nbus_12119[0] ), .A(addrshft[2]), .B(n_36925), .Z
		(n_40437));
	notech_reg addrshft_reg_3(.CP(n_62255), .D(n_40443), .CD(n_60987), .Q(addrshft
		[3]));
	notech_mux2 i_53460(.S(\nbus_12119[0] ), .A(addrshft[3]), .B(n_36931), .Z
		(n_40443));
	notech_reg addrshft_reg_4(.CP(n_62255), .D(n_40449), .CD(n_60987), .Q(addrshft
		[4]));
	notech_mux2 i_53468(.S(\nbus_12119[0] ), .A(addrshft[4]), .B(n_20596673)
		, .Z(n_40449));
	notech_reg addrshft_reg_5(.CP(n_62255), .D(n_40455), .CD(n_60988), .Q(addrshft
		[5]));
	notech_mux2 i_53476(.S(\nbus_12119[0] ), .A(addrshft[5]), .B(n_52296990)
		, .Z(n_40455));
	notech_reg wptr_reg_0(.CP(n_62255), .D(n_40461), .CD(n_60987), .Q(wptr[0
		]));
	notech_mux2 i_53484(.S(n_42171), .A(wptr[0]), .B(n_30496772), .Z(n_40461
		));
	notech_reg wptr_reg_1(.CP(n_62255), .D(n_40467), .CD(n_60987), .Q(wptr[1
		]));
	notech_mux2 i_53492(.S(n_42171), .A(n_60277), .B(n_35007), .Z(n_40467)
		);
	notech_reg fault_wptr_reg_0(.CP(n_62255), .D(n_40473), .CD(n_60987), .Q(fault_wptr
		[0]));
	notech_mux2 i_53500(.S(\nbus_12115[0] ), .A(fault_wptr[0]), .B(n_42172),
		 .Z(n_40473));
	notech_reg fault_wptr_reg_1(.CP(n_62255), .D(n_40479), .CD(n_60982), .Q(fault_wptr
		[1]));
	notech_mux2 i_53508(.S(\nbus_12115[0] ), .A(fault_wptr[1]), .B(n_42173),
		 .Z(n_40479));
	notech_or2 i_49178200(.A(n_58247), .B(n_42193), .Z(n_1378));
	notech_reg pc_pg_fault_reg(.CP(n_62255), .D(n_40485), .CD(n_60982), .Q(pc_pg_fault
		));
	notech_mux2 i_53516(.S(n_42174), .A(pc_pg_fault), .B(n_42167), .Z(n_40485
		));
	notech_reg purge_cnt_reg_0(.CP(n_62255), .D(n_40491), .CD(n_60982), .Q(purge_cnt
		[0]));
	notech_mux2 i_53524(.S(\nbus_12118[0] ), .A(purge_cnt[0]), .B(n_29396761
		), .Z(n_40491));
	notech_reg purge_cnt_reg_1(.CP(n_62255), .D(n_40497), .CD(n_60982), .Q(purge_cnt
		[1]));
	notech_mux2 i_53532(.S(\nbus_12118[0] ), .A(purge_cnt[1]), .B(n_29496762
		), .Z(n_40497));
	notech_and4 i_1624995(.A(n_2182), .B(n_2181), .C(n_2176), .D(n_2180), .Z
		(squeue_1597090));
	notech_reg purge_cnt_reg_2(.CP(n_62255), .D(n_40503), .CD(n_60982), .Q(purge_cnt
		[2]));
	notech_mux2 i_53540(.S(\nbus_12118[0] ), .A(purge_cnt[2]), .B(n_29596763
		), .Z(n_40503));
	notech_nand3 i_47378218(.A(n_57935), .B(n_58206), .C(queue[15]), .Z(n_1375
		));
	notech_reg purge_cnt_reg_3(.CP(n_62255), .D(n_40509), .CD(n_60983), .Q(purge_cnt
		[3]));
	notech_mux2 i_53548(.S(\nbus_12118[0] ), .A(purge_cnt[3]), .B(n_29696764
		), .Z(n_40509));
	notech_reg purge_cnt_reg_4(.CP(n_62255), .D(n_40515), .CD(n_60983), .Q(purge_cnt
		[4]));
	notech_mux2 i_53556(.S(\nbus_12118[0] ), .A(purge_cnt[4]), .B(n_29796765
		), .Z(n_40515));
	notech_reg purge_cnt_reg_5(.CP(n_62179), .D(n_40521), .CD(n_60983), .Q(purge_cnt
		[5]));
	notech_mux2 i_53564(.S(\nbus_12118[0] ), .A(purge_cnt[5]), .B(n_29896766
		), .Z(n_40521));
	notech_reg purge_cnt_reg_6(.CP(n_62179), .D(n_40527), .CD(n_60982), .Q(purge_cnt
		[6]));
	notech_mux2 i_53572(.S(\nbus_12118[0] ), .A(purge_cnt[6]), .B(n_29996767
		), .Z(n_40527));
	notech_reg purge_cnt_reg_7(.CP(n_62179), .D(n_40533), .CD(n_60982), .Q(purge_cnt
		[7]));
	notech_mux2 i_53580(.S(\nbus_12118[0] ), .A(purge_cnt[7]), .B(n_30096768
		), .Z(n_40533));
	notech_reg purge_cnt_reg_8(.CP(n_62179), .D(n_40539), .CD(n_60982), .Q(purge_cnt
		[8]));
	notech_mux2 i_53588(.S(\nbus_12118[0] ), .A(purge_cnt[8]), .B(n_30196769
		), .Z(n_40539));
	notech_reg purge_cnt_reg_9(.CP(n_62179), .D(n_40545), .CD(n_60981), .Q(purge_cnt
		[9]));
	notech_mux2 i_53596(.S(\nbus_12118[0] ), .A(purge_cnt[9]), .B(n_30296770
		), .Z(n_40545));
	notech_reg purge_cnt_reg_10(.CP(n_62179), .D(n_40551), .CD(n_60982), .Q(purge_cnt
		[10]));
	notech_mux2 i_53604(.S(\nbus_12118[0] ), .A(purge_cnt[10]), .B(n_30396771
		), .Z(n_40551));
	notech_reg_set purge_reg(.CP(n_62179), .D(n_40557), .SD(n_60981), .Q(purge
		));
	notech_mux2 i_53612(.S(n_36952), .A(purge), .B(pc_pg_fault), .Z(n_40557)
		);
	notech_reg addrf_reg_0(.CP(n_62179), .D(iaddr[0]), .CD(n_60981), .Q(addrf
		[0]));
	notech_reg addrf_reg_1(.CP(n_62179), .D(iaddr[1]), .CD(n_60981), .Q(addrf
		[1]));
	notech_reg addrf_reg_2(.CP(n_62255), .D(iaddr[2]), .CD(n_60982), .Q(addrf
		[2]));
	notech_reg addrf_reg_3(.CP(n_62251), .D(iaddr[3]), .CD(n_60982), .Q(addrf
		[3]));
	notech_reg addrf_reg_4(.CP(n_62177), .D(iaddr[4]), .CD(n_60982), .Q(addrf
		[4]));
	notech_reg addrf_reg_5(.CP(n_62251), .D(iaddr[5]), .CD(n_60982), .Q(addrf
		[5]));
	notech_reg addrf_reg_6(.CP(n_62251), .D(iaddr[6]), .CD(n_60982), .Q(addrf
		[6]));
	notech_reg addrf_reg_7(.CP(n_62251), .D(iaddr[7]), .CD(n_60983), .Q(addrf
		[7]));
	notech_reg addrf_reg_8(.CP(n_62251), .D(iaddr[8]), .CD(n_60985), .Q(addrf
		[8]));
	notech_reg addrf_reg_9(.CP(n_62251), .D(iaddr[9]), .CD(n_60985), .Q(addrf
		[9]));
	notech_reg addrf_reg_10(.CP(n_62251), .D(iaddr[10]), .CD(n_60985), .Q(addrf
		[10]));
	notech_reg addrf_reg_11(.CP(n_62251), .D(iaddr[11]), .CD(n_60985), .Q(addrf
		[11]));
	notech_reg addrf_reg_12(.CP(n_62251), .D(iaddr[12]), .CD(n_60985), .Q(addrf
		[12]));
	notech_reg addrf_reg_13(.CP(n_62251), .D(iaddr[13]), .CD(n_60985), .Q(addrf
		[13]));
	notech_reg addrf_reg_14(.CP(n_62251), .D(iaddr[14]), .CD(n_60985), .Q(addrf
		[14]));
	notech_reg addrf_reg_15(.CP(n_62331), .D(iaddr[15]), .CD(n_60985), .Q(addrf
		[15]));
	notech_reg addrf_reg_16(.CP(n_62331), .D(iaddr[16]), .CD(n_60985), .Q(addrf
		[16]));
	notech_reg addrf_reg_17(.CP(n_62331), .D(iaddr[17]), .CD(n_60985), .Q(addrf
		[17]));
	notech_reg addrf_reg_18(.CP(n_62331), .D(iaddr[18]), .CD(n_60985), .Q(addrf
		[18]));
	notech_reg addrf_reg_19(.CP(n_62331), .D(iaddr[19]), .CD(n_60983), .Q(addrf
		[19]));
	notech_reg addrf_reg_20(.CP(n_62331), .D(iaddr[20]), .CD(n_60983), .Q(addrf
		[20]));
	notech_reg addrf_reg_21(.CP(n_62331), .D(iaddr[21]), .CD(n_60983), .Q(addrf
		[21]));
	notech_reg addrf_reg_22(.CP(n_62331), .D(iaddr[22]), .CD(n_60983), .Q(addrf
		[22]));
	notech_reg addrf_reg_23(.CP(n_62331), .D(iaddr[23]), .CD(n_60983), .Q(addrf
		[23]));
	notech_reg addrf_reg_24(.CP(n_62331), .D(iaddr[24]), .CD(n_60983), .Q(addrf
		[24]));
	notech_reg addrf_reg_25(.CP(n_62331), .D(iaddr[25]), .CD(n_60983), .Q(addrf
		[25]));
	notech_reg addrf_reg_26(.CP(n_62331), .D(iaddr[26]), .CD(n_60983), .Q(addrf
		[26]));
	notech_reg addrf_reg_27(.CP(n_62331), .D(iaddr[27]), .CD(n_60983), .Q(addrf
		[27]));
	notech_reg addrf_reg_28(.CP(n_62331), .D(iaddr[28]), .CD(n_60983), .Q(addrf
		[28]));
	notech_reg addrf_reg_29(.CP(n_62331), .D(iaddr[29]), .CD(n_60993), .Q(addrf
		[29]));
	notech_reg addrf_reg_30(.CP(n_62331), .D(iaddr[30]), .CD(n_60994), .Q(addrf
		[30]));
	notech_reg addrf_reg_31(.CP(n_62331), .D(iaddr[31]), .CD(n_60993), .Q(addrf
		[31]));
	notech_reg queue_reg_0(.CP(n_62331), .D(n_40627), .CD(n_60993), .Q(queue
		[0]));
	notech_mux2 i_53748(.S(n_54326), .A(queue[0]), .B(n_35075), .Z(n_40627)
		);
	notech_reg queue_reg_1(.CP(n_62251), .D(n_40633), .CD(n_60993), .Q(queue
		[1]));
	notech_mux2 i_53756(.S(n_54326), .A(queue[1]), .B(n_35081), .Z(n_40633)
		);
	notech_reg queue_reg_2(.CP(n_62177), .D(n_40639), .CD(n_60994), .Q(queue
		[2]));
	notech_mux2 i_53764(.S(n_54326), .A(queue[2]), .B(n_35087), .Z(n_40639)
		);
	notech_reg queue_reg_3(.CP(n_62253), .D(n_40645), .CD(n_60994), .Q(queue
		[3]));
	notech_mux2 i_53772(.S(n_54326), .A(queue[3]), .B(n_35093), .Z(n_40645)
		);
	notech_or2 i_46078231(.A(n_58266), .B(n_42184), .Z(n_1362));
	notech_reg queue_reg_4(.CP(n_62253), .D(n_40651), .CD(n_60994), .Q(queue
		[4]));
	notech_mux2 i_53780(.S(n_54326), .A(queue[4]), .B(n_35099), .Z(n_40651)
		);
	notech_reg queue_reg_5(.CP(n_62253), .D(n_40657), .CD(n_60994), .Q(queue
		[5]));
	notech_mux2 i_53788(.S(n_54326), .A(queue[5]), .B(n_35105), .Z(n_40657)
		);
	notech_reg queue_reg_6(.CP(n_62253), .D(n_40663), .CD(n_60994), .Q(queue
		[6]));
	notech_mux2 i_53796(.S(n_54326), .A(queue[6]), .B(n_35111), .Z(n_40663)
		);
	notech_and4 i_1424993(.A(n_2168), .B(n_2167), .C(n_2162), .D(n_2166), .Z
		(squeue_1397091));
	notech_reg queue_reg_7(.CP(n_62253), .D(n_40669), .CD(n_60993), .Q(queue
		[7]));
	notech_mux2 i_53804(.S(n_54326), .A(queue[7]), .B(n_35117), .Z(n_40669)
		);
	notech_nand3 i_44278249(.A(n_57935), .B(n_58206), .C(queue[13]), .Z(n_1359
		));
	notech_reg queue_reg_8(.CP(n_62253), .D(n_40675), .CD(n_60993), .Q(queue
		[8]));
	notech_mux2 i_53812(.S(n_54326), .A(queue[8]), .B(n_35123), .Z(n_40675)
		);
	notech_reg queue_reg_9(.CP(n_62253), .D(n_40681), .CD(n_60993), .Q(queue
		[9]));
	notech_mux2 i_53820(.S(n_54326), .A(queue[9]), .B(n_35129), .Z(n_40681)
		);
	notech_reg queue_reg_10(.CP(n_62253), .D(n_40687), .CD(n_60993), .Q(queue
		[10]));
	notech_mux2 i_53828(.S(n_54326), .A(queue[10]), .B(n_35135), .Z(n_40687)
		);
	notech_reg queue_reg_11(.CP(n_62253), .D(n_40693), .CD(n_60992), .Q(queue
		[11]));
	notech_mux2 i_53836(.S(n_54326), .A(queue[11]), .B(n_35141), .Z(n_40693)
		);
	notech_reg queue_reg_12(.CP(n_62253), .D(n_40699), .CD(n_60993), .Q(queue
		[12]));
	notech_mux2 i_53844(.S(n_54326), .A(queue[12]), .B(n_35147), .Z(n_40699)
		);
	notech_reg queue_reg_13(.CP(n_62253), .D(n_40705), .CD(n_60993), .Q(queue
		[13]));
	notech_mux2 i_53852(.S(n_54326), .A(queue[13]), .B(n_35153), .Z(n_40705)
		);
	notech_reg queue_reg_14(.CP(n_62253), .D(n_40711), .CD(n_60993), .Q(queue
		[14]));
	notech_mux2 i_53860(.S(n_54326), .A(queue[14]), .B(n_35159), .Z(n_40711)
		);
	notech_reg queue_reg_15(.CP(n_62253), .D(n_40717), .CD(n_60993), .Q(queue
		[15]));
	notech_mux2 i_53868(.S(n_54326), .A(queue[15]), .B(n_35165), .Z(n_40717)
		);
	notech_reg queue_reg_16(.CP(n_62253), .D(n_40723), .CD(n_60993), .Q(queue
		[16]));
	notech_mux2 i_53876(.S(n_54324), .A(queue[16]), .B(n_35171), .Z(n_40723)
		);
	notech_reg queue_reg_17(.CP(n_62253), .D(n_40729), .CD(n_60993), .Q(queue
		[17]));
	notech_mux2 i_53884(.S(n_54324), .A(queue[17]), .B(n_35177), .Z(n_40729)
		);
	notech_reg queue_reg_18(.CP(n_62253), .D(n_40735), .CD(n_60994), .Q(queue
		[18]));
	notech_mux2 i_53892(.S(n_54324), .A(queue[18]), .B(n_35183), .Z(n_40735)
		);
	notech_reg queue_reg_19(.CP(n_62253), .D(n_40741), .CD(n_60995), .Q(queue
		[19]));
	notech_mux2 i_53900(.S(n_54324), .A(queue[19]), .B(n_35189), .Z(n_40741)
		);
	notech_reg queue_reg_20(.CP(n_62253), .D(n_40747), .CD(n_60995), .Q(queue
		[20]));
	notech_mux2 i_53908(.S(n_54324), .A(queue[20]), .B(n_35195), .Z(n_40747)
		);
	notech_nand3 i_42978262(.A(n_60258), .B(n_58375), .C(queue[21]), .Z(n_1346
		));
	notech_reg queue_reg_21(.CP(n_62253), .D(n_40753), .CD(n_60995), .Q(queue
		[21]));
	notech_mux2 i_53916(.S(n_54324), .A(queue[21]), .B(n_35201), .Z(n_40753)
		);
	notech_reg queue_reg_22(.CP(n_62177), .D(n_40759), .CD(n_60995), .Q(queue
		[22]));
	notech_mux2 i_53924(.S(n_54324), .A(queue[22]), .B(n_35207), .Z(n_40759)
		);
	notech_reg queue_reg_23(.CP(n_62177), .D(n_40765), .CD(n_60995), .Q(queue
		[23]));
	notech_mux2 i_53932(.S(n_54324), .A(queue[23]), .B(n_35213), .Z(n_40765)
		);
	notech_and4 i_1324992(.A(n_2154), .B(n_2153), .C(n_2148), .D(n_2152), .Z
		(squeue_1297092));
	notech_reg queue_reg_24(.CP(n_62177), .D(n_40771), .CD(n_60995), .Q(queue
		[24]));
	notech_mux2 i_53940(.S(n_54324), .A(queue[24]), .B(n_35219), .Z(n_40771)
		);
	notech_nand3 i_41178280(.A(n_57935), .B(n_58206), .C(queue[12]), .Z(n_1343
		));
	notech_reg queue_reg_25(.CP(n_62177), .D(n_40777), .CD(n_60995), .Q(queue
		[25]));
	notech_mux2 i_53948(.S(n_54324), .A(queue[25]), .B(n_35225), .Z(n_40777)
		);
	notech_reg queue_reg_26(.CP(n_62177), .D(n_40783), .CD(n_60995), .Q(queue
		[26]));
	notech_mux2 i_53956(.S(n_54324), .A(queue[26]), .B(n_35231), .Z(n_40783)
		);
	notech_reg queue_reg_27(.CP(n_62177), .D(n_40789), .CD(n_60995), .Q(queue
		[27]));
	notech_mux2 i_53964(.S(n_54324), .A(queue[27]), .B(n_35237), .Z(n_40789)
		);
	notech_reg queue_reg_28(.CP(n_62177), .D(n_40795), .CD(n_60995), .Q(queue
		[28]));
	notech_mux2 i_53972(.S(n_54324), .A(queue[28]), .B(n_35243), .Z(n_40795)
		);
	notech_reg queue_reg_29(.CP(n_62177), .D(n_40801), .CD(n_60995), .Q(queue
		[29]));
	notech_mux2 i_53980(.S(n_54324), .A(queue[29]), .B(n_35249), .Z(n_40801)
		);
	notech_reg queue_reg_30(.CP(n_62177), .D(n_40807), .CD(n_60994), .Q(queue
		[30]));
	notech_mux2 i_53988(.S(n_54324), .A(queue[30]), .B(n_35255), .Z(n_40807)
		);
	notech_reg queue_reg_31(.CP(n_62331), .D(n_40813), .CD(n_60994), .Q(queue
		[31]));
	notech_mux2 i_53996(.S(n_54324), .A(queue[31]), .B(n_35261), .Z(n_40813)
		);
	notech_reg queue_reg_32(.CP(n_62245), .D(n_40819), .CD(n_60994), .Q(queue
		[32]));
	notech_mux2 i_54004(.S(n_54331), .A(queue[32]), .B(n_35267), .Z(n_40819)
		);
	notech_reg queue_reg_33(.CP(n_62245), .D(n_40825), .CD(n_60994), .Q(queue
		[33]));
	notech_mux2 i_54012(.S(n_54331), .A(queue[33]), .B(n_35273), .Z(n_40825)
		);
	notech_reg queue_reg_34(.CP(n_62245), .D(n_40831), .CD(n_60994), .Q(queue
		[34]));
	notech_mux2 i_54020(.S(n_54331), .A(queue[34]), .B(n_35279), .Z(n_40831)
		);
	notech_reg queue_reg_35(.CP(n_62245), .D(n_40837), .CD(n_60995), .Q(queue
		[35]));
	notech_mux2 i_54028(.S(n_54331), .A(queue[35]), .B(n_35285), .Z(n_40837)
		);
	notech_reg queue_reg_36(.CP(n_62245), .D(n_40843), .CD(n_60995), .Q(queue
		[36]));
	notech_mux2 i_54036(.S(n_54331), .A(queue[36]), .B(n_35291), .Z(n_40843)
		);
	notech_reg queue_reg_37(.CP(n_62245), .D(n_40849), .CD(n_60995), .Q(queue
		[37]));
	notech_mux2 i_54044(.S(n_54331), .A(queue[37]), .B(n_35297), .Z(n_40849)
		);
	notech_nand3 i_39878293(.A(n_60258), .B(n_58379), .C(queue[20]), .Z(n_1330
		));
	notech_reg queue_reg_38(.CP(n_62245), .D(n_40855), .CD(n_60994), .Q(queue
		[38]));
	notech_mux2 i_54052(.S(n_54331), .A(queue[38]), .B(n_35303), .Z(n_40855)
		);
	notech_reg queue_reg_39(.CP(n_62245), .D(n_40861), .CD(n_60994), .Q(queue
		[39]));
	notech_mux2 i_54060(.S(n_54331), .A(queue[39]), .B(n_35309), .Z(n_40861)
		);
	notech_reg queue_reg_40(.CP(n_62245), .D(n_40867), .CD(n_60989), .Q(queue
		[40]));
	notech_mux2 i_54068(.S(n_54331), .A(queue[40]), .B(n_35315), .Z(n_40867)
		);
	notech_and4 i_1224991(.A(n_2140), .B(n_2139), .C(n_2134), .D(n_2138), .Z
		(squeue_1197093));
	notech_reg queue_reg_41(.CP(n_62245), .D(n_40873), .CD(n_60989), .Q(queue
		[41]));
	notech_mux2 i_54076(.S(n_54331), .A(queue[41]), .B(n_35321), .Z(n_40873)
		);
	notech_nand3 i_38078311(.A(n_57935), .B(n_58206), .C(queue[11]), .Z(n_1327
		));
	notech_reg queue_reg_42(.CP(n_62245), .D(n_40879), .CD(n_60989), .Q(queue
		[42]));
	notech_mux2 i_54084(.S(n_54331), .A(queue[42]), .B(n_35327), .Z(n_40879)
		);
	notech_reg queue_reg_43(.CP(n_62327), .D(n_40885), .CD(n_60989), .Q(queue
		[43]));
	notech_mux2 i_54092(.S(n_54331), .A(queue[43]), .B(n_35333), .Z(n_40885)
		);
	notech_reg queue_reg_44(.CP(n_62327), .D(n_40891), .CD(n_60989), .Q(queue
		[44]));
	notech_mux2 i_54100(.S(n_54331), .A(queue[44]), .B(n_35339), .Z(n_40891)
		);
	notech_reg queue_reg_45(.CP(n_62327), .D(n_40897), .CD(n_60991), .Q(queue
		[45]));
	notech_mux2 i_54108(.S(n_54331), .A(queue[45]), .B(n_35345), .Z(n_40897)
		);
	notech_reg queue_reg_46(.CP(n_62327), .D(n_40903), .CD(n_60991), .Q(queue
		[46]));
	notech_mux2 i_54116(.S(n_54331), .A(queue[46]), .B(n_35351), .Z(n_40903)
		);
	notech_reg queue_reg_47(.CP(n_62327), .D(n_40909), .CD(n_60991), .Q(queue
		[47]));
	notech_mux2 i_54124(.S(n_54331), .A(queue[47]), .B(n_35357), .Z(n_40909)
		);
	notech_reg queue_reg_48(.CP(n_62327), .D(n_40915), .CD(n_60991), .Q(queue
		[48]));
	notech_mux2 i_54132(.S(n_54329), .A(queue[48]), .B(n_35363), .Z(n_40915)
		);
	notech_reg queue_reg_49(.CP(n_62327), .D(n_40921), .CD(n_60991), .Q(queue
		[49]));
	notech_mux2 i_54140(.S(n_54329), .A(queue[49]), .B(n_35369), .Z(n_40921)
		);
	notech_reg queue_reg_50(.CP(n_62327), .D(n_40927), .CD(n_60989), .Q(queue
		[50]));
	notech_mux2 i_54148(.S(n_54329), .A(queue[50]), .B(n_35375), .Z(n_40927)
		);
	notech_reg queue_reg_51(.CP(n_62327), .D(n_40933), .CD(n_60989), .Q(queue
		[51]));
	notech_mux2 i_54156(.S(n_54329), .A(queue[51]), .B(n_35381), .Z(n_40933)
		);
	notech_reg queue_reg_52(.CP(n_62327), .D(n_40939), .CD(n_60989), .Q(queue
		[52]));
	notech_mux2 i_54164(.S(n_54329), .A(queue[52]), .B(n_35387), .Z(n_40939)
		);
	notech_reg queue_reg_53(.CP(n_62327), .D(n_40945), .CD(n_60989), .Q(queue
		[53]));
	notech_mux2 i_54172(.S(n_54329), .A(queue[53]), .B(n_35393), .Z(n_40945)
		);
	notech_reg queue_reg_54(.CP(n_62327), .D(n_40951), .CD(n_60988), .Q(queue
		[54]));
	notech_mux2 i_54180(.S(n_54329), .A(queue[54]), .B(n_35399), .Z(n_40951)
		);
	notech_nand3 i_36778324(.A(n_60262), .B(n_58379), .C(queue[19]), .Z(n_1308
		));
	notech_reg queue_reg_55(.CP(n_62327), .D(n_40957), .CD(n_60988), .Q(queue
		[55]));
	notech_mux2 i_54188(.S(n_54329), .A(queue[55]), .B(n_35405), .Z(n_40957)
		);
	notech_reg queue_reg_56(.CP(n_62327), .D(n_40963), .CD(n_60989), .Q(queue
		[56]));
	notech_mux2 i_54196(.S(n_54329), .A(queue[56]), .B(n_35411), .Z(n_40963)
		);
	notech_reg queue_reg_57(.CP(n_62327), .D(n_40969), .CD(n_60989), .Q(queue
		[57]));
	notech_mux2 i_54204(.S(n_54329), .A(queue[57]), .B(n_35417), .Z(n_40969)
		);
	notech_and4 i_1124990(.A(n_2126), .B(n_2125), .C(n_2120), .D(n_2124), .Z
		(squeue_1097094));
	notech_reg queue_reg_58(.CP(n_62327), .D(n_40975), .CD(n_60989), .Q(queue
		[58]));
	notech_mux2 i_54212(.S(n_54329), .A(queue[58]), .B(n_35423), .Z(n_40975)
		);
	notech_nand3 i_34978342(.A(n_57935), .B(n_58206), .C(queue[10]), .Z(n_1303
		));
	notech_reg queue_reg_59(.CP(n_62327), .D(n_40981), .CD(n_60989), .Q(queue
		[59]));
	notech_mux2 i_54220(.S(n_54329), .A(queue[59]), .B(n_35429), .Z(n_40981)
		);
	notech_reg queue_reg_60(.CP(n_62327), .D(n_40987), .CD(n_60989), .Q(queue
		[60]));
	notech_mux2 i_54228(.S(n_54329), .A(queue[60]), .B(n_35435), .Z(n_40987)
		);
	notech_reg queue_reg_61(.CP(n_62327), .D(n_40993), .CD(n_60991), .Q(queue
		[61]));
	notech_mux2 i_54236(.S(n_54329), .A(queue[61]), .B(n_35441), .Z(n_40993)
		);
	notech_reg queue_reg_62(.CP(n_62375), .D(n_40999), .CD(n_60992), .Q(queue
		[62]));
	notech_mux2 i_54244(.S(n_54329), .A(queue[62]), .B(n_35447), .Z(n_40999)
		);
	notech_reg queue_reg_63(.CP(n_62375), .D(n_41005), .CD(n_60992), .Q(queue
		[63]));
	notech_mux2 i_54252(.S(n_54329), .A(queue[63]), .B(n_35453), .Z(n_41005)
		);
	notech_reg queue_reg_64(.CP(n_62375), .D(n_41011), .CD(n_60992), .Q(queue
		[64]));
	notech_mux2 i_54260(.S(n_54316), .A(queue[64]), .B(n_35459), .Z(n_41011)
		);
	notech_reg queue_reg_65(.CP(n_62375), .D(n_41017), .CD(n_60992), .Q(queue
		[65]));
	notech_mux2 i_54268(.S(n_54316), .A(queue[65]), .B(n_35465), .Z(n_41017)
		);
	notech_reg queue_reg_66(.CP(n_62375), .D(n_41023), .CD(n_60992), .Q(queue
		[66]));
	notech_mux2 i_54276(.S(n_54316), .A(queue[66]), .B(n_35471), .Z(n_41023)
		);
	notech_reg queue_reg_67(.CP(n_62375), .D(n_41029), .CD(n_60992), .Q(queue
		[67]));
	notech_mux2 i_54284(.S(n_54316), .A(queue[67]), .B(n_35477), .Z(n_41029)
		);
	notech_reg queue_reg_68(.CP(n_62375), .D(n_41035), .CD(n_60992), .Q(queue
		[68]));
	notech_mux2 i_54292(.S(n_54316), .A(queue[68]), .B(n_35483), .Z(n_41035)
		);
	notech_reg queue_reg_69(.CP(n_62375), .D(n_41041), .CD(n_60992), .Q(queue
		[69]));
	notech_mux2 i_54300(.S(n_54316), .A(queue[69]), .B(n_35489), .Z(n_41041)
		);
	notech_reg queue_reg_70(.CP(n_62375), .D(n_41047), .CD(n_60992), .Q(queue
		[70]));
	notech_mux2 i_54308(.S(n_54316), .A(queue[70]), .B(n_35495), .Z(n_41047)
		);
	notech_reg queue_reg_71(.CP(n_62375), .D(n_41053), .CD(n_60992), .Q(queue
		[71]));
	notech_mux2 i_54316(.S(n_54316), .A(queue[71]), .B(n_35501), .Z(n_41053)
		);
	notech_nand3 i_33678355(.A(n_60262), .B(n_58379), .C(queue[18]), .Z(n_1282
		));
	notech_reg queue_reg_72(.CP(n_62375), .D(n_41059), .CD(n_60992), .Q(queue
		[72]));
	notech_mux2 i_54324(.S(n_54316), .A(queue[72]), .B(n_35507), .Z(n_41059)
		);
	notech_reg queue_reg_73(.CP(n_62375), .D(n_41065), .CD(n_60991), .Q(queue
		[73]));
	notech_mux2 i_54332(.S(n_54316), .A(queue[73]), .B(n_35513), .Z(n_41065)
		);
	notech_reg queue_reg_74(.CP(n_62375), .D(n_41071), .CD(n_60991), .Q(queue
		[74]));
	notech_mux2 i_54340(.S(n_54316), .A(queue[74]), .B(n_35519), .Z(n_41071)
		);
	notech_and4 i_1024989(.A(n_2112), .B(n_2111), .C(n_2106), .D(n_2110), .Z
		(squeue_997095));
	notech_reg queue_reg_75(.CP(n_62375), .D(n_41077), .CD(n_60991), .Q(queue
		[75]));
	notech_mux2 i_54348(.S(n_54316), .A(queue[75]), .B(n_35525), .Z(n_41077)
		);
	notech_nand3 i_31878373(.A(n_57935), .B(n_58206), .C(queue[9]), .Z(n_1279
		));
	notech_reg queue_reg_76(.CP(n_62375), .D(n_41083), .CD(n_60991), .Q(queue
		[76]));
	notech_mux2 i_54356(.S(n_54316), .A(queue[76]), .B(n_35531), .Z(n_41083)
		);
	notech_reg queue_reg_77(.CP(n_62375), .D(n_41089), .CD(n_60991), .Q(queue
		[77]));
	notech_mux2 i_54364(.S(n_54316), .A(queue[77]), .B(n_35537), .Z(n_41089)
		);
	notech_reg queue_reg_78(.CP(n_62375), .D(n_41095), .CD(n_60992), .Q(queue
		[78]));
	notech_mux2 i_54372(.S(n_54316), .A(queue[78]), .B(n_35543), .Z(n_41095)
		);
	notech_reg queue_reg_79(.CP(n_62375), .D(n_41101), .CD(n_60992), .Q(queue
		[79]));
	notech_mux2 i_54380(.S(n_54316), .A(queue[79]), .B(n_35549), .Z(n_41101)
		);
	notech_reg queue_reg_80(.CP(n_62375), .D(n_41107), .CD(n_60991), .Q(queue
		[80]));
	notech_mux2 i_54388(.S(n_54314), .A(queue[80]), .B(n_35555), .Z(n_41107)
		);
	notech_reg queue_reg_81(.CP(n_62375), .D(n_41113), .CD(n_60991), .Q(queue
		[81]));
	notech_mux2 i_54396(.S(n_54314), .A(queue[81]), .B(n_35561), .Z(n_41113)
		);
	notech_reg queue_reg_82(.CP(n_62325), .D(n_41119), .CD(n_60991), .Q(queue
		[82]));
	notech_mux2 i_54404(.S(n_54314), .A(queue[82]), .B(n_35567), .Z(n_41119)
		);
	notech_reg queue_reg_83(.CP(n_62325), .D(n_41125), .CD(n_60981), .Q(queue
		[83]));
	notech_mux2 i_54412(.S(n_54314), .A(queue[83]), .B(n_35573), .Z(n_41125)
		);
	notech_reg queue_reg_84(.CP(n_62325), .D(n_41131), .CD(n_60971), .Q(queue
		[84]));
	notech_mux2 i_54420(.S(n_54314), .A(queue[84]), .B(n_35579), .Z(n_41131)
		);
	notech_reg queue_reg_85(.CP(n_62325), .D(n_41137), .CD(n_60971), .Q(queue
		[85]));
	notech_mux2 i_54428(.S(n_54314), .A(queue[85]), .B(n_35585), .Z(n_41137)
		);
	notech_reg queue_reg_86(.CP(n_62325), .D(n_41143), .CD(n_60971), .Q(queue
		[86]));
	notech_mux2 i_54436(.S(n_54314), .A(queue[86]), .B(n_35591), .Z(n_41143)
		);
	notech_reg queue_reg_87(.CP(n_62325), .D(n_41149), .CD(n_60971), .Q(queue
		[87]));
	notech_mux2 i_54444(.S(n_54314), .A(queue[87]), .B(n_35597), .Z(n_41149)
		);
	notech_reg queue_reg_88(.CP(n_62325), .D(n_41155), .CD(n_60971), .Q(queue
		[88]));
	notech_mux2 i_54452(.S(n_54314), .A(queue[88]), .B(n_35603), .Z(n_41155)
		);
	notech_nand3 i_30578386(.A(n_60262), .B(n_58379), .C(queue[17]), .Z(n_1266
		));
	notech_reg queue_reg_89(.CP(n_62325), .D(n_41161), .CD(n_60971), .Q(queue
		[89]));
	notech_mux2 i_54460(.S(n_54314), .A(queue[89]), .B(n_35609), .Z(n_41161)
		);
	notech_reg queue_reg_90(.CP(n_62325), .D(n_41167), .CD(n_60971), .Q(queue
		[90]));
	notech_mux2 i_54468(.S(n_54314), .A(queue[90]), .B(n_35615), .Z(n_41167)
		);
	notech_reg queue_reg_91(.CP(n_62325), .D(n_41173), .CD(n_60971), .Q(queue
		[91]));
	notech_mux2 i_54476(.S(n_54314), .A(queue[91]), .B(n_35621), .Z(n_41173)
		);
	notech_and4 i_924988(.A(n_2098), .B(n_2097), .C(n_2092), .D(n_2096), .Z(squeue_897096
		));
	notech_reg queue_reg_92(.CP(n_62325), .D(n_41179), .CD(n_60971), .Q(queue
		[92]));
	notech_mux2 i_54484(.S(n_54314), .A(queue[92]), .B(n_35627), .Z(n_41179)
		);
	notech_nand3 i_28778404(.A(n_57935), .B(n_58209), .C(queue[8]), .Z(n_1263
		));
	notech_reg queue_reg_93(.CP(n_62325), .D(n_41185), .CD(n_60971), .Q(queue
		[93]));
	notech_mux2 i_54492(.S(n_54314), .A(queue[93]), .B(n_35633), .Z(n_41185)
		);
	notech_reg queue_reg_94(.CP(n_62329), .D(n_41191), .CD(n_60971), .Q(queue
		[94]));
	notech_mux2 i_54500(.S(n_54314), .A(queue[94]), .B(n_35639), .Z(n_41191)
		);
	notech_reg queue_reg_95(.CP(n_62247), .D(n_41197), .CD(n_60970), .Q(queue
		[95]));
	notech_mux2 i_54508(.S(n_54314), .A(queue[95]), .B(n_35645), .Z(n_41197)
		);
	notech_reg queue_reg_96(.CP(n_62247), .D(n_41203), .CD(n_60970), .Q(queue
		[96]));
	notech_mux2 i_54516(.S(n_54321), .A(queue[96]), .B(n_35651), .Z(n_41203)
		);
	notech_reg queue_reg_97(.CP(n_62247), .D(n_41209), .CD(n_60970), .Q(queue
		[97]));
	notech_mux2 i_54524(.S(n_54321), .A(queue[97]), .B(n_35657), .Z(n_41209)
		);
	notech_reg queue_reg_98(.CP(n_62247), .D(n_41215), .CD(n_60970), .Q(queue
		[98]));
	notech_mux2 i_54532(.S(n_54321), .A(queue[98]), .B(n_35663), .Z(n_41215)
		);
	notech_reg queue_reg_99(.CP(n_62247), .D(n_41221), .CD(n_60970), .Q(queue
		[99]));
	notech_mux2 i_54540(.S(n_54321), .A(queue[99]), .B(n_35669), .Z(n_41221)
		);
	notech_reg queue_reg_100(.CP(n_62247), .D(n_41227), .CD(n_60970), .Q(queue
		[100]));
	notech_mux2 i_54548(.S(n_54321), .A(queue[100]), .B(n_35675), .Z(n_41227
		));
	notech_reg queue_reg_101(.CP(n_62247), .D(n_41233), .CD(n_60971), .Q(queue
		[101]));
	notech_mux2 i_54556(.S(n_54321), .A(queue[101]), .B(n_35681), .Z(n_41233
		));
	notech_reg queue_reg_102(.CP(n_62247), .D(n_41239), .CD(n_60970), .Q(queue
		[102]));
	notech_mux2 i_54564(.S(n_54321), .A(queue[102]), .B(n_35687), .Z(n_41239
		));
	notech_reg queue_reg_103(.CP(n_62247), .D(n_41245), .CD(n_60970), .Q(queue
		[103]));
	notech_mux2 i_54572(.S(n_54321), .A(queue[103]), .B(n_35693), .Z(n_41245
		));
	notech_reg queue_reg_104(.CP(n_62329), .D(n_41251), .CD(n_60970), .Q(queue
		[104]));
	notech_mux2 i_54580(.S(n_54321), .A(queue[104]), .B(n_35699), .Z(n_41251
		));
	notech_reg queue_reg_105(.CP(n_62329), .D(n_41257), .CD(n_60971), .Q(queue
		[105]));
	notech_mux2 i_54588(.S(n_54321), .A(queue[105]), .B(n_35705), .Z(n_41257
		));
	notech_or2 i_27478417(.A(n_58228), .B(n_42193), .Z(n_1250));
	notech_reg queue_reg_106(.CP(n_62329), .D(n_41263), .CD(n_60974), .Q(queue
		[106]));
	notech_mux2 i_54596(.S(n_54321), .A(queue[106]), .B(n_35711), .Z(n_41263
		));
	notech_reg queue_reg_107(.CP(n_62329), .D(n_41269), .CD(n_60974), .Q(queue
		[107]));
	notech_mux2 i_54604(.S(n_54321), .A(queue[107]), .B(n_35717), .Z(n_41269
		));
	notech_reg queue_reg_108(.CP(n_62329), .D(n_41275), .CD(n_60973), .Q(queue
		[108]));
	notech_mux2 i_54612(.S(n_54321), .A(queue[108]), .B(n_35723), .Z(n_41275
		));
	notech_and4 i_724986(.A(n_2084), .B(n_2083), .C(n_2078), .D(n_2082), .Z(squeue_697097
		));
	notech_reg queue_reg_109(.CP(n_62329), .D(n_41281), .CD(n_60973), .Q(queue
		[109]));
	notech_mux2 i_54620(.S(n_54321), .A(queue[109]), .B(n_35729), .Z(n_41281
		));
	notech_nand3 i_25678435(.A(n_57935), .B(n_58209), .C(queue[6]), .Z(n_1247
		));
	notech_reg queue_reg_110(.CP(n_62329), .D(n_41287), .CD(n_60973), .Q(queue
		[110]));
	notech_mux2 i_54628(.S(n_54321), .A(queue[110]), .B(n_35735), .Z(n_41287
		));
	notech_reg queue_reg_111(.CP(n_62329), .D(n_41293), .CD(n_60974), .Q(queue
		[111]));
	notech_mux2 i_54636(.S(n_54321), .A(queue[111]), .B(n_35741), .Z(n_41293
		));
	notech_reg queue_reg_112(.CP(n_62329), .D(n_41299), .CD(n_60974), .Q(queue
		[112]));
	notech_mux2 i_54644(.S(n_54319), .A(queue[112]), .B(n_35747), .Z(n_41299
		));
	notech_reg queue_reg_113(.CP(n_62329), .D(n_41305), .CD(n_60974), .Q(queue
		[113]));
	notech_mux2 i_54652(.S(n_54319), .A(queue[113]), .B(n_35753), .Z(n_41305
		));
	notech_reg queue_reg_114(.CP(n_62329), .D(n_41311), .CD(n_60974), .Q(queue
		[114]));
	notech_mux2 i_54660(.S(n_54319), .A(queue[114]), .B(n_35759), .Z(n_41311
		));
	notech_reg queue_reg_115(.CP(n_62329), .D(n_41317), .CD(n_60974), .Q(queue
		[115]));
	notech_mux2 i_54668(.S(n_54319), .A(queue[115]), .B(n_35765), .Z(n_41317
		));
	notech_reg queue_reg_116(.CP(n_62329), .D(n_41323), .CD(n_60973), .Q(queue
		[116]));
	notech_mux2 i_54676(.S(n_54319), .A(queue[116]), .B(n_35771), .Z(n_41323
		));
	notech_reg queue_reg_117(.CP(n_62329), .D(n_41329), .CD(n_60973), .Q(queue
		[117]));
	notech_mux2 i_54684(.S(n_54319), .A(queue[117]), .B(n_35777), .Z(n_41329
		));
	notech_reg queue_reg_118(.CP(n_62329), .D(n_41335), .CD(n_60973), .Q(queue
		[118]));
	notech_mux2 i_54692(.S(n_54319), .A(queue[118]), .B(n_35783), .Z(n_41335
		));
	notech_reg queue_reg_119(.CP(n_62329), .D(n_41341), .CD(n_60973), .Q(queue
		[119]));
	notech_mux2 i_54700(.S(n_54319), .A(queue[119]), .B(n_35789), .Z(n_41341
		));
	notech_reg queue_reg_120(.CP(n_62329), .D(n_41347), .CD(n_60973), .Q(queue
		[120]));
	notech_mux2 i_54708(.S(n_54319), .A(queue[120]), .B(n_35795), .Z(n_41347
		));
	notech_reg queue_reg_121(.CP(n_62329), .D(n_41353), .CD(n_60973), .Q(queue
		[121]));
	notech_mux2 i_54716(.S(n_54319), .A(queue[121]), .B(n_35801), .Z(n_41353
		));
	notech_reg queue_reg_122(.CP(n_62247), .D(n_41359), .CD(n_60973), .Q(queue
		[122]));
	notech_mux2 i_54724(.S(n_54319), .A(queue[122]), .B(n_35807), .Z(n_41359
		));
	notech_nand3 i_24378448(.A(queue[14]), .B(n_60262), .C(n_58379), .Z(n_1234
		));
	notech_reg queue_reg_123(.CP(n_62247), .D(n_41365), .CD(n_60973), .Q(queue
		[123]));
	notech_mux2 i_54732(.S(n_54319), .A(queue[123]), .B(n_35813), .Z(n_41365
		));
	notech_reg queue_reg_124(.CP(n_62249), .D(n_41371), .CD(n_60973), .Q(queue
		[124]));
	notech_mux2 i_54740(.S(n_54319), .A(queue[124]), .B(n_35819), .Z(n_41371
		));
	notech_reg queue_reg_125(.CP(n_62249), .D(n_41377), .CD(n_60973), .Q(queue
		[125]));
	notech_mux2 i_54748(.S(n_54319), .A(queue[125]), .B(n_35825), .Z(n_41377
		));
	notech_and4 i_624985(.A(n_2070), .B(n_2069), .C(n_2064), .D(n_2068), .Z(squeue_597098
		));
	notech_reg queue_reg_126(.CP(n_62249), .D(n_41383), .CD(n_60973), .Q(queue
		[126]));
	notech_mux2 i_54756(.S(n_54319), .A(queue[126]), .B(n_35831), .Z(n_41383
		));
	notech_nand3 i_22578466(.A(n_57935), .B(n_58209), .C(queue[5]), .Z(n_1231
		));
	notech_reg queue_reg_127(.CP(n_62249), .D(n_41389), .CD(n_60968), .Q(queue
		[127]));
	notech_mux2 i_54764(.S(n_54319), .A(queue[127]), .B(n_35837), .Z(n_41389
		));
	notech_reg queue_reg_128(.CP(n_62249), .D(n_41395), .CD(n_60968), .Q(queue
		[128]));
	notech_mux2 i_54772(.S(n_54305), .A(queue[128]), .B(n_42290), .Z(n_41395
		));
	notech_reg queue_reg_129(.CP(n_62249), .D(n_41401), .CD(n_60968), .Q(queue
		[129]));
	notech_mux2 i_54780(.S(n_54305), .A(queue[129]), .B(n_42292), .Z(n_41401
		));
	notech_reg queue_reg_130(.CP(n_62249), .D(n_41407), .CD(n_60967), .Q(queue
		[130]));
	notech_mux2 i_54788(.S(n_54305), .A(queue[130]), .B(n_42294), .Z(n_41407
		));
	notech_reg queue_reg_131(.CP(n_62249), .D(n_41413), .CD(n_60967), .Q(queue
		[131]));
	notech_mux2 i_54796(.S(n_54305), .A(queue[131]), .B(n_42296), .Z(n_41413
		));
	notech_reg queue_reg_132(.CP(n_62249), .D(n_41419), .CD(n_60968), .Q(queue
		[132]));
	notech_mux2 i_54804(.S(n_54305), .A(queue[132]), .B(n_42298), .Z(n_41419
		));
	notech_reg queue_reg_133(.CP(n_62249), .D(n_41425), .CD(n_60968), .Q(queue
		[133]));
	notech_mux2 i_54812(.S(n_54305), .A(queue[133]), .B(n_42300), .Z(n_41425
		));
	notech_reg queue_reg_134(.CP(n_62249), .D(n_41431), .CD(n_60968), .Q(queue
		[134]));
	notech_mux2 i_54820(.S(n_54305), .A(queue[134]), .B(n_42302), .Z(n_41431
		));
	notech_reg queue_reg_135(.CP(n_62249), .D(n_41437), .CD(n_60968), .Q(queue
		[135]));
	notech_mux2 i_54828(.S(n_54305), .A(queue[135]), .B(n_42304), .Z(n_41437
		));
	notech_reg queue_reg_136(.CP(n_62249), .D(n_41443), .CD(n_60968), .Q(queue
		[136]));
	notech_mux2 i_54836(.S(n_54305), .A(queue[136]), .B(n_42306), .Z(n_41443
		));
	notech_reg queue_reg_137(.CP(n_62249), .D(n_41449), .CD(n_60967), .Q(queue
		[137]));
	notech_mux2 i_54844(.S(n_54305), .A(queue[137]), .B(n_42308), .Z(n_41449
		));
	notech_reg queue_reg_138(.CP(n_62249), .D(n_41455), .CD(n_60967), .Q(queue
		[138]));
	notech_mux2 i_54852(.S(n_54305), .A(queue[138]), .B(n_42310), .Z(n_41455
		));
	notech_reg queue_reg_139(.CP(n_62249), .D(n_41461), .CD(n_60967), .Q(queue
		[139]));
	notech_mux2 i_54860(.S(n_54305), .A(queue[139]), .B(n_42312), .Z(n_41461
		));
	notech_nand3 i_21278479(.A(n_60262), .B(n_58379), .C(queue[13]), .Z(n_1218
		));
	notech_reg queue_reg_140(.CP(n_62249), .D(n_41467), .CD(n_60967), .Q(queue
		[140]));
	notech_mux2 i_54868(.S(n_54305), .A(queue[140]), .B(n_42314), .Z(n_41467
		));
	notech_reg queue_reg_141(.CP(n_62249), .D(n_41473), .CD(n_60967), .Q(queue
		[141]));
	notech_mux2 i_54876(.S(n_54305), .A(queue[141]), .B(n_42316), .Z(n_41473
		));
	notech_reg queue_reg_142(.CP(n_62249), .D(n_41479), .CD(n_60967), .Q(queue
		[142]));
	notech_mux2 i_54884(.S(n_54305), .A(queue[142]), .B(n_42318), .Z(n_41479
		));
	notech_and4 i_524984(.A(n_2056), .B(n_2055), .C(n_2050), .D(n_2054), .Z(squeue_497099
		));
	notech_reg queue_reg_143(.CP(n_62175), .D(n_41485), .CD(n_60967), .Q(queue
		[143]));
	notech_mux2 i_54892(.S(n_54305), .A(queue[143]), .B(n_42320), .Z(n_41485
		));
	notech_nand3 i_19478497(.A(n_57935), .B(n_58209), .C(queue[4]), .Z(n_1215
		));
	notech_reg queue_reg_144(.CP(n_62175), .D(n_41491), .CD(n_60967), .Q(queue
		[144]));
	notech_mux2 i_54900(.S(n_54303), .A(queue[144]), .B(n_42322), .Z(n_41491
		));
	notech_reg queue_reg_145(.CP(n_62175), .D(n_41497), .CD(n_60967), .Q(queue
		[145]));
	notech_mux2 i_54908(.S(n_54303), .A(queue[145]), .B(n_42324), .Z(n_41497
		));
	notech_reg queue_reg_146(.CP(n_62175), .D(n_41503), .CD(n_60967), .Q(queue
		[146]));
	notech_mux2 i_54916(.S(n_54303), .A(queue[146]), .B(n_42326), .Z(n_41503
		));
	notech_reg queue_reg_147(.CP(n_62175), .D(n_41509), .CD(n_60967), .Q(queue
		[147]));
	notech_mux2 i_54924(.S(n_54303), .A(queue[147]), .B(n_42328), .Z(n_41509
		));
	notech_reg queue_reg_148(.CP(n_62175), .D(n_41515), .CD(n_60968), .Q(queue
		[148]));
	notech_mux2 i_54932(.S(n_54303), .A(queue[148]), .B(n_42330), .Z(n_41515
		));
	notech_reg queue_reg_149(.CP(n_62175), .D(n_41521), .CD(n_60969), .Q(queue
		[149]));
	notech_mux2 i_54940(.S(n_54303), .A(queue[149]), .B(n_42332), .Z(n_41521
		));
	notech_reg queue_reg_150(.CP(n_62175), .D(n_41527), .CD(n_60969), .Q(queue
		[150]));
	notech_mux2 i_54948(.S(n_54303), .A(queue[150]), .B(n_42334), .Z(n_41527
		));
	notech_reg queue_reg_151(.CP(n_62175), .D(n_41533), .CD(n_60969), .Q(queue
		[151]));
	notech_mux2 i_54956(.S(n_54303), .A(queue[151]), .B(n_42336), .Z(n_41533
		));
	notech_reg queue_reg_152(.CP(n_62175), .D(n_41539), .CD(n_60969), .Q(queue
		[152]));
	notech_mux2 i_54964(.S(n_54303), .A(queue[152]), .B(n_42338), .Z(n_41539
		));
	notech_reg queue_reg_153(.CP(n_62175), .D(n_41545), .CD(n_60969), .Q(queue
		[153]));
	notech_mux2 i_54972(.S(n_54303), .A(queue[153]), .B(n_42340), .Z(n_41545
		));
	notech_reg queue_reg_154(.CP(n_62257), .D(n_41551), .CD(n_60970), .Q(queue
		[154]));
	notech_mux2 i_54980(.S(n_54303), .A(queue[154]), .B(n_42342), .Z(n_41551
		));
	notech_reg queue_reg_155(.CP(clk), .D(n_41557), .CD(n_60970), .Q(queue[
		155]));
	notech_mux2 i_54988(.S(n_54303), .A(queue[155]), .B(n_42344), .Z(n_41557
		));
	notech_reg queue_reg_156(.CP(clk), .D(n_41563), .CD(n_60970), .Q(queue[
		156]));
	notech_mux2 i_54996(.S(n_54303), .A(queue[156]), .B(n_42346), .Z(n_41563
		));
	notech_nand3 i_18178510(.A(n_60262), .B(n_58379), .C(queue[12]), .Z(n_1201
		));
	notech_reg queue_reg_157(.CP(clk), .D(n_41569), .CD(n_60969), .Q(queue[
		157]));
	notech_mux2 i_55004(.S(n_54303), .A(queue[157]), .B(n_42348), .Z(n_41569
		));
	notech_reg queue_reg_158(.CP(clk), .D(n_41575), .CD(n_60970), .Q(queue[
		158]));
	notech_mux2 i_55012(.S(n_54303), .A(queue[158]), .B(n_42350), .Z(n_41575
		));
	notech_reg queue_reg_159(.CP(n_62187), .D(n_41581), .CD(n_60969), .Q(queue
		[159]));
	notech_mux2 i_55020(.S(n_54303), .A(queue[159]), .B(n_42352), .Z(n_41581
		));
	notech_and4 i_424983(.A(n_2042), .B(n_2041), .C(n_2036), .D(n_2040), .Z(squeue_397100
		));
	notech_reg queue_reg_160(.CP(n_62187), .D(n_41587), .CD(n_60968), .Q(queue
		[160]));
	notech_mux2 i_55028(.S(n_54310), .A(queue[160]), .B(n_42354), .Z(n_41587
		));
	notech_nand3 i_16378528(.A(n_57935), .B(n_58206), .C(queue[3]), .Z(n_1198
		));
	notech_reg queue_reg_161(.CP(n_62187), .D(n_41593), .CD(n_60969), .Q(queue
		[161]));
	notech_mux2 i_55036(.S(n_54310), .A(queue[161]), .B(n_42356), .Z(n_41593
		));
	notech_reg queue_reg_162(.CP(n_62187), .D(n_41599), .CD(n_60968), .Q(queue
		[162]));
	notech_mux2 i_55044(.S(n_54310), .A(queue[162]), .B(n_42358), .Z(n_41599
		));
	notech_reg queue_reg_163(.CP(n_62187), .D(n_41605), .CD(n_60968), .Q(queue
		[163]));
	notech_mux2 i_55052(.S(n_54310), .A(queue[163]), .B(n_42360), .Z(n_41605
		));
	notech_reg queue_reg_164(.CP(n_62187), .D(n_41611), .CD(n_60968), .Q(queue
		[164]));
	notech_mux2 i_55060(.S(n_54310), .A(queue[164]), .B(n_42362), .Z(n_41611
		));
	notech_reg queue_reg_165(.CP(n_62187), .D(n_41617), .CD(n_60969), .Q(queue
		[165]));
	notech_mux2 i_55068(.S(n_54310), .A(queue[165]), .B(n_42364), .Z(n_41617
		));
	notech_reg queue_reg_166(.CP(n_62187), .D(n_41623), .CD(n_60969), .Q(queue
		[166]));
	notech_mux2 i_55076(.S(n_54310), .A(queue[166]), .B(n_42366), .Z(n_41623
		));
	notech_reg queue_reg_167(.CP(n_62187), .D(n_41629), .CD(n_60969), .Q(queue
		[167]));
	notech_mux2 i_55084(.S(n_54310), .A(queue[167]), .B(n_42368), .Z(n_41629
		));
	notech_reg queue_reg_168(.CP(n_62187), .D(n_41635), .CD(n_60969), .Q(queue
		[168]));
	notech_mux2 i_55092(.S(n_54310), .A(queue[168]), .B(n_42370), .Z(n_41635
		));
	notech_reg queue_reg_169(.CP(n_62187), .D(n_41641), .CD(n_60969), .Q(queue
		[169]));
	notech_mux2 i_55100(.S(n_54310), .A(queue[169]), .B(n_42372), .Z(n_41641
		));
	notech_reg queue_reg_170(.CP(n_62187), .D(n_41647), .CD(n_60979), .Q(queue
		[170]));
	notech_mux2 i_55108(.S(n_54310), .A(queue[170]), .B(n_42374), .Z(n_41647
		));
	notech_reg queue_reg_171(.CP(n_62187), .D(n_41653), .CD(n_60979), .Q(queue
		[171]));
	notech_mux2 i_55116(.S(n_54310), .A(queue[171]), .B(n_42376), .Z(n_41653
		));
	notech_reg queue_reg_172(.CP(n_62187), .D(n_41659), .CD(n_60979), .Q(queue
		[172]));
	notech_mux2 i_55124(.S(n_54310), .A(queue[172]), .B(n_42378), .Z(n_41659
		));
	notech_reg queue_reg_173(.CP(n_62187), .D(n_41665), .CD(n_60979), .Q(queue
		[173]));
	notech_mux2 i_55132(.S(n_54310), .A(queue[173]), .B(n_42380), .Z(n_41665
		));
	notech_nand3 i_15078541(.A(n_60262), .B(n_58379), .C(queue[11]), .Z(n_1185
		));
	notech_reg queue_reg_174(.CP(n_62187), .D(n_41671), .CD(n_60979), .Q(queue
		[174]));
	notech_mux2 i_55140(.S(n_54310), .A(queue[174]), .B(n_42382), .Z(n_41671
		));
	notech_reg queue_reg_175(.CP(n_62187), .D(n_41677), .CD(n_60979), .Q(queue
		[175]));
	notech_mux2 i_55148(.S(n_54310), .A(queue[175]), .B(n_42384), .Z(n_41677
		));
	notech_reg queue_reg_176(.CP(n_62187), .D(n_41683), .CD(n_60980), .Q(queue
		[176]));
	notech_mux2 i_55156(.S(n_54308), .A(queue[176]), .B(n_42386), .Z(n_41683
		));
	notech_and4 i_324982(.A(n_2028), .B(n_2027), .C(n_2022), .D(n_2026), .Z(squeue_297101
		));
	notech_reg queue_reg_177(.CP(n_62187), .D(n_41689), .CD(n_60979), .Q(queue
		[177]));
	notech_mux2 i_55164(.S(n_54308), .A(queue[177]), .B(n_42388), .Z(n_41689
		));
	notech_nand3 i_13278559(.A(n_57935), .B(n_58206), .C(queue[2]), .Z(n_1182
		));
	notech_reg queue_reg_178(.CP(n_62261), .D(n_41695), .CD(n_60979), .Q(queue
		[178]));
	notech_mux2 i_55172(.S(n_54308), .A(queue[178]), .B(n_42390), .Z(n_41695
		));
	notech_reg queue_reg_179(.CP(n_62185), .D(n_41701), .CD(n_60979), .Q(queue
		[179]));
	notech_mux2 i_55180(.S(n_54308), .A(queue[179]), .B(n_42392), .Z(n_41701
		));
	notech_reg queue_reg_180(.CP(n_62261), .D(n_41707), .CD(n_60979), .Q(queue
		[180]));
	notech_mux2 i_55188(.S(n_54308), .A(queue[180]), .B(n_42394), .Z(n_41707
		));
	notech_reg queue_reg_181(.CP(n_62261), .D(n_41713), .CD(n_60977), .Q(queue
		[181]));
	notech_mux2 i_55196(.S(n_54308), .A(queue[181]), .B(n_42396), .Z(n_41713
		));
	notech_reg queue_reg_182(.CP(n_62261), .D(n_41719), .CD(n_60977), .Q(queue
		[182]));
	notech_mux2 i_55204(.S(n_54308), .A(queue[182]), .B(n_42398), .Z(n_41719
		));
	notech_reg queue_reg_183(.CP(n_62261), .D(n_41725), .CD(n_60977), .Q(queue
		[183]));
	notech_mux2 i_55212(.S(n_54308), .A(queue[183]), .B(n_42400), .Z(n_41725
		));
	notech_reg queue_reg_184(.CP(n_62261), .D(n_41731), .CD(n_60977), .Q(queue
		[184]));
	notech_mux2 i_55220(.S(n_54308), .A(queue[184]), .B(n_42402), .Z(n_41731
		));
	notech_reg queue_reg_185(.CP(n_62261), .D(n_41737), .CD(n_60977), .Q(queue
		[185]));
	notech_mux2 i_55228(.S(n_54308), .A(queue[185]), .B(n_42404), .Z(n_41737
		));
	notech_reg queue_reg_186(.CP(n_62261), .D(n_41743), .CD(n_60979), .Q(queue
		[186]));
	notech_mux2 i_55236(.S(n_54308), .A(queue[186]), .B(n_42406), .Z(n_41743
		));
	notech_reg queue_reg_187(.CP(n_62261), .D(n_41749), .CD(n_60979), .Q(queue
		[187]));
	notech_mux2 i_55244(.S(n_54308), .A(queue[187]), .B(n_42408), .Z(n_41749
		));
	notech_reg queue_reg_188(.CP(n_62261), .D(n_41755), .CD(n_60979), .Q(queue
		[188]));
	notech_mux2 i_55252(.S(n_54308), .A(queue[188]), .B(n_42410), .Z(n_41755
		));
	notech_reg queue_reg_189(.CP(n_62261), .D(n_41761), .CD(n_60977), .Q(queue
		[189]));
	notech_mux2 i_55260(.S(n_54308), .A(queue[189]), .B(n_42412), .Z(n_41761
		));
	notech_reg queue_reg_190(.CP(n_62261), .D(n_41767), .CD(n_60979), .Q(queue
		[190]));
	notech_mux2 i_55268(.S(n_54308), .A(queue[190]), .B(n_42414), .Z(n_41767
		));
	notech_nand3 i_11978572(.A(n_60262), .B(n_58379), .C(queue[10]), .Z(n_1169
		));
	notech_reg queue_reg_191(.CP(n_62261), .D(n_41773), .CD(n_60980), .Q(queue
		[191]));
	notech_mux2 i_55276(.S(n_54308), .A(queue[191]), .B(n_42416), .Z(n_41773
		));
	notech_reg queue_reg_192(.CP(n_62261), .D(n_41779), .CD(n_60981), .Q(queue
		[192]));
	notech_mux2 i_55284(.S(n_54295), .A(queue[192]), .B(n_42418), .Z(n_41779
		));
	notech_reg queue_reg_193(.CP(n_62261), .D(n_41785), .CD(n_60981), .Q(queue
		[193]));
	notech_mux2 i_55292(.S(n_54295), .A(queue[193]), .B(n_42420), .Z(n_41785
		));
	notech_and4 i_224981(.A(n_2014), .B(n_2013), .C(n_2008), .D(n_2012), .Z(squeue_197102
		));
	notech_reg queue_reg_194(.CP(n_62261), .D(n_41791), .CD(n_60981), .Q(queue
		[194]));
	notech_mux2 i_55300(.S(n_54295), .A(queue[194]), .B(n_42422), .Z(n_41791
		));
	notech_nand3 i_10178590(.A(n_57935), .B(n_58209), .C(queue[1]), .Z(n_1166
		));
	notech_reg queue_reg_195(.CP(n_62261), .D(n_41797), .CD(n_60980), .Q(queue
		[195]));
	notech_mux2 i_55308(.S(n_54295), .A(queue[195]), .B(n_42424), .Z(n_41797
		));
	notech_reg queue_reg_196(.CP(n_62261), .D(n_41803), .CD(n_60981), .Q(queue
		[196]));
	notech_mux2 i_55316(.S(n_54295), .A(queue[196]), .B(n_42426), .Z(n_41803
		));
	notech_reg queue_reg_197(.CP(n_62261), .D(n_41809), .CD(n_60981), .Q(queue
		[197]));
	notech_mux2 i_55324(.S(n_54295), .A(queue[197]), .B(n_42428), .Z(n_41809
		));
	notech_reg queue_reg_198(.CP(n_62185), .D(n_41815), .CD(n_60981), .Q(queue
		[198]));
	notech_mux2 i_55332(.S(n_54295), .A(queue[198]), .B(n_42430), .Z(n_41815
		));
	notech_reg queue_reg_199(.CP(n_62185), .D(n_41821), .CD(n_60981), .Q(queue
		[199]));
	notech_mux2 i_55340(.S(n_54295), .A(queue[199]), .B(n_42432), .Z(n_41821
		));
	notech_reg queue_reg_200(.CP(n_62185), .D(n_41827), .CD(n_60981), .Q(queue
		[200]));
	notech_mux2 i_55348(.S(n_54295), .A(queue[200]), .B(n_42434), .Z(n_41827
		));
	notech_reg queue_reg_201(.CP(n_62185), .D(n_41833), .CD(n_60981), .Q(queue
		[201]));
	notech_mux2 i_55356(.S(n_54295), .A(queue[201]), .B(n_42436), .Z(n_41833
		));
	notech_reg queue_reg_202(.CP(n_62185), .D(n_41839), .CD(n_60980), .Q(queue
		[202]));
	notech_mux2 i_55364(.S(n_54295), .A(queue[202]), .B(n_42438), .Z(n_41839
		));
	notech_reg queue_reg_203(.CP(n_62185), .D(n_41845), .CD(n_60980), .Q(queue
		[203]));
	notech_mux2 i_55372(.S(n_54295), .A(queue[203]), .B(n_42440), .Z(n_41845
		));
	notech_reg queue_reg_204(.CP(clk), .D(n_41851), .CD(n_60980), .Q(queue[
		204]));
	notech_mux2 i_55380(.S(n_54295), .A(queue[204]), .B(n_42442), .Z(n_41851
		));
	notech_reg queue_reg_205(.CP(n_62183), .D(n_41857), .CD(n_60980), .Q(queue
		[205]));
	notech_mux2 i_55388(.S(n_54295), .A(queue[205]), .B(n_42444), .Z(n_41857
		));
	notech_reg queue_reg_206(.CP(n_62257), .D(n_41863), .CD(n_60980), .Q(queue
		[206]));
	notech_mux2 i_55396(.S(n_54295), .A(queue[206]), .B(n_42446), .Z(n_41863
		));
	notech_reg queue_reg_207(.CP(n_62257), .D(n_41869), .CD(n_60980), .Q(queue
		[207]));
	notech_mux2 i_55404(.S(n_54295), .A(queue[207]), .B(n_42448), .Z(n_41869
		));
	notech_nand3 i_8878603(.A(n_60262), .B(n_58379), .C(queue[9]), .Z(n_1153
		));
	notech_reg queue_reg_208(.CP(n_62257), .D(n_41875), .CD(n_60980), .Q(queue
		[208]));
	notech_mux2 i_55412(.S(n_54293), .A(queue[208]), .B(n_42450), .Z(n_41875
		));
	notech_reg queue_reg_209(.CP(n_62257), .D(n_41881), .CD(n_60980), .Q(queue
		[209]));
	notech_mux2 i_55420(.S(n_54293), .A(queue[209]), .B(n_42452), .Z(n_41881
		));
	notech_reg queue_reg_210(.CP(n_62257), .D(n_41887), .CD(n_60980), .Q(queue
		[210]));
	notech_mux2 i_55428(.S(n_54293), .A(queue[210]), .B(n_42454), .Z(n_41887
		));
	notech_and4 i_124980(.A(n_2000), .B(n_1997), .C(n_1986), .D(n_1994), .Z(squeue_097103
		));
	notech_reg queue_reg_211(.CP(n_62333), .D(n_41893), .CD(n_60980), .Q(queue
		[211]));
	notech_mux2 i_55436(.S(n_54293), .A(queue[211]), .B(n_42456), .Z(n_41893
		));
	notech_nand3 i_6678621(.A(n_57935), .B(n_58209), .C(queue[0]), .Z(n_1150
		));
	notech_reg queue_reg_212(.CP(n_62333), .D(n_41899), .CD(n_60980), .Q(queue
		[212]));
	notech_mux2 i_55444(.S(n_54293), .A(queue[212]), .B(n_42458), .Z(n_41899
		));
	notech_reg queue_reg_213(.CP(n_62333), .D(n_41905), .CD(n_60975), .Q(queue
		[213]));
	notech_mux2 i_55452(.S(n_54293), .A(queue[213]), .B(n_42460), .Z(n_41905
		));
	notech_reg queue_reg_214(.CP(n_62333), .D(n_41911), .CD(n_60975), .Q(queue
		[214]));
	notech_mux2 i_55460(.S(n_54293), .A(queue[214]), .B(n_42462), .Z(n_41911
		));
	notech_reg queue_reg_215(.CP(n_62333), .D(n_41917), .CD(n_60975), .Q(queue
		[215]));
	notech_mux2 i_55468(.S(n_54293), .A(queue[215]), .B(n_42464), .Z(n_41917
		));
	notech_reg queue_reg_216(.CP(n_62333), .D(n_41923), .CD(n_60975), .Q(queue
		[216]));
	notech_mux2 i_55476(.S(n_54293), .A(queue[216]), .B(n_42466), .Z(n_41923
		));
	notech_reg queue_reg_217(.CP(n_62333), .D(n_41929), .CD(n_60975), .Q(queue
		[217]));
	notech_mux2 i_55484(.S(n_54293), .A(queue[217]), .B(n_42468), .Z(n_41929
		));
	notech_reg queue_reg_218(.CP(n_62333), .D(n_41935), .CD(n_60975), .Q(queue
		[218]));
	notech_mux2 i_55492(.S(n_54293), .A(queue[218]), .B(n_42470), .Z(n_41935
		));
	notech_reg queue_reg_219(.CP(n_62333), .D(n_41941), .CD(n_60975), .Q(queue
		[219]));
	notech_mux2 i_55500(.S(n_54293), .A(queue[219]), .B(n_42472), .Z(n_41941
		));
	notech_reg queue_reg_220(.CP(n_62333), .D(n_41947), .CD(n_60975), .Q(queue
		[220]));
	notech_mux2 i_55508(.S(n_54293), .A(queue[220]), .B(n_42474), .Z(n_41947
		));
	notech_reg queue_reg_221(.CP(n_62333), .D(n_41953), .CD(n_60975), .Q(queue
		[221]));
	notech_mux2 i_55516(.S(n_54293), .A(queue[221]), .B(n_42476), .Z(n_41953
		));
	notech_reg queue_reg_222(.CP(n_62333), .D(n_41959), .CD(n_60975), .Q(queue
		[222]));
	notech_mux2 i_55524(.S(n_54293), .A(queue[222]), .B(n_42478), .Z(n_41959
		));
	notech_reg queue_reg_223(.CP(n_62333), .D(n_41965), .CD(n_60975), .Q(queue
		[223]));
	notech_mux2 i_55532(.S(n_54293), .A(queue[223]), .B(n_42480), .Z(n_41965
		));
	notech_reg queue_reg_224(.CP(n_62333), .D(n_41971), .CD(n_60974), .Q(queue
		[224]));
	notech_mux2 i_55540(.S(n_54300), .A(queue[224]), .B(n_42482), .Z(n_41971
		));
	notech_nand3 i_5278634(.A(n_60262), .B(n_58379), .C(queue[8]), .Z(n_113293395
		));
	notech_reg queue_reg_225(.CP(n_62333), .D(n_41977), .CD(n_60974), .Q(queue
		[225]));
	notech_mux2 i_55548(.S(n_54300), .A(queue[225]), .B(n_42484), .Z(n_41977
		));
	notech_reg queue_reg_226(.CP(n_62333), .D(n_41983), .CD(n_60974), .Q(queue
		[226]));
	notech_mux2 i_55556(.S(n_54300), .A(queue[226]), .B(n_42486), .Z(n_41983
		));
	notech_reg queue_reg_227(.CP(n_62333), .D(n_41989), .CD(n_60974), .Q(queue
		[227]));
	notech_mux2 i_55564(.S(n_54300), .A(queue[227]), .B(n_42488), .Z(n_41989
		));
	notech_reg queue_reg_228(.CP(n_62333), .D(n_41995), .CD(n_60974), .Q(queue
		[228]));
	notech_mux2 i_55572(.S(n_54300), .A(queue[228]), .B(n_42490), .Z(n_41995
		));
	notech_reg queue_reg_229(.CP(n_62257), .D(n_42001), .CD(n_60975), .Q(queue
		[229]));
	notech_mux2 i_55580(.S(n_54300), .A(queue[229]), .B(n_42492), .Z(n_42001
		));
	notech_nand3 i_44778776(.A(addrshft[3]), .B(n_42548), .C(n_42549), .Z(n_112793393
		));
	notech_reg queue_reg_230(.CP(n_62333), .D(n_42007), .CD(n_60975), .Q(queue
		[230]));
	notech_mux2 i_55588(.S(n_54300), .A(queue[230]), .B(n_42494), .Z(n_42007
		));
	notech_nor2 i_3131103(.A(addrshft[0]), .B(addrshft[1]), .Z(n_1126));
	notech_reg queue_reg_231(.CP(n_62259), .D(n_42013), .CD(n_60975), .Q(queue
		[231]));
	notech_mux2 i_55596(.S(n_54300), .A(queue[231]), .B(n_42496), .Z(n_42013
		));
	notech_or2 i_44878775(.A(addrshft[0]), .B(n_42548), .Z(n_112593392));
	notech_reg queue_reg_232(.CP(n_62259), .D(n_42019), .CD(n_60974), .Q(queue
		[232]));
	notech_mux2 i_55604(.S(n_54300), .A(queue[232]), .B(n_42498), .Z(n_42019
		));
	notech_nand3 i_6179187(.A(wptr[0]), .B(n_3062), .C(n_42170), .Z(n_112493391
		));
	notech_reg queue_reg_233(.CP(n_62259), .D(n_42025), .CD(n_60974), .Q(queue
		[233]));
	notech_mux2 i_55612(.S(n_54300), .A(queue[233]), .B(n_42500), .Z(n_42025
		));
	notech_reg queue_reg_234(.CP(n_62259), .D(n_42031), .CD(n_60976), .Q(queue
		[234]));
	notech_mux2 i_55620(.S(n_54300), .A(queue[234]), .B(n_42502), .Z(n_42031
		));
	notech_reg queue_reg_235(.CP(n_62259), .D(n_42037), .CD(n_60977), .Q(queue
		[235]));
	notech_mux2 i_55628(.S(n_54300), .A(queue[235]), .B(n_42504), .Z(n_42037
		));
	notech_ao4 i_3479184(.A(wptr[0]), .B(n_42170), .C(n_112493391), .D(n_42547
		), .Z(n_1119));
	notech_reg queue_reg_236(.CP(n_62259), .D(n_42043), .CD(n_60977), .Q(queue
		[236]));
	notech_mux2 i_55636(.S(n_54300), .A(queue[236]), .B(n_42506), .Z(n_42043
		));
	notech_reg queue_reg_237(.CP(n_62259), .D(n_42049), .CD(n_60977), .Q(queue
		[237]));
	notech_mux2 i_55644(.S(n_54300), .A(queue[237]), .B(n_42508), .Z(n_42049
		));
	notech_reg queue_reg_238(.CP(n_62259), .D(n_42055), .CD(n_60976), .Q(queue
		[238]));
	notech_mux2 i_55652(.S(n_54300), .A(queue[238]), .B(n_42510), .Z(n_42055
		));
	notech_reg queue_reg_239(.CP(n_62259), .D(n_42061), .CD(n_60976), .Q(queue
		[239]));
	notech_mux2 i_55660(.S(n_54300), .A(queue[239]), .B(n_42512), .Z(n_42061
		));
	notech_reg queue_reg_240(.CP(n_62259), .D(n_42067), .CD(n_60977), .Q(queue
		[240]));
	notech_mux2 i_55668(.S(n_54298), .A(queue[240]), .B(n_42514), .Z(n_42067
		));
	notech_reg queue_reg_241(.CP(n_62259), .D(n_42073), .CD(n_60977), .Q(queue
		[241]));
	notech_mux2 i_55676(.S(n_54298), .A(queue[241]), .B(n_42516), .Z(n_42073
		));
	notech_xor2 i_3779181(.A(n_1126), .B(addrshft[2]), .Z(n_1112));
	notech_reg queue_reg_242(.CP(n_62259), .D(n_42079), .CD(n_60977), .Q(queue
		[242]));
	notech_mux2 i_55684(.S(n_54298), .A(queue[242]), .B(n_42518), .Z(n_42079
		));
	notech_reg queue_reg_243(.CP(n_62259), .D(n_42085), .CD(n_60977), .Q(queue
		[243]));
	notech_mux2 i_55692(.S(n_54298), .A(queue[243]), .B(n_42520), .Z(n_42085
		));
	notech_reg queue_reg_244(.CP(n_62259), .D(n_42091), .CD(n_60977), .Q(queue
		[244]));
	notech_mux2 i_55700(.S(n_54298), .A(queue[244]), .B(n_42522), .Z(n_42091
		));
	notech_reg queue_reg_245(.CP(n_62259), .D(n_42097), .CD(n_60976), .Q(queue
		[245]));
	notech_mux2 i_55708(.S(n_54298), .A(queue[245]), .B(n_42524), .Z(n_42097
		));
	notech_reg queue_reg_246(.CP(n_62259), .D(n_42103), .CD(n_60976), .Q(queue
		[246]));
	notech_mux2 i_55716(.S(n_54298), .A(queue[246]), .B(n_42526), .Z(n_42103
		));
	notech_ao4 i_3879180(.A(n_60262), .B(addrshft[3]), .C(addrshft[0]), .D(n_112793393
		), .Z(n_1107));
	notech_reg queue_reg_247(.CP(n_62259), .D(n_42109), .CD(n_60976), .Q(queue
		[247]));
	notech_mux2 i_55724(.S(n_54298), .A(queue[247]), .B(n_42528), .Z(n_42109
		));
	notech_reg queue_reg_248(.CP(n_62259), .D(n_42115), .CD(n_60976), .Q(queue
		[248]));
	notech_mux2 i_55732(.S(n_54298), .A(queue[248]), .B(n_42530), .Z(n_42115
		));
	notech_reg queue_reg_249(.CP(n_62259), .D(n_42121), .CD(n_60976), .Q(queue
		[249]));
	notech_mux2 i_55740(.S(n_54298), .A(queue[249]), .B(n_42532), .Z(n_42121
		));
	notech_reg queue_reg_250(.CP(n_62183), .D(n_42127), .CD(n_60976), .Q(queue
		[250]));
	notech_mux2 i_55748(.S(n_54298), .A(queue[250]), .B(n_42534), .Z(n_42127
		));
	notech_reg queue_reg_251(.CP(n_62183), .D(n_42133), .CD(n_60976), .Q(queue
		[251]));
	notech_mux2 i_55756(.S(n_54298), .A(queue[251]), .B(n_42536), .Z(n_42133
		));
	notech_reg queue_reg_252(.CP(n_62183), .D(n_42139), .CD(n_60976), .Q(queue
		[252]));
	notech_mux2 i_55764(.S(n_54298), .A(queue[252]), .B(n_42538), .Z(n_42139
		));
	notech_reg queue_reg_253(.CP(n_62183), .D(n_42145), .CD(n_60976), .Q(queue
		[253]));
	notech_mux2 i_55772(.S(n_54298), .A(queue[253]), .B(n_42540), .Z(n_42145
		));
	notech_reg queue_reg_254(.CP(clk), .D(n_42151), .CD(n_60976), .Q(queue[
		254]));
	notech_mux2 i_55780(.S(n_54298), .A(queue[254]), .B(n_42542), .Z(n_42151
		));
	notech_reg queue_reg_255(.CP(n_62183), .D(n_42157), .CD(n_60976), .Q(queue
		[255]));
	notech_mux2 i_55788(.S(n_54298), .A(queue[255]), .B(n_42544), .Z(n_42157
		));
	notech_inv i_58839(.A(n_7790), .Z(n_42163));
	notech_inv i_58840(.A(n_8288), .Z(n_42164));
	notech_inv i_58841(.A(n_3855342), .Z(n_42165));
	notech_inv i_58843(.A(n_309596466), .Z(n_42167));
	notech_inv i_58844(.A(n_8293), .Z(n_42168));
	notech_inv i_58845(.A(wptr[0]), .Z(n_42169));
	notech_inv i_58846(.A(n_60277), .Z(n_42170));
	notech_inv i_58847(.A(\nbus_12114[0] ), .Z(n_42171));
	notech_inv i_58848(.A(n_35031), .Z(n_42172));
	notech_inv i_58849(.A(n_35037), .Z(n_42173));
	notech_inv i_58850(.A(n_35044), .Z(n_42174));
	notech_inv i_58851(.A(purge), .Z(cacheD[148]));
	notech_inv i_58852(.A(queue[15]), .Z(n_42176));
	notech_inv i_58853(.A(queue[16]), .Z(n_42177));
	notech_inv i_58854(.A(queue[17]), .Z(n_42178));
	notech_inv i_58855(.A(queue[18]), .Z(n_42179));
	notech_inv i_58856(.A(queue[19]), .Z(n_42180));
	notech_inv i_58857(.A(queue[20]), .Z(n_42181));
	notech_inv i_58858(.A(queue[21]), .Z(n_42182));
	notech_inv i_58859(.A(queue[22]), .Z(n_42183));
	notech_inv i_58860(.A(queue[23]), .Z(n_42184));
	notech_inv i_58861(.A(queue[24]), .Z(n_42185));
	notech_inv i_58862(.A(queue[25]), .Z(n_42186));
	notech_inv i_58863(.A(queue[26]), .Z(n_42187));
	notech_inv i_58864(.A(queue[27]), .Z(n_42188));
	notech_inv i_58865(.A(queue[28]), .Z(n_42189));
	notech_inv i_58866(.A(queue[29]), .Z(n_42190));
	notech_inv i_58867(.A(queue[30]), .Z(n_42191));
	notech_inv i_58868(.A(queue[31]), .Z(n_42192));
	notech_inv i_58869(.A(queue[32]), .Z(n_42193));
	notech_inv i_58870(.A(queue[33]), .Z(n_42194));
	notech_inv i_58871(.A(queue[34]), .Z(n_42195));
	notech_inv i_58872(.A(queue[35]), .Z(n_42196));
	notech_inv i_58873(.A(queue[36]), .Z(n_42197));
	notech_inv i_58874(.A(queue[37]), .Z(n_42198));
	notech_inv i_58875(.A(queue[38]), .Z(n_42199));
	notech_inv i_58876(.A(queue[39]), .Z(n_42200));
	notech_inv i_58877(.A(queue[40]), .Z(n_42201));
	notech_inv i_58878(.A(queue[41]), .Z(n_42202));
	notech_inv i_58879(.A(queue[42]), .Z(n_42203));
	notech_inv i_58880(.A(queue[43]), .Z(n_42204));
	notech_inv i_58881(.A(queue[44]), .Z(n_42205));
	notech_inv i_58882(.A(queue[45]), .Z(n_42206));
	notech_inv i_58883(.A(queue[46]), .Z(n_42207));
	notech_inv i_58884(.A(queue[47]), .Z(n_42208));
	notech_inv i_58885(.A(queue[48]), .Z(n_42209));
	notech_inv i_58886(.A(queue[49]), .Z(n_42210));
	notech_inv i_58887(.A(queue[50]), .Z(n_42211));
	notech_inv i_58888(.A(queue[51]), .Z(n_42212));
	notech_inv i_58889(.A(queue[52]), .Z(n_42213));
	notech_inv i_58890(.A(queue[53]), .Z(n_42214));
	notech_inv i_58891(.A(queue[54]), .Z(n_42215));
	notech_inv i_58892(.A(queue[55]), .Z(n_42216));
	notech_inv i_58893(.A(queue[56]), .Z(n_42217));
	notech_inv i_58894(.A(queue[57]), .Z(n_42218));
	notech_inv i_58895(.A(queue[58]), .Z(n_42219));
	notech_inv i_58896(.A(queue[59]), .Z(n_42220));
	notech_inv i_58897(.A(queue[60]), .Z(n_42221));
	notech_inv i_58898(.A(queue[61]), .Z(n_42222));
	notech_inv i_58899(.A(queue[62]), .Z(n_42223));
	notech_inv i_58900(.A(queue[63]), .Z(n_42224));
	notech_inv i_58901(.A(queue[64]), .Z(n_42225));
	notech_inv i_58902(.A(queue[65]), .Z(n_42226));
	notech_inv i_58903(.A(queue[66]), .Z(n_42227));
	notech_inv i_58904(.A(queue[67]), .Z(n_42228));
	notech_inv i_58905(.A(queue[68]), .Z(n_42229));
	notech_inv i_58906(.A(queue[69]), .Z(n_42230));
	notech_inv i_58907(.A(queue[70]), .Z(n_42231));
	notech_inv i_58908(.A(queue[71]), .Z(n_42232));
	notech_inv i_58909(.A(queue[72]), .Z(n_42233));
	notech_inv i_58910(.A(queue[73]), .Z(n_42234));
	notech_inv i_58911(.A(queue[74]), .Z(n_42235));
	notech_inv i_58912(.A(queue[75]), .Z(n_42236));
	notech_inv i_58913(.A(queue[76]), .Z(n_42237));
	notech_inv i_58914(.A(queue[77]), .Z(n_42238));
	notech_inv i_58915(.A(queue[78]), .Z(n_42239));
	notech_inv i_58916(.A(queue[79]), .Z(n_42240));
	notech_inv i_58917(.A(queue[80]), .Z(n_42241));
	notech_inv i_58918(.A(queue[81]), .Z(n_42242));
	notech_inv i_58919(.A(queue[82]), .Z(n_42243));
	notech_inv i_58920(.A(queue[83]), .Z(n_42244));
	notech_inv i_58921(.A(queue[84]), .Z(n_42245));
	notech_inv i_58922(.A(queue[85]), .Z(n_42246));
	notech_inv i_58923(.A(queue[86]), .Z(n_42247));
	notech_inv i_58924(.A(queue[87]), .Z(n_42248));
	notech_inv i_58925(.A(queue[88]), .Z(n_42249));
	notech_inv i_58926(.A(queue[89]), .Z(n_42250));
	notech_inv i_58927(.A(queue[90]), .Z(n_42251));
	notech_inv i_58928(.A(queue[91]), .Z(n_42252));
	notech_inv i_58929(.A(queue[92]), .Z(n_42253));
	notech_inv i_58930(.A(queue[93]), .Z(n_42254));
	notech_inv i_58931(.A(queue[94]), .Z(n_42255));
	notech_inv i_58932(.A(queue[95]), .Z(n_42256));
	notech_inv i_58933(.A(queue[96]), .Z(n_42257));
	notech_inv i_58934(.A(queue[97]), .Z(n_42258));
	notech_inv i_58935(.A(queue[98]), .Z(n_42259));
	notech_inv i_58936(.A(queue[99]), .Z(n_42260));
	notech_inv i_58937(.A(queue[100]), .Z(n_42261));
	notech_inv i_58938(.A(queue[101]), .Z(n_42262));
	notech_inv i_58939(.A(queue[102]), .Z(n_42263));
	notech_inv i_58940(.A(queue[103]), .Z(n_42264));
	notech_inv i_58941(.A(queue[104]), .Z(n_42265));
	notech_inv i_58942(.A(queue[105]), .Z(n_42266));
	notech_inv i_58943(.A(queue[106]), .Z(n_42267));
	notech_inv i_58944(.A(queue[107]), .Z(n_42268));
	notech_inv i_58945(.A(queue[108]), .Z(n_42269));
	notech_inv i_58946(.A(queue[109]), .Z(n_42270));
	notech_inv i_58947(.A(queue[110]), .Z(n_42271));
	notech_inv i_58948(.A(queue[111]), .Z(n_42272));
	notech_inv i_58949(.A(queue[112]), .Z(n_42273));
	notech_inv i_58950(.A(queue[113]), .Z(n_42274));
	notech_inv i_58951(.A(queue[114]), .Z(n_42275));
	notech_inv i_58952(.A(queue[115]), .Z(n_42276));
	notech_inv i_58953(.A(queue[116]), .Z(n_42277));
	notech_inv i_58954(.A(queue[117]), .Z(n_42278));
	notech_inv i_58955(.A(queue[118]), .Z(n_42279));
	notech_inv i_58956(.A(queue[119]), .Z(n_42280));
	notech_inv i_58957(.A(queue[120]), .Z(n_42281));
	notech_inv i_58958(.A(queue[121]), .Z(n_42282));
	notech_inv i_58959(.A(queue[122]), .Z(n_42283));
	notech_inv i_58960(.A(queue[123]), .Z(n_42284));
	notech_inv i_58961(.A(queue[124]), .Z(n_42285));
	notech_inv i_58962(.A(queue[125]), .Z(n_42286));
	notech_inv i_58963(.A(queue[126]), .Z(n_42287));
	notech_inv i_58964(.A(queue[127]), .Z(n_42288));
	notech_inv i_58966(.A(n_35843), .Z(n_42290));
	notech_inv i_58967(.A(queue[128]), .Z(n_42291));
	notech_inv i_58968(.A(n_35849), .Z(n_42292));
	notech_inv i_58969(.A(queue[129]), .Z(n_42293));
	notech_inv i_58970(.A(n_35855), .Z(n_42294));
	notech_inv i_58971(.A(queue[130]), .Z(n_42295));
	notech_inv i_58972(.A(n_35861), .Z(n_42296));
	notech_inv i_58973(.A(queue[131]), .Z(n_42297));
	notech_inv i_58974(.A(n_35867), .Z(n_42298));
	notech_inv i_58975(.A(queue[132]), .Z(n_42299));
	notech_inv i_58976(.A(n_35873), .Z(n_42300));
	notech_inv i_58977(.A(queue[133]), .Z(n_42301));
	notech_inv i_58978(.A(n_35879), .Z(n_42302));
	notech_inv i_58979(.A(queue[134]), .Z(n_42303));
	notech_inv i_58980(.A(n_35885), .Z(n_42304));
	notech_inv i_58981(.A(queue[135]), .Z(n_42305));
	notech_inv i_58982(.A(n_35891), .Z(n_42306));
	notech_inv i_58983(.A(queue[136]), .Z(n_42307));
	notech_inv i_58984(.A(n_35897), .Z(n_42308));
	notech_inv i_58985(.A(queue[137]), .Z(n_42309));
	notech_inv i_58986(.A(n_35903), .Z(n_42310));
	notech_inv i_58987(.A(queue[138]), .Z(n_42311));
	notech_inv i_58988(.A(n_35909), .Z(n_42312));
	notech_inv i_58989(.A(queue[139]), .Z(n_42313));
	notech_inv i_58990(.A(n_35915), .Z(n_42314));
	notech_inv i_58991(.A(queue[140]), .Z(n_42315));
	notech_inv i_58992(.A(n_35921), .Z(n_42316));
	notech_inv i_58993(.A(queue[141]), .Z(n_42317));
	notech_inv i_58994(.A(n_35927), .Z(n_42318));
	notech_inv i_58995(.A(queue[142]), .Z(n_42319));
	notech_inv i_58996(.A(n_35933), .Z(n_42320));
	notech_inv i_58997(.A(queue[143]), .Z(n_42321));
	notech_inv i_58998(.A(n_35939), .Z(n_42322));
	notech_inv i_58999(.A(queue[144]), .Z(n_42323));
	notech_inv i_59000(.A(n_35945), .Z(n_42324));
	notech_inv i_59001(.A(queue[145]), .Z(n_42325));
	notech_inv i_59002(.A(n_35951), .Z(n_42326));
	notech_inv i_59003(.A(queue[146]), .Z(n_42327));
	notech_inv i_59004(.A(n_35957), .Z(n_42328));
	notech_inv i_59005(.A(queue[147]), .Z(n_42329));
	notech_inv i_59006(.A(n_35963), .Z(n_42330));
	notech_inv i_59007(.A(queue[148]), .Z(n_42331));
	notech_inv i_59008(.A(n_35969), .Z(n_42332));
	notech_inv i_59009(.A(queue[149]), .Z(n_42333));
	notech_inv i_59010(.A(n_35975), .Z(n_42334));
	notech_inv i_59011(.A(queue[150]), .Z(n_42335));
	notech_inv i_59012(.A(n_35981), .Z(n_42336));
	notech_inv i_59013(.A(queue[151]), .Z(n_42337));
	notech_inv i_59014(.A(n_35987), .Z(n_42338));
	notech_inv i_59015(.A(queue[152]), .Z(n_42339));
	notech_inv i_59016(.A(n_35993), .Z(n_42340));
	notech_inv i_59017(.A(queue[153]), .Z(n_42341));
	notech_inv i_59018(.A(n_35999), .Z(n_42342));
	notech_inv i_59019(.A(queue[154]), .Z(n_42343));
	notech_inv i_59020(.A(n_36005), .Z(n_42344));
	notech_inv i_59021(.A(queue[155]), .Z(n_42345));
	notech_inv i_59022(.A(n_36011), .Z(n_42346));
	notech_inv i_59023(.A(queue[156]), .Z(n_42347));
	notech_inv i_59024(.A(n_36017), .Z(n_42348));
	notech_inv i_59025(.A(queue[157]), .Z(n_42349));
	notech_inv i_59026(.A(n_36023), .Z(n_42350));
	notech_inv i_59027(.A(queue[158]), .Z(n_42351));
	notech_inv i_59028(.A(n_36029), .Z(n_42352));
	notech_inv i_59029(.A(queue[159]), .Z(n_42353));
	notech_inv i_59030(.A(n_36035), .Z(n_42354));
	notech_inv i_59031(.A(queue[160]), .Z(n_42355));
	notech_inv i_59032(.A(n_36041), .Z(n_42356));
	notech_inv i_59033(.A(queue[161]), .Z(n_42357));
	notech_inv i_59034(.A(n_36047), .Z(n_42358));
	notech_inv i_59035(.A(queue[162]), .Z(n_42359));
	notech_inv i_59036(.A(n_36053), .Z(n_42360));
	notech_inv i_59037(.A(queue[163]), .Z(n_42361));
	notech_inv i_59038(.A(n_36059), .Z(n_42362));
	notech_inv i_59039(.A(queue[164]), .Z(n_42363));
	notech_inv i_59040(.A(n_36065), .Z(n_42364));
	notech_inv i_59041(.A(queue[165]), .Z(n_42365));
	notech_inv i_59042(.A(n_36071), .Z(n_42366));
	notech_inv i_59043(.A(queue[166]), .Z(n_42367));
	notech_inv i_59044(.A(n_36077), .Z(n_42368));
	notech_inv i_59045(.A(queue[167]), .Z(n_42369));
	notech_inv i_59046(.A(n_36083), .Z(n_42370));
	notech_inv i_59047(.A(queue[168]), .Z(n_42371));
	notech_inv i_59048(.A(n_36089), .Z(n_42372));
	notech_inv i_59049(.A(queue[169]), .Z(n_42373));
	notech_inv i_59050(.A(n_36095), .Z(n_42374));
	notech_inv i_59051(.A(queue[170]), .Z(n_42375));
	notech_inv i_59052(.A(n_36101), .Z(n_42376));
	notech_inv i_59053(.A(queue[171]), .Z(n_42377));
	notech_inv i_59054(.A(n_36107), .Z(n_42378));
	notech_inv i_59055(.A(queue[172]), .Z(n_42379));
	notech_inv i_59056(.A(n_36113), .Z(n_42380));
	notech_inv i_59057(.A(queue[173]), .Z(n_42381));
	notech_inv i_59058(.A(n_36119), .Z(n_42382));
	notech_inv i_59059(.A(queue[174]), .Z(n_42383));
	notech_inv i_59060(.A(n_36125), .Z(n_42384));
	notech_inv i_59061(.A(queue[175]), .Z(n_42385));
	notech_inv i_59062(.A(n_36131), .Z(n_42386));
	notech_inv i_59063(.A(queue[176]), .Z(n_42387));
	notech_inv i_59064(.A(n_36137), .Z(n_42388));
	notech_inv i_59065(.A(queue[177]), .Z(n_42389));
	notech_inv i_59066(.A(n_36143), .Z(n_42390));
	notech_inv i_59067(.A(queue[178]), .Z(n_42391));
	notech_inv i_59068(.A(n_36149), .Z(n_42392));
	notech_inv i_59069(.A(queue[179]), .Z(n_42393));
	notech_inv i_59070(.A(n_36155), .Z(n_42394));
	notech_inv i_59071(.A(queue[180]), .Z(n_42395));
	notech_inv i_59072(.A(n_36161), .Z(n_42396));
	notech_inv i_59073(.A(queue[181]), .Z(n_42397));
	notech_inv i_59074(.A(n_36167), .Z(n_42398));
	notech_inv i_59075(.A(queue[182]), .Z(n_42399));
	notech_inv i_59076(.A(n_36173), .Z(n_42400));
	notech_inv i_59077(.A(queue[183]), .Z(n_42401));
	notech_inv i_59078(.A(n_36179), .Z(n_42402));
	notech_inv i_59079(.A(queue[184]), .Z(n_42403));
	notech_inv i_59080(.A(n_36185), .Z(n_42404));
	notech_inv i_59081(.A(queue[185]), .Z(n_42405));
	notech_inv i_59082(.A(n_36191), .Z(n_42406));
	notech_inv i_59083(.A(queue[186]), .Z(n_42407));
	notech_inv i_59084(.A(n_36197), .Z(n_42408));
	notech_inv i_59085(.A(queue[187]), .Z(n_42409));
	notech_inv i_59086(.A(n_36203), .Z(n_42410));
	notech_inv i_59087(.A(queue[188]), .Z(n_42411));
	notech_inv i_59088(.A(n_36209), .Z(n_42412));
	notech_inv i_59089(.A(queue[189]), .Z(n_42413));
	notech_inv i_59090(.A(n_36215), .Z(n_42414));
	notech_inv i_59091(.A(queue[190]), .Z(n_42415));
	notech_inv i_59092(.A(n_36221), .Z(n_42416));
	notech_inv i_59093(.A(queue[191]), .Z(n_42417));
	notech_inv i_59094(.A(n_36227), .Z(n_42418));
	notech_inv i_59095(.A(queue[192]), .Z(n_42419));
	notech_inv i_59096(.A(n_36233), .Z(n_42420));
	notech_inv i_59097(.A(queue[193]), .Z(n_42421));
	notech_inv i_59098(.A(n_36239), .Z(n_42422));
	notech_inv i_59099(.A(queue[194]), .Z(n_42423));
	notech_inv i_59100(.A(n_36245), .Z(n_42424));
	notech_inv i_59101(.A(queue[195]), .Z(n_42425));
	notech_inv i_59102(.A(n_36251), .Z(n_42426));
	notech_inv i_59103(.A(queue[196]), .Z(n_42427));
	notech_inv i_59104(.A(n_36257), .Z(n_42428));
	notech_inv i_59105(.A(queue[197]), .Z(n_42429));
	notech_inv i_59106(.A(n_36263), .Z(n_42430));
	notech_inv i_59107(.A(queue[198]), .Z(n_42431));
	notech_inv i_59108(.A(n_36269), .Z(n_42432));
	notech_inv i_59109(.A(queue[199]), .Z(n_42433));
	notech_inv i_59110(.A(n_36275), .Z(n_42434));
	notech_inv i_59111(.A(queue[200]), .Z(n_42435));
	notech_inv i_59112(.A(n_36281), .Z(n_42436));
	notech_inv i_59113(.A(queue[201]), .Z(n_42437));
	notech_inv i_59114(.A(n_36287), .Z(n_42438));
	notech_inv i_59115(.A(queue[202]), .Z(n_42439));
	notech_inv i_59116(.A(n_36293), .Z(n_42440));
	notech_inv i_59117(.A(queue[203]), .Z(n_42441));
	notech_inv i_59118(.A(n_36299), .Z(n_42442));
	notech_inv i_59119(.A(queue[204]), .Z(n_42443));
	notech_inv i_59120(.A(n_36305), .Z(n_42444));
	notech_inv i_59121(.A(queue[205]), .Z(n_42445));
	notech_inv i_59122(.A(n_36311), .Z(n_42446));
	notech_inv i_59123(.A(queue[206]), .Z(n_42447));
	notech_inv i_59124(.A(n_36317), .Z(n_42448));
	notech_inv i_59125(.A(queue[207]), .Z(n_42449));
	notech_inv i_59126(.A(n_36323), .Z(n_42450));
	notech_inv i_59127(.A(queue[208]), .Z(n_42451));
	notech_inv i_59128(.A(n_36329), .Z(n_42452));
	notech_inv i_59129(.A(queue[209]), .Z(n_42453));
	notech_inv i_59130(.A(n_36335), .Z(n_42454));
	notech_inv i_59131(.A(queue[210]), .Z(n_42455));
	notech_inv i_59132(.A(n_36341), .Z(n_42456));
	notech_inv i_59133(.A(queue[211]), .Z(n_42457));
	notech_inv i_59134(.A(n_36347), .Z(n_42458));
	notech_inv i_59135(.A(queue[212]), .Z(n_42459));
	notech_inv i_59136(.A(n_36353), .Z(n_42460));
	notech_inv i_59137(.A(queue[213]), .Z(n_42461));
	notech_inv i_59138(.A(n_36359), .Z(n_42462));
	notech_inv i_59139(.A(queue[214]), .Z(n_42463));
	notech_inv i_59140(.A(n_36365), .Z(n_42464));
	notech_inv i_59141(.A(queue[215]), .Z(n_42465));
	notech_inv i_59142(.A(n_36371), .Z(n_42466));
	notech_inv i_59143(.A(queue[216]), .Z(n_42467));
	notech_inv i_59144(.A(n_36377), .Z(n_42468));
	notech_inv i_59145(.A(queue[217]), .Z(n_42469));
	notech_inv i_59146(.A(n_36383), .Z(n_42470));
	notech_inv i_59147(.A(queue[218]), .Z(n_42471));
	notech_inv i_59148(.A(n_36389), .Z(n_42472));
	notech_inv i_59149(.A(queue[219]), .Z(n_42473));
	notech_inv i_59150(.A(n_36395), .Z(n_42474));
	notech_inv i_59151(.A(queue[220]), .Z(n_42475));
	notech_inv i_59152(.A(n_36401), .Z(n_42476));
	notech_inv i_59153(.A(queue[221]), .Z(n_42477));
	notech_inv i_59154(.A(n_36407), .Z(n_42478));
	notech_inv i_59155(.A(queue[222]), .Z(n_42479));
	notech_inv i_59156(.A(n_36413), .Z(n_42480));
	notech_inv i_59157(.A(queue[223]), .Z(n_42481));
	notech_inv i_59158(.A(n_36419), .Z(n_42482));
	notech_inv i_59159(.A(queue[224]), .Z(n_42483));
	notech_inv i_59160(.A(n_36425), .Z(n_42484));
	notech_inv i_59161(.A(queue[225]), .Z(n_42485));
	notech_inv i_59162(.A(n_36431), .Z(n_42486));
	notech_inv i_59163(.A(queue[226]), .Z(n_42487));
	notech_inv i_59164(.A(n_36437), .Z(n_42488));
	notech_inv i_59165(.A(queue[227]), .Z(n_42489));
	notech_inv i_59166(.A(n_36443), .Z(n_42490));
	notech_inv i_59167(.A(queue[228]), .Z(n_42491));
	notech_inv i_59168(.A(n_36449), .Z(n_42492));
	notech_inv i_59169(.A(queue[229]), .Z(n_42493));
	notech_inv i_59170(.A(n_36455), .Z(n_42494));
	notech_inv i_59171(.A(queue[230]), .Z(n_42495));
	notech_inv i_59172(.A(n_36461), .Z(n_42496));
	notech_inv i_59173(.A(queue[231]), .Z(n_42497));
	notech_inv i_59174(.A(n_36467), .Z(n_42498));
	notech_inv i_59175(.A(queue[232]), .Z(n_42499));
	notech_inv i_59176(.A(n_36473), .Z(n_42500));
	notech_inv i_59177(.A(queue[233]), .Z(n_42501));
	notech_inv i_59178(.A(n_36479), .Z(n_42502));
	notech_inv i_59179(.A(queue[234]), .Z(n_42503));
	notech_inv i_59180(.A(n_36485), .Z(n_42504));
	notech_inv i_59181(.A(queue[235]), .Z(n_42505));
	notech_inv i_59182(.A(n_36491), .Z(n_42506));
	notech_inv i_59183(.A(queue[236]), .Z(n_42507));
	notech_inv i_59184(.A(n_36497), .Z(n_42508));
	notech_inv i_59185(.A(queue[237]), .Z(n_42509));
	notech_inv i_59186(.A(n_36503), .Z(n_42510));
	notech_inv i_59187(.A(queue[238]), .Z(n_42511));
	notech_inv i_59188(.A(n_36509), .Z(n_42512));
	notech_inv i_59189(.A(queue[239]), .Z(n_42513));
	notech_inv i_59190(.A(n_36515), .Z(n_42514));
	notech_inv i_59191(.A(queue[240]), .Z(n_42515));
	notech_inv i_59192(.A(n_36521), .Z(n_42516));
	notech_inv i_59193(.A(queue[241]), .Z(n_42517));
	notech_inv i_59194(.A(n_36527), .Z(n_42518));
	notech_inv i_59195(.A(queue[242]), .Z(n_42519));
	notech_inv i_59196(.A(n_36533), .Z(n_42520));
	notech_inv i_59197(.A(queue[243]), .Z(n_42521));
	notech_inv i_59198(.A(n_36539), .Z(n_42522));
	notech_inv i_59199(.A(queue[244]), .Z(n_42523));
	notech_inv i_59200(.A(n_36545), .Z(n_42524));
	notech_inv i_59201(.A(queue[245]), .Z(n_42525));
	notech_inv i_59202(.A(n_36551), .Z(n_42526));
	notech_inv i_59203(.A(queue[246]), .Z(n_42527));
	notech_inv i_59204(.A(n_36557), .Z(n_42528));
	notech_inv i_59205(.A(queue[247]), .Z(n_42529));
	notech_inv i_59206(.A(n_36563), .Z(n_42530));
	notech_inv i_59207(.A(queue[248]), .Z(n_42531));
	notech_inv i_59208(.A(n_36569), .Z(n_42532));
	notech_inv i_59209(.A(queue[249]), .Z(n_42533));
	notech_inv i_59210(.A(n_36575), .Z(n_42534));
	notech_inv i_59211(.A(queue[250]), .Z(n_42535));
	notech_inv i_59212(.A(n_36581), .Z(n_42536));
	notech_inv i_59213(.A(queue[251]), .Z(n_42537));
	notech_inv i_59214(.A(n_36587), .Z(n_42538));
	notech_inv i_59215(.A(queue[252]), .Z(n_42539));
	notech_inv i_59216(.A(n_36593), .Z(n_42540));
	notech_inv i_59217(.A(queue[253]), .Z(n_42541));
	notech_inv i_59218(.A(n_36599), .Z(n_42542));
	notech_inv i_59219(.A(queue[254]), .Z(n_42543));
	notech_inv i_59220(.A(n_36605), .Z(n_42544));
	notech_inv i_59221(.A(queue[255]), .Z(n_42545));
	notech_inv i_59223(.A(addrshft[0]), .Z(n_42547));
	notech_inv i_59224(.A(addrshft[1]), .Z(n_42548));
	notech_inv i_59225(.A(addrshft[2]), .Z(n_42549));
	notech_inv i_59226(.A(squeue_097103), .Z(squeue[0]));
	notech_inv i_59227(.A(squeue_197102), .Z(squeue[1]));
	notech_inv i_59228(.A(squeue_297101), .Z(squeue[2]));
	notech_inv i_59229(.A(squeue_397100), .Z(squeue[3]));
	notech_inv i_59230(.A(squeue_497099), .Z(squeue[4]));
	notech_inv i_59231(.A(squeue_597098), .Z(squeue[5]));
	notech_inv i_59232(.A(squeue_697097), .Z(squeue[6]));
	notech_inv i_59233(.A(squeue_897096), .Z(squeue[8]));
	notech_inv i_59234(.A(squeue_997095), .Z(squeue[9]));
	notech_inv i_59235(.A(squeue_1097094), .Z(squeue[10]));
	notech_inv i_59236(.A(squeue_1197093), .Z(squeue[11]));
	notech_inv i_59237(.A(squeue_1297092), .Z(squeue[12]));
	notech_inv i_59238(.A(squeue_1397091), .Z(squeue[13]));
	notech_inv i_59239(.A(squeue_1597090), .Z(squeue[15]));
	notech_inv i_59240(.A(squeue_1697089), .Z(squeue[16]));
	notech_inv i_59241(.A(squeue_1797088), .Z(squeue[17]));
	notech_inv i_59242(.A(squeue_1897087), .Z(squeue[18]));
	notech_inv i_59243(.A(squeue_1997086), .Z(squeue[19]));
	notech_inv i_59244(.A(squeue_2097085), .Z(squeue[20]));
	notech_inv i_59245(.A(squeue_2197084), .Z(squeue[21]));
	notech_inv i_59246(.A(squeue_2297083), .Z(squeue[22]));
	notech_inv i_59247(.A(squeue_2397082), .Z(squeue[23]));
	notech_inv i_59248(.A(squeue_2497081), .Z(squeue[24]));
	notech_inv i_59249(.A(squeue_2597080), .Z(squeue[25]));
	notech_inv i_59250(.A(squeue_2697079), .Z(squeue[26]));
	notech_inv i_59251(.A(squeue_2797078), .Z(squeue[27]));
	notech_inv i_59252(.A(squeue_2897077), .Z(squeue[28]));
	notech_inv i_59253(.A(squeue_3097076), .Z(squeue[30]));
	notech_inv i_59254(.A(squeue_3197075), .Z(squeue[31]));
	notech_inv i_59255(.A(squeue_3297074), .Z(squeue[32]));
	notech_inv i_59256(.A(squeue_3397073), .Z(squeue[33]));
	notech_inv i_59257(.A(squeue_3497072), .Z(squeue[34]));
	notech_inv i_59258(.A(squeue_3597071), .Z(squeue[35]));
	notech_inv i_59259(.A(squeue_3697070), .Z(squeue[36]));
	notech_inv i_59260(.A(squeue_3897069), .Z(squeue[38]));
	notech_inv i_59261(.A(squeue_3997068), .Z(squeue[39]));
	notech_inv i_59262(.A(squeue_4097067), .Z(squeue[40]));
	notech_inv i_59263(.A(squeue_4197066), .Z(squeue[41]));
	notech_inv i_59264(.A(squeue_4297065), .Z(squeue[42]));
	notech_inv i_59265(.A(squeue_4397064), .Z(squeue[43]));
	notech_inv i_59266(.A(squeue_4497063), .Z(squeue[44]));
	notech_inv i_59267(.A(squeue_4597062), .Z(squeue[45]));
	notech_inv i_59268(.A(squeue_4697061), .Z(squeue[46]));
	notech_inv i_59269(.A(squeue_4797060), .Z(squeue[47]));
	notech_inv i_59270(.A(squeue_4897059), .Z(squeue[48]));
	notech_inv i_59271(.A(squeue_4997058), .Z(squeue[49]));
	notech_inv i_59272(.A(squeue_5097057), .Z(squeue[50]));
	notech_inv i_59273(.A(squeue_5197056), .Z(squeue[51]));
	notech_inv i_59274(.A(squeue_5297055), .Z(squeue[52]));
	notech_inv i_59275(.A(squeue_5397054), .Z(squeue[53]));
	notech_inv i_59276(.A(squeue_6597053), .Z(squeue[65]));
	notech_inv i_59277(.A(nbus_12105[4]), .Z(n_42601));
	notech_inv i_59278(.A(nbus_12105[5]), .Z(n_42602));
	notech_inv i_59279(.A(idata[0]), .Z(n_42603));
	notech_inv i_59280(.A(idata[1]), .Z(n_42604));
	notech_inv i_59281(.A(idata[2]), .Z(n_42605));
	notech_inv i_59282(.A(idata[3]), .Z(n_42606));
	notech_inv i_59283(.A(idata[4]), .Z(n_42607));
	notech_inv i_59284(.A(idata[5]), .Z(n_42608));
	notech_inv i_59285(.A(idata[6]), .Z(n_42609));
	notech_inv i_59286(.A(idata[7]), .Z(n_42610));
	notech_inv i_59287(.A(idata[8]), .Z(n_42611));
	notech_inv i_59288(.A(idata[9]), .Z(n_42612));
	notech_inv i_59289(.A(idata[10]), .Z(n_42613));
	notech_inv i_59290(.A(idata[11]), .Z(n_42614));
	notech_inv i_59291(.A(idata[12]), .Z(n_42615));
	notech_inv i_59292(.A(idata[13]), .Z(n_42616));
	notech_inv i_59293(.A(idata[14]), .Z(n_42617));
	notech_inv i_59294(.A(idata[15]), .Z(n_42618));
	notech_inv i_59295(.A(idata[16]), .Z(n_42619));
	notech_inv i_59296(.A(idata[17]), .Z(n_42620));
	notech_inv i_59297(.A(idata[18]), .Z(n_42621));
	notech_inv i_59298(.A(idata[19]), .Z(n_42622));
	notech_inv i_59299(.A(idata[20]), .Z(n_42623));
	notech_inv i_59300(.A(idata[21]), .Z(n_42624));
	notech_inv i_59301(.A(idata[22]), .Z(n_42625));
	notech_inv i_59302(.A(idata[23]), .Z(n_42626));
	notech_inv i_59303(.A(idata[24]), .Z(n_42627));
	notech_inv i_59304(.A(idata[25]), .Z(n_42628));
	notech_inv i_59305(.A(idata[26]), .Z(n_42629));
	notech_inv i_59306(.A(idata[27]), .Z(n_42630));
	notech_inv i_59307(.A(idata[28]), .Z(n_42631));
	notech_inv i_59308(.A(idata[29]), .Z(n_42632));
	notech_inv i_59309(.A(idata[30]), .Z(n_42633));
	notech_inv i_59310(.A(idata[31]), .Z(n_42634));
	notech_inv i_59311(.A(idata[32]), .Z(n_42635));
	notech_inv i_59312(.A(idata[33]), .Z(n_42636));
	notech_inv i_59313(.A(idata[34]), .Z(n_42637));
	notech_inv i_59314(.A(idata[35]), .Z(n_42638));
	notech_inv i_59315(.A(idata[36]), .Z(n_42639));
	notech_inv i_59316(.A(idata[37]), .Z(n_42640));
	notech_inv i_59317(.A(idata[38]), .Z(n_42641));
	notech_inv i_59318(.A(idata[39]), .Z(n_42642));
	notech_inv i_59319(.A(idata[40]), .Z(n_42643));
	notech_inv i_59320(.A(idata[41]), .Z(n_42644));
	notech_inv i_59321(.A(idata[42]), .Z(n_42645));
	notech_inv i_59322(.A(idata[43]), .Z(n_42646));
	notech_inv i_59323(.A(idata[44]), .Z(n_42647));
	notech_inv i_59324(.A(idata[45]), .Z(n_42648));
	notech_inv i_59325(.A(idata[46]), .Z(n_42649));
	notech_inv i_59326(.A(idata[47]), .Z(n_42650));
	notech_inv i_59327(.A(idata[48]), .Z(n_42651));
	notech_inv i_59328(.A(idata[49]), .Z(n_42652));
	notech_inv i_59329(.A(idata[50]), .Z(n_42653));
	notech_inv i_59330(.A(idata[51]), .Z(n_42654));
	notech_inv i_59331(.A(idata[52]), .Z(n_42655));
	notech_inv i_59332(.A(idata[53]), .Z(n_42656));
	notech_inv i_59333(.A(idata[54]), .Z(n_42657));
	notech_inv i_59334(.A(idata[55]), .Z(n_42658));
	notech_inv i_59335(.A(idata[56]), .Z(n_42659));
	notech_inv i_59336(.A(idata[57]), .Z(n_42660));
	notech_inv i_59337(.A(idata[58]), .Z(n_42661));
	notech_inv i_59338(.A(idata[59]), .Z(n_42662));
	notech_inv i_59339(.A(idata[60]), .Z(n_42663));
	notech_inv i_59340(.A(idata[61]), .Z(n_42664));
	notech_inv i_59341(.A(idata[62]), .Z(n_42665));
	notech_inv i_59342(.A(idata[63]), .Z(n_42666));
	notech_inv i_59343(.A(idata[64]), .Z(n_42667));
	notech_inv i_59344(.A(idata[65]), .Z(n_42668));
	notech_inv i_59345(.A(idata[66]), .Z(n_42669));
	notech_inv i_59346(.A(idata[67]), .Z(n_42670));
	notech_inv i_59347(.A(idata[68]), .Z(n_42671));
	notech_inv i_59348(.A(idata[69]), .Z(n_42672));
	notech_inv i_59349(.A(idata[70]), .Z(n_42673));
	notech_inv i_59350(.A(idata[71]), .Z(n_42674));
	notech_inv i_59351(.A(idata[72]), .Z(n_42675));
	notech_inv i_59352(.A(idata[73]), .Z(n_42676));
	notech_inv i_59353(.A(idata[74]), .Z(n_42677));
	notech_inv i_59354(.A(idata[75]), .Z(n_42678));
	notech_inv i_59355(.A(idata[76]), .Z(n_42679));
	notech_inv i_59356(.A(idata[77]), .Z(n_42680));
	notech_inv i_59357(.A(idata[78]), .Z(n_42681));
	notech_inv i_59358(.A(idata[79]), .Z(n_42682));
	notech_inv i_59359(.A(idata[80]), .Z(n_42683));
	notech_inv i_59360(.A(idata[81]), .Z(n_42684));
	notech_inv i_59361(.A(idata[82]), .Z(n_42685));
	notech_inv i_59362(.A(idata[83]), .Z(n_42686));
	notech_inv i_59363(.A(idata[84]), .Z(n_42687));
	notech_inv i_59364(.A(idata[85]), .Z(n_42688));
	notech_inv i_59365(.A(idata[86]), .Z(n_42689));
	notech_inv i_59366(.A(idata[87]), .Z(n_42690));
	notech_inv i_59367(.A(idata[88]), .Z(n_42691));
	notech_inv i_59368(.A(idata[89]), .Z(n_42692));
	notech_inv i_59369(.A(idata[90]), .Z(n_42693));
	notech_inv i_59370(.A(idata[91]), .Z(n_42694));
	notech_inv i_59371(.A(idata[92]), .Z(n_42695));
	notech_inv i_59372(.A(idata[93]), .Z(n_42696));
	notech_inv i_59373(.A(idata[94]), .Z(n_42697));
	notech_inv i_59374(.A(idata[95]), .Z(n_42698));
	notech_inv i_59375(.A(idata[96]), .Z(n_42699));
	notech_inv i_59376(.A(idata[97]), .Z(n_42700));
	notech_inv i_59377(.A(idata[98]), .Z(n_42701));
	notech_inv i_59378(.A(idata[99]), .Z(n_42702));
	notech_inv i_59379(.A(idata[100]), .Z(n_42703));
	notech_inv i_59380(.A(idata[101]), .Z(n_42704));
	notech_inv i_59381(.A(idata[102]), .Z(n_42705));
	notech_inv i_59382(.A(idata[103]), .Z(n_42706));
	notech_inv i_59383(.A(idata[104]), .Z(n_42707));
	notech_inv i_59384(.A(idata[105]), .Z(n_42708));
	notech_inv i_59385(.A(idata[106]), .Z(n_42709));
	notech_inv i_59386(.A(idata[107]), .Z(n_42710));
	notech_inv i_59387(.A(idata[108]), .Z(n_42711));
	notech_inv i_59388(.A(idata[109]), .Z(n_42712));
	notech_inv i_59389(.A(idata[110]), .Z(n_42713));
	notech_inv i_59390(.A(idata[111]), .Z(n_42714));
	notech_inv i_59391(.A(idata[112]), .Z(n_42715));
	notech_inv i_59392(.A(idata[113]), .Z(n_42716));
	notech_inv i_59393(.A(idata[114]), .Z(n_42717));
	notech_inv i_59394(.A(idata[115]), .Z(n_42718));
	notech_inv i_59395(.A(idata[116]), .Z(n_42719));
	notech_inv i_59396(.A(idata[117]), .Z(n_42720));
	notech_inv i_59397(.A(idata[118]), .Z(n_42721));
	notech_inv i_59398(.A(idata[119]), .Z(n_42722));
	notech_inv i_59399(.A(idata[120]), .Z(n_42723));
	notech_inv i_59400(.A(idata[121]), .Z(n_42724));
	notech_inv i_59401(.A(idata[122]), .Z(n_42725));
	notech_inv i_59402(.A(idata[123]), .Z(n_42726));
	notech_inv i_59403(.A(idata[124]), .Z(n_42727));
	notech_inv i_59404(.A(idata[125]), .Z(n_42728));
	notech_inv i_59405(.A(idata[126]), .Z(n_42729));
	notech_inv i_59406(.A(idata[127]), .Z(n_42730));
	notech_inv i_59407(.A(valid_len_097049), .Z(valid_len[0]));
	notech_inv i_59408(.A(valid_len_197052), .Z(valid_len[1]));
	notech_inv i_59409(.A(valid_len_297051), .Z(valid_len[2]));
	notech_inv i_59410(.A(valid_len_397050), .Z(valid_len[3]));
	notech_inv i_59411(.A(valid_len_497048), .Z(valid_len[4]));
	notech_inv i_59412(.A(\queue_0[26] ), .Z(n_42736));
	notech_inv i_59413(.A(\queue_0[18] ), .Z(n_42737));
	notech_inv i_59414(.A(\queue_0[10] ), .Z(n_42738));
	notech_inv i_59415(.A(\queue_0[2] ), .Z(n_42739));
	notech_inv i_59416(.A(busy_ram), .Z(n_42740));
	notech_inv i_59417(.A(n_60396), .Z(n_42741));
	notech_inv i_59418(.A(pc_pg_fault), .Z(n_42742));
	notech_inv i_59419(.A(n_61549), .Z(n_42743));
	notech_inv i_59420(.A(\queue_0[126] ), .Z(n_42744));
	notech_inv i_59421(.A(\queue_0[124] ), .Z(n_42745));
	notech_inv i_59422(.A(\queue_0[123] ), .Z(n_42746));
	notech_inv i_59423(.A(\queue_0[122] ), .Z(n_42747));
	notech_inv i_59424(.A(\queue_0[121] ), .Z(n_42748));
	notech_inv i_59425(.A(\queue_0[120] ), .Z(n_42749));
	notech_inv i_59426(.A(\queue_0[119] ), .Z(n_42750));
	notech_inv i_59427(.A(\queue_0[118] ), .Z(n_42751));
	notech_inv i_59428(.A(\queue_0[117] ), .Z(n_42752));
	notech_inv i_59429(.A(\queue_0[116] ), .Z(n_42753));
	notech_inv i_59430(.A(\queue_0[115] ), .Z(n_42754));
	notech_inv i_59431(.A(\queue_0[114] ), .Z(n_42755));
	notech_inv i_59432(.A(\queue_0[113] ), .Z(n_42756));
	notech_inv i_59433(.A(\queue_0[112] ), .Z(n_42757));
	notech_inv i_59434(.A(\queue_0[111] ), .Z(n_42758));
	notech_inv i_59435(.A(\queue_0[110] ), .Z(n_42759));
	notech_inv i_59436(.A(\queue_0[109] ), .Z(n_42760));
	notech_inv i_59437(.A(\queue_0[108] ), .Z(n_42761));
	notech_inv i_59438(.A(\queue_0[107] ), .Z(n_42762));
	notech_inv i_59439(.A(\queue_0[106] ), .Z(n_42763));
	notech_inv i_59440(.A(\queue_0[105] ), .Z(n_42764));
	notech_inv i_59441(.A(\queue_0[104] ), .Z(n_42765));
	notech_inv i_59442(.A(\queue_0[103] ), .Z(n_42766));
	notech_inv i_59443(.A(\queue_0[102] ), .Z(n_42767));
	notech_inv i_59444(.A(\queue_0[101] ), .Z(n_42768));
	notech_inv i_59445(.A(\queue_0[100] ), .Z(n_42769));
	notech_inv i_59446(.A(\queue_0[99] ), .Z(n_42770));
	notech_inv i_59447(.A(\queue_0[98] ), .Z(n_42771));
	notech_inv i_59448(.A(\queue_0[97] ), .Z(n_42772));
	notech_inv i_59449(.A(\queue_0[96] ), .Z(n_42773));
	notech_inv i_59450(.A(\queue_0[95] ), .Z(n_42774));
	notech_inv i_59451(.A(\queue_0[94] ), .Z(n_42775));
	notech_inv i_59452(.A(\queue_0[93] ), .Z(n_42776));
	notech_inv i_59453(.A(\queue_0[92] ), .Z(n_42777));
	notech_inv i_59454(.A(\queue_0[91] ), .Z(n_42778));
	notech_inv i_59455(.A(\queue_0[90] ), .Z(n_42779));
	notech_inv i_59456(.A(\queue_0[89] ), .Z(n_42780));
	notech_inv i_59457(.A(\queue_0[87] ), .Z(n_42781));
	notech_inv i_59458(.A(\queue_0[86] ), .Z(n_42782));
	notech_inv i_59459(.A(\queue_0[85] ), .Z(n_42783));
	notech_inv i_59460(.A(\queue_0[84] ), .Z(n_42784));
	notech_inv i_59461(.A(\queue_0[83] ), .Z(n_42785));
	notech_inv i_59462(.A(\queue_0[82] ), .Z(n_42786));
	notech_inv i_59463(.A(\queue_0[81] ), .Z(n_42787));
	notech_inv i_59464(.A(\queue_0[80] ), .Z(n_42788));
	notech_inv i_59465(.A(\queue_0[79] ), .Z(n_42789));
	notech_inv i_59466(.A(\queue_0[78] ), .Z(n_42790));
	notech_inv i_59467(.A(\queue_0[77] ), .Z(n_42791));
	notech_inv i_59468(.A(\queue_0[76] ), .Z(n_42792));
	notech_inv i_59469(.A(\queue_0[75] ), .Z(n_42793));
	notech_inv i_59470(.A(\queue_0[74] ), .Z(n_42794));
	notech_inv i_59471(.A(\queue_0[73] ), .Z(n_42795));
	notech_inv i_59472(.A(\queue_0[72] ), .Z(n_42796));
	notech_inv i_59473(.A(\queue_0[71] ), .Z(n_42797));
	notech_inv i_59474(.A(\queue_0[69] ), .Z(n_42798));
	notech_inv i_59475(.A(\queue_0[68] ), .Z(n_42799));
	notech_inv i_59476(.A(\queue_0[67] ), .Z(n_42800));
	notech_inv i_59477(.A(\queue_0[66] ), .Z(n_42801));
	notech_inv i_59478(.A(\queue_0[65] ), .Z(n_42802));
	notech_inv i_59479(.A(\queue_0[64] ), .Z(n_42803));
	notech_inv i_59480(.A(\queue_0[63] ), .Z(n_42804));
	notech_inv i_59481(.A(\queue_0[62] ), .Z(n_42805));
	notech_inv i_59482(.A(\queue_0[61] ), .Z(n_42806));
	notech_inv i_59483(.A(\queue_0[60] ), .Z(n_42807));
	notech_inv i_59484(.A(\queue_0[59] ), .Z(n_42808));
	notech_inv i_59485(.A(\queue_0[57] ), .Z(n_42809));
	notech_inv i_59486(.A(\queue_0[56] ), .Z(n_42810));
	notech_inv i_59487(.A(\queue_0[55] ), .Z(n_42811));
	notech_inv i_59488(.A(\queue_0[54] ), .Z(n_42812));
	notech_inv i_59489(.A(\queue_0[53] ), .Z(n_42813));
	notech_inv i_59490(.A(\queue_0[52] ), .Z(n_42814));
	notech_inv i_59491(.A(\queue_0[51] ), .Z(n_42815));
	notech_inv i_59492(.A(\queue_0[50] ), .Z(n_42816));
	notech_inv i_59493(.A(\queue_0[49] ), .Z(n_42817));
	notech_inv i_59494(.A(\queue_0[48] ), .Z(n_42818));
	notech_inv i_59495(.A(\queue_0[47] ), .Z(n_42819));
	notech_inv i_59496(.A(\queue_0[46] ), .Z(n_42820));
	notech_inv i_59497(.A(\queue_0[45] ), .Z(n_42821));
	notech_inv i_59498(.A(\queue_0[44] ), .Z(n_42822));
	notech_inv i_59499(.A(\queue_0[43] ), .Z(n_42823));
	notech_inv i_59500(.A(\queue_0[42] ), .Z(n_42824));
	notech_inv i_59501(.A(\queue_0[41] ), .Z(n_42825));
	notech_inv i_59502(.A(\queue_0[40] ), .Z(n_42826));
	notech_inv i_59503(.A(\queue_0[39] ), .Z(n_42827));
	notech_inv i_59504(.A(\queue_0[38] ), .Z(n_42828));
	notech_inv i_59505(.A(\queue_0[37] ), .Z(n_42829));
	notech_inv i_59506(.A(\queue_0[36] ), .Z(n_42830));
	notech_inv i_59507(.A(\queue_0[35] ), .Z(n_42831));
	notech_inv i_59508(.A(\queue_0[34] ), .Z(n_42832));
	notech_inv i_59509(.A(\queue_0[33] ), .Z(n_42833));
	notech_inv i_59510(.A(\queue_0[32] ), .Z(n_42834));
	notech_inv i_59511(.A(\queue_0[31] ), .Z(n_42835));
	notech_inv i_59512(.A(\queue_0[30] ), .Z(n_42836));
	notech_inv i_59513(.A(\queue_0[29] ), .Z(n_42837));
	notech_inv i_59514(.A(\queue_0[28] ), .Z(n_42838));
	notech_inv i_59515(.A(\queue_0[27] ), .Z(n_42839));
	notech_inv i_59516(.A(\queue_0[25] ), .Z(n_42840));
	notech_inv i_59517(.A(\queue_0[24] ), .Z(n_42841));
	notech_inv i_59518(.A(\queue_0[23] ), .Z(n_42842));
	notech_inv i_59519(.A(\queue_0[22] ), .Z(n_42843));
	notech_inv i_59520(.A(\queue_0[21] ), .Z(n_42844));
	notech_inv i_59521(.A(\queue_0[20] ), .Z(n_42845));
	notech_inv i_59522(.A(\queue_0[19] ), .Z(n_42846));
	notech_inv i_59523(.A(\queue_0[17] ), .Z(n_42847));
	notech_inv i_59524(.A(\queue_0[16] ), .Z(n_42848));
	notech_inv i_59525(.A(\queue_0[15] ), .Z(n_42849));
	notech_inv i_59526(.A(\queue_0[14] ), .Z(n_42850));
	notech_inv i_59527(.A(\queue_0[13] ), .Z(n_42851));
	notech_inv i_59528(.A(\queue_0[12] ), .Z(n_42852));
	notech_inv i_59529(.A(\queue_0[11] ), .Z(n_42853));
	notech_inv i_59530(.A(\queue_0[9] ), .Z(n_42854));
	notech_inv i_59531(.A(\queue_0[8] ), .Z(n_42855));
	notech_inv i_59532(.A(\queue_0[7] ), .Z(n_42856));
	notech_inv i_59533(.A(\queue_0[6] ), .Z(n_42857));
	notech_inv i_59534(.A(\queue_0[5] ), .Z(n_42858));
	notech_inv i_59535(.A(\queue_0[4] ), .Z(n_42859));
	notech_inv i_59536(.A(\queue_0[3] ), .Z(n_42860));
	notech_inv i_59537(.A(\queue_0[1] ), .Z(n_42861));
	notech_inv i_59538(.A(\queue_0[0] ), .Z(n_42862));
	notech_inv i_59539(.A(\queue_0[58] ), .Z(n_42863));
	notech_inv i_59540(.A(\queue_0[70] ), .Z(n_42864));
	notech_inv i_59541(.A(\queue_0[125] ), .Z(n_42865));
	notech_inv i_59542(.A(\queue_0[127] ), .Z(n_42866));
	notech_inv i_59543(.A(\queue_0[88] ), .Z(n_42867));
	AWDP_ADD_2 i_64381(.O0(addr_0), .addr(iaddr));
	AWDP_EQ_46 i_64380(.O0({n_34674}), .addr(iaddr), .addrf(addrf));
	AWDP_EQ_715217 i_64375(.O0({n_35018}), .tagA(tagA), .addr({iaddr[31], iaddr
		[30], iaddr[29], iaddr[28], iaddr[27], iaddr[26], iaddr[25], iaddr
		[24], iaddr[23], iaddr[22], iaddr[21], iaddr[20], iaddr[19], iaddr
		[18], iaddr[17], iaddr[16], iaddr[15], iaddr[14]}));
	AWDP_ADD_12 i_64362(.O0(nbus_12105), .addrshft(addrshft), .useq_ptr(useq_ptr
		));
	AWDP_INC_1 i_64347(.O0({n_34650, n_34648, n_34646, n_34644, n_34642, n_34640
		, n_34638, n_34636, n_34634, n_34632, n_34630}), .purge_cnt(purge_cnt
		));
	datacache c1(.clk(clk), .A(cacheA), .D({AMBIT_GND, cacheD[148], 
		AMBIT_GND, AMBIT_GND, cacheD[145], cacheD[144], cacheD[143], cacheD
		[142], cacheD[141], cacheD[140], cacheD[139], cacheD[138], cacheD
		[137], cacheD[136], cacheD[135], cacheD[134], cacheD[133], cacheD
		[132], cacheD[131], cacheD[130], cacheD[129], cacheD[128], cacheD
		[127], cacheD[126], cacheD[125], cacheD[124], cacheD[123], cacheD
		[122], cacheD[121], cacheD[120], cacheD[119], cacheD[118], cacheD
		[117], cacheD[116], cacheD[115], cacheD[114], cacheD[113], cacheD
		[112], cacheD[111], cacheD[110], cacheD[109], cacheD[108], cacheD
		[107], cacheD[106], cacheD[105], cacheD[104], cacheD[103], cacheD
		[102], cacheD[101], cacheD[100], cacheD[99], cacheD[98], cacheD[
		97], cacheD[96], cacheD[95], cacheD[94], cacheD[93], cacheD[92],
		 cacheD[91], cacheD[90], cacheD[89], cacheD[88], cacheD[87], cacheD
		[86], cacheD[85], cacheD[84], cacheD[83], cacheD[82], cacheD[81]
		, cacheD[80], cacheD[79], cacheD[78], cacheD[77], cacheD[76], cacheD
		[75], cacheD[74], cacheD[73], cacheD[72], cacheD[71], cacheD[70]
		, cacheD[69], cacheD[68], cacheD[67], cacheD[66], cacheD[65], cacheD
		[64], cacheD[63], cacheD[62], cacheD[61], cacheD[60], cacheD[59]
		, cacheD[58], cacheD[57], cacheD[56], cacheD[55], cacheD[54], cacheD
		[53], cacheD[52], cacheD[51], cacheD[50], cacheD[49], cacheD[48]
		, cacheD[47], cacheD[46], cacheD[45], cacheD[44], cacheD[43], cacheD
		[42], cacheD[41], cacheD[40], cacheD[39], cacheD[38], cacheD[37]
		, cacheD[36], cacheD[35], cacheD[34], cacheD[33], cacheD[32], cacheD
		[31], cacheD[30], cacheD[29], cacheD[28], cacheD[27], cacheD[26]
		, cacheD[25], cacheD[24], cacheD[23], cacheD[22], cacheD[21], cacheD
		[20], cacheD[19], cacheD[18], cacheD[17], cacheD[16], cacheD[15]
		, cacheD[14], cacheD[13], cacheD[12], cacheD[11], cacheD[10], cacheD
		[9], cacheD[8], cacheD[7], cacheD[6], cacheD[5], cacheD[4], cacheD
		[3], cacheD[2], cacheD[1], cacheD[0]}), .Q({tagV[3], tagV[2], tagV
		[1], tagV[0], tagA[17], tagA[16], tagA[15], tagA[14], tagA[13], tagA
		[12], tagA[11], tagA[10], tagA[9], tagA[8], tagA[7], tagA[6], tagA
		[5], tagA[4], tagA[3], tagA[2], tagA[1], tagA[0], \queue_0[127] 
		, \queue_0[126] , \queue_0[125] , \queue_0[124] , \queue_0[123] 
		, \queue_0[122] , \queue_0[121] , \queue_0[120] , \queue_0[119] 
		, \queue_0[118] , \queue_0[117] , \queue_0[116] , \queue_0[115] 
		, \queue_0[114] , \queue_0[113] , \queue_0[112] , \queue_0[111] 
		, \queue_0[110] , \queue_0[109] , \queue_0[108] , \queue_0[107] 
		, \queue_0[106] , \queue_0[105] , \queue_0[104] , \queue_0[103] 
		, \queue_0[102] , \queue_0[101] , \queue_0[100] , \queue_0[99] ,
		 \queue_0[98] , \queue_0[97] , \queue_0[96] , \queue_0[95] , \queue_0[94] 
		, \queue_0[93] , \queue_0[92] , \queue_0[91] , \queue_0[90] , \queue_0[89] 
		, \queue_0[88] , \queue_0[87] , \queue_0[86] , \queue_0[85] , \queue_0[84] 
		, \queue_0[83] , \queue_0[82] , \queue_0[81] , \queue_0[80] , \queue_0[79] 
		, \queue_0[78] , \queue_0[77] , \queue_0[76] , \queue_0[75] , \queue_0[74] 
		, \queue_0[73] , \queue_0[72] , \queue_0[71] , \queue_0[70] , \queue_0[69] 
		, \queue_0[68] , \queue_0[67] , \queue_0[66] , \queue_0[65] , \queue_0[64] 
		, \queue_0[63] , \queue_0[62] , \queue_0[61] , \queue_0[60] , \queue_0[59] 
		, \queue_0[58] , \queue_0[57] , \queue_0[56] , \queue_0[55] , \queue_0[54] 
		, \queue_0[53] , \queue_0[52] , \queue_0[51] , \queue_0[50] , \queue_0[49] 
		, \queue_0[48] , \queue_0[47] , \queue_0[46] , \queue_0[45] , \queue_0[44] 
		, \queue_0[43] , \queue_0[42] , \queue_0[41] , \queue_0[40] , \queue_0[39] 
		, \queue_0[38] , \queue_0[37] , \queue_0[36] , \queue_0[35] , \queue_0[34] 
		, \queue_0[33] , \queue_0[32] , \queue_0[31] , \queue_0[30] , \queue_0[29] 
		, \queue_0[28] , \queue_0[27] , \queue_0[26] , \queue_0[25] , \queue_0[24] 
		, \queue_0[23] , \queue_0[22] , \queue_0[21] , \queue_0[20] , \queue_0[19] 
		, \queue_0[18] , \queue_0[17] , \queue_0[16] , \queue_0[15] , \queue_0[14] 
		, \queue_0[13] , \queue_0[12] , \queue_0[11] , \queue_0[10] , \queue_0[9] 
		, \queue_0[8] , \queue_0[7] , \queue_0[6] , \queue_0[5] , \queue_0[4] 
		, \queue_0[3] , \queue_0[2] , \queue_0[1] , \queue_0[0] }), .WEN
		(codeWEN), .M({AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, 
		AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD
		, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, AMBIT_VDD, 
		AMBIT_VDD}));
endmodule
module core(clk, rstn, ivect, int_main, iack, code_addr, code_data, code_req, code_ack
		, code_wreq, code_wack, code_wdata, readio_data, io_add, writeio_data
		, writeio_req, readio_req, writeio_ack, readio_ack, write_req, write_ack
		, write_data, write_sz, read_sz, write_msk, read_req, read_ack, read_data
		, Daddr, busy_ram, ipg_fault, outstanding);

	input clk;
	input rstn;
	input [7:0] ivect;
	input int_main;
	output iack;
	output [31:0] code_addr;
	input [127:0] code_data;
	output code_req;
	input code_ack;
	output code_wreq;
	input code_wack;
	output [31:0] code_wdata;
	input [31:0] readio_data;
	output [31:0] io_add;
	output [31:0] writeio_data;
	output writeio_req;
	output readio_req;
	input writeio_ack;
	input readio_ack;
	output write_req;
	input write_ack;
	output [31:0] write_data;
	output [1:0] write_sz;
	output [1:0] read_sz;
	output [3:0] write_msk;
	output read_req;
	input read_ack;
	input [31:0] read_data;
	output [31:0] Daddr;
	input busy_ram;
	output ipg_fault;
	output outstanding;

	wire [31:0] write_data_realign;
	wire [31:0] read_data_realign;
	wire [31:0] Daddr_realign;
	wire [5:0] valid_len;
	wire [1:0] int_write_sz;
	wire [31:0] iwrite_data;
	wire [31:0] int_code_addr;
	wire [31:0] icr2;
	wire [31:0] cr2;
	wire [31:0] pc_out;
	wire [31:0] int_Daddr;
	wire [3:0] useq_ptr;
	wire [127:0] queue;
	wire [1:0] nbus_14525;



	realign i_realign(.clk(clk), .rstn(rstn), .write_msk_out(write_msk), .addr_in
		(Daddr_realign), .addr_out({Daddr[31], Daddr[30], Daddr[29], Daddr
		[28], Daddr[27], Daddr[26], Daddr[25], Daddr[24], Daddr[23], Daddr
		[22], Daddr[21], Daddr[20], Daddr[19], Daddr[18], Daddr[17], Daddr
		[16], Daddr[15], Daddr[14], Daddr[13], Daddr[12], Daddr[11], Daddr
		[10], Daddr[9], Daddr[8], Daddr[7], Daddr[6], Daddr[5], Daddr[4]
		, Daddr[3], Daddr[2], UNCONNECTED_000, UNCONNECTED_001}), .write_sz_in
		(nbus_14525), .write_req_in(write_req_realign), .write_req_out(write_req
		), .write_ack_in(write_ack), .write_ack_out(write_ack_realign), 
		.read_req_in(read_req_realign), .read_req_out(read_req), .read_ack_in
		(read_ack), .read_ack_out(read_ack_realign), .read_data_in(read_data
		), .read_data_out(read_data_realign), .write_data_in(write_data_realign
		), .write_data_out(write_data));
	Itlb i_Itlb(.clk(clk), .rstn(rstn), .addr_phys({code_addr[31], code_addr
		[30], code_addr[29], code_addr[28], code_addr[27], code_addr[26]
		, code_addr[25], code_addr[24], code_addr[23], code_addr[22], code_addr
		[21], code_addr[20], code_addr[19], code_addr[18], code_addr[17]
		, code_addr[16], code_addr[15], code_addr[14], code_addr[13], code_addr
		[12], code_addr[11], code_addr[10], code_addr[9], code_addr[8], code_addr
		[7], code_addr[6], code_addr[5], code_addr[4], code_addr[3], code_addr
		[2], UNCONNECTED_002, UNCONNECTED_003}), .cr3({\cr3[31] , \cr3[30] 
		, \cr3[29] , \cr3[28] , \cr3[27] , \cr3[26] , \cr3[25] , \cr3[24] 
		, \cr3[23] , \cr3[22] , \cr3[21] , \cr3[20] , \cr3[19] , \cr3[18] 
		, \cr3[17] , \cr3[16] , \cr3[15] , \cr3[14] , \cr3[13] , \cr3[12] 
		, UNCONNECTED_004, UNCONNECTED_005, UNCONNECTED_006, 
		UNCONNECTED_007, UNCONNECTED_008, UNCONNECTED_009, 
		UNCONNECTED_010, UNCONNECTED_011, UNCONNECTED_012, 
		UNCONNECTED_013, UNCONNECTED_014, UNCONNECTED_015}), .data_miss(
		{code_data[31], code_data[30], code_data[29], code_data[28], code_data
		[27], code_data[26], code_data[25], code_data[24], code_data[23]
		, code_data[22], code_data[21], code_data[20], code_data[19], code_data
		[18], code_data[17], code_data[16], code_data[15], code_data[14]
		, code_data[13], code_data[12], UNCONNECTED_016, UNCONNECTED_017
		, UNCONNECTED_018, UNCONNECTED_019, code_data[7], code_data[6], code_data
		[5], code_data[4], code_data[3], code_data[2], code_data[1], code_data
		[0]}), .iDaddr(int_code_addr), .pg_en(pg_en), .owrite_data({
		UNCONNECTED_020, UNCONNECTED_021, UNCONNECTED_022, 
		UNCONNECTED_023, UNCONNECTED_024, UNCONNECTED_025, 
		UNCONNECTED_026, UNCONNECTED_027, UNCONNECTED_028, 
		UNCONNECTED_029, UNCONNECTED_030, UNCONNECTED_031, 
		UNCONNECTED_032, UNCONNECTED_033, UNCONNECTED_034, 
		UNCONNECTED_035, UNCONNECTED_036, UNCONNECTED_037, 
		UNCONNECTED_038, UNCONNECTED_039, UNCONNECTED_040, 
		UNCONNECTED_041, UNCONNECTED_042, UNCONNECTED_043, code_wdata[7]
		, code_wdata[6], code_wdata[5], code_wdata[4], code_wdata[3], code_wdata
		[2], code_wdata[1], code_wdata[0]}), .iread_req(int_code_req), .iread_ack
		(code_ack), .iwrite_ack(code_wack), .oread_req(code_req), .oread_ack
		(int_code_ack), .owrite_req(code_wreq), .pg_fault(n_3135), .cr2(icr2
		), .flush_tlb(flush_Itlb), .busy_ram(busy_ram));
	Dtlb i_Dtlb(.clk(clk), .rstn(rstn), .addr_phys(Daddr_realign), .cr3({\cr3[31] 
		, \cr3[30] , \cr3[29] , \cr3[28] , \cr3[27] , \cr3[26] , \cr3[25] 
		, \cr3[24] , \cr3[23] , \cr3[22] , \cr3[21] , \cr3[20] , \cr3[19] 
		, \cr3[18] , \cr3[17] , \cr3[16] , \cr3[15] , \cr3[14] , \cr3[13] 
		, \cr3[12] , UNCONNECTED_044, UNCONNECTED_045, UNCONNECTED_046, 
		UNCONNECTED_047, UNCONNECTED_048, UNCONNECTED_049, 
		UNCONNECTED_050, UNCONNECTED_051, UNCONNECTED_052, 
		UNCONNECTED_053, UNCONNECTED_054, UNCONNECTED_055}), .cr0({
		UNCONNECTED_056, UNCONNECTED_057, UNCONNECTED_058, 
		UNCONNECTED_059, UNCONNECTED_060, UNCONNECTED_061, 
		UNCONNECTED_062, UNCONNECTED_063, UNCONNECTED_064, 
		UNCONNECTED_065, UNCONNECTED_066, UNCONNECTED_067, 
		UNCONNECTED_068, UNCONNECTED_069, UNCONNECTED_070, \cr0[16] , 
		UNCONNECTED_071, UNCONNECTED_072, UNCONNECTED_073, 
		UNCONNECTED_074, UNCONNECTED_075, UNCONNECTED_076, 
		UNCONNECTED_077, UNCONNECTED_078, UNCONNECTED_079, 
		UNCONNECTED_080, UNCONNECTED_081, UNCONNECTED_082, 
		UNCONNECTED_083, UNCONNECTED_084, UNCONNECTED_085, 
		UNCONNECTED_086}), .data_miss(read_data_realign), .iDaddr(int_Daddr
		), .pg_en(pg_en), .iwrite_data(iwrite_data), .owrite_data(write_data_realign
		), .iread_req(int_read_req), .iread_ack(read_ack_realign), .iwrite_req
		(int_write_req), .iwrite_ack(write_ack_realign), .iwrite_sz(int_write_sz
		), .owrite_sz(nbus_14525), .oread_req(read_req_realign), .oread_ack
		(int_read_ack), .owrite_req(write_req_realign), .owrite_ack(int_write_ack
		), .pg_fault(pg_fault), .wr_fault(wr_fault), .cr2(cr2), .flush_tlb
		(flush_Dtlb), .cs({UNCONNECTED_087, UNCONNECTED_088, 
		UNCONNECTED_089, UNCONNECTED_090, UNCONNECTED_091, 
		UNCONNECTED_092, UNCONNECTED_093, UNCONNECTED_094, 
		UNCONNECTED_095, UNCONNECTED_096, UNCONNECTED_097, 
		UNCONNECTED_098, UNCONNECTED_099, UNCONNECTED_100, 
		UNCONNECTED_101, UNCONNECTED_102, UNCONNECTED_103, 
		UNCONNECTED_104, UNCONNECTED_105, UNCONNECTED_106, 
		UNCONNECTED_107, UNCONNECTED_108, UNCONNECTED_109, 
		UNCONNECTED_110, UNCONNECTED_111, UNCONNECTED_112, 
		UNCONNECTED_113, UNCONNECTED_114, UNCONNECTED_115, 
		UNCONNECTED_116, \cs[1] , \cs[0] }), .pt_fault(pt_fault), .busy_ram
		(busy_ram));
	cpu i_cpu(.clk(clk), .rstn(rstn), .iack(iack), .int_cpu(int_main), .ivect
		(ivect), .cr0({UNCONNECTED_117, UNCONNECTED_118, UNCONNECTED_119
		, UNCONNECTED_120, UNCONNECTED_121, UNCONNECTED_122, 
		UNCONNECTED_123, UNCONNECTED_124, UNCONNECTED_125, 
		UNCONNECTED_126, UNCONNECTED_127, UNCONNECTED_128, 
		UNCONNECTED_129, UNCONNECTED_130, UNCONNECTED_131, \cr0[16] , 
		UNCONNECTED_132, UNCONNECTED_133, UNCONNECTED_134, 
		UNCONNECTED_135, UNCONNECTED_136, UNCONNECTED_137, 
		UNCONNECTED_138, UNCONNECTED_139, UNCONNECTED_140, 
		UNCONNECTED_141, UNCONNECTED_142, UNCONNECTED_143, 
		UNCONNECTED_144, UNCONNECTED_145, UNCONNECTED_146, 
		UNCONNECTED_147}), .cr2(cr2), .icr2(icr2), .cr3({\cr3[31] , \cr3[30] 
		, \cr3[29] , \cr3[28] , \cr3[27] , \cr3[26] , \cr3[25] , \cr3[24] 
		, \cr3[23] , \cr3[22] , \cr3[21] , \cr3[20] , \cr3[19] , \cr3[18] 
		, \cr3[17] , \cr3[16] , \cr3[15] , \cr3[14] , \cr3[13] , \cr3[12] 
		, UNCONNECTED_148, UNCONNECTED_149, UNCONNECTED_150, 
		UNCONNECTED_151, UNCONNECTED_152, UNCONNECTED_153, 
		UNCONNECTED_154, UNCONNECTED_155, UNCONNECTED_156, 
		UNCONNECTED_157, UNCONNECTED_158, UNCONNECTED_159}), .cs({
		UNCONNECTED_160, UNCONNECTED_161, UNCONNECTED_162, 
		UNCONNECTED_163, UNCONNECTED_164, UNCONNECTED_165, 
		UNCONNECTED_166, UNCONNECTED_167, UNCONNECTED_168, 
		UNCONNECTED_169, UNCONNECTED_170, UNCONNECTED_171, 
		UNCONNECTED_172, UNCONNECTED_173, UNCONNECTED_174, 
		UNCONNECTED_175, UNCONNECTED_176, UNCONNECTED_177, 
		UNCONNECTED_178, UNCONNECTED_179, UNCONNECTED_180, 
		UNCONNECTED_181, UNCONNECTED_182, UNCONNECTED_183, 
		UNCONNECTED_184, UNCONNECTED_185, UNCONNECTED_186, 
		UNCONNECTED_187, UNCONNECTED_188, UNCONNECTED_189, \cs[1] , \cs[0] 
		}), .pg_fault(pg_fault), .ipg_fault(pc_pg_fault), .useq_ptr(useq_ptr
		), .valid_len(valid_len), .queue(queue), .pg_en(pg_en), .pc_out(pc_out
		), .pc_req(pc_req), .read_req(int_read_req), .write_req(int_write_req
		), .read_ack(int_read_ack), .write_ack(int_write_ack), .flush_Itlb
		(flush_Itlb), .flush_Dtlb(flush_Dtlb), .readio_req(readio_req), 
		.writeio_req(writeio_req), .readio_ack(readio_ack), .writeio_ack
		(writeio_ack), .write_data(iwrite_data), .writeio_data(writeio_data
		), .read_data(read_data_realign), .readio_data(readio_data), .write_sz
		(int_write_sz), .io_add({UNCONNECTED_190, UNCONNECTED_191, 
		UNCONNECTED_192, UNCONNECTED_193, UNCONNECTED_194, 
		UNCONNECTED_195, UNCONNECTED_196, UNCONNECTED_197, 
		UNCONNECTED_198, UNCONNECTED_199, UNCONNECTED_200, 
		UNCONNECTED_201, UNCONNECTED_202, UNCONNECTED_203, 
		UNCONNECTED_204, UNCONNECTED_205, io_add[15], io_add[14], io_add
		[13], io_add[12], io_add[11], io_add[10], io_add[9], io_add[8], io_add
		[7], io_add[6], io_add[5], io_add[4], io_add[3], io_add[2], io_add
		[1], io_add[0]}), .Daddr(int_Daddr), .pt_fault(pt_fault), .wr_fault
		(wr_fault));
	useq i_useq(.iaddr(int_code_addr), .idata(code_data), .code_req(int_code_req
		), .code_ack(int_code_ack), .clk(clk), .rstn(rstn), .useq_ptr(useq_ptr
		), .squeue(queue), .pc_in(pc_out), .pc_req(pc_req), .pg_fault(n_3135
		), .pc_pg_fault(pc_pg_fault), .valid_len(valid_len), .busy_ram(busy_ram
		));
endmodule
module v586(m00_AXI_RSTN, m00_AXI_CLK, m00_AXI_AWADDR, m00_AXI_AWVALID, m00_AXI_AWREADY
		, m00_AXI_AWBURST, m00_AXI_AWLEN, m00_AXI_AWSIZE, m00_AXI_ARADDR
		, m00_AXI_ARVALID, m00_AXI_ARREADY, m00_AXI_ARBURST, m00_AXI_ARLEN
		, m00_AXI_ARSIZE, m00_AXI_WDATA, m00_AXI_WVALID, m00_AXI_WREADY,
		 m00_AXI_WSTRB, m00_AXI_WLAST, m00_AXI_RDATA, m00_AXI_RVALID, m00_AXI_RREADY
		, m00_AXI_RLAST, m00_AXI_BVALID, m00_AXI_BREADY, m01_AXI_AWADDR,
		 m01_AXI_AWVALID, m01_AXI_AWREADY, m01_AXI_AWBURST, m01_AXI_AWLEN
		, m01_AXI_AWSIZE, m01_AXI_ARADDR, m01_AXI_ARVALID, m01_AXI_ARREADY
		, m01_AXI_ARBURST, m01_AXI_ARLEN, m01_AXI_ARSIZE, m01_AXI_WDATA,
		 m01_AXI_WVALID, m01_AXI_WREADY, m01_AXI_WSTRB, m01_AXI_WLAST, m01_AXI_RDATA
		, m01_AXI_RVALID, m01_AXI_RREADY, m01_AXI_RLAST, m01_AXI_BVALID,
		 m01_AXI_BREADY, int_pic, iack, ivect, debug);

	input m00_AXI_RSTN;
	input m00_AXI_CLK;
	output [31:0] m00_AXI_AWADDR;
	output m00_AXI_AWVALID;
	input m00_AXI_AWREADY;
	output [1:0] m00_AXI_AWBURST;
	output [7:0] m00_AXI_AWLEN;
	output [2:0] m00_AXI_AWSIZE;
	output [31:0] m00_AXI_ARADDR;
	output m00_AXI_ARVALID;
	input m00_AXI_ARREADY;
	output [1:0] m00_AXI_ARBURST;
	output [7:0] m00_AXI_ARLEN;
	output [2:0] m00_AXI_ARSIZE;
	output [31:0] m00_AXI_WDATA;
	output m00_AXI_WVALID;
	input m00_AXI_WREADY;
	output [3:0] m00_AXI_WSTRB;
	output m00_AXI_WLAST;
	input [31:0] m00_AXI_RDATA;
	input m00_AXI_RVALID;
	output m00_AXI_RREADY;
	input m00_AXI_RLAST;
	input m00_AXI_BVALID;
	output m00_AXI_BREADY;
	output [31:0] m01_AXI_AWADDR;
	output m01_AXI_AWVALID;
	input m01_AXI_AWREADY;
	output [1:0] m01_AXI_AWBURST;
	output [7:0] m01_AXI_AWLEN;
	output [2:0] m01_AXI_AWSIZE;
	output [31:0] m01_AXI_ARADDR;
	output m01_AXI_ARVALID;
	input m01_AXI_ARREADY;
	output [1:0] m01_AXI_ARBURST;
	output [7:0] m01_AXI_ARLEN;
	output [2:0] m01_AXI_ARSIZE;
	output [31:0] m01_AXI_WDATA;
	output m01_AXI_WVALID;
	input m01_AXI_WREADY;
	output [3:0] m01_AXI_WSTRB;
	output m01_AXI_WLAST;
	input [31:0] m01_AXI_RDATA;
	input m01_AXI_RVALID;
	output m01_AXI_RREADY;
	input m01_AXI_RLAST;
	input m01_AXI_BVALID;
	output m01_AXI_BREADY;
	input int_pic;
	output iack;
	input [7:0] ivect;
	output [4:0] debug;

	wire [3:0] write_msk;
	wire [31:0] writeio_data;
	wire [31:0] readio_data;
	wire [31:0] read_data;
	wire [31:0] write_data;
	wire [127:0] code_data;

	assign m00_AXI_BREADY = 1'b1;
	assign m01_AXI_AWBURST[1] = 1'b0;
	assign m01_AXI_AWBURST[0] = 1'b1;
	assign m01_AXI_AWLEN[7] = 1'b0;
	assign m01_AXI_AWLEN[6] = 1'b0;
	assign m01_AXI_AWLEN[5] = 1'b0;
	assign m01_AXI_AWLEN[4] = 1'b0;
	assign m01_AXI_AWLEN[3] = 1'b0;
	assign m01_AXI_AWLEN[2] = 1'b0;
	assign m01_AXI_AWLEN[1] = 1'b0;
	assign m01_AXI_AWLEN[0] = 1'b0;
	assign m01_AXI_AWSIZE[2] = 1'b0;
	assign m01_AXI_AWSIZE[1] = 1'b1;
	assign m01_AXI_AWSIZE[0] = 1'b0;
	assign m01_AXI_ARBURST[1] = 1'b0;
	assign m01_AXI_ARBURST[0] = 1'b1;
	assign m01_AXI_ARLEN[7] = 1'b0;
	assign m01_AXI_ARLEN[6] = 1'b0;
	assign m01_AXI_ARLEN[5] = 1'b0;
	assign m01_AXI_ARLEN[4] = 1'b0;
	assign m01_AXI_ARLEN[3] = 1'b0;
	assign m01_AXI_ARLEN[2] = 1'b0;
	assign m01_AXI_ARLEN[1] = 1'b0;
	assign m01_AXI_ARLEN[0] = 1'b0;
	assign m01_AXI_ARSIZE[2] = 1'b0;
	assign m01_AXI_ARSIZE[1] = 1'b1;
	assign m01_AXI_ARSIZE[0] = 1'b0;
	assign m01_AXI_WSTRB[3] = 1'b0;
	assign m01_AXI_WSTRB[2] = 1'b0;
	assign m01_AXI_WSTRB[1] = 1'b0;
	assign m01_AXI_WSTRB[0] = 1'b1;


	notech_inv i_15642(.A(n_61975), .Z(n_61977));
	notech_inv i_15641(.A(n_61975), .Z(n_61976));
	notech_inv i_15640(.A(m00_AXI_CLK), .Z(n_61975));
	biu32_axi ubiu(.rstn(m00_AXI_RSTN), .clk(n_61976), .write_req(write_req)
		, .write_ack(write_ack), .write_data(write_data), .write_msk(write_msk
		), .read_req(read_req), .read_ack(read_ack), .read_data(read_data
		), .Daddr({\Daddr[31] , \Daddr[30] , \Daddr[29] , \Daddr[28] , \Daddr[27] 
		, \Daddr[26] , \Daddr[25] , \Daddr[24] , \Daddr[23] , \Daddr[22] 
		, \Daddr[21] , \Daddr[20] , \Daddr[19] , \Daddr[18] , \Daddr[17] 
		, \Daddr[16] , \Daddr[15] , \Daddr[14] , \Daddr[13] , \Daddr[12] 
		, \Daddr[11] , \Daddr[10] , \Daddr[9] , \Daddr[8] , \Daddr[7] , \Daddr[6] 
		, \Daddr[5] , \Daddr[4] , \Daddr[3] , \Daddr[2] , 
		UNCONNECTED_000, UNCONNECTED_001}), .code_req(code_req), .code_ack
		(code_ack), .code_data(code_data), .code_addr({\code_addr[31] , \code_addr[30] 
		, \code_addr[29] , \code_addr[28] , \code_addr[27] , \code_addr[26] 
		, \code_addr[25] , \code_addr[24] , \code_addr[23] , \code_addr[22] 
		, \code_addr[21] , \code_addr[20] , \code_addr[19] , \code_addr[18] 
		, \code_addr[17] , \code_addr[16] , \code_addr[15] , \code_addr[14] 
		, \code_addr[13] , \code_addr[12] , \code_addr[11] , \code_addr[10] 
		, \code_addr[9] , \code_addr[8] , \code_addr[7] , \code_addr[6] 
		, \code_addr[5] , \code_addr[4] , \code_addr[3] , \code_addr[2] 
		, UNCONNECTED_002, UNCONNECTED_003}), .code_wreq(code_wreq), .code_wack
		(code_wack), .code_wdata({UNCONNECTED_004, UNCONNECTED_005, 
		UNCONNECTED_006, UNCONNECTED_007, UNCONNECTED_008, 
		UNCONNECTED_009, UNCONNECTED_010, UNCONNECTED_011, 
		UNCONNECTED_012, UNCONNECTED_013, UNCONNECTED_014, 
		UNCONNECTED_015, UNCONNECTED_016, UNCONNECTED_017, 
		UNCONNECTED_018, UNCONNECTED_019, UNCONNECTED_020, 
		UNCONNECTED_021, UNCONNECTED_022, UNCONNECTED_023, 
		UNCONNECTED_024, UNCONNECTED_025, UNCONNECTED_026, 
		UNCONNECTED_027, \code_wdata[7] , \code_wdata[6] , \code_wdata[5] 
		, \code_wdata[4] , \code_wdata[3] , \code_wdata[2] , \code_wdata[1] 
		, \code_wdata[0] }), .readio_req(readio_req), .writeio_req(writeio_req
		), .readio_ack(readio_ack), .writeio_ack(writeio_ack), .writeio_data
		(writeio_data), .readio_data(readio_data), .io_add({
		UNCONNECTED_028, UNCONNECTED_029, UNCONNECTED_030, 
		UNCONNECTED_031, UNCONNECTED_032, UNCONNECTED_033, 
		UNCONNECTED_034, UNCONNECTED_035, UNCONNECTED_036, 
		UNCONNECTED_037, UNCONNECTED_038, UNCONNECTED_039, 
		UNCONNECTED_040, UNCONNECTED_041, UNCONNECTED_042, 
		UNCONNECTED_043, \io_add[15] , \io_add[14] , \io_add[13] , \io_add[12] 
		, \io_add[11] , \io_add[10] , \io_add[9] , \io_add[8] , \io_add[7] 
		, \io_add[6] , \io_add[5] , \io_add[4] , \io_add[3] , \io_add[2] 
		, \io_add[1] , \io_add[0] }), .axi_AW(m00_AXI_AWADDR), .axi_AWVALID
		(m00_AXI_AWVALID), .axi_AWREADY(m00_AXI_AWREADY), .axi_AWBURST(m00_AXI_AWBURST
		), .axi_AWLEN(m00_AXI_AWLEN), .axi_AWSIZE(m00_AXI_AWSIZE), .axi_W
		(m00_AXI_WDATA), .axi_WVALID(m00_AXI_WVALID), .axi_WREADY(m00_AXI_WREADY
		), .axi_WSTRB(m00_AXI_WSTRB), .axi_WLAST(m00_AXI_WLAST), .axi_AR
		(m00_AXI_ARADDR), .axi_ARVALID(m00_AXI_ARVALID), .axi_ARREADY(m00_AXI_ARREADY
		), .axi_ARBURST(m00_AXI_ARBURST), .axi_ARLEN(m00_AXI_ARLEN), .axi_ARSIZE
		(m00_AXI_ARSIZE), .axi_R(m00_AXI_RDATA), .axi_RVALID(m00_AXI_RVALID
		), .axi_RREADY(m00_AXI_RREADY), .axi_RLAST(m00_AXI_RLAST), .axi_io_AW
		(m01_AXI_AWADDR), .axi_io_AWVALID(m01_AXI_AWVALID), .axi_io_AWREADY
		(m01_AXI_AWREADY), .axi_io_W(m01_AXI_WDATA), .axi_io_WVALID(m01_AXI_WVALID
		), .axi_io_WREADY(m01_AXI_WREADY), .axi_io_WLAST(m01_AXI_WLAST),
		 .axi_io_AR(m01_AXI_ARADDR), .axi_io_ARVALID(m01_AXI_ARVALID), .axi_io_ARREADY
		(m01_AXI_ARREADY), .axi_io_R(m01_AXI_RDATA), .axi_io_RVALID(m01_AXI_RVALID
		), .axi_io_RREADY(m01_AXI_RREADY), .busy(busy_ram));
	core ucore(.clk(n_61977), .rstn(m00_AXI_RSTN), .ivect(ivect), .int_main(int_pic
		), .iack(iack), .code_addr({\code_addr[31] , \code_addr[30] , \code_addr[29] 
		, \code_addr[28] , \code_addr[27] , \code_addr[26] , \code_addr[25] 
		, \code_addr[24] , \code_addr[23] , \code_addr[22] , \code_addr[21] 
		, \code_addr[20] , \code_addr[19] , \code_addr[18] , \code_addr[17] 
		, \code_addr[16] , \code_addr[15] , \code_addr[14] , \code_addr[13] 
		, \code_addr[12] , \code_addr[11] , \code_addr[10] , \code_addr[9] 
		, \code_addr[8] , \code_addr[7] , \code_addr[6] , \code_addr[5] 
		, \code_addr[4] , \code_addr[3] , \code_addr[2] , 
		UNCONNECTED_044, UNCONNECTED_045}), .code_data(code_data), .code_req
		(code_req), .code_ack(code_ack), .code_wreq(code_wreq), .code_wack
		(code_wack), .code_wdata({UNCONNECTED_046, UNCONNECTED_047, 
		UNCONNECTED_048, UNCONNECTED_049, UNCONNECTED_050, 
		UNCONNECTED_051, UNCONNECTED_052, UNCONNECTED_053, 
		UNCONNECTED_054, UNCONNECTED_055, UNCONNECTED_056, 
		UNCONNECTED_057, UNCONNECTED_058, UNCONNECTED_059, 
		UNCONNECTED_060, UNCONNECTED_061, UNCONNECTED_062, 
		UNCONNECTED_063, UNCONNECTED_064, UNCONNECTED_065, 
		UNCONNECTED_066, UNCONNECTED_067, UNCONNECTED_068, 
		UNCONNECTED_069, \code_wdata[7] , \code_wdata[6] , \code_wdata[5] 
		, \code_wdata[4] , \code_wdata[3] , \code_wdata[2] , \code_wdata[1] 
		, \code_wdata[0] }), .readio_data(readio_data), .io_add({
		UNCONNECTED_070, UNCONNECTED_071, UNCONNECTED_072, 
		UNCONNECTED_073, UNCONNECTED_074, UNCONNECTED_075, 
		UNCONNECTED_076, UNCONNECTED_077, UNCONNECTED_078, 
		UNCONNECTED_079, UNCONNECTED_080, UNCONNECTED_081, 
		UNCONNECTED_082, UNCONNECTED_083, UNCONNECTED_084, 
		UNCONNECTED_085, \io_add[15] , \io_add[14] , \io_add[13] , \io_add[12] 
		, \io_add[11] , \io_add[10] , \io_add[9] , \io_add[8] , \io_add[7] 
		, \io_add[6] , \io_add[5] , \io_add[4] , \io_add[3] , \io_add[2] 
		, \io_add[1] , \io_add[0] }), .writeio_data(writeio_data), .writeio_req
		(writeio_req), .readio_req(readio_req), .writeio_ack(writeio_ack
		), .readio_ack(readio_ack), .write_req(write_req), .write_ack(write_ack
		), .write_data(write_data), .write_msk(write_msk), .read_req(read_req
		), .read_ack(read_ack), .read_data(read_data), .Daddr({\Daddr[31] 
		, \Daddr[30] , \Daddr[29] , \Daddr[28] , \Daddr[27] , \Daddr[26] 
		, \Daddr[25] , \Daddr[24] , \Daddr[23] , \Daddr[22] , \Daddr[21] 
		, \Daddr[20] , \Daddr[19] , \Daddr[18] , \Daddr[17] , \Daddr[16] 
		, \Daddr[15] , \Daddr[14] , \Daddr[13] , \Daddr[12] , \Daddr[11] 
		, \Daddr[10] , \Daddr[9] , \Daddr[8] , \Daddr[7] , \Daddr[6] , \Daddr[5] 
		, \Daddr[4] , \Daddr[3] , \Daddr[2] , UNCONNECTED_086, 
		UNCONNECTED_087}), .busy_ram(busy_ram));
endmodule
